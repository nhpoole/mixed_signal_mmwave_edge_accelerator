magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect 8500 -31610 42469 5732
<< nwell >>
rect 15390 -1694 24486 2310
rect 25972 1912 31856 2230
rect 25972 -1694 32316 1912
<< pwell >>
rect 15400 4184 24476 4336
rect 15400 2636 15552 4184
rect 24324 2636 24476 4184
rect 15400 2484 24476 2636
rect 25982 4184 31478 4336
rect 25982 2556 26134 4184
rect 31326 2556 31478 4184
rect 25982 2404 31478 2556
<< psubdiff >>
rect 15426 4277 24450 4310
rect 15426 4243 15603 4277
rect 15637 4243 15671 4277
rect 15705 4243 15739 4277
rect 15773 4243 15807 4277
rect 15841 4243 15875 4277
rect 15909 4243 15943 4277
rect 15977 4243 16011 4277
rect 16045 4243 16079 4277
rect 16113 4243 16147 4277
rect 16181 4243 16215 4277
rect 16249 4243 16283 4277
rect 16317 4243 16351 4277
rect 16385 4243 16419 4277
rect 16453 4243 16487 4277
rect 16521 4243 16555 4277
rect 16589 4243 16623 4277
rect 16657 4243 16691 4277
rect 16725 4243 16759 4277
rect 16793 4243 16827 4277
rect 16861 4243 16895 4277
rect 16929 4243 16963 4277
rect 16997 4243 17031 4277
rect 17065 4243 17099 4277
rect 17133 4243 17167 4277
rect 17201 4243 17235 4277
rect 17269 4243 17303 4277
rect 17337 4243 17371 4277
rect 17405 4243 17439 4277
rect 17473 4243 17507 4277
rect 17541 4243 17575 4277
rect 17609 4243 17643 4277
rect 17677 4243 17711 4277
rect 17745 4243 17779 4277
rect 17813 4243 17847 4277
rect 17881 4243 17915 4277
rect 17949 4243 17983 4277
rect 18017 4243 18051 4277
rect 18085 4243 18119 4277
rect 18153 4243 18187 4277
rect 18221 4243 18255 4277
rect 18289 4243 18323 4277
rect 18357 4243 18391 4277
rect 18425 4243 18459 4277
rect 18493 4243 18527 4277
rect 18561 4243 18595 4277
rect 18629 4243 18663 4277
rect 18697 4243 18731 4277
rect 18765 4243 18799 4277
rect 18833 4243 18867 4277
rect 18901 4243 18935 4277
rect 18969 4243 19003 4277
rect 19037 4243 19071 4277
rect 19105 4243 19139 4277
rect 19173 4243 19207 4277
rect 19241 4243 19275 4277
rect 19309 4243 19343 4277
rect 19377 4243 19411 4277
rect 19445 4243 19479 4277
rect 19513 4243 19547 4277
rect 19581 4243 19615 4277
rect 19649 4243 19683 4277
rect 19717 4243 19751 4277
rect 19785 4243 19819 4277
rect 19853 4243 19887 4277
rect 19921 4243 19955 4277
rect 19989 4243 20023 4277
rect 20057 4243 20091 4277
rect 20125 4243 20159 4277
rect 20193 4243 20227 4277
rect 20261 4243 20295 4277
rect 20329 4243 20363 4277
rect 20397 4243 20431 4277
rect 20465 4243 20499 4277
rect 20533 4243 20567 4277
rect 20601 4243 20635 4277
rect 20669 4243 20703 4277
rect 20737 4243 20771 4277
rect 20805 4243 20839 4277
rect 20873 4243 20907 4277
rect 20941 4243 20975 4277
rect 21009 4243 21043 4277
rect 21077 4243 21111 4277
rect 21145 4243 21179 4277
rect 21213 4243 21247 4277
rect 21281 4243 21315 4277
rect 21349 4243 21383 4277
rect 21417 4243 21451 4277
rect 21485 4243 21519 4277
rect 21553 4243 21587 4277
rect 21621 4243 21655 4277
rect 21689 4243 21723 4277
rect 21757 4243 21791 4277
rect 21825 4243 21859 4277
rect 21893 4243 21927 4277
rect 21961 4243 21995 4277
rect 22029 4243 22063 4277
rect 22097 4243 22131 4277
rect 22165 4243 22199 4277
rect 22233 4243 22267 4277
rect 22301 4243 22335 4277
rect 22369 4243 22403 4277
rect 22437 4243 22471 4277
rect 22505 4243 22539 4277
rect 22573 4243 22607 4277
rect 22641 4243 22675 4277
rect 22709 4243 22743 4277
rect 22777 4243 22811 4277
rect 22845 4243 22879 4277
rect 22913 4243 22947 4277
rect 22981 4243 23015 4277
rect 23049 4243 23083 4277
rect 23117 4243 23151 4277
rect 23185 4243 23219 4277
rect 23253 4243 23287 4277
rect 23321 4243 23355 4277
rect 23389 4243 23423 4277
rect 23457 4243 23491 4277
rect 23525 4243 23559 4277
rect 23593 4243 23627 4277
rect 23661 4243 23695 4277
rect 23729 4243 23763 4277
rect 23797 4243 23831 4277
rect 23865 4243 23899 4277
rect 23933 4243 23967 4277
rect 24001 4243 24035 4277
rect 24069 4243 24103 4277
rect 24137 4243 24171 4277
rect 24205 4243 24239 4277
rect 24273 4243 24450 4277
rect 15426 4210 24450 4243
rect 15426 4141 15526 4210
rect 15426 4107 15459 4141
rect 15493 4107 15526 4141
rect 15426 4073 15526 4107
rect 15426 4039 15459 4073
rect 15493 4039 15526 4073
rect 15426 4005 15526 4039
rect 15426 3971 15459 4005
rect 15493 3971 15526 4005
rect 15426 3937 15526 3971
rect 15426 3903 15459 3937
rect 15493 3903 15526 3937
rect 15426 3869 15526 3903
rect 15426 3835 15459 3869
rect 15493 3835 15526 3869
rect 15426 3801 15526 3835
rect 15426 3767 15459 3801
rect 15493 3767 15526 3801
rect 15426 3733 15526 3767
rect 15426 3699 15459 3733
rect 15493 3699 15526 3733
rect 15426 3665 15526 3699
rect 15426 3631 15459 3665
rect 15493 3631 15526 3665
rect 15426 3597 15526 3631
rect 15426 3563 15459 3597
rect 15493 3563 15526 3597
rect 15426 3529 15526 3563
rect 15426 3495 15459 3529
rect 15493 3495 15526 3529
rect 15426 3461 15526 3495
rect 15426 3427 15459 3461
rect 15493 3427 15526 3461
rect 15426 3393 15526 3427
rect 15426 3359 15459 3393
rect 15493 3359 15526 3393
rect 15426 3325 15526 3359
rect 15426 3291 15459 3325
rect 15493 3291 15526 3325
rect 15426 3257 15526 3291
rect 15426 3223 15459 3257
rect 15493 3223 15526 3257
rect 15426 3189 15526 3223
rect 15426 3155 15459 3189
rect 15493 3155 15526 3189
rect 15426 3121 15526 3155
rect 15426 3087 15459 3121
rect 15493 3087 15526 3121
rect 15426 3053 15526 3087
rect 15426 3019 15459 3053
rect 15493 3019 15526 3053
rect 15426 2985 15526 3019
rect 15426 2951 15459 2985
rect 15493 2951 15526 2985
rect 15426 2917 15526 2951
rect 15426 2883 15459 2917
rect 15493 2883 15526 2917
rect 15426 2849 15526 2883
rect 15426 2815 15459 2849
rect 15493 2815 15526 2849
rect 15426 2781 15526 2815
rect 15426 2747 15459 2781
rect 15493 2747 15526 2781
rect 15426 2713 15526 2747
rect 15426 2679 15459 2713
rect 15493 2679 15526 2713
rect 15426 2610 15526 2679
rect 24350 4141 24450 4210
rect 24350 4107 24383 4141
rect 24417 4107 24450 4141
rect 24350 4073 24450 4107
rect 24350 4039 24383 4073
rect 24417 4039 24450 4073
rect 24350 4005 24450 4039
rect 24350 3971 24383 4005
rect 24417 3971 24450 4005
rect 24350 3937 24450 3971
rect 24350 3903 24383 3937
rect 24417 3903 24450 3937
rect 24350 3869 24450 3903
rect 24350 3835 24383 3869
rect 24417 3835 24450 3869
rect 24350 3801 24450 3835
rect 24350 3767 24383 3801
rect 24417 3767 24450 3801
rect 24350 3733 24450 3767
rect 24350 3699 24383 3733
rect 24417 3699 24450 3733
rect 24350 3665 24450 3699
rect 24350 3631 24383 3665
rect 24417 3631 24450 3665
rect 24350 3597 24450 3631
rect 24350 3563 24383 3597
rect 24417 3563 24450 3597
rect 24350 3529 24450 3563
rect 24350 3495 24383 3529
rect 24417 3495 24450 3529
rect 24350 3461 24450 3495
rect 24350 3427 24383 3461
rect 24417 3427 24450 3461
rect 24350 3393 24450 3427
rect 24350 3359 24383 3393
rect 24417 3359 24450 3393
rect 24350 3325 24450 3359
rect 24350 3291 24383 3325
rect 24417 3291 24450 3325
rect 24350 3257 24450 3291
rect 24350 3223 24383 3257
rect 24417 3223 24450 3257
rect 24350 3189 24450 3223
rect 24350 3155 24383 3189
rect 24417 3155 24450 3189
rect 24350 3121 24450 3155
rect 24350 3087 24383 3121
rect 24417 3087 24450 3121
rect 24350 3053 24450 3087
rect 24350 3019 24383 3053
rect 24417 3019 24450 3053
rect 24350 2985 24450 3019
rect 24350 2951 24383 2985
rect 24417 2951 24450 2985
rect 24350 2917 24450 2951
rect 24350 2883 24383 2917
rect 24417 2883 24450 2917
rect 24350 2849 24450 2883
rect 24350 2815 24383 2849
rect 24417 2815 24450 2849
rect 24350 2781 24450 2815
rect 24350 2747 24383 2781
rect 24417 2747 24450 2781
rect 24350 2713 24450 2747
rect 24350 2679 24383 2713
rect 24417 2679 24450 2713
rect 24350 2610 24450 2679
rect 15426 2577 24450 2610
rect 15426 2543 15603 2577
rect 15637 2543 15671 2577
rect 15705 2543 15739 2577
rect 15773 2543 15807 2577
rect 15841 2543 15875 2577
rect 15909 2543 15943 2577
rect 15977 2543 16011 2577
rect 16045 2543 16079 2577
rect 16113 2543 16147 2577
rect 16181 2543 16215 2577
rect 16249 2543 16283 2577
rect 16317 2543 16351 2577
rect 16385 2543 16419 2577
rect 16453 2543 16487 2577
rect 16521 2543 16555 2577
rect 16589 2543 16623 2577
rect 16657 2543 16691 2577
rect 16725 2543 16759 2577
rect 16793 2543 16827 2577
rect 16861 2543 16895 2577
rect 16929 2543 16963 2577
rect 16997 2543 17031 2577
rect 17065 2543 17099 2577
rect 17133 2543 17167 2577
rect 17201 2543 17235 2577
rect 17269 2543 17303 2577
rect 17337 2543 17371 2577
rect 17405 2543 17439 2577
rect 17473 2543 17507 2577
rect 17541 2543 17575 2577
rect 17609 2543 17643 2577
rect 17677 2543 17711 2577
rect 17745 2543 17779 2577
rect 17813 2543 17847 2577
rect 17881 2543 17915 2577
rect 17949 2543 17983 2577
rect 18017 2543 18051 2577
rect 18085 2543 18119 2577
rect 18153 2543 18187 2577
rect 18221 2543 18255 2577
rect 18289 2543 18323 2577
rect 18357 2543 18391 2577
rect 18425 2543 18459 2577
rect 18493 2543 18527 2577
rect 18561 2543 18595 2577
rect 18629 2543 18663 2577
rect 18697 2543 18731 2577
rect 18765 2543 18799 2577
rect 18833 2543 18867 2577
rect 18901 2543 18935 2577
rect 18969 2543 19003 2577
rect 19037 2543 19071 2577
rect 19105 2543 19139 2577
rect 19173 2543 19207 2577
rect 19241 2543 19275 2577
rect 19309 2543 19343 2577
rect 19377 2543 19411 2577
rect 19445 2543 19479 2577
rect 19513 2543 19547 2577
rect 19581 2543 19615 2577
rect 19649 2543 19683 2577
rect 19717 2543 19751 2577
rect 19785 2543 19819 2577
rect 19853 2543 19887 2577
rect 19921 2543 19955 2577
rect 19989 2543 20023 2577
rect 20057 2543 20091 2577
rect 20125 2543 20159 2577
rect 20193 2543 20227 2577
rect 20261 2543 20295 2577
rect 20329 2543 20363 2577
rect 20397 2543 20431 2577
rect 20465 2543 20499 2577
rect 20533 2543 20567 2577
rect 20601 2543 20635 2577
rect 20669 2543 20703 2577
rect 20737 2543 20771 2577
rect 20805 2543 20839 2577
rect 20873 2543 20907 2577
rect 20941 2543 20975 2577
rect 21009 2543 21043 2577
rect 21077 2543 21111 2577
rect 21145 2543 21179 2577
rect 21213 2543 21247 2577
rect 21281 2543 21315 2577
rect 21349 2543 21383 2577
rect 21417 2543 21451 2577
rect 21485 2543 21519 2577
rect 21553 2543 21587 2577
rect 21621 2543 21655 2577
rect 21689 2543 21723 2577
rect 21757 2543 21791 2577
rect 21825 2543 21859 2577
rect 21893 2543 21927 2577
rect 21961 2543 21995 2577
rect 22029 2543 22063 2577
rect 22097 2543 22131 2577
rect 22165 2543 22199 2577
rect 22233 2543 22267 2577
rect 22301 2543 22335 2577
rect 22369 2543 22403 2577
rect 22437 2543 22471 2577
rect 22505 2543 22539 2577
rect 22573 2543 22607 2577
rect 22641 2543 22675 2577
rect 22709 2543 22743 2577
rect 22777 2543 22811 2577
rect 22845 2543 22879 2577
rect 22913 2543 22947 2577
rect 22981 2543 23015 2577
rect 23049 2543 23083 2577
rect 23117 2543 23151 2577
rect 23185 2543 23219 2577
rect 23253 2543 23287 2577
rect 23321 2543 23355 2577
rect 23389 2543 23423 2577
rect 23457 2543 23491 2577
rect 23525 2543 23559 2577
rect 23593 2543 23627 2577
rect 23661 2543 23695 2577
rect 23729 2543 23763 2577
rect 23797 2543 23831 2577
rect 23865 2543 23899 2577
rect 23933 2543 23967 2577
rect 24001 2543 24035 2577
rect 24069 2543 24103 2577
rect 24137 2543 24171 2577
rect 24205 2543 24239 2577
rect 24273 2543 24450 2577
rect 15426 2510 24450 2543
rect 26008 4277 31452 4310
rect 26008 4243 26197 4277
rect 26231 4243 26265 4277
rect 26299 4243 26333 4277
rect 26367 4243 26401 4277
rect 26435 4243 26469 4277
rect 26503 4243 26537 4277
rect 26571 4243 26605 4277
rect 26639 4243 26673 4277
rect 26707 4243 26741 4277
rect 26775 4243 26809 4277
rect 26843 4243 26877 4277
rect 26911 4243 26945 4277
rect 26979 4243 27013 4277
rect 27047 4243 27081 4277
rect 27115 4243 27149 4277
rect 27183 4243 27217 4277
rect 27251 4243 27285 4277
rect 27319 4243 27353 4277
rect 27387 4243 27421 4277
rect 27455 4243 27489 4277
rect 27523 4243 27557 4277
rect 27591 4243 27625 4277
rect 27659 4243 27693 4277
rect 27727 4243 27761 4277
rect 27795 4243 27829 4277
rect 27863 4243 27897 4277
rect 27931 4243 27965 4277
rect 27999 4243 28033 4277
rect 28067 4243 28101 4277
rect 28135 4243 28169 4277
rect 28203 4243 28237 4277
rect 28271 4243 28305 4277
rect 28339 4243 28373 4277
rect 28407 4243 28441 4277
rect 28475 4243 28509 4277
rect 28543 4243 28577 4277
rect 28611 4243 28645 4277
rect 28679 4243 28713 4277
rect 28747 4243 28781 4277
rect 28815 4243 28849 4277
rect 28883 4243 28917 4277
rect 28951 4243 28985 4277
rect 29019 4243 29053 4277
rect 29087 4243 29121 4277
rect 29155 4243 29189 4277
rect 29223 4243 29257 4277
rect 29291 4243 29325 4277
rect 29359 4243 29393 4277
rect 29427 4243 29461 4277
rect 29495 4243 29529 4277
rect 29563 4243 29597 4277
rect 29631 4243 29665 4277
rect 29699 4243 29733 4277
rect 29767 4243 29801 4277
rect 29835 4243 29869 4277
rect 29903 4243 29937 4277
rect 29971 4243 30005 4277
rect 30039 4243 30073 4277
rect 30107 4243 30141 4277
rect 30175 4243 30209 4277
rect 30243 4243 30277 4277
rect 30311 4243 30345 4277
rect 30379 4243 30413 4277
rect 30447 4243 30481 4277
rect 30515 4243 30549 4277
rect 30583 4243 30617 4277
rect 30651 4243 30685 4277
rect 30719 4243 30753 4277
rect 30787 4243 30821 4277
rect 30855 4243 30889 4277
rect 30923 4243 30957 4277
rect 30991 4243 31025 4277
rect 31059 4243 31093 4277
rect 31127 4243 31161 4277
rect 31195 4243 31229 4277
rect 31263 4243 31452 4277
rect 26008 4210 31452 4243
rect 26008 4135 26108 4210
rect 26008 4101 26041 4135
rect 26075 4101 26108 4135
rect 26008 4067 26108 4101
rect 26008 4033 26041 4067
rect 26075 4033 26108 4067
rect 26008 3999 26108 4033
rect 26008 3965 26041 3999
rect 26075 3965 26108 3999
rect 26008 3931 26108 3965
rect 26008 3897 26041 3931
rect 26075 3897 26108 3931
rect 26008 3863 26108 3897
rect 26008 3829 26041 3863
rect 26075 3829 26108 3863
rect 26008 3795 26108 3829
rect 26008 3761 26041 3795
rect 26075 3761 26108 3795
rect 26008 3727 26108 3761
rect 26008 3693 26041 3727
rect 26075 3693 26108 3727
rect 26008 3659 26108 3693
rect 26008 3625 26041 3659
rect 26075 3625 26108 3659
rect 26008 3591 26108 3625
rect 26008 3557 26041 3591
rect 26075 3557 26108 3591
rect 26008 3523 26108 3557
rect 26008 3489 26041 3523
rect 26075 3489 26108 3523
rect 26008 3455 26108 3489
rect 26008 3421 26041 3455
rect 26075 3421 26108 3455
rect 26008 3387 26108 3421
rect 26008 3353 26041 3387
rect 26075 3353 26108 3387
rect 26008 3319 26108 3353
rect 26008 3285 26041 3319
rect 26075 3285 26108 3319
rect 26008 3251 26108 3285
rect 26008 3217 26041 3251
rect 26075 3217 26108 3251
rect 26008 3183 26108 3217
rect 26008 3149 26041 3183
rect 26075 3149 26108 3183
rect 26008 3115 26108 3149
rect 26008 3081 26041 3115
rect 26075 3081 26108 3115
rect 26008 3047 26108 3081
rect 26008 3013 26041 3047
rect 26075 3013 26108 3047
rect 26008 2979 26108 3013
rect 26008 2945 26041 2979
rect 26075 2945 26108 2979
rect 26008 2911 26108 2945
rect 26008 2877 26041 2911
rect 26075 2877 26108 2911
rect 26008 2843 26108 2877
rect 26008 2809 26041 2843
rect 26075 2809 26108 2843
rect 26008 2775 26108 2809
rect 26008 2741 26041 2775
rect 26075 2741 26108 2775
rect 26008 2707 26108 2741
rect 26008 2673 26041 2707
rect 26075 2673 26108 2707
rect 26008 2639 26108 2673
rect 26008 2605 26041 2639
rect 26075 2605 26108 2639
rect 26008 2530 26108 2605
rect 31352 4135 31452 4210
rect 31352 4101 31385 4135
rect 31419 4101 31452 4135
rect 31352 4067 31452 4101
rect 31352 4033 31385 4067
rect 31419 4033 31452 4067
rect 31352 3999 31452 4033
rect 31352 3965 31385 3999
rect 31419 3965 31452 3999
rect 31352 3931 31452 3965
rect 31352 3897 31385 3931
rect 31419 3897 31452 3931
rect 31352 3863 31452 3897
rect 31352 3829 31385 3863
rect 31419 3829 31452 3863
rect 31352 3795 31452 3829
rect 31352 3761 31385 3795
rect 31419 3761 31452 3795
rect 31352 3727 31452 3761
rect 31352 3693 31385 3727
rect 31419 3693 31452 3727
rect 31352 3659 31452 3693
rect 31352 3625 31385 3659
rect 31419 3625 31452 3659
rect 31352 3591 31452 3625
rect 31352 3557 31385 3591
rect 31419 3557 31452 3591
rect 31352 3523 31452 3557
rect 31352 3489 31385 3523
rect 31419 3489 31452 3523
rect 31352 3455 31452 3489
rect 31352 3421 31385 3455
rect 31419 3421 31452 3455
rect 31352 3387 31452 3421
rect 31352 3353 31385 3387
rect 31419 3353 31452 3387
rect 31352 3319 31452 3353
rect 31352 3285 31385 3319
rect 31419 3285 31452 3319
rect 31352 3251 31452 3285
rect 31352 3217 31385 3251
rect 31419 3217 31452 3251
rect 31352 3183 31452 3217
rect 31352 3149 31385 3183
rect 31419 3149 31452 3183
rect 31352 3115 31452 3149
rect 31352 3081 31385 3115
rect 31419 3081 31452 3115
rect 31352 3047 31452 3081
rect 31352 3013 31385 3047
rect 31419 3013 31452 3047
rect 31352 2979 31452 3013
rect 31352 2945 31385 2979
rect 31419 2945 31452 2979
rect 31352 2911 31452 2945
rect 31352 2877 31385 2911
rect 31419 2877 31452 2911
rect 31352 2843 31452 2877
rect 31352 2809 31385 2843
rect 31419 2809 31452 2843
rect 31352 2775 31452 2809
rect 31352 2741 31385 2775
rect 31419 2741 31452 2775
rect 31352 2707 31452 2741
rect 31352 2673 31385 2707
rect 31419 2673 31452 2707
rect 31352 2639 31452 2673
rect 31352 2605 31385 2639
rect 31419 2605 31452 2639
rect 31352 2530 31452 2605
rect 26008 2497 31452 2530
rect 26008 2463 26197 2497
rect 26231 2463 26265 2497
rect 26299 2463 26333 2497
rect 26367 2463 26401 2497
rect 26435 2463 26469 2497
rect 26503 2463 26537 2497
rect 26571 2463 26605 2497
rect 26639 2463 26673 2497
rect 26707 2463 26741 2497
rect 26775 2463 26809 2497
rect 26843 2463 26877 2497
rect 26911 2463 26945 2497
rect 26979 2463 27013 2497
rect 27047 2463 27081 2497
rect 27115 2463 27149 2497
rect 27183 2463 27217 2497
rect 27251 2463 27285 2497
rect 27319 2463 27353 2497
rect 27387 2463 27421 2497
rect 27455 2463 27489 2497
rect 27523 2463 27557 2497
rect 27591 2463 27625 2497
rect 27659 2463 27693 2497
rect 27727 2463 27761 2497
rect 27795 2463 27829 2497
rect 27863 2463 27897 2497
rect 27931 2463 27965 2497
rect 27999 2463 28033 2497
rect 28067 2463 28101 2497
rect 28135 2463 28169 2497
rect 28203 2463 28237 2497
rect 28271 2463 28305 2497
rect 28339 2463 28373 2497
rect 28407 2463 28441 2497
rect 28475 2463 28509 2497
rect 28543 2463 28577 2497
rect 28611 2463 28645 2497
rect 28679 2463 28713 2497
rect 28747 2463 28781 2497
rect 28815 2463 28849 2497
rect 28883 2463 28917 2497
rect 28951 2463 28985 2497
rect 29019 2463 29053 2497
rect 29087 2463 29121 2497
rect 29155 2463 29189 2497
rect 29223 2463 29257 2497
rect 29291 2463 29325 2497
rect 29359 2463 29393 2497
rect 29427 2463 29461 2497
rect 29495 2463 29529 2497
rect 29563 2463 29597 2497
rect 29631 2463 29665 2497
rect 29699 2463 29733 2497
rect 29767 2463 29801 2497
rect 29835 2463 29869 2497
rect 29903 2463 29937 2497
rect 29971 2463 30005 2497
rect 30039 2463 30073 2497
rect 30107 2463 30141 2497
rect 30175 2463 30209 2497
rect 30243 2463 30277 2497
rect 30311 2463 30345 2497
rect 30379 2463 30413 2497
rect 30447 2463 30481 2497
rect 30515 2463 30549 2497
rect 30583 2463 30617 2497
rect 30651 2463 30685 2497
rect 30719 2463 30753 2497
rect 30787 2463 30821 2497
rect 30855 2463 30889 2497
rect 30923 2463 30957 2497
rect 30991 2463 31025 2497
rect 31059 2463 31093 2497
rect 31127 2463 31161 2497
rect 31195 2463 31229 2497
rect 31263 2463 31452 2497
rect 26008 2430 31452 2463
<< nsubdiff >>
rect 15426 2241 24450 2274
rect 15426 2207 15603 2241
rect 15637 2207 15671 2241
rect 15705 2207 15739 2241
rect 15773 2207 15807 2241
rect 15841 2207 15875 2241
rect 15909 2207 15943 2241
rect 15977 2207 16011 2241
rect 16045 2207 16079 2241
rect 16113 2207 16147 2241
rect 16181 2207 16215 2241
rect 16249 2207 16283 2241
rect 16317 2207 16351 2241
rect 16385 2207 16419 2241
rect 16453 2207 16487 2241
rect 16521 2207 16555 2241
rect 16589 2207 16623 2241
rect 16657 2207 16691 2241
rect 16725 2207 16759 2241
rect 16793 2207 16827 2241
rect 16861 2207 16895 2241
rect 16929 2207 16963 2241
rect 16997 2207 17031 2241
rect 17065 2207 17099 2241
rect 17133 2207 17167 2241
rect 17201 2207 17235 2241
rect 17269 2207 17303 2241
rect 17337 2207 17371 2241
rect 17405 2207 17439 2241
rect 17473 2207 17507 2241
rect 17541 2207 17575 2241
rect 17609 2207 17643 2241
rect 17677 2207 17711 2241
rect 17745 2207 17779 2241
rect 17813 2207 17847 2241
rect 17881 2207 17915 2241
rect 17949 2207 17983 2241
rect 18017 2207 18051 2241
rect 18085 2207 18119 2241
rect 18153 2207 18187 2241
rect 18221 2207 18255 2241
rect 18289 2207 18323 2241
rect 18357 2207 18391 2241
rect 18425 2207 18459 2241
rect 18493 2207 18527 2241
rect 18561 2207 18595 2241
rect 18629 2207 18663 2241
rect 18697 2207 18731 2241
rect 18765 2207 18799 2241
rect 18833 2207 18867 2241
rect 18901 2207 18935 2241
rect 18969 2207 19003 2241
rect 19037 2207 19071 2241
rect 19105 2207 19139 2241
rect 19173 2207 19207 2241
rect 19241 2207 19275 2241
rect 19309 2207 19343 2241
rect 19377 2207 19411 2241
rect 19445 2207 19479 2241
rect 19513 2207 19547 2241
rect 19581 2207 19615 2241
rect 19649 2207 19683 2241
rect 19717 2207 19751 2241
rect 19785 2207 19819 2241
rect 19853 2207 19887 2241
rect 19921 2207 19955 2241
rect 19989 2207 20023 2241
rect 20057 2207 20091 2241
rect 20125 2207 20159 2241
rect 20193 2207 20227 2241
rect 20261 2207 20295 2241
rect 20329 2207 20363 2241
rect 20397 2207 20431 2241
rect 20465 2207 20499 2241
rect 20533 2207 20567 2241
rect 20601 2207 20635 2241
rect 20669 2207 20703 2241
rect 20737 2207 20771 2241
rect 20805 2207 20839 2241
rect 20873 2207 20907 2241
rect 20941 2207 20975 2241
rect 21009 2207 21043 2241
rect 21077 2207 21111 2241
rect 21145 2207 21179 2241
rect 21213 2207 21247 2241
rect 21281 2207 21315 2241
rect 21349 2207 21383 2241
rect 21417 2207 21451 2241
rect 21485 2207 21519 2241
rect 21553 2207 21587 2241
rect 21621 2207 21655 2241
rect 21689 2207 21723 2241
rect 21757 2207 21791 2241
rect 21825 2207 21859 2241
rect 21893 2207 21927 2241
rect 21961 2207 21995 2241
rect 22029 2207 22063 2241
rect 22097 2207 22131 2241
rect 22165 2207 22199 2241
rect 22233 2207 22267 2241
rect 22301 2207 22335 2241
rect 22369 2207 22403 2241
rect 22437 2207 22471 2241
rect 22505 2207 22539 2241
rect 22573 2207 22607 2241
rect 22641 2207 22675 2241
rect 22709 2207 22743 2241
rect 22777 2207 22811 2241
rect 22845 2207 22879 2241
rect 22913 2207 22947 2241
rect 22981 2207 23015 2241
rect 23049 2207 23083 2241
rect 23117 2207 23151 2241
rect 23185 2207 23219 2241
rect 23253 2207 23287 2241
rect 23321 2207 23355 2241
rect 23389 2207 23423 2241
rect 23457 2207 23491 2241
rect 23525 2207 23559 2241
rect 23593 2207 23627 2241
rect 23661 2207 23695 2241
rect 23729 2207 23763 2241
rect 23797 2207 23831 2241
rect 23865 2207 23899 2241
rect 23933 2207 23967 2241
rect 24001 2207 24035 2241
rect 24069 2207 24103 2241
rect 24137 2207 24171 2241
rect 24205 2207 24239 2241
rect 24273 2207 24450 2241
rect 15426 2174 24450 2207
rect 15426 2093 15526 2174
rect 15426 2059 15459 2093
rect 15493 2059 15526 2093
rect 15426 2025 15526 2059
rect 15426 1991 15459 2025
rect 15493 1991 15526 2025
rect 15426 1957 15526 1991
rect 15426 1923 15459 1957
rect 15493 1923 15526 1957
rect 15426 1889 15526 1923
rect 15426 1855 15459 1889
rect 15493 1855 15526 1889
rect 15426 1821 15526 1855
rect 15426 1787 15459 1821
rect 15493 1787 15526 1821
rect 15426 1753 15526 1787
rect 15426 1719 15459 1753
rect 15493 1719 15526 1753
rect 15426 1685 15526 1719
rect 15426 1651 15459 1685
rect 15493 1651 15526 1685
rect 15426 1617 15526 1651
rect 15426 1583 15459 1617
rect 15493 1583 15526 1617
rect 15426 1549 15526 1583
rect 15426 1515 15459 1549
rect 15493 1515 15526 1549
rect 15426 1481 15526 1515
rect 15426 1447 15459 1481
rect 15493 1447 15526 1481
rect 15426 1413 15526 1447
rect 15426 1379 15459 1413
rect 15493 1379 15526 1413
rect 15426 1345 15526 1379
rect 15426 1311 15459 1345
rect 15493 1311 15526 1345
rect 15426 1277 15526 1311
rect 15426 1243 15459 1277
rect 15493 1243 15526 1277
rect 15426 1209 15526 1243
rect 15426 1175 15459 1209
rect 15493 1175 15526 1209
rect 15426 1141 15526 1175
rect 15426 1107 15459 1141
rect 15493 1107 15526 1141
rect 15426 1073 15526 1107
rect 15426 1039 15459 1073
rect 15493 1039 15526 1073
rect 15426 1005 15526 1039
rect 15426 971 15459 1005
rect 15493 971 15526 1005
rect 15426 937 15526 971
rect 15426 903 15459 937
rect 15493 903 15526 937
rect 15426 869 15526 903
rect 15426 835 15459 869
rect 15493 835 15526 869
rect 15426 801 15526 835
rect 15426 767 15459 801
rect 15493 767 15526 801
rect 15426 733 15526 767
rect 15426 699 15459 733
rect 15493 699 15526 733
rect 15426 665 15526 699
rect 15426 631 15459 665
rect 15493 631 15526 665
rect 15426 597 15526 631
rect 15426 563 15459 597
rect 15493 563 15526 597
rect 15426 529 15526 563
rect 15426 495 15459 529
rect 15493 495 15526 529
rect 15426 461 15526 495
rect 15426 427 15459 461
rect 15493 427 15526 461
rect 15426 393 15526 427
rect 15426 359 15459 393
rect 15493 359 15526 393
rect 15426 325 15526 359
rect 15426 291 15459 325
rect 15493 291 15526 325
rect 15426 257 15526 291
rect 15426 223 15459 257
rect 15493 223 15526 257
rect 15426 189 15526 223
rect 15426 155 15459 189
rect 15493 155 15526 189
rect 15426 121 15526 155
rect 15426 87 15459 121
rect 15493 87 15526 121
rect 15426 53 15526 87
rect 15426 19 15459 53
rect 15493 19 15526 53
rect 15426 -15 15526 19
rect 15426 -49 15459 -15
rect 15493 -49 15526 -15
rect 15426 -83 15526 -49
rect 15426 -117 15459 -83
rect 15493 -117 15526 -83
rect 15426 -151 15526 -117
rect 15426 -185 15459 -151
rect 15493 -185 15526 -151
rect 15426 -219 15526 -185
rect 15426 -253 15459 -219
rect 15493 -253 15526 -219
rect 15426 -287 15526 -253
rect 15426 -321 15459 -287
rect 15493 -321 15526 -287
rect 15426 -355 15526 -321
rect 15426 -389 15459 -355
rect 15493 -389 15526 -355
rect 15426 -423 15526 -389
rect 15426 -457 15459 -423
rect 15493 -457 15526 -423
rect 15426 -491 15526 -457
rect 15426 -525 15459 -491
rect 15493 -525 15526 -491
rect 15426 -559 15526 -525
rect 15426 -593 15459 -559
rect 15493 -593 15526 -559
rect 15426 -627 15526 -593
rect 15426 -661 15459 -627
rect 15493 -661 15526 -627
rect 15426 -695 15526 -661
rect 15426 -729 15459 -695
rect 15493 -729 15526 -695
rect 15426 -763 15526 -729
rect 15426 -797 15459 -763
rect 15493 -797 15526 -763
rect 15426 -831 15526 -797
rect 15426 -865 15459 -831
rect 15493 -865 15526 -831
rect 15426 -899 15526 -865
rect 15426 -933 15459 -899
rect 15493 -933 15526 -899
rect 15426 -967 15526 -933
rect 15426 -1001 15459 -967
rect 15493 -1001 15526 -967
rect 15426 -1035 15526 -1001
rect 15426 -1069 15459 -1035
rect 15493 -1069 15526 -1035
rect 15426 -1103 15526 -1069
rect 15426 -1137 15459 -1103
rect 15493 -1137 15526 -1103
rect 15426 -1171 15526 -1137
rect 15426 -1205 15459 -1171
rect 15493 -1205 15526 -1171
rect 15426 -1239 15526 -1205
rect 15426 -1273 15459 -1239
rect 15493 -1273 15526 -1239
rect 15426 -1307 15526 -1273
rect 15426 -1341 15459 -1307
rect 15493 -1341 15526 -1307
rect 15426 -1375 15526 -1341
rect 15426 -1409 15459 -1375
rect 15493 -1409 15526 -1375
rect 15426 -1443 15526 -1409
rect 15426 -1477 15459 -1443
rect 15493 -1477 15526 -1443
rect 15426 -1558 15526 -1477
rect 24350 2093 24450 2174
rect 24350 2059 24383 2093
rect 24417 2059 24450 2093
rect 24350 2025 24450 2059
rect 24350 1991 24383 2025
rect 24417 1991 24450 2025
rect 24350 1957 24450 1991
rect 24350 1923 24383 1957
rect 24417 1923 24450 1957
rect 24350 1889 24450 1923
rect 24350 1855 24383 1889
rect 24417 1855 24450 1889
rect 24350 1821 24450 1855
rect 24350 1787 24383 1821
rect 24417 1787 24450 1821
rect 24350 1753 24450 1787
rect 24350 1719 24383 1753
rect 24417 1719 24450 1753
rect 24350 1685 24450 1719
rect 24350 1651 24383 1685
rect 24417 1651 24450 1685
rect 24350 1617 24450 1651
rect 24350 1583 24383 1617
rect 24417 1583 24450 1617
rect 24350 1549 24450 1583
rect 24350 1515 24383 1549
rect 24417 1515 24450 1549
rect 24350 1481 24450 1515
rect 24350 1447 24383 1481
rect 24417 1447 24450 1481
rect 24350 1413 24450 1447
rect 24350 1379 24383 1413
rect 24417 1379 24450 1413
rect 24350 1345 24450 1379
rect 24350 1311 24383 1345
rect 24417 1311 24450 1345
rect 24350 1277 24450 1311
rect 24350 1243 24383 1277
rect 24417 1243 24450 1277
rect 24350 1209 24450 1243
rect 24350 1175 24383 1209
rect 24417 1175 24450 1209
rect 24350 1141 24450 1175
rect 24350 1107 24383 1141
rect 24417 1107 24450 1141
rect 24350 1073 24450 1107
rect 24350 1039 24383 1073
rect 24417 1039 24450 1073
rect 24350 1005 24450 1039
rect 24350 971 24383 1005
rect 24417 971 24450 1005
rect 24350 937 24450 971
rect 24350 903 24383 937
rect 24417 903 24450 937
rect 24350 869 24450 903
rect 24350 835 24383 869
rect 24417 835 24450 869
rect 24350 801 24450 835
rect 24350 767 24383 801
rect 24417 767 24450 801
rect 24350 733 24450 767
rect 24350 699 24383 733
rect 24417 699 24450 733
rect 24350 665 24450 699
rect 24350 631 24383 665
rect 24417 631 24450 665
rect 24350 597 24450 631
rect 24350 563 24383 597
rect 24417 563 24450 597
rect 24350 529 24450 563
rect 24350 495 24383 529
rect 24417 495 24450 529
rect 24350 461 24450 495
rect 24350 427 24383 461
rect 24417 427 24450 461
rect 24350 393 24450 427
rect 24350 359 24383 393
rect 24417 359 24450 393
rect 24350 325 24450 359
rect 24350 291 24383 325
rect 24417 291 24450 325
rect 24350 257 24450 291
rect 24350 223 24383 257
rect 24417 223 24450 257
rect 24350 189 24450 223
rect 24350 155 24383 189
rect 24417 155 24450 189
rect 24350 121 24450 155
rect 24350 87 24383 121
rect 24417 87 24450 121
rect 24350 53 24450 87
rect 24350 19 24383 53
rect 24417 19 24450 53
rect 24350 -15 24450 19
rect 24350 -49 24383 -15
rect 24417 -49 24450 -15
rect 24350 -83 24450 -49
rect 24350 -117 24383 -83
rect 24417 -117 24450 -83
rect 24350 -151 24450 -117
rect 24350 -185 24383 -151
rect 24417 -185 24450 -151
rect 24350 -219 24450 -185
rect 24350 -253 24383 -219
rect 24417 -253 24450 -219
rect 24350 -287 24450 -253
rect 24350 -321 24383 -287
rect 24417 -321 24450 -287
rect 24350 -355 24450 -321
rect 24350 -389 24383 -355
rect 24417 -389 24450 -355
rect 24350 -423 24450 -389
rect 24350 -457 24383 -423
rect 24417 -457 24450 -423
rect 24350 -491 24450 -457
rect 24350 -525 24383 -491
rect 24417 -525 24450 -491
rect 24350 -559 24450 -525
rect 24350 -593 24383 -559
rect 24417 -593 24450 -559
rect 24350 -627 24450 -593
rect 24350 -661 24383 -627
rect 24417 -661 24450 -627
rect 24350 -695 24450 -661
rect 24350 -729 24383 -695
rect 24417 -729 24450 -695
rect 24350 -763 24450 -729
rect 24350 -797 24383 -763
rect 24417 -797 24450 -763
rect 24350 -831 24450 -797
rect 24350 -865 24383 -831
rect 24417 -865 24450 -831
rect 24350 -899 24450 -865
rect 24350 -933 24383 -899
rect 24417 -933 24450 -899
rect 24350 -967 24450 -933
rect 24350 -1001 24383 -967
rect 24417 -1001 24450 -967
rect 24350 -1035 24450 -1001
rect 24350 -1069 24383 -1035
rect 24417 -1069 24450 -1035
rect 24350 -1103 24450 -1069
rect 24350 -1137 24383 -1103
rect 24417 -1137 24450 -1103
rect 24350 -1171 24450 -1137
rect 24350 -1205 24383 -1171
rect 24417 -1205 24450 -1171
rect 24350 -1239 24450 -1205
rect 24350 -1273 24383 -1239
rect 24417 -1273 24450 -1239
rect 24350 -1307 24450 -1273
rect 24350 -1341 24383 -1307
rect 24417 -1341 24450 -1307
rect 24350 -1375 24450 -1341
rect 24350 -1409 24383 -1375
rect 24417 -1409 24450 -1375
rect 24350 -1443 24450 -1409
rect 24350 -1477 24383 -1443
rect 24417 -1477 24450 -1443
rect 24350 -1558 24450 -1477
rect 15426 -1591 24450 -1558
rect 15426 -1625 15603 -1591
rect 15637 -1625 15671 -1591
rect 15705 -1625 15739 -1591
rect 15773 -1625 15807 -1591
rect 15841 -1625 15875 -1591
rect 15909 -1625 15943 -1591
rect 15977 -1625 16011 -1591
rect 16045 -1625 16079 -1591
rect 16113 -1625 16147 -1591
rect 16181 -1625 16215 -1591
rect 16249 -1625 16283 -1591
rect 16317 -1625 16351 -1591
rect 16385 -1625 16419 -1591
rect 16453 -1625 16487 -1591
rect 16521 -1625 16555 -1591
rect 16589 -1625 16623 -1591
rect 16657 -1625 16691 -1591
rect 16725 -1625 16759 -1591
rect 16793 -1625 16827 -1591
rect 16861 -1625 16895 -1591
rect 16929 -1625 16963 -1591
rect 16997 -1625 17031 -1591
rect 17065 -1625 17099 -1591
rect 17133 -1625 17167 -1591
rect 17201 -1625 17235 -1591
rect 17269 -1625 17303 -1591
rect 17337 -1625 17371 -1591
rect 17405 -1625 17439 -1591
rect 17473 -1625 17507 -1591
rect 17541 -1625 17575 -1591
rect 17609 -1625 17643 -1591
rect 17677 -1625 17711 -1591
rect 17745 -1625 17779 -1591
rect 17813 -1625 17847 -1591
rect 17881 -1625 17915 -1591
rect 17949 -1625 17983 -1591
rect 18017 -1625 18051 -1591
rect 18085 -1625 18119 -1591
rect 18153 -1625 18187 -1591
rect 18221 -1625 18255 -1591
rect 18289 -1625 18323 -1591
rect 18357 -1625 18391 -1591
rect 18425 -1625 18459 -1591
rect 18493 -1625 18527 -1591
rect 18561 -1625 18595 -1591
rect 18629 -1625 18663 -1591
rect 18697 -1625 18731 -1591
rect 18765 -1625 18799 -1591
rect 18833 -1625 18867 -1591
rect 18901 -1625 18935 -1591
rect 18969 -1625 19003 -1591
rect 19037 -1625 19071 -1591
rect 19105 -1625 19139 -1591
rect 19173 -1625 19207 -1591
rect 19241 -1625 19275 -1591
rect 19309 -1625 19343 -1591
rect 19377 -1625 19411 -1591
rect 19445 -1625 19479 -1591
rect 19513 -1625 19547 -1591
rect 19581 -1625 19615 -1591
rect 19649 -1625 19683 -1591
rect 19717 -1625 19751 -1591
rect 19785 -1625 19819 -1591
rect 19853 -1625 19887 -1591
rect 19921 -1625 19955 -1591
rect 19989 -1625 20023 -1591
rect 20057 -1625 20091 -1591
rect 20125 -1625 20159 -1591
rect 20193 -1625 20227 -1591
rect 20261 -1625 20295 -1591
rect 20329 -1625 20363 -1591
rect 20397 -1625 20431 -1591
rect 20465 -1625 20499 -1591
rect 20533 -1625 20567 -1591
rect 20601 -1625 20635 -1591
rect 20669 -1625 20703 -1591
rect 20737 -1625 20771 -1591
rect 20805 -1625 20839 -1591
rect 20873 -1625 20907 -1591
rect 20941 -1625 20975 -1591
rect 21009 -1625 21043 -1591
rect 21077 -1625 21111 -1591
rect 21145 -1625 21179 -1591
rect 21213 -1625 21247 -1591
rect 21281 -1625 21315 -1591
rect 21349 -1625 21383 -1591
rect 21417 -1625 21451 -1591
rect 21485 -1625 21519 -1591
rect 21553 -1625 21587 -1591
rect 21621 -1625 21655 -1591
rect 21689 -1625 21723 -1591
rect 21757 -1625 21791 -1591
rect 21825 -1625 21859 -1591
rect 21893 -1625 21927 -1591
rect 21961 -1625 21995 -1591
rect 22029 -1625 22063 -1591
rect 22097 -1625 22131 -1591
rect 22165 -1625 22199 -1591
rect 22233 -1625 22267 -1591
rect 22301 -1625 22335 -1591
rect 22369 -1625 22403 -1591
rect 22437 -1625 22471 -1591
rect 22505 -1625 22539 -1591
rect 22573 -1625 22607 -1591
rect 22641 -1625 22675 -1591
rect 22709 -1625 22743 -1591
rect 22777 -1625 22811 -1591
rect 22845 -1625 22879 -1591
rect 22913 -1625 22947 -1591
rect 22981 -1625 23015 -1591
rect 23049 -1625 23083 -1591
rect 23117 -1625 23151 -1591
rect 23185 -1625 23219 -1591
rect 23253 -1625 23287 -1591
rect 23321 -1625 23355 -1591
rect 23389 -1625 23423 -1591
rect 23457 -1625 23491 -1591
rect 23525 -1625 23559 -1591
rect 23593 -1625 23627 -1591
rect 23661 -1625 23695 -1591
rect 23729 -1625 23763 -1591
rect 23797 -1625 23831 -1591
rect 23865 -1625 23899 -1591
rect 23933 -1625 23967 -1591
rect 24001 -1625 24035 -1591
rect 24069 -1625 24103 -1591
rect 24137 -1625 24171 -1591
rect 24205 -1625 24239 -1591
rect 24273 -1625 24450 -1591
rect 15426 -1658 24450 -1625
rect 26008 2161 31452 2194
rect 26008 2127 26197 2161
rect 26231 2127 26265 2161
rect 26299 2127 26333 2161
rect 26367 2127 26401 2161
rect 26435 2127 26469 2161
rect 26503 2127 26537 2161
rect 26571 2127 26605 2161
rect 26639 2127 26673 2161
rect 26707 2127 26741 2161
rect 26775 2127 26809 2161
rect 26843 2127 26877 2161
rect 26911 2127 26945 2161
rect 26979 2127 27013 2161
rect 27047 2127 27081 2161
rect 27115 2127 27149 2161
rect 27183 2127 27217 2161
rect 27251 2127 27285 2161
rect 27319 2127 27353 2161
rect 27387 2127 27421 2161
rect 27455 2127 27489 2161
rect 27523 2127 27557 2161
rect 27591 2127 27625 2161
rect 27659 2127 27693 2161
rect 27727 2127 27761 2161
rect 27795 2127 27829 2161
rect 27863 2127 27897 2161
rect 27931 2127 27965 2161
rect 27999 2127 28033 2161
rect 28067 2127 28101 2161
rect 28135 2127 28169 2161
rect 28203 2127 28237 2161
rect 28271 2127 28305 2161
rect 28339 2127 28373 2161
rect 28407 2127 28441 2161
rect 28475 2127 28509 2161
rect 28543 2127 28577 2161
rect 28611 2127 28645 2161
rect 28679 2127 28713 2161
rect 28747 2127 28781 2161
rect 28815 2127 28849 2161
rect 28883 2127 28917 2161
rect 28951 2127 28985 2161
rect 29019 2127 29053 2161
rect 29087 2127 29121 2161
rect 29155 2127 29189 2161
rect 29223 2127 29257 2161
rect 29291 2127 29325 2161
rect 29359 2127 29393 2161
rect 29427 2127 29461 2161
rect 29495 2127 29529 2161
rect 29563 2127 29597 2161
rect 29631 2127 29665 2161
rect 29699 2127 29733 2161
rect 29767 2127 29801 2161
rect 29835 2127 29869 2161
rect 29903 2127 29937 2161
rect 29971 2127 30005 2161
rect 30039 2127 30073 2161
rect 30107 2127 30141 2161
rect 30175 2127 30209 2161
rect 30243 2127 30277 2161
rect 30311 2127 30345 2161
rect 30379 2127 30413 2161
rect 30447 2127 30481 2161
rect 30515 2127 30549 2161
rect 30583 2127 30617 2161
rect 30651 2127 30685 2161
rect 30719 2127 30753 2161
rect 30787 2127 30821 2161
rect 30855 2127 30889 2161
rect 30923 2127 30957 2161
rect 30991 2127 31025 2161
rect 31059 2127 31093 2161
rect 31127 2127 31161 2161
rect 31195 2127 31229 2161
rect 31263 2127 31452 2161
rect 26008 2094 31452 2127
rect 26008 2019 26108 2094
rect 26008 1985 26041 2019
rect 26075 1985 26108 2019
rect 26008 1951 26108 1985
rect 26008 1917 26041 1951
rect 26075 1917 26108 1951
rect 26008 1883 26108 1917
rect 26008 1849 26041 1883
rect 26075 1849 26108 1883
rect 26008 1815 26108 1849
rect 26008 1781 26041 1815
rect 26075 1781 26108 1815
rect 26008 1747 26108 1781
rect 26008 1713 26041 1747
rect 26075 1713 26108 1747
rect 26008 1679 26108 1713
rect 26008 1645 26041 1679
rect 26075 1645 26108 1679
rect 26008 1611 26108 1645
rect 26008 1577 26041 1611
rect 26075 1577 26108 1611
rect 26008 1543 26108 1577
rect 26008 1509 26041 1543
rect 26075 1509 26108 1543
rect 26008 1475 26108 1509
rect 26008 1441 26041 1475
rect 26075 1441 26108 1475
rect 26008 1407 26108 1441
rect 26008 1373 26041 1407
rect 26075 1373 26108 1407
rect 26008 1339 26108 1373
rect 26008 1305 26041 1339
rect 26075 1305 26108 1339
rect 26008 1271 26108 1305
rect 26008 1237 26041 1271
rect 26075 1237 26108 1271
rect 26008 1203 26108 1237
rect 26008 1169 26041 1203
rect 26075 1169 26108 1203
rect 26008 1135 26108 1169
rect 26008 1101 26041 1135
rect 26075 1101 26108 1135
rect 26008 1067 26108 1101
rect 26008 1033 26041 1067
rect 26075 1033 26108 1067
rect 26008 999 26108 1033
rect 26008 965 26041 999
rect 26075 965 26108 999
rect 26008 931 26108 965
rect 26008 897 26041 931
rect 26075 897 26108 931
rect 26008 863 26108 897
rect 26008 829 26041 863
rect 26075 829 26108 863
rect 26008 795 26108 829
rect 26008 761 26041 795
rect 26075 761 26108 795
rect 26008 727 26108 761
rect 26008 693 26041 727
rect 26075 693 26108 727
rect 26008 659 26108 693
rect 26008 625 26041 659
rect 26075 625 26108 659
rect 26008 591 26108 625
rect 26008 557 26041 591
rect 26075 557 26108 591
rect 26008 523 26108 557
rect 26008 489 26041 523
rect 26075 489 26108 523
rect 26008 455 26108 489
rect 26008 421 26041 455
rect 26075 421 26108 455
rect 26008 387 26108 421
rect 26008 353 26041 387
rect 26075 353 26108 387
rect 26008 319 26108 353
rect 26008 285 26041 319
rect 26075 285 26108 319
rect 26008 251 26108 285
rect 26008 217 26041 251
rect 26075 217 26108 251
rect 26008 183 26108 217
rect 26008 149 26041 183
rect 26075 149 26108 183
rect 26008 115 26108 149
rect 26008 81 26041 115
rect 26075 81 26108 115
rect 26008 47 26108 81
rect 26008 13 26041 47
rect 26075 13 26108 47
rect 26008 -21 26108 13
rect 26008 -55 26041 -21
rect 26075 -55 26108 -21
rect 26008 -89 26108 -55
rect 26008 -123 26041 -89
rect 26075 -123 26108 -89
rect 26008 -157 26108 -123
rect 26008 -191 26041 -157
rect 26075 -191 26108 -157
rect 26008 -225 26108 -191
rect 26008 -259 26041 -225
rect 26075 -259 26108 -225
rect 26008 -293 26108 -259
rect 26008 -327 26041 -293
rect 26075 -327 26108 -293
rect 26008 -361 26108 -327
rect 26008 -395 26041 -361
rect 26075 -395 26108 -361
rect 26008 -429 26108 -395
rect 26008 -463 26041 -429
rect 26075 -463 26108 -429
rect 26008 -497 26108 -463
rect 26008 -531 26041 -497
rect 26075 -531 26108 -497
rect 26008 -565 26108 -531
rect 26008 -599 26041 -565
rect 26075 -599 26108 -565
rect 26008 -633 26108 -599
rect 26008 -667 26041 -633
rect 26075 -667 26108 -633
rect 26008 -701 26108 -667
rect 26008 -735 26041 -701
rect 26075 -735 26108 -701
rect 26008 -769 26108 -735
rect 26008 -803 26041 -769
rect 26075 -803 26108 -769
rect 26008 -837 26108 -803
rect 26008 -871 26041 -837
rect 26075 -871 26108 -837
rect 26008 -905 26108 -871
rect 26008 -939 26041 -905
rect 26075 -939 26108 -905
rect 26008 -973 26108 -939
rect 26008 -1007 26041 -973
rect 26075 -1007 26108 -973
rect 26008 -1041 26108 -1007
rect 26008 -1075 26041 -1041
rect 26075 -1075 26108 -1041
rect 26008 -1109 26108 -1075
rect 26008 -1143 26041 -1109
rect 26075 -1143 26108 -1109
rect 26008 -1177 26108 -1143
rect 26008 -1211 26041 -1177
rect 26075 -1211 26108 -1177
rect 26008 -1245 26108 -1211
rect 26008 -1279 26041 -1245
rect 26075 -1279 26108 -1245
rect 26008 -1313 26108 -1279
rect 26008 -1347 26041 -1313
rect 26075 -1347 26108 -1313
rect 26008 -1381 26108 -1347
rect 26008 -1415 26041 -1381
rect 26075 -1415 26108 -1381
rect 26008 -1449 26108 -1415
rect 26008 -1483 26041 -1449
rect 26075 -1483 26108 -1449
rect 26008 -1558 26108 -1483
rect 31352 2019 31452 2094
rect 31352 1985 31385 2019
rect 31419 1985 31452 2019
rect 31352 1951 31452 1985
rect 31352 1917 31385 1951
rect 31419 1917 31452 1951
rect 31352 1883 31452 1917
rect 31352 1849 31385 1883
rect 31419 1849 31452 1883
rect 31352 1815 31452 1849
rect 31352 1781 31385 1815
rect 31419 1781 31452 1815
rect 31352 1747 31452 1781
rect 31352 1713 31385 1747
rect 31419 1713 31452 1747
rect 31352 1679 31452 1713
rect 31352 1645 31385 1679
rect 31419 1645 31452 1679
rect 31352 1611 31452 1645
rect 31352 1577 31385 1611
rect 31419 1577 31452 1611
rect 31352 1543 31452 1577
rect 31352 1509 31385 1543
rect 31419 1509 31452 1543
rect 31352 1475 31452 1509
rect 31352 1441 31385 1475
rect 31419 1441 31452 1475
rect 31352 1407 31452 1441
rect 31352 1373 31385 1407
rect 31419 1373 31452 1407
rect 31352 1339 31452 1373
rect 31352 1305 31385 1339
rect 31419 1305 31452 1339
rect 31352 1271 31452 1305
rect 31352 1237 31385 1271
rect 31419 1237 31452 1271
rect 31352 1203 31452 1237
rect 31352 1169 31385 1203
rect 31419 1169 31452 1203
rect 31352 1135 31452 1169
rect 31352 1101 31385 1135
rect 31419 1101 31452 1135
rect 31352 1067 31452 1101
rect 31352 1033 31385 1067
rect 31419 1033 31452 1067
rect 31352 999 31452 1033
rect 31352 965 31385 999
rect 31419 965 31452 999
rect 31352 931 31452 965
rect 31352 897 31385 931
rect 31419 897 31452 931
rect 31352 863 31452 897
rect 31352 829 31385 863
rect 31419 829 31452 863
rect 31352 795 31452 829
rect 31352 761 31385 795
rect 31419 761 31452 795
rect 31352 727 31452 761
rect 31352 693 31385 727
rect 31419 693 31452 727
rect 31352 659 31452 693
rect 31352 625 31385 659
rect 31419 625 31452 659
rect 31352 591 31452 625
rect 31352 557 31385 591
rect 31419 557 31452 591
rect 31352 523 31452 557
rect 31352 489 31385 523
rect 31419 489 31452 523
rect 31352 455 31452 489
rect 31352 421 31385 455
rect 31419 421 31452 455
rect 31352 387 31452 421
rect 31352 353 31385 387
rect 31419 353 31452 387
rect 31352 319 31452 353
rect 31352 285 31385 319
rect 31419 285 31452 319
rect 31352 251 31452 285
rect 31352 217 31385 251
rect 31419 217 31452 251
rect 31352 183 31452 217
rect 31352 149 31385 183
rect 31419 149 31452 183
rect 31352 115 31452 149
rect 31352 81 31385 115
rect 31419 81 31452 115
rect 31352 47 31452 81
rect 31352 13 31385 47
rect 31419 13 31452 47
rect 31352 -21 31452 13
rect 31352 -55 31385 -21
rect 31419 -55 31452 -21
rect 31352 -89 31452 -55
rect 31352 -123 31385 -89
rect 31419 -123 31452 -89
rect 31352 -157 31452 -123
rect 31352 -191 31385 -157
rect 31419 -191 31452 -157
rect 31352 -225 31452 -191
rect 31352 -259 31385 -225
rect 31419 -259 31452 -225
rect 31352 -293 31452 -259
rect 31352 -327 31385 -293
rect 31419 -327 31452 -293
rect 31352 -361 31452 -327
rect 31352 -395 31385 -361
rect 31419 -395 31452 -361
rect 31352 -429 31452 -395
rect 31352 -463 31385 -429
rect 31419 -463 31452 -429
rect 31352 -497 31452 -463
rect 31352 -531 31385 -497
rect 31419 -531 31452 -497
rect 31352 -565 31452 -531
rect 31352 -599 31385 -565
rect 31419 -599 31452 -565
rect 31352 -633 31452 -599
rect 31352 -667 31385 -633
rect 31419 -667 31452 -633
rect 31352 -701 31452 -667
rect 31352 -735 31385 -701
rect 31419 -735 31452 -701
rect 31352 -769 31452 -735
rect 31352 -803 31385 -769
rect 31419 -803 31452 -769
rect 31352 -837 31452 -803
rect 31352 -871 31385 -837
rect 31419 -871 31452 -837
rect 31352 -905 31452 -871
rect 31352 -939 31385 -905
rect 31419 -939 31452 -905
rect 31352 -973 31452 -939
rect 31352 -1007 31385 -973
rect 31419 -1007 31452 -973
rect 31352 -1041 31452 -1007
rect 31352 -1075 31385 -1041
rect 31419 -1075 31452 -1041
rect 31352 -1109 31452 -1075
rect 31352 -1143 31385 -1109
rect 31419 -1143 31452 -1109
rect 31352 -1177 31452 -1143
rect 31352 -1211 31385 -1177
rect 31419 -1211 31452 -1177
rect 31352 -1245 31452 -1211
rect 31352 -1279 31385 -1245
rect 31419 -1279 31452 -1245
rect 31352 -1313 31452 -1279
rect 31352 -1347 31385 -1313
rect 31419 -1347 31452 -1313
rect 31352 -1381 31452 -1347
rect 31352 -1415 31385 -1381
rect 31419 -1415 31452 -1381
rect 31352 -1449 31452 -1415
rect 31352 -1483 31385 -1449
rect 31419 -1483 31452 -1449
rect 31352 -1558 31452 -1483
rect 26008 -1591 31452 -1558
rect 26008 -1625 26197 -1591
rect 26231 -1625 26265 -1591
rect 26299 -1625 26333 -1591
rect 26367 -1625 26401 -1591
rect 26435 -1625 26469 -1591
rect 26503 -1625 26537 -1591
rect 26571 -1625 26605 -1591
rect 26639 -1625 26673 -1591
rect 26707 -1625 26741 -1591
rect 26775 -1625 26809 -1591
rect 26843 -1625 26877 -1591
rect 26911 -1625 26945 -1591
rect 26979 -1625 27013 -1591
rect 27047 -1625 27081 -1591
rect 27115 -1625 27149 -1591
rect 27183 -1625 27217 -1591
rect 27251 -1625 27285 -1591
rect 27319 -1625 27353 -1591
rect 27387 -1625 27421 -1591
rect 27455 -1625 27489 -1591
rect 27523 -1625 27557 -1591
rect 27591 -1625 27625 -1591
rect 27659 -1625 27693 -1591
rect 27727 -1625 27761 -1591
rect 27795 -1625 27829 -1591
rect 27863 -1625 27897 -1591
rect 27931 -1625 27965 -1591
rect 27999 -1625 28033 -1591
rect 28067 -1625 28101 -1591
rect 28135 -1625 28169 -1591
rect 28203 -1625 28237 -1591
rect 28271 -1625 28305 -1591
rect 28339 -1625 28373 -1591
rect 28407 -1625 28441 -1591
rect 28475 -1625 28509 -1591
rect 28543 -1625 28577 -1591
rect 28611 -1625 28645 -1591
rect 28679 -1625 28713 -1591
rect 28747 -1625 28781 -1591
rect 28815 -1625 28849 -1591
rect 28883 -1625 28917 -1591
rect 28951 -1625 28985 -1591
rect 29019 -1625 29053 -1591
rect 29087 -1625 29121 -1591
rect 29155 -1625 29189 -1591
rect 29223 -1625 29257 -1591
rect 29291 -1625 29325 -1591
rect 29359 -1625 29393 -1591
rect 29427 -1625 29461 -1591
rect 29495 -1625 29529 -1591
rect 29563 -1625 29597 -1591
rect 29631 -1625 29665 -1591
rect 29699 -1625 29733 -1591
rect 29767 -1625 29801 -1591
rect 29835 -1625 29869 -1591
rect 29903 -1625 29937 -1591
rect 29971 -1625 30005 -1591
rect 30039 -1625 30073 -1591
rect 30107 -1625 30141 -1591
rect 30175 -1625 30209 -1591
rect 30243 -1625 30277 -1591
rect 30311 -1625 30345 -1591
rect 30379 -1625 30413 -1591
rect 30447 -1625 30481 -1591
rect 30515 -1625 30549 -1591
rect 30583 -1625 30617 -1591
rect 30651 -1625 30685 -1591
rect 30719 -1625 30753 -1591
rect 30787 -1625 30821 -1591
rect 30855 -1625 30889 -1591
rect 30923 -1625 30957 -1591
rect 30991 -1625 31025 -1591
rect 31059 -1625 31093 -1591
rect 31127 -1625 31161 -1591
rect 31195 -1625 31229 -1591
rect 31263 -1625 31452 -1591
rect 26008 -1658 31452 -1625
<< psubdiffcont >>
rect 15603 4243 15637 4277
rect 15671 4243 15705 4277
rect 15739 4243 15773 4277
rect 15807 4243 15841 4277
rect 15875 4243 15909 4277
rect 15943 4243 15977 4277
rect 16011 4243 16045 4277
rect 16079 4243 16113 4277
rect 16147 4243 16181 4277
rect 16215 4243 16249 4277
rect 16283 4243 16317 4277
rect 16351 4243 16385 4277
rect 16419 4243 16453 4277
rect 16487 4243 16521 4277
rect 16555 4243 16589 4277
rect 16623 4243 16657 4277
rect 16691 4243 16725 4277
rect 16759 4243 16793 4277
rect 16827 4243 16861 4277
rect 16895 4243 16929 4277
rect 16963 4243 16997 4277
rect 17031 4243 17065 4277
rect 17099 4243 17133 4277
rect 17167 4243 17201 4277
rect 17235 4243 17269 4277
rect 17303 4243 17337 4277
rect 17371 4243 17405 4277
rect 17439 4243 17473 4277
rect 17507 4243 17541 4277
rect 17575 4243 17609 4277
rect 17643 4243 17677 4277
rect 17711 4243 17745 4277
rect 17779 4243 17813 4277
rect 17847 4243 17881 4277
rect 17915 4243 17949 4277
rect 17983 4243 18017 4277
rect 18051 4243 18085 4277
rect 18119 4243 18153 4277
rect 18187 4243 18221 4277
rect 18255 4243 18289 4277
rect 18323 4243 18357 4277
rect 18391 4243 18425 4277
rect 18459 4243 18493 4277
rect 18527 4243 18561 4277
rect 18595 4243 18629 4277
rect 18663 4243 18697 4277
rect 18731 4243 18765 4277
rect 18799 4243 18833 4277
rect 18867 4243 18901 4277
rect 18935 4243 18969 4277
rect 19003 4243 19037 4277
rect 19071 4243 19105 4277
rect 19139 4243 19173 4277
rect 19207 4243 19241 4277
rect 19275 4243 19309 4277
rect 19343 4243 19377 4277
rect 19411 4243 19445 4277
rect 19479 4243 19513 4277
rect 19547 4243 19581 4277
rect 19615 4243 19649 4277
rect 19683 4243 19717 4277
rect 19751 4243 19785 4277
rect 19819 4243 19853 4277
rect 19887 4243 19921 4277
rect 19955 4243 19989 4277
rect 20023 4243 20057 4277
rect 20091 4243 20125 4277
rect 20159 4243 20193 4277
rect 20227 4243 20261 4277
rect 20295 4243 20329 4277
rect 20363 4243 20397 4277
rect 20431 4243 20465 4277
rect 20499 4243 20533 4277
rect 20567 4243 20601 4277
rect 20635 4243 20669 4277
rect 20703 4243 20737 4277
rect 20771 4243 20805 4277
rect 20839 4243 20873 4277
rect 20907 4243 20941 4277
rect 20975 4243 21009 4277
rect 21043 4243 21077 4277
rect 21111 4243 21145 4277
rect 21179 4243 21213 4277
rect 21247 4243 21281 4277
rect 21315 4243 21349 4277
rect 21383 4243 21417 4277
rect 21451 4243 21485 4277
rect 21519 4243 21553 4277
rect 21587 4243 21621 4277
rect 21655 4243 21689 4277
rect 21723 4243 21757 4277
rect 21791 4243 21825 4277
rect 21859 4243 21893 4277
rect 21927 4243 21961 4277
rect 21995 4243 22029 4277
rect 22063 4243 22097 4277
rect 22131 4243 22165 4277
rect 22199 4243 22233 4277
rect 22267 4243 22301 4277
rect 22335 4243 22369 4277
rect 22403 4243 22437 4277
rect 22471 4243 22505 4277
rect 22539 4243 22573 4277
rect 22607 4243 22641 4277
rect 22675 4243 22709 4277
rect 22743 4243 22777 4277
rect 22811 4243 22845 4277
rect 22879 4243 22913 4277
rect 22947 4243 22981 4277
rect 23015 4243 23049 4277
rect 23083 4243 23117 4277
rect 23151 4243 23185 4277
rect 23219 4243 23253 4277
rect 23287 4243 23321 4277
rect 23355 4243 23389 4277
rect 23423 4243 23457 4277
rect 23491 4243 23525 4277
rect 23559 4243 23593 4277
rect 23627 4243 23661 4277
rect 23695 4243 23729 4277
rect 23763 4243 23797 4277
rect 23831 4243 23865 4277
rect 23899 4243 23933 4277
rect 23967 4243 24001 4277
rect 24035 4243 24069 4277
rect 24103 4243 24137 4277
rect 24171 4243 24205 4277
rect 24239 4243 24273 4277
rect 15459 4107 15493 4141
rect 15459 4039 15493 4073
rect 15459 3971 15493 4005
rect 15459 3903 15493 3937
rect 15459 3835 15493 3869
rect 15459 3767 15493 3801
rect 15459 3699 15493 3733
rect 15459 3631 15493 3665
rect 15459 3563 15493 3597
rect 15459 3495 15493 3529
rect 15459 3427 15493 3461
rect 15459 3359 15493 3393
rect 15459 3291 15493 3325
rect 15459 3223 15493 3257
rect 15459 3155 15493 3189
rect 15459 3087 15493 3121
rect 15459 3019 15493 3053
rect 15459 2951 15493 2985
rect 15459 2883 15493 2917
rect 15459 2815 15493 2849
rect 15459 2747 15493 2781
rect 15459 2679 15493 2713
rect 24383 4107 24417 4141
rect 24383 4039 24417 4073
rect 24383 3971 24417 4005
rect 24383 3903 24417 3937
rect 24383 3835 24417 3869
rect 24383 3767 24417 3801
rect 24383 3699 24417 3733
rect 24383 3631 24417 3665
rect 24383 3563 24417 3597
rect 24383 3495 24417 3529
rect 24383 3427 24417 3461
rect 24383 3359 24417 3393
rect 24383 3291 24417 3325
rect 24383 3223 24417 3257
rect 24383 3155 24417 3189
rect 24383 3087 24417 3121
rect 24383 3019 24417 3053
rect 24383 2951 24417 2985
rect 24383 2883 24417 2917
rect 24383 2815 24417 2849
rect 24383 2747 24417 2781
rect 24383 2679 24417 2713
rect 15603 2543 15637 2577
rect 15671 2543 15705 2577
rect 15739 2543 15773 2577
rect 15807 2543 15841 2577
rect 15875 2543 15909 2577
rect 15943 2543 15977 2577
rect 16011 2543 16045 2577
rect 16079 2543 16113 2577
rect 16147 2543 16181 2577
rect 16215 2543 16249 2577
rect 16283 2543 16317 2577
rect 16351 2543 16385 2577
rect 16419 2543 16453 2577
rect 16487 2543 16521 2577
rect 16555 2543 16589 2577
rect 16623 2543 16657 2577
rect 16691 2543 16725 2577
rect 16759 2543 16793 2577
rect 16827 2543 16861 2577
rect 16895 2543 16929 2577
rect 16963 2543 16997 2577
rect 17031 2543 17065 2577
rect 17099 2543 17133 2577
rect 17167 2543 17201 2577
rect 17235 2543 17269 2577
rect 17303 2543 17337 2577
rect 17371 2543 17405 2577
rect 17439 2543 17473 2577
rect 17507 2543 17541 2577
rect 17575 2543 17609 2577
rect 17643 2543 17677 2577
rect 17711 2543 17745 2577
rect 17779 2543 17813 2577
rect 17847 2543 17881 2577
rect 17915 2543 17949 2577
rect 17983 2543 18017 2577
rect 18051 2543 18085 2577
rect 18119 2543 18153 2577
rect 18187 2543 18221 2577
rect 18255 2543 18289 2577
rect 18323 2543 18357 2577
rect 18391 2543 18425 2577
rect 18459 2543 18493 2577
rect 18527 2543 18561 2577
rect 18595 2543 18629 2577
rect 18663 2543 18697 2577
rect 18731 2543 18765 2577
rect 18799 2543 18833 2577
rect 18867 2543 18901 2577
rect 18935 2543 18969 2577
rect 19003 2543 19037 2577
rect 19071 2543 19105 2577
rect 19139 2543 19173 2577
rect 19207 2543 19241 2577
rect 19275 2543 19309 2577
rect 19343 2543 19377 2577
rect 19411 2543 19445 2577
rect 19479 2543 19513 2577
rect 19547 2543 19581 2577
rect 19615 2543 19649 2577
rect 19683 2543 19717 2577
rect 19751 2543 19785 2577
rect 19819 2543 19853 2577
rect 19887 2543 19921 2577
rect 19955 2543 19989 2577
rect 20023 2543 20057 2577
rect 20091 2543 20125 2577
rect 20159 2543 20193 2577
rect 20227 2543 20261 2577
rect 20295 2543 20329 2577
rect 20363 2543 20397 2577
rect 20431 2543 20465 2577
rect 20499 2543 20533 2577
rect 20567 2543 20601 2577
rect 20635 2543 20669 2577
rect 20703 2543 20737 2577
rect 20771 2543 20805 2577
rect 20839 2543 20873 2577
rect 20907 2543 20941 2577
rect 20975 2543 21009 2577
rect 21043 2543 21077 2577
rect 21111 2543 21145 2577
rect 21179 2543 21213 2577
rect 21247 2543 21281 2577
rect 21315 2543 21349 2577
rect 21383 2543 21417 2577
rect 21451 2543 21485 2577
rect 21519 2543 21553 2577
rect 21587 2543 21621 2577
rect 21655 2543 21689 2577
rect 21723 2543 21757 2577
rect 21791 2543 21825 2577
rect 21859 2543 21893 2577
rect 21927 2543 21961 2577
rect 21995 2543 22029 2577
rect 22063 2543 22097 2577
rect 22131 2543 22165 2577
rect 22199 2543 22233 2577
rect 22267 2543 22301 2577
rect 22335 2543 22369 2577
rect 22403 2543 22437 2577
rect 22471 2543 22505 2577
rect 22539 2543 22573 2577
rect 22607 2543 22641 2577
rect 22675 2543 22709 2577
rect 22743 2543 22777 2577
rect 22811 2543 22845 2577
rect 22879 2543 22913 2577
rect 22947 2543 22981 2577
rect 23015 2543 23049 2577
rect 23083 2543 23117 2577
rect 23151 2543 23185 2577
rect 23219 2543 23253 2577
rect 23287 2543 23321 2577
rect 23355 2543 23389 2577
rect 23423 2543 23457 2577
rect 23491 2543 23525 2577
rect 23559 2543 23593 2577
rect 23627 2543 23661 2577
rect 23695 2543 23729 2577
rect 23763 2543 23797 2577
rect 23831 2543 23865 2577
rect 23899 2543 23933 2577
rect 23967 2543 24001 2577
rect 24035 2543 24069 2577
rect 24103 2543 24137 2577
rect 24171 2543 24205 2577
rect 24239 2543 24273 2577
rect 26197 4243 26231 4277
rect 26265 4243 26299 4277
rect 26333 4243 26367 4277
rect 26401 4243 26435 4277
rect 26469 4243 26503 4277
rect 26537 4243 26571 4277
rect 26605 4243 26639 4277
rect 26673 4243 26707 4277
rect 26741 4243 26775 4277
rect 26809 4243 26843 4277
rect 26877 4243 26911 4277
rect 26945 4243 26979 4277
rect 27013 4243 27047 4277
rect 27081 4243 27115 4277
rect 27149 4243 27183 4277
rect 27217 4243 27251 4277
rect 27285 4243 27319 4277
rect 27353 4243 27387 4277
rect 27421 4243 27455 4277
rect 27489 4243 27523 4277
rect 27557 4243 27591 4277
rect 27625 4243 27659 4277
rect 27693 4243 27727 4277
rect 27761 4243 27795 4277
rect 27829 4243 27863 4277
rect 27897 4243 27931 4277
rect 27965 4243 27999 4277
rect 28033 4243 28067 4277
rect 28101 4243 28135 4277
rect 28169 4243 28203 4277
rect 28237 4243 28271 4277
rect 28305 4243 28339 4277
rect 28373 4243 28407 4277
rect 28441 4243 28475 4277
rect 28509 4243 28543 4277
rect 28577 4243 28611 4277
rect 28645 4243 28679 4277
rect 28713 4243 28747 4277
rect 28781 4243 28815 4277
rect 28849 4243 28883 4277
rect 28917 4243 28951 4277
rect 28985 4243 29019 4277
rect 29053 4243 29087 4277
rect 29121 4243 29155 4277
rect 29189 4243 29223 4277
rect 29257 4243 29291 4277
rect 29325 4243 29359 4277
rect 29393 4243 29427 4277
rect 29461 4243 29495 4277
rect 29529 4243 29563 4277
rect 29597 4243 29631 4277
rect 29665 4243 29699 4277
rect 29733 4243 29767 4277
rect 29801 4243 29835 4277
rect 29869 4243 29903 4277
rect 29937 4243 29971 4277
rect 30005 4243 30039 4277
rect 30073 4243 30107 4277
rect 30141 4243 30175 4277
rect 30209 4243 30243 4277
rect 30277 4243 30311 4277
rect 30345 4243 30379 4277
rect 30413 4243 30447 4277
rect 30481 4243 30515 4277
rect 30549 4243 30583 4277
rect 30617 4243 30651 4277
rect 30685 4243 30719 4277
rect 30753 4243 30787 4277
rect 30821 4243 30855 4277
rect 30889 4243 30923 4277
rect 30957 4243 30991 4277
rect 31025 4243 31059 4277
rect 31093 4243 31127 4277
rect 31161 4243 31195 4277
rect 31229 4243 31263 4277
rect 26041 4101 26075 4135
rect 26041 4033 26075 4067
rect 26041 3965 26075 3999
rect 26041 3897 26075 3931
rect 26041 3829 26075 3863
rect 26041 3761 26075 3795
rect 26041 3693 26075 3727
rect 26041 3625 26075 3659
rect 26041 3557 26075 3591
rect 26041 3489 26075 3523
rect 26041 3421 26075 3455
rect 26041 3353 26075 3387
rect 26041 3285 26075 3319
rect 26041 3217 26075 3251
rect 26041 3149 26075 3183
rect 26041 3081 26075 3115
rect 26041 3013 26075 3047
rect 26041 2945 26075 2979
rect 26041 2877 26075 2911
rect 26041 2809 26075 2843
rect 26041 2741 26075 2775
rect 26041 2673 26075 2707
rect 26041 2605 26075 2639
rect 31385 4101 31419 4135
rect 31385 4033 31419 4067
rect 31385 3965 31419 3999
rect 31385 3897 31419 3931
rect 31385 3829 31419 3863
rect 31385 3761 31419 3795
rect 31385 3693 31419 3727
rect 31385 3625 31419 3659
rect 31385 3557 31419 3591
rect 31385 3489 31419 3523
rect 31385 3421 31419 3455
rect 31385 3353 31419 3387
rect 31385 3285 31419 3319
rect 31385 3217 31419 3251
rect 31385 3149 31419 3183
rect 31385 3081 31419 3115
rect 31385 3013 31419 3047
rect 31385 2945 31419 2979
rect 31385 2877 31419 2911
rect 31385 2809 31419 2843
rect 31385 2741 31419 2775
rect 31385 2673 31419 2707
rect 31385 2605 31419 2639
rect 26197 2463 26231 2497
rect 26265 2463 26299 2497
rect 26333 2463 26367 2497
rect 26401 2463 26435 2497
rect 26469 2463 26503 2497
rect 26537 2463 26571 2497
rect 26605 2463 26639 2497
rect 26673 2463 26707 2497
rect 26741 2463 26775 2497
rect 26809 2463 26843 2497
rect 26877 2463 26911 2497
rect 26945 2463 26979 2497
rect 27013 2463 27047 2497
rect 27081 2463 27115 2497
rect 27149 2463 27183 2497
rect 27217 2463 27251 2497
rect 27285 2463 27319 2497
rect 27353 2463 27387 2497
rect 27421 2463 27455 2497
rect 27489 2463 27523 2497
rect 27557 2463 27591 2497
rect 27625 2463 27659 2497
rect 27693 2463 27727 2497
rect 27761 2463 27795 2497
rect 27829 2463 27863 2497
rect 27897 2463 27931 2497
rect 27965 2463 27999 2497
rect 28033 2463 28067 2497
rect 28101 2463 28135 2497
rect 28169 2463 28203 2497
rect 28237 2463 28271 2497
rect 28305 2463 28339 2497
rect 28373 2463 28407 2497
rect 28441 2463 28475 2497
rect 28509 2463 28543 2497
rect 28577 2463 28611 2497
rect 28645 2463 28679 2497
rect 28713 2463 28747 2497
rect 28781 2463 28815 2497
rect 28849 2463 28883 2497
rect 28917 2463 28951 2497
rect 28985 2463 29019 2497
rect 29053 2463 29087 2497
rect 29121 2463 29155 2497
rect 29189 2463 29223 2497
rect 29257 2463 29291 2497
rect 29325 2463 29359 2497
rect 29393 2463 29427 2497
rect 29461 2463 29495 2497
rect 29529 2463 29563 2497
rect 29597 2463 29631 2497
rect 29665 2463 29699 2497
rect 29733 2463 29767 2497
rect 29801 2463 29835 2497
rect 29869 2463 29903 2497
rect 29937 2463 29971 2497
rect 30005 2463 30039 2497
rect 30073 2463 30107 2497
rect 30141 2463 30175 2497
rect 30209 2463 30243 2497
rect 30277 2463 30311 2497
rect 30345 2463 30379 2497
rect 30413 2463 30447 2497
rect 30481 2463 30515 2497
rect 30549 2463 30583 2497
rect 30617 2463 30651 2497
rect 30685 2463 30719 2497
rect 30753 2463 30787 2497
rect 30821 2463 30855 2497
rect 30889 2463 30923 2497
rect 30957 2463 30991 2497
rect 31025 2463 31059 2497
rect 31093 2463 31127 2497
rect 31161 2463 31195 2497
rect 31229 2463 31263 2497
<< nsubdiffcont >>
rect 15603 2207 15637 2241
rect 15671 2207 15705 2241
rect 15739 2207 15773 2241
rect 15807 2207 15841 2241
rect 15875 2207 15909 2241
rect 15943 2207 15977 2241
rect 16011 2207 16045 2241
rect 16079 2207 16113 2241
rect 16147 2207 16181 2241
rect 16215 2207 16249 2241
rect 16283 2207 16317 2241
rect 16351 2207 16385 2241
rect 16419 2207 16453 2241
rect 16487 2207 16521 2241
rect 16555 2207 16589 2241
rect 16623 2207 16657 2241
rect 16691 2207 16725 2241
rect 16759 2207 16793 2241
rect 16827 2207 16861 2241
rect 16895 2207 16929 2241
rect 16963 2207 16997 2241
rect 17031 2207 17065 2241
rect 17099 2207 17133 2241
rect 17167 2207 17201 2241
rect 17235 2207 17269 2241
rect 17303 2207 17337 2241
rect 17371 2207 17405 2241
rect 17439 2207 17473 2241
rect 17507 2207 17541 2241
rect 17575 2207 17609 2241
rect 17643 2207 17677 2241
rect 17711 2207 17745 2241
rect 17779 2207 17813 2241
rect 17847 2207 17881 2241
rect 17915 2207 17949 2241
rect 17983 2207 18017 2241
rect 18051 2207 18085 2241
rect 18119 2207 18153 2241
rect 18187 2207 18221 2241
rect 18255 2207 18289 2241
rect 18323 2207 18357 2241
rect 18391 2207 18425 2241
rect 18459 2207 18493 2241
rect 18527 2207 18561 2241
rect 18595 2207 18629 2241
rect 18663 2207 18697 2241
rect 18731 2207 18765 2241
rect 18799 2207 18833 2241
rect 18867 2207 18901 2241
rect 18935 2207 18969 2241
rect 19003 2207 19037 2241
rect 19071 2207 19105 2241
rect 19139 2207 19173 2241
rect 19207 2207 19241 2241
rect 19275 2207 19309 2241
rect 19343 2207 19377 2241
rect 19411 2207 19445 2241
rect 19479 2207 19513 2241
rect 19547 2207 19581 2241
rect 19615 2207 19649 2241
rect 19683 2207 19717 2241
rect 19751 2207 19785 2241
rect 19819 2207 19853 2241
rect 19887 2207 19921 2241
rect 19955 2207 19989 2241
rect 20023 2207 20057 2241
rect 20091 2207 20125 2241
rect 20159 2207 20193 2241
rect 20227 2207 20261 2241
rect 20295 2207 20329 2241
rect 20363 2207 20397 2241
rect 20431 2207 20465 2241
rect 20499 2207 20533 2241
rect 20567 2207 20601 2241
rect 20635 2207 20669 2241
rect 20703 2207 20737 2241
rect 20771 2207 20805 2241
rect 20839 2207 20873 2241
rect 20907 2207 20941 2241
rect 20975 2207 21009 2241
rect 21043 2207 21077 2241
rect 21111 2207 21145 2241
rect 21179 2207 21213 2241
rect 21247 2207 21281 2241
rect 21315 2207 21349 2241
rect 21383 2207 21417 2241
rect 21451 2207 21485 2241
rect 21519 2207 21553 2241
rect 21587 2207 21621 2241
rect 21655 2207 21689 2241
rect 21723 2207 21757 2241
rect 21791 2207 21825 2241
rect 21859 2207 21893 2241
rect 21927 2207 21961 2241
rect 21995 2207 22029 2241
rect 22063 2207 22097 2241
rect 22131 2207 22165 2241
rect 22199 2207 22233 2241
rect 22267 2207 22301 2241
rect 22335 2207 22369 2241
rect 22403 2207 22437 2241
rect 22471 2207 22505 2241
rect 22539 2207 22573 2241
rect 22607 2207 22641 2241
rect 22675 2207 22709 2241
rect 22743 2207 22777 2241
rect 22811 2207 22845 2241
rect 22879 2207 22913 2241
rect 22947 2207 22981 2241
rect 23015 2207 23049 2241
rect 23083 2207 23117 2241
rect 23151 2207 23185 2241
rect 23219 2207 23253 2241
rect 23287 2207 23321 2241
rect 23355 2207 23389 2241
rect 23423 2207 23457 2241
rect 23491 2207 23525 2241
rect 23559 2207 23593 2241
rect 23627 2207 23661 2241
rect 23695 2207 23729 2241
rect 23763 2207 23797 2241
rect 23831 2207 23865 2241
rect 23899 2207 23933 2241
rect 23967 2207 24001 2241
rect 24035 2207 24069 2241
rect 24103 2207 24137 2241
rect 24171 2207 24205 2241
rect 24239 2207 24273 2241
rect 15459 2059 15493 2093
rect 15459 1991 15493 2025
rect 15459 1923 15493 1957
rect 15459 1855 15493 1889
rect 15459 1787 15493 1821
rect 15459 1719 15493 1753
rect 15459 1651 15493 1685
rect 15459 1583 15493 1617
rect 15459 1515 15493 1549
rect 15459 1447 15493 1481
rect 15459 1379 15493 1413
rect 15459 1311 15493 1345
rect 15459 1243 15493 1277
rect 15459 1175 15493 1209
rect 15459 1107 15493 1141
rect 15459 1039 15493 1073
rect 15459 971 15493 1005
rect 15459 903 15493 937
rect 15459 835 15493 869
rect 15459 767 15493 801
rect 15459 699 15493 733
rect 15459 631 15493 665
rect 15459 563 15493 597
rect 15459 495 15493 529
rect 15459 427 15493 461
rect 15459 359 15493 393
rect 15459 291 15493 325
rect 15459 223 15493 257
rect 15459 155 15493 189
rect 15459 87 15493 121
rect 15459 19 15493 53
rect 15459 -49 15493 -15
rect 15459 -117 15493 -83
rect 15459 -185 15493 -151
rect 15459 -253 15493 -219
rect 15459 -321 15493 -287
rect 15459 -389 15493 -355
rect 15459 -457 15493 -423
rect 15459 -525 15493 -491
rect 15459 -593 15493 -559
rect 15459 -661 15493 -627
rect 15459 -729 15493 -695
rect 15459 -797 15493 -763
rect 15459 -865 15493 -831
rect 15459 -933 15493 -899
rect 15459 -1001 15493 -967
rect 15459 -1069 15493 -1035
rect 15459 -1137 15493 -1103
rect 15459 -1205 15493 -1171
rect 15459 -1273 15493 -1239
rect 15459 -1341 15493 -1307
rect 15459 -1409 15493 -1375
rect 15459 -1477 15493 -1443
rect 24383 2059 24417 2093
rect 24383 1991 24417 2025
rect 24383 1923 24417 1957
rect 24383 1855 24417 1889
rect 24383 1787 24417 1821
rect 24383 1719 24417 1753
rect 24383 1651 24417 1685
rect 24383 1583 24417 1617
rect 24383 1515 24417 1549
rect 24383 1447 24417 1481
rect 24383 1379 24417 1413
rect 24383 1311 24417 1345
rect 24383 1243 24417 1277
rect 24383 1175 24417 1209
rect 24383 1107 24417 1141
rect 24383 1039 24417 1073
rect 24383 971 24417 1005
rect 24383 903 24417 937
rect 24383 835 24417 869
rect 24383 767 24417 801
rect 24383 699 24417 733
rect 24383 631 24417 665
rect 24383 563 24417 597
rect 24383 495 24417 529
rect 24383 427 24417 461
rect 24383 359 24417 393
rect 24383 291 24417 325
rect 24383 223 24417 257
rect 24383 155 24417 189
rect 24383 87 24417 121
rect 24383 19 24417 53
rect 24383 -49 24417 -15
rect 24383 -117 24417 -83
rect 24383 -185 24417 -151
rect 24383 -253 24417 -219
rect 24383 -321 24417 -287
rect 24383 -389 24417 -355
rect 24383 -457 24417 -423
rect 24383 -525 24417 -491
rect 24383 -593 24417 -559
rect 24383 -661 24417 -627
rect 24383 -729 24417 -695
rect 24383 -797 24417 -763
rect 24383 -865 24417 -831
rect 24383 -933 24417 -899
rect 24383 -1001 24417 -967
rect 24383 -1069 24417 -1035
rect 24383 -1137 24417 -1103
rect 24383 -1205 24417 -1171
rect 24383 -1273 24417 -1239
rect 24383 -1341 24417 -1307
rect 24383 -1409 24417 -1375
rect 24383 -1477 24417 -1443
rect 15603 -1625 15637 -1591
rect 15671 -1625 15705 -1591
rect 15739 -1625 15773 -1591
rect 15807 -1625 15841 -1591
rect 15875 -1625 15909 -1591
rect 15943 -1625 15977 -1591
rect 16011 -1625 16045 -1591
rect 16079 -1625 16113 -1591
rect 16147 -1625 16181 -1591
rect 16215 -1625 16249 -1591
rect 16283 -1625 16317 -1591
rect 16351 -1625 16385 -1591
rect 16419 -1625 16453 -1591
rect 16487 -1625 16521 -1591
rect 16555 -1625 16589 -1591
rect 16623 -1625 16657 -1591
rect 16691 -1625 16725 -1591
rect 16759 -1625 16793 -1591
rect 16827 -1625 16861 -1591
rect 16895 -1625 16929 -1591
rect 16963 -1625 16997 -1591
rect 17031 -1625 17065 -1591
rect 17099 -1625 17133 -1591
rect 17167 -1625 17201 -1591
rect 17235 -1625 17269 -1591
rect 17303 -1625 17337 -1591
rect 17371 -1625 17405 -1591
rect 17439 -1625 17473 -1591
rect 17507 -1625 17541 -1591
rect 17575 -1625 17609 -1591
rect 17643 -1625 17677 -1591
rect 17711 -1625 17745 -1591
rect 17779 -1625 17813 -1591
rect 17847 -1625 17881 -1591
rect 17915 -1625 17949 -1591
rect 17983 -1625 18017 -1591
rect 18051 -1625 18085 -1591
rect 18119 -1625 18153 -1591
rect 18187 -1625 18221 -1591
rect 18255 -1625 18289 -1591
rect 18323 -1625 18357 -1591
rect 18391 -1625 18425 -1591
rect 18459 -1625 18493 -1591
rect 18527 -1625 18561 -1591
rect 18595 -1625 18629 -1591
rect 18663 -1625 18697 -1591
rect 18731 -1625 18765 -1591
rect 18799 -1625 18833 -1591
rect 18867 -1625 18901 -1591
rect 18935 -1625 18969 -1591
rect 19003 -1625 19037 -1591
rect 19071 -1625 19105 -1591
rect 19139 -1625 19173 -1591
rect 19207 -1625 19241 -1591
rect 19275 -1625 19309 -1591
rect 19343 -1625 19377 -1591
rect 19411 -1625 19445 -1591
rect 19479 -1625 19513 -1591
rect 19547 -1625 19581 -1591
rect 19615 -1625 19649 -1591
rect 19683 -1625 19717 -1591
rect 19751 -1625 19785 -1591
rect 19819 -1625 19853 -1591
rect 19887 -1625 19921 -1591
rect 19955 -1625 19989 -1591
rect 20023 -1625 20057 -1591
rect 20091 -1625 20125 -1591
rect 20159 -1625 20193 -1591
rect 20227 -1625 20261 -1591
rect 20295 -1625 20329 -1591
rect 20363 -1625 20397 -1591
rect 20431 -1625 20465 -1591
rect 20499 -1625 20533 -1591
rect 20567 -1625 20601 -1591
rect 20635 -1625 20669 -1591
rect 20703 -1625 20737 -1591
rect 20771 -1625 20805 -1591
rect 20839 -1625 20873 -1591
rect 20907 -1625 20941 -1591
rect 20975 -1625 21009 -1591
rect 21043 -1625 21077 -1591
rect 21111 -1625 21145 -1591
rect 21179 -1625 21213 -1591
rect 21247 -1625 21281 -1591
rect 21315 -1625 21349 -1591
rect 21383 -1625 21417 -1591
rect 21451 -1625 21485 -1591
rect 21519 -1625 21553 -1591
rect 21587 -1625 21621 -1591
rect 21655 -1625 21689 -1591
rect 21723 -1625 21757 -1591
rect 21791 -1625 21825 -1591
rect 21859 -1625 21893 -1591
rect 21927 -1625 21961 -1591
rect 21995 -1625 22029 -1591
rect 22063 -1625 22097 -1591
rect 22131 -1625 22165 -1591
rect 22199 -1625 22233 -1591
rect 22267 -1625 22301 -1591
rect 22335 -1625 22369 -1591
rect 22403 -1625 22437 -1591
rect 22471 -1625 22505 -1591
rect 22539 -1625 22573 -1591
rect 22607 -1625 22641 -1591
rect 22675 -1625 22709 -1591
rect 22743 -1625 22777 -1591
rect 22811 -1625 22845 -1591
rect 22879 -1625 22913 -1591
rect 22947 -1625 22981 -1591
rect 23015 -1625 23049 -1591
rect 23083 -1625 23117 -1591
rect 23151 -1625 23185 -1591
rect 23219 -1625 23253 -1591
rect 23287 -1625 23321 -1591
rect 23355 -1625 23389 -1591
rect 23423 -1625 23457 -1591
rect 23491 -1625 23525 -1591
rect 23559 -1625 23593 -1591
rect 23627 -1625 23661 -1591
rect 23695 -1625 23729 -1591
rect 23763 -1625 23797 -1591
rect 23831 -1625 23865 -1591
rect 23899 -1625 23933 -1591
rect 23967 -1625 24001 -1591
rect 24035 -1625 24069 -1591
rect 24103 -1625 24137 -1591
rect 24171 -1625 24205 -1591
rect 24239 -1625 24273 -1591
rect 26197 2127 26231 2161
rect 26265 2127 26299 2161
rect 26333 2127 26367 2161
rect 26401 2127 26435 2161
rect 26469 2127 26503 2161
rect 26537 2127 26571 2161
rect 26605 2127 26639 2161
rect 26673 2127 26707 2161
rect 26741 2127 26775 2161
rect 26809 2127 26843 2161
rect 26877 2127 26911 2161
rect 26945 2127 26979 2161
rect 27013 2127 27047 2161
rect 27081 2127 27115 2161
rect 27149 2127 27183 2161
rect 27217 2127 27251 2161
rect 27285 2127 27319 2161
rect 27353 2127 27387 2161
rect 27421 2127 27455 2161
rect 27489 2127 27523 2161
rect 27557 2127 27591 2161
rect 27625 2127 27659 2161
rect 27693 2127 27727 2161
rect 27761 2127 27795 2161
rect 27829 2127 27863 2161
rect 27897 2127 27931 2161
rect 27965 2127 27999 2161
rect 28033 2127 28067 2161
rect 28101 2127 28135 2161
rect 28169 2127 28203 2161
rect 28237 2127 28271 2161
rect 28305 2127 28339 2161
rect 28373 2127 28407 2161
rect 28441 2127 28475 2161
rect 28509 2127 28543 2161
rect 28577 2127 28611 2161
rect 28645 2127 28679 2161
rect 28713 2127 28747 2161
rect 28781 2127 28815 2161
rect 28849 2127 28883 2161
rect 28917 2127 28951 2161
rect 28985 2127 29019 2161
rect 29053 2127 29087 2161
rect 29121 2127 29155 2161
rect 29189 2127 29223 2161
rect 29257 2127 29291 2161
rect 29325 2127 29359 2161
rect 29393 2127 29427 2161
rect 29461 2127 29495 2161
rect 29529 2127 29563 2161
rect 29597 2127 29631 2161
rect 29665 2127 29699 2161
rect 29733 2127 29767 2161
rect 29801 2127 29835 2161
rect 29869 2127 29903 2161
rect 29937 2127 29971 2161
rect 30005 2127 30039 2161
rect 30073 2127 30107 2161
rect 30141 2127 30175 2161
rect 30209 2127 30243 2161
rect 30277 2127 30311 2161
rect 30345 2127 30379 2161
rect 30413 2127 30447 2161
rect 30481 2127 30515 2161
rect 30549 2127 30583 2161
rect 30617 2127 30651 2161
rect 30685 2127 30719 2161
rect 30753 2127 30787 2161
rect 30821 2127 30855 2161
rect 30889 2127 30923 2161
rect 30957 2127 30991 2161
rect 31025 2127 31059 2161
rect 31093 2127 31127 2161
rect 31161 2127 31195 2161
rect 31229 2127 31263 2161
rect 26041 1985 26075 2019
rect 26041 1917 26075 1951
rect 26041 1849 26075 1883
rect 26041 1781 26075 1815
rect 26041 1713 26075 1747
rect 26041 1645 26075 1679
rect 26041 1577 26075 1611
rect 26041 1509 26075 1543
rect 26041 1441 26075 1475
rect 26041 1373 26075 1407
rect 26041 1305 26075 1339
rect 26041 1237 26075 1271
rect 26041 1169 26075 1203
rect 26041 1101 26075 1135
rect 26041 1033 26075 1067
rect 26041 965 26075 999
rect 26041 897 26075 931
rect 26041 829 26075 863
rect 26041 761 26075 795
rect 26041 693 26075 727
rect 26041 625 26075 659
rect 26041 557 26075 591
rect 26041 489 26075 523
rect 26041 421 26075 455
rect 26041 353 26075 387
rect 26041 285 26075 319
rect 26041 217 26075 251
rect 26041 149 26075 183
rect 26041 81 26075 115
rect 26041 13 26075 47
rect 26041 -55 26075 -21
rect 26041 -123 26075 -89
rect 26041 -191 26075 -157
rect 26041 -259 26075 -225
rect 26041 -327 26075 -293
rect 26041 -395 26075 -361
rect 26041 -463 26075 -429
rect 26041 -531 26075 -497
rect 26041 -599 26075 -565
rect 26041 -667 26075 -633
rect 26041 -735 26075 -701
rect 26041 -803 26075 -769
rect 26041 -871 26075 -837
rect 26041 -939 26075 -905
rect 26041 -1007 26075 -973
rect 26041 -1075 26075 -1041
rect 26041 -1143 26075 -1109
rect 26041 -1211 26075 -1177
rect 26041 -1279 26075 -1245
rect 26041 -1347 26075 -1313
rect 26041 -1415 26075 -1381
rect 26041 -1483 26075 -1449
rect 31385 1985 31419 2019
rect 31385 1917 31419 1951
rect 31385 1849 31419 1883
rect 31385 1781 31419 1815
rect 31385 1713 31419 1747
rect 31385 1645 31419 1679
rect 31385 1577 31419 1611
rect 31385 1509 31419 1543
rect 31385 1441 31419 1475
rect 31385 1373 31419 1407
rect 31385 1305 31419 1339
rect 31385 1237 31419 1271
rect 31385 1169 31419 1203
rect 31385 1101 31419 1135
rect 31385 1033 31419 1067
rect 31385 965 31419 999
rect 31385 897 31419 931
rect 31385 829 31419 863
rect 31385 761 31419 795
rect 31385 693 31419 727
rect 31385 625 31419 659
rect 31385 557 31419 591
rect 31385 489 31419 523
rect 31385 421 31419 455
rect 31385 353 31419 387
rect 31385 285 31419 319
rect 31385 217 31419 251
rect 31385 149 31419 183
rect 31385 81 31419 115
rect 31385 13 31419 47
rect 31385 -55 31419 -21
rect 31385 -123 31419 -89
rect 31385 -191 31419 -157
rect 31385 -259 31419 -225
rect 31385 -327 31419 -293
rect 31385 -395 31419 -361
rect 31385 -463 31419 -429
rect 31385 -531 31419 -497
rect 31385 -599 31419 -565
rect 31385 -667 31419 -633
rect 31385 -735 31419 -701
rect 31385 -803 31419 -769
rect 31385 -871 31419 -837
rect 31385 -939 31419 -905
rect 31385 -1007 31419 -973
rect 31385 -1075 31419 -1041
rect 31385 -1143 31419 -1109
rect 31385 -1211 31419 -1177
rect 31385 -1279 31419 -1245
rect 31385 -1347 31419 -1313
rect 31385 -1415 31419 -1381
rect 31385 -1483 31419 -1449
rect 26197 -1625 26231 -1591
rect 26265 -1625 26299 -1591
rect 26333 -1625 26367 -1591
rect 26401 -1625 26435 -1591
rect 26469 -1625 26503 -1591
rect 26537 -1625 26571 -1591
rect 26605 -1625 26639 -1591
rect 26673 -1625 26707 -1591
rect 26741 -1625 26775 -1591
rect 26809 -1625 26843 -1591
rect 26877 -1625 26911 -1591
rect 26945 -1625 26979 -1591
rect 27013 -1625 27047 -1591
rect 27081 -1625 27115 -1591
rect 27149 -1625 27183 -1591
rect 27217 -1625 27251 -1591
rect 27285 -1625 27319 -1591
rect 27353 -1625 27387 -1591
rect 27421 -1625 27455 -1591
rect 27489 -1625 27523 -1591
rect 27557 -1625 27591 -1591
rect 27625 -1625 27659 -1591
rect 27693 -1625 27727 -1591
rect 27761 -1625 27795 -1591
rect 27829 -1625 27863 -1591
rect 27897 -1625 27931 -1591
rect 27965 -1625 27999 -1591
rect 28033 -1625 28067 -1591
rect 28101 -1625 28135 -1591
rect 28169 -1625 28203 -1591
rect 28237 -1625 28271 -1591
rect 28305 -1625 28339 -1591
rect 28373 -1625 28407 -1591
rect 28441 -1625 28475 -1591
rect 28509 -1625 28543 -1591
rect 28577 -1625 28611 -1591
rect 28645 -1625 28679 -1591
rect 28713 -1625 28747 -1591
rect 28781 -1625 28815 -1591
rect 28849 -1625 28883 -1591
rect 28917 -1625 28951 -1591
rect 28985 -1625 29019 -1591
rect 29053 -1625 29087 -1591
rect 29121 -1625 29155 -1591
rect 29189 -1625 29223 -1591
rect 29257 -1625 29291 -1591
rect 29325 -1625 29359 -1591
rect 29393 -1625 29427 -1591
rect 29461 -1625 29495 -1591
rect 29529 -1625 29563 -1591
rect 29597 -1625 29631 -1591
rect 29665 -1625 29699 -1591
rect 29733 -1625 29767 -1591
rect 29801 -1625 29835 -1591
rect 29869 -1625 29903 -1591
rect 29937 -1625 29971 -1591
rect 30005 -1625 30039 -1591
rect 30073 -1625 30107 -1591
rect 30141 -1625 30175 -1591
rect 30209 -1625 30243 -1591
rect 30277 -1625 30311 -1591
rect 30345 -1625 30379 -1591
rect 30413 -1625 30447 -1591
rect 30481 -1625 30515 -1591
rect 30549 -1625 30583 -1591
rect 30617 -1625 30651 -1591
rect 30685 -1625 30719 -1591
rect 30753 -1625 30787 -1591
rect 30821 -1625 30855 -1591
rect 30889 -1625 30923 -1591
rect 30957 -1625 30991 -1591
rect 31025 -1625 31059 -1591
rect 31093 -1625 31127 -1591
rect 31161 -1625 31195 -1591
rect 31229 -1625 31263 -1591
<< locali >>
rect 15426 4277 24450 4310
rect 15426 4243 15529 4277
rect 15563 4243 15601 4277
rect 15637 4243 15671 4277
rect 15707 4243 15739 4277
rect 15779 4243 15807 4277
rect 15851 4243 15875 4277
rect 15923 4243 15943 4277
rect 15995 4243 16011 4277
rect 16067 4243 16079 4277
rect 16139 4243 16147 4277
rect 16211 4243 16215 4277
rect 16317 4243 16321 4277
rect 16385 4243 16393 4277
rect 16453 4243 16465 4277
rect 16521 4243 16537 4277
rect 16589 4243 16609 4277
rect 16657 4243 16681 4277
rect 16725 4243 16753 4277
rect 16793 4243 16825 4277
rect 16861 4243 16895 4277
rect 16931 4243 16963 4277
rect 17003 4243 17031 4277
rect 17075 4243 17099 4277
rect 17147 4243 17167 4277
rect 17219 4243 17235 4277
rect 17291 4243 17303 4277
rect 17363 4243 17371 4277
rect 17435 4243 17439 4277
rect 17541 4243 17545 4277
rect 17609 4243 17617 4277
rect 17677 4243 17689 4277
rect 17745 4243 17761 4277
rect 17813 4243 17833 4277
rect 17881 4243 17905 4277
rect 17949 4243 17977 4277
rect 18017 4243 18049 4277
rect 18085 4243 18119 4277
rect 18155 4243 18187 4277
rect 18227 4243 18255 4277
rect 18299 4243 18323 4277
rect 18371 4243 18391 4277
rect 18443 4243 18459 4277
rect 18515 4243 18527 4277
rect 18587 4243 18595 4277
rect 18659 4243 18663 4277
rect 18765 4243 18769 4277
rect 18833 4243 18841 4277
rect 18901 4243 18913 4277
rect 18969 4243 18985 4277
rect 19037 4243 19057 4277
rect 19105 4243 19129 4277
rect 19173 4243 19201 4277
rect 19241 4243 19273 4277
rect 19309 4243 19343 4277
rect 19379 4243 19411 4277
rect 19451 4243 19479 4277
rect 19523 4243 19547 4277
rect 19595 4243 19615 4277
rect 19667 4243 19683 4277
rect 19739 4243 19751 4277
rect 19811 4243 19819 4277
rect 19883 4243 19887 4277
rect 19989 4243 19993 4277
rect 20057 4243 20065 4277
rect 20125 4243 20137 4277
rect 20193 4243 20209 4277
rect 20261 4243 20281 4277
rect 20329 4243 20353 4277
rect 20397 4243 20425 4277
rect 20465 4243 20497 4277
rect 20533 4243 20567 4277
rect 20603 4243 20635 4277
rect 20675 4243 20703 4277
rect 20747 4243 20771 4277
rect 20819 4243 20839 4277
rect 20891 4243 20907 4277
rect 20963 4243 20975 4277
rect 21035 4243 21043 4277
rect 21107 4243 21111 4277
rect 21213 4243 21217 4277
rect 21281 4243 21289 4277
rect 21349 4243 21361 4277
rect 21417 4243 21433 4277
rect 21485 4243 21505 4277
rect 21553 4243 21577 4277
rect 21621 4243 21649 4277
rect 21689 4243 21721 4277
rect 21757 4243 21791 4277
rect 21827 4243 21859 4277
rect 21899 4243 21927 4277
rect 21971 4243 21995 4277
rect 22043 4243 22063 4277
rect 22115 4243 22131 4277
rect 22187 4243 22199 4277
rect 22259 4243 22267 4277
rect 22331 4243 22335 4277
rect 22437 4243 22441 4277
rect 22505 4243 22513 4277
rect 22573 4243 22585 4277
rect 22641 4243 22657 4277
rect 22709 4243 22729 4277
rect 22777 4243 22801 4277
rect 22845 4243 22873 4277
rect 22913 4243 22945 4277
rect 22981 4243 23015 4277
rect 23051 4243 23083 4277
rect 23123 4243 23151 4277
rect 23195 4243 23219 4277
rect 23267 4243 23287 4277
rect 23339 4243 23355 4277
rect 23411 4243 23423 4277
rect 23483 4243 23491 4277
rect 23555 4243 23559 4277
rect 23661 4243 23665 4277
rect 23729 4243 23737 4277
rect 23797 4243 23809 4277
rect 23865 4243 23881 4277
rect 23933 4243 23953 4277
rect 24001 4243 24025 4277
rect 24069 4243 24097 4277
rect 24137 4243 24169 4277
rect 24205 4243 24239 4277
rect 24275 4243 24313 4277
rect 24347 4243 24450 4277
rect 15426 4210 24450 4243
rect 15426 4141 15526 4210
rect 15426 4077 15459 4141
rect 15493 4077 15526 4141
rect 15426 4073 15526 4077
rect 15426 3971 15459 4073
rect 15493 3971 15526 4073
rect 15426 3967 15526 3971
rect 15426 3903 15459 3967
rect 15493 3903 15526 3967
rect 15426 3895 15526 3903
rect 15426 3835 15459 3895
rect 15493 3835 15526 3895
rect 15426 3823 15526 3835
rect 15426 3767 15459 3823
rect 15493 3767 15526 3823
rect 15426 3751 15526 3767
rect 15426 3699 15459 3751
rect 15493 3699 15526 3751
rect 15426 3679 15526 3699
rect 15426 3631 15459 3679
rect 15493 3631 15526 3679
rect 15426 3607 15526 3631
rect 15426 3563 15459 3607
rect 15493 3563 15526 3607
rect 15426 3535 15526 3563
rect 15426 3495 15459 3535
rect 15493 3495 15526 3535
rect 15426 3463 15526 3495
rect 15426 3427 15459 3463
rect 15493 3427 15526 3463
rect 15426 3393 15526 3427
rect 15426 3357 15459 3393
rect 15493 3357 15526 3393
rect 15426 3325 15526 3357
rect 15426 3285 15459 3325
rect 15493 3285 15526 3325
rect 15426 3257 15526 3285
rect 15426 3213 15459 3257
rect 15493 3213 15526 3257
rect 15426 3189 15526 3213
rect 15426 3141 15459 3189
rect 15493 3141 15526 3189
rect 15426 3121 15526 3141
rect 15426 3069 15459 3121
rect 15493 3069 15526 3121
rect 15426 3053 15526 3069
rect 15426 2997 15459 3053
rect 15493 2997 15526 3053
rect 15426 2985 15526 2997
rect 15426 2925 15459 2985
rect 15493 2925 15526 2985
rect 15426 2917 15526 2925
rect 15426 2853 15459 2917
rect 15493 2853 15526 2917
rect 15426 2849 15526 2853
rect 15426 2747 15459 2849
rect 15493 2747 15526 2849
rect 15426 2743 15526 2747
rect 15426 2679 15459 2743
rect 15493 2679 15526 2743
rect 15426 2610 15526 2679
rect 24350 4141 24450 4210
rect 24350 4077 24383 4141
rect 24417 4077 24450 4141
rect 24350 4073 24450 4077
rect 24350 3971 24383 4073
rect 24417 3971 24450 4073
rect 24350 3967 24450 3971
rect 24350 3903 24383 3967
rect 24417 3903 24450 3967
rect 24350 3895 24450 3903
rect 24350 3835 24383 3895
rect 24417 3835 24450 3895
rect 24350 3823 24450 3835
rect 24350 3767 24383 3823
rect 24417 3767 24450 3823
rect 24350 3751 24450 3767
rect 24350 3699 24383 3751
rect 24417 3699 24450 3751
rect 24350 3679 24450 3699
rect 24350 3631 24383 3679
rect 24417 3631 24450 3679
rect 24350 3607 24450 3631
rect 24350 3563 24383 3607
rect 24417 3563 24450 3607
rect 24350 3535 24450 3563
rect 24350 3495 24383 3535
rect 24417 3495 24450 3535
rect 24350 3463 24450 3495
rect 24350 3427 24383 3463
rect 24417 3427 24450 3463
rect 24350 3393 24450 3427
rect 24350 3357 24383 3393
rect 24417 3357 24450 3393
rect 24350 3325 24450 3357
rect 24350 3285 24383 3325
rect 24417 3285 24450 3325
rect 24350 3257 24450 3285
rect 24350 3213 24383 3257
rect 24417 3213 24450 3257
rect 24350 3189 24450 3213
rect 24350 3141 24383 3189
rect 24417 3141 24450 3189
rect 24350 3121 24450 3141
rect 24350 3069 24383 3121
rect 24417 3069 24450 3121
rect 24350 3053 24450 3069
rect 24350 2997 24383 3053
rect 24417 2997 24450 3053
rect 24350 2985 24450 2997
rect 24350 2925 24383 2985
rect 24417 2925 24450 2985
rect 24350 2917 24450 2925
rect 24350 2853 24383 2917
rect 24417 2853 24450 2917
rect 24350 2849 24450 2853
rect 24350 2747 24383 2849
rect 24417 2747 24450 2849
rect 24350 2743 24450 2747
rect 24350 2679 24383 2743
rect 24417 2679 24450 2743
rect 24350 2610 24450 2679
rect 15426 2577 24450 2610
rect 15426 2543 15529 2577
rect 15563 2543 15601 2577
rect 15637 2543 15671 2577
rect 15707 2543 15739 2577
rect 15779 2543 15807 2577
rect 15851 2543 15875 2577
rect 15923 2543 15943 2577
rect 15995 2543 16011 2577
rect 16067 2543 16079 2577
rect 16139 2543 16147 2577
rect 16211 2543 16215 2577
rect 16317 2543 16321 2577
rect 16385 2543 16393 2577
rect 16453 2543 16465 2577
rect 16521 2543 16537 2577
rect 16589 2543 16609 2577
rect 16657 2543 16681 2577
rect 16725 2543 16753 2577
rect 16793 2543 16825 2577
rect 16861 2543 16895 2577
rect 16931 2543 16963 2577
rect 17003 2543 17031 2577
rect 17075 2543 17099 2577
rect 17147 2543 17167 2577
rect 17219 2543 17235 2577
rect 17291 2543 17303 2577
rect 17363 2543 17371 2577
rect 17435 2543 17439 2577
rect 17541 2543 17545 2577
rect 17609 2543 17617 2577
rect 17677 2543 17689 2577
rect 17745 2543 17761 2577
rect 17813 2543 17833 2577
rect 17881 2543 17905 2577
rect 17949 2543 17977 2577
rect 18017 2543 18049 2577
rect 18085 2543 18119 2577
rect 18155 2543 18187 2577
rect 18227 2543 18255 2577
rect 18299 2543 18323 2577
rect 18371 2543 18391 2577
rect 18443 2543 18459 2577
rect 18515 2543 18527 2577
rect 18587 2543 18595 2577
rect 18659 2543 18663 2577
rect 18765 2543 18769 2577
rect 18833 2543 18841 2577
rect 18901 2543 18913 2577
rect 18969 2543 18985 2577
rect 19037 2543 19057 2577
rect 19105 2543 19129 2577
rect 19173 2543 19201 2577
rect 19241 2543 19273 2577
rect 19309 2543 19343 2577
rect 19379 2543 19411 2577
rect 19451 2543 19479 2577
rect 19523 2543 19547 2577
rect 19595 2543 19615 2577
rect 19667 2543 19683 2577
rect 19739 2543 19751 2577
rect 19811 2543 19819 2577
rect 19883 2543 19887 2577
rect 19989 2543 19993 2577
rect 20057 2543 20065 2577
rect 20125 2543 20137 2577
rect 20193 2543 20209 2577
rect 20261 2543 20281 2577
rect 20329 2543 20353 2577
rect 20397 2543 20425 2577
rect 20465 2543 20497 2577
rect 20533 2543 20567 2577
rect 20603 2543 20635 2577
rect 20675 2543 20703 2577
rect 20747 2543 20771 2577
rect 20819 2543 20839 2577
rect 20891 2543 20907 2577
rect 20963 2543 20975 2577
rect 21035 2543 21043 2577
rect 21107 2543 21111 2577
rect 21213 2543 21217 2577
rect 21281 2543 21289 2577
rect 21349 2543 21361 2577
rect 21417 2543 21433 2577
rect 21485 2543 21505 2577
rect 21553 2543 21577 2577
rect 21621 2543 21649 2577
rect 21689 2543 21721 2577
rect 21757 2543 21791 2577
rect 21827 2543 21859 2577
rect 21899 2543 21927 2577
rect 21971 2543 21995 2577
rect 22043 2543 22063 2577
rect 22115 2543 22131 2577
rect 22187 2543 22199 2577
rect 22259 2543 22267 2577
rect 22331 2543 22335 2577
rect 22437 2543 22441 2577
rect 22505 2543 22513 2577
rect 22573 2543 22585 2577
rect 22641 2543 22657 2577
rect 22709 2543 22729 2577
rect 22777 2543 22801 2577
rect 22845 2543 22873 2577
rect 22913 2543 22945 2577
rect 22981 2543 23015 2577
rect 23051 2543 23083 2577
rect 23123 2543 23151 2577
rect 23195 2543 23219 2577
rect 23267 2543 23287 2577
rect 23339 2543 23355 2577
rect 23411 2543 23423 2577
rect 23483 2543 23491 2577
rect 23555 2543 23559 2577
rect 23661 2543 23665 2577
rect 23729 2543 23737 2577
rect 23797 2543 23809 2577
rect 23865 2543 23881 2577
rect 23933 2543 23953 2577
rect 24001 2543 24025 2577
rect 24069 2543 24097 2577
rect 24137 2543 24169 2577
rect 24205 2543 24239 2577
rect 24275 2543 24313 2577
rect 24347 2543 24450 2577
rect 15426 2510 24450 2543
rect 26008 4277 31452 4310
rect 26008 4243 26121 4277
rect 26155 4243 26193 4277
rect 26231 4243 26265 4277
rect 26299 4243 26333 4277
rect 26371 4243 26401 4277
rect 26443 4243 26469 4277
rect 26515 4243 26537 4277
rect 26587 4243 26605 4277
rect 26659 4243 26673 4277
rect 26731 4243 26741 4277
rect 26803 4243 26809 4277
rect 26875 4243 26877 4277
rect 26911 4243 26913 4277
rect 26979 4243 26985 4277
rect 27047 4243 27057 4277
rect 27115 4243 27129 4277
rect 27183 4243 27201 4277
rect 27251 4243 27273 4277
rect 27319 4243 27345 4277
rect 27387 4243 27417 4277
rect 27455 4243 27489 4277
rect 27523 4243 27557 4277
rect 27595 4243 27625 4277
rect 27667 4243 27693 4277
rect 27739 4243 27761 4277
rect 27811 4243 27829 4277
rect 27883 4243 27897 4277
rect 27955 4243 27965 4277
rect 28027 4243 28033 4277
rect 28099 4243 28101 4277
rect 28135 4243 28137 4277
rect 28203 4243 28209 4277
rect 28271 4243 28281 4277
rect 28339 4243 28353 4277
rect 28407 4243 28425 4277
rect 28475 4243 28497 4277
rect 28543 4243 28569 4277
rect 28611 4243 28641 4277
rect 28679 4243 28713 4277
rect 28747 4243 28781 4277
rect 28819 4243 28849 4277
rect 28891 4243 28917 4277
rect 28963 4243 28985 4277
rect 29035 4243 29053 4277
rect 29107 4243 29121 4277
rect 29179 4243 29189 4277
rect 29251 4243 29257 4277
rect 29323 4243 29325 4277
rect 29359 4243 29361 4277
rect 29427 4243 29433 4277
rect 29495 4243 29505 4277
rect 29563 4243 29577 4277
rect 29631 4243 29649 4277
rect 29699 4243 29721 4277
rect 29767 4243 29793 4277
rect 29835 4243 29865 4277
rect 29903 4243 29937 4277
rect 29971 4243 30005 4277
rect 30043 4243 30073 4277
rect 30115 4243 30141 4277
rect 30187 4243 30209 4277
rect 30259 4243 30277 4277
rect 30331 4243 30345 4277
rect 30403 4243 30413 4277
rect 30475 4243 30481 4277
rect 30547 4243 30549 4277
rect 30583 4243 30585 4277
rect 30651 4243 30657 4277
rect 30719 4243 30729 4277
rect 30787 4243 30801 4277
rect 30855 4243 30873 4277
rect 30923 4243 30945 4277
rect 30991 4243 31017 4277
rect 31059 4243 31089 4277
rect 31127 4243 31161 4277
rect 31195 4243 31229 4277
rect 31267 4243 31305 4277
rect 31339 4243 31452 4277
rect 26008 4210 31452 4243
rect 26008 4135 26108 4210
rect 26008 4073 26041 4135
rect 26075 4073 26108 4135
rect 26008 4067 26108 4073
rect 26008 4001 26041 4067
rect 26075 4001 26108 4067
rect 26008 3999 26108 4001
rect 26008 3965 26041 3999
rect 26075 3965 26108 3999
rect 26008 3963 26108 3965
rect 26008 3897 26041 3963
rect 26075 3897 26108 3963
rect 26008 3891 26108 3897
rect 26008 3829 26041 3891
rect 26075 3829 26108 3891
rect 26008 3819 26108 3829
rect 26008 3761 26041 3819
rect 26075 3761 26108 3819
rect 26008 3747 26108 3761
rect 26008 3693 26041 3747
rect 26075 3693 26108 3747
rect 26008 3675 26108 3693
rect 26008 3625 26041 3675
rect 26075 3625 26108 3675
rect 26008 3603 26108 3625
rect 26008 3557 26041 3603
rect 26075 3557 26108 3603
rect 26008 3531 26108 3557
rect 26008 3489 26041 3531
rect 26075 3489 26108 3531
rect 26008 3459 26108 3489
rect 26008 3421 26041 3459
rect 26075 3421 26108 3459
rect 26008 3387 26108 3421
rect 26008 3353 26041 3387
rect 26075 3353 26108 3387
rect 26008 3319 26108 3353
rect 26008 3281 26041 3319
rect 26075 3281 26108 3319
rect 26008 3251 26108 3281
rect 26008 3209 26041 3251
rect 26075 3209 26108 3251
rect 26008 3183 26108 3209
rect 26008 3137 26041 3183
rect 26075 3137 26108 3183
rect 26008 3115 26108 3137
rect 26008 3065 26041 3115
rect 26075 3065 26108 3115
rect 26008 3047 26108 3065
rect 26008 2993 26041 3047
rect 26075 2993 26108 3047
rect 26008 2979 26108 2993
rect 26008 2921 26041 2979
rect 26075 2921 26108 2979
rect 26008 2911 26108 2921
rect 26008 2849 26041 2911
rect 26075 2849 26108 2911
rect 26008 2843 26108 2849
rect 26008 2777 26041 2843
rect 26075 2777 26108 2843
rect 26008 2775 26108 2777
rect 26008 2741 26041 2775
rect 26075 2741 26108 2775
rect 26008 2739 26108 2741
rect 26008 2673 26041 2739
rect 26075 2673 26108 2739
rect 26008 2667 26108 2673
rect 26008 2605 26041 2667
rect 26075 2605 26108 2667
rect 26008 2530 26108 2605
rect 31352 4135 31452 4210
rect 31352 4073 31385 4135
rect 31419 4073 31452 4135
rect 31352 4067 31452 4073
rect 31352 4001 31385 4067
rect 31419 4001 31452 4067
rect 31352 3999 31452 4001
rect 31352 3965 31385 3999
rect 31419 3965 31452 3999
rect 31352 3963 31452 3965
rect 31352 3897 31385 3963
rect 31419 3897 31452 3963
rect 31352 3891 31452 3897
rect 31352 3829 31385 3891
rect 31419 3829 31452 3891
rect 31352 3819 31452 3829
rect 31352 3761 31385 3819
rect 31419 3761 31452 3819
rect 31352 3747 31452 3761
rect 31352 3693 31385 3747
rect 31419 3693 31452 3747
rect 31352 3675 31452 3693
rect 31352 3625 31385 3675
rect 31419 3625 31452 3675
rect 31352 3603 31452 3625
rect 31352 3557 31385 3603
rect 31419 3557 31452 3603
rect 31352 3531 31452 3557
rect 31352 3489 31385 3531
rect 31419 3489 31452 3531
rect 31352 3459 31452 3489
rect 31352 3421 31385 3459
rect 31419 3421 31452 3459
rect 31352 3387 31452 3421
rect 31352 3353 31385 3387
rect 31419 3353 31452 3387
rect 31352 3319 31452 3353
rect 31352 3281 31385 3319
rect 31419 3281 31452 3319
rect 31352 3251 31452 3281
rect 31352 3209 31385 3251
rect 31419 3209 31452 3251
rect 31352 3183 31452 3209
rect 31352 3137 31385 3183
rect 31419 3137 31452 3183
rect 31352 3115 31452 3137
rect 31352 3065 31385 3115
rect 31419 3065 31452 3115
rect 31352 3047 31452 3065
rect 31352 2993 31385 3047
rect 31419 2993 31452 3047
rect 31352 2979 31452 2993
rect 31352 2921 31385 2979
rect 31419 2921 31452 2979
rect 31352 2911 31452 2921
rect 31352 2849 31385 2911
rect 31419 2849 31452 2911
rect 31352 2843 31452 2849
rect 31352 2777 31385 2843
rect 31419 2777 31452 2843
rect 31352 2775 31452 2777
rect 31352 2741 31385 2775
rect 31419 2741 31452 2775
rect 31352 2739 31452 2741
rect 31352 2673 31385 2739
rect 31419 2673 31452 2739
rect 31352 2667 31452 2673
rect 31352 2605 31385 2667
rect 31419 2605 31452 2667
rect 31352 2530 31452 2605
rect 26008 2497 31452 2530
rect 26008 2463 26121 2497
rect 26155 2463 26193 2497
rect 26231 2463 26265 2497
rect 26299 2463 26333 2497
rect 26371 2463 26401 2497
rect 26443 2463 26469 2497
rect 26515 2463 26537 2497
rect 26587 2463 26605 2497
rect 26659 2463 26673 2497
rect 26731 2463 26741 2497
rect 26803 2463 26809 2497
rect 26875 2463 26877 2497
rect 26911 2463 26913 2497
rect 26979 2463 26985 2497
rect 27047 2463 27057 2497
rect 27115 2463 27129 2497
rect 27183 2463 27201 2497
rect 27251 2463 27273 2497
rect 27319 2463 27345 2497
rect 27387 2463 27417 2497
rect 27455 2463 27489 2497
rect 27523 2463 27557 2497
rect 27595 2463 27625 2497
rect 27667 2463 27693 2497
rect 27739 2463 27761 2497
rect 27811 2463 27829 2497
rect 27883 2463 27897 2497
rect 27955 2463 27965 2497
rect 28027 2463 28033 2497
rect 28099 2463 28101 2497
rect 28135 2463 28137 2497
rect 28203 2463 28209 2497
rect 28271 2463 28281 2497
rect 28339 2463 28353 2497
rect 28407 2463 28425 2497
rect 28475 2463 28497 2497
rect 28543 2463 28569 2497
rect 28611 2463 28641 2497
rect 28679 2463 28713 2497
rect 28747 2463 28781 2497
rect 28819 2463 28849 2497
rect 28891 2463 28917 2497
rect 28963 2463 28985 2497
rect 29035 2463 29053 2497
rect 29107 2463 29121 2497
rect 29179 2463 29189 2497
rect 29251 2463 29257 2497
rect 29323 2463 29325 2497
rect 29359 2463 29361 2497
rect 29427 2463 29433 2497
rect 29495 2463 29505 2497
rect 29563 2463 29577 2497
rect 29631 2463 29649 2497
rect 29699 2463 29721 2497
rect 29767 2463 29793 2497
rect 29835 2463 29865 2497
rect 29903 2463 29937 2497
rect 29971 2463 30005 2497
rect 30043 2463 30073 2497
rect 30115 2463 30141 2497
rect 30187 2463 30209 2497
rect 30259 2463 30277 2497
rect 30331 2463 30345 2497
rect 30403 2463 30413 2497
rect 30475 2463 30481 2497
rect 30547 2463 30549 2497
rect 30583 2463 30585 2497
rect 30651 2463 30657 2497
rect 30719 2463 30729 2497
rect 30787 2463 30801 2497
rect 30855 2463 30873 2497
rect 30923 2463 30945 2497
rect 30991 2463 31017 2497
rect 31059 2463 31089 2497
rect 31127 2463 31161 2497
rect 31195 2463 31229 2497
rect 31267 2463 31305 2497
rect 31339 2463 31452 2497
rect 26008 2430 31452 2463
rect 15426 2241 24450 2274
rect 15426 2207 15529 2241
rect 15563 2207 15601 2241
rect 15637 2207 15671 2241
rect 15707 2207 15739 2241
rect 15779 2207 15807 2241
rect 15851 2207 15875 2241
rect 15923 2207 15943 2241
rect 15995 2207 16011 2241
rect 16067 2207 16079 2241
rect 16139 2207 16147 2241
rect 16211 2207 16215 2241
rect 16317 2207 16321 2241
rect 16385 2207 16393 2241
rect 16453 2207 16465 2241
rect 16521 2207 16537 2241
rect 16589 2207 16609 2241
rect 16657 2207 16681 2241
rect 16725 2207 16753 2241
rect 16793 2207 16825 2241
rect 16861 2207 16895 2241
rect 16931 2207 16963 2241
rect 17003 2207 17031 2241
rect 17075 2207 17099 2241
rect 17147 2207 17167 2241
rect 17219 2207 17235 2241
rect 17291 2207 17303 2241
rect 17363 2207 17371 2241
rect 17435 2207 17439 2241
rect 17541 2207 17545 2241
rect 17609 2207 17617 2241
rect 17677 2207 17689 2241
rect 17745 2207 17761 2241
rect 17813 2207 17833 2241
rect 17881 2207 17905 2241
rect 17949 2207 17977 2241
rect 18017 2207 18049 2241
rect 18085 2207 18119 2241
rect 18155 2207 18187 2241
rect 18227 2207 18255 2241
rect 18299 2207 18323 2241
rect 18371 2207 18391 2241
rect 18443 2207 18459 2241
rect 18515 2207 18527 2241
rect 18587 2207 18595 2241
rect 18659 2207 18663 2241
rect 18765 2207 18769 2241
rect 18833 2207 18841 2241
rect 18901 2207 18913 2241
rect 18969 2207 18985 2241
rect 19037 2207 19057 2241
rect 19105 2207 19129 2241
rect 19173 2207 19201 2241
rect 19241 2207 19273 2241
rect 19309 2207 19343 2241
rect 19379 2207 19411 2241
rect 19451 2207 19479 2241
rect 19523 2207 19547 2241
rect 19595 2207 19615 2241
rect 19667 2207 19683 2241
rect 19739 2207 19751 2241
rect 19811 2207 19819 2241
rect 19883 2207 19887 2241
rect 19989 2207 19993 2241
rect 20057 2207 20065 2241
rect 20125 2207 20137 2241
rect 20193 2207 20209 2241
rect 20261 2207 20281 2241
rect 20329 2207 20353 2241
rect 20397 2207 20425 2241
rect 20465 2207 20497 2241
rect 20533 2207 20567 2241
rect 20603 2207 20635 2241
rect 20675 2207 20703 2241
rect 20747 2207 20771 2241
rect 20819 2207 20839 2241
rect 20891 2207 20907 2241
rect 20963 2207 20975 2241
rect 21035 2207 21043 2241
rect 21107 2207 21111 2241
rect 21213 2207 21217 2241
rect 21281 2207 21289 2241
rect 21349 2207 21361 2241
rect 21417 2207 21433 2241
rect 21485 2207 21505 2241
rect 21553 2207 21577 2241
rect 21621 2207 21649 2241
rect 21689 2207 21721 2241
rect 21757 2207 21791 2241
rect 21827 2207 21859 2241
rect 21899 2207 21927 2241
rect 21971 2207 21995 2241
rect 22043 2207 22063 2241
rect 22115 2207 22131 2241
rect 22187 2207 22199 2241
rect 22259 2207 22267 2241
rect 22331 2207 22335 2241
rect 22437 2207 22441 2241
rect 22505 2207 22513 2241
rect 22573 2207 22585 2241
rect 22641 2207 22657 2241
rect 22709 2207 22729 2241
rect 22777 2207 22801 2241
rect 22845 2207 22873 2241
rect 22913 2207 22945 2241
rect 22981 2207 23015 2241
rect 23051 2207 23083 2241
rect 23123 2207 23151 2241
rect 23195 2207 23219 2241
rect 23267 2207 23287 2241
rect 23339 2207 23355 2241
rect 23411 2207 23423 2241
rect 23483 2207 23491 2241
rect 23555 2207 23559 2241
rect 23661 2207 23665 2241
rect 23729 2207 23737 2241
rect 23797 2207 23809 2241
rect 23865 2207 23881 2241
rect 23933 2207 23953 2241
rect 24001 2207 24025 2241
rect 24069 2207 24097 2241
rect 24137 2207 24169 2241
rect 24205 2207 24239 2241
rect 24275 2207 24313 2241
rect 24347 2207 24450 2241
rect 31606 2267 31654 2274
rect 31606 2233 31613 2267
rect 31647 2233 31654 2267
rect 31606 2226 31654 2233
rect 31712 2269 31760 2276
rect 31712 2235 31719 2269
rect 31753 2235 31760 2269
rect 31712 2228 31760 2235
rect 31848 2269 31896 2276
rect 31848 2235 31855 2269
rect 31889 2235 31896 2269
rect 31848 2228 31896 2235
rect 32204 2269 32252 2276
rect 32204 2235 32211 2269
rect 32245 2235 32252 2269
rect 32204 2228 32252 2235
rect 15426 2174 24450 2207
rect 15426 2093 15526 2174
rect 15426 2059 15459 2093
rect 15493 2059 15526 2093
rect 15426 2025 15526 2059
rect 15426 1991 15459 2025
rect 15493 1991 15526 2025
rect 15426 1957 15526 1991
rect 15426 1911 15459 1957
rect 15493 1911 15526 1957
rect 15426 1889 15526 1911
rect 15426 1839 15459 1889
rect 15493 1839 15526 1889
rect 15426 1821 15526 1839
rect 15426 1767 15459 1821
rect 15493 1767 15526 1821
rect 15426 1753 15526 1767
rect 15426 1695 15459 1753
rect 15493 1695 15526 1753
rect 15426 1685 15526 1695
rect 15426 1623 15459 1685
rect 15493 1623 15526 1685
rect 15426 1617 15526 1623
rect 15426 1551 15459 1617
rect 15493 1551 15526 1617
rect 15426 1549 15526 1551
rect 15426 1515 15459 1549
rect 15493 1515 15526 1549
rect 15426 1513 15526 1515
rect 15426 1447 15459 1513
rect 15493 1447 15526 1513
rect 15426 1441 15526 1447
rect 15426 1379 15459 1441
rect 15493 1379 15526 1441
rect 15426 1369 15526 1379
rect 15426 1311 15459 1369
rect 15493 1311 15526 1369
rect 15426 1297 15526 1311
rect 15426 1243 15459 1297
rect 15493 1243 15526 1297
rect 15426 1225 15526 1243
rect 15426 1175 15459 1225
rect 15493 1175 15526 1225
rect 15426 1153 15526 1175
rect 15426 1107 15459 1153
rect 15493 1107 15526 1153
rect 15426 1081 15526 1107
rect 15426 1039 15459 1081
rect 15493 1039 15526 1081
rect 15426 1009 15526 1039
rect 15426 971 15459 1009
rect 15493 971 15526 1009
rect 15426 937 15526 971
rect 15426 903 15459 937
rect 15493 903 15526 937
rect 15426 869 15526 903
rect 15426 831 15459 869
rect 15493 831 15526 869
rect 15426 801 15526 831
rect 15426 759 15459 801
rect 15493 759 15526 801
rect 15426 733 15526 759
rect 15426 687 15459 733
rect 15493 687 15526 733
rect 15426 665 15526 687
rect 15426 615 15459 665
rect 15493 615 15526 665
rect 15426 597 15526 615
rect 15426 543 15459 597
rect 15493 543 15526 597
rect 15426 529 15526 543
rect 15426 471 15459 529
rect 15493 471 15526 529
rect 15426 461 15526 471
rect 15426 399 15459 461
rect 15493 399 15526 461
rect 15426 393 15526 399
rect 15426 327 15459 393
rect 15493 327 15526 393
rect 15426 325 15526 327
rect 15426 291 15459 325
rect 15493 291 15526 325
rect 15426 289 15526 291
rect 15426 223 15459 289
rect 15493 223 15526 289
rect 15426 217 15526 223
rect 15426 155 15459 217
rect 15493 155 15526 217
rect 15426 145 15526 155
rect 15426 87 15459 145
rect 15493 87 15526 145
rect 15426 73 15526 87
rect 15426 19 15459 73
rect 15493 19 15526 73
rect 15426 1 15526 19
rect 15426 -49 15459 1
rect 15493 -49 15526 1
rect 15426 -71 15526 -49
rect 15426 -117 15459 -71
rect 15493 -117 15526 -71
rect 15426 -143 15526 -117
rect 15426 -185 15459 -143
rect 15493 -185 15526 -143
rect 15426 -215 15526 -185
rect 15426 -253 15459 -215
rect 15493 -253 15526 -215
rect 15426 -287 15526 -253
rect 15426 -321 15459 -287
rect 15493 -321 15526 -287
rect 15426 -355 15526 -321
rect 15426 -393 15459 -355
rect 15493 -393 15526 -355
rect 15426 -423 15526 -393
rect 15426 -465 15459 -423
rect 15493 -465 15526 -423
rect 15426 -491 15526 -465
rect 15426 -537 15459 -491
rect 15493 -537 15526 -491
rect 15426 -559 15526 -537
rect 15426 -609 15459 -559
rect 15493 -609 15526 -559
rect 15426 -627 15526 -609
rect 15426 -681 15459 -627
rect 15493 -681 15526 -627
rect 15426 -695 15526 -681
rect 15426 -753 15459 -695
rect 15493 -753 15526 -695
rect 15426 -763 15526 -753
rect 15426 -825 15459 -763
rect 15493 -825 15526 -763
rect 15426 -831 15526 -825
rect 15426 -897 15459 -831
rect 15493 -897 15526 -831
rect 15426 -899 15526 -897
rect 15426 -933 15459 -899
rect 15493 -933 15526 -899
rect 15426 -935 15526 -933
rect 15426 -1001 15459 -935
rect 15493 -1001 15526 -935
rect 15426 -1007 15526 -1001
rect 15426 -1069 15459 -1007
rect 15493 -1069 15526 -1007
rect 15426 -1079 15526 -1069
rect 15426 -1137 15459 -1079
rect 15493 -1137 15526 -1079
rect 15426 -1151 15526 -1137
rect 15426 -1205 15459 -1151
rect 15493 -1205 15526 -1151
rect 15426 -1223 15526 -1205
rect 15426 -1273 15459 -1223
rect 15493 -1273 15526 -1223
rect 15426 -1295 15526 -1273
rect 15426 -1341 15459 -1295
rect 15493 -1341 15526 -1295
rect 15426 -1375 15526 -1341
rect 15426 -1409 15459 -1375
rect 15493 -1409 15526 -1375
rect 15426 -1443 15526 -1409
rect 15426 -1477 15459 -1443
rect 15493 -1477 15526 -1443
rect 15426 -1558 15526 -1477
rect 24350 2093 24450 2174
rect 24350 2059 24383 2093
rect 24417 2059 24450 2093
rect 24350 2025 24450 2059
rect 24350 1991 24383 2025
rect 24417 1991 24450 2025
rect 24350 1957 24450 1991
rect 24350 1911 24383 1957
rect 24417 1911 24450 1957
rect 24350 1889 24450 1911
rect 24350 1839 24383 1889
rect 24417 1839 24450 1889
rect 24350 1821 24450 1839
rect 24350 1767 24383 1821
rect 24417 1767 24450 1821
rect 24350 1753 24450 1767
rect 24350 1695 24383 1753
rect 24417 1695 24450 1753
rect 24350 1685 24450 1695
rect 24350 1623 24383 1685
rect 24417 1623 24450 1685
rect 24350 1617 24450 1623
rect 24350 1551 24383 1617
rect 24417 1551 24450 1617
rect 24350 1549 24450 1551
rect 24350 1515 24383 1549
rect 24417 1515 24450 1549
rect 24350 1513 24450 1515
rect 24350 1447 24383 1513
rect 24417 1447 24450 1513
rect 24350 1441 24450 1447
rect 24350 1379 24383 1441
rect 24417 1379 24450 1441
rect 24350 1369 24450 1379
rect 24350 1311 24383 1369
rect 24417 1311 24450 1369
rect 24350 1297 24450 1311
rect 24350 1243 24383 1297
rect 24417 1243 24450 1297
rect 24350 1225 24450 1243
rect 24350 1175 24383 1225
rect 24417 1175 24450 1225
rect 24350 1153 24450 1175
rect 24350 1107 24383 1153
rect 24417 1107 24450 1153
rect 24350 1081 24450 1107
rect 24350 1039 24383 1081
rect 24417 1039 24450 1081
rect 24350 1009 24450 1039
rect 24350 971 24383 1009
rect 24417 971 24450 1009
rect 24350 937 24450 971
rect 24350 903 24383 937
rect 24417 903 24450 937
rect 24350 869 24450 903
rect 24350 831 24383 869
rect 24417 831 24450 869
rect 24350 801 24450 831
rect 24350 759 24383 801
rect 24417 759 24450 801
rect 24350 733 24450 759
rect 24350 687 24383 733
rect 24417 687 24450 733
rect 24350 665 24450 687
rect 24350 615 24383 665
rect 24417 615 24450 665
rect 24350 597 24450 615
rect 24350 543 24383 597
rect 24417 543 24450 597
rect 24350 529 24450 543
rect 24350 471 24383 529
rect 24417 471 24450 529
rect 24350 461 24450 471
rect 24350 399 24383 461
rect 24417 399 24450 461
rect 24350 393 24450 399
rect 24350 327 24383 393
rect 24417 327 24450 393
rect 24350 325 24450 327
rect 24350 291 24383 325
rect 24417 291 24450 325
rect 24350 289 24450 291
rect 24350 223 24383 289
rect 24417 223 24450 289
rect 24350 217 24450 223
rect 24350 155 24383 217
rect 24417 155 24450 217
rect 24350 145 24450 155
rect 24350 87 24383 145
rect 24417 87 24450 145
rect 24350 73 24450 87
rect 24350 19 24383 73
rect 24417 19 24450 73
rect 24350 1 24450 19
rect 24350 -49 24383 1
rect 24417 -49 24450 1
rect 24350 -71 24450 -49
rect 24350 -117 24383 -71
rect 24417 -117 24450 -71
rect 24350 -143 24450 -117
rect 24350 -185 24383 -143
rect 24417 -185 24450 -143
rect 24350 -215 24450 -185
rect 24350 -253 24383 -215
rect 24417 -253 24450 -215
rect 24350 -287 24450 -253
rect 24350 -321 24383 -287
rect 24417 -321 24450 -287
rect 24350 -355 24450 -321
rect 24350 -393 24383 -355
rect 24417 -393 24450 -355
rect 24350 -423 24450 -393
rect 24350 -465 24383 -423
rect 24417 -465 24450 -423
rect 24350 -491 24450 -465
rect 24350 -537 24383 -491
rect 24417 -537 24450 -491
rect 24350 -559 24450 -537
rect 24350 -609 24383 -559
rect 24417 -609 24450 -559
rect 24350 -627 24450 -609
rect 24350 -681 24383 -627
rect 24417 -681 24450 -627
rect 24350 -695 24450 -681
rect 24350 -753 24383 -695
rect 24417 -753 24450 -695
rect 24350 -763 24450 -753
rect 24350 -825 24383 -763
rect 24417 -825 24450 -763
rect 24350 -831 24450 -825
rect 24350 -897 24383 -831
rect 24417 -897 24450 -831
rect 24350 -899 24450 -897
rect 24350 -933 24383 -899
rect 24417 -933 24450 -899
rect 24350 -935 24450 -933
rect 24350 -1001 24383 -935
rect 24417 -1001 24450 -935
rect 24350 -1007 24450 -1001
rect 24350 -1069 24383 -1007
rect 24417 -1069 24450 -1007
rect 24350 -1079 24450 -1069
rect 24350 -1137 24383 -1079
rect 24417 -1137 24450 -1079
rect 24350 -1151 24450 -1137
rect 24350 -1205 24383 -1151
rect 24417 -1205 24450 -1151
rect 24350 -1223 24450 -1205
rect 24350 -1273 24383 -1223
rect 24417 -1273 24450 -1223
rect 24350 -1295 24450 -1273
rect 24350 -1341 24383 -1295
rect 24417 -1341 24450 -1295
rect 24350 -1375 24450 -1341
rect 24350 -1409 24383 -1375
rect 24417 -1409 24450 -1375
rect 24350 -1443 24450 -1409
rect 24350 -1477 24383 -1443
rect 24417 -1477 24450 -1443
rect 24350 -1558 24450 -1477
rect 15426 -1591 24450 -1558
rect 15426 -1625 15529 -1591
rect 15563 -1625 15601 -1591
rect 15637 -1625 15671 -1591
rect 15707 -1625 15739 -1591
rect 15779 -1625 15807 -1591
rect 15851 -1625 15875 -1591
rect 15923 -1625 15943 -1591
rect 15995 -1625 16011 -1591
rect 16067 -1625 16079 -1591
rect 16139 -1625 16147 -1591
rect 16211 -1625 16215 -1591
rect 16317 -1625 16321 -1591
rect 16385 -1625 16393 -1591
rect 16453 -1625 16465 -1591
rect 16521 -1625 16537 -1591
rect 16589 -1625 16609 -1591
rect 16657 -1625 16681 -1591
rect 16725 -1625 16753 -1591
rect 16793 -1625 16825 -1591
rect 16861 -1625 16895 -1591
rect 16931 -1625 16963 -1591
rect 17003 -1625 17031 -1591
rect 17075 -1625 17099 -1591
rect 17147 -1625 17167 -1591
rect 17219 -1625 17235 -1591
rect 17291 -1625 17303 -1591
rect 17363 -1625 17371 -1591
rect 17435 -1625 17439 -1591
rect 17541 -1625 17545 -1591
rect 17609 -1625 17617 -1591
rect 17677 -1625 17689 -1591
rect 17745 -1625 17761 -1591
rect 17813 -1625 17833 -1591
rect 17881 -1625 17905 -1591
rect 17949 -1625 17977 -1591
rect 18017 -1625 18049 -1591
rect 18085 -1625 18119 -1591
rect 18155 -1625 18187 -1591
rect 18227 -1625 18255 -1591
rect 18299 -1625 18323 -1591
rect 18371 -1625 18391 -1591
rect 18443 -1625 18459 -1591
rect 18515 -1625 18527 -1591
rect 18587 -1625 18595 -1591
rect 18659 -1625 18663 -1591
rect 18765 -1625 18769 -1591
rect 18833 -1625 18841 -1591
rect 18901 -1625 18913 -1591
rect 18969 -1625 18985 -1591
rect 19037 -1625 19057 -1591
rect 19105 -1625 19129 -1591
rect 19173 -1625 19201 -1591
rect 19241 -1625 19273 -1591
rect 19309 -1625 19343 -1591
rect 19379 -1625 19411 -1591
rect 19451 -1625 19479 -1591
rect 19523 -1625 19547 -1591
rect 19595 -1625 19615 -1591
rect 19667 -1625 19683 -1591
rect 19739 -1625 19751 -1591
rect 19811 -1625 19819 -1591
rect 19883 -1625 19887 -1591
rect 19989 -1625 19993 -1591
rect 20057 -1625 20065 -1591
rect 20125 -1625 20137 -1591
rect 20193 -1625 20209 -1591
rect 20261 -1625 20281 -1591
rect 20329 -1625 20353 -1591
rect 20397 -1625 20425 -1591
rect 20465 -1625 20497 -1591
rect 20533 -1625 20567 -1591
rect 20603 -1625 20635 -1591
rect 20675 -1625 20703 -1591
rect 20747 -1625 20771 -1591
rect 20819 -1625 20839 -1591
rect 20891 -1625 20907 -1591
rect 20963 -1625 20975 -1591
rect 21035 -1625 21043 -1591
rect 21107 -1625 21111 -1591
rect 21213 -1625 21217 -1591
rect 21281 -1625 21289 -1591
rect 21349 -1625 21361 -1591
rect 21417 -1625 21433 -1591
rect 21485 -1625 21505 -1591
rect 21553 -1625 21577 -1591
rect 21621 -1625 21649 -1591
rect 21689 -1625 21721 -1591
rect 21757 -1625 21791 -1591
rect 21827 -1625 21859 -1591
rect 21899 -1625 21927 -1591
rect 21971 -1625 21995 -1591
rect 22043 -1625 22063 -1591
rect 22115 -1625 22131 -1591
rect 22187 -1625 22199 -1591
rect 22259 -1625 22267 -1591
rect 22331 -1625 22335 -1591
rect 22437 -1625 22441 -1591
rect 22505 -1625 22513 -1591
rect 22573 -1625 22585 -1591
rect 22641 -1625 22657 -1591
rect 22709 -1625 22729 -1591
rect 22777 -1625 22801 -1591
rect 22845 -1625 22873 -1591
rect 22913 -1625 22945 -1591
rect 22981 -1625 23015 -1591
rect 23051 -1625 23083 -1591
rect 23123 -1625 23151 -1591
rect 23195 -1625 23219 -1591
rect 23267 -1625 23287 -1591
rect 23339 -1625 23355 -1591
rect 23411 -1625 23423 -1591
rect 23483 -1625 23491 -1591
rect 23555 -1625 23559 -1591
rect 23661 -1625 23665 -1591
rect 23729 -1625 23737 -1591
rect 23797 -1625 23809 -1591
rect 23865 -1625 23881 -1591
rect 23933 -1625 23953 -1591
rect 24001 -1625 24025 -1591
rect 24069 -1625 24097 -1591
rect 24137 -1625 24169 -1591
rect 24205 -1625 24239 -1591
rect 24275 -1625 24313 -1591
rect 24347 -1625 24450 -1591
rect 15426 -1658 24450 -1625
rect 26008 2161 31452 2194
rect 26008 2127 26121 2161
rect 26155 2127 26193 2161
rect 26231 2127 26265 2161
rect 26299 2127 26333 2161
rect 26371 2127 26401 2161
rect 26443 2127 26469 2161
rect 26515 2127 26537 2161
rect 26587 2127 26605 2161
rect 26659 2127 26673 2161
rect 26731 2127 26741 2161
rect 26803 2127 26809 2161
rect 26875 2127 26877 2161
rect 26911 2127 26913 2161
rect 26979 2127 26985 2161
rect 27047 2127 27057 2161
rect 27115 2127 27129 2161
rect 27183 2127 27201 2161
rect 27251 2127 27273 2161
rect 27319 2127 27345 2161
rect 27387 2127 27417 2161
rect 27455 2127 27489 2161
rect 27523 2127 27557 2161
rect 27595 2127 27625 2161
rect 27667 2127 27693 2161
rect 27739 2127 27761 2161
rect 27811 2127 27829 2161
rect 27883 2127 27897 2161
rect 27955 2127 27965 2161
rect 28027 2127 28033 2161
rect 28099 2127 28101 2161
rect 28135 2127 28137 2161
rect 28203 2127 28209 2161
rect 28271 2127 28281 2161
rect 28339 2127 28353 2161
rect 28407 2127 28425 2161
rect 28475 2127 28497 2161
rect 28543 2127 28569 2161
rect 28611 2127 28641 2161
rect 28679 2127 28713 2161
rect 28747 2127 28781 2161
rect 28819 2127 28849 2161
rect 28891 2127 28917 2161
rect 28963 2127 28985 2161
rect 29035 2127 29053 2161
rect 29107 2127 29121 2161
rect 29179 2127 29189 2161
rect 29251 2127 29257 2161
rect 29323 2127 29325 2161
rect 29359 2127 29361 2161
rect 29427 2127 29433 2161
rect 29495 2127 29505 2161
rect 29563 2127 29577 2161
rect 29631 2127 29649 2161
rect 29699 2127 29721 2161
rect 29767 2127 29793 2161
rect 29835 2127 29865 2161
rect 29903 2127 29937 2161
rect 29971 2127 30005 2161
rect 30043 2127 30073 2161
rect 30115 2127 30141 2161
rect 30187 2127 30209 2161
rect 30259 2127 30277 2161
rect 30331 2127 30345 2161
rect 30403 2127 30413 2161
rect 30475 2127 30481 2161
rect 30547 2127 30549 2161
rect 30583 2127 30585 2161
rect 30651 2127 30657 2161
rect 30719 2127 30729 2161
rect 30787 2127 30801 2161
rect 30855 2127 30873 2161
rect 30923 2127 30945 2161
rect 30991 2127 31017 2161
rect 31059 2127 31089 2161
rect 31127 2127 31161 2161
rect 31195 2127 31229 2161
rect 31267 2127 31305 2161
rect 31339 2127 31452 2161
rect 26008 2094 31452 2127
rect 26008 2019 26108 2094
rect 26008 1985 26041 2019
rect 26075 1985 26108 2019
rect 26008 1951 26108 1985
rect 26008 1917 26041 1951
rect 26075 1917 26108 1951
rect 26008 1905 26108 1917
rect 26008 1849 26041 1905
rect 26075 1849 26108 1905
rect 26008 1833 26108 1849
rect 26008 1781 26041 1833
rect 26075 1781 26108 1833
rect 26008 1761 26108 1781
rect 26008 1713 26041 1761
rect 26075 1713 26108 1761
rect 26008 1689 26108 1713
rect 26008 1645 26041 1689
rect 26075 1645 26108 1689
rect 26008 1617 26108 1645
rect 26008 1577 26041 1617
rect 26075 1577 26108 1617
rect 26008 1545 26108 1577
rect 26008 1509 26041 1545
rect 26075 1509 26108 1545
rect 26008 1475 26108 1509
rect 26008 1439 26041 1475
rect 26075 1439 26108 1475
rect 26008 1407 26108 1439
rect 26008 1367 26041 1407
rect 26075 1367 26108 1407
rect 26008 1339 26108 1367
rect 26008 1295 26041 1339
rect 26075 1295 26108 1339
rect 26008 1271 26108 1295
rect 26008 1223 26041 1271
rect 26075 1223 26108 1271
rect 26008 1203 26108 1223
rect 26008 1151 26041 1203
rect 26075 1151 26108 1203
rect 26008 1135 26108 1151
rect 26008 1079 26041 1135
rect 26075 1079 26108 1135
rect 26008 1067 26108 1079
rect 26008 1007 26041 1067
rect 26075 1007 26108 1067
rect 26008 999 26108 1007
rect 26008 935 26041 999
rect 26075 935 26108 999
rect 26008 931 26108 935
rect 26008 829 26041 931
rect 26075 829 26108 931
rect 26008 825 26108 829
rect 26008 761 26041 825
rect 26075 761 26108 825
rect 26008 753 26108 761
rect 26008 693 26041 753
rect 26075 693 26108 753
rect 26008 681 26108 693
rect 26008 625 26041 681
rect 26075 625 26108 681
rect 26008 609 26108 625
rect 26008 557 26041 609
rect 26075 557 26108 609
rect 26008 537 26108 557
rect 26008 489 26041 537
rect 26075 489 26108 537
rect 26008 465 26108 489
rect 26008 421 26041 465
rect 26075 421 26108 465
rect 26008 393 26108 421
rect 26008 353 26041 393
rect 26075 353 26108 393
rect 26008 321 26108 353
rect 26008 285 26041 321
rect 26075 285 26108 321
rect 26008 251 26108 285
rect 26008 215 26041 251
rect 26075 215 26108 251
rect 26008 183 26108 215
rect 26008 143 26041 183
rect 26075 143 26108 183
rect 26008 115 26108 143
rect 26008 71 26041 115
rect 26075 71 26108 115
rect 26008 47 26108 71
rect 26008 -1 26041 47
rect 26075 -1 26108 47
rect 26008 -21 26108 -1
rect 26008 -73 26041 -21
rect 26075 -73 26108 -21
rect 26008 -89 26108 -73
rect 26008 -145 26041 -89
rect 26075 -145 26108 -89
rect 26008 -157 26108 -145
rect 26008 -217 26041 -157
rect 26075 -217 26108 -157
rect 26008 -225 26108 -217
rect 26008 -289 26041 -225
rect 26075 -289 26108 -225
rect 26008 -293 26108 -289
rect 26008 -395 26041 -293
rect 26075 -395 26108 -293
rect 26008 -399 26108 -395
rect 26008 -463 26041 -399
rect 26075 -463 26108 -399
rect 26008 -471 26108 -463
rect 26008 -531 26041 -471
rect 26075 -531 26108 -471
rect 26008 -543 26108 -531
rect 26008 -599 26041 -543
rect 26075 -599 26108 -543
rect 26008 -615 26108 -599
rect 26008 -667 26041 -615
rect 26075 -667 26108 -615
rect 26008 -687 26108 -667
rect 26008 -735 26041 -687
rect 26075 -735 26108 -687
rect 26008 -759 26108 -735
rect 26008 -803 26041 -759
rect 26075 -803 26108 -759
rect 26008 -831 26108 -803
rect 26008 -871 26041 -831
rect 26075 -871 26108 -831
rect 26008 -903 26108 -871
rect 26008 -939 26041 -903
rect 26075 -939 26108 -903
rect 26008 -973 26108 -939
rect 26008 -1009 26041 -973
rect 26075 -1009 26108 -973
rect 26008 -1041 26108 -1009
rect 26008 -1081 26041 -1041
rect 26075 -1081 26108 -1041
rect 26008 -1109 26108 -1081
rect 26008 -1153 26041 -1109
rect 26075 -1153 26108 -1109
rect 26008 -1177 26108 -1153
rect 26008 -1225 26041 -1177
rect 26075 -1225 26108 -1177
rect 26008 -1245 26108 -1225
rect 26008 -1297 26041 -1245
rect 26075 -1297 26108 -1245
rect 26008 -1313 26108 -1297
rect 26008 -1369 26041 -1313
rect 26075 -1369 26108 -1313
rect 26008 -1381 26108 -1369
rect 26008 -1415 26041 -1381
rect 26075 -1415 26108 -1381
rect 26008 -1449 26108 -1415
rect 26008 -1483 26041 -1449
rect 26075 -1483 26108 -1449
rect 26008 -1558 26108 -1483
rect 31352 2019 31452 2094
rect 31352 1985 31385 2019
rect 31419 1985 31452 2019
rect 31352 1951 31452 1985
rect 31352 1917 31385 1951
rect 31419 1917 31452 1951
rect 31352 1905 31452 1917
rect 31352 1849 31385 1905
rect 31419 1849 31452 1905
rect 31352 1833 31452 1849
rect 31352 1781 31385 1833
rect 31419 1781 31452 1833
rect 31352 1761 31452 1781
rect 31352 1713 31385 1761
rect 31419 1713 31452 1761
rect 31352 1689 31452 1713
rect 31352 1645 31385 1689
rect 31419 1645 31452 1689
rect 31352 1617 31452 1645
rect 31352 1577 31385 1617
rect 31419 1577 31452 1617
rect 31352 1545 31452 1577
rect 31352 1509 31385 1545
rect 31419 1509 31452 1545
rect 31352 1475 31452 1509
rect 31352 1439 31385 1475
rect 31419 1439 31452 1475
rect 31352 1407 31452 1439
rect 31352 1367 31385 1407
rect 31419 1367 31452 1407
rect 31352 1339 31452 1367
rect 31352 1295 31385 1339
rect 31419 1295 31452 1339
rect 31352 1271 31452 1295
rect 31352 1223 31385 1271
rect 31419 1223 31452 1271
rect 31352 1203 31452 1223
rect 31352 1151 31385 1203
rect 31419 1151 31452 1203
rect 31352 1135 31452 1151
rect 31352 1079 31385 1135
rect 31419 1079 31452 1135
rect 31352 1067 31452 1079
rect 31352 1007 31385 1067
rect 31419 1007 31452 1067
rect 31352 999 31452 1007
rect 31352 935 31385 999
rect 31419 935 31452 999
rect 31352 931 31452 935
rect 31352 829 31385 931
rect 31419 829 31452 931
rect 31352 825 31452 829
rect 31352 761 31385 825
rect 31419 761 31452 825
rect 31352 753 31452 761
rect 31352 693 31385 753
rect 31419 693 31452 753
rect 31352 681 31452 693
rect 31352 625 31385 681
rect 31419 625 31452 681
rect 31352 609 31452 625
rect 31352 557 31385 609
rect 31419 557 31452 609
rect 31352 537 31452 557
rect 31352 489 31385 537
rect 31419 489 31452 537
rect 31352 465 31452 489
rect 31352 421 31385 465
rect 31419 421 31452 465
rect 31352 393 31452 421
rect 31352 353 31385 393
rect 31419 353 31452 393
rect 31352 321 31452 353
rect 31352 285 31385 321
rect 31419 285 31452 321
rect 31352 251 31452 285
rect 31352 215 31385 251
rect 31419 215 31452 251
rect 31352 183 31452 215
rect 31352 143 31385 183
rect 31419 143 31452 183
rect 31352 115 31452 143
rect 31352 71 31385 115
rect 31419 71 31452 115
rect 31352 47 31452 71
rect 31352 -1 31385 47
rect 31419 -1 31452 47
rect 31352 -21 31452 -1
rect 31352 -73 31385 -21
rect 31419 -73 31452 -21
rect 31352 -89 31452 -73
rect 31352 -145 31385 -89
rect 31419 -145 31452 -89
rect 31352 -157 31452 -145
rect 31352 -217 31385 -157
rect 31419 -217 31452 -157
rect 31352 -225 31452 -217
rect 31352 -289 31385 -225
rect 31419 -289 31452 -225
rect 31352 -293 31452 -289
rect 31352 -395 31385 -293
rect 31419 -395 31452 -293
rect 31352 -399 31452 -395
rect 31352 -463 31385 -399
rect 31419 -463 31452 -399
rect 31352 -471 31452 -463
rect 31352 -531 31385 -471
rect 31419 -531 31452 -471
rect 31352 -543 31452 -531
rect 31352 -599 31385 -543
rect 31419 -599 31452 -543
rect 31352 -615 31452 -599
rect 31352 -667 31385 -615
rect 31419 -667 31452 -615
rect 31352 -687 31452 -667
rect 31352 -735 31385 -687
rect 31419 -735 31452 -687
rect 31352 -759 31452 -735
rect 31352 -803 31385 -759
rect 31419 -803 31452 -759
rect 31352 -831 31452 -803
rect 31352 -871 31385 -831
rect 31419 -871 31452 -831
rect 31352 -903 31452 -871
rect 31352 -939 31385 -903
rect 31419 -939 31452 -903
rect 31352 -973 31452 -939
rect 31352 -1009 31385 -973
rect 31419 -1009 31452 -973
rect 31352 -1041 31452 -1009
rect 31352 -1081 31385 -1041
rect 31419 -1081 31452 -1041
rect 31352 -1109 31452 -1081
rect 31352 -1153 31385 -1109
rect 31419 -1153 31452 -1109
rect 31352 -1177 31452 -1153
rect 31352 -1225 31385 -1177
rect 31419 -1225 31452 -1177
rect 31352 -1245 31452 -1225
rect 31352 -1297 31385 -1245
rect 31419 -1297 31452 -1245
rect 31352 -1313 31452 -1297
rect 31352 -1369 31385 -1313
rect 31419 -1369 31452 -1313
rect 31352 -1381 31452 -1369
rect 31352 -1415 31385 -1381
rect 31419 -1415 31452 -1381
rect 31352 -1449 31452 -1415
rect 31352 -1483 31385 -1449
rect 31419 -1483 31452 -1449
rect 31352 -1558 31452 -1483
rect 26008 -1591 31452 -1558
rect 26008 -1625 26121 -1591
rect 26155 -1625 26193 -1591
rect 26231 -1625 26265 -1591
rect 26299 -1625 26333 -1591
rect 26371 -1625 26401 -1591
rect 26443 -1625 26469 -1591
rect 26515 -1625 26537 -1591
rect 26587 -1625 26605 -1591
rect 26659 -1625 26673 -1591
rect 26731 -1625 26741 -1591
rect 26803 -1625 26809 -1591
rect 26875 -1625 26877 -1591
rect 26911 -1625 26913 -1591
rect 26979 -1625 26985 -1591
rect 27047 -1625 27057 -1591
rect 27115 -1625 27129 -1591
rect 27183 -1625 27201 -1591
rect 27251 -1625 27273 -1591
rect 27319 -1625 27345 -1591
rect 27387 -1625 27417 -1591
rect 27455 -1625 27489 -1591
rect 27523 -1625 27557 -1591
rect 27595 -1625 27625 -1591
rect 27667 -1625 27693 -1591
rect 27739 -1625 27761 -1591
rect 27811 -1625 27829 -1591
rect 27883 -1625 27897 -1591
rect 27955 -1625 27965 -1591
rect 28027 -1625 28033 -1591
rect 28099 -1625 28101 -1591
rect 28135 -1625 28137 -1591
rect 28203 -1625 28209 -1591
rect 28271 -1625 28281 -1591
rect 28339 -1625 28353 -1591
rect 28407 -1625 28425 -1591
rect 28475 -1625 28497 -1591
rect 28543 -1625 28569 -1591
rect 28611 -1625 28641 -1591
rect 28679 -1625 28713 -1591
rect 28747 -1625 28781 -1591
rect 28819 -1625 28849 -1591
rect 28891 -1625 28917 -1591
rect 28963 -1625 28985 -1591
rect 29035 -1625 29053 -1591
rect 29107 -1625 29121 -1591
rect 29179 -1625 29189 -1591
rect 29251 -1625 29257 -1591
rect 29323 -1625 29325 -1591
rect 29359 -1625 29361 -1591
rect 29427 -1625 29433 -1591
rect 29495 -1625 29505 -1591
rect 29563 -1625 29577 -1591
rect 29631 -1625 29649 -1591
rect 29699 -1625 29721 -1591
rect 29767 -1625 29793 -1591
rect 29835 -1625 29865 -1591
rect 29903 -1625 29937 -1591
rect 29971 -1625 30005 -1591
rect 30043 -1625 30073 -1591
rect 30115 -1625 30141 -1591
rect 30187 -1625 30209 -1591
rect 30259 -1625 30277 -1591
rect 30331 -1625 30345 -1591
rect 30403 -1625 30413 -1591
rect 30475 -1625 30481 -1591
rect 30547 -1625 30549 -1591
rect 30583 -1625 30585 -1591
rect 30651 -1625 30657 -1591
rect 30719 -1625 30729 -1591
rect 30787 -1625 30801 -1591
rect 30855 -1625 30873 -1591
rect 30923 -1625 30945 -1591
rect 30991 -1625 31017 -1591
rect 31059 -1625 31089 -1591
rect 31127 -1625 31161 -1591
rect 31195 -1625 31229 -1591
rect 31267 -1625 31305 -1591
rect 31339 -1625 31452 -1591
rect 26008 -1658 31452 -1625
<< viali >>
rect 15529 4243 15563 4277
rect 15601 4243 15603 4277
rect 15603 4243 15635 4277
rect 15673 4243 15705 4277
rect 15705 4243 15707 4277
rect 15745 4243 15773 4277
rect 15773 4243 15779 4277
rect 15817 4243 15841 4277
rect 15841 4243 15851 4277
rect 15889 4243 15909 4277
rect 15909 4243 15923 4277
rect 15961 4243 15977 4277
rect 15977 4243 15995 4277
rect 16033 4243 16045 4277
rect 16045 4243 16067 4277
rect 16105 4243 16113 4277
rect 16113 4243 16139 4277
rect 16177 4243 16181 4277
rect 16181 4243 16211 4277
rect 16249 4243 16283 4277
rect 16321 4243 16351 4277
rect 16351 4243 16355 4277
rect 16393 4243 16419 4277
rect 16419 4243 16427 4277
rect 16465 4243 16487 4277
rect 16487 4243 16499 4277
rect 16537 4243 16555 4277
rect 16555 4243 16571 4277
rect 16609 4243 16623 4277
rect 16623 4243 16643 4277
rect 16681 4243 16691 4277
rect 16691 4243 16715 4277
rect 16753 4243 16759 4277
rect 16759 4243 16787 4277
rect 16825 4243 16827 4277
rect 16827 4243 16859 4277
rect 16897 4243 16929 4277
rect 16929 4243 16931 4277
rect 16969 4243 16997 4277
rect 16997 4243 17003 4277
rect 17041 4243 17065 4277
rect 17065 4243 17075 4277
rect 17113 4243 17133 4277
rect 17133 4243 17147 4277
rect 17185 4243 17201 4277
rect 17201 4243 17219 4277
rect 17257 4243 17269 4277
rect 17269 4243 17291 4277
rect 17329 4243 17337 4277
rect 17337 4243 17363 4277
rect 17401 4243 17405 4277
rect 17405 4243 17435 4277
rect 17473 4243 17507 4277
rect 17545 4243 17575 4277
rect 17575 4243 17579 4277
rect 17617 4243 17643 4277
rect 17643 4243 17651 4277
rect 17689 4243 17711 4277
rect 17711 4243 17723 4277
rect 17761 4243 17779 4277
rect 17779 4243 17795 4277
rect 17833 4243 17847 4277
rect 17847 4243 17867 4277
rect 17905 4243 17915 4277
rect 17915 4243 17939 4277
rect 17977 4243 17983 4277
rect 17983 4243 18011 4277
rect 18049 4243 18051 4277
rect 18051 4243 18083 4277
rect 18121 4243 18153 4277
rect 18153 4243 18155 4277
rect 18193 4243 18221 4277
rect 18221 4243 18227 4277
rect 18265 4243 18289 4277
rect 18289 4243 18299 4277
rect 18337 4243 18357 4277
rect 18357 4243 18371 4277
rect 18409 4243 18425 4277
rect 18425 4243 18443 4277
rect 18481 4243 18493 4277
rect 18493 4243 18515 4277
rect 18553 4243 18561 4277
rect 18561 4243 18587 4277
rect 18625 4243 18629 4277
rect 18629 4243 18659 4277
rect 18697 4243 18731 4277
rect 18769 4243 18799 4277
rect 18799 4243 18803 4277
rect 18841 4243 18867 4277
rect 18867 4243 18875 4277
rect 18913 4243 18935 4277
rect 18935 4243 18947 4277
rect 18985 4243 19003 4277
rect 19003 4243 19019 4277
rect 19057 4243 19071 4277
rect 19071 4243 19091 4277
rect 19129 4243 19139 4277
rect 19139 4243 19163 4277
rect 19201 4243 19207 4277
rect 19207 4243 19235 4277
rect 19273 4243 19275 4277
rect 19275 4243 19307 4277
rect 19345 4243 19377 4277
rect 19377 4243 19379 4277
rect 19417 4243 19445 4277
rect 19445 4243 19451 4277
rect 19489 4243 19513 4277
rect 19513 4243 19523 4277
rect 19561 4243 19581 4277
rect 19581 4243 19595 4277
rect 19633 4243 19649 4277
rect 19649 4243 19667 4277
rect 19705 4243 19717 4277
rect 19717 4243 19739 4277
rect 19777 4243 19785 4277
rect 19785 4243 19811 4277
rect 19849 4243 19853 4277
rect 19853 4243 19883 4277
rect 19921 4243 19955 4277
rect 19993 4243 20023 4277
rect 20023 4243 20027 4277
rect 20065 4243 20091 4277
rect 20091 4243 20099 4277
rect 20137 4243 20159 4277
rect 20159 4243 20171 4277
rect 20209 4243 20227 4277
rect 20227 4243 20243 4277
rect 20281 4243 20295 4277
rect 20295 4243 20315 4277
rect 20353 4243 20363 4277
rect 20363 4243 20387 4277
rect 20425 4243 20431 4277
rect 20431 4243 20459 4277
rect 20497 4243 20499 4277
rect 20499 4243 20531 4277
rect 20569 4243 20601 4277
rect 20601 4243 20603 4277
rect 20641 4243 20669 4277
rect 20669 4243 20675 4277
rect 20713 4243 20737 4277
rect 20737 4243 20747 4277
rect 20785 4243 20805 4277
rect 20805 4243 20819 4277
rect 20857 4243 20873 4277
rect 20873 4243 20891 4277
rect 20929 4243 20941 4277
rect 20941 4243 20963 4277
rect 21001 4243 21009 4277
rect 21009 4243 21035 4277
rect 21073 4243 21077 4277
rect 21077 4243 21107 4277
rect 21145 4243 21179 4277
rect 21217 4243 21247 4277
rect 21247 4243 21251 4277
rect 21289 4243 21315 4277
rect 21315 4243 21323 4277
rect 21361 4243 21383 4277
rect 21383 4243 21395 4277
rect 21433 4243 21451 4277
rect 21451 4243 21467 4277
rect 21505 4243 21519 4277
rect 21519 4243 21539 4277
rect 21577 4243 21587 4277
rect 21587 4243 21611 4277
rect 21649 4243 21655 4277
rect 21655 4243 21683 4277
rect 21721 4243 21723 4277
rect 21723 4243 21755 4277
rect 21793 4243 21825 4277
rect 21825 4243 21827 4277
rect 21865 4243 21893 4277
rect 21893 4243 21899 4277
rect 21937 4243 21961 4277
rect 21961 4243 21971 4277
rect 22009 4243 22029 4277
rect 22029 4243 22043 4277
rect 22081 4243 22097 4277
rect 22097 4243 22115 4277
rect 22153 4243 22165 4277
rect 22165 4243 22187 4277
rect 22225 4243 22233 4277
rect 22233 4243 22259 4277
rect 22297 4243 22301 4277
rect 22301 4243 22331 4277
rect 22369 4243 22403 4277
rect 22441 4243 22471 4277
rect 22471 4243 22475 4277
rect 22513 4243 22539 4277
rect 22539 4243 22547 4277
rect 22585 4243 22607 4277
rect 22607 4243 22619 4277
rect 22657 4243 22675 4277
rect 22675 4243 22691 4277
rect 22729 4243 22743 4277
rect 22743 4243 22763 4277
rect 22801 4243 22811 4277
rect 22811 4243 22835 4277
rect 22873 4243 22879 4277
rect 22879 4243 22907 4277
rect 22945 4243 22947 4277
rect 22947 4243 22979 4277
rect 23017 4243 23049 4277
rect 23049 4243 23051 4277
rect 23089 4243 23117 4277
rect 23117 4243 23123 4277
rect 23161 4243 23185 4277
rect 23185 4243 23195 4277
rect 23233 4243 23253 4277
rect 23253 4243 23267 4277
rect 23305 4243 23321 4277
rect 23321 4243 23339 4277
rect 23377 4243 23389 4277
rect 23389 4243 23411 4277
rect 23449 4243 23457 4277
rect 23457 4243 23483 4277
rect 23521 4243 23525 4277
rect 23525 4243 23555 4277
rect 23593 4243 23627 4277
rect 23665 4243 23695 4277
rect 23695 4243 23699 4277
rect 23737 4243 23763 4277
rect 23763 4243 23771 4277
rect 23809 4243 23831 4277
rect 23831 4243 23843 4277
rect 23881 4243 23899 4277
rect 23899 4243 23915 4277
rect 23953 4243 23967 4277
rect 23967 4243 23987 4277
rect 24025 4243 24035 4277
rect 24035 4243 24059 4277
rect 24097 4243 24103 4277
rect 24103 4243 24131 4277
rect 24169 4243 24171 4277
rect 24171 4243 24203 4277
rect 24241 4243 24273 4277
rect 24273 4243 24275 4277
rect 24313 4243 24347 4277
rect 15459 4107 15493 4111
rect 15459 4077 15493 4107
rect 15459 4005 15493 4039
rect 15459 3937 15493 3967
rect 15459 3933 15493 3937
rect 15459 3869 15493 3895
rect 15459 3861 15493 3869
rect 15459 3801 15493 3823
rect 15459 3789 15493 3801
rect 15459 3733 15493 3751
rect 15459 3717 15493 3733
rect 15459 3665 15493 3679
rect 15459 3645 15493 3665
rect 15459 3597 15493 3607
rect 15459 3573 15493 3597
rect 15459 3529 15493 3535
rect 15459 3501 15493 3529
rect 15459 3461 15493 3463
rect 15459 3429 15493 3461
rect 15459 3359 15493 3391
rect 15459 3357 15493 3359
rect 15459 3291 15493 3319
rect 15459 3285 15493 3291
rect 15459 3223 15493 3247
rect 15459 3213 15493 3223
rect 15459 3155 15493 3175
rect 15459 3141 15493 3155
rect 15459 3087 15493 3103
rect 15459 3069 15493 3087
rect 15459 3019 15493 3031
rect 15459 2997 15493 3019
rect 15459 2951 15493 2959
rect 15459 2925 15493 2951
rect 15459 2883 15493 2887
rect 15459 2853 15493 2883
rect 15459 2781 15493 2815
rect 15459 2713 15493 2743
rect 15459 2709 15493 2713
rect 24383 4107 24417 4111
rect 24383 4077 24417 4107
rect 24383 4005 24417 4039
rect 24383 3937 24417 3967
rect 24383 3933 24417 3937
rect 24383 3869 24417 3895
rect 24383 3861 24417 3869
rect 24383 3801 24417 3823
rect 24383 3789 24417 3801
rect 24383 3733 24417 3751
rect 24383 3717 24417 3733
rect 24383 3665 24417 3679
rect 24383 3645 24417 3665
rect 24383 3597 24417 3607
rect 24383 3573 24417 3597
rect 24383 3529 24417 3535
rect 24383 3501 24417 3529
rect 24383 3461 24417 3463
rect 24383 3429 24417 3461
rect 24383 3359 24417 3391
rect 24383 3357 24417 3359
rect 24383 3291 24417 3319
rect 24383 3285 24417 3291
rect 24383 3223 24417 3247
rect 24383 3213 24417 3223
rect 24383 3155 24417 3175
rect 24383 3141 24417 3155
rect 24383 3087 24417 3103
rect 24383 3069 24417 3087
rect 24383 3019 24417 3031
rect 24383 2997 24417 3019
rect 24383 2951 24417 2959
rect 24383 2925 24417 2951
rect 24383 2883 24417 2887
rect 24383 2853 24417 2883
rect 24383 2781 24417 2815
rect 24383 2713 24417 2743
rect 24383 2709 24417 2713
rect 15529 2543 15563 2577
rect 15601 2543 15603 2577
rect 15603 2543 15635 2577
rect 15673 2543 15705 2577
rect 15705 2543 15707 2577
rect 15745 2543 15773 2577
rect 15773 2543 15779 2577
rect 15817 2543 15841 2577
rect 15841 2543 15851 2577
rect 15889 2543 15909 2577
rect 15909 2543 15923 2577
rect 15961 2543 15977 2577
rect 15977 2543 15995 2577
rect 16033 2543 16045 2577
rect 16045 2543 16067 2577
rect 16105 2543 16113 2577
rect 16113 2543 16139 2577
rect 16177 2543 16181 2577
rect 16181 2543 16211 2577
rect 16249 2543 16283 2577
rect 16321 2543 16351 2577
rect 16351 2543 16355 2577
rect 16393 2543 16419 2577
rect 16419 2543 16427 2577
rect 16465 2543 16487 2577
rect 16487 2543 16499 2577
rect 16537 2543 16555 2577
rect 16555 2543 16571 2577
rect 16609 2543 16623 2577
rect 16623 2543 16643 2577
rect 16681 2543 16691 2577
rect 16691 2543 16715 2577
rect 16753 2543 16759 2577
rect 16759 2543 16787 2577
rect 16825 2543 16827 2577
rect 16827 2543 16859 2577
rect 16897 2543 16929 2577
rect 16929 2543 16931 2577
rect 16969 2543 16997 2577
rect 16997 2543 17003 2577
rect 17041 2543 17065 2577
rect 17065 2543 17075 2577
rect 17113 2543 17133 2577
rect 17133 2543 17147 2577
rect 17185 2543 17201 2577
rect 17201 2543 17219 2577
rect 17257 2543 17269 2577
rect 17269 2543 17291 2577
rect 17329 2543 17337 2577
rect 17337 2543 17363 2577
rect 17401 2543 17405 2577
rect 17405 2543 17435 2577
rect 17473 2543 17507 2577
rect 17545 2543 17575 2577
rect 17575 2543 17579 2577
rect 17617 2543 17643 2577
rect 17643 2543 17651 2577
rect 17689 2543 17711 2577
rect 17711 2543 17723 2577
rect 17761 2543 17779 2577
rect 17779 2543 17795 2577
rect 17833 2543 17847 2577
rect 17847 2543 17867 2577
rect 17905 2543 17915 2577
rect 17915 2543 17939 2577
rect 17977 2543 17983 2577
rect 17983 2543 18011 2577
rect 18049 2543 18051 2577
rect 18051 2543 18083 2577
rect 18121 2543 18153 2577
rect 18153 2543 18155 2577
rect 18193 2543 18221 2577
rect 18221 2543 18227 2577
rect 18265 2543 18289 2577
rect 18289 2543 18299 2577
rect 18337 2543 18357 2577
rect 18357 2543 18371 2577
rect 18409 2543 18425 2577
rect 18425 2543 18443 2577
rect 18481 2543 18493 2577
rect 18493 2543 18515 2577
rect 18553 2543 18561 2577
rect 18561 2543 18587 2577
rect 18625 2543 18629 2577
rect 18629 2543 18659 2577
rect 18697 2543 18731 2577
rect 18769 2543 18799 2577
rect 18799 2543 18803 2577
rect 18841 2543 18867 2577
rect 18867 2543 18875 2577
rect 18913 2543 18935 2577
rect 18935 2543 18947 2577
rect 18985 2543 19003 2577
rect 19003 2543 19019 2577
rect 19057 2543 19071 2577
rect 19071 2543 19091 2577
rect 19129 2543 19139 2577
rect 19139 2543 19163 2577
rect 19201 2543 19207 2577
rect 19207 2543 19235 2577
rect 19273 2543 19275 2577
rect 19275 2543 19307 2577
rect 19345 2543 19377 2577
rect 19377 2543 19379 2577
rect 19417 2543 19445 2577
rect 19445 2543 19451 2577
rect 19489 2543 19513 2577
rect 19513 2543 19523 2577
rect 19561 2543 19581 2577
rect 19581 2543 19595 2577
rect 19633 2543 19649 2577
rect 19649 2543 19667 2577
rect 19705 2543 19717 2577
rect 19717 2543 19739 2577
rect 19777 2543 19785 2577
rect 19785 2543 19811 2577
rect 19849 2543 19853 2577
rect 19853 2543 19883 2577
rect 19921 2543 19955 2577
rect 19993 2543 20023 2577
rect 20023 2543 20027 2577
rect 20065 2543 20091 2577
rect 20091 2543 20099 2577
rect 20137 2543 20159 2577
rect 20159 2543 20171 2577
rect 20209 2543 20227 2577
rect 20227 2543 20243 2577
rect 20281 2543 20295 2577
rect 20295 2543 20315 2577
rect 20353 2543 20363 2577
rect 20363 2543 20387 2577
rect 20425 2543 20431 2577
rect 20431 2543 20459 2577
rect 20497 2543 20499 2577
rect 20499 2543 20531 2577
rect 20569 2543 20601 2577
rect 20601 2543 20603 2577
rect 20641 2543 20669 2577
rect 20669 2543 20675 2577
rect 20713 2543 20737 2577
rect 20737 2543 20747 2577
rect 20785 2543 20805 2577
rect 20805 2543 20819 2577
rect 20857 2543 20873 2577
rect 20873 2543 20891 2577
rect 20929 2543 20941 2577
rect 20941 2543 20963 2577
rect 21001 2543 21009 2577
rect 21009 2543 21035 2577
rect 21073 2543 21077 2577
rect 21077 2543 21107 2577
rect 21145 2543 21179 2577
rect 21217 2543 21247 2577
rect 21247 2543 21251 2577
rect 21289 2543 21315 2577
rect 21315 2543 21323 2577
rect 21361 2543 21383 2577
rect 21383 2543 21395 2577
rect 21433 2543 21451 2577
rect 21451 2543 21467 2577
rect 21505 2543 21519 2577
rect 21519 2543 21539 2577
rect 21577 2543 21587 2577
rect 21587 2543 21611 2577
rect 21649 2543 21655 2577
rect 21655 2543 21683 2577
rect 21721 2543 21723 2577
rect 21723 2543 21755 2577
rect 21793 2543 21825 2577
rect 21825 2543 21827 2577
rect 21865 2543 21893 2577
rect 21893 2543 21899 2577
rect 21937 2543 21961 2577
rect 21961 2543 21971 2577
rect 22009 2543 22029 2577
rect 22029 2543 22043 2577
rect 22081 2543 22097 2577
rect 22097 2543 22115 2577
rect 22153 2543 22165 2577
rect 22165 2543 22187 2577
rect 22225 2543 22233 2577
rect 22233 2543 22259 2577
rect 22297 2543 22301 2577
rect 22301 2543 22331 2577
rect 22369 2543 22403 2577
rect 22441 2543 22471 2577
rect 22471 2543 22475 2577
rect 22513 2543 22539 2577
rect 22539 2543 22547 2577
rect 22585 2543 22607 2577
rect 22607 2543 22619 2577
rect 22657 2543 22675 2577
rect 22675 2543 22691 2577
rect 22729 2543 22743 2577
rect 22743 2543 22763 2577
rect 22801 2543 22811 2577
rect 22811 2543 22835 2577
rect 22873 2543 22879 2577
rect 22879 2543 22907 2577
rect 22945 2543 22947 2577
rect 22947 2543 22979 2577
rect 23017 2543 23049 2577
rect 23049 2543 23051 2577
rect 23089 2543 23117 2577
rect 23117 2543 23123 2577
rect 23161 2543 23185 2577
rect 23185 2543 23195 2577
rect 23233 2543 23253 2577
rect 23253 2543 23267 2577
rect 23305 2543 23321 2577
rect 23321 2543 23339 2577
rect 23377 2543 23389 2577
rect 23389 2543 23411 2577
rect 23449 2543 23457 2577
rect 23457 2543 23483 2577
rect 23521 2543 23525 2577
rect 23525 2543 23555 2577
rect 23593 2543 23627 2577
rect 23665 2543 23695 2577
rect 23695 2543 23699 2577
rect 23737 2543 23763 2577
rect 23763 2543 23771 2577
rect 23809 2543 23831 2577
rect 23831 2543 23843 2577
rect 23881 2543 23899 2577
rect 23899 2543 23915 2577
rect 23953 2543 23967 2577
rect 23967 2543 23987 2577
rect 24025 2543 24035 2577
rect 24035 2543 24059 2577
rect 24097 2543 24103 2577
rect 24103 2543 24131 2577
rect 24169 2543 24171 2577
rect 24171 2543 24203 2577
rect 24241 2543 24273 2577
rect 24273 2543 24275 2577
rect 24313 2543 24347 2577
rect 26121 4243 26155 4277
rect 26193 4243 26197 4277
rect 26197 4243 26227 4277
rect 26265 4243 26299 4277
rect 26337 4243 26367 4277
rect 26367 4243 26371 4277
rect 26409 4243 26435 4277
rect 26435 4243 26443 4277
rect 26481 4243 26503 4277
rect 26503 4243 26515 4277
rect 26553 4243 26571 4277
rect 26571 4243 26587 4277
rect 26625 4243 26639 4277
rect 26639 4243 26659 4277
rect 26697 4243 26707 4277
rect 26707 4243 26731 4277
rect 26769 4243 26775 4277
rect 26775 4243 26803 4277
rect 26841 4243 26843 4277
rect 26843 4243 26875 4277
rect 26913 4243 26945 4277
rect 26945 4243 26947 4277
rect 26985 4243 27013 4277
rect 27013 4243 27019 4277
rect 27057 4243 27081 4277
rect 27081 4243 27091 4277
rect 27129 4243 27149 4277
rect 27149 4243 27163 4277
rect 27201 4243 27217 4277
rect 27217 4243 27235 4277
rect 27273 4243 27285 4277
rect 27285 4243 27307 4277
rect 27345 4243 27353 4277
rect 27353 4243 27379 4277
rect 27417 4243 27421 4277
rect 27421 4243 27451 4277
rect 27489 4243 27523 4277
rect 27561 4243 27591 4277
rect 27591 4243 27595 4277
rect 27633 4243 27659 4277
rect 27659 4243 27667 4277
rect 27705 4243 27727 4277
rect 27727 4243 27739 4277
rect 27777 4243 27795 4277
rect 27795 4243 27811 4277
rect 27849 4243 27863 4277
rect 27863 4243 27883 4277
rect 27921 4243 27931 4277
rect 27931 4243 27955 4277
rect 27993 4243 27999 4277
rect 27999 4243 28027 4277
rect 28065 4243 28067 4277
rect 28067 4243 28099 4277
rect 28137 4243 28169 4277
rect 28169 4243 28171 4277
rect 28209 4243 28237 4277
rect 28237 4243 28243 4277
rect 28281 4243 28305 4277
rect 28305 4243 28315 4277
rect 28353 4243 28373 4277
rect 28373 4243 28387 4277
rect 28425 4243 28441 4277
rect 28441 4243 28459 4277
rect 28497 4243 28509 4277
rect 28509 4243 28531 4277
rect 28569 4243 28577 4277
rect 28577 4243 28603 4277
rect 28641 4243 28645 4277
rect 28645 4243 28675 4277
rect 28713 4243 28747 4277
rect 28785 4243 28815 4277
rect 28815 4243 28819 4277
rect 28857 4243 28883 4277
rect 28883 4243 28891 4277
rect 28929 4243 28951 4277
rect 28951 4243 28963 4277
rect 29001 4243 29019 4277
rect 29019 4243 29035 4277
rect 29073 4243 29087 4277
rect 29087 4243 29107 4277
rect 29145 4243 29155 4277
rect 29155 4243 29179 4277
rect 29217 4243 29223 4277
rect 29223 4243 29251 4277
rect 29289 4243 29291 4277
rect 29291 4243 29323 4277
rect 29361 4243 29393 4277
rect 29393 4243 29395 4277
rect 29433 4243 29461 4277
rect 29461 4243 29467 4277
rect 29505 4243 29529 4277
rect 29529 4243 29539 4277
rect 29577 4243 29597 4277
rect 29597 4243 29611 4277
rect 29649 4243 29665 4277
rect 29665 4243 29683 4277
rect 29721 4243 29733 4277
rect 29733 4243 29755 4277
rect 29793 4243 29801 4277
rect 29801 4243 29827 4277
rect 29865 4243 29869 4277
rect 29869 4243 29899 4277
rect 29937 4243 29971 4277
rect 30009 4243 30039 4277
rect 30039 4243 30043 4277
rect 30081 4243 30107 4277
rect 30107 4243 30115 4277
rect 30153 4243 30175 4277
rect 30175 4243 30187 4277
rect 30225 4243 30243 4277
rect 30243 4243 30259 4277
rect 30297 4243 30311 4277
rect 30311 4243 30331 4277
rect 30369 4243 30379 4277
rect 30379 4243 30403 4277
rect 30441 4243 30447 4277
rect 30447 4243 30475 4277
rect 30513 4243 30515 4277
rect 30515 4243 30547 4277
rect 30585 4243 30617 4277
rect 30617 4243 30619 4277
rect 30657 4243 30685 4277
rect 30685 4243 30691 4277
rect 30729 4243 30753 4277
rect 30753 4243 30763 4277
rect 30801 4243 30821 4277
rect 30821 4243 30835 4277
rect 30873 4243 30889 4277
rect 30889 4243 30907 4277
rect 30945 4243 30957 4277
rect 30957 4243 30979 4277
rect 31017 4243 31025 4277
rect 31025 4243 31051 4277
rect 31089 4243 31093 4277
rect 31093 4243 31123 4277
rect 31161 4243 31195 4277
rect 31233 4243 31263 4277
rect 31263 4243 31267 4277
rect 31305 4243 31339 4277
rect 26041 4101 26075 4107
rect 26041 4073 26075 4101
rect 26041 4033 26075 4035
rect 26041 4001 26075 4033
rect 26041 3931 26075 3963
rect 26041 3929 26075 3931
rect 26041 3863 26075 3891
rect 26041 3857 26075 3863
rect 26041 3795 26075 3819
rect 26041 3785 26075 3795
rect 26041 3727 26075 3747
rect 26041 3713 26075 3727
rect 26041 3659 26075 3675
rect 26041 3641 26075 3659
rect 26041 3591 26075 3603
rect 26041 3569 26075 3591
rect 26041 3523 26075 3531
rect 26041 3497 26075 3523
rect 26041 3455 26075 3459
rect 26041 3425 26075 3455
rect 26041 3353 26075 3387
rect 26041 3285 26075 3315
rect 26041 3281 26075 3285
rect 26041 3217 26075 3243
rect 26041 3209 26075 3217
rect 26041 3149 26075 3171
rect 26041 3137 26075 3149
rect 26041 3081 26075 3099
rect 26041 3065 26075 3081
rect 26041 3013 26075 3027
rect 26041 2993 26075 3013
rect 26041 2945 26075 2955
rect 26041 2921 26075 2945
rect 26041 2877 26075 2883
rect 26041 2849 26075 2877
rect 26041 2809 26075 2811
rect 26041 2777 26075 2809
rect 26041 2707 26075 2739
rect 26041 2705 26075 2707
rect 26041 2639 26075 2667
rect 26041 2633 26075 2639
rect 31385 4101 31419 4107
rect 31385 4073 31419 4101
rect 31385 4033 31419 4035
rect 31385 4001 31419 4033
rect 31385 3931 31419 3963
rect 31385 3929 31419 3931
rect 31385 3863 31419 3891
rect 31385 3857 31419 3863
rect 31385 3795 31419 3819
rect 31385 3785 31419 3795
rect 31385 3727 31419 3747
rect 31385 3713 31419 3727
rect 31385 3659 31419 3675
rect 31385 3641 31419 3659
rect 31385 3591 31419 3603
rect 31385 3569 31419 3591
rect 31385 3523 31419 3531
rect 31385 3497 31419 3523
rect 31385 3455 31419 3459
rect 31385 3425 31419 3455
rect 31385 3353 31419 3387
rect 31385 3285 31419 3315
rect 31385 3281 31419 3285
rect 31385 3217 31419 3243
rect 31385 3209 31419 3217
rect 31385 3149 31419 3171
rect 31385 3137 31419 3149
rect 31385 3081 31419 3099
rect 31385 3065 31419 3081
rect 31385 3013 31419 3027
rect 31385 2993 31419 3013
rect 31385 2945 31419 2955
rect 31385 2921 31419 2945
rect 31385 2877 31419 2883
rect 31385 2849 31419 2877
rect 31385 2809 31419 2811
rect 31385 2777 31419 2809
rect 31385 2707 31419 2739
rect 31385 2705 31419 2707
rect 31385 2639 31419 2667
rect 31385 2633 31419 2639
rect 26121 2463 26155 2497
rect 26193 2463 26197 2497
rect 26197 2463 26227 2497
rect 26265 2463 26299 2497
rect 26337 2463 26367 2497
rect 26367 2463 26371 2497
rect 26409 2463 26435 2497
rect 26435 2463 26443 2497
rect 26481 2463 26503 2497
rect 26503 2463 26515 2497
rect 26553 2463 26571 2497
rect 26571 2463 26587 2497
rect 26625 2463 26639 2497
rect 26639 2463 26659 2497
rect 26697 2463 26707 2497
rect 26707 2463 26731 2497
rect 26769 2463 26775 2497
rect 26775 2463 26803 2497
rect 26841 2463 26843 2497
rect 26843 2463 26875 2497
rect 26913 2463 26945 2497
rect 26945 2463 26947 2497
rect 26985 2463 27013 2497
rect 27013 2463 27019 2497
rect 27057 2463 27081 2497
rect 27081 2463 27091 2497
rect 27129 2463 27149 2497
rect 27149 2463 27163 2497
rect 27201 2463 27217 2497
rect 27217 2463 27235 2497
rect 27273 2463 27285 2497
rect 27285 2463 27307 2497
rect 27345 2463 27353 2497
rect 27353 2463 27379 2497
rect 27417 2463 27421 2497
rect 27421 2463 27451 2497
rect 27489 2463 27523 2497
rect 27561 2463 27591 2497
rect 27591 2463 27595 2497
rect 27633 2463 27659 2497
rect 27659 2463 27667 2497
rect 27705 2463 27727 2497
rect 27727 2463 27739 2497
rect 27777 2463 27795 2497
rect 27795 2463 27811 2497
rect 27849 2463 27863 2497
rect 27863 2463 27883 2497
rect 27921 2463 27931 2497
rect 27931 2463 27955 2497
rect 27993 2463 27999 2497
rect 27999 2463 28027 2497
rect 28065 2463 28067 2497
rect 28067 2463 28099 2497
rect 28137 2463 28169 2497
rect 28169 2463 28171 2497
rect 28209 2463 28237 2497
rect 28237 2463 28243 2497
rect 28281 2463 28305 2497
rect 28305 2463 28315 2497
rect 28353 2463 28373 2497
rect 28373 2463 28387 2497
rect 28425 2463 28441 2497
rect 28441 2463 28459 2497
rect 28497 2463 28509 2497
rect 28509 2463 28531 2497
rect 28569 2463 28577 2497
rect 28577 2463 28603 2497
rect 28641 2463 28645 2497
rect 28645 2463 28675 2497
rect 28713 2463 28747 2497
rect 28785 2463 28815 2497
rect 28815 2463 28819 2497
rect 28857 2463 28883 2497
rect 28883 2463 28891 2497
rect 28929 2463 28951 2497
rect 28951 2463 28963 2497
rect 29001 2463 29019 2497
rect 29019 2463 29035 2497
rect 29073 2463 29087 2497
rect 29087 2463 29107 2497
rect 29145 2463 29155 2497
rect 29155 2463 29179 2497
rect 29217 2463 29223 2497
rect 29223 2463 29251 2497
rect 29289 2463 29291 2497
rect 29291 2463 29323 2497
rect 29361 2463 29393 2497
rect 29393 2463 29395 2497
rect 29433 2463 29461 2497
rect 29461 2463 29467 2497
rect 29505 2463 29529 2497
rect 29529 2463 29539 2497
rect 29577 2463 29597 2497
rect 29597 2463 29611 2497
rect 29649 2463 29665 2497
rect 29665 2463 29683 2497
rect 29721 2463 29733 2497
rect 29733 2463 29755 2497
rect 29793 2463 29801 2497
rect 29801 2463 29827 2497
rect 29865 2463 29869 2497
rect 29869 2463 29899 2497
rect 29937 2463 29971 2497
rect 30009 2463 30039 2497
rect 30039 2463 30043 2497
rect 30081 2463 30107 2497
rect 30107 2463 30115 2497
rect 30153 2463 30175 2497
rect 30175 2463 30187 2497
rect 30225 2463 30243 2497
rect 30243 2463 30259 2497
rect 30297 2463 30311 2497
rect 30311 2463 30331 2497
rect 30369 2463 30379 2497
rect 30379 2463 30403 2497
rect 30441 2463 30447 2497
rect 30447 2463 30475 2497
rect 30513 2463 30515 2497
rect 30515 2463 30547 2497
rect 30585 2463 30617 2497
rect 30617 2463 30619 2497
rect 30657 2463 30685 2497
rect 30685 2463 30691 2497
rect 30729 2463 30753 2497
rect 30753 2463 30763 2497
rect 30801 2463 30821 2497
rect 30821 2463 30835 2497
rect 30873 2463 30889 2497
rect 30889 2463 30907 2497
rect 30945 2463 30957 2497
rect 30957 2463 30979 2497
rect 31017 2463 31025 2497
rect 31025 2463 31051 2497
rect 31089 2463 31093 2497
rect 31093 2463 31123 2497
rect 31161 2463 31195 2497
rect 31233 2463 31263 2497
rect 31263 2463 31267 2497
rect 31305 2463 31339 2497
rect 15529 2207 15563 2241
rect 15601 2207 15603 2241
rect 15603 2207 15635 2241
rect 15673 2207 15705 2241
rect 15705 2207 15707 2241
rect 15745 2207 15773 2241
rect 15773 2207 15779 2241
rect 15817 2207 15841 2241
rect 15841 2207 15851 2241
rect 15889 2207 15909 2241
rect 15909 2207 15923 2241
rect 15961 2207 15977 2241
rect 15977 2207 15995 2241
rect 16033 2207 16045 2241
rect 16045 2207 16067 2241
rect 16105 2207 16113 2241
rect 16113 2207 16139 2241
rect 16177 2207 16181 2241
rect 16181 2207 16211 2241
rect 16249 2207 16283 2241
rect 16321 2207 16351 2241
rect 16351 2207 16355 2241
rect 16393 2207 16419 2241
rect 16419 2207 16427 2241
rect 16465 2207 16487 2241
rect 16487 2207 16499 2241
rect 16537 2207 16555 2241
rect 16555 2207 16571 2241
rect 16609 2207 16623 2241
rect 16623 2207 16643 2241
rect 16681 2207 16691 2241
rect 16691 2207 16715 2241
rect 16753 2207 16759 2241
rect 16759 2207 16787 2241
rect 16825 2207 16827 2241
rect 16827 2207 16859 2241
rect 16897 2207 16929 2241
rect 16929 2207 16931 2241
rect 16969 2207 16997 2241
rect 16997 2207 17003 2241
rect 17041 2207 17065 2241
rect 17065 2207 17075 2241
rect 17113 2207 17133 2241
rect 17133 2207 17147 2241
rect 17185 2207 17201 2241
rect 17201 2207 17219 2241
rect 17257 2207 17269 2241
rect 17269 2207 17291 2241
rect 17329 2207 17337 2241
rect 17337 2207 17363 2241
rect 17401 2207 17405 2241
rect 17405 2207 17435 2241
rect 17473 2207 17507 2241
rect 17545 2207 17575 2241
rect 17575 2207 17579 2241
rect 17617 2207 17643 2241
rect 17643 2207 17651 2241
rect 17689 2207 17711 2241
rect 17711 2207 17723 2241
rect 17761 2207 17779 2241
rect 17779 2207 17795 2241
rect 17833 2207 17847 2241
rect 17847 2207 17867 2241
rect 17905 2207 17915 2241
rect 17915 2207 17939 2241
rect 17977 2207 17983 2241
rect 17983 2207 18011 2241
rect 18049 2207 18051 2241
rect 18051 2207 18083 2241
rect 18121 2207 18153 2241
rect 18153 2207 18155 2241
rect 18193 2207 18221 2241
rect 18221 2207 18227 2241
rect 18265 2207 18289 2241
rect 18289 2207 18299 2241
rect 18337 2207 18357 2241
rect 18357 2207 18371 2241
rect 18409 2207 18425 2241
rect 18425 2207 18443 2241
rect 18481 2207 18493 2241
rect 18493 2207 18515 2241
rect 18553 2207 18561 2241
rect 18561 2207 18587 2241
rect 18625 2207 18629 2241
rect 18629 2207 18659 2241
rect 18697 2207 18731 2241
rect 18769 2207 18799 2241
rect 18799 2207 18803 2241
rect 18841 2207 18867 2241
rect 18867 2207 18875 2241
rect 18913 2207 18935 2241
rect 18935 2207 18947 2241
rect 18985 2207 19003 2241
rect 19003 2207 19019 2241
rect 19057 2207 19071 2241
rect 19071 2207 19091 2241
rect 19129 2207 19139 2241
rect 19139 2207 19163 2241
rect 19201 2207 19207 2241
rect 19207 2207 19235 2241
rect 19273 2207 19275 2241
rect 19275 2207 19307 2241
rect 19345 2207 19377 2241
rect 19377 2207 19379 2241
rect 19417 2207 19445 2241
rect 19445 2207 19451 2241
rect 19489 2207 19513 2241
rect 19513 2207 19523 2241
rect 19561 2207 19581 2241
rect 19581 2207 19595 2241
rect 19633 2207 19649 2241
rect 19649 2207 19667 2241
rect 19705 2207 19717 2241
rect 19717 2207 19739 2241
rect 19777 2207 19785 2241
rect 19785 2207 19811 2241
rect 19849 2207 19853 2241
rect 19853 2207 19883 2241
rect 19921 2207 19955 2241
rect 19993 2207 20023 2241
rect 20023 2207 20027 2241
rect 20065 2207 20091 2241
rect 20091 2207 20099 2241
rect 20137 2207 20159 2241
rect 20159 2207 20171 2241
rect 20209 2207 20227 2241
rect 20227 2207 20243 2241
rect 20281 2207 20295 2241
rect 20295 2207 20315 2241
rect 20353 2207 20363 2241
rect 20363 2207 20387 2241
rect 20425 2207 20431 2241
rect 20431 2207 20459 2241
rect 20497 2207 20499 2241
rect 20499 2207 20531 2241
rect 20569 2207 20601 2241
rect 20601 2207 20603 2241
rect 20641 2207 20669 2241
rect 20669 2207 20675 2241
rect 20713 2207 20737 2241
rect 20737 2207 20747 2241
rect 20785 2207 20805 2241
rect 20805 2207 20819 2241
rect 20857 2207 20873 2241
rect 20873 2207 20891 2241
rect 20929 2207 20941 2241
rect 20941 2207 20963 2241
rect 21001 2207 21009 2241
rect 21009 2207 21035 2241
rect 21073 2207 21077 2241
rect 21077 2207 21107 2241
rect 21145 2207 21179 2241
rect 21217 2207 21247 2241
rect 21247 2207 21251 2241
rect 21289 2207 21315 2241
rect 21315 2207 21323 2241
rect 21361 2207 21383 2241
rect 21383 2207 21395 2241
rect 21433 2207 21451 2241
rect 21451 2207 21467 2241
rect 21505 2207 21519 2241
rect 21519 2207 21539 2241
rect 21577 2207 21587 2241
rect 21587 2207 21611 2241
rect 21649 2207 21655 2241
rect 21655 2207 21683 2241
rect 21721 2207 21723 2241
rect 21723 2207 21755 2241
rect 21793 2207 21825 2241
rect 21825 2207 21827 2241
rect 21865 2207 21893 2241
rect 21893 2207 21899 2241
rect 21937 2207 21961 2241
rect 21961 2207 21971 2241
rect 22009 2207 22029 2241
rect 22029 2207 22043 2241
rect 22081 2207 22097 2241
rect 22097 2207 22115 2241
rect 22153 2207 22165 2241
rect 22165 2207 22187 2241
rect 22225 2207 22233 2241
rect 22233 2207 22259 2241
rect 22297 2207 22301 2241
rect 22301 2207 22331 2241
rect 22369 2207 22403 2241
rect 22441 2207 22471 2241
rect 22471 2207 22475 2241
rect 22513 2207 22539 2241
rect 22539 2207 22547 2241
rect 22585 2207 22607 2241
rect 22607 2207 22619 2241
rect 22657 2207 22675 2241
rect 22675 2207 22691 2241
rect 22729 2207 22743 2241
rect 22743 2207 22763 2241
rect 22801 2207 22811 2241
rect 22811 2207 22835 2241
rect 22873 2207 22879 2241
rect 22879 2207 22907 2241
rect 22945 2207 22947 2241
rect 22947 2207 22979 2241
rect 23017 2207 23049 2241
rect 23049 2207 23051 2241
rect 23089 2207 23117 2241
rect 23117 2207 23123 2241
rect 23161 2207 23185 2241
rect 23185 2207 23195 2241
rect 23233 2207 23253 2241
rect 23253 2207 23267 2241
rect 23305 2207 23321 2241
rect 23321 2207 23339 2241
rect 23377 2207 23389 2241
rect 23389 2207 23411 2241
rect 23449 2207 23457 2241
rect 23457 2207 23483 2241
rect 23521 2207 23525 2241
rect 23525 2207 23555 2241
rect 23593 2207 23627 2241
rect 23665 2207 23695 2241
rect 23695 2207 23699 2241
rect 23737 2207 23763 2241
rect 23763 2207 23771 2241
rect 23809 2207 23831 2241
rect 23831 2207 23843 2241
rect 23881 2207 23899 2241
rect 23899 2207 23915 2241
rect 23953 2207 23967 2241
rect 23967 2207 23987 2241
rect 24025 2207 24035 2241
rect 24035 2207 24059 2241
rect 24097 2207 24103 2241
rect 24103 2207 24131 2241
rect 24169 2207 24171 2241
rect 24171 2207 24203 2241
rect 24241 2207 24273 2241
rect 24273 2207 24275 2241
rect 24313 2207 24347 2241
rect 31613 2233 31647 2267
rect 31719 2235 31753 2269
rect 31855 2235 31889 2269
rect 32211 2235 32245 2269
rect 15459 1923 15493 1945
rect 15459 1911 15493 1923
rect 15459 1855 15493 1873
rect 15459 1839 15493 1855
rect 15459 1787 15493 1801
rect 15459 1767 15493 1787
rect 15459 1719 15493 1729
rect 15459 1695 15493 1719
rect 15459 1651 15493 1657
rect 15459 1623 15493 1651
rect 15459 1583 15493 1585
rect 15459 1551 15493 1583
rect 15459 1481 15493 1513
rect 15459 1479 15493 1481
rect 15459 1413 15493 1441
rect 15459 1407 15493 1413
rect 15459 1345 15493 1369
rect 15459 1335 15493 1345
rect 15459 1277 15493 1297
rect 15459 1263 15493 1277
rect 15459 1209 15493 1225
rect 15459 1191 15493 1209
rect 15459 1141 15493 1153
rect 15459 1119 15493 1141
rect 15459 1073 15493 1081
rect 15459 1047 15493 1073
rect 15459 1005 15493 1009
rect 15459 975 15493 1005
rect 15459 903 15493 937
rect 15459 835 15493 865
rect 15459 831 15493 835
rect 15459 767 15493 793
rect 15459 759 15493 767
rect 15459 699 15493 721
rect 15459 687 15493 699
rect 15459 631 15493 649
rect 15459 615 15493 631
rect 15459 563 15493 577
rect 15459 543 15493 563
rect 15459 495 15493 505
rect 15459 471 15493 495
rect 15459 427 15493 433
rect 15459 399 15493 427
rect 15459 359 15493 361
rect 15459 327 15493 359
rect 15459 257 15493 289
rect 15459 255 15493 257
rect 15459 189 15493 217
rect 15459 183 15493 189
rect 15459 121 15493 145
rect 15459 111 15493 121
rect 15459 53 15493 73
rect 15459 39 15493 53
rect 15459 -15 15493 1
rect 15459 -33 15493 -15
rect 15459 -83 15493 -71
rect 15459 -105 15493 -83
rect 15459 -151 15493 -143
rect 15459 -177 15493 -151
rect 15459 -219 15493 -215
rect 15459 -249 15493 -219
rect 15459 -321 15493 -287
rect 15459 -389 15493 -359
rect 15459 -393 15493 -389
rect 15459 -457 15493 -431
rect 15459 -465 15493 -457
rect 15459 -525 15493 -503
rect 15459 -537 15493 -525
rect 15459 -593 15493 -575
rect 15459 -609 15493 -593
rect 15459 -661 15493 -647
rect 15459 -681 15493 -661
rect 15459 -729 15493 -719
rect 15459 -753 15493 -729
rect 15459 -797 15493 -791
rect 15459 -825 15493 -797
rect 15459 -865 15493 -863
rect 15459 -897 15493 -865
rect 15459 -967 15493 -935
rect 15459 -969 15493 -967
rect 15459 -1035 15493 -1007
rect 15459 -1041 15493 -1035
rect 15459 -1103 15493 -1079
rect 15459 -1113 15493 -1103
rect 15459 -1171 15493 -1151
rect 15459 -1185 15493 -1171
rect 15459 -1239 15493 -1223
rect 15459 -1257 15493 -1239
rect 15459 -1307 15493 -1295
rect 15459 -1329 15493 -1307
rect 24383 1923 24417 1945
rect 24383 1911 24417 1923
rect 24383 1855 24417 1873
rect 24383 1839 24417 1855
rect 24383 1787 24417 1801
rect 24383 1767 24417 1787
rect 24383 1719 24417 1729
rect 24383 1695 24417 1719
rect 24383 1651 24417 1657
rect 24383 1623 24417 1651
rect 24383 1583 24417 1585
rect 24383 1551 24417 1583
rect 24383 1481 24417 1513
rect 24383 1479 24417 1481
rect 24383 1413 24417 1441
rect 24383 1407 24417 1413
rect 24383 1345 24417 1369
rect 24383 1335 24417 1345
rect 24383 1277 24417 1297
rect 24383 1263 24417 1277
rect 24383 1209 24417 1225
rect 24383 1191 24417 1209
rect 24383 1141 24417 1153
rect 24383 1119 24417 1141
rect 24383 1073 24417 1081
rect 24383 1047 24417 1073
rect 24383 1005 24417 1009
rect 24383 975 24417 1005
rect 24383 903 24417 937
rect 24383 835 24417 865
rect 24383 831 24417 835
rect 24383 767 24417 793
rect 24383 759 24417 767
rect 24383 699 24417 721
rect 24383 687 24417 699
rect 24383 631 24417 649
rect 24383 615 24417 631
rect 24383 563 24417 577
rect 24383 543 24417 563
rect 24383 495 24417 505
rect 24383 471 24417 495
rect 24383 427 24417 433
rect 24383 399 24417 427
rect 24383 359 24417 361
rect 24383 327 24417 359
rect 24383 257 24417 289
rect 24383 255 24417 257
rect 24383 189 24417 217
rect 24383 183 24417 189
rect 24383 121 24417 145
rect 24383 111 24417 121
rect 24383 53 24417 73
rect 24383 39 24417 53
rect 24383 -15 24417 1
rect 24383 -33 24417 -15
rect 24383 -83 24417 -71
rect 24383 -105 24417 -83
rect 24383 -151 24417 -143
rect 24383 -177 24417 -151
rect 24383 -219 24417 -215
rect 24383 -249 24417 -219
rect 24383 -321 24417 -287
rect 24383 -389 24417 -359
rect 24383 -393 24417 -389
rect 24383 -457 24417 -431
rect 24383 -465 24417 -457
rect 24383 -525 24417 -503
rect 24383 -537 24417 -525
rect 24383 -593 24417 -575
rect 24383 -609 24417 -593
rect 24383 -661 24417 -647
rect 24383 -681 24417 -661
rect 24383 -729 24417 -719
rect 24383 -753 24417 -729
rect 24383 -797 24417 -791
rect 24383 -825 24417 -797
rect 24383 -865 24417 -863
rect 24383 -897 24417 -865
rect 24383 -967 24417 -935
rect 24383 -969 24417 -967
rect 24383 -1035 24417 -1007
rect 24383 -1041 24417 -1035
rect 24383 -1103 24417 -1079
rect 24383 -1113 24417 -1103
rect 24383 -1171 24417 -1151
rect 24383 -1185 24417 -1171
rect 24383 -1239 24417 -1223
rect 24383 -1257 24417 -1239
rect 24383 -1307 24417 -1295
rect 24383 -1329 24417 -1307
rect 15529 -1625 15563 -1591
rect 15601 -1625 15603 -1591
rect 15603 -1625 15635 -1591
rect 15673 -1625 15705 -1591
rect 15705 -1625 15707 -1591
rect 15745 -1625 15773 -1591
rect 15773 -1625 15779 -1591
rect 15817 -1625 15841 -1591
rect 15841 -1625 15851 -1591
rect 15889 -1625 15909 -1591
rect 15909 -1625 15923 -1591
rect 15961 -1625 15977 -1591
rect 15977 -1625 15995 -1591
rect 16033 -1625 16045 -1591
rect 16045 -1625 16067 -1591
rect 16105 -1625 16113 -1591
rect 16113 -1625 16139 -1591
rect 16177 -1625 16181 -1591
rect 16181 -1625 16211 -1591
rect 16249 -1625 16283 -1591
rect 16321 -1625 16351 -1591
rect 16351 -1625 16355 -1591
rect 16393 -1625 16419 -1591
rect 16419 -1625 16427 -1591
rect 16465 -1625 16487 -1591
rect 16487 -1625 16499 -1591
rect 16537 -1625 16555 -1591
rect 16555 -1625 16571 -1591
rect 16609 -1625 16623 -1591
rect 16623 -1625 16643 -1591
rect 16681 -1625 16691 -1591
rect 16691 -1625 16715 -1591
rect 16753 -1625 16759 -1591
rect 16759 -1625 16787 -1591
rect 16825 -1625 16827 -1591
rect 16827 -1625 16859 -1591
rect 16897 -1625 16929 -1591
rect 16929 -1625 16931 -1591
rect 16969 -1625 16997 -1591
rect 16997 -1625 17003 -1591
rect 17041 -1625 17065 -1591
rect 17065 -1625 17075 -1591
rect 17113 -1625 17133 -1591
rect 17133 -1625 17147 -1591
rect 17185 -1625 17201 -1591
rect 17201 -1625 17219 -1591
rect 17257 -1625 17269 -1591
rect 17269 -1625 17291 -1591
rect 17329 -1625 17337 -1591
rect 17337 -1625 17363 -1591
rect 17401 -1625 17405 -1591
rect 17405 -1625 17435 -1591
rect 17473 -1625 17507 -1591
rect 17545 -1625 17575 -1591
rect 17575 -1625 17579 -1591
rect 17617 -1625 17643 -1591
rect 17643 -1625 17651 -1591
rect 17689 -1625 17711 -1591
rect 17711 -1625 17723 -1591
rect 17761 -1625 17779 -1591
rect 17779 -1625 17795 -1591
rect 17833 -1625 17847 -1591
rect 17847 -1625 17867 -1591
rect 17905 -1625 17915 -1591
rect 17915 -1625 17939 -1591
rect 17977 -1625 17983 -1591
rect 17983 -1625 18011 -1591
rect 18049 -1625 18051 -1591
rect 18051 -1625 18083 -1591
rect 18121 -1625 18153 -1591
rect 18153 -1625 18155 -1591
rect 18193 -1625 18221 -1591
rect 18221 -1625 18227 -1591
rect 18265 -1625 18289 -1591
rect 18289 -1625 18299 -1591
rect 18337 -1625 18357 -1591
rect 18357 -1625 18371 -1591
rect 18409 -1625 18425 -1591
rect 18425 -1625 18443 -1591
rect 18481 -1625 18493 -1591
rect 18493 -1625 18515 -1591
rect 18553 -1625 18561 -1591
rect 18561 -1625 18587 -1591
rect 18625 -1625 18629 -1591
rect 18629 -1625 18659 -1591
rect 18697 -1625 18731 -1591
rect 18769 -1625 18799 -1591
rect 18799 -1625 18803 -1591
rect 18841 -1625 18867 -1591
rect 18867 -1625 18875 -1591
rect 18913 -1625 18935 -1591
rect 18935 -1625 18947 -1591
rect 18985 -1625 19003 -1591
rect 19003 -1625 19019 -1591
rect 19057 -1625 19071 -1591
rect 19071 -1625 19091 -1591
rect 19129 -1625 19139 -1591
rect 19139 -1625 19163 -1591
rect 19201 -1625 19207 -1591
rect 19207 -1625 19235 -1591
rect 19273 -1625 19275 -1591
rect 19275 -1625 19307 -1591
rect 19345 -1625 19377 -1591
rect 19377 -1625 19379 -1591
rect 19417 -1625 19445 -1591
rect 19445 -1625 19451 -1591
rect 19489 -1625 19513 -1591
rect 19513 -1625 19523 -1591
rect 19561 -1625 19581 -1591
rect 19581 -1625 19595 -1591
rect 19633 -1625 19649 -1591
rect 19649 -1625 19667 -1591
rect 19705 -1625 19717 -1591
rect 19717 -1625 19739 -1591
rect 19777 -1625 19785 -1591
rect 19785 -1625 19811 -1591
rect 19849 -1625 19853 -1591
rect 19853 -1625 19883 -1591
rect 19921 -1625 19955 -1591
rect 19993 -1625 20023 -1591
rect 20023 -1625 20027 -1591
rect 20065 -1625 20091 -1591
rect 20091 -1625 20099 -1591
rect 20137 -1625 20159 -1591
rect 20159 -1625 20171 -1591
rect 20209 -1625 20227 -1591
rect 20227 -1625 20243 -1591
rect 20281 -1625 20295 -1591
rect 20295 -1625 20315 -1591
rect 20353 -1625 20363 -1591
rect 20363 -1625 20387 -1591
rect 20425 -1625 20431 -1591
rect 20431 -1625 20459 -1591
rect 20497 -1625 20499 -1591
rect 20499 -1625 20531 -1591
rect 20569 -1625 20601 -1591
rect 20601 -1625 20603 -1591
rect 20641 -1625 20669 -1591
rect 20669 -1625 20675 -1591
rect 20713 -1625 20737 -1591
rect 20737 -1625 20747 -1591
rect 20785 -1625 20805 -1591
rect 20805 -1625 20819 -1591
rect 20857 -1625 20873 -1591
rect 20873 -1625 20891 -1591
rect 20929 -1625 20941 -1591
rect 20941 -1625 20963 -1591
rect 21001 -1625 21009 -1591
rect 21009 -1625 21035 -1591
rect 21073 -1625 21077 -1591
rect 21077 -1625 21107 -1591
rect 21145 -1625 21179 -1591
rect 21217 -1625 21247 -1591
rect 21247 -1625 21251 -1591
rect 21289 -1625 21315 -1591
rect 21315 -1625 21323 -1591
rect 21361 -1625 21383 -1591
rect 21383 -1625 21395 -1591
rect 21433 -1625 21451 -1591
rect 21451 -1625 21467 -1591
rect 21505 -1625 21519 -1591
rect 21519 -1625 21539 -1591
rect 21577 -1625 21587 -1591
rect 21587 -1625 21611 -1591
rect 21649 -1625 21655 -1591
rect 21655 -1625 21683 -1591
rect 21721 -1625 21723 -1591
rect 21723 -1625 21755 -1591
rect 21793 -1625 21825 -1591
rect 21825 -1625 21827 -1591
rect 21865 -1625 21893 -1591
rect 21893 -1625 21899 -1591
rect 21937 -1625 21961 -1591
rect 21961 -1625 21971 -1591
rect 22009 -1625 22029 -1591
rect 22029 -1625 22043 -1591
rect 22081 -1625 22097 -1591
rect 22097 -1625 22115 -1591
rect 22153 -1625 22165 -1591
rect 22165 -1625 22187 -1591
rect 22225 -1625 22233 -1591
rect 22233 -1625 22259 -1591
rect 22297 -1625 22301 -1591
rect 22301 -1625 22331 -1591
rect 22369 -1625 22403 -1591
rect 22441 -1625 22471 -1591
rect 22471 -1625 22475 -1591
rect 22513 -1625 22539 -1591
rect 22539 -1625 22547 -1591
rect 22585 -1625 22607 -1591
rect 22607 -1625 22619 -1591
rect 22657 -1625 22675 -1591
rect 22675 -1625 22691 -1591
rect 22729 -1625 22743 -1591
rect 22743 -1625 22763 -1591
rect 22801 -1625 22811 -1591
rect 22811 -1625 22835 -1591
rect 22873 -1625 22879 -1591
rect 22879 -1625 22907 -1591
rect 22945 -1625 22947 -1591
rect 22947 -1625 22979 -1591
rect 23017 -1625 23049 -1591
rect 23049 -1625 23051 -1591
rect 23089 -1625 23117 -1591
rect 23117 -1625 23123 -1591
rect 23161 -1625 23185 -1591
rect 23185 -1625 23195 -1591
rect 23233 -1625 23253 -1591
rect 23253 -1625 23267 -1591
rect 23305 -1625 23321 -1591
rect 23321 -1625 23339 -1591
rect 23377 -1625 23389 -1591
rect 23389 -1625 23411 -1591
rect 23449 -1625 23457 -1591
rect 23457 -1625 23483 -1591
rect 23521 -1625 23525 -1591
rect 23525 -1625 23555 -1591
rect 23593 -1625 23627 -1591
rect 23665 -1625 23695 -1591
rect 23695 -1625 23699 -1591
rect 23737 -1625 23763 -1591
rect 23763 -1625 23771 -1591
rect 23809 -1625 23831 -1591
rect 23831 -1625 23843 -1591
rect 23881 -1625 23899 -1591
rect 23899 -1625 23915 -1591
rect 23953 -1625 23967 -1591
rect 23967 -1625 23987 -1591
rect 24025 -1625 24035 -1591
rect 24035 -1625 24059 -1591
rect 24097 -1625 24103 -1591
rect 24103 -1625 24131 -1591
rect 24169 -1625 24171 -1591
rect 24171 -1625 24203 -1591
rect 24241 -1625 24273 -1591
rect 24273 -1625 24275 -1591
rect 24313 -1625 24347 -1591
rect 26121 2127 26155 2161
rect 26193 2127 26197 2161
rect 26197 2127 26227 2161
rect 26265 2127 26299 2161
rect 26337 2127 26367 2161
rect 26367 2127 26371 2161
rect 26409 2127 26435 2161
rect 26435 2127 26443 2161
rect 26481 2127 26503 2161
rect 26503 2127 26515 2161
rect 26553 2127 26571 2161
rect 26571 2127 26587 2161
rect 26625 2127 26639 2161
rect 26639 2127 26659 2161
rect 26697 2127 26707 2161
rect 26707 2127 26731 2161
rect 26769 2127 26775 2161
rect 26775 2127 26803 2161
rect 26841 2127 26843 2161
rect 26843 2127 26875 2161
rect 26913 2127 26945 2161
rect 26945 2127 26947 2161
rect 26985 2127 27013 2161
rect 27013 2127 27019 2161
rect 27057 2127 27081 2161
rect 27081 2127 27091 2161
rect 27129 2127 27149 2161
rect 27149 2127 27163 2161
rect 27201 2127 27217 2161
rect 27217 2127 27235 2161
rect 27273 2127 27285 2161
rect 27285 2127 27307 2161
rect 27345 2127 27353 2161
rect 27353 2127 27379 2161
rect 27417 2127 27421 2161
rect 27421 2127 27451 2161
rect 27489 2127 27523 2161
rect 27561 2127 27591 2161
rect 27591 2127 27595 2161
rect 27633 2127 27659 2161
rect 27659 2127 27667 2161
rect 27705 2127 27727 2161
rect 27727 2127 27739 2161
rect 27777 2127 27795 2161
rect 27795 2127 27811 2161
rect 27849 2127 27863 2161
rect 27863 2127 27883 2161
rect 27921 2127 27931 2161
rect 27931 2127 27955 2161
rect 27993 2127 27999 2161
rect 27999 2127 28027 2161
rect 28065 2127 28067 2161
rect 28067 2127 28099 2161
rect 28137 2127 28169 2161
rect 28169 2127 28171 2161
rect 28209 2127 28237 2161
rect 28237 2127 28243 2161
rect 28281 2127 28305 2161
rect 28305 2127 28315 2161
rect 28353 2127 28373 2161
rect 28373 2127 28387 2161
rect 28425 2127 28441 2161
rect 28441 2127 28459 2161
rect 28497 2127 28509 2161
rect 28509 2127 28531 2161
rect 28569 2127 28577 2161
rect 28577 2127 28603 2161
rect 28641 2127 28645 2161
rect 28645 2127 28675 2161
rect 28713 2127 28747 2161
rect 28785 2127 28815 2161
rect 28815 2127 28819 2161
rect 28857 2127 28883 2161
rect 28883 2127 28891 2161
rect 28929 2127 28951 2161
rect 28951 2127 28963 2161
rect 29001 2127 29019 2161
rect 29019 2127 29035 2161
rect 29073 2127 29087 2161
rect 29087 2127 29107 2161
rect 29145 2127 29155 2161
rect 29155 2127 29179 2161
rect 29217 2127 29223 2161
rect 29223 2127 29251 2161
rect 29289 2127 29291 2161
rect 29291 2127 29323 2161
rect 29361 2127 29393 2161
rect 29393 2127 29395 2161
rect 29433 2127 29461 2161
rect 29461 2127 29467 2161
rect 29505 2127 29529 2161
rect 29529 2127 29539 2161
rect 29577 2127 29597 2161
rect 29597 2127 29611 2161
rect 29649 2127 29665 2161
rect 29665 2127 29683 2161
rect 29721 2127 29733 2161
rect 29733 2127 29755 2161
rect 29793 2127 29801 2161
rect 29801 2127 29827 2161
rect 29865 2127 29869 2161
rect 29869 2127 29899 2161
rect 29937 2127 29971 2161
rect 30009 2127 30039 2161
rect 30039 2127 30043 2161
rect 30081 2127 30107 2161
rect 30107 2127 30115 2161
rect 30153 2127 30175 2161
rect 30175 2127 30187 2161
rect 30225 2127 30243 2161
rect 30243 2127 30259 2161
rect 30297 2127 30311 2161
rect 30311 2127 30331 2161
rect 30369 2127 30379 2161
rect 30379 2127 30403 2161
rect 30441 2127 30447 2161
rect 30447 2127 30475 2161
rect 30513 2127 30515 2161
rect 30515 2127 30547 2161
rect 30585 2127 30617 2161
rect 30617 2127 30619 2161
rect 30657 2127 30685 2161
rect 30685 2127 30691 2161
rect 30729 2127 30753 2161
rect 30753 2127 30763 2161
rect 30801 2127 30821 2161
rect 30821 2127 30835 2161
rect 30873 2127 30889 2161
rect 30889 2127 30907 2161
rect 30945 2127 30957 2161
rect 30957 2127 30979 2161
rect 31017 2127 31025 2161
rect 31025 2127 31051 2161
rect 31089 2127 31093 2161
rect 31093 2127 31123 2161
rect 31161 2127 31195 2161
rect 31233 2127 31263 2161
rect 31263 2127 31267 2161
rect 31305 2127 31339 2161
rect 26041 1883 26075 1905
rect 26041 1871 26075 1883
rect 26041 1815 26075 1833
rect 26041 1799 26075 1815
rect 26041 1747 26075 1761
rect 26041 1727 26075 1747
rect 26041 1679 26075 1689
rect 26041 1655 26075 1679
rect 26041 1611 26075 1617
rect 26041 1583 26075 1611
rect 26041 1543 26075 1545
rect 26041 1511 26075 1543
rect 26041 1441 26075 1473
rect 26041 1439 26075 1441
rect 26041 1373 26075 1401
rect 26041 1367 26075 1373
rect 26041 1305 26075 1329
rect 26041 1295 26075 1305
rect 26041 1237 26075 1257
rect 26041 1223 26075 1237
rect 26041 1169 26075 1185
rect 26041 1151 26075 1169
rect 26041 1101 26075 1113
rect 26041 1079 26075 1101
rect 26041 1033 26075 1041
rect 26041 1007 26075 1033
rect 26041 965 26075 969
rect 26041 935 26075 965
rect 26041 863 26075 897
rect 26041 795 26075 825
rect 26041 791 26075 795
rect 26041 727 26075 753
rect 26041 719 26075 727
rect 26041 659 26075 681
rect 26041 647 26075 659
rect 26041 591 26075 609
rect 26041 575 26075 591
rect 26041 523 26075 537
rect 26041 503 26075 523
rect 26041 455 26075 465
rect 26041 431 26075 455
rect 26041 387 26075 393
rect 26041 359 26075 387
rect 26041 319 26075 321
rect 26041 287 26075 319
rect 26041 217 26075 249
rect 26041 215 26075 217
rect 26041 149 26075 177
rect 26041 143 26075 149
rect 26041 81 26075 105
rect 26041 71 26075 81
rect 26041 13 26075 33
rect 26041 -1 26075 13
rect 26041 -55 26075 -39
rect 26041 -73 26075 -55
rect 26041 -123 26075 -111
rect 26041 -145 26075 -123
rect 26041 -191 26075 -183
rect 26041 -217 26075 -191
rect 26041 -259 26075 -255
rect 26041 -289 26075 -259
rect 26041 -361 26075 -327
rect 26041 -429 26075 -399
rect 26041 -433 26075 -429
rect 26041 -497 26075 -471
rect 26041 -505 26075 -497
rect 26041 -565 26075 -543
rect 26041 -577 26075 -565
rect 26041 -633 26075 -615
rect 26041 -649 26075 -633
rect 26041 -701 26075 -687
rect 26041 -721 26075 -701
rect 26041 -769 26075 -759
rect 26041 -793 26075 -769
rect 26041 -837 26075 -831
rect 26041 -865 26075 -837
rect 26041 -905 26075 -903
rect 26041 -937 26075 -905
rect 26041 -1007 26075 -975
rect 26041 -1009 26075 -1007
rect 26041 -1075 26075 -1047
rect 26041 -1081 26075 -1075
rect 26041 -1143 26075 -1119
rect 26041 -1153 26075 -1143
rect 26041 -1211 26075 -1191
rect 26041 -1225 26075 -1211
rect 26041 -1279 26075 -1263
rect 26041 -1297 26075 -1279
rect 26041 -1347 26075 -1335
rect 26041 -1369 26075 -1347
rect 31385 1883 31419 1905
rect 31385 1871 31419 1883
rect 31385 1815 31419 1833
rect 31385 1799 31419 1815
rect 31385 1747 31419 1761
rect 31385 1727 31419 1747
rect 31385 1679 31419 1689
rect 31385 1655 31419 1679
rect 31385 1611 31419 1617
rect 31385 1583 31419 1611
rect 31385 1543 31419 1545
rect 31385 1511 31419 1543
rect 31385 1441 31419 1473
rect 31385 1439 31419 1441
rect 31385 1373 31419 1401
rect 31385 1367 31419 1373
rect 31385 1305 31419 1329
rect 31385 1295 31419 1305
rect 31385 1237 31419 1257
rect 31385 1223 31419 1237
rect 31385 1169 31419 1185
rect 31385 1151 31419 1169
rect 31385 1101 31419 1113
rect 31385 1079 31419 1101
rect 31385 1033 31419 1041
rect 31385 1007 31419 1033
rect 31385 965 31419 969
rect 31385 935 31419 965
rect 31385 863 31419 897
rect 31385 795 31419 825
rect 31385 791 31419 795
rect 31385 727 31419 753
rect 31385 719 31419 727
rect 31385 659 31419 681
rect 31385 647 31419 659
rect 31385 591 31419 609
rect 31385 575 31419 591
rect 31385 523 31419 537
rect 31385 503 31419 523
rect 31385 455 31419 465
rect 31385 431 31419 455
rect 31385 387 31419 393
rect 31385 359 31419 387
rect 31385 319 31419 321
rect 31385 287 31419 319
rect 31385 217 31419 249
rect 31385 215 31419 217
rect 31385 149 31419 177
rect 31385 143 31419 149
rect 31385 81 31419 105
rect 31385 71 31419 81
rect 31385 13 31419 33
rect 31385 -1 31419 13
rect 31385 -55 31419 -39
rect 31385 -73 31419 -55
rect 31385 -123 31419 -111
rect 31385 -145 31419 -123
rect 31385 -191 31419 -183
rect 31385 -217 31419 -191
rect 31385 -259 31419 -255
rect 31385 -289 31419 -259
rect 31385 -361 31419 -327
rect 31385 -429 31419 -399
rect 31385 -433 31419 -429
rect 31385 -497 31419 -471
rect 31385 -505 31419 -497
rect 31385 -565 31419 -543
rect 31385 -577 31419 -565
rect 31385 -633 31419 -615
rect 31385 -649 31419 -633
rect 31385 -701 31419 -687
rect 31385 -721 31419 -701
rect 31385 -769 31419 -759
rect 31385 -793 31419 -769
rect 31385 -837 31419 -831
rect 31385 -865 31419 -837
rect 31385 -905 31419 -903
rect 31385 -937 31419 -905
rect 31385 -1007 31419 -975
rect 31385 -1009 31419 -1007
rect 31385 -1075 31419 -1047
rect 31385 -1081 31419 -1075
rect 31385 -1143 31419 -1119
rect 31385 -1153 31419 -1143
rect 31385 -1211 31419 -1191
rect 31385 -1225 31419 -1211
rect 31385 -1279 31419 -1263
rect 31385 -1297 31419 -1279
rect 31385 -1347 31419 -1335
rect 31385 -1369 31419 -1347
rect 26121 -1625 26155 -1591
rect 26193 -1625 26197 -1591
rect 26197 -1625 26227 -1591
rect 26265 -1625 26299 -1591
rect 26337 -1625 26367 -1591
rect 26367 -1625 26371 -1591
rect 26409 -1625 26435 -1591
rect 26435 -1625 26443 -1591
rect 26481 -1625 26503 -1591
rect 26503 -1625 26515 -1591
rect 26553 -1625 26571 -1591
rect 26571 -1625 26587 -1591
rect 26625 -1625 26639 -1591
rect 26639 -1625 26659 -1591
rect 26697 -1625 26707 -1591
rect 26707 -1625 26731 -1591
rect 26769 -1625 26775 -1591
rect 26775 -1625 26803 -1591
rect 26841 -1625 26843 -1591
rect 26843 -1625 26875 -1591
rect 26913 -1625 26945 -1591
rect 26945 -1625 26947 -1591
rect 26985 -1625 27013 -1591
rect 27013 -1625 27019 -1591
rect 27057 -1625 27081 -1591
rect 27081 -1625 27091 -1591
rect 27129 -1625 27149 -1591
rect 27149 -1625 27163 -1591
rect 27201 -1625 27217 -1591
rect 27217 -1625 27235 -1591
rect 27273 -1625 27285 -1591
rect 27285 -1625 27307 -1591
rect 27345 -1625 27353 -1591
rect 27353 -1625 27379 -1591
rect 27417 -1625 27421 -1591
rect 27421 -1625 27451 -1591
rect 27489 -1625 27523 -1591
rect 27561 -1625 27591 -1591
rect 27591 -1625 27595 -1591
rect 27633 -1625 27659 -1591
rect 27659 -1625 27667 -1591
rect 27705 -1625 27727 -1591
rect 27727 -1625 27739 -1591
rect 27777 -1625 27795 -1591
rect 27795 -1625 27811 -1591
rect 27849 -1625 27863 -1591
rect 27863 -1625 27883 -1591
rect 27921 -1625 27931 -1591
rect 27931 -1625 27955 -1591
rect 27993 -1625 27999 -1591
rect 27999 -1625 28027 -1591
rect 28065 -1625 28067 -1591
rect 28067 -1625 28099 -1591
rect 28137 -1625 28169 -1591
rect 28169 -1625 28171 -1591
rect 28209 -1625 28237 -1591
rect 28237 -1625 28243 -1591
rect 28281 -1625 28305 -1591
rect 28305 -1625 28315 -1591
rect 28353 -1625 28373 -1591
rect 28373 -1625 28387 -1591
rect 28425 -1625 28441 -1591
rect 28441 -1625 28459 -1591
rect 28497 -1625 28509 -1591
rect 28509 -1625 28531 -1591
rect 28569 -1625 28577 -1591
rect 28577 -1625 28603 -1591
rect 28641 -1625 28645 -1591
rect 28645 -1625 28675 -1591
rect 28713 -1625 28747 -1591
rect 28785 -1625 28815 -1591
rect 28815 -1625 28819 -1591
rect 28857 -1625 28883 -1591
rect 28883 -1625 28891 -1591
rect 28929 -1625 28951 -1591
rect 28951 -1625 28963 -1591
rect 29001 -1625 29019 -1591
rect 29019 -1625 29035 -1591
rect 29073 -1625 29087 -1591
rect 29087 -1625 29107 -1591
rect 29145 -1625 29155 -1591
rect 29155 -1625 29179 -1591
rect 29217 -1625 29223 -1591
rect 29223 -1625 29251 -1591
rect 29289 -1625 29291 -1591
rect 29291 -1625 29323 -1591
rect 29361 -1625 29393 -1591
rect 29393 -1625 29395 -1591
rect 29433 -1625 29461 -1591
rect 29461 -1625 29467 -1591
rect 29505 -1625 29529 -1591
rect 29529 -1625 29539 -1591
rect 29577 -1625 29597 -1591
rect 29597 -1625 29611 -1591
rect 29649 -1625 29665 -1591
rect 29665 -1625 29683 -1591
rect 29721 -1625 29733 -1591
rect 29733 -1625 29755 -1591
rect 29793 -1625 29801 -1591
rect 29801 -1625 29827 -1591
rect 29865 -1625 29869 -1591
rect 29869 -1625 29899 -1591
rect 29937 -1625 29971 -1591
rect 30009 -1625 30039 -1591
rect 30039 -1625 30043 -1591
rect 30081 -1625 30107 -1591
rect 30107 -1625 30115 -1591
rect 30153 -1625 30175 -1591
rect 30175 -1625 30187 -1591
rect 30225 -1625 30243 -1591
rect 30243 -1625 30259 -1591
rect 30297 -1625 30311 -1591
rect 30311 -1625 30331 -1591
rect 30369 -1625 30379 -1591
rect 30379 -1625 30403 -1591
rect 30441 -1625 30447 -1591
rect 30447 -1625 30475 -1591
rect 30513 -1625 30515 -1591
rect 30515 -1625 30547 -1591
rect 30585 -1625 30617 -1591
rect 30617 -1625 30619 -1591
rect 30657 -1625 30685 -1591
rect 30685 -1625 30691 -1591
rect 30729 -1625 30753 -1591
rect 30753 -1625 30763 -1591
rect 30801 -1625 30821 -1591
rect 30821 -1625 30835 -1591
rect 30873 -1625 30889 -1591
rect 30889 -1625 30907 -1591
rect 30945 -1625 30957 -1591
rect 30957 -1625 30979 -1591
rect 31017 -1625 31025 -1591
rect 31025 -1625 31051 -1591
rect 31089 -1625 31093 -1591
rect 31093 -1625 31123 -1591
rect 31161 -1625 31195 -1591
rect 31233 -1625 31263 -1591
rect 31263 -1625 31267 -1591
rect 31305 -1625 31339 -1591
<< metal1 >>
rect 15420 4277 24456 4316
rect 15420 4243 15529 4277
rect 15563 4243 15601 4277
rect 15635 4243 15673 4277
rect 15707 4243 15745 4277
rect 15779 4243 15817 4277
rect 15851 4243 15889 4277
rect 15923 4243 15961 4277
rect 15995 4243 16033 4277
rect 16067 4243 16105 4277
rect 16139 4243 16177 4277
rect 16211 4243 16249 4277
rect 16283 4243 16321 4277
rect 16355 4243 16393 4277
rect 16427 4243 16465 4277
rect 16499 4243 16537 4277
rect 16571 4243 16609 4277
rect 16643 4243 16681 4277
rect 16715 4243 16753 4277
rect 16787 4243 16825 4277
rect 16859 4243 16897 4277
rect 16931 4243 16969 4277
rect 17003 4243 17041 4277
rect 17075 4243 17113 4277
rect 17147 4243 17185 4277
rect 17219 4243 17257 4277
rect 17291 4243 17329 4277
rect 17363 4243 17401 4277
rect 17435 4243 17473 4277
rect 17507 4243 17545 4277
rect 17579 4243 17617 4277
rect 17651 4243 17689 4277
rect 17723 4243 17761 4277
rect 17795 4243 17833 4277
rect 17867 4243 17905 4277
rect 17939 4243 17977 4277
rect 18011 4243 18049 4277
rect 18083 4243 18121 4277
rect 18155 4243 18193 4277
rect 18227 4243 18265 4277
rect 18299 4243 18337 4277
rect 18371 4243 18409 4277
rect 18443 4243 18481 4277
rect 18515 4243 18553 4277
rect 18587 4243 18625 4277
rect 18659 4243 18697 4277
rect 18731 4243 18769 4277
rect 18803 4243 18841 4277
rect 18875 4243 18913 4277
rect 18947 4243 18985 4277
rect 19019 4243 19057 4277
rect 19091 4243 19129 4277
rect 19163 4243 19201 4277
rect 19235 4243 19273 4277
rect 19307 4243 19345 4277
rect 19379 4243 19417 4277
rect 19451 4243 19489 4277
rect 19523 4243 19561 4277
rect 19595 4243 19633 4277
rect 19667 4243 19705 4277
rect 19739 4243 19777 4277
rect 19811 4243 19849 4277
rect 19883 4243 19921 4277
rect 19955 4243 19993 4277
rect 20027 4243 20065 4277
rect 20099 4243 20137 4277
rect 20171 4243 20209 4277
rect 20243 4243 20281 4277
rect 20315 4243 20353 4277
rect 20387 4243 20425 4277
rect 20459 4243 20497 4277
rect 20531 4243 20569 4277
rect 20603 4243 20641 4277
rect 20675 4243 20713 4277
rect 20747 4243 20785 4277
rect 20819 4243 20857 4277
rect 20891 4243 20929 4277
rect 20963 4243 21001 4277
rect 21035 4243 21073 4277
rect 21107 4243 21145 4277
rect 21179 4243 21217 4277
rect 21251 4243 21289 4277
rect 21323 4243 21361 4277
rect 21395 4243 21433 4277
rect 21467 4243 21505 4277
rect 21539 4243 21577 4277
rect 21611 4243 21649 4277
rect 21683 4243 21721 4277
rect 21755 4243 21793 4277
rect 21827 4243 21865 4277
rect 21899 4243 21937 4277
rect 21971 4243 22009 4277
rect 22043 4243 22081 4277
rect 22115 4243 22153 4277
rect 22187 4243 22225 4277
rect 22259 4243 22297 4277
rect 22331 4243 22369 4277
rect 22403 4243 22441 4277
rect 22475 4243 22513 4277
rect 22547 4243 22585 4277
rect 22619 4243 22657 4277
rect 22691 4243 22729 4277
rect 22763 4243 22801 4277
rect 22835 4243 22873 4277
rect 22907 4243 22945 4277
rect 22979 4243 23017 4277
rect 23051 4243 23089 4277
rect 23123 4243 23161 4277
rect 23195 4243 23233 4277
rect 23267 4243 23305 4277
rect 23339 4243 23377 4277
rect 23411 4243 23449 4277
rect 23483 4243 23521 4277
rect 23555 4243 23593 4277
rect 23627 4243 23665 4277
rect 23699 4243 23737 4277
rect 23771 4243 23809 4277
rect 23843 4243 23881 4277
rect 23915 4243 23953 4277
rect 23987 4243 24025 4277
rect 24059 4243 24097 4277
rect 24131 4243 24169 4277
rect 24203 4243 24241 4277
rect 24275 4243 24313 4277
rect 24347 4243 24456 4277
rect 15420 4204 24456 4243
rect 15420 4176 15924 4204
rect 15420 4111 15537 4176
rect 15420 4077 15459 4111
rect 15493 4077 15537 4111
rect 15420 4039 15537 4077
rect 15420 4005 15459 4039
rect 15493 4005 15537 4039
rect 15420 3967 15537 4005
rect 15420 3933 15459 3967
rect 15493 3933 15537 3967
rect 15420 3932 15537 3933
rect 15909 3932 15924 4176
rect 15420 3904 15924 3932
rect 23656 4176 24456 4204
rect 23656 3932 23691 4176
rect 24319 4111 24456 4176
rect 24319 4077 24383 4111
rect 24417 4077 24456 4111
rect 24319 4039 24456 4077
rect 24319 4005 24383 4039
rect 24417 4005 24456 4039
rect 24319 3967 24456 4005
rect 24319 3933 24383 3967
rect 24417 3933 24456 3967
rect 24319 3932 24456 3933
rect 23656 3904 24456 3932
rect 15420 3895 15532 3904
rect 15420 3861 15459 3895
rect 15493 3861 15532 3895
rect 15420 3823 15532 3861
rect 15420 3789 15459 3823
rect 15493 3789 15532 3823
rect 15420 3751 15532 3789
rect 24344 3895 24456 3904
rect 24344 3861 24383 3895
rect 24417 3861 24456 3895
rect 24344 3823 24456 3861
rect 24344 3789 24383 3823
rect 24417 3789 24456 3823
rect 15420 3717 15459 3751
rect 15493 3717 15532 3751
rect 15420 3679 15532 3717
rect 15420 3645 15459 3679
rect 15493 3645 15532 3679
rect 15420 3607 15532 3645
rect 17550 3709 22522 3756
rect 17550 3657 17622 3709
rect 17674 3657 18202 3709
rect 18254 3657 18802 3709
rect 18854 3657 19402 3709
rect 19454 3657 20002 3709
rect 20054 3657 20602 3709
rect 20654 3657 21202 3709
rect 21254 3657 21802 3709
rect 21854 3657 22402 3709
rect 22454 3657 22522 3709
rect 17550 3612 22522 3657
rect 24344 3751 24456 3789
rect 24344 3717 24383 3751
rect 24417 3717 24456 3751
rect 24344 3679 24456 3717
rect 24344 3645 24383 3679
rect 24417 3645 24456 3679
rect 15420 3573 15459 3607
rect 15493 3573 15532 3607
rect 15420 3535 15532 3573
rect 15420 3501 15459 3535
rect 15493 3501 15532 3535
rect 15420 3463 15532 3501
rect 15420 3429 15459 3463
rect 15493 3429 15532 3463
rect 15420 3391 15532 3429
rect 15420 3357 15459 3391
rect 15493 3357 15532 3391
rect 15420 3319 15532 3357
rect 15420 3285 15459 3319
rect 15493 3285 15532 3319
rect 15420 3247 15532 3285
rect 15420 3213 15459 3247
rect 15493 3213 15532 3247
rect 15420 3175 15532 3213
rect 17614 3202 17674 3612
rect 17854 3282 17914 3612
rect 18304 3444 21580 3448
rect 18304 3392 21518 3444
rect 21570 3392 21580 3444
rect 18304 3388 21580 3392
rect 18304 3282 18364 3388
rect 18766 3292 18826 3388
rect 19220 3286 19280 3388
rect 19682 3286 19742 3388
rect 20136 3286 20196 3388
rect 20586 3292 20646 3388
rect 21052 3298 21112 3388
rect 21508 3292 21568 3388
rect 21742 3204 21802 3612
rect 21968 3280 22028 3612
rect 15420 3141 15459 3175
rect 15493 3141 15532 3175
rect 15420 3103 15532 3141
rect 15420 3069 15459 3103
rect 15493 3069 15532 3103
rect 15420 3031 15532 3069
rect 15420 2997 15459 3031
rect 15493 2997 15532 3031
rect 15420 2959 15532 2997
rect 15420 2925 15459 2959
rect 15493 2925 15532 2959
rect 15420 2887 15532 2925
rect 15420 2853 15459 2887
rect 15493 2853 15532 2887
rect 15420 2815 15532 2853
rect 15420 2781 15459 2815
rect 15493 2781 15532 2815
rect 15420 2743 15532 2781
rect 15420 2709 15459 2743
rect 15493 2709 15532 2743
rect 15420 2616 15532 2709
rect 17622 2616 17682 3076
rect 17850 2616 17910 3006
rect 18078 2764 18138 3084
rect 18310 2894 18376 3006
rect 18772 2894 18838 3006
rect 19226 2894 19292 3006
rect 19688 2894 19754 3006
rect 20142 2894 20208 3006
rect 20592 2894 20658 3006
rect 21058 2894 21124 3006
rect 21514 2894 21580 3006
rect 18310 2828 21580 2894
rect 18078 2712 18082 2764
rect 18134 2712 18138 2764
rect 18078 2702 18138 2712
rect 21748 2616 21808 3076
rect 21976 2616 22036 3008
rect 22208 2616 22268 3612
rect 24344 3607 24456 3645
rect 24344 3573 24383 3607
rect 24417 3573 24456 3607
rect 24344 3535 24456 3573
rect 24344 3501 24383 3535
rect 24417 3501 24456 3535
rect 24344 3463 24456 3501
rect 24344 3429 24383 3463
rect 24417 3429 24456 3463
rect 24344 3391 24456 3429
rect 24344 3357 24383 3391
rect 24417 3357 24456 3391
rect 24344 3319 24456 3357
rect 24344 3285 24383 3319
rect 24417 3285 24456 3319
rect 24344 3247 24456 3285
rect 24344 3213 24383 3247
rect 24417 3213 24456 3247
rect 24344 3175 24456 3213
rect 24344 3141 24383 3175
rect 24417 3141 24456 3175
rect 24344 3103 24456 3141
rect 24344 3069 24383 3103
rect 24417 3069 24456 3103
rect 24344 3031 24456 3069
rect 24344 2997 24383 3031
rect 24417 2997 24456 3031
rect 24344 2959 24456 2997
rect 24344 2925 24383 2959
rect 24417 2925 24456 2959
rect 24344 2887 24456 2925
rect 24344 2853 24383 2887
rect 24417 2853 24456 2887
rect 24344 2815 24456 2853
rect 24344 2781 24383 2815
rect 24417 2781 24456 2815
rect 24344 2743 24456 2781
rect 24344 2709 24383 2743
rect 24417 2709 24456 2743
rect 24344 2616 24456 2709
rect 15420 2577 24456 2616
rect 15420 2543 15529 2577
rect 15563 2543 15601 2577
rect 15635 2543 15673 2577
rect 15707 2543 15745 2577
rect 15779 2543 15817 2577
rect 15851 2543 15889 2577
rect 15923 2543 15961 2577
rect 15995 2543 16033 2577
rect 16067 2543 16105 2577
rect 16139 2543 16177 2577
rect 16211 2543 16249 2577
rect 16283 2543 16321 2577
rect 16355 2543 16393 2577
rect 16427 2543 16465 2577
rect 16499 2543 16537 2577
rect 16571 2543 16609 2577
rect 16643 2543 16681 2577
rect 16715 2543 16753 2577
rect 16787 2543 16825 2577
rect 16859 2543 16897 2577
rect 16931 2543 16969 2577
rect 17003 2543 17041 2577
rect 17075 2543 17113 2577
rect 17147 2543 17185 2577
rect 17219 2543 17257 2577
rect 17291 2543 17329 2577
rect 17363 2543 17401 2577
rect 17435 2543 17473 2577
rect 17507 2543 17545 2577
rect 17579 2543 17617 2577
rect 17651 2543 17689 2577
rect 17723 2543 17761 2577
rect 17795 2543 17833 2577
rect 17867 2543 17905 2577
rect 17939 2543 17977 2577
rect 18011 2543 18049 2577
rect 18083 2543 18121 2577
rect 18155 2543 18193 2577
rect 18227 2543 18265 2577
rect 18299 2543 18337 2577
rect 18371 2543 18409 2577
rect 18443 2543 18481 2577
rect 18515 2543 18553 2577
rect 18587 2543 18625 2577
rect 18659 2543 18697 2577
rect 18731 2543 18769 2577
rect 18803 2543 18841 2577
rect 18875 2543 18913 2577
rect 18947 2543 18985 2577
rect 19019 2543 19057 2577
rect 19091 2543 19129 2577
rect 19163 2543 19201 2577
rect 19235 2543 19273 2577
rect 19307 2543 19345 2577
rect 19379 2543 19417 2577
rect 19451 2543 19489 2577
rect 19523 2543 19561 2577
rect 19595 2543 19633 2577
rect 19667 2543 19705 2577
rect 19739 2543 19777 2577
rect 19811 2543 19849 2577
rect 19883 2543 19921 2577
rect 19955 2543 19993 2577
rect 20027 2543 20065 2577
rect 20099 2543 20137 2577
rect 20171 2543 20209 2577
rect 20243 2543 20281 2577
rect 20315 2543 20353 2577
rect 20387 2543 20425 2577
rect 20459 2543 20497 2577
rect 20531 2543 20569 2577
rect 20603 2543 20641 2577
rect 20675 2543 20713 2577
rect 20747 2543 20785 2577
rect 20819 2543 20857 2577
rect 20891 2543 20929 2577
rect 20963 2543 21001 2577
rect 21035 2543 21073 2577
rect 21107 2543 21145 2577
rect 21179 2543 21217 2577
rect 21251 2543 21289 2577
rect 21323 2543 21361 2577
rect 21395 2543 21433 2577
rect 21467 2543 21505 2577
rect 21539 2543 21577 2577
rect 21611 2543 21649 2577
rect 21683 2543 21721 2577
rect 21755 2543 21793 2577
rect 21827 2543 21865 2577
rect 21899 2543 21937 2577
rect 21971 2543 22009 2577
rect 22043 2543 22081 2577
rect 22115 2543 22153 2577
rect 22187 2543 22225 2577
rect 22259 2543 22297 2577
rect 22331 2543 22369 2577
rect 22403 2543 22441 2577
rect 22475 2543 22513 2577
rect 22547 2543 22585 2577
rect 22619 2543 22657 2577
rect 22691 2543 22729 2577
rect 22763 2543 22801 2577
rect 22835 2543 22873 2577
rect 22907 2543 22945 2577
rect 22979 2543 23017 2577
rect 23051 2543 23089 2577
rect 23123 2543 23161 2577
rect 23195 2543 23233 2577
rect 23267 2543 23305 2577
rect 23339 2543 23377 2577
rect 23411 2543 23449 2577
rect 23483 2543 23521 2577
rect 23555 2543 23593 2577
rect 23627 2543 23665 2577
rect 23699 2543 23737 2577
rect 23771 2543 23809 2577
rect 23843 2543 23881 2577
rect 23915 2543 23953 2577
rect 23987 2543 24025 2577
rect 24059 2543 24097 2577
rect 24131 2543 24169 2577
rect 24203 2543 24241 2577
rect 24275 2543 24313 2577
rect 24347 2543 24456 2577
rect 15420 2504 24456 2543
rect 26002 4277 31458 4316
rect 26002 4243 26121 4277
rect 26155 4243 26193 4277
rect 26227 4243 26265 4277
rect 26299 4243 26337 4277
rect 26371 4243 26409 4277
rect 26443 4243 26481 4277
rect 26515 4243 26553 4277
rect 26587 4243 26625 4277
rect 26659 4243 26697 4277
rect 26731 4243 26769 4277
rect 26803 4243 26841 4277
rect 26875 4243 26913 4277
rect 26947 4243 26985 4277
rect 27019 4243 27057 4277
rect 27091 4243 27129 4277
rect 27163 4243 27201 4277
rect 27235 4243 27273 4277
rect 27307 4243 27345 4277
rect 27379 4243 27417 4277
rect 27451 4243 27489 4277
rect 27523 4243 27561 4277
rect 27595 4243 27633 4277
rect 27667 4243 27705 4277
rect 27739 4243 27777 4277
rect 27811 4243 27849 4277
rect 27883 4243 27921 4277
rect 27955 4243 27993 4277
rect 28027 4243 28065 4277
rect 28099 4243 28137 4277
rect 28171 4243 28209 4277
rect 28243 4243 28281 4277
rect 28315 4243 28353 4277
rect 28387 4243 28425 4277
rect 28459 4243 28497 4277
rect 28531 4243 28569 4277
rect 28603 4243 28641 4277
rect 28675 4243 28713 4277
rect 28747 4243 28785 4277
rect 28819 4243 28857 4277
rect 28891 4243 28929 4277
rect 28963 4243 29001 4277
rect 29035 4243 29073 4277
rect 29107 4243 29145 4277
rect 29179 4243 29217 4277
rect 29251 4243 29289 4277
rect 29323 4243 29361 4277
rect 29395 4243 29433 4277
rect 29467 4243 29505 4277
rect 29539 4243 29577 4277
rect 29611 4243 29649 4277
rect 29683 4243 29721 4277
rect 29755 4243 29793 4277
rect 29827 4243 29865 4277
rect 29899 4243 29937 4277
rect 29971 4243 30009 4277
rect 30043 4243 30081 4277
rect 30115 4243 30153 4277
rect 30187 4243 30225 4277
rect 30259 4243 30297 4277
rect 30331 4243 30369 4277
rect 30403 4243 30441 4277
rect 30475 4243 30513 4277
rect 30547 4243 30585 4277
rect 30619 4243 30657 4277
rect 30691 4243 30729 4277
rect 30763 4243 30801 4277
rect 30835 4243 30873 4277
rect 30907 4243 30945 4277
rect 30979 4243 31017 4277
rect 31051 4243 31089 4277
rect 31123 4243 31161 4277
rect 31195 4243 31233 4277
rect 31267 4243 31305 4277
rect 31339 4243 31458 4277
rect 26002 4204 31458 4243
rect 26002 4176 26724 4204
rect 26002 4107 26132 4176
rect 26002 4073 26041 4107
rect 26075 4073 26132 4107
rect 26002 4035 26132 4073
rect 26002 4001 26041 4035
rect 26075 4001 26132 4035
rect 26002 3963 26132 4001
rect 26002 3929 26041 3963
rect 26075 3932 26132 3963
rect 26696 3932 26724 4176
rect 26075 3929 26724 3932
rect 26002 3904 26724 3929
rect 30736 4176 31458 4204
rect 30736 3932 30764 4176
rect 31328 4107 31458 4176
rect 31328 4073 31385 4107
rect 31419 4073 31458 4107
rect 31328 4035 31458 4073
rect 31328 4001 31385 4035
rect 31419 4001 31458 4035
rect 31328 3963 31458 4001
rect 31328 3932 31385 3963
rect 30736 3929 31385 3932
rect 31419 3929 31458 3963
rect 30736 3904 31458 3929
rect 26002 3891 26114 3904
rect 26002 3857 26041 3891
rect 26075 3857 26114 3891
rect 26002 3819 26114 3857
rect 26002 3785 26041 3819
rect 26075 3785 26114 3819
rect 26002 3747 26114 3785
rect 31346 3891 31458 3904
rect 31346 3857 31385 3891
rect 31419 3857 31458 3891
rect 31346 3819 31458 3857
rect 31346 3785 31385 3819
rect 31419 3785 31458 3819
rect 26002 3713 26041 3747
rect 26075 3713 26114 3747
rect 26002 3675 26114 3713
rect 26002 3641 26041 3675
rect 26075 3641 26114 3675
rect 26002 3603 26114 3641
rect 26312 3709 31284 3756
rect 26312 3657 26384 3709
rect 26436 3657 26964 3709
rect 27016 3657 27564 3709
rect 27616 3657 28164 3709
rect 28216 3657 28764 3709
rect 28816 3657 29364 3709
rect 29416 3657 29964 3709
rect 30016 3657 30564 3709
rect 30616 3657 31164 3709
rect 31216 3657 31284 3709
rect 26312 3612 31284 3657
rect 31346 3747 31458 3785
rect 31346 3713 31385 3747
rect 31419 3713 31458 3747
rect 31346 3675 31458 3713
rect 31346 3641 31385 3675
rect 31419 3641 31458 3675
rect 26002 3569 26041 3603
rect 26075 3569 26114 3603
rect 26002 3531 26114 3569
rect 26002 3497 26041 3531
rect 26075 3497 26114 3531
rect 26002 3459 26114 3497
rect 26002 3425 26041 3459
rect 26075 3425 26114 3459
rect 26002 3387 26114 3425
rect 26002 3353 26041 3387
rect 26075 3353 26114 3387
rect 26002 3315 26114 3353
rect 26002 3281 26041 3315
rect 26075 3281 26114 3315
rect 26002 3243 26114 3281
rect 26002 3209 26041 3243
rect 26075 3209 26114 3243
rect 26002 3171 26114 3209
rect 26376 3202 26436 3612
rect 26616 3282 26676 3612
rect 26002 3137 26041 3171
rect 26075 3137 26114 3171
rect 26002 3099 26114 3137
rect 26002 3065 26041 3099
rect 26075 3065 26114 3099
rect 26002 3027 26114 3065
rect 26002 2993 26041 3027
rect 26075 2993 26114 3027
rect 26002 2955 26114 2993
rect 26002 2921 26041 2955
rect 26075 2921 26114 2955
rect 26002 2883 26114 2921
rect 26002 2849 26041 2883
rect 26075 2849 26114 2883
rect 26002 2811 26114 2849
rect 26002 2777 26041 2811
rect 26075 2777 26114 2811
rect 26002 2739 26114 2777
rect 26002 2705 26041 2739
rect 26075 2705 26114 2739
rect 26002 2667 26114 2705
rect 26002 2633 26041 2667
rect 26075 2633 26114 2667
rect 26002 2536 26114 2633
rect 26384 2536 26444 3076
rect 26612 2536 26672 3006
rect 26840 2536 26900 3612
rect 27066 3388 30330 3448
rect 27066 3282 27126 3388
rect 27528 3292 27588 3388
rect 27982 3286 28042 3388
rect 28444 3286 28504 3388
rect 28898 3286 28958 3388
rect 29348 3292 29408 3388
rect 29814 3298 29874 3388
rect 30270 3292 30330 3388
rect 30730 3280 30790 3612
rect 27066 2894 27126 3002
rect 27528 2894 27588 3004
rect 27982 2896 28042 3004
rect 27976 2894 28048 2896
rect 28444 2894 28504 3006
rect 28898 2894 28958 3006
rect 29348 2894 29408 3006
rect 29814 2894 29874 3002
rect 30270 2894 30330 3006
rect 27059 2892 30337 2894
rect 27059 2890 27986 2892
rect 27059 2838 27070 2890
rect 27122 2838 27532 2890
rect 27584 2840 27986 2890
rect 28038 2890 30337 2892
rect 28038 2840 28448 2890
rect 27584 2838 28448 2840
rect 28500 2838 28902 2890
rect 28954 2838 29352 2890
rect 29404 2838 29818 2890
rect 29870 2838 30274 2890
rect 30326 2838 30337 2890
rect 27059 2828 30337 2838
rect 30504 2686 30564 3110
rect 30498 2682 30570 2686
rect 30498 2630 30508 2682
rect 30560 2630 30570 2682
rect 30498 2626 30570 2630
rect 30738 2536 30798 3008
rect 30970 2536 31030 3612
rect 31346 3603 31458 3641
rect 31346 3569 31385 3603
rect 31419 3569 31458 3603
rect 31346 3531 31458 3569
rect 31346 3497 31385 3531
rect 31419 3497 31458 3531
rect 31346 3459 31458 3497
rect 31346 3425 31385 3459
rect 31419 3425 31458 3459
rect 31346 3387 31458 3425
rect 31346 3353 31385 3387
rect 31419 3353 31458 3387
rect 31346 3315 31458 3353
rect 31346 3281 31385 3315
rect 31419 3281 31458 3315
rect 31346 3243 31458 3281
rect 31346 3209 31385 3243
rect 31419 3209 31458 3243
rect 31346 3171 31458 3209
rect 31346 3137 31385 3171
rect 31419 3137 31458 3171
rect 31346 3099 31458 3137
rect 31346 3065 31385 3099
rect 31419 3065 31458 3099
rect 31346 3027 31458 3065
rect 31346 2993 31385 3027
rect 31419 2993 31458 3027
rect 31346 2955 31458 2993
rect 31346 2921 31385 2955
rect 31419 2921 31458 2955
rect 31346 2883 31458 2921
rect 31346 2849 31385 2883
rect 31419 2849 31458 2883
rect 31346 2811 31458 2849
rect 31346 2777 31385 2811
rect 31419 2777 31458 2811
rect 31346 2739 31458 2777
rect 31346 2705 31385 2739
rect 31419 2705 31458 2739
rect 31346 2667 31458 2705
rect 31346 2633 31385 2667
rect 31419 2633 31458 2667
rect 31346 2538 31458 2633
rect 31346 2536 31542 2538
rect 26002 2497 31542 2536
rect 26002 2463 26121 2497
rect 26155 2463 26193 2497
rect 26227 2463 26265 2497
rect 26299 2463 26337 2497
rect 26371 2463 26409 2497
rect 26443 2463 26481 2497
rect 26515 2463 26553 2497
rect 26587 2463 26625 2497
rect 26659 2463 26697 2497
rect 26731 2463 26769 2497
rect 26803 2463 26841 2497
rect 26875 2463 26913 2497
rect 26947 2463 26985 2497
rect 27019 2463 27057 2497
rect 27091 2463 27129 2497
rect 27163 2463 27201 2497
rect 27235 2463 27273 2497
rect 27307 2463 27345 2497
rect 27379 2463 27417 2497
rect 27451 2463 27489 2497
rect 27523 2463 27561 2497
rect 27595 2463 27633 2497
rect 27667 2463 27705 2497
rect 27739 2463 27777 2497
rect 27811 2463 27849 2497
rect 27883 2463 27921 2497
rect 27955 2463 27993 2497
rect 28027 2463 28065 2497
rect 28099 2463 28137 2497
rect 28171 2463 28209 2497
rect 28243 2463 28281 2497
rect 28315 2463 28353 2497
rect 28387 2463 28425 2497
rect 28459 2463 28497 2497
rect 28531 2463 28569 2497
rect 28603 2463 28641 2497
rect 28675 2463 28713 2497
rect 28747 2463 28785 2497
rect 28819 2463 28857 2497
rect 28891 2463 28929 2497
rect 28963 2463 29001 2497
rect 29035 2463 29073 2497
rect 29107 2463 29145 2497
rect 29179 2463 29217 2497
rect 29251 2463 29289 2497
rect 29323 2463 29361 2497
rect 29395 2463 29433 2497
rect 29467 2463 29505 2497
rect 29539 2463 29577 2497
rect 29611 2463 29649 2497
rect 29683 2463 29721 2497
rect 29755 2463 29793 2497
rect 29827 2463 29865 2497
rect 29899 2463 29937 2497
rect 29971 2463 30009 2497
rect 30043 2463 30081 2497
rect 30115 2463 30153 2497
rect 30187 2463 30225 2497
rect 30259 2463 30297 2497
rect 30331 2463 30369 2497
rect 30403 2463 30441 2497
rect 30475 2463 30513 2497
rect 30547 2463 30585 2497
rect 30619 2463 30657 2497
rect 30691 2463 30729 2497
rect 30763 2463 30801 2497
rect 30835 2463 30873 2497
rect 30907 2463 30945 2497
rect 30979 2463 31017 2497
rect 31051 2463 31089 2497
rect 31123 2463 31161 2497
rect 31195 2463 31233 2497
rect 31267 2463 31305 2497
rect 31339 2463 31542 2497
rect 26002 2442 31542 2463
rect 26002 2424 31458 2442
rect 30504 2344 30564 2350
rect 25234 2340 31566 2344
rect 25234 2288 30508 2340
rect 30560 2288 31566 2340
rect 25234 2284 31566 2288
rect 15420 2241 24456 2280
rect 15420 2207 15529 2241
rect 15563 2207 15601 2241
rect 15635 2207 15673 2241
rect 15707 2207 15745 2241
rect 15779 2207 15817 2241
rect 15851 2207 15889 2241
rect 15923 2207 15961 2241
rect 15995 2207 16033 2241
rect 16067 2207 16105 2241
rect 16139 2207 16177 2241
rect 16211 2207 16249 2241
rect 16283 2207 16321 2241
rect 16355 2207 16393 2241
rect 16427 2207 16465 2241
rect 16499 2207 16537 2241
rect 16571 2207 16609 2241
rect 16643 2207 16681 2241
rect 16715 2207 16753 2241
rect 16787 2207 16825 2241
rect 16859 2207 16897 2241
rect 16931 2207 16969 2241
rect 17003 2207 17041 2241
rect 17075 2207 17113 2241
rect 17147 2207 17185 2241
rect 17219 2207 17257 2241
rect 17291 2207 17329 2241
rect 17363 2207 17401 2241
rect 17435 2207 17473 2241
rect 17507 2207 17545 2241
rect 17579 2207 17617 2241
rect 17651 2207 17689 2241
rect 17723 2207 17761 2241
rect 17795 2207 17833 2241
rect 17867 2207 17905 2241
rect 17939 2207 17977 2241
rect 18011 2207 18049 2241
rect 18083 2207 18121 2241
rect 18155 2207 18193 2241
rect 18227 2207 18265 2241
rect 18299 2207 18337 2241
rect 18371 2207 18409 2241
rect 18443 2207 18481 2241
rect 18515 2207 18553 2241
rect 18587 2207 18625 2241
rect 18659 2207 18697 2241
rect 18731 2207 18769 2241
rect 18803 2207 18841 2241
rect 18875 2207 18913 2241
rect 18947 2207 18985 2241
rect 19019 2207 19057 2241
rect 19091 2207 19129 2241
rect 19163 2207 19201 2241
rect 19235 2207 19273 2241
rect 19307 2207 19345 2241
rect 19379 2207 19417 2241
rect 19451 2207 19489 2241
rect 19523 2207 19561 2241
rect 19595 2207 19633 2241
rect 19667 2207 19705 2241
rect 19739 2207 19777 2241
rect 19811 2207 19849 2241
rect 19883 2207 19921 2241
rect 19955 2207 19993 2241
rect 20027 2207 20065 2241
rect 20099 2207 20137 2241
rect 20171 2207 20209 2241
rect 20243 2207 20281 2241
rect 20315 2207 20353 2241
rect 20387 2207 20425 2241
rect 20459 2207 20497 2241
rect 20531 2207 20569 2241
rect 20603 2207 20641 2241
rect 20675 2207 20713 2241
rect 20747 2207 20785 2241
rect 20819 2207 20857 2241
rect 20891 2207 20929 2241
rect 20963 2207 21001 2241
rect 21035 2207 21073 2241
rect 21107 2207 21145 2241
rect 21179 2207 21217 2241
rect 21251 2207 21289 2241
rect 21323 2207 21361 2241
rect 21395 2207 21433 2241
rect 21467 2207 21505 2241
rect 21539 2207 21577 2241
rect 21611 2207 21649 2241
rect 21683 2207 21721 2241
rect 21755 2207 21793 2241
rect 21827 2207 21865 2241
rect 21899 2207 21937 2241
rect 21971 2207 22009 2241
rect 22043 2207 22081 2241
rect 22115 2207 22153 2241
rect 22187 2207 22225 2241
rect 22259 2207 22297 2241
rect 22331 2207 22369 2241
rect 22403 2207 22441 2241
rect 22475 2207 22513 2241
rect 22547 2207 22585 2241
rect 22619 2207 22657 2241
rect 22691 2207 22729 2241
rect 22763 2207 22801 2241
rect 22835 2207 22873 2241
rect 22907 2207 22945 2241
rect 22979 2207 23017 2241
rect 23051 2207 23089 2241
rect 23123 2207 23161 2241
rect 23195 2207 23233 2241
rect 23267 2207 23305 2241
rect 23339 2207 23377 2241
rect 23411 2207 23449 2241
rect 23483 2207 23521 2241
rect 23555 2207 23593 2241
rect 23627 2207 23665 2241
rect 23699 2207 23737 2241
rect 23771 2207 23809 2241
rect 23843 2207 23881 2241
rect 23915 2207 23953 2241
rect 23987 2207 24025 2241
rect 24059 2207 24097 2241
rect 24131 2207 24169 2241
rect 24203 2207 24241 2241
rect 24275 2207 24313 2241
rect 24347 2207 24456 2241
rect 15420 2168 24456 2207
rect 15420 1945 15532 2168
rect 15420 1911 15459 1945
rect 15493 1911 15532 1945
rect 15420 1873 15532 1911
rect 15420 1839 15459 1873
rect 15493 1839 15532 1873
rect 15420 1801 15532 1839
rect 15420 1767 15459 1801
rect 15493 1767 15532 1801
rect 15420 1729 15532 1767
rect 15420 1695 15459 1729
rect 15493 1695 15532 1729
rect 15420 1657 15532 1695
rect 15420 1623 15459 1657
rect 15493 1623 15532 1657
rect 15420 1614 15532 1623
rect 15790 1614 15850 2168
rect 16018 1614 16078 2168
rect 16244 1614 16304 2168
rect 16702 2026 23178 2086
rect 15420 1585 16304 1614
rect 15420 1551 15459 1585
rect 15493 1554 16304 1585
rect 16468 1610 16540 1614
rect 16468 1558 16478 1610
rect 16530 1558 16540 1610
rect 16468 1554 16540 1558
rect 15493 1551 15532 1554
rect 15420 1513 15532 1551
rect 15420 1479 15459 1513
rect 15493 1479 15532 1513
rect 15420 1441 15532 1479
rect 15420 1407 15459 1441
rect 15493 1407 15532 1441
rect 15420 1369 15532 1407
rect 15420 1335 15459 1369
rect 15493 1335 15532 1369
rect 15420 1297 15532 1335
rect 15790 1322 15850 1554
rect 16018 1438 16078 1554
rect 16244 1338 16304 1554
rect 16474 1446 16534 1554
rect 16702 1298 16762 2026
rect 17620 1902 22264 1962
rect 16924 1610 16996 1614
rect 16924 1558 16934 1610
rect 16986 1558 16996 1610
rect 16924 1554 16996 1558
rect 17384 1610 17456 1614
rect 17384 1558 17394 1610
rect 17446 1558 17456 1610
rect 17384 1554 17456 1558
rect 16930 1448 16990 1554
rect 17390 1442 17450 1554
rect 17620 1304 17680 1902
rect 18528 1778 21344 1838
rect 17840 1610 17912 1614
rect 17840 1558 17850 1610
rect 17902 1558 17912 1610
rect 17840 1554 17912 1558
rect 18298 1610 18370 1614
rect 18298 1558 18308 1610
rect 18360 1558 18370 1610
rect 18298 1554 18370 1558
rect 17846 1448 17906 1554
rect 18304 1448 18364 1554
rect 18528 1310 18588 1778
rect 19452 1662 20430 1722
rect 18762 1610 18834 1614
rect 18762 1558 18772 1610
rect 18824 1558 18834 1610
rect 18762 1554 18834 1558
rect 19216 1610 19288 1614
rect 19216 1558 19226 1610
rect 19278 1558 19288 1610
rect 19216 1554 19288 1558
rect 18768 1444 18828 1554
rect 19222 1442 19282 1554
rect 19452 1302 19512 1662
rect 19676 1610 19748 1614
rect 19676 1558 19686 1610
rect 19738 1558 19748 1610
rect 19676 1554 19748 1558
rect 19906 1610 19978 1614
rect 19906 1558 19916 1610
rect 19968 1558 19978 1610
rect 19906 1554 19978 1558
rect 20134 1610 20206 1614
rect 20134 1558 20144 1610
rect 20196 1558 20206 1610
rect 20134 1554 20206 1558
rect 19682 1444 19742 1554
rect 19912 1332 19972 1554
rect 20140 1436 20200 1554
rect 20370 1354 20430 1662
rect 20590 1610 20662 1614
rect 20590 1558 20600 1610
rect 20652 1558 20662 1610
rect 20590 1554 20662 1558
rect 21050 1610 21122 1614
rect 21050 1558 21060 1610
rect 21112 1558 21122 1610
rect 21050 1554 21122 1558
rect 20596 1442 20656 1554
rect 21056 1448 21116 1554
rect 21284 1350 21344 1778
rect 21506 1610 21578 1614
rect 21506 1558 21516 1610
rect 21568 1558 21578 1610
rect 21506 1554 21578 1558
rect 21962 1610 22034 1614
rect 21962 1558 21972 1610
rect 22024 1558 22034 1610
rect 21962 1554 22034 1558
rect 21512 1448 21572 1554
rect 21968 1448 22028 1554
rect 22204 1314 22264 1902
rect 22418 1610 22490 1614
rect 22418 1558 22428 1610
rect 22480 1558 22490 1610
rect 22418 1554 22490 1558
rect 22876 1610 22948 1614
rect 22876 1558 22886 1610
rect 22938 1558 22948 1610
rect 22876 1554 22948 1558
rect 22424 1452 22484 1554
rect 22882 1448 22942 1554
rect 23118 1322 23178 2026
rect 23572 1614 23632 2168
rect 23804 1614 23864 2168
rect 24030 1614 24090 2168
rect 24344 1945 24456 2168
rect 24344 1911 24383 1945
rect 24417 1911 24456 1945
rect 24344 1873 24456 1911
rect 24344 1839 24383 1873
rect 24417 1839 24456 1873
rect 24344 1801 24456 1839
rect 24344 1767 24383 1801
rect 24417 1767 24456 1801
rect 24344 1729 24456 1767
rect 24344 1695 24383 1729
rect 24417 1695 24456 1729
rect 24344 1657 24456 1695
rect 24344 1623 24383 1657
rect 24417 1623 24456 1657
rect 24344 1614 24456 1623
rect 23336 1610 23408 1614
rect 23336 1558 23346 1610
rect 23398 1558 23408 1610
rect 23336 1554 23408 1558
rect 23572 1585 24456 1614
rect 23572 1554 24383 1585
rect 23342 1444 23402 1554
rect 23572 1320 23632 1554
rect 23804 1440 23864 1554
rect 24030 1338 24090 1554
rect 24344 1551 24383 1554
rect 24417 1551 24456 1585
rect 24344 1513 24456 1551
rect 24344 1479 24383 1513
rect 24417 1479 24456 1513
rect 24344 1441 24456 1479
rect 24344 1407 24383 1441
rect 24417 1407 24456 1441
rect 24344 1369 24456 1407
rect 24344 1335 24383 1369
rect 24417 1335 24456 1369
rect 15420 1263 15459 1297
rect 15493 1263 15532 1297
rect 15420 1225 15532 1263
rect 15420 1191 15459 1225
rect 15493 1191 15532 1225
rect 15420 1153 15532 1191
rect 15420 1119 15459 1153
rect 15493 1119 15532 1153
rect 15420 1081 15532 1119
rect 15420 1047 15459 1081
rect 15493 1047 15532 1081
rect 15420 1009 15532 1047
rect 15420 975 15459 1009
rect 15493 975 15532 1009
rect 15420 937 15532 975
rect 15420 903 15459 937
rect 15493 903 15532 937
rect 15420 865 15532 903
rect 15420 831 15459 865
rect 15493 831 15532 865
rect 15420 793 15532 831
rect 15420 759 15459 793
rect 15493 759 15532 793
rect 15420 721 15532 759
rect 15420 687 15459 721
rect 15493 687 15532 721
rect 15420 649 15532 687
rect 15420 615 15459 649
rect 15493 615 15532 649
rect 15420 577 15532 615
rect 15420 543 15459 577
rect 15493 543 15532 577
rect 15420 505 15532 543
rect 15420 471 15459 505
rect 15493 471 15532 505
rect 15420 433 15532 471
rect 15420 399 15459 433
rect 15493 399 15532 433
rect 15420 361 15532 399
rect 15420 327 15459 361
rect 15493 327 15532 361
rect 15420 289 15532 327
rect 15420 255 15459 289
rect 15493 255 15532 289
rect 15420 217 15532 255
rect 15420 183 15459 217
rect 15493 183 15532 217
rect 15420 145 15532 183
rect 15420 111 15459 145
rect 15493 111 15532 145
rect 15420 73 15532 111
rect 15420 39 15459 73
rect 15493 39 15532 73
rect 15420 1 15532 39
rect 15420 -33 15459 1
rect 15493 -33 15532 1
rect 15420 -71 15532 -33
rect 15420 -105 15459 -71
rect 15493 -105 15532 -71
rect 15420 -143 15532 -105
rect 24344 1297 24456 1335
rect 24344 1263 24383 1297
rect 24417 1263 24456 1297
rect 24344 1225 24456 1263
rect 24344 1191 24383 1225
rect 24417 1191 24456 1225
rect 24344 1153 24456 1191
rect 24344 1119 24383 1153
rect 24417 1119 24456 1153
rect 24344 1081 24456 1119
rect 24344 1047 24383 1081
rect 24417 1047 24456 1081
rect 24344 1009 24456 1047
rect 24344 975 24383 1009
rect 24417 975 24456 1009
rect 24344 937 24456 975
rect 24344 903 24383 937
rect 24417 903 24456 937
rect 24344 865 24456 903
rect 24344 831 24383 865
rect 24417 831 24456 865
rect 24344 793 24456 831
rect 24344 759 24383 793
rect 24417 759 24456 793
rect 24344 721 24456 759
rect 24344 687 24383 721
rect 24417 687 24456 721
rect 24344 649 24456 687
rect 24344 615 24383 649
rect 24417 615 24456 649
rect 24344 577 24456 615
rect 24344 543 24383 577
rect 24417 543 24456 577
rect 24344 505 24456 543
rect 24344 471 24383 505
rect 24417 471 24456 505
rect 24344 433 24456 471
rect 24344 399 24383 433
rect 24417 399 24456 433
rect 24344 361 24456 399
rect 24344 327 24383 361
rect 24417 327 24456 361
rect 24344 289 24456 327
rect 24344 255 24383 289
rect 24417 255 24456 289
rect 24344 217 24456 255
rect 24344 183 24383 217
rect 24417 183 24456 217
rect 24344 145 24456 183
rect 24344 111 24383 145
rect 24417 111 24456 145
rect 24344 73 24456 111
rect 24344 39 24383 73
rect 24417 39 24456 73
rect 24344 1 24456 39
rect 24344 -33 24383 1
rect 24417 -33 24456 1
rect 24344 -71 24456 -33
rect 24344 -105 24383 -71
rect 24417 -105 24456 -71
rect 15420 -177 15459 -143
rect 15493 -177 15532 -143
rect 15420 -215 15532 -177
rect 15420 -249 15459 -215
rect 15493 -249 15532 -215
rect 15420 -287 15532 -249
rect 15420 -321 15459 -287
rect 15493 -321 15532 -287
rect 15420 -359 15532 -321
rect 15420 -393 15459 -359
rect 15493 -393 15532 -359
rect 15420 -431 15532 -393
rect 15420 -465 15459 -431
rect 15493 -465 15532 -431
rect 15420 -503 15532 -465
rect 15420 -537 15459 -503
rect 15493 -537 15532 -503
rect 15420 -575 15532 -537
rect 15420 -609 15459 -575
rect 15493 -609 15532 -575
rect 15420 -647 15532 -609
rect 15420 -681 15459 -647
rect 15493 -681 15532 -647
rect 15420 -719 15532 -681
rect 15420 -753 15459 -719
rect 15493 -753 15532 -719
rect 15420 -791 15532 -753
rect 15420 -825 15459 -791
rect 15493 -825 15532 -791
rect 15420 -863 15532 -825
rect 15420 -897 15459 -863
rect 15493 -897 15532 -863
rect 15420 -935 15532 -897
rect 15420 -969 15459 -935
rect 15493 -969 15532 -935
rect 15420 -1007 15532 -969
rect 15788 -982 15848 -162
rect 16020 -982 16080 -254
rect 16246 -982 16306 -130
rect 16478 -360 16538 -252
rect 16934 -360 16994 -254
rect 16472 -364 16544 -360
rect 16472 -416 16482 -364
rect 16534 -416 16544 -364
rect 16472 -420 16544 -416
rect 16928 -364 17000 -360
rect 16928 -416 16938 -364
rect 16990 -416 17000 -364
rect 16928 -420 17000 -416
rect 17162 -728 17222 -136
rect 17394 -360 17454 -248
rect 17850 -360 17910 -254
rect 17388 -364 17460 -360
rect 17388 -416 17398 -364
rect 17450 -416 17460 -364
rect 17388 -420 17460 -416
rect 17844 -364 17916 -360
rect 17844 -416 17854 -364
rect 17906 -416 17916 -364
rect 17844 -420 17916 -416
rect 18078 -594 18138 -134
rect 18308 -360 18368 -254
rect 18772 -360 18832 -250
rect 18302 -364 18374 -360
rect 18302 -416 18312 -364
rect 18364 -416 18374 -364
rect 18302 -420 18374 -416
rect 18766 -364 18838 -360
rect 18766 -416 18776 -364
rect 18828 -416 18838 -364
rect 18766 -420 18838 -416
rect 18994 -470 19054 -116
rect 19222 -360 19282 -256
rect 19678 -360 19738 -256
rect 20146 -360 20206 -256
rect 20604 -360 20664 -260
rect 19216 -364 19288 -360
rect 19216 -416 19226 -364
rect 19278 -416 19288 -364
rect 19216 -420 19288 -416
rect 19672 -364 19744 -360
rect 19672 -416 19682 -364
rect 19734 -416 19744 -364
rect 19672 -420 19744 -416
rect 20140 -364 20212 -360
rect 20140 -416 20150 -364
rect 20202 -416 20212 -364
rect 20140 -420 20212 -416
rect 20598 -364 20670 -360
rect 20598 -416 20608 -364
rect 20660 -416 20670 -364
rect 20598 -420 20670 -416
rect 20824 -470 20884 -150
rect 21060 -360 21120 -254
rect 21516 -360 21576 -254
rect 21054 -364 21126 -360
rect 21054 -416 21064 -364
rect 21116 -416 21126 -364
rect 21054 -420 21126 -416
rect 21510 -364 21582 -360
rect 21510 -416 21520 -364
rect 21572 -416 21582 -364
rect 21510 -420 21582 -416
rect 18994 -530 20884 -470
rect 21740 -594 21800 -136
rect 21972 -360 22032 -254
rect 22428 -360 22488 -258
rect 21966 -364 22038 -360
rect 21966 -416 21976 -364
rect 22028 -416 22038 -364
rect 21966 -420 22038 -416
rect 22422 -364 22494 -360
rect 22422 -416 22432 -364
rect 22484 -416 22494 -364
rect 22422 -420 22494 -416
rect 18078 -654 21800 -594
rect 22660 -728 22720 -138
rect 22886 -360 22946 -254
rect 23346 -360 23406 -250
rect 22880 -364 22952 -360
rect 22880 -416 22890 -364
rect 22942 -416 22952 -364
rect 22880 -420 22952 -416
rect 23340 -364 23412 -360
rect 23340 -416 23350 -364
rect 23402 -416 23412 -364
rect 23340 -420 23412 -416
rect 17162 -788 22720 -728
rect 23576 -982 23636 -118
rect 23806 -982 23866 -252
rect 24034 -982 24094 -124
rect 24344 -143 24456 -105
rect 24344 -177 24383 -143
rect 24417 -177 24456 -143
rect 24344 -215 24456 -177
rect 24344 -249 24383 -215
rect 24417 -249 24456 -215
rect 24344 -287 24456 -249
rect 24344 -321 24383 -287
rect 24417 -321 24456 -287
rect 24344 -359 24456 -321
rect 24344 -393 24383 -359
rect 24417 -393 24456 -359
rect 24344 -431 24456 -393
rect 24344 -465 24383 -431
rect 24417 -465 24456 -431
rect 24344 -503 24456 -465
rect 24344 -537 24383 -503
rect 24417 -537 24456 -503
rect 24344 -575 24456 -537
rect 24344 -609 24383 -575
rect 24417 -609 24456 -575
rect 24344 -647 24456 -609
rect 24344 -681 24383 -647
rect 24417 -681 24456 -647
rect 24344 -719 24456 -681
rect 24344 -753 24383 -719
rect 24417 -753 24456 -719
rect 24344 -791 24456 -753
rect 24344 -825 24383 -791
rect 24417 -825 24456 -791
rect 24344 -863 24456 -825
rect 24344 -897 24383 -863
rect 24417 -897 24456 -863
rect 24344 -935 24456 -897
rect 24344 -969 24383 -935
rect 24417 -969 24456 -935
rect 24344 -982 24456 -969
rect 15420 -1041 15459 -1007
rect 15493 -1041 15532 -1007
rect 15420 -1079 15532 -1041
rect 15420 -1113 15459 -1079
rect 15493 -1113 15532 -1079
rect 15760 -1007 24458 -982
rect 15760 -1009 24383 -1007
rect 15760 -1061 15796 -1009
rect 15848 -1061 16396 -1009
rect 16448 -1061 16996 -1009
rect 17048 -1061 17596 -1009
rect 17648 -1061 18196 -1009
rect 18248 -1061 18796 -1009
rect 18848 -1061 19396 -1009
rect 19448 -1061 19996 -1009
rect 20048 -1061 20596 -1009
rect 20648 -1061 21196 -1009
rect 21248 -1061 21796 -1009
rect 21848 -1061 22396 -1009
rect 22448 -1061 22996 -1009
rect 23048 -1061 23596 -1009
rect 23648 -1061 24016 -1009
rect 24068 -1041 24383 -1009
rect 24417 -1041 24458 -1007
rect 24068 -1061 24458 -1041
rect 15760 -1079 24458 -1061
rect 15760 -1092 24383 -1079
rect 15420 -1151 15532 -1113
rect 15420 -1185 15459 -1151
rect 15493 -1185 15532 -1151
rect 15420 -1223 15532 -1185
rect 15420 -1257 15459 -1223
rect 15493 -1252 15532 -1223
rect 24344 -1113 24383 -1092
rect 24417 -1092 24458 -1079
rect 24417 -1113 24456 -1092
rect 24344 -1151 24456 -1113
rect 24344 -1185 24383 -1151
rect 24417 -1185 24456 -1151
rect 24344 -1223 24456 -1185
rect 24344 -1252 24383 -1223
rect 15493 -1257 15924 -1252
rect 15420 -1280 15924 -1257
rect 15420 -1295 15537 -1280
rect 15420 -1329 15459 -1295
rect 15493 -1329 15537 -1295
rect 15420 -1524 15537 -1329
rect 15909 -1524 15924 -1280
rect 15420 -1552 15924 -1524
rect 23656 -1257 24383 -1252
rect 24417 -1257 24456 -1223
rect 23656 -1280 24456 -1257
rect 23656 -1524 23691 -1280
rect 24319 -1295 24456 -1280
rect 24319 -1329 24383 -1295
rect 24417 -1329 24456 -1295
rect 24319 -1524 24456 -1329
rect 23656 -1552 24456 -1524
rect 15420 -1591 24456 -1552
rect 15420 -1625 15529 -1591
rect 15563 -1625 15601 -1591
rect 15635 -1625 15673 -1591
rect 15707 -1625 15745 -1591
rect 15779 -1625 15817 -1591
rect 15851 -1625 15889 -1591
rect 15923 -1625 15961 -1591
rect 15995 -1625 16033 -1591
rect 16067 -1625 16105 -1591
rect 16139 -1625 16177 -1591
rect 16211 -1625 16249 -1591
rect 16283 -1625 16321 -1591
rect 16355 -1625 16393 -1591
rect 16427 -1625 16465 -1591
rect 16499 -1625 16537 -1591
rect 16571 -1625 16609 -1591
rect 16643 -1625 16681 -1591
rect 16715 -1625 16753 -1591
rect 16787 -1625 16825 -1591
rect 16859 -1625 16897 -1591
rect 16931 -1625 16969 -1591
rect 17003 -1625 17041 -1591
rect 17075 -1625 17113 -1591
rect 17147 -1625 17185 -1591
rect 17219 -1625 17257 -1591
rect 17291 -1625 17329 -1591
rect 17363 -1625 17401 -1591
rect 17435 -1625 17473 -1591
rect 17507 -1625 17545 -1591
rect 17579 -1625 17617 -1591
rect 17651 -1625 17689 -1591
rect 17723 -1625 17761 -1591
rect 17795 -1625 17833 -1591
rect 17867 -1625 17905 -1591
rect 17939 -1625 17977 -1591
rect 18011 -1625 18049 -1591
rect 18083 -1625 18121 -1591
rect 18155 -1625 18193 -1591
rect 18227 -1625 18265 -1591
rect 18299 -1625 18337 -1591
rect 18371 -1625 18409 -1591
rect 18443 -1625 18481 -1591
rect 18515 -1625 18553 -1591
rect 18587 -1625 18625 -1591
rect 18659 -1625 18697 -1591
rect 18731 -1625 18769 -1591
rect 18803 -1625 18841 -1591
rect 18875 -1625 18913 -1591
rect 18947 -1625 18985 -1591
rect 19019 -1625 19057 -1591
rect 19091 -1625 19129 -1591
rect 19163 -1625 19201 -1591
rect 19235 -1625 19273 -1591
rect 19307 -1625 19345 -1591
rect 19379 -1625 19417 -1591
rect 19451 -1625 19489 -1591
rect 19523 -1625 19561 -1591
rect 19595 -1625 19633 -1591
rect 19667 -1625 19705 -1591
rect 19739 -1625 19777 -1591
rect 19811 -1625 19849 -1591
rect 19883 -1625 19921 -1591
rect 19955 -1625 19993 -1591
rect 20027 -1625 20065 -1591
rect 20099 -1625 20137 -1591
rect 20171 -1625 20209 -1591
rect 20243 -1625 20281 -1591
rect 20315 -1625 20353 -1591
rect 20387 -1625 20425 -1591
rect 20459 -1625 20497 -1591
rect 20531 -1625 20569 -1591
rect 20603 -1625 20641 -1591
rect 20675 -1625 20713 -1591
rect 20747 -1625 20785 -1591
rect 20819 -1625 20857 -1591
rect 20891 -1625 20929 -1591
rect 20963 -1625 21001 -1591
rect 21035 -1625 21073 -1591
rect 21107 -1625 21145 -1591
rect 21179 -1625 21217 -1591
rect 21251 -1625 21289 -1591
rect 21323 -1625 21361 -1591
rect 21395 -1625 21433 -1591
rect 21467 -1625 21505 -1591
rect 21539 -1625 21577 -1591
rect 21611 -1625 21649 -1591
rect 21683 -1625 21721 -1591
rect 21755 -1625 21793 -1591
rect 21827 -1625 21865 -1591
rect 21899 -1625 21937 -1591
rect 21971 -1625 22009 -1591
rect 22043 -1625 22081 -1591
rect 22115 -1625 22153 -1591
rect 22187 -1625 22225 -1591
rect 22259 -1625 22297 -1591
rect 22331 -1625 22369 -1591
rect 22403 -1625 22441 -1591
rect 22475 -1625 22513 -1591
rect 22547 -1625 22585 -1591
rect 22619 -1625 22657 -1591
rect 22691 -1625 22729 -1591
rect 22763 -1625 22801 -1591
rect 22835 -1625 22873 -1591
rect 22907 -1625 22945 -1591
rect 22979 -1625 23017 -1591
rect 23051 -1625 23089 -1591
rect 23123 -1625 23161 -1591
rect 23195 -1625 23233 -1591
rect 23267 -1625 23305 -1591
rect 23339 -1625 23377 -1591
rect 23411 -1625 23449 -1591
rect 23483 -1625 23521 -1591
rect 23555 -1625 23593 -1591
rect 23627 -1625 23665 -1591
rect 23699 -1625 23737 -1591
rect 23771 -1625 23809 -1591
rect 23843 -1625 23881 -1591
rect 23915 -1625 23953 -1591
rect 23987 -1625 24025 -1591
rect 24059 -1625 24097 -1591
rect 24131 -1625 24169 -1591
rect 24203 -1625 24241 -1591
rect 24275 -1625 24313 -1591
rect 24347 -1625 24456 -1591
rect 15420 -1664 24456 -1625
rect 25234 -5664 25294 2284
rect 30504 2278 30564 2284
rect 31506 2280 31566 2284
rect 31506 2267 31666 2280
rect 31506 2233 31613 2267
rect 31647 2233 31666 2267
rect 31506 2220 31666 2233
rect 31700 2269 31908 2282
rect 31700 2235 31719 2269
rect 31753 2235 31855 2269
rect 31889 2235 31908 2269
rect 31700 2222 31908 2235
rect 32192 2269 32478 2282
rect 32192 2235 32211 2269
rect 32245 2235 32478 2269
rect 32192 2222 32478 2235
rect 25546 2196 25606 2206
rect 25546 2144 25550 2196
rect 25602 2144 25606 2196
rect 25400 -364 25472 -360
rect 25400 -416 25410 -364
rect 25462 -416 25472 -364
rect 25400 -420 25472 -416
rect 25406 -3260 25466 -420
rect 25406 -3270 25468 -3260
rect 25406 -3322 25412 -3270
rect 25464 -3322 25468 -3270
rect 25406 -3332 25468 -3322
rect 25228 -5668 25300 -5664
rect 25228 -5720 25238 -5668
rect 25290 -5720 25300 -5668
rect 25228 -5724 25300 -5720
rect 15000 -5932 15190 -5928
rect 15000 -5984 15128 -5932
rect 15180 -5984 15190 -5932
rect 15000 -5988 15190 -5984
rect 15010 -9654 15182 -9650
rect 15010 -9706 15120 -9654
rect 15172 -9706 15182 -9654
rect 15010 -9710 15182 -9706
rect 23994 -11898 24128 -11894
rect 23994 -11950 24066 -11898
rect 24118 -11950 24128 -11898
rect 23994 -11954 24128 -11950
rect 25406 -16308 25466 -3332
rect 25546 -9650 25606 2144
rect 26002 2161 31458 2200
rect 26002 2127 26121 2161
rect 26155 2127 26193 2161
rect 26227 2127 26265 2161
rect 26299 2127 26337 2161
rect 26371 2127 26409 2161
rect 26443 2127 26481 2161
rect 26515 2127 26553 2161
rect 26587 2127 26625 2161
rect 26659 2127 26697 2161
rect 26731 2127 26769 2161
rect 26803 2127 26841 2161
rect 26875 2127 26913 2161
rect 26947 2127 26985 2161
rect 27019 2127 27057 2161
rect 27091 2127 27129 2161
rect 27163 2127 27201 2161
rect 27235 2127 27273 2161
rect 27307 2127 27345 2161
rect 27379 2127 27417 2161
rect 27451 2127 27489 2161
rect 27523 2127 27561 2161
rect 27595 2127 27633 2161
rect 27667 2127 27705 2161
rect 27739 2127 27777 2161
rect 27811 2127 27849 2161
rect 27883 2127 27921 2161
rect 27955 2127 27993 2161
rect 28027 2127 28065 2161
rect 28099 2127 28137 2161
rect 28171 2127 28209 2161
rect 28243 2127 28281 2161
rect 28315 2127 28353 2161
rect 28387 2127 28425 2161
rect 28459 2127 28497 2161
rect 28531 2127 28569 2161
rect 28603 2127 28641 2161
rect 28675 2127 28713 2161
rect 28747 2127 28785 2161
rect 28819 2127 28857 2161
rect 28891 2127 28929 2161
rect 28963 2127 29001 2161
rect 29035 2127 29073 2161
rect 29107 2127 29145 2161
rect 29179 2127 29217 2161
rect 29251 2127 29289 2161
rect 29323 2127 29361 2161
rect 29395 2127 29433 2161
rect 29467 2127 29505 2161
rect 29539 2127 29577 2161
rect 29611 2127 29649 2161
rect 29683 2127 29721 2161
rect 29755 2127 29793 2161
rect 29827 2127 29865 2161
rect 29899 2127 29937 2161
rect 29971 2127 30009 2161
rect 30043 2127 30081 2161
rect 30115 2127 30153 2161
rect 30187 2127 30225 2161
rect 30259 2127 30297 2161
rect 30331 2127 30369 2161
rect 30403 2127 30441 2161
rect 30475 2127 30513 2161
rect 30547 2127 30585 2161
rect 30619 2127 30657 2161
rect 30691 2127 30729 2161
rect 30763 2127 30801 2161
rect 30835 2127 30873 2161
rect 30907 2127 30945 2161
rect 30979 2127 31017 2161
rect 31051 2127 31089 2161
rect 31123 2127 31161 2161
rect 31195 2127 31233 2161
rect 31267 2127 31305 2161
rect 31339 2127 31458 2161
rect 26002 2088 31458 2127
rect 26002 1905 26114 2088
rect 26002 1871 26041 1905
rect 26075 1871 26114 1905
rect 26002 1833 26114 1871
rect 26002 1799 26041 1833
rect 26075 1799 26114 1833
rect 26002 1761 26114 1799
rect 26384 1778 26444 2088
rect 26612 1858 26672 2088
rect 26002 1727 26041 1761
rect 26075 1727 26114 1761
rect 26002 1689 26114 1727
rect 26002 1655 26041 1689
rect 26075 1655 26114 1689
rect 26002 1617 26114 1655
rect 26002 1583 26041 1617
rect 26075 1583 26114 1617
rect 26002 1545 26114 1583
rect 26002 1511 26041 1545
rect 26075 1511 26114 1545
rect 26002 1473 26114 1511
rect 26002 1439 26041 1473
rect 26075 1439 26114 1473
rect 26002 1401 26114 1439
rect 26002 1367 26041 1401
rect 26075 1367 26114 1401
rect 26002 1329 26114 1367
rect 26002 1295 26041 1329
rect 26075 1295 26114 1329
rect 26002 1257 26114 1295
rect 26002 1223 26041 1257
rect 26075 1223 26114 1257
rect 26002 1185 26114 1223
rect 26002 1151 26041 1185
rect 26075 1151 26114 1185
rect 26002 1113 26114 1151
rect 26002 1079 26041 1113
rect 26075 1079 26114 1113
rect 26002 1041 26114 1079
rect 26002 1007 26041 1041
rect 26075 1007 26114 1041
rect 26002 969 26114 1007
rect 26002 935 26041 969
rect 26075 935 26114 969
rect 26002 897 26114 935
rect 26002 863 26041 897
rect 26075 863 26114 897
rect 26002 825 26114 863
rect 26002 791 26041 825
rect 26075 791 26114 825
rect 26002 753 26114 791
rect 26002 719 26041 753
rect 26075 719 26114 753
rect 26002 681 26114 719
rect 26002 647 26041 681
rect 26075 647 26114 681
rect 26002 609 26114 647
rect 26002 575 26041 609
rect 26075 575 26114 609
rect 26002 537 26114 575
rect 26002 503 26041 537
rect 26075 503 26114 537
rect 26002 465 26114 503
rect 26002 431 26041 465
rect 26075 431 26114 465
rect 26002 420 26114 431
rect 26384 420 26444 670
rect 26612 420 26672 562
rect 26842 420 26902 2088
rect 27066 2026 27126 2032
rect 27528 2026 27588 2032
rect 27982 2026 28042 2032
rect 28444 2026 28504 2032
rect 28898 2026 28958 2032
rect 29348 2026 29408 2032
rect 29814 2026 29874 2032
rect 30270 2026 30330 2032
rect 30504 2028 30564 2038
rect 27060 2022 30336 2026
rect 27060 1970 27070 2022
rect 27122 1970 27532 2022
rect 27584 1970 27986 2022
rect 28038 1970 28448 2022
rect 28500 1970 28902 2022
rect 28954 1970 29352 2022
rect 29404 1970 29818 2022
rect 29870 1970 30274 2022
rect 30326 1970 30336 2022
rect 27060 1966 30336 1970
rect 30504 1976 30508 2028
rect 30560 1976 30564 2028
rect 27066 1854 27126 1966
rect 27528 1870 27588 1966
rect 27982 1864 28042 1966
rect 28444 1864 28504 1966
rect 28898 1864 28958 1966
rect 29348 1870 29408 1966
rect 29814 1876 29874 1966
rect 30270 1870 30330 1966
rect 30504 1732 30564 1976
rect 30734 1856 30794 2088
rect 30962 1764 31022 2088
rect 31346 1994 31458 2088
rect 31346 1905 31542 1994
rect 31346 1871 31385 1905
rect 31419 1898 31542 1905
rect 31419 1871 31458 1898
rect 31346 1833 31458 1871
rect 31346 1799 31385 1833
rect 31419 1799 31458 1833
rect 31346 1761 31458 1799
rect 31346 1727 31385 1761
rect 31419 1727 31458 1761
rect 31346 1689 31458 1727
rect 31346 1655 31385 1689
rect 31419 1655 31458 1689
rect 31346 1617 31458 1655
rect 31346 1583 31385 1617
rect 31419 1583 31458 1617
rect 31346 1545 31458 1583
rect 31346 1511 31385 1545
rect 31419 1511 31458 1545
rect 31346 1473 31458 1511
rect 31346 1439 31385 1473
rect 31419 1439 31458 1473
rect 31346 1401 31458 1439
rect 31346 1367 31385 1401
rect 31419 1367 31458 1401
rect 31346 1329 31458 1367
rect 31346 1295 31385 1329
rect 31419 1295 31458 1329
rect 31346 1257 31458 1295
rect 31346 1223 31385 1257
rect 31419 1223 31458 1257
rect 31346 1185 31458 1223
rect 31346 1151 31385 1185
rect 31419 1151 31458 1185
rect 31346 1113 31458 1151
rect 31346 1079 31385 1113
rect 31419 1079 31458 1113
rect 31346 1041 31458 1079
rect 31346 1007 31385 1041
rect 31419 1007 31458 1041
rect 31346 969 31458 1007
rect 31346 935 31385 969
rect 31419 935 31458 969
rect 31346 897 31458 935
rect 31346 863 31385 897
rect 31419 863 31458 897
rect 31346 825 31458 863
rect 31346 791 31385 825
rect 31419 791 31458 825
rect 31346 753 31458 791
rect 31346 719 31385 753
rect 31419 719 31458 753
rect 31346 681 31458 719
rect 31346 647 31385 681
rect 31419 647 31458 681
rect 26002 393 26902 420
rect 27074 454 27134 566
rect 27536 454 27596 550
rect 27990 454 28050 556
rect 28452 454 28512 556
rect 28906 454 28966 556
rect 29356 454 29416 550
rect 29822 454 29882 544
rect 30278 454 30338 550
rect 30734 472 30794 562
rect 30964 472 31024 638
rect 31346 609 31458 647
rect 31346 575 31385 609
rect 31419 575 31458 609
rect 31346 537 31458 575
rect 31346 503 31385 537
rect 31419 503 31458 537
rect 31346 472 31458 503
rect 30734 465 31458 472
rect 27074 450 30344 454
rect 27074 398 30282 450
rect 30334 398 30344 450
rect 27074 394 30344 398
rect 30734 431 31385 465
rect 31419 431 31458 465
rect 30734 412 31458 431
rect 26002 359 26041 393
rect 26075 360 26902 393
rect 26075 359 26114 360
rect 26002 321 26114 359
rect 26002 287 26041 321
rect 26075 287 26114 321
rect 26002 249 26114 287
rect 26002 215 26041 249
rect 26075 215 26114 249
rect 26002 177 26114 215
rect 26002 143 26041 177
rect 26075 143 26114 177
rect 26002 105 26114 143
rect 26002 71 26041 105
rect 26075 71 26114 105
rect 26002 33 26114 71
rect 26002 -1 26041 33
rect 26075 -1 26114 33
rect 26002 -39 26114 -1
rect 26002 -73 26041 -39
rect 26075 -73 26114 -39
rect 26002 -111 26114 -73
rect 26002 -145 26041 -111
rect 26075 -145 26114 -111
rect 26002 -183 26114 -145
rect 26002 -217 26041 -183
rect 26075 -217 26114 -183
rect 26002 -255 26114 -217
rect 26002 -289 26041 -255
rect 26075 -289 26114 -255
rect 26002 -327 26114 -289
rect 26002 -361 26041 -327
rect 26075 -361 26114 -327
rect 26002 -399 26114 -361
rect 26002 -433 26041 -399
rect 26075 -433 26114 -399
rect 26002 -471 26114 -433
rect 26002 -505 26041 -471
rect 26075 -505 26114 -471
rect 26002 -543 26114 -505
rect 26002 -577 26041 -543
rect 26075 -577 26114 -543
rect 26002 -615 26114 -577
rect 26002 -649 26041 -615
rect 26075 -649 26114 -615
rect 26002 -687 26114 -649
rect 26002 -721 26041 -687
rect 26075 -721 26114 -687
rect 26002 -759 26114 -721
rect 26002 -793 26041 -759
rect 26075 -793 26114 -759
rect 26002 -831 26114 -793
rect 26002 -865 26041 -831
rect 26075 -865 26114 -831
rect 26002 -903 26114 -865
rect 26002 -937 26041 -903
rect 26075 -937 26114 -903
rect 26002 -975 26114 -937
rect 26002 -982 26041 -975
rect 26000 -1009 26041 -982
rect 26075 -982 26114 -975
rect 26384 -982 26444 360
rect 26612 -982 26672 360
rect 26842 -982 26902 360
rect 30734 -982 30794 412
rect 30964 -982 31024 412
rect 31346 393 31458 412
rect 31346 359 31385 393
rect 31419 359 31458 393
rect 31346 321 31458 359
rect 31346 287 31385 321
rect 31419 287 31458 321
rect 31346 249 31458 287
rect 31346 215 31385 249
rect 31419 215 31458 249
rect 31346 177 31458 215
rect 31346 143 31385 177
rect 31419 143 31458 177
rect 31346 105 31458 143
rect 31346 71 31385 105
rect 31419 71 31458 105
rect 31346 33 31458 71
rect 31346 -1 31385 33
rect 31419 -1 31458 33
rect 31346 -39 31458 -1
rect 31346 -73 31385 -39
rect 31419 -73 31458 -39
rect 31346 -111 31458 -73
rect 31346 -145 31385 -111
rect 31419 -145 31458 -111
rect 31346 -183 31458 -145
rect 31346 -217 31385 -183
rect 31419 -217 31458 -183
rect 31346 -255 31458 -217
rect 31346 -289 31385 -255
rect 31419 -289 31458 -255
rect 31346 -327 31458 -289
rect 31346 -361 31385 -327
rect 31419 -361 31458 -327
rect 31346 -399 31458 -361
rect 31346 -433 31385 -399
rect 31419 -433 31458 -399
rect 31346 -471 31458 -433
rect 31346 -505 31385 -471
rect 31419 -505 31458 -471
rect 31346 -543 31458 -505
rect 31346 -577 31385 -543
rect 31419 -577 31458 -543
rect 31346 -615 31458 -577
rect 31346 -649 31385 -615
rect 31419 -649 31458 -615
rect 31346 -687 31458 -649
rect 31346 -721 31385 -687
rect 31419 -721 31458 -687
rect 31346 -759 31458 -721
rect 31346 -793 31385 -759
rect 31419 -793 31458 -759
rect 31346 -831 31458 -793
rect 31346 -865 31385 -831
rect 31419 -865 31458 -831
rect 31346 -903 31458 -865
rect 31346 -937 31385 -903
rect 31419 -937 31458 -903
rect 31346 -975 31458 -937
rect 26075 -1009 31274 -982
rect 26000 -1047 26312 -1009
rect 26000 -1081 26041 -1047
rect 26075 -1061 26312 -1047
rect 26364 -1061 26912 -1009
rect 26964 -1061 27512 -1009
rect 27564 -1061 28112 -1009
rect 28164 -1061 28712 -1009
rect 28764 -1061 29312 -1009
rect 29364 -1061 29912 -1009
rect 29964 -1061 30512 -1009
rect 30564 -1061 31112 -1009
rect 31164 -1061 31274 -1009
rect 26075 -1081 31274 -1061
rect 26000 -1092 31274 -1081
rect 31346 -1009 31385 -975
rect 31419 -1009 31458 -975
rect 31346 -1047 31458 -1009
rect 31346 -1081 31385 -1047
rect 31419 -1081 31458 -1047
rect 26002 -1119 26114 -1092
rect 26002 -1153 26041 -1119
rect 26075 -1153 26114 -1119
rect 26002 -1191 26114 -1153
rect 26002 -1225 26041 -1191
rect 26075 -1225 26114 -1191
rect 26002 -1252 26114 -1225
rect 31346 -1119 31458 -1081
rect 31346 -1153 31385 -1119
rect 31419 -1153 31458 -1119
rect 31346 -1191 31458 -1153
rect 31346 -1225 31385 -1191
rect 31419 -1225 31458 -1191
rect 31346 -1252 31458 -1225
rect 26002 -1263 26724 -1252
rect 26002 -1297 26041 -1263
rect 26075 -1280 26724 -1263
rect 26075 -1297 26132 -1280
rect 26002 -1335 26132 -1297
rect 26002 -1369 26041 -1335
rect 26075 -1369 26132 -1335
rect 26002 -1524 26132 -1369
rect 26696 -1524 26724 -1280
rect 26002 -1552 26724 -1524
rect 30736 -1263 31458 -1252
rect 30736 -1280 31385 -1263
rect 30736 -1524 30764 -1280
rect 31328 -1297 31385 -1280
rect 31419 -1297 31458 -1263
rect 31328 -1335 31458 -1297
rect 31328 -1369 31385 -1335
rect 31419 -1369 31458 -1335
rect 31328 -1524 31458 -1369
rect 30736 -1552 31458 -1524
rect 26002 -1591 31458 -1552
rect 26002 -1625 26121 -1591
rect 26155 -1625 26193 -1591
rect 26227 -1625 26265 -1591
rect 26299 -1625 26337 -1591
rect 26371 -1625 26409 -1591
rect 26443 -1625 26481 -1591
rect 26515 -1625 26553 -1591
rect 26587 -1625 26625 -1591
rect 26659 -1625 26697 -1591
rect 26731 -1625 26769 -1591
rect 26803 -1625 26841 -1591
rect 26875 -1625 26913 -1591
rect 26947 -1625 26985 -1591
rect 27019 -1625 27057 -1591
rect 27091 -1625 27129 -1591
rect 27163 -1625 27201 -1591
rect 27235 -1625 27273 -1591
rect 27307 -1625 27345 -1591
rect 27379 -1625 27417 -1591
rect 27451 -1625 27489 -1591
rect 27523 -1625 27561 -1591
rect 27595 -1625 27633 -1591
rect 27667 -1625 27705 -1591
rect 27739 -1625 27777 -1591
rect 27811 -1625 27849 -1591
rect 27883 -1625 27921 -1591
rect 27955 -1625 27993 -1591
rect 28027 -1625 28065 -1591
rect 28099 -1625 28137 -1591
rect 28171 -1625 28209 -1591
rect 28243 -1625 28281 -1591
rect 28315 -1625 28353 -1591
rect 28387 -1625 28425 -1591
rect 28459 -1625 28497 -1591
rect 28531 -1625 28569 -1591
rect 28603 -1625 28641 -1591
rect 28675 -1625 28713 -1591
rect 28747 -1625 28785 -1591
rect 28819 -1625 28857 -1591
rect 28891 -1625 28929 -1591
rect 28963 -1625 29001 -1591
rect 29035 -1625 29073 -1591
rect 29107 -1625 29145 -1591
rect 29179 -1625 29217 -1591
rect 29251 -1625 29289 -1591
rect 29323 -1625 29361 -1591
rect 29395 -1625 29433 -1591
rect 29467 -1625 29505 -1591
rect 29539 -1625 29577 -1591
rect 29611 -1625 29649 -1591
rect 29683 -1625 29721 -1591
rect 29755 -1625 29793 -1591
rect 29827 -1625 29865 -1591
rect 29899 -1625 29937 -1591
rect 29971 -1625 30009 -1591
rect 30043 -1625 30081 -1591
rect 30115 -1625 30153 -1591
rect 30187 -1625 30225 -1591
rect 30259 -1625 30297 -1591
rect 30331 -1625 30369 -1591
rect 30403 -1625 30441 -1591
rect 30475 -1625 30513 -1591
rect 30547 -1625 30585 -1591
rect 30619 -1625 30657 -1591
rect 30691 -1625 30729 -1591
rect 30763 -1625 30801 -1591
rect 30835 -1625 30873 -1591
rect 30907 -1625 30945 -1591
rect 30979 -1625 31017 -1591
rect 31051 -1625 31089 -1591
rect 31123 -1625 31161 -1591
rect 31195 -1625 31233 -1591
rect 31267 -1625 31305 -1591
rect 31339 -1625 31458 -1591
rect 26002 -1664 31458 -1625
rect 25540 -9654 25612 -9650
rect 25540 -9706 25550 -9654
rect 25602 -9706 25612 -9654
rect 25540 -9710 25612 -9706
rect 26914 -9654 26974 -9644
rect 26914 -9706 26918 -9654
rect 26970 -9706 26974 -9654
rect 25406 -16360 25410 -16308
rect 25462 -16360 25466 -16308
rect 25406 -23240 25466 -16360
rect 25546 -11898 25606 -9710
rect 26914 -9716 26974 -9706
rect 25546 -11950 25550 -11898
rect 25602 -11950 25606 -11898
rect 25400 -23244 25472 -23240
rect 25400 -23296 25410 -23244
rect 25462 -23296 25472 -23244
rect 25400 -23300 25472 -23296
rect 15118 -27654 15178 -27644
rect 25546 -27650 25606 -11950
rect 35856 -11894 35916 -11888
rect 35856 -11898 36076 -11894
rect 35856 -11950 35860 -11898
rect 35912 -11950 36076 -11898
rect 35856 -11954 36076 -11950
rect 35856 -11960 35916 -11954
rect 15118 -27706 15122 -27654
rect 15174 -27706 15178 -27654
rect 15118 -27716 15178 -27706
rect 25540 -27654 25612 -27650
rect 25540 -27706 25550 -27654
rect 25602 -27706 25612 -27654
rect 25540 -27710 25612 -27706
rect 26908 -27654 27050 -27650
rect 26908 -27706 26918 -27654
rect 26970 -27706 27050 -27654
rect 26908 -27710 27050 -27706
<< via1 >>
rect 15537 3932 15909 4176
rect 23691 3932 24319 4176
rect 17622 3657 17674 3709
rect 18202 3657 18254 3709
rect 18802 3657 18854 3709
rect 19402 3657 19454 3709
rect 20002 3657 20054 3709
rect 20602 3657 20654 3709
rect 21202 3657 21254 3709
rect 21802 3657 21854 3709
rect 22402 3657 22454 3709
rect 21518 3392 21570 3444
rect 18082 2712 18134 2764
rect 26132 3932 26696 4176
rect 30764 3932 31328 4176
rect 26384 3657 26436 3709
rect 26964 3657 27016 3709
rect 27564 3657 27616 3709
rect 28164 3657 28216 3709
rect 28764 3657 28816 3709
rect 29364 3657 29416 3709
rect 29964 3657 30016 3709
rect 30564 3657 30616 3709
rect 31164 3657 31216 3709
rect 27070 2838 27122 2890
rect 27532 2838 27584 2890
rect 27986 2840 28038 2892
rect 28448 2838 28500 2890
rect 28902 2838 28954 2890
rect 29352 2838 29404 2890
rect 29818 2838 29870 2890
rect 30274 2838 30326 2890
rect 30508 2630 30560 2682
rect 30508 2288 30560 2340
rect 16478 1558 16530 1610
rect 16934 1558 16986 1610
rect 17394 1558 17446 1610
rect 17850 1558 17902 1610
rect 18308 1558 18360 1610
rect 18772 1558 18824 1610
rect 19226 1558 19278 1610
rect 19686 1558 19738 1610
rect 19916 1558 19968 1610
rect 20144 1558 20196 1610
rect 20600 1558 20652 1610
rect 21060 1558 21112 1610
rect 21516 1558 21568 1610
rect 21972 1558 22024 1610
rect 22428 1558 22480 1610
rect 22886 1558 22938 1610
rect 23346 1558 23398 1610
rect 16482 -416 16534 -364
rect 16938 -416 16990 -364
rect 17398 -416 17450 -364
rect 17854 -416 17906 -364
rect 18312 -416 18364 -364
rect 18776 -416 18828 -364
rect 19226 -416 19278 -364
rect 19682 -416 19734 -364
rect 20150 -416 20202 -364
rect 20608 -416 20660 -364
rect 21064 -416 21116 -364
rect 21520 -416 21572 -364
rect 21976 -416 22028 -364
rect 22432 -416 22484 -364
rect 22890 -416 22942 -364
rect 23350 -416 23402 -364
rect 15796 -1061 15848 -1009
rect 16396 -1061 16448 -1009
rect 16996 -1061 17048 -1009
rect 17596 -1061 17648 -1009
rect 18196 -1061 18248 -1009
rect 18796 -1061 18848 -1009
rect 19396 -1061 19448 -1009
rect 19996 -1061 20048 -1009
rect 20596 -1061 20648 -1009
rect 21196 -1061 21248 -1009
rect 21796 -1061 21848 -1009
rect 22396 -1061 22448 -1009
rect 22996 -1061 23048 -1009
rect 23596 -1061 23648 -1009
rect 24016 -1061 24068 -1009
rect 15537 -1524 15909 -1280
rect 23691 -1524 24319 -1280
rect 25550 2144 25602 2196
rect 25410 -416 25462 -364
rect 25412 -3322 25464 -3270
rect 25238 -5720 25290 -5668
rect 15128 -5984 15180 -5932
rect 15120 -9706 15172 -9654
rect 24066 -11950 24118 -11898
rect 27070 1970 27122 2022
rect 27532 1970 27584 2022
rect 27986 1970 28038 2022
rect 28448 1970 28500 2022
rect 28902 1970 28954 2022
rect 29352 1970 29404 2022
rect 29818 1970 29870 2022
rect 30274 1970 30326 2022
rect 30508 1976 30560 2028
rect 30282 398 30334 450
rect 26312 -1061 26364 -1009
rect 26912 -1061 26964 -1009
rect 27512 -1061 27564 -1009
rect 28112 -1061 28164 -1009
rect 28712 -1061 28764 -1009
rect 29312 -1061 29364 -1009
rect 29912 -1061 29964 -1009
rect 30512 -1061 30564 -1009
rect 31112 -1061 31164 -1009
rect 26132 -1524 26696 -1280
rect 30764 -1524 31328 -1280
rect 25550 -9706 25602 -9654
rect 26918 -9706 26970 -9654
rect 25410 -16360 25462 -16308
rect 25550 -11950 25602 -11898
rect 25410 -23296 25462 -23244
rect 35860 -11950 35912 -11898
rect 15122 -27706 15174 -27654
rect 25550 -27706 25602 -27654
rect 26918 -27706 26970 -27654
<< metal2 >>
rect 15532 4202 15914 4214
rect 15532 3906 15535 4202
rect 15911 3906 15914 4202
rect 15532 3894 15914 3906
rect 23666 4202 24344 4214
rect 23666 4176 23697 4202
rect 24313 4176 24344 4202
rect 23666 3932 23691 4176
rect 24319 3932 24344 4176
rect 23666 3906 23697 3932
rect 24313 3906 24344 3932
rect 23666 3894 24344 3906
rect 26114 4202 26714 4214
rect 26114 4176 26146 4202
rect 26682 4176 26714 4202
rect 26114 3932 26132 4176
rect 26696 3932 26714 4176
rect 26114 3906 26146 3932
rect 26682 3906 26714 3932
rect 26114 3894 26714 3906
rect 30746 4202 31346 4214
rect 30746 4176 30778 4202
rect 31314 4176 31346 4202
rect 30746 3932 30764 4176
rect 31328 3932 31346 4176
rect 30746 3906 30778 3932
rect 31314 3906 31346 3932
rect 30746 3894 31346 3906
rect 17550 3711 22522 3756
rect 17550 3655 17620 3711
rect 17676 3655 18200 3711
rect 18256 3655 18800 3711
rect 18856 3655 19400 3711
rect 19456 3655 20000 3711
rect 20056 3655 20600 3711
rect 20656 3655 21200 3711
rect 21256 3655 21800 3711
rect 21856 3655 22400 3711
rect 22456 3655 22522 3711
rect 17550 3612 22522 3655
rect 26312 3711 31284 3756
rect 26312 3655 26382 3711
rect 26438 3655 26962 3711
rect 27018 3655 27562 3711
rect 27618 3655 28162 3711
rect 28218 3655 28762 3711
rect 28818 3655 29362 3711
rect 29418 3655 29962 3711
rect 30018 3655 30562 3711
rect 30618 3655 31162 3711
rect 31218 3655 31284 3711
rect 26312 3612 31284 3655
rect 21514 3448 21574 3454
rect 21514 3444 25606 3448
rect 21514 3392 21518 3444
rect 21570 3392 25606 3444
rect 21514 3388 25606 3392
rect 21514 3382 21574 3388
rect 18072 2764 18144 2768
rect 18072 2712 18082 2764
rect 18134 2712 18144 2764
rect 18072 2708 18144 2712
rect 16474 1614 16534 1620
rect 16930 1614 16990 1620
rect 17390 1614 17450 1620
rect 17846 1614 17906 1620
rect 18078 1614 18138 2708
rect 25546 2200 25606 3388
rect 27066 2890 27126 2900
rect 27066 2838 27070 2890
rect 27122 2838 27126 2890
rect 25540 2196 25612 2200
rect 25540 2144 25550 2196
rect 25602 2144 25612 2196
rect 25540 2140 25612 2144
rect 27066 2022 27126 2838
rect 27066 1970 27070 2022
rect 27122 1970 27126 2022
rect 27066 1960 27126 1970
rect 27528 2890 27588 2900
rect 27528 2838 27532 2890
rect 27584 2838 27588 2890
rect 27528 2022 27588 2838
rect 27982 2892 28042 2902
rect 27982 2840 27986 2892
rect 28038 2840 28042 2892
rect 27982 2026 28042 2840
rect 28444 2890 28504 2900
rect 28444 2838 28448 2890
rect 28500 2838 28504 2890
rect 28444 2026 28504 2838
rect 28898 2890 28958 2900
rect 28898 2838 28902 2890
rect 28954 2838 28958 2890
rect 27528 1970 27532 2022
rect 27584 1970 27588 2022
rect 27528 1960 27588 1970
rect 27976 2022 28048 2026
rect 27976 1970 27986 2022
rect 28038 1970 28048 2022
rect 27976 1966 28048 1970
rect 28438 2022 28510 2026
rect 28438 1970 28448 2022
rect 28500 1970 28510 2022
rect 28438 1966 28510 1970
rect 28898 2022 28958 2838
rect 29348 2890 29408 2900
rect 29348 2838 29352 2890
rect 29404 2838 29408 2890
rect 29348 2026 29408 2838
rect 29814 2890 29874 2900
rect 29814 2838 29818 2890
rect 29870 2838 29874 2890
rect 29814 2026 29874 2838
rect 30270 2890 30330 2900
rect 30270 2838 30274 2890
rect 30326 2838 30330 2890
rect 28898 1970 28902 2022
rect 28954 1970 28958 2022
rect 28898 1960 28958 1970
rect 29342 2022 29414 2026
rect 29342 1970 29352 2022
rect 29404 1970 29414 2022
rect 29342 1966 29414 1970
rect 29808 2022 29880 2026
rect 29808 1970 29818 2022
rect 29870 1970 29880 2022
rect 29808 1966 29880 1970
rect 30270 2022 30330 2838
rect 30504 2682 30564 2692
rect 30504 2630 30508 2682
rect 30560 2630 30564 2682
rect 30504 2344 30564 2630
rect 30498 2340 30570 2344
rect 30498 2288 30508 2340
rect 30560 2288 30570 2340
rect 30498 2284 30570 2288
rect 30504 2032 30564 2284
rect 30270 1970 30274 2022
rect 30326 1970 30330 2022
rect 30498 2028 30570 2032
rect 30498 1976 30508 2028
rect 30560 1976 30570 2028
rect 30498 1972 30570 1976
rect 30270 1960 30330 1970
rect 18304 1614 18364 1620
rect 18768 1614 18828 1620
rect 19222 1614 19282 1620
rect 19682 1614 19742 1620
rect 19912 1614 19972 1620
rect 20140 1614 20200 1620
rect 20596 1614 20656 1620
rect 21056 1614 21116 1620
rect 21512 1614 21572 1620
rect 21968 1614 22028 1620
rect 22424 1614 22484 1620
rect 22882 1614 22942 1620
rect 23342 1614 23402 1620
rect 16474 1610 23402 1614
rect 16474 1558 16478 1610
rect 16530 1558 16934 1610
rect 16986 1558 17394 1610
rect 17446 1558 17850 1610
rect 17902 1558 18308 1610
rect 18360 1558 18772 1610
rect 18824 1558 19226 1610
rect 19278 1558 19686 1610
rect 19738 1558 19916 1610
rect 19968 1558 20144 1610
rect 20196 1558 20600 1610
rect 20652 1558 21060 1610
rect 21112 1558 21516 1610
rect 21568 1558 21972 1610
rect 22024 1558 22428 1610
rect 22480 1558 22886 1610
rect 22938 1558 23346 1610
rect 23398 1558 23402 1610
rect 16474 1554 23402 1558
rect 16474 1548 16534 1554
rect 16930 1548 16990 1554
rect 17390 1548 17450 1554
rect 17846 1548 17906 1554
rect 18304 1548 18364 1554
rect 18768 1548 18828 1554
rect 19222 1548 19282 1554
rect 19682 1548 19742 1554
rect 19912 1548 19972 1554
rect 20140 1548 20200 1554
rect 20596 1548 20656 1554
rect 21056 1548 21116 1554
rect 21512 1548 21572 1554
rect 21968 1548 22028 1554
rect 22424 1548 22484 1554
rect 22882 1548 22942 1554
rect 23342 1548 23402 1554
rect 30278 454 30338 460
rect 30278 450 31902 454
rect 30278 398 30282 450
rect 30334 398 31902 450
rect 30278 394 31902 398
rect 30278 388 30338 394
rect 16478 -360 16538 -354
rect 16934 -360 16994 -354
rect 17394 -360 17454 -354
rect 17850 -360 17910 -354
rect 18308 -360 18368 -354
rect 18772 -360 18832 -354
rect 19222 -360 19282 -354
rect 19678 -360 19738 -354
rect 20146 -360 20206 -354
rect 20604 -360 20664 -354
rect 21060 -360 21120 -354
rect 21516 -360 21576 -354
rect 21972 -360 22032 -354
rect 22428 -360 22488 -354
rect 22886 -360 22946 -354
rect 23346 -360 23406 -354
rect 25406 -360 25466 -354
rect 16478 -364 25466 -360
rect 16478 -416 16482 -364
rect 16534 -416 16938 -364
rect 16990 -416 17398 -364
rect 17450 -416 17854 -364
rect 17906 -416 18312 -364
rect 18364 -416 18776 -364
rect 18828 -416 19226 -364
rect 19278 -416 19682 -364
rect 19734 -416 20150 -364
rect 20202 -416 20608 -364
rect 20660 -416 21064 -364
rect 21116 -416 21520 -364
rect 21572 -416 21976 -364
rect 22028 -416 22432 -364
rect 22484 -416 22890 -364
rect 22942 -416 23350 -364
rect 23402 -416 25410 -364
rect 25462 -416 25466 -364
rect 16478 -420 25466 -416
rect 16478 -426 16538 -420
rect 16934 -426 16994 -420
rect 17394 -426 17454 -420
rect 17850 -426 17910 -420
rect 18308 -426 18368 -420
rect 18772 -426 18832 -420
rect 19222 -426 19282 -420
rect 19678 -426 19738 -420
rect 20146 -426 20206 -420
rect 20604 -426 20664 -420
rect 21060 -426 21120 -420
rect 21516 -426 21576 -420
rect 21972 -426 22032 -420
rect 22428 -426 22488 -420
rect 22886 -426 22946 -420
rect 23346 -426 23406 -420
rect 25406 -426 25466 -420
rect 31802 -948 31902 394
rect 15760 -1007 24116 -982
rect 15760 -1063 15794 -1007
rect 15850 -1063 16394 -1007
rect 16450 -1063 16994 -1007
rect 17050 -1063 17594 -1007
rect 17650 -1063 18194 -1007
rect 18250 -1063 18794 -1007
rect 18850 -1063 19394 -1007
rect 19450 -1063 19994 -1007
rect 20050 -1063 20594 -1007
rect 20650 -1063 21194 -1007
rect 21250 -1063 21794 -1007
rect 21850 -1063 22394 -1007
rect 22450 -1063 22994 -1007
rect 23050 -1063 23594 -1007
rect 23650 -1063 24014 -1007
rect 24070 -1063 24116 -1007
rect 15760 -1092 24116 -1063
rect 26276 -1007 31274 -982
rect 26276 -1063 26310 -1007
rect 26366 -1063 26910 -1007
rect 26966 -1063 27510 -1007
rect 27566 -1063 28110 -1007
rect 28166 -1063 28710 -1007
rect 28766 -1063 29310 -1007
rect 29366 -1063 29910 -1007
rect 29966 -1063 30510 -1007
rect 30566 -1063 31110 -1007
rect 31166 -1063 31274 -1007
rect 31802 -1048 36438 -948
rect 26276 -1092 31274 -1063
rect 15532 -1254 15914 -1242
rect 15532 -1550 15535 -1254
rect 15911 -1550 15914 -1254
rect 15532 -1562 15914 -1550
rect 23666 -1254 24344 -1242
rect 23666 -1280 23697 -1254
rect 24313 -1280 24344 -1254
rect 23666 -1524 23691 -1280
rect 24319 -1524 24344 -1280
rect 23666 -1550 23697 -1524
rect 24313 -1550 24344 -1524
rect 23666 -1562 24344 -1550
rect 26114 -1254 26714 -1242
rect 26114 -1280 26146 -1254
rect 26682 -1280 26714 -1254
rect 26114 -1524 26132 -1280
rect 26696 -1524 26714 -1280
rect 26114 -1550 26146 -1524
rect 26682 -1550 26714 -1524
rect 26114 -1562 26714 -1550
rect 30746 -1254 31346 -1242
rect 30746 -1280 30778 -1254
rect 31314 -1280 31346 -1254
rect 30746 -1524 30764 -1280
rect 31328 -1524 31346 -1280
rect 30746 -1550 30778 -1524
rect 31314 -1550 31346 -1524
rect 30746 -1562 31346 -1550
rect 19242 -3270 27720 -3266
rect 19242 -3322 25412 -3270
rect 25464 -3322 27720 -3270
rect 19242 -3326 27720 -3322
rect 25234 -5664 25294 -5658
rect 16180 -5668 25294 -5664
rect 16180 -5720 25238 -5668
rect 25290 -5720 25294 -5668
rect 16180 -5724 25294 -5720
rect 15124 -5928 15184 -5922
rect 16180 -5928 16240 -5724
rect 25234 -5730 25294 -5724
rect 15124 -5932 16240 -5928
rect 15124 -5984 15128 -5932
rect 15180 -5984 16240 -5932
rect 15124 -5988 16240 -5984
rect 15124 -5994 15184 -5988
rect 25616 -7958 25676 -7949
rect 25616 -7960 27308 -7958
rect 25616 -8016 25618 -7960
rect 25674 -8016 27308 -7960
rect 25616 -8018 27308 -8016
rect 25616 -8027 25676 -8018
rect 36338 -8128 36438 -1048
rect 15116 -9650 15176 -9644
rect 25546 -9650 25606 -9644
rect 15116 -9654 26980 -9650
rect 15116 -9706 15120 -9654
rect 15172 -9706 25550 -9654
rect 25602 -9706 26918 -9654
rect 26970 -9706 26980 -9654
rect 15116 -9710 26980 -9706
rect 15116 -9716 15176 -9710
rect 25546 -9716 25606 -9710
rect 24062 -11894 24122 -11888
rect 24062 -11898 35922 -11894
rect 24062 -11950 24066 -11898
rect 24118 -11950 25550 -11898
rect 25602 -11950 35860 -11898
rect 35912 -11950 35922 -11898
rect 24062 -11954 35922 -11950
rect 24062 -11960 24122 -11954
rect 10630 -13357 10690 -13352
rect 10600 -13374 10708 -13357
rect 10600 -13430 10626 -13374
rect 10682 -13430 10708 -13374
rect 10600 -13447 10708 -13430
rect 10630 -25958 10690 -13447
rect 25300 -13586 25360 -13577
rect 23754 -13588 25360 -13586
rect 23754 -13644 25302 -13588
rect 25358 -13644 25360 -13588
rect 23754 -13646 25360 -13644
rect 38988 -13646 40380 -13586
rect 25300 -13655 25360 -13646
rect 23180 -16308 32052 -16304
rect 23180 -16360 25410 -16308
rect 25462 -16360 32052 -16308
rect 23180 -16364 32052 -16360
rect 25406 -23240 25466 -23234
rect 19246 -23244 27852 -23240
rect 19246 -23296 25410 -23244
rect 25462 -23296 27852 -23244
rect 19246 -23300 27852 -23296
rect 25406 -23306 25466 -23300
rect 10630 -26018 12078 -25958
rect 25420 -26018 27060 -25958
rect 25420 -26157 25480 -26018
rect 40320 -26157 40380 -13646
rect 25398 -26174 25506 -26157
rect 25398 -26230 25424 -26174
rect 25480 -26230 25506 -26174
rect 25398 -26247 25506 -26230
rect 40296 -26174 40404 -26157
rect 40296 -26230 40322 -26174
rect 40378 -26230 40404 -26174
rect 40296 -26247 40404 -26230
rect 25420 -26252 25480 -26247
rect 40320 -26252 40380 -26247
rect 25546 -27650 25606 -27644
rect 26914 -27650 26974 -27644
rect 15112 -27654 26974 -27650
rect 15112 -27706 15122 -27654
rect 15174 -27706 25550 -27654
rect 25602 -27706 26918 -27654
rect 26970 -27706 26974 -27654
rect 15112 -27710 26974 -27706
rect 25546 -27716 25606 -27710
rect 26914 -27716 26974 -27710
<< via2 >>
rect 15535 4176 15911 4202
rect 15535 3932 15537 4176
rect 15537 3932 15909 4176
rect 15909 3932 15911 4176
rect 15535 3906 15911 3932
rect 23697 4176 24313 4202
rect 23697 3932 24313 4176
rect 23697 3906 24313 3932
rect 26146 4176 26682 4202
rect 26146 3932 26682 4176
rect 26146 3906 26682 3932
rect 30778 4176 31314 4202
rect 30778 3932 31314 4176
rect 30778 3906 31314 3932
rect 17620 3709 17676 3711
rect 17620 3657 17622 3709
rect 17622 3657 17674 3709
rect 17674 3657 17676 3709
rect 17620 3655 17676 3657
rect 18200 3709 18256 3711
rect 18200 3657 18202 3709
rect 18202 3657 18254 3709
rect 18254 3657 18256 3709
rect 18200 3655 18256 3657
rect 18800 3709 18856 3711
rect 18800 3657 18802 3709
rect 18802 3657 18854 3709
rect 18854 3657 18856 3709
rect 18800 3655 18856 3657
rect 19400 3709 19456 3711
rect 19400 3657 19402 3709
rect 19402 3657 19454 3709
rect 19454 3657 19456 3709
rect 19400 3655 19456 3657
rect 20000 3709 20056 3711
rect 20000 3657 20002 3709
rect 20002 3657 20054 3709
rect 20054 3657 20056 3709
rect 20000 3655 20056 3657
rect 20600 3709 20656 3711
rect 20600 3657 20602 3709
rect 20602 3657 20654 3709
rect 20654 3657 20656 3709
rect 20600 3655 20656 3657
rect 21200 3709 21256 3711
rect 21200 3657 21202 3709
rect 21202 3657 21254 3709
rect 21254 3657 21256 3709
rect 21200 3655 21256 3657
rect 21800 3709 21856 3711
rect 21800 3657 21802 3709
rect 21802 3657 21854 3709
rect 21854 3657 21856 3709
rect 21800 3655 21856 3657
rect 22400 3709 22456 3711
rect 22400 3657 22402 3709
rect 22402 3657 22454 3709
rect 22454 3657 22456 3709
rect 22400 3655 22456 3657
rect 26382 3709 26438 3711
rect 26382 3657 26384 3709
rect 26384 3657 26436 3709
rect 26436 3657 26438 3709
rect 26382 3655 26438 3657
rect 26962 3709 27018 3711
rect 26962 3657 26964 3709
rect 26964 3657 27016 3709
rect 27016 3657 27018 3709
rect 26962 3655 27018 3657
rect 27562 3709 27618 3711
rect 27562 3657 27564 3709
rect 27564 3657 27616 3709
rect 27616 3657 27618 3709
rect 27562 3655 27618 3657
rect 28162 3709 28218 3711
rect 28162 3657 28164 3709
rect 28164 3657 28216 3709
rect 28216 3657 28218 3709
rect 28162 3655 28218 3657
rect 28762 3709 28818 3711
rect 28762 3657 28764 3709
rect 28764 3657 28816 3709
rect 28816 3657 28818 3709
rect 28762 3655 28818 3657
rect 29362 3709 29418 3711
rect 29362 3657 29364 3709
rect 29364 3657 29416 3709
rect 29416 3657 29418 3709
rect 29362 3655 29418 3657
rect 29962 3709 30018 3711
rect 29962 3657 29964 3709
rect 29964 3657 30016 3709
rect 30016 3657 30018 3709
rect 29962 3655 30018 3657
rect 30562 3709 30618 3711
rect 30562 3657 30564 3709
rect 30564 3657 30616 3709
rect 30616 3657 30618 3709
rect 30562 3655 30618 3657
rect 31162 3709 31218 3711
rect 31162 3657 31164 3709
rect 31164 3657 31216 3709
rect 31216 3657 31218 3709
rect 31162 3655 31218 3657
rect 15794 -1009 15850 -1007
rect 15794 -1061 15796 -1009
rect 15796 -1061 15848 -1009
rect 15848 -1061 15850 -1009
rect 15794 -1063 15850 -1061
rect 16394 -1009 16450 -1007
rect 16394 -1061 16396 -1009
rect 16396 -1061 16448 -1009
rect 16448 -1061 16450 -1009
rect 16394 -1063 16450 -1061
rect 16994 -1009 17050 -1007
rect 16994 -1061 16996 -1009
rect 16996 -1061 17048 -1009
rect 17048 -1061 17050 -1009
rect 16994 -1063 17050 -1061
rect 17594 -1009 17650 -1007
rect 17594 -1061 17596 -1009
rect 17596 -1061 17648 -1009
rect 17648 -1061 17650 -1009
rect 17594 -1063 17650 -1061
rect 18194 -1009 18250 -1007
rect 18194 -1061 18196 -1009
rect 18196 -1061 18248 -1009
rect 18248 -1061 18250 -1009
rect 18194 -1063 18250 -1061
rect 18794 -1009 18850 -1007
rect 18794 -1061 18796 -1009
rect 18796 -1061 18848 -1009
rect 18848 -1061 18850 -1009
rect 18794 -1063 18850 -1061
rect 19394 -1009 19450 -1007
rect 19394 -1061 19396 -1009
rect 19396 -1061 19448 -1009
rect 19448 -1061 19450 -1009
rect 19394 -1063 19450 -1061
rect 19994 -1009 20050 -1007
rect 19994 -1061 19996 -1009
rect 19996 -1061 20048 -1009
rect 20048 -1061 20050 -1009
rect 19994 -1063 20050 -1061
rect 20594 -1009 20650 -1007
rect 20594 -1061 20596 -1009
rect 20596 -1061 20648 -1009
rect 20648 -1061 20650 -1009
rect 20594 -1063 20650 -1061
rect 21194 -1009 21250 -1007
rect 21194 -1061 21196 -1009
rect 21196 -1061 21248 -1009
rect 21248 -1061 21250 -1009
rect 21194 -1063 21250 -1061
rect 21794 -1009 21850 -1007
rect 21794 -1061 21796 -1009
rect 21796 -1061 21848 -1009
rect 21848 -1061 21850 -1009
rect 21794 -1063 21850 -1061
rect 22394 -1009 22450 -1007
rect 22394 -1061 22396 -1009
rect 22396 -1061 22448 -1009
rect 22448 -1061 22450 -1009
rect 22394 -1063 22450 -1061
rect 22994 -1009 23050 -1007
rect 22994 -1061 22996 -1009
rect 22996 -1061 23048 -1009
rect 23048 -1061 23050 -1009
rect 22994 -1063 23050 -1061
rect 23594 -1009 23650 -1007
rect 23594 -1061 23596 -1009
rect 23596 -1061 23648 -1009
rect 23648 -1061 23650 -1009
rect 23594 -1063 23650 -1061
rect 24014 -1009 24070 -1007
rect 24014 -1061 24016 -1009
rect 24016 -1061 24068 -1009
rect 24068 -1061 24070 -1009
rect 24014 -1063 24070 -1061
rect 26310 -1009 26366 -1007
rect 26310 -1061 26312 -1009
rect 26312 -1061 26364 -1009
rect 26364 -1061 26366 -1009
rect 26310 -1063 26366 -1061
rect 26910 -1009 26966 -1007
rect 26910 -1061 26912 -1009
rect 26912 -1061 26964 -1009
rect 26964 -1061 26966 -1009
rect 26910 -1063 26966 -1061
rect 27510 -1009 27566 -1007
rect 27510 -1061 27512 -1009
rect 27512 -1061 27564 -1009
rect 27564 -1061 27566 -1009
rect 27510 -1063 27566 -1061
rect 28110 -1009 28166 -1007
rect 28110 -1061 28112 -1009
rect 28112 -1061 28164 -1009
rect 28164 -1061 28166 -1009
rect 28110 -1063 28166 -1061
rect 28710 -1009 28766 -1007
rect 28710 -1061 28712 -1009
rect 28712 -1061 28764 -1009
rect 28764 -1061 28766 -1009
rect 28710 -1063 28766 -1061
rect 29310 -1009 29366 -1007
rect 29310 -1061 29312 -1009
rect 29312 -1061 29364 -1009
rect 29364 -1061 29366 -1009
rect 29310 -1063 29366 -1061
rect 29910 -1009 29966 -1007
rect 29910 -1061 29912 -1009
rect 29912 -1061 29964 -1009
rect 29964 -1061 29966 -1009
rect 29910 -1063 29966 -1061
rect 30510 -1009 30566 -1007
rect 30510 -1061 30512 -1009
rect 30512 -1061 30564 -1009
rect 30564 -1061 30566 -1009
rect 30510 -1063 30566 -1061
rect 31110 -1009 31166 -1007
rect 31110 -1061 31112 -1009
rect 31112 -1061 31164 -1009
rect 31164 -1061 31166 -1009
rect 31110 -1063 31166 -1061
rect 15535 -1280 15911 -1254
rect 15535 -1524 15537 -1280
rect 15537 -1524 15909 -1280
rect 15909 -1524 15911 -1280
rect 15535 -1550 15911 -1524
rect 23697 -1280 24313 -1254
rect 23697 -1524 24313 -1280
rect 23697 -1550 24313 -1524
rect 26146 -1280 26682 -1254
rect 26146 -1524 26682 -1280
rect 26146 -1550 26682 -1524
rect 30778 -1280 31314 -1254
rect 30778 -1524 31314 -1280
rect 30778 -1550 31314 -1524
rect 25618 -8016 25674 -7960
rect 10626 -13430 10682 -13374
rect 25302 -13644 25358 -13588
rect 25424 -26230 25480 -26174
rect 40322 -26230 40378 -26174
<< metal3 >>
rect 15522 4202 15924 4209
rect 15522 3906 15535 4202
rect 15911 3906 15924 4202
rect 15522 3899 15924 3906
rect 23656 4202 24354 4209
rect 23656 4166 23697 4202
rect 24313 4166 24354 4202
rect 23656 3942 23693 4166
rect 24317 3942 24354 4166
rect 23656 3906 23697 3942
rect 24313 3906 24354 3942
rect 23656 3899 24354 3906
rect 26104 4202 26724 4209
rect 26104 4166 26146 4202
rect 26682 4166 26724 4202
rect 26104 3942 26142 4166
rect 26686 3942 26724 4166
rect 26104 3906 26146 3942
rect 26682 3906 26724 3942
rect 26104 3899 26724 3906
rect 30736 4202 31356 4209
rect 30736 4166 30778 4202
rect 31314 4166 31356 4202
rect 30736 3942 30774 4166
rect 31318 3942 31356 4166
rect 30736 3906 30778 3942
rect 31314 3906 31356 3942
rect 30736 3899 31356 3906
rect 17550 3715 22522 3756
rect 17550 3651 17616 3715
rect 17680 3651 18196 3715
rect 18260 3651 18796 3715
rect 18860 3651 19396 3715
rect 19460 3651 19996 3715
rect 20060 3651 20596 3715
rect 20660 3651 21196 3715
rect 21260 3651 21796 3715
rect 21860 3651 22396 3715
rect 22460 3651 22522 3715
rect 17550 3612 22522 3651
rect 26312 3715 31284 3756
rect 26312 3651 26378 3715
rect 26442 3651 26958 3715
rect 27022 3651 27558 3715
rect 27622 3651 28158 3715
rect 28222 3651 28758 3715
rect 28822 3651 29358 3715
rect 29422 3651 29958 3715
rect 30022 3651 30558 3715
rect 30622 3651 31158 3715
rect 31222 3651 31284 3715
rect 26312 3612 31284 3651
rect 15760 -1007 24116 -982
rect 15760 -1063 15794 -1007
rect 15850 -1063 16394 -1007
rect 16450 -1063 16994 -1007
rect 17050 -1063 17594 -1007
rect 17650 -1063 18194 -1007
rect 18250 -1063 18794 -1007
rect 18850 -1063 19394 -1007
rect 19450 -1063 19994 -1007
rect 20050 -1063 20594 -1007
rect 20650 -1063 21194 -1007
rect 21250 -1063 21794 -1007
rect 21850 -1063 22394 -1007
rect 22450 -1063 22994 -1007
rect 23050 -1063 23594 -1007
rect 23650 -1063 24014 -1007
rect 24070 -1063 24116 -1007
rect 15760 -1092 24116 -1063
rect 26276 -1007 31274 -982
rect 26276 -1063 26310 -1007
rect 26366 -1063 26910 -1007
rect 26966 -1063 27510 -1007
rect 27566 -1063 28110 -1007
rect 28166 -1063 28710 -1007
rect 28766 -1063 29310 -1007
rect 29366 -1063 29910 -1007
rect 29966 -1063 30510 -1007
rect 30566 -1063 31110 -1007
rect 31166 -1063 31274 -1007
rect 26276 -1092 31274 -1063
rect 15522 -1254 15924 -1247
rect 15522 -1550 15535 -1254
rect 15911 -1550 15924 -1254
rect 15522 -1557 15924 -1550
rect 23656 -1254 24354 -1247
rect 23656 -1290 23697 -1254
rect 24313 -1290 24354 -1254
rect 23656 -1514 23693 -1290
rect 24317 -1514 24354 -1290
rect 23656 -1550 23697 -1514
rect 24313 -1550 24354 -1514
rect 23656 -1557 24354 -1550
rect 26104 -1254 26724 -1247
rect 26104 -1290 26146 -1254
rect 26682 -1290 26724 -1254
rect 26104 -1514 26142 -1290
rect 26686 -1514 26724 -1290
rect 26104 -1550 26146 -1514
rect 26682 -1550 26724 -1514
rect 26104 -1557 26724 -1550
rect 30736 -1254 31356 -1247
rect 30736 -1290 30778 -1254
rect 31314 -1290 31356 -1254
rect 30736 -1514 30774 -1290
rect 31318 -1514 31356 -1290
rect 30736 -1550 30778 -1514
rect 31314 -1550 31356 -1514
rect 30736 -1557 31356 -1550
rect 25611 -7958 25681 -7953
rect 25596 -7960 25696 -7958
rect 25596 -8016 25618 -7960
rect 25674 -8016 25696 -7960
rect 25272 -8153 25372 -8152
rect 25267 -8170 25377 -8153
rect 25267 -8234 25290 -8170
rect 25354 -8234 25377 -8170
rect 25267 -8251 25377 -8234
rect 10604 -13353 10704 -13352
rect 10599 -13370 10709 -13353
rect 10599 -13434 10622 -13370
rect 10686 -13434 10709 -13370
rect 10599 -13451 10709 -13434
rect 10604 -13452 10704 -13451
rect 25272 -13588 25372 -8251
rect 25596 -13353 25696 -8016
rect 25591 -13370 25701 -13353
rect 25591 -13434 25614 -13370
rect 25678 -13434 25701 -13370
rect 25591 -13451 25701 -13434
rect 25596 -13452 25696 -13451
rect 25272 -13644 25302 -13588
rect 25358 -13644 25372 -13588
rect 25272 -13662 25372 -13644
rect 25402 -26153 25502 -26152
rect 40300 -26153 40400 -26152
rect 25397 -26170 25507 -26153
rect 25397 -26234 25420 -26170
rect 25484 -26234 25507 -26170
rect 25397 -26251 25507 -26234
rect 40295 -26170 40405 -26153
rect 40295 -26234 40318 -26170
rect 40382 -26234 40405 -26170
rect 40295 -26251 40405 -26234
rect 25402 -26252 25502 -26251
rect 40300 -26252 40400 -26251
<< via3 >>
rect 15571 3942 15875 4166
rect 23693 3942 23697 4166
rect 23697 3942 24313 4166
rect 24313 3942 24317 4166
rect 26142 3942 26146 4166
rect 26146 3942 26682 4166
rect 26682 3942 26686 4166
rect 30774 3942 30778 4166
rect 30778 3942 31314 4166
rect 31314 3942 31318 4166
rect 17616 3711 17680 3715
rect 17616 3655 17620 3711
rect 17620 3655 17676 3711
rect 17676 3655 17680 3711
rect 17616 3651 17680 3655
rect 18196 3711 18260 3715
rect 18196 3655 18200 3711
rect 18200 3655 18256 3711
rect 18256 3655 18260 3711
rect 18196 3651 18260 3655
rect 18796 3711 18860 3715
rect 18796 3655 18800 3711
rect 18800 3655 18856 3711
rect 18856 3655 18860 3711
rect 18796 3651 18860 3655
rect 19396 3711 19460 3715
rect 19396 3655 19400 3711
rect 19400 3655 19456 3711
rect 19456 3655 19460 3711
rect 19396 3651 19460 3655
rect 19996 3711 20060 3715
rect 19996 3655 20000 3711
rect 20000 3655 20056 3711
rect 20056 3655 20060 3711
rect 19996 3651 20060 3655
rect 20596 3711 20660 3715
rect 20596 3655 20600 3711
rect 20600 3655 20656 3711
rect 20656 3655 20660 3711
rect 20596 3651 20660 3655
rect 21196 3711 21260 3715
rect 21196 3655 21200 3711
rect 21200 3655 21256 3711
rect 21256 3655 21260 3711
rect 21196 3651 21260 3655
rect 21796 3711 21860 3715
rect 21796 3655 21800 3711
rect 21800 3655 21856 3711
rect 21856 3655 21860 3711
rect 21796 3651 21860 3655
rect 22396 3711 22460 3715
rect 22396 3655 22400 3711
rect 22400 3655 22456 3711
rect 22456 3655 22460 3711
rect 22396 3651 22460 3655
rect 26378 3711 26442 3715
rect 26378 3655 26382 3711
rect 26382 3655 26438 3711
rect 26438 3655 26442 3711
rect 26378 3651 26442 3655
rect 26958 3711 27022 3715
rect 26958 3655 26962 3711
rect 26962 3655 27018 3711
rect 27018 3655 27022 3711
rect 26958 3651 27022 3655
rect 27558 3711 27622 3715
rect 27558 3655 27562 3711
rect 27562 3655 27618 3711
rect 27618 3655 27622 3711
rect 27558 3651 27622 3655
rect 28158 3711 28222 3715
rect 28158 3655 28162 3711
rect 28162 3655 28218 3711
rect 28218 3655 28222 3711
rect 28158 3651 28222 3655
rect 28758 3711 28822 3715
rect 28758 3655 28762 3711
rect 28762 3655 28818 3711
rect 28818 3655 28822 3711
rect 28758 3651 28822 3655
rect 29358 3711 29422 3715
rect 29358 3655 29362 3711
rect 29362 3655 29418 3711
rect 29418 3655 29422 3711
rect 29358 3651 29422 3655
rect 29958 3711 30022 3715
rect 29958 3655 29962 3711
rect 29962 3655 30018 3711
rect 30018 3655 30022 3711
rect 29958 3651 30022 3655
rect 30558 3711 30622 3715
rect 30558 3655 30562 3711
rect 30562 3655 30618 3711
rect 30618 3655 30622 3711
rect 30558 3651 30622 3655
rect 31158 3711 31222 3715
rect 31158 3655 31162 3711
rect 31162 3655 31218 3711
rect 31218 3655 31222 3711
rect 31158 3651 31222 3655
rect 15571 -1514 15875 -1290
rect 23693 -1514 23697 -1290
rect 23697 -1514 24313 -1290
rect 24313 -1514 24317 -1290
rect 26142 -1514 26146 -1290
rect 26146 -1514 26682 -1290
rect 26682 -1514 26686 -1290
rect 30774 -1514 30778 -1290
rect 30778 -1514 31314 -1290
rect 31314 -1514 31318 -1290
rect 25290 -8234 25354 -8170
rect 10622 -13374 10686 -13370
rect 10622 -13430 10626 -13374
rect 10626 -13430 10682 -13374
rect 10682 -13430 10686 -13374
rect 10622 -13434 10686 -13430
rect 25614 -13434 25678 -13370
rect 25420 -26174 25484 -26170
rect 25420 -26230 25424 -26174
rect 25424 -26230 25480 -26174
rect 25480 -26230 25484 -26174
rect 25420 -26234 25484 -26230
rect 40318 -26174 40382 -26170
rect 40318 -26230 40322 -26174
rect 40322 -26230 40378 -26174
rect 40378 -26230 40382 -26174
rect 40318 -26234 40382 -26230
<< metal4 >>
rect 9784 4266 40288 4388
rect 9784 3710 9906 4266
rect 10462 4166 40288 4266
rect 10462 3942 15571 4166
rect 15875 3942 23693 4166
rect 24317 3942 26142 4166
rect 26686 3942 30774 4166
rect 31318 3942 40288 4166
rect 10462 3715 40288 3942
rect 10462 3710 17616 3715
rect 9784 3651 17616 3710
rect 17680 3651 18196 3715
rect 18260 3651 18796 3715
rect 18860 3651 19396 3715
rect 19460 3651 19996 3715
rect 20060 3651 20596 3715
rect 20660 3651 21196 3715
rect 21260 3651 21796 3715
rect 21860 3651 22396 3715
rect 22460 3651 26378 3715
rect 26442 3651 26958 3715
rect 27022 3651 27558 3715
rect 27622 3651 28158 3715
rect 28222 3651 28758 3715
rect 28822 3651 29358 3715
rect 29422 3651 29958 3715
rect 30022 3651 30558 3715
rect 30622 3651 31158 3715
rect 31222 3651 40288 3715
rect 9784 3588 40288 3651
rect 15348 -940 31530 -936
rect 10744 -1090 41209 -940
rect 10744 -1290 40527 -1090
rect 10744 -1514 15571 -1290
rect 15875 -1514 23693 -1290
rect 24317 -1514 26142 -1290
rect 26686 -1514 30774 -1290
rect 31318 -1514 40527 -1290
rect 10744 -2606 40527 -1514
rect 41083 -2606 41209 -1090
rect 10744 -2750 41209 -2606
rect 25158 -8170 25372 -8152
rect 25158 -8234 25290 -8170
rect 25354 -8234 25372 -8170
rect 25158 -8252 25372 -8234
rect 9780 -9856 12644 -9850
rect 24250 -9856 26734 -9850
rect 9780 -9882 40292 -9856
rect 9780 -11718 9903 -9882
rect 10459 -11718 40292 -9882
rect 9780 -11754 40292 -11718
rect 10604 -13370 10844 -13352
rect 10604 -13434 10622 -13370
rect 10686 -13434 10844 -13370
rect 10604 -13452 10844 -13434
rect 25596 -13370 25860 -13352
rect 25596 -13434 25614 -13370
rect 25678 -13434 25860 -13370
rect 25596 -13452 25860 -13434
rect 10740 -18885 41204 -18850
rect 10740 -20721 40521 -18885
rect 41077 -20721 41204 -18885
rect 10740 -20752 41204 -20721
rect 25190 -26170 25502 -26152
rect 25190 -26234 25420 -26170
rect 25484 -26234 25502 -26170
rect 25190 -26252 25502 -26234
rect 40190 -26170 40400 -26152
rect 40190 -26234 40318 -26170
rect 40382 -26234 40400 -26170
rect 40190 -26252 40400 -26234
rect 9786 -27972 11168 -27850
rect 9786 -28528 9908 -27972
rect 10464 -28528 11168 -27972
rect 9786 -28650 11168 -28528
rect 24488 -28650 26804 -27850
<< via4 >>
rect 9906 3710 10462 4266
rect 40527 -2606 41083 -1090
rect 9903 -11718 10459 -9882
rect 40521 -20721 41077 -18885
rect 9908 -28528 10464 -27972
<< metal5 >>
rect 9786 4412 10586 4472
rect 9760 4266 10608 4412
rect 9760 3710 9906 4266
rect 10462 3710 10608 4266
rect 9760 3564 10608 3710
rect 9786 -9882 10586 3564
rect 9786 -11718 9903 -9882
rect 10459 -11718 10586 -9882
rect 9786 -27826 10586 -11718
rect 40402 -1090 41202 4472
rect 40402 -2606 40527 -1090
rect 41083 -2606 41202 -1090
rect 40402 -18885 41202 -2606
rect 40402 -20721 40521 -18885
rect 41077 -20721 41202 -18885
rect 9762 -27972 10610 -27826
rect 9762 -28528 9908 -27972
rect 10464 -28528 10610 -27972
rect 9762 -28674 10610 -28528
rect 9786 -28686 10586 -28674
rect 40402 -28686 41202 -20721
use cs_ring_osc_stage  cs_ring_osc_stage_5
timestamp 1626065694
transform 1 0 30840 0 1 -12350
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_4
timestamp 1626065694
transform 1 0 15840 0 1 -12350
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_3
timestamp 1626065694
transform -1 0 35194 0 -1 -9254
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_2
timestamp 1626065694
transform -1 0 20194 0 -1 -9254
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_1
timestamp 1626065694
transform 1 0 30840 0 1 -30350
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_0
timestamp 1626065694
transform 1 0 15840 0 1 -30350
box -5100 1696 9450 10400
use sky130_fd_pr__pfet_01v8_hvt_GK2P2M  sky130_fd_pr__pfet_01v8_hvt_GK2P2M_0
timestamp 1626065694
transform 1 0 19941 0 -1 593
box -4187 -900 4187 900
use sky130_fd_pr__pfet_01v8_hvt_8Q5PU3  sky130_fd_pr__pfet_01v8_hvt_8Q5PU3_0
timestamp 1626065694
transform 1 0 28704 0 -1 1213
box -2355 -700 2355 700
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_1
timestamp 1626065694
transform 1 0 28703 0 -1 3144
box -2345 -188 2345 188
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_0
timestamp 1626065694
transform 1 0 19941 0 -1 3144
box -2345 -188 2345 188
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626065694
transform 1 0 31542 0 -1 2490
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1626065694
transform 1 0 31818 0 -1 2490
box -38 -48 498 592
<< labels >>
flabel metal2 s 16596 1582 16604 1588 5 FreeSans 600 0 0 0 vpbias
flabel metal1 s 18498 3414 18504 3422 5 FreeSans 600 0 0 0 vctrl
flabel metal1 s 32398 2246 32414 2260 1 FreeSans 600 0 0 0 voscbuf
flabel metal1 s 31098 2304 31114 2316 1 FreeSans 600 0 0 0 vosc
flabel metal1 s 31796 2256 31804 2260 1 FreeSans 600 0 0 0 vosc2
flabel metal4 s 13612 3930 13632 3948 1 FreeSans 600 0 0 0 VSS
flabel metal4 s 13272 -1542 13284 -1524 1 FreeSans 600 0 0 0 VDD
<< properties >>
string FIXED_BBOX 20128 1902 25472 3682
<< end >>
