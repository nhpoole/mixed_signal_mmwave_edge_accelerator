magic
tech sky130A
magscale 1 2
timestamp 1623983327
use sky130_fd_pr__res_generic_m1_6PYWN2  sky130_fd_pr__res_generic_m1_6PYWN2_0
timestamp 1623983327
transform 1 0 78 0 1 87
box -100 -87 100 87
<< labels >>
flabel space 74 148 76 154 1 FreeSans 480 0 0 0 term1
flabel space 72 16 76 20 1 FreeSans 480 0 0 0 term2
<< end >>
