magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal1 >>
rect 102319 120005 104783 120033
rect 102195 119903 103615 119931
<< metal2 >>
rect 102181 117628 102209 119917
rect 102305 119118 102333 120019
rect 103601 119917 103629 121292
rect 104769 120019 104797 121292
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 104751 0 1 119987
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 102287 0 1 119086
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 102287 0 1 119987
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 103583 0 1 119885
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 102163 0 1 117596
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 102163 0 1 119885
box 0 0 64 64
<< properties >>
string FIXED_BBOX 102163 117596 104815 121292
<< end >>
