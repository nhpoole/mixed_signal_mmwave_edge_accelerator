magic
tech sky130A
magscale 1 2
timestamp 1621999597
<< nwell >>
rect 15390 -1694 24486 2310
rect 25972 2229 31856 2230
rect 25972 1908 32316 2229
rect 25972 -1694 31488 1908
rect 10782 -8068 21298 -1992
rect 25782 -8068 36298 -1992
rect 14736 -19612 25252 -13536
rect 29736 -19612 40252 -13536
rect 10782 -26068 21298 -19992
rect 25782 -26068 36298 -19992
<< pwell >>
rect 15390 2474 24486 4420
rect 25972 2394 31488 4346
rect 31571 2473 31605 2507
rect 31584 2469 31605 2473
rect 31847 2469 31881 2507
rect 31584 2287 31770 2469
rect 31829 2287 32267 2469
rect 10782 -10598 21298 -8232
rect 25782 -10598 36298 -8232
rect 14736 -13372 25252 -11006
rect 29736 -13372 40252 -11006
rect 10782 -28598 21298 -26232
rect 25782 -28598 36298 -26232
<< nmos >>
rect 17680 3044 18080 3244
rect 18138 3044 18538 3244
rect 18596 3044 18996 3244
rect 19054 3044 19454 3244
rect 19512 3044 19912 3244
rect 19970 3044 20370 3244
rect 20428 3044 20828 3244
rect 20886 3044 21286 3244
rect 21344 3044 21744 3244
rect 21802 3044 22202 3244
rect 26442 3044 26842 3244
rect 26900 3044 27300 3244
rect 27358 3044 27758 3244
rect 27816 3044 28216 3244
rect 28274 3044 28674 3244
rect 28732 3044 29132 3244
rect 29190 3044 29590 3244
rect 29648 3044 30048 3244
rect 30106 3044 30506 3244
rect 30564 3044 30964 3244
rect 11290 -8838 11690 -8638
rect 11748 -8838 12148 -8638
rect 12206 -8838 12606 -8638
rect 12664 -8838 13064 -8638
rect 13122 -8838 13522 -8638
rect 13580 -8838 13980 -8638
rect 14038 -8838 14438 -8638
rect 14496 -8838 14896 -8638
rect 14954 -8838 15354 -8638
rect 15412 -8838 15812 -8638
rect 16290 -8838 16690 -8638
rect 16748 -8838 17148 -8638
rect 17206 -8838 17606 -8638
rect 17664 -8838 18064 -8638
rect 18122 -8838 18522 -8638
rect 18580 -8838 18980 -8638
rect 19038 -8838 19438 -8638
rect 19496 -8838 19896 -8638
rect 19954 -8838 20354 -8638
rect 20412 -8838 20812 -8638
rect 11290 -9506 11690 -9306
rect 11748 -9506 12148 -9306
rect 12206 -9506 12606 -9306
rect 12664 -9506 13064 -9306
rect 13122 -9506 13522 -9306
rect 13580 -9506 13980 -9306
rect 14038 -9506 14438 -9306
rect 14496 -9506 14896 -9306
rect 14954 -9506 15354 -9306
rect 15412 -9506 15812 -9306
rect 26290 -8838 26690 -8638
rect 26748 -8838 27148 -8638
rect 27206 -8838 27606 -8638
rect 27664 -8838 28064 -8638
rect 28122 -8838 28522 -8638
rect 28580 -8838 28980 -8638
rect 29038 -8838 29438 -8638
rect 29496 -8838 29896 -8638
rect 29954 -8838 30354 -8638
rect 30412 -8838 30812 -8638
rect 31290 -8838 31690 -8638
rect 31748 -8838 32148 -8638
rect 32206 -8838 32606 -8638
rect 32664 -8838 33064 -8638
rect 33122 -8838 33522 -8638
rect 33580 -8838 33980 -8638
rect 34038 -8838 34438 -8638
rect 34496 -8838 34896 -8638
rect 34954 -8838 35354 -8638
rect 35412 -8838 35812 -8638
rect 26290 -9506 26690 -9306
rect 26748 -9506 27148 -9306
rect 27206 -9506 27606 -9306
rect 27664 -9506 28064 -9306
rect 28122 -9506 28522 -9306
rect 28580 -9506 28980 -9306
rect 29038 -9506 29438 -9306
rect 29496 -9506 29896 -9306
rect 29954 -9506 30354 -9306
rect 30412 -9506 30812 -9306
rect 20222 -12298 20622 -12098
rect 20680 -12298 21080 -12098
rect 21138 -12298 21538 -12098
rect 21596 -12298 21996 -12098
rect 22054 -12298 22454 -12098
rect 22512 -12298 22912 -12098
rect 22970 -12298 23370 -12098
rect 23428 -12298 23828 -12098
rect 23886 -12298 24286 -12098
rect 24344 -12298 24744 -12098
rect 15222 -12966 15622 -12766
rect 15680 -12966 16080 -12766
rect 16138 -12966 16538 -12766
rect 16596 -12966 16996 -12766
rect 17054 -12966 17454 -12766
rect 17512 -12966 17912 -12766
rect 17970 -12966 18370 -12766
rect 18428 -12966 18828 -12766
rect 18886 -12966 19286 -12766
rect 19344 -12966 19744 -12766
rect 20222 -12966 20622 -12766
rect 20680 -12966 21080 -12766
rect 21138 -12966 21538 -12766
rect 21596 -12966 21996 -12766
rect 22054 -12966 22454 -12766
rect 22512 -12966 22912 -12766
rect 22970 -12966 23370 -12766
rect 23428 -12966 23828 -12766
rect 23886 -12966 24286 -12766
rect 24344 -12966 24744 -12766
rect 35222 -12298 35622 -12098
rect 35680 -12298 36080 -12098
rect 36138 -12298 36538 -12098
rect 36596 -12298 36996 -12098
rect 37054 -12298 37454 -12098
rect 37512 -12298 37912 -12098
rect 37970 -12298 38370 -12098
rect 38428 -12298 38828 -12098
rect 38886 -12298 39286 -12098
rect 39344 -12298 39744 -12098
rect 30222 -12966 30622 -12766
rect 30680 -12966 31080 -12766
rect 31138 -12966 31538 -12766
rect 31596 -12966 31996 -12766
rect 32054 -12966 32454 -12766
rect 32512 -12966 32912 -12766
rect 32970 -12966 33370 -12766
rect 33428 -12966 33828 -12766
rect 33886 -12966 34286 -12766
rect 34344 -12966 34744 -12766
rect 35222 -12966 35622 -12766
rect 35680 -12966 36080 -12766
rect 36138 -12966 36538 -12766
rect 36596 -12966 36996 -12766
rect 37054 -12966 37454 -12766
rect 37512 -12966 37912 -12766
rect 37970 -12966 38370 -12766
rect 38428 -12966 38828 -12766
rect 38886 -12966 39286 -12766
rect 39344 -12966 39744 -12766
rect 11290 -26838 11690 -26638
rect 11748 -26838 12148 -26638
rect 12206 -26838 12606 -26638
rect 12664 -26838 13064 -26638
rect 13122 -26838 13522 -26638
rect 13580 -26838 13980 -26638
rect 14038 -26838 14438 -26638
rect 14496 -26838 14896 -26638
rect 14954 -26838 15354 -26638
rect 15412 -26838 15812 -26638
rect 16290 -26838 16690 -26638
rect 16748 -26838 17148 -26638
rect 17206 -26838 17606 -26638
rect 17664 -26838 18064 -26638
rect 18122 -26838 18522 -26638
rect 18580 -26838 18980 -26638
rect 19038 -26838 19438 -26638
rect 19496 -26838 19896 -26638
rect 19954 -26838 20354 -26638
rect 20412 -26838 20812 -26638
rect 11290 -27506 11690 -27306
rect 11748 -27506 12148 -27306
rect 12206 -27506 12606 -27306
rect 12664 -27506 13064 -27306
rect 13122 -27506 13522 -27306
rect 13580 -27506 13980 -27306
rect 14038 -27506 14438 -27306
rect 14496 -27506 14896 -27306
rect 14954 -27506 15354 -27306
rect 15412 -27506 15812 -27306
rect 26290 -26838 26690 -26638
rect 26748 -26838 27148 -26638
rect 27206 -26838 27606 -26638
rect 27664 -26838 28064 -26638
rect 28122 -26838 28522 -26638
rect 28580 -26838 28980 -26638
rect 29038 -26838 29438 -26638
rect 29496 -26838 29896 -26638
rect 29954 -26838 30354 -26638
rect 30412 -26838 30812 -26638
rect 31290 -26838 31690 -26638
rect 31748 -26838 32148 -26638
rect 32206 -26838 32606 -26638
rect 32664 -26838 33064 -26638
rect 33122 -26838 33522 -26638
rect 33580 -26838 33980 -26638
rect 34038 -26838 34438 -26638
rect 34496 -26838 34896 -26638
rect 34954 -26838 35354 -26638
rect 35412 -26838 35812 -26638
rect 26290 -27506 26690 -27306
rect 26748 -27506 27148 -27306
rect 27206 -27506 27606 -27306
rect 27664 -27506 28064 -27306
rect 28122 -27506 28522 -27306
rect 28580 -27506 28980 -27306
rect 29038 -27506 29438 -27306
rect 29496 -27506 29896 -27306
rect 29954 -27506 30354 -27306
rect 30412 -27506 30812 -27306
<< scnmos >>
rect 31662 2313 31692 2443
rect 31907 2313 31937 2443
rect 31991 2313 32021 2443
rect 32075 2313 32105 2443
rect 32159 2313 32189 2443
<< scpmoshvt >>
rect 31662 1993 31692 2193
rect 31907 1993 31937 2193
rect 31991 1993 32021 2193
rect 32075 1993 32105 2193
rect 32159 1993 32189 2193
<< pmoshvt >>
rect 15848 -207 16248 1393
rect 16306 -207 16706 1393
rect 16764 -207 17164 1393
rect 17222 -207 17622 1393
rect 17680 -207 18080 1393
rect 18138 -207 18538 1393
rect 18596 -207 18996 1393
rect 19054 -207 19454 1393
rect 19512 -207 19912 1393
rect 19970 -207 20370 1393
rect 20428 -207 20828 1393
rect 20886 -207 21286 1393
rect 21344 -207 21744 1393
rect 21802 -207 22202 1393
rect 22260 -207 22660 1393
rect 22718 -207 23118 1393
rect 23176 -207 23576 1393
rect 23634 -207 24034 1393
rect 26443 613 26843 1813
rect 26901 613 27301 1813
rect 27359 613 27759 1813
rect 27817 613 28217 1813
rect 28275 613 28675 1813
rect 28733 613 29133 1813
rect 29191 613 29591 1813
rect 29649 613 30049 1813
rect 30107 613 30507 1813
rect 30565 613 30965 1813
rect 11850 -5080 12250 -3480
rect 12308 -5080 12708 -3480
rect 12766 -5080 13166 -3480
rect 13224 -5080 13624 -3480
rect 13682 -5080 14082 -3480
rect 14140 -5080 14540 -3480
rect 14598 -5080 14998 -3480
rect 15056 -5080 15456 -3480
rect 15514 -5080 15914 -3480
rect 15972 -5080 16372 -3480
rect 16430 -5080 16830 -3480
rect 16888 -5080 17288 -3480
rect 17346 -5080 17746 -3480
rect 17804 -5080 18204 -3480
rect 18262 -5080 18662 -3480
rect 18720 -5080 19120 -3480
rect 19178 -5080 19578 -3480
rect 19636 -5080 20036 -3480
rect 11291 -7345 11691 -6145
rect 11749 -7345 12149 -6145
rect 12207 -7345 12607 -6145
rect 12665 -7345 13065 -6145
rect 13123 -7345 13523 -6145
rect 13581 -7345 13981 -6145
rect 14039 -7345 14439 -6145
rect 14497 -7345 14897 -6145
rect 14955 -7345 15355 -6145
rect 15413 -7345 15813 -6145
rect 16291 -7345 16691 -6145
rect 16749 -7345 17149 -6145
rect 17207 -7345 17607 -6145
rect 17665 -7345 18065 -6145
rect 18123 -7345 18523 -6145
rect 18581 -7345 18981 -6145
rect 19039 -7345 19439 -6145
rect 19497 -7345 19897 -6145
rect 19955 -7345 20355 -6145
rect 20413 -7345 20813 -6145
rect 26850 -5080 27250 -3480
rect 27308 -5080 27708 -3480
rect 27766 -5080 28166 -3480
rect 28224 -5080 28624 -3480
rect 28682 -5080 29082 -3480
rect 29140 -5080 29540 -3480
rect 29598 -5080 29998 -3480
rect 30056 -5080 30456 -3480
rect 30514 -5080 30914 -3480
rect 30972 -5080 31372 -3480
rect 31430 -5080 31830 -3480
rect 31888 -5080 32288 -3480
rect 32346 -5080 32746 -3480
rect 32804 -5080 33204 -3480
rect 33262 -5080 33662 -3480
rect 33720 -5080 34120 -3480
rect 34178 -5080 34578 -3480
rect 34636 -5080 35036 -3480
rect 26291 -7345 26691 -6145
rect 26749 -7345 27149 -6145
rect 27207 -7345 27607 -6145
rect 27665 -7345 28065 -6145
rect 28123 -7345 28523 -6145
rect 28581 -7345 28981 -6145
rect 29039 -7345 29439 -6145
rect 29497 -7345 29897 -6145
rect 29955 -7345 30355 -6145
rect 30413 -7345 30813 -6145
rect 31291 -7345 31691 -6145
rect 31749 -7345 32149 -6145
rect 32207 -7345 32607 -6145
rect 32665 -7345 33065 -6145
rect 33123 -7345 33523 -6145
rect 33581 -7345 33981 -6145
rect 34039 -7345 34439 -6145
rect 34497 -7345 34897 -6145
rect 34955 -7345 35355 -6145
rect 35413 -7345 35813 -6145
rect 15221 -15459 15621 -14259
rect 15679 -15459 16079 -14259
rect 16137 -15459 16537 -14259
rect 16595 -15459 16995 -14259
rect 17053 -15459 17453 -14259
rect 17511 -15459 17911 -14259
rect 17969 -15459 18369 -14259
rect 18427 -15459 18827 -14259
rect 18885 -15459 19285 -14259
rect 19343 -15459 19743 -14259
rect 20221 -15459 20621 -14259
rect 20679 -15459 21079 -14259
rect 21137 -15459 21537 -14259
rect 21595 -15459 21995 -14259
rect 22053 -15459 22453 -14259
rect 22511 -15459 22911 -14259
rect 22969 -15459 23369 -14259
rect 23427 -15459 23827 -14259
rect 23885 -15459 24285 -14259
rect 24343 -15459 24743 -14259
rect 15998 -18124 16398 -16524
rect 16456 -18124 16856 -16524
rect 16914 -18124 17314 -16524
rect 17372 -18124 17772 -16524
rect 17830 -18124 18230 -16524
rect 18288 -18124 18688 -16524
rect 18746 -18124 19146 -16524
rect 19204 -18124 19604 -16524
rect 19662 -18124 20062 -16524
rect 20120 -18124 20520 -16524
rect 20578 -18124 20978 -16524
rect 21036 -18124 21436 -16524
rect 21494 -18124 21894 -16524
rect 21952 -18124 22352 -16524
rect 22410 -18124 22810 -16524
rect 22868 -18124 23268 -16524
rect 23326 -18124 23726 -16524
rect 23784 -18124 24184 -16524
rect 30221 -15459 30621 -14259
rect 30679 -15459 31079 -14259
rect 31137 -15459 31537 -14259
rect 31595 -15459 31995 -14259
rect 32053 -15459 32453 -14259
rect 32511 -15459 32911 -14259
rect 32969 -15459 33369 -14259
rect 33427 -15459 33827 -14259
rect 33885 -15459 34285 -14259
rect 34343 -15459 34743 -14259
rect 35221 -15459 35621 -14259
rect 35679 -15459 36079 -14259
rect 36137 -15459 36537 -14259
rect 36595 -15459 36995 -14259
rect 37053 -15459 37453 -14259
rect 37511 -15459 37911 -14259
rect 37969 -15459 38369 -14259
rect 38427 -15459 38827 -14259
rect 38885 -15459 39285 -14259
rect 39343 -15459 39743 -14259
rect 30998 -18124 31398 -16524
rect 31456 -18124 31856 -16524
rect 31914 -18124 32314 -16524
rect 32372 -18124 32772 -16524
rect 32830 -18124 33230 -16524
rect 33288 -18124 33688 -16524
rect 33746 -18124 34146 -16524
rect 34204 -18124 34604 -16524
rect 34662 -18124 35062 -16524
rect 35120 -18124 35520 -16524
rect 35578 -18124 35978 -16524
rect 36036 -18124 36436 -16524
rect 36494 -18124 36894 -16524
rect 36952 -18124 37352 -16524
rect 37410 -18124 37810 -16524
rect 37868 -18124 38268 -16524
rect 38326 -18124 38726 -16524
rect 38784 -18124 39184 -16524
rect 11850 -23080 12250 -21480
rect 12308 -23080 12708 -21480
rect 12766 -23080 13166 -21480
rect 13224 -23080 13624 -21480
rect 13682 -23080 14082 -21480
rect 14140 -23080 14540 -21480
rect 14598 -23080 14998 -21480
rect 15056 -23080 15456 -21480
rect 15514 -23080 15914 -21480
rect 15972 -23080 16372 -21480
rect 16430 -23080 16830 -21480
rect 16888 -23080 17288 -21480
rect 17346 -23080 17746 -21480
rect 17804 -23080 18204 -21480
rect 18262 -23080 18662 -21480
rect 18720 -23080 19120 -21480
rect 19178 -23080 19578 -21480
rect 19636 -23080 20036 -21480
rect 11291 -25345 11691 -24145
rect 11749 -25345 12149 -24145
rect 12207 -25345 12607 -24145
rect 12665 -25345 13065 -24145
rect 13123 -25345 13523 -24145
rect 13581 -25345 13981 -24145
rect 14039 -25345 14439 -24145
rect 14497 -25345 14897 -24145
rect 14955 -25345 15355 -24145
rect 15413 -25345 15813 -24145
rect 16291 -25345 16691 -24145
rect 16749 -25345 17149 -24145
rect 17207 -25345 17607 -24145
rect 17665 -25345 18065 -24145
rect 18123 -25345 18523 -24145
rect 18581 -25345 18981 -24145
rect 19039 -25345 19439 -24145
rect 19497 -25345 19897 -24145
rect 19955 -25345 20355 -24145
rect 20413 -25345 20813 -24145
rect 26850 -23080 27250 -21480
rect 27308 -23080 27708 -21480
rect 27766 -23080 28166 -21480
rect 28224 -23080 28624 -21480
rect 28682 -23080 29082 -21480
rect 29140 -23080 29540 -21480
rect 29598 -23080 29998 -21480
rect 30056 -23080 30456 -21480
rect 30514 -23080 30914 -21480
rect 30972 -23080 31372 -21480
rect 31430 -23080 31830 -21480
rect 31888 -23080 32288 -21480
rect 32346 -23080 32746 -21480
rect 32804 -23080 33204 -21480
rect 33262 -23080 33662 -21480
rect 33720 -23080 34120 -21480
rect 34178 -23080 34578 -21480
rect 34636 -23080 35036 -21480
rect 26291 -25345 26691 -24145
rect 26749 -25345 27149 -24145
rect 27207 -25345 27607 -24145
rect 27665 -25345 28065 -24145
rect 28123 -25345 28523 -24145
rect 28581 -25345 28981 -24145
rect 29039 -25345 29439 -24145
rect 29497 -25345 29897 -24145
rect 29955 -25345 30355 -24145
rect 30413 -25345 30813 -24145
rect 31291 -25345 31691 -24145
rect 31749 -25345 32149 -24145
rect 32207 -25345 32607 -24145
rect 32665 -25345 33065 -24145
rect 33123 -25345 33523 -24145
rect 33581 -25345 33981 -24145
rect 34039 -25345 34439 -24145
rect 34497 -25345 34897 -24145
rect 34955 -25345 35355 -24145
rect 35413 -25345 35813 -24145
<< ndiff >>
rect 17622 3232 17680 3244
rect 17622 3056 17634 3232
rect 17668 3056 17680 3232
rect 17622 3044 17680 3056
rect 18080 3232 18138 3244
rect 18080 3056 18092 3232
rect 18126 3056 18138 3232
rect 18080 3044 18138 3056
rect 18538 3232 18596 3244
rect 18538 3056 18550 3232
rect 18584 3056 18596 3232
rect 18538 3044 18596 3056
rect 18996 3232 19054 3244
rect 18996 3056 19008 3232
rect 19042 3056 19054 3232
rect 18996 3044 19054 3056
rect 19454 3232 19512 3244
rect 19454 3056 19466 3232
rect 19500 3056 19512 3232
rect 19454 3044 19512 3056
rect 19912 3232 19970 3244
rect 19912 3056 19924 3232
rect 19958 3056 19970 3232
rect 19912 3044 19970 3056
rect 20370 3232 20428 3244
rect 20370 3056 20382 3232
rect 20416 3056 20428 3232
rect 20370 3044 20428 3056
rect 20828 3232 20886 3244
rect 20828 3056 20840 3232
rect 20874 3056 20886 3232
rect 20828 3044 20886 3056
rect 21286 3232 21344 3244
rect 21286 3056 21298 3232
rect 21332 3056 21344 3232
rect 21286 3044 21344 3056
rect 21744 3232 21802 3244
rect 21744 3056 21756 3232
rect 21790 3056 21802 3232
rect 21744 3044 21802 3056
rect 22202 3232 22260 3244
rect 22202 3056 22214 3232
rect 22248 3056 22260 3232
rect 22202 3044 22260 3056
rect 26384 3232 26442 3244
rect 26384 3056 26396 3232
rect 26430 3056 26442 3232
rect 26384 3044 26442 3056
rect 26842 3232 26900 3244
rect 26842 3056 26854 3232
rect 26888 3056 26900 3232
rect 26842 3044 26900 3056
rect 27300 3232 27358 3244
rect 27300 3056 27312 3232
rect 27346 3056 27358 3232
rect 27300 3044 27358 3056
rect 27758 3232 27816 3244
rect 27758 3056 27770 3232
rect 27804 3056 27816 3232
rect 27758 3044 27816 3056
rect 28216 3232 28274 3244
rect 28216 3056 28228 3232
rect 28262 3056 28274 3232
rect 28216 3044 28274 3056
rect 28674 3232 28732 3244
rect 28674 3056 28686 3232
rect 28720 3056 28732 3232
rect 28674 3044 28732 3056
rect 29132 3232 29190 3244
rect 29132 3056 29144 3232
rect 29178 3056 29190 3232
rect 29132 3044 29190 3056
rect 29590 3232 29648 3244
rect 29590 3056 29602 3232
rect 29636 3056 29648 3232
rect 29590 3044 29648 3056
rect 30048 3232 30106 3244
rect 30048 3056 30060 3232
rect 30094 3056 30106 3232
rect 30048 3044 30106 3056
rect 30506 3232 30564 3244
rect 30506 3056 30518 3232
rect 30552 3056 30564 3232
rect 30506 3044 30564 3056
rect 30964 3232 31022 3244
rect 30964 3056 30976 3232
rect 31010 3056 31022 3232
rect 30964 3044 31022 3056
rect 31610 2427 31662 2443
rect 31610 2393 31618 2427
rect 31652 2393 31662 2427
rect 31610 2359 31662 2393
rect 31610 2325 31618 2359
rect 31652 2325 31662 2359
rect 31610 2313 31662 2325
rect 31692 2427 31744 2443
rect 31692 2393 31702 2427
rect 31736 2393 31744 2427
rect 31692 2359 31744 2393
rect 31692 2325 31702 2359
rect 31736 2325 31744 2359
rect 31692 2313 31744 2325
rect 31855 2431 31907 2443
rect 31855 2397 31863 2431
rect 31897 2397 31907 2431
rect 31855 2313 31907 2397
rect 31937 2423 31991 2443
rect 31937 2389 31947 2423
rect 31981 2389 31991 2423
rect 31937 2313 31991 2389
rect 32021 2431 32075 2443
rect 32021 2397 32031 2431
rect 32065 2397 32075 2431
rect 32021 2313 32075 2397
rect 32105 2423 32159 2443
rect 32105 2389 32115 2423
rect 32149 2389 32159 2423
rect 32105 2313 32159 2389
rect 32189 2430 32241 2443
rect 32189 2396 32199 2430
rect 32233 2396 32241 2430
rect 32189 2313 32241 2396
rect 11232 -8650 11290 -8638
rect 11232 -8826 11244 -8650
rect 11278 -8826 11290 -8650
rect 11232 -8838 11290 -8826
rect 11690 -8650 11748 -8638
rect 11690 -8826 11702 -8650
rect 11736 -8826 11748 -8650
rect 11690 -8838 11748 -8826
rect 12148 -8650 12206 -8638
rect 12148 -8826 12160 -8650
rect 12194 -8826 12206 -8650
rect 12148 -8838 12206 -8826
rect 12606 -8650 12664 -8638
rect 12606 -8826 12618 -8650
rect 12652 -8826 12664 -8650
rect 12606 -8838 12664 -8826
rect 13064 -8650 13122 -8638
rect 13064 -8826 13076 -8650
rect 13110 -8826 13122 -8650
rect 13064 -8838 13122 -8826
rect 13522 -8650 13580 -8638
rect 13522 -8826 13534 -8650
rect 13568 -8826 13580 -8650
rect 13522 -8838 13580 -8826
rect 13980 -8650 14038 -8638
rect 13980 -8826 13992 -8650
rect 14026 -8826 14038 -8650
rect 13980 -8838 14038 -8826
rect 14438 -8650 14496 -8638
rect 14438 -8826 14450 -8650
rect 14484 -8826 14496 -8650
rect 14438 -8838 14496 -8826
rect 14896 -8650 14954 -8638
rect 14896 -8826 14908 -8650
rect 14942 -8826 14954 -8650
rect 14896 -8838 14954 -8826
rect 15354 -8650 15412 -8638
rect 15354 -8826 15366 -8650
rect 15400 -8826 15412 -8650
rect 15354 -8838 15412 -8826
rect 15812 -8650 15870 -8638
rect 15812 -8826 15824 -8650
rect 15858 -8826 15870 -8650
rect 15812 -8838 15870 -8826
rect 16232 -8650 16290 -8638
rect 16232 -8826 16244 -8650
rect 16278 -8826 16290 -8650
rect 16232 -8838 16290 -8826
rect 16690 -8650 16748 -8638
rect 16690 -8826 16702 -8650
rect 16736 -8826 16748 -8650
rect 16690 -8838 16748 -8826
rect 17148 -8650 17206 -8638
rect 17148 -8826 17160 -8650
rect 17194 -8826 17206 -8650
rect 17148 -8838 17206 -8826
rect 17606 -8650 17664 -8638
rect 17606 -8826 17618 -8650
rect 17652 -8826 17664 -8650
rect 17606 -8838 17664 -8826
rect 18064 -8650 18122 -8638
rect 18064 -8826 18076 -8650
rect 18110 -8826 18122 -8650
rect 18064 -8838 18122 -8826
rect 18522 -8650 18580 -8638
rect 18522 -8826 18534 -8650
rect 18568 -8826 18580 -8650
rect 18522 -8838 18580 -8826
rect 18980 -8650 19038 -8638
rect 18980 -8826 18992 -8650
rect 19026 -8826 19038 -8650
rect 18980 -8838 19038 -8826
rect 19438 -8650 19496 -8638
rect 19438 -8826 19450 -8650
rect 19484 -8826 19496 -8650
rect 19438 -8838 19496 -8826
rect 19896 -8650 19954 -8638
rect 19896 -8826 19908 -8650
rect 19942 -8826 19954 -8650
rect 19896 -8838 19954 -8826
rect 20354 -8650 20412 -8638
rect 20354 -8826 20366 -8650
rect 20400 -8826 20412 -8650
rect 20354 -8838 20412 -8826
rect 20812 -8650 20870 -8638
rect 20812 -8826 20824 -8650
rect 20858 -8826 20870 -8650
rect 20812 -8838 20870 -8826
rect 11232 -9318 11290 -9306
rect 11232 -9494 11244 -9318
rect 11278 -9494 11290 -9318
rect 11232 -9506 11290 -9494
rect 11690 -9318 11748 -9306
rect 11690 -9494 11702 -9318
rect 11736 -9494 11748 -9318
rect 11690 -9506 11748 -9494
rect 12148 -9318 12206 -9306
rect 12148 -9494 12160 -9318
rect 12194 -9494 12206 -9318
rect 12148 -9506 12206 -9494
rect 12606 -9318 12664 -9306
rect 12606 -9494 12618 -9318
rect 12652 -9494 12664 -9318
rect 12606 -9506 12664 -9494
rect 13064 -9318 13122 -9306
rect 13064 -9494 13076 -9318
rect 13110 -9494 13122 -9318
rect 13064 -9506 13122 -9494
rect 13522 -9318 13580 -9306
rect 13522 -9494 13534 -9318
rect 13568 -9494 13580 -9318
rect 13522 -9506 13580 -9494
rect 13980 -9318 14038 -9306
rect 13980 -9494 13992 -9318
rect 14026 -9494 14038 -9318
rect 13980 -9506 14038 -9494
rect 14438 -9318 14496 -9306
rect 14438 -9494 14450 -9318
rect 14484 -9494 14496 -9318
rect 14438 -9506 14496 -9494
rect 14896 -9318 14954 -9306
rect 14896 -9494 14908 -9318
rect 14942 -9494 14954 -9318
rect 14896 -9506 14954 -9494
rect 15354 -9318 15412 -9306
rect 15354 -9494 15366 -9318
rect 15400 -9494 15412 -9318
rect 15354 -9506 15412 -9494
rect 15812 -9318 15870 -9306
rect 15812 -9494 15824 -9318
rect 15858 -9494 15870 -9318
rect 15812 -9506 15870 -9494
rect 26232 -8650 26290 -8638
rect 26232 -8826 26244 -8650
rect 26278 -8826 26290 -8650
rect 26232 -8838 26290 -8826
rect 26690 -8650 26748 -8638
rect 26690 -8826 26702 -8650
rect 26736 -8826 26748 -8650
rect 26690 -8838 26748 -8826
rect 27148 -8650 27206 -8638
rect 27148 -8826 27160 -8650
rect 27194 -8826 27206 -8650
rect 27148 -8838 27206 -8826
rect 27606 -8650 27664 -8638
rect 27606 -8826 27618 -8650
rect 27652 -8826 27664 -8650
rect 27606 -8838 27664 -8826
rect 28064 -8650 28122 -8638
rect 28064 -8826 28076 -8650
rect 28110 -8826 28122 -8650
rect 28064 -8838 28122 -8826
rect 28522 -8650 28580 -8638
rect 28522 -8826 28534 -8650
rect 28568 -8826 28580 -8650
rect 28522 -8838 28580 -8826
rect 28980 -8650 29038 -8638
rect 28980 -8826 28992 -8650
rect 29026 -8826 29038 -8650
rect 28980 -8838 29038 -8826
rect 29438 -8650 29496 -8638
rect 29438 -8826 29450 -8650
rect 29484 -8826 29496 -8650
rect 29438 -8838 29496 -8826
rect 29896 -8650 29954 -8638
rect 29896 -8826 29908 -8650
rect 29942 -8826 29954 -8650
rect 29896 -8838 29954 -8826
rect 30354 -8650 30412 -8638
rect 30354 -8826 30366 -8650
rect 30400 -8826 30412 -8650
rect 30354 -8838 30412 -8826
rect 30812 -8650 30870 -8638
rect 30812 -8826 30824 -8650
rect 30858 -8826 30870 -8650
rect 30812 -8838 30870 -8826
rect 31232 -8650 31290 -8638
rect 31232 -8826 31244 -8650
rect 31278 -8826 31290 -8650
rect 31232 -8838 31290 -8826
rect 31690 -8650 31748 -8638
rect 31690 -8826 31702 -8650
rect 31736 -8826 31748 -8650
rect 31690 -8838 31748 -8826
rect 32148 -8650 32206 -8638
rect 32148 -8826 32160 -8650
rect 32194 -8826 32206 -8650
rect 32148 -8838 32206 -8826
rect 32606 -8650 32664 -8638
rect 32606 -8826 32618 -8650
rect 32652 -8826 32664 -8650
rect 32606 -8838 32664 -8826
rect 33064 -8650 33122 -8638
rect 33064 -8826 33076 -8650
rect 33110 -8826 33122 -8650
rect 33064 -8838 33122 -8826
rect 33522 -8650 33580 -8638
rect 33522 -8826 33534 -8650
rect 33568 -8826 33580 -8650
rect 33522 -8838 33580 -8826
rect 33980 -8650 34038 -8638
rect 33980 -8826 33992 -8650
rect 34026 -8826 34038 -8650
rect 33980 -8838 34038 -8826
rect 34438 -8650 34496 -8638
rect 34438 -8826 34450 -8650
rect 34484 -8826 34496 -8650
rect 34438 -8838 34496 -8826
rect 34896 -8650 34954 -8638
rect 34896 -8826 34908 -8650
rect 34942 -8826 34954 -8650
rect 34896 -8838 34954 -8826
rect 35354 -8650 35412 -8638
rect 35354 -8826 35366 -8650
rect 35400 -8826 35412 -8650
rect 35354 -8838 35412 -8826
rect 35812 -8650 35870 -8638
rect 35812 -8826 35824 -8650
rect 35858 -8826 35870 -8650
rect 35812 -8838 35870 -8826
rect 26232 -9318 26290 -9306
rect 26232 -9494 26244 -9318
rect 26278 -9494 26290 -9318
rect 26232 -9506 26290 -9494
rect 26690 -9318 26748 -9306
rect 26690 -9494 26702 -9318
rect 26736 -9494 26748 -9318
rect 26690 -9506 26748 -9494
rect 27148 -9318 27206 -9306
rect 27148 -9494 27160 -9318
rect 27194 -9494 27206 -9318
rect 27148 -9506 27206 -9494
rect 27606 -9318 27664 -9306
rect 27606 -9494 27618 -9318
rect 27652 -9494 27664 -9318
rect 27606 -9506 27664 -9494
rect 28064 -9318 28122 -9306
rect 28064 -9494 28076 -9318
rect 28110 -9494 28122 -9318
rect 28064 -9506 28122 -9494
rect 28522 -9318 28580 -9306
rect 28522 -9494 28534 -9318
rect 28568 -9494 28580 -9318
rect 28522 -9506 28580 -9494
rect 28980 -9318 29038 -9306
rect 28980 -9494 28992 -9318
rect 29026 -9494 29038 -9318
rect 28980 -9506 29038 -9494
rect 29438 -9318 29496 -9306
rect 29438 -9494 29450 -9318
rect 29484 -9494 29496 -9318
rect 29438 -9506 29496 -9494
rect 29896 -9318 29954 -9306
rect 29896 -9494 29908 -9318
rect 29942 -9494 29954 -9318
rect 29896 -9506 29954 -9494
rect 30354 -9318 30412 -9306
rect 30354 -9494 30366 -9318
rect 30400 -9494 30412 -9318
rect 30354 -9506 30412 -9494
rect 30812 -9318 30870 -9306
rect 30812 -9494 30824 -9318
rect 30858 -9494 30870 -9318
rect 30812 -9506 30870 -9494
rect 20164 -12110 20222 -12098
rect 20164 -12286 20176 -12110
rect 20210 -12286 20222 -12110
rect 20164 -12298 20222 -12286
rect 20622 -12110 20680 -12098
rect 20622 -12286 20634 -12110
rect 20668 -12286 20680 -12110
rect 20622 -12298 20680 -12286
rect 21080 -12110 21138 -12098
rect 21080 -12286 21092 -12110
rect 21126 -12286 21138 -12110
rect 21080 -12298 21138 -12286
rect 21538 -12110 21596 -12098
rect 21538 -12286 21550 -12110
rect 21584 -12286 21596 -12110
rect 21538 -12298 21596 -12286
rect 21996 -12110 22054 -12098
rect 21996 -12286 22008 -12110
rect 22042 -12286 22054 -12110
rect 21996 -12298 22054 -12286
rect 22454 -12110 22512 -12098
rect 22454 -12286 22466 -12110
rect 22500 -12286 22512 -12110
rect 22454 -12298 22512 -12286
rect 22912 -12110 22970 -12098
rect 22912 -12286 22924 -12110
rect 22958 -12286 22970 -12110
rect 22912 -12298 22970 -12286
rect 23370 -12110 23428 -12098
rect 23370 -12286 23382 -12110
rect 23416 -12286 23428 -12110
rect 23370 -12298 23428 -12286
rect 23828 -12110 23886 -12098
rect 23828 -12286 23840 -12110
rect 23874 -12286 23886 -12110
rect 23828 -12298 23886 -12286
rect 24286 -12110 24344 -12098
rect 24286 -12286 24298 -12110
rect 24332 -12286 24344 -12110
rect 24286 -12298 24344 -12286
rect 24744 -12110 24802 -12098
rect 24744 -12286 24756 -12110
rect 24790 -12286 24802 -12110
rect 24744 -12298 24802 -12286
rect 15164 -12778 15222 -12766
rect 15164 -12954 15176 -12778
rect 15210 -12954 15222 -12778
rect 15164 -12966 15222 -12954
rect 15622 -12778 15680 -12766
rect 15622 -12954 15634 -12778
rect 15668 -12954 15680 -12778
rect 15622 -12966 15680 -12954
rect 16080 -12778 16138 -12766
rect 16080 -12954 16092 -12778
rect 16126 -12954 16138 -12778
rect 16080 -12966 16138 -12954
rect 16538 -12778 16596 -12766
rect 16538 -12954 16550 -12778
rect 16584 -12954 16596 -12778
rect 16538 -12966 16596 -12954
rect 16996 -12778 17054 -12766
rect 16996 -12954 17008 -12778
rect 17042 -12954 17054 -12778
rect 16996 -12966 17054 -12954
rect 17454 -12778 17512 -12766
rect 17454 -12954 17466 -12778
rect 17500 -12954 17512 -12778
rect 17454 -12966 17512 -12954
rect 17912 -12778 17970 -12766
rect 17912 -12954 17924 -12778
rect 17958 -12954 17970 -12778
rect 17912 -12966 17970 -12954
rect 18370 -12778 18428 -12766
rect 18370 -12954 18382 -12778
rect 18416 -12954 18428 -12778
rect 18370 -12966 18428 -12954
rect 18828 -12778 18886 -12766
rect 18828 -12954 18840 -12778
rect 18874 -12954 18886 -12778
rect 18828 -12966 18886 -12954
rect 19286 -12778 19344 -12766
rect 19286 -12954 19298 -12778
rect 19332 -12954 19344 -12778
rect 19286 -12966 19344 -12954
rect 19744 -12778 19802 -12766
rect 19744 -12954 19756 -12778
rect 19790 -12954 19802 -12778
rect 19744 -12966 19802 -12954
rect 20164 -12778 20222 -12766
rect 20164 -12954 20176 -12778
rect 20210 -12954 20222 -12778
rect 20164 -12966 20222 -12954
rect 20622 -12778 20680 -12766
rect 20622 -12954 20634 -12778
rect 20668 -12954 20680 -12778
rect 20622 -12966 20680 -12954
rect 21080 -12778 21138 -12766
rect 21080 -12954 21092 -12778
rect 21126 -12954 21138 -12778
rect 21080 -12966 21138 -12954
rect 21538 -12778 21596 -12766
rect 21538 -12954 21550 -12778
rect 21584 -12954 21596 -12778
rect 21538 -12966 21596 -12954
rect 21996 -12778 22054 -12766
rect 21996 -12954 22008 -12778
rect 22042 -12954 22054 -12778
rect 21996 -12966 22054 -12954
rect 22454 -12778 22512 -12766
rect 22454 -12954 22466 -12778
rect 22500 -12954 22512 -12778
rect 22454 -12966 22512 -12954
rect 22912 -12778 22970 -12766
rect 22912 -12954 22924 -12778
rect 22958 -12954 22970 -12778
rect 22912 -12966 22970 -12954
rect 23370 -12778 23428 -12766
rect 23370 -12954 23382 -12778
rect 23416 -12954 23428 -12778
rect 23370 -12966 23428 -12954
rect 23828 -12778 23886 -12766
rect 23828 -12954 23840 -12778
rect 23874 -12954 23886 -12778
rect 23828 -12966 23886 -12954
rect 24286 -12778 24344 -12766
rect 24286 -12954 24298 -12778
rect 24332 -12954 24344 -12778
rect 24286 -12966 24344 -12954
rect 24744 -12778 24802 -12766
rect 24744 -12954 24756 -12778
rect 24790 -12954 24802 -12778
rect 24744 -12966 24802 -12954
rect 35164 -12110 35222 -12098
rect 35164 -12286 35176 -12110
rect 35210 -12286 35222 -12110
rect 35164 -12298 35222 -12286
rect 35622 -12110 35680 -12098
rect 35622 -12286 35634 -12110
rect 35668 -12286 35680 -12110
rect 35622 -12298 35680 -12286
rect 36080 -12110 36138 -12098
rect 36080 -12286 36092 -12110
rect 36126 -12286 36138 -12110
rect 36080 -12298 36138 -12286
rect 36538 -12110 36596 -12098
rect 36538 -12286 36550 -12110
rect 36584 -12286 36596 -12110
rect 36538 -12298 36596 -12286
rect 36996 -12110 37054 -12098
rect 36996 -12286 37008 -12110
rect 37042 -12286 37054 -12110
rect 36996 -12298 37054 -12286
rect 37454 -12110 37512 -12098
rect 37454 -12286 37466 -12110
rect 37500 -12286 37512 -12110
rect 37454 -12298 37512 -12286
rect 37912 -12110 37970 -12098
rect 37912 -12286 37924 -12110
rect 37958 -12286 37970 -12110
rect 37912 -12298 37970 -12286
rect 38370 -12110 38428 -12098
rect 38370 -12286 38382 -12110
rect 38416 -12286 38428 -12110
rect 38370 -12298 38428 -12286
rect 38828 -12110 38886 -12098
rect 38828 -12286 38840 -12110
rect 38874 -12286 38886 -12110
rect 38828 -12298 38886 -12286
rect 39286 -12110 39344 -12098
rect 39286 -12286 39298 -12110
rect 39332 -12286 39344 -12110
rect 39286 -12298 39344 -12286
rect 39744 -12110 39802 -12098
rect 39744 -12286 39756 -12110
rect 39790 -12286 39802 -12110
rect 39744 -12298 39802 -12286
rect 30164 -12778 30222 -12766
rect 30164 -12954 30176 -12778
rect 30210 -12954 30222 -12778
rect 30164 -12966 30222 -12954
rect 30622 -12778 30680 -12766
rect 30622 -12954 30634 -12778
rect 30668 -12954 30680 -12778
rect 30622 -12966 30680 -12954
rect 31080 -12778 31138 -12766
rect 31080 -12954 31092 -12778
rect 31126 -12954 31138 -12778
rect 31080 -12966 31138 -12954
rect 31538 -12778 31596 -12766
rect 31538 -12954 31550 -12778
rect 31584 -12954 31596 -12778
rect 31538 -12966 31596 -12954
rect 31996 -12778 32054 -12766
rect 31996 -12954 32008 -12778
rect 32042 -12954 32054 -12778
rect 31996 -12966 32054 -12954
rect 32454 -12778 32512 -12766
rect 32454 -12954 32466 -12778
rect 32500 -12954 32512 -12778
rect 32454 -12966 32512 -12954
rect 32912 -12778 32970 -12766
rect 32912 -12954 32924 -12778
rect 32958 -12954 32970 -12778
rect 32912 -12966 32970 -12954
rect 33370 -12778 33428 -12766
rect 33370 -12954 33382 -12778
rect 33416 -12954 33428 -12778
rect 33370 -12966 33428 -12954
rect 33828 -12778 33886 -12766
rect 33828 -12954 33840 -12778
rect 33874 -12954 33886 -12778
rect 33828 -12966 33886 -12954
rect 34286 -12778 34344 -12766
rect 34286 -12954 34298 -12778
rect 34332 -12954 34344 -12778
rect 34286 -12966 34344 -12954
rect 34744 -12778 34802 -12766
rect 34744 -12954 34756 -12778
rect 34790 -12954 34802 -12778
rect 34744 -12966 34802 -12954
rect 35164 -12778 35222 -12766
rect 35164 -12954 35176 -12778
rect 35210 -12954 35222 -12778
rect 35164 -12966 35222 -12954
rect 35622 -12778 35680 -12766
rect 35622 -12954 35634 -12778
rect 35668 -12954 35680 -12778
rect 35622 -12966 35680 -12954
rect 36080 -12778 36138 -12766
rect 36080 -12954 36092 -12778
rect 36126 -12954 36138 -12778
rect 36080 -12966 36138 -12954
rect 36538 -12778 36596 -12766
rect 36538 -12954 36550 -12778
rect 36584 -12954 36596 -12778
rect 36538 -12966 36596 -12954
rect 36996 -12778 37054 -12766
rect 36996 -12954 37008 -12778
rect 37042 -12954 37054 -12778
rect 36996 -12966 37054 -12954
rect 37454 -12778 37512 -12766
rect 37454 -12954 37466 -12778
rect 37500 -12954 37512 -12778
rect 37454 -12966 37512 -12954
rect 37912 -12778 37970 -12766
rect 37912 -12954 37924 -12778
rect 37958 -12954 37970 -12778
rect 37912 -12966 37970 -12954
rect 38370 -12778 38428 -12766
rect 38370 -12954 38382 -12778
rect 38416 -12954 38428 -12778
rect 38370 -12966 38428 -12954
rect 38828 -12778 38886 -12766
rect 38828 -12954 38840 -12778
rect 38874 -12954 38886 -12778
rect 38828 -12966 38886 -12954
rect 39286 -12778 39344 -12766
rect 39286 -12954 39298 -12778
rect 39332 -12954 39344 -12778
rect 39286 -12966 39344 -12954
rect 39744 -12778 39802 -12766
rect 39744 -12954 39756 -12778
rect 39790 -12954 39802 -12778
rect 39744 -12966 39802 -12954
rect 11232 -26650 11290 -26638
rect 11232 -26826 11244 -26650
rect 11278 -26826 11290 -26650
rect 11232 -26838 11290 -26826
rect 11690 -26650 11748 -26638
rect 11690 -26826 11702 -26650
rect 11736 -26826 11748 -26650
rect 11690 -26838 11748 -26826
rect 12148 -26650 12206 -26638
rect 12148 -26826 12160 -26650
rect 12194 -26826 12206 -26650
rect 12148 -26838 12206 -26826
rect 12606 -26650 12664 -26638
rect 12606 -26826 12618 -26650
rect 12652 -26826 12664 -26650
rect 12606 -26838 12664 -26826
rect 13064 -26650 13122 -26638
rect 13064 -26826 13076 -26650
rect 13110 -26826 13122 -26650
rect 13064 -26838 13122 -26826
rect 13522 -26650 13580 -26638
rect 13522 -26826 13534 -26650
rect 13568 -26826 13580 -26650
rect 13522 -26838 13580 -26826
rect 13980 -26650 14038 -26638
rect 13980 -26826 13992 -26650
rect 14026 -26826 14038 -26650
rect 13980 -26838 14038 -26826
rect 14438 -26650 14496 -26638
rect 14438 -26826 14450 -26650
rect 14484 -26826 14496 -26650
rect 14438 -26838 14496 -26826
rect 14896 -26650 14954 -26638
rect 14896 -26826 14908 -26650
rect 14942 -26826 14954 -26650
rect 14896 -26838 14954 -26826
rect 15354 -26650 15412 -26638
rect 15354 -26826 15366 -26650
rect 15400 -26826 15412 -26650
rect 15354 -26838 15412 -26826
rect 15812 -26650 15870 -26638
rect 15812 -26826 15824 -26650
rect 15858 -26826 15870 -26650
rect 15812 -26838 15870 -26826
rect 16232 -26650 16290 -26638
rect 16232 -26826 16244 -26650
rect 16278 -26826 16290 -26650
rect 16232 -26838 16290 -26826
rect 16690 -26650 16748 -26638
rect 16690 -26826 16702 -26650
rect 16736 -26826 16748 -26650
rect 16690 -26838 16748 -26826
rect 17148 -26650 17206 -26638
rect 17148 -26826 17160 -26650
rect 17194 -26826 17206 -26650
rect 17148 -26838 17206 -26826
rect 17606 -26650 17664 -26638
rect 17606 -26826 17618 -26650
rect 17652 -26826 17664 -26650
rect 17606 -26838 17664 -26826
rect 18064 -26650 18122 -26638
rect 18064 -26826 18076 -26650
rect 18110 -26826 18122 -26650
rect 18064 -26838 18122 -26826
rect 18522 -26650 18580 -26638
rect 18522 -26826 18534 -26650
rect 18568 -26826 18580 -26650
rect 18522 -26838 18580 -26826
rect 18980 -26650 19038 -26638
rect 18980 -26826 18992 -26650
rect 19026 -26826 19038 -26650
rect 18980 -26838 19038 -26826
rect 19438 -26650 19496 -26638
rect 19438 -26826 19450 -26650
rect 19484 -26826 19496 -26650
rect 19438 -26838 19496 -26826
rect 19896 -26650 19954 -26638
rect 19896 -26826 19908 -26650
rect 19942 -26826 19954 -26650
rect 19896 -26838 19954 -26826
rect 20354 -26650 20412 -26638
rect 20354 -26826 20366 -26650
rect 20400 -26826 20412 -26650
rect 20354 -26838 20412 -26826
rect 20812 -26650 20870 -26638
rect 20812 -26826 20824 -26650
rect 20858 -26826 20870 -26650
rect 20812 -26838 20870 -26826
rect 11232 -27318 11290 -27306
rect 11232 -27494 11244 -27318
rect 11278 -27494 11290 -27318
rect 11232 -27506 11290 -27494
rect 11690 -27318 11748 -27306
rect 11690 -27494 11702 -27318
rect 11736 -27494 11748 -27318
rect 11690 -27506 11748 -27494
rect 12148 -27318 12206 -27306
rect 12148 -27494 12160 -27318
rect 12194 -27494 12206 -27318
rect 12148 -27506 12206 -27494
rect 12606 -27318 12664 -27306
rect 12606 -27494 12618 -27318
rect 12652 -27494 12664 -27318
rect 12606 -27506 12664 -27494
rect 13064 -27318 13122 -27306
rect 13064 -27494 13076 -27318
rect 13110 -27494 13122 -27318
rect 13064 -27506 13122 -27494
rect 13522 -27318 13580 -27306
rect 13522 -27494 13534 -27318
rect 13568 -27494 13580 -27318
rect 13522 -27506 13580 -27494
rect 13980 -27318 14038 -27306
rect 13980 -27494 13992 -27318
rect 14026 -27494 14038 -27318
rect 13980 -27506 14038 -27494
rect 14438 -27318 14496 -27306
rect 14438 -27494 14450 -27318
rect 14484 -27494 14496 -27318
rect 14438 -27506 14496 -27494
rect 14896 -27318 14954 -27306
rect 14896 -27494 14908 -27318
rect 14942 -27494 14954 -27318
rect 14896 -27506 14954 -27494
rect 15354 -27318 15412 -27306
rect 15354 -27494 15366 -27318
rect 15400 -27494 15412 -27318
rect 15354 -27506 15412 -27494
rect 15812 -27318 15870 -27306
rect 15812 -27494 15824 -27318
rect 15858 -27494 15870 -27318
rect 15812 -27506 15870 -27494
rect 26232 -26650 26290 -26638
rect 26232 -26826 26244 -26650
rect 26278 -26826 26290 -26650
rect 26232 -26838 26290 -26826
rect 26690 -26650 26748 -26638
rect 26690 -26826 26702 -26650
rect 26736 -26826 26748 -26650
rect 26690 -26838 26748 -26826
rect 27148 -26650 27206 -26638
rect 27148 -26826 27160 -26650
rect 27194 -26826 27206 -26650
rect 27148 -26838 27206 -26826
rect 27606 -26650 27664 -26638
rect 27606 -26826 27618 -26650
rect 27652 -26826 27664 -26650
rect 27606 -26838 27664 -26826
rect 28064 -26650 28122 -26638
rect 28064 -26826 28076 -26650
rect 28110 -26826 28122 -26650
rect 28064 -26838 28122 -26826
rect 28522 -26650 28580 -26638
rect 28522 -26826 28534 -26650
rect 28568 -26826 28580 -26650
rect 28522 -26838 28580 -26826
rect 28980 -26650 29038 -26638
rect 28980 -26826 28992 -26650
rect 29026 -26826 29038 -26650
rect 28980 -26838 29038 -26826
rect 29438 -26650 29496 -26638
rect 29438 -26826 29450 -26650
rect 29484 -26826 29496 -26650
rect 29438 -26838 29496 -26826
rect 29896 -26650 29954 -26638
rect 29896 -26826 29908 -26650
rect 29942 -26826 29954 -26650
rect 29896 -26838 29954 -26826
rect 30354 -26650 30412 -26638
rect 30354 -26826 30366 -26650
rect 30400 -26826 30412 -26650
rect 30354 -26838 30412 -26826
rect 30812 -26650 30870 -26638
rect 30812 -26826 30824 -26650
rect 30858 -26826 30870 -26650
rect 30812 -26838 30870 -26826
rect 31232 -26650 31290 -26638
rect 31232 -26826 31244 -26650
rect 31278 -26826 31290 -26650
rect 31232 -26838 31290 -26826
rect 31690 -26650 31748 -26638
rect 31690 -26826 31702 -26650
rect 31736 -26826 31748 -26650
rect 31690 -26838 31748 -26826
rect 32148 -26650 32206 -26638
rect 32148 -26826 32160 -26650
rect 32194 -26826 32206 -26650
rect 32148 -26838 32206 -26826
rect 32606 -26650 32664 -26638
rect 32606 -26826 32618 -26650
rect 32652 -26826 32664 -26650
rect 32606 -26838 32664 -26826
rect 33064 -26650 33122 -26638
rect 33064 -26826 33076 -26650
rect 33110 -26826 33122 -26650
rect 33064 -26838 33122 -26826
rect 33522 -26650 33580 -26638
rect 33522 -26826 33534 -26650
rect 33568 -26826 33580 -26650
rect 33522 -26838 33580 -26826
rect 33980 -26650 34038 -26638
rect 33980 -26826 33992 -26650
rect 34026 -26826 34038 -26650
rect 33980 -26838 34038 -26826
rect 34438 -26650 34496 -26638
rect 34438 -26826 34450 -26650
rect 34484 -26826 34496 -26650
rect 34438 -26838 34496 -26826
rect 34896 -26650 34954 -26638
rect 34896 -26826 34908 -26650
rect 34942 -26826 34954 -26650
rect 34896 -26838 34954 -26826
rect 35354 -26650 35412 -26638
rect 35354 -26826 35366 -26650
rect 35400 -26826 35412 -26650
rect 35354 -26838 35412 -26826
rect 35812 -26650 35870 -26638
rect 35812 -26826 35824 -26650
rect 35858 -26826 35870 -26650
rect 35812 -26838 35870 -26826
rect 26232 -27318 26290 -27306
rect 26232 -27494 26244 -27318
rect 26278 -27494 26290 -27318
rect 26232 -27506 26290 -27494
rect 26690 -27318 26748 -27306
rect 26690 -27494 26702 -27318
rect 26736 -27494 26748 -27318
rect 26690 -27506 26748 -27494
rect 27148 -27318 27206 -27306
rect 27148 -27494 27160 -27318
rect 27194 -27494 27206 -27318
rect 27148 -27506 27206 -27494
rect 27606 -27318 27664 -27306
rect 27606 -27494 27618 -27318
rect 27652 -27494 27664 -27318
rect 27606 -27506 27664 -27494
rect 28064 -27318 28122 -27306
rect 28064 -27494 28076 -27318
rect 28110 -27494 28122 -27318
rect 28064 -27506 28122 -27494
rect 28522 -27318 28580 -27306
rect 28522 -27494 28534 -27318
rect 28568 -27494 28580 -27318
rect 28522 -27506 28580 -27494
rect 28980 -27318 29038 -27306
rect 28980 -27494 28992 -27318
rect 29026 -27494 29038 -27318
rect 28980 -27506 29038 -27494
rect 29438 -27318 29496 -27306
rect 29438 -27494 29450 -27318
rect 29484 -27494 29496 -27318
rect 29438 -27506 29496 -27494
rect 29896 -27318 29954 -27306
rect 29896 -27494 29908 -27318
rect 29942 -27494 29954 -27318
rect 29896 -27506 29954 -27494
rect 30354 -27318 30412 -27306
rect 30354 -27494 30366 -27318
rect 30400 -27494 30412 -27318
rect 30354 -27506 30412 -27494
rect 30812 -27318 30870 -27306
rect 30812 -27494 30824 -27318
rect 30858 -27494 30870 -27318
rect 30812 -27506 30870 -27494
<< pdiff >>
rect 15790 1381 15848 1393
rect 15790 -195 15802 1381
rect 15836 -195 15848 1381
rect 15790 -207 15848 -195
rect 16248 1381 16306 1393
rect 16248 -195 16260 1381
rect 16294 -195 16306 1381
rect 16248 -207 16306 -195
rect 16706 1381 16764 1393
rect 16706 -195 16718 1381
rect 16752 -195 16764 1381
rect 16706 -207 16764 -195
rect 17164 1381 17222 1393
rect 17164 -195 17176 1381
rect 17210 -195 17222 1381
rect 17164 -207 17222 -195
rect 17622 1381 17680 1393
rect 17622 -195 17634 1381
rect 17668 -195 17680 1381
rect 17622 -207 17680 -195
rect 18080 1381 18138 1393
rect 18080 -195 18092 1381
rect 18126 -195 18138 1381
rect 18080 -207 18138 -195
rect 18538 1381 18596 1393
rect 18538 -195 18550 1381
rect 18584 -195 18596 1381
rect 18538 -207 18596 -195
rect 18996 1381 19054 1393
rect 18996 -195 19008 1381
rect 19042 -195 19054 1381
rect 18996 -207 19054 -195
rect 19454 1381 19512 1393
rect 19454 -195 19466 1381
rect 19500 -195 19512 1381
rect 19454 -207 19512 -195
rect 19912 1381 19970 1393
rect 19912 -195 19924 1381
rect 19958 -195 19970 1381
rect 19912 -207 19970 -195
rect 20370 1381 20428 1393
rect 20370 -195 20382 1381
rect 20416 -195 20428 1381
rect 20370 -207 20428 -195
rect 20828 1381 20886 1393
rect 20828 -195 20840 1381
rect 20874 -195 20886 1381
rect 20828 -207 20886 -195
rect 21286 1381 21344 1393
rect 21286 -195 21298 1381
rect 21332 -195 21344 1381
rect 21286 -207 21344 -195
rect 21744 1381 21802 1393
rect 21744 -195 21756 1381
rect 21790 -195 21802 1381
rect 21744 -207 21802 -195
rect 22202 1381 22260 1393
rect 22202 -195 22214 1381
rect 22248 -195 22260 1381
rect 22202 -207 22260 -195
rect 22660 1381 22718 1393
rect 22660 -195 22672 1381
rect 22706 -195 22718 1381
rect 22660 -207 22718 -195
rect 23118 1381 23176 1393
rect 23118 -195 23130 1381
rect 23164 -195 23176 1381
rect 23118 -207 23176 -195
rect 23576 1381 23634 1393
rect 23576 -195 23588 1381
rect 23622 -195 23634 1381
rect 23576 -207 23634 -195
rect 24034 1381 24092 1393
rect 24034 -195 24046 1381
rect 24080 -195 24092 1381
rect 24034 -207 24092 -195
rect 26385 1801 26443 1813
rect 26385 625 26397 1801
rect 26431 625 26443 1801
rect 26385 613 26443 625
rect 26843 1801 26901 1813
rect 26843 625 26855 1801
rect 26889 625 26901 1801
rect 26843 613 26901 625
rect 27301 1801 27359 1813
rect 27301 625 27313 1801
rect 27347 625 27359 1801
rect 27301 613 27359 625
rect 27759 1801 27817 1813
rect 27759 625 27771 1801
rect 27805 625 27817 1801
rect 27759 613 27817 625
rect 28217 1801 28275 1813
rect 28217 625 28229 1801
rect 28263 625 28275 1801
rect 28217 613 28275 625
rect 28675 1801 28733 1813
rect 28675 625 28687 1801
rect 28721 625 28733 1801
rect 28675 613 28733 625
rect 29133 1801 29191 1813
rect 29133 625 29145 1801
rect 29179 625 29191 1801
rect 29133 613 29191 625
rect 29591 1801 29649 1813
rect 29591 625 29603 1801
rect 29637 625 29649 1801
rect 29591 613 29649 625
rect 30049 1801 30107 1813
rect 30049 625 30061 1801
rect 30095 625 30107 1801
rect 30049 613 30107 625
rect 30507 1801 30565 1813
rect 30507 625 30519 1801
rect 30553 625 30565 1801
rect 30507 613 30565 625
rect 30965 1801 31023 1813
rect 30965 625 30977 1801
rect 31011 625 31023 1801
rect 30965 613 31023 625
rect 31610 2175 31662 2193
rect 31610 2141 31618 2175
rect 31652 2141 31662 2175
rect 31610 2107 31662 2141
rect 31610 2073 31618 2107
rect 31652 2073 31662 2107
rect 31610 2039 31662 2073
rect 31610 2005 31618 2039
rect 31652 2005 31662 2039
rect 31610 1993 31662 2005
rect 31692 2175 31744 2193
rect 31692 2141 31702 2175
rect 31736 2141 31744 2175
rect 31692 2107 31744 2141
rect 31692 2073 31702 2107
rect 31736 2073 31744 2107
rect 31692 2039 31744 2073
rect 31692 2005 31702 2039
rect 31736 2005 31744 2039
rect 31692 1993 31744 2005
rect 31855 2175 31907 2193
rect 31855 2141 31863 2175
rect 31897 2141 31907 2175
rect 31855 2107 31907 2141
rect 31855 2073 31863 2107
rect 31897 2073 31907 2107
rect 31855 2039 31907 2073
rect 31855 2005 31863 2039
rect 31897 2005 31907 2039
rect 31855 1993 31907 2005
rect 31937 2175 31991 2193
rect 31937 2141 31947 2175
rect 31981 2141 31991 2175
rect 31937 2107 31991 2141
rect 31937 2073 31947 2107
rect 31981 2073 31991 2107
rect 31937 2039 31991 2073
rect 31937 2005 31947 2039
rect 31981 2005 31991 2039
rect 31937 1993 31991 2005
rect 32021 2107 32075 2193
rect 32021 2073 32031 2107
rect 32065 2073 32075 2107
rect 32021 2039 32075 2073
rect 32021 2005 32031 2039
rect 32065 2005 32075 2039
rect 32021 1993 32075 2005
rect 32105 2175 32159 2193
rect 32105 2141 32115 2175
rect 32149 2141 32159 2175
rect 32105 2107 32159 2141
rect 32105 2073 32115 2107
rect 32149 2073 32159 2107
rect 32105 2039 32159 2073
rect 32105 2005 32115 2039
rect 32149 2005 32159 2039
rect 32105 1993 32159 2005
rect 32189 2039 32241 2193
rect 32189 2005 32199 2039
rect 32233 2005 32241 2039
rect 32189 1993 32241 2005
rect 11792 -3492 11850 -3480
rect 11792 -5068 11804 -3492
rect 11838 -5068 11850 -3492
rect 11792 -5080 11850 -5068
rect 12250 -3492 12308 -3480
rect 12250 -5068 12262 -3492
rect 12296 -5068 12308 -3492
rect 12250 -5080 12308 -5068
rect 12708 -3492 12766 -3480
rect 12708 -5068 12720 -3492
rect 12754 -5068 12766 -3492
rect 12708 -5080 12766 -5068
rect 13166 -3492 13224 -3480
rect 13166 -5068 13178 -3492
rect 13212 -5068 13224 -3492
rect 13166 -5080 13224 -5068
rect 13624 -3492 13682 -3480
rect 13624 -5068 13636 -3492
rect 13670 -5068 13682 -3492
rect 13624 -5080 13682 -5068
rect 14082 -3492 14140 -3480
rect 14082 -5068 14094 -3492
rect 14128 -5068 14140 -3492
rect 14082 -5080 14140 -5068
rect 14540 -3492 14598 -3480
rect 14540 -5068 14552 -3492
rect 14586 -5068 14598 -3492
rect 14540 -5080 14598 -5068
rect 14998 -3492 15056 -3480
rect 14998 -5068 15010 -3492
rect 15044 -5068 15056 -3492
rect 14998 -5080 15056 -5068
rect 15456 -3492 15514 -3480
rect 15456 -5068 15468 -3492
rect 15502 -5068 15514 -3492
rect 15456 -5080 15514 -5068
rect 15914 -3492 15972 -3480
rect 15914 -5068 15926 -3492
rect 15960 -5068 15972 -3492
rect 15914 -5080 15972 -5068
rect 16372 -3492 16430 -3480
rect 16372 -5068 16384 -3492
rect 16418 -5068 16430 -3492
rect 16372 -5080 16430 -5068
rect 16830 -3492 16888 -3480
rect 16830 -5068 16842 -3492
rect 16876 -5068 16888 -3492
rect 16830 -5080 16888 -5068
rect 17288 -3492 17346 -3480
rect 17288 -5068 17300 -3492
rect 17334 -5068 17346 -3492
rect 17288 -5080 17346 -5068
rect 17746 -3492 17804 -3480
rect 17746 -5068 17758 -3492
rect 17792 -5068 17804 -3492
rect 17746 -5080 17804 -5068
rect 18204 -3492 18262 -3480
rect 18204 -5068 18216 -3492
rect 18250 -5068 18262 -3492
rect 18204 -5080 18262 -5068
rect 18662 -3492 18720 -3480
rect 18662 -5068 18674 -3492
rect 18708 -5068 18720 -3492
rect 18662 -5080 18720 -5068
rect 19120 -3492 19178 -3480
rect 19120 -5068 19132 -3492
rect 19166 -5068 19178 -3492
rect 19120 -5080 19178 -5068
rect 19578 -3492 19636 -3480
rect 19578 -5068 19590 -3492
rect 19624 -5068 19636 -3492
rect 19578 -5080 19636 -5068
rect 20036 -3492 20094 -3480
rect 20036 -5068 20048 -3492
rect 20082 -5068 20094 -3492
rect 20036 -5080 20094 -5068
rect 11233 -6157 11291 -6145
rect 11233 -7333 11245 -6157
rect 11279 -7333 11291 -6157
rect 11233 -7345 11291 -7333
rect 11691 -6157 11749 -6145
rect 11691 -7333 11703 -6157
rect 11737 -7333 11749 -6157
rect 11691 -7345 11749 -7333
rect 12149 -6157 12207 -6145
rect 12149 -7333 12161 -6157
rect 12195 -7333 12207 -6157
rect 12149 -7345 12207 -7333
rect 12607 -6157 12665 -6145
rect 12607 -7333 12619 -6157
rect 12653 -7333 12665 -6157
rect 12607 -7345 12665 -7333
rect 13065 -6157 13123 -6145
rect 13065 -7333 13077 -6157
rect 13111 -7333 13123 -6157
rect 13065 -7345 13123 -7333
rect 13523 -6157 13581 -6145
rect 13523 -7333 13535 -6157
rect 13569 -7333 13581 -6157
rect 13523 -7345 13581 -7333
rect 13981 -6157 14039 -6145
rect 13981 -7333 13993 -6157
rect 14027 -7333 14039 -6157
rect 13981 -7345 14039 -7333
rect 14439 -6157 14497 -6145
rect 14439 -7333 14451 -6157
rect 14485 -7333 14497 -6157
rect 14439 -7345 14497 -7333
rect 14897 -6157 14955 -6145
rect 14897 -7333 14909 -6157
rect 14943 -7333 14955 -6157
rect 14897 -7345 14955 -7333
rect 15355 -6157 15413 -6145
rect 15355 -7333 15367 -6157
rect 15401 -7333 15413 -6157
rect 15355 -7345 15413 -7333
rect 15813 -6157 15871 -6145
rect 15813 -7333 15825 -6157
rect 15859 -7333 15871 -6157
rect 15813 -7345 15871 -7333
rect 16233 -6157 16291 -6145
rect 16233 -7333 16245 -6157
rect 16279 -7333 16291 -6157
rect 16233 -7345 16291 -7333
rect 16691 -6157 16749 -6145
rect 16691 -7333 16703 -6157
rect 16737 -7333 16749 -6157
rect 16691 -7345 16749 -7333
rect 17149 -6157 17207 -6145
rect 17149 -7333 17161 -6157
rect 17195 -7333 17207 -6157
rect 17149 -7345 17207 -7333
rect 17607 -6157 17665 -6145
rect 17607 -7333 17619 -6157
rect 17653 -7333 17665 -6157
rect 17607 -7345 17665 -7333
rect 18065 -6157 18123 -6145
rect 18065 -7333 18077 -6157
rect 18111 -7333 18123 -6157
rect 18065 -7345 18123 -7333
rect 18523 -6157 18581 -6145
rect 18523 -7333 18535 -6157
rect 18569 -7333 18581 -6157
rect 18523 -7345 18581 -7333
rect 18981 -6157 19039 -6145
rect 18981 -7333 18993 -6157
rect 19027 -7333 19039 -6157
rect 18981 -7345 19039 -7333
rect 19439 -6157 19497 -6145
rect 19439 -7333 19451 -6157
rect 19485 -7333 19497 -6157
rect 19439 -7345 19497 -7333
rect 19897 -6157 19955 -6145
rect 19897 -7333 19909 -6157
rect 19943 -7333 19955 -6157
rect 19897 -7345 19955 -7333
rect 20355 -6157 20413 -6145
rect 20355 -7333 20367 -6157
rect 20401 -7333 20413 -6157
rect 20355 -7345 20413 -7333
rect 20813 -6157 20871 -6145
rect 20813 -7333 20825 -6157
rect 20859 -7333 20871 -6157
rect 20813 -7345 20871 -7333
rect 26792 -3492 26850 -3480
rect 26792 -5068 26804 -3492
rect 26838 -5068 26850 -3492
rect 26792 -5080 26850 -5068
rect 27250 -3492 27308 -3480
rect 27250 -5068 27262 -3492
rect 27296 -5068 27308 -3492
rect 27250 -5080 27308 -5068
rect 27708 -3492 27766 -3480
rect 27708 -5068 27720 -3492
rect 27754 -5068 27766 -3492
rect 27708 -5080 27766 -5068
rect 28166 -3492 28224 -3480
rect 28166 -5068 28178 -3492
rect 28212 -5068 28224 -3492
rect 28166 -5080 28224 -5068
rect 28624 -3492 28682 -3480
rect 28624 -5068 28636 -3492
rect 28670 -5068 28682 -3492
rect 28624 -5080 28682 -5068
rect 29082 -3492 29140 -3480
rect 29082 -5068 29094 -3492
rect 29128 -5068 29140 -3492
rect 29082 -5080 29140 -5068
rect 29540 -3492 29598 -3480
rect 29540 -5068 29552 -3492
rect 29586 -5068 29598 -3492
rect 29540 -5080 29598 -5068
rect 29998 -3492 30056 -3480
rect 29998 -5068 30010 -3492
rect 30044 -5068 30056 -3492
rect 29998 -5080 30056 -5068
rect 30456 -3492 30514 -3480
rect 30456 -5068 30468 -3492
rect 30502 -5068 30514 -3492
rect 30456 -5080 30514 -5068
rect 30914 -3492 30972 -3480
rect 30914 -5068 30926 -3492
rect 30960 -5068 30972 -3492
rect 30914 -5080 30972 -5068
rect 31372 -3492 31430 -3480
rect 31372 -5068 31384 -3492
rect 31418 -5068 31430 -3492
rect 31372 -5080 31430 -5068
rect 31830 -3492 31888 -3480
rect 31830 -5068 31842 -3492
rect 31876 -5068 31888 -3492
rect 31830 -5080 31888 -5068
rect 32288 -3492 32346 -3480
rect 32288 -5068 32300 -3492
rect 32334 -5068 32346 -3492
rect 32288 -5080 32346 -5068
rect 32746 -3492 32804 -3480
rect 32746 -5068 32758 -3492
rect 32792 -5068 32804 -3492
rect 32746 -5080 32804 -5068
rect 33204 -3492 33262 -3480
rect 33204 -5068 33216 -3492
rect 33250 -5068 33262 -3492
rect 33204 -5080 33262 -5068
rect 33662 -3492 33720 -3480
rect 33662 -5068 33674 -3492
rect 33708 -5068 33720 -3492
rect 33662 -5080 33720 -5068
rect 34120 -3492 34178 -3480
rect 34120 -5068 34132 -3492
rect 34166 -5068 34178 -3492
rect 34120 -5080 34178 -5068
rect 34578 -3492 34636 -3480
rect 34578 -5068 34590 -3492
rect 34624 -5068 34636 -3492
rect 34578 -5080 34636 -5068
rect 35036 -3492 35094 -3480
rect 35036 -5068 35048 -3492
rect 35082 -5068 35094 -3492
rect 35036 -5080 35094 -5068
rect 26233 -6157 26291 -6145
rect 26233 -7333 26245 -6157
rect 26279 -7333 26291 -6157
rect 26233 -7345 26291 -7333
rect 26691 -6157 26749 -6145
rect 26691 -7333 26703 -6157
rect 26737 -7333 26749 -6157
rect 26691 -7345 26749 -7333
rect 27149 -6157 27207 -6145
rect 27149 -7333 27161 -6157
rect 27195 -7333 27207 -6157
rect 27149 -7345 27207 -7333
rect 27607 -6157 27665 -6145
rect 27607 -7333 27619 -6157
rect 27653 -7333 27665 -6157
rect 27607 -7345 27665 -7333
rect 28065 -6157 28123 -6145
rect 28065 -7333 28077 -6157
rect 28111 -7333 28123 -6157
rect 28065 -7345 28123 -7333
rect 28523 -6157 28581 -6145
rect 28523 -7333 28535 -6157
rect 28569 -7333 28581 -6157
rect 28523 -7345 28581 -7333
rect 28981 -6157 29039 -6145
rect 28981 -7333 28993 -6157
rect 29027 -7333 29039 -6157
rect 28981 -7345 29039 -7333
rect 29439 -6157 29497 -6145
rect 29439 -7333 29451 -6157
rect 29485 -7333 29497 -6157
rect 29439 -7345 29497 -7333
rect 29897 -6157 29955 -6145
rect 29897 -7333 29909 -6157
rect 29943 -7333 29955 -6157
rect 29897 -7345 29955 -7333
rect 30355 -6157 30413 -6145
rect 30355 -7333 30367 -6157
rect 30401 -7333 30413 -6157
rect 30355 -7345 30413 -7333
rect 30813 -6157 30871 -6145
rect 30813 -7333 30825 -6157
rect 30859 -7333 30871 -6157
rect 30813 -7345 30871 -7333
rect 31233 -6157 31291 -6145
rect 31233 -7333 31245 -6157
rect 31279 -7333 31291 -6157
rect 31233 -7345 31291 -7333
rect 31691 -6157 31749 -6145
rect 31691 -7333 31703 -6157
rect 31737 -7333 31749 -6157
rect 31691 -7345 31749 -7333
rect 32149 -6157 32207 -6145
rect 32149 -7333 32161 -6157
rect 32195 -7333 32207 -6157
rect 32149 -7345 32207 -7333
rect 32607 -6157 32665 -6145
rect 32607 -7333 32619 -6157
rect 32653 -7333 32665 -6157
rect 32607 -7345 32665 -7333
rect 33065 -6157 33123 -6145
rect 33065 -7333 33077 -6157
rect 33111 -7333 33123 -6157
rect 33065 -7345 33123 -7333
rect 33523 -6157 33581 -6145
rect 33523 -7333 33535 -6157
rect 33569 -7333 33581 -6157
rect 33523 -7345 33581 -7333
rect 33981 -6157 34039 -6145
rect 33981 -7333 33993 -6157
rect 34027 -7333 34039 -6157
rect 33981 -7345 34039 -7333
rect 34439 -6157 34497 -6145
rect 34439 -7333 34451 -6157
rect 34485 -7333 34497 -6157
rect 34439 -7345 34497 -7333
rect 34897 -6157 34955 -6145
rect 34897 -7333 34909 -6157
rect 34943 -7333 34955 -6157
rect 34897 -7345 34955 -7333
rect 35355 -6157 35413 -6145
rect 35355 -7333 35367 -6157
rect 35401 -7333 35413 -6157
rect 35355 -7345 35413 -7333
rect 35813 -6157 35871 -6145
rect 35813 -7333 35825 -6157
rect 35859 -7333 35871 -6157
rect 35813 -7345 35871 -7333
rect 15163 -14271 15221 -14259
rect 15163 -15447 15175 -14271
rect 15209 -15447 15221 -14271
rect 15163 -15459 15221 -15447
rect 15621 -14271 15679 -14259
rect 15621 -15447 15633 -14271
rect 15667 -15447 15679 -14271
rect 15621 -15459 15679 -15447
rect 16079 -14271 16137 -14259
rect 16079 -15447 16091 -14271
rect 16125 -15447 16137 -14271
rect 16079 -15459 16137 -15447
rect 16537 -14271 16595 -14259
rect 16537 -15447 16549 -14271
rect 16583 -15447 16595 -14271
rect 16537 -15459 16595 -15447
rect 16995 -14271 17053 -14259
rect 16995 -15447 17007 -14271
rect 17041 -15447 17053 -14271
rect 16995 -15459 17053 -15447
rect 17453 -14271 17511 -14259
rect 17453 -15447 17465 -14271
rect 17499 -15447 17511 -14271
rect 17453 -15459 17511 -15447
rect 17911 -14271 17969 -14259
rect 17911 -15447 17923 -14271
rect 17957 -15447 17969 -14271
rect 17911 -15459 17969 -15447
rect 18369 -14271 18427 -14259
rect 18369 -15447 18381 -14271
rect 18415 -15447 18427 -14271
rect 18369 -15459 18427 -15447
rect 18827 -14271 18885 -14259
rect 18827 -15447 18839 -14271
rect 18873 -15447 18885 -14271
rect 18827 -15459 18885 -15447
rect 19285 -14271 19343 -14259
rect 19285 -15447 19297 -14271
rect 19331 -15447 19343 -14271
rect 19285 -15459 19343 -15447
rect 19743 -14271 19801 -14259
rect 19743 -15447 19755 -14271
rect 19789 -15447 19801 -14271
rect 19743 -15459 19801 -15447
rect 20163 -14271 20221 -14259
rect 20163 -15447 20175 -14271
rect 20209 -15447 20221 -14271
rect 20163 -15459 20221 -15447
rect 20621 -14271 20679 -14259
rect 20621 -15447 20633 -14271
rect 20667 -15447 20679 -14271
rect 20621 -15459 20679 -15447
rect 21079 -14271 21137 -14259
rect 21079 -15447 21091 -14271
rect 21125 -15447 21137 -14271
rect 21079 -15459 21137 -15447
rect 21537 -14271 21595 -14259
rect 21537 -15447 21549 -14271
rect 21583 -15447 21595 -14271
rect 21537 -15459 21595 -15447
rect 21995 -14271 22053 -14259
rect 21995 -15447 22007 -14271
rect 22041 -15447 22053 -14271
rect 21995 -15459 22053 -15447
rect 22453 -14271 22511 -14259
rect 22453 -15447 22465 -14271
rect 22499 -15447 22511 -14271
rect 22453 -15459 22511 -15447
rect 22911 -14271 22969 -14259
rect 22911 -15447 22923 -14271
rect 22957 -15447 22969 -14271
rect 22911 -15459 22969 -15447
rect 23369 -14271 23427 -14259
rect 23369 -15447 23381 -14271
rect 23415 -15447 23427 -14271
rect 23369 -15459 23427 -15447
rect 23827 -14271 23885 -14259
rect 23827 -15447 23839 -14271
rect 23873 -15447 23885 -14271
rect 23827 -15459 23885 -15447
rect 24285 -14271 24343 -14259
rect 24285 -15447 24297 -14271
rect 24331 -15447 24343 -14271
rect 24285 -15459 24343 -15447
rect 24743 -14271 24801 -14259
rect 24743 -15447 24755 -14271
rect 24789 -15447 24801 -14271
rect 24743 -15459 24801 -15447
rect 15940 -16536 15998 -16524
rect 15940 -18112 15952 -16536
rect 15986 -18112 15998 -16536
rect 15940 -18124 15998 -18112
rect 16398 -16536 16456 -16524
rect 16398 -18112 16410 -16536
rect 16444 -18112 16456 -16536
rect 16398 -18124 16456 -18112
rect 16856 -16536 16914 -16524
rect 16856 -18112 16868 -16536
rect 16902 -18112 16914 -16536
rect 16856 -18124 16914 -18112
rect 17314 -16536 17372 -16524
rect 17314 -18112 17326 -16536
rect 17360 -18112 17372 -16536
rect 17314 -18124 17372 -18112
rect 17772 -16536 17830 -16524
rect 17772 -18112 17784 -16536
rect 17818 -18112 17830 -16536
rect 17772 -18124 17830 -18112
rect 18230 -16536 18288 -16524
rect 18230 -18112 18242 -16536
rect 18276 -18112 18288 -16536
rect 18230 -18124 18288 -18112
rect 18688 -16536 18746 -16524
rect 18688 -18112 18700 -16536
rect 18734 -18112 18746 -16536
rect 18688 -18124 18746 -18112
rect 19146 -16536 19204 -16524
rect 19146 -18112 19158 -16536
rect 19192 -18112 19204 -16536
rect 19146 -18124 19204 -18112
rect 19604 -16536 19662 -16524
rect 19604 -18112 19616 -16536
rect 19650 -18112 19662 -16536
rect 19604 -18124 19662 -18112
rect 20062 -16536 20120 -16524
rect 20062 -18112 20074 -16536
rect 20108 -18112 20120 -16536
rect 20062 -18124 20120 -18112
rect 20520 -16536 20578 -16524
rect 20520 -18112 20532 -16536
rect 20566 -18112 20578 -16536
rect 20520 -18124 20578 -18112
rect 20978 -16536 21036 -16524
rect 20978 -18112 20990 -16536
rect 21024 -18112 21036 -16536
rect 20978 -18124 21036 -18112
rect 21436 -16536 21494 -16524
rect 21436 -18112 21448 -16536
rect 21482 -18112 21494 -16536
rect 21436 -18124 21494 -18112
rect 21894 -16536 21952 -16524
rect 21894 -18112 21906 -16536
rect 21940 -18112 21952 -16536
rect 21894 -18124 21952 -18112
rect 22352 -16536 22410 -16524
rect 22352 -18112 22364 -16536
rect 22398 -18112 22410 -16536
rect 22352 -18124 22410 -18112
rect 22810 -16536 22868 -16524
rect 22810 -18112 22822 -16536
rect 22856 -18112 22868 -16536
rect 22810 -18124 22868 -18112
rect 23268 -16536 23326 -16524
rect 23268 -18112 23280 -16536
rect 23314 -18112 23326 -16536
rect 23268 -18124 23326 -18112
rect 23726 -16536 23784 -16524
rect 23726 -18112 23738 -16536
rect 23772 -18112 23784 -16536
rect 23726 -18124 23784 -18112
rect 24184 -16536 24242 -16524
rect 24184 -18112 24196 -16536
rect 24230 -18112 24242 -16536
rect 24184 -18124 24242 -18112
rect 30163 -14271 30221 -14259
rect 30163 -15447 30175 -14271
rect 30209 -15447 30221 -14271
rect 30163 -15459 30221 -15447
rect 30621 -14271 30679 -14259
rect 30621 -15447 30633 -14271
rect 30667 -15447 30679 -14271
rect 30621 -15459 30679 -15447
rect 31079 -14271 31137 -14259
rect 31079 -15447 31091 -14271
rect 31125 -15447 31137 -14271
rect 31079 -15459 31137 -15447
rect 31537 -14271 31595 -14259
rect 31537 -15447 31549 -14271
rect 31583 -15447 31595 -14271
rect 31537 -15459 31595 -15447
rect 31995 -14271 32053 -14259
rect 31995 -15447 32007 -14271
rect 32041 -15447 32053 -14271
rect 31995 -15459 32053 -15447
rect 32453 -14271 32511 -14259
rect 32453 -15447 32465 -14271
rect 32499 -15447 32511 -14271
rect 32453 -15459 32511 -15447
rect 32911 -14271 32969 -14259
rect 32911 -15447 32923 -14271
rect 32957 -15447 32969 -14271
rect 32911 -15459 32969 -15447
rect 33369 -14271 33427 -14259
rect 33369 -15447 33381 -14271
rect 33415 -15447 33427 -14271
rect 33369 -15459 33427 -15447
rect 33827 -14271 33885 -14259
rect 33827 -15447 33839 -14271
rect 33873 -15447 33885 -14271
rect 33827 -15459 33885 -15447
rect 34285 -14271 34343 -14259
rect 34285 -15447 34297 -14271
rect 34331 -15447 34343 -14271
rect 34285 -15459 34343 -15447
rect 34743 -14271 34801 -14259
rect 34743 -15447 34755 -14271
rect 34789 -15447 34801 -14271
rect 34743 -15459 34801 -15447
rect 35163 -14271 35221 -14259
rect 35163 -15447 35175 -14271
rect 35209 -15447 35221 -14271
rect 35163 -15459 35221 -15447
rect 35621 -14271 35679 -14259
rect 35621 -15447 35633 -14271
rect 35667 -15447 35679 -14271
rect 35621 -15459 35679 -15447
rect 36079 -14271 36137 -14259
rect 36079 -15447 36091 -14271
rect 36125 -15447 36137 -14271
rect 36079 -15459 36137 -15447
rect 36537 -14271 36595 -14259
rect 36537 -15447 36549 -14271
rect 36583 -15447 36595 -14271
rect 36537 -15459 36595 -15447
rect 36995 -14271 37053 -14259
rect 36995 -15447 37007 -14271
rect 37041 -15447 37053 -14271
rect 36995 -15459 37053 -15447
rect 37453 -14271 37511 -14259
rect 37453 -15447 37465 -14271
rect 37499 -15447 37511 -14271
rect 37453 -15459 37511 -15447
rect 37911 -14271 37969 -14259
rect 37911 -15447 37923 -14271
rect 37957 -15447 37969 -14271
rect 37911 -15459 37969 -15447
rect 38369 -14271 38427 -14259
rect 38369 -15447 38381 -14271
rect 38415 -15447 38427 -14271
rect 38369 -15459 38427 -15447
rect 38827 -14271 38885 -14259
rect 38827 -15447 38839 -14271
rect 38873 -15447 38885 -14271
rect 38827 -15459 38885 -15447
rect 39285 -14271 39343 -14259
rect 39285 -15447 39297 -14271
rect 39331 -15447 39343 -14271
rect 39285 -15459 39343 -15447
rect 39743 -14271 39801 -14259
rect 39743 -15447 39755 -14271
rect 39789 -15447 39801 -14271
rect 39743 -15459 39801 -15447
rect 30940 -16536 30998 -16524
rect 30940 -18112 30952 -16536
rect 30986 -18112 30998 -16536
rect 30940 -18124 30998 -18112
rect 31398 -16536 31456 -16524
rect 31398 -18112 31410 -16536
rect 31444 -18112 31456 -16536
rect 31398 -18124 31456 -18112
rect 31856 -16536 31914 -16524
rect 31856 -18112 31868 -16536
rect 31902 -18112 31914 -16536
rect 31856 -18124 31914 -18112
rect 32314 -16536 32372 -16524
rect 32314 -18112 32326 -16536
rect 32360 -18112 32372 -16536
rect 32314 -18124 32372 -18112
rect 32772 -16536 32830 -16524
rect 32772 -18112 32784 -16536
rect 32818 -18112 32830 -16536
rect 32772 -18124 32830 -18112
rect 33230 -16536 33288 -16524
rect 33230 -18112 33242 -16536
rect 33276 -18112 33288 -16536
rect 33230 -18124 33288 -18112
rect 33688 -16536 33746 -16524
rect 33688 -18112 33700 -16536
rect 33734 -18112 33746 -16536
rect 33688 -18124 33746 -18112
rect 34146 -16536 34204 -16524
rect 34146 -18112 34158 -16536
rect 34192 -18112 34204 -16536
rect 34146 -18124 34204 -18112
rect 34604 -16536 34662 -16524
rect 34604 -18112 34616 -16536
rect 34650 -18112 34662 -16536
rect 34604 -18124 34662 -18112
rect 35062 -16536 35120 -16524
rect 35062 -18112 35074 -16536
rect 35108 -18112 35120 -16536
rect 35062 -18124 35120 -18112
rect 35520 -16536 35578 -16524
rect 35520 -18112 35532 -16536
rect 35566 -18112 35578 -16536
rect 35520 -18124 35578 -18112
rect 35978 -16536 36036 -16524
rect 35978 -18112 35990 -16536
rect 36024 -18112 36036 -16536
rect 35978 -18124 36036 -18112
rect 36436 -16536 36494 -16524
rect 36436 -18112 36448 -16536
rect 36482 -18112 36494 -16536
rect 36436 -18124 36494 -18112
rect 36894 -16536 36952 -16524
rect 36894 -18112 36906 -16536
rect 36940 -18112 36952 -16536
rect 36894 -18124 36952 -18112
rect 37352 -16536 37410 -16524
rect 37352 -18112 37364 -16536
rect 37398 -18112 37410 -16536
rect 37352 -18124 37410 -18112
rect 37810 -16536 37868 -16524
rect 37810 -18112 37822 -16536
rect 37856 -18112 37868 -16536
rect 37810 -18124 37868 -18112
rect 38268 -16536 38326 -16524
rect 38268 -18112 38280 -16536
rect 38314 -18112 38326 -16536
rect 38268 -18124 38326 -18112
rect 38726 -16536 38784 -16524
rect 38726 -18112 38738 -16536
rect 38772 -18112 38784 -16536
rect 38726 -18124 38784 -18112
rect 39184 -16536 39242 -16524
rect 39184 -18112 39196 -16536
rect 39230 -18112 39242 -16536
rect 39184 -18124 39242 -18112
rect 11792 -21492 11850 -21480
rect 11792 -23068 11804 -21492
rect 11838 -23068 11850 -21492
rect 11792 -23080 11850 -23068
rect 12250 -21492 12308 -21480
rect 12250 -23068 12262 -21492
rect 12296 -23068 12308 -21492
rect 12250 -23080 12308 -23068
rect 12708 -21492 12766 -21480
rect 12708 -23068 12720 -21492
rect 12754 -23068 12766 -21492
rect 12708 -23080 12766 -23068
rect 13166 -21492 13224 -21480
rect 13166 -23068 13178 -21492
rect 13212 -23068 13224 -21492
rect 13166 -23080 13224 -23068
rect 13624 -21492 13682 -21480
rect 13624 -23068 13636 -21492
rect 13670 -23068 13682 -21492
rect 13624 -23080 13682 -23068
rect 14082 -21492 14140 -21480
rect 14082 -23068 14094 -21492
rect 14128 -23068 14140 -21492
rect 14082 -23080 14140 -23068
rect 14540 -21492 14598 -21480
rect 14540 -23068 14552 -21492
rect 14586 -23068 14598 -21492
rect 14540 -23080 14598 -23068
rect 14998 -21492 15056 -21480
rect 14998 -23068 15010 -21492
rect 15044 -23068 15056 -21492
rect 14998 -23080 15056 -23068
rect 15456 -21492 15514 -21480
rect 15456 -23068 15468 -21492
rect 15502 -23068 15514 -21492
rect 15456 -23080 15514 -23068
rect 15914 -21492 15972 -21480
rect 15914 -23068 15926 -21492
rect 15960 -23068 15972 -21492
rect 15914 -23080 15972 -23068
rect 16372 -21492 16430 -21480
rect 16372 -23068 16384 -21492
rect 16418 -23068 16430 -21492
rect 16372 -23080 16430 -23068
rect 16830 -21492 16888 -21480
rect 16830 -23068 16842 -21492
rect 16876 -23068 16888 -21492
rect 16830 -23080 16888 -23068
rect 17288 -21492 17346 -21480
rect 17288 -23068 17300 -21492
rect 17334 -23068 17346 -21492
rect 17288 -23080 17346 -23068
rect 17746 -21492 17804 -21480
rect 17746 -23068 17758 -21492
rect 17792 -23068 17804 -21492
rect 17746 -23080 17804 -23068
rect 18204 -21492 18262 -21480
rect 18204 -23068 18216 -21492
rect 18250 -23068 18262 -21492
rect 18204 -23080 18262 -23068
rect 18662 -21492 18720 -21480
rect 18662 -23068 18674 -21492
rect 18708 -23068 18720 -21492
rect 18662 -23080 18720 -23068
rect 19120 -21492 19178 -21480
rect 19120 -23068 19132 -21492
rect 19166 -23068 19178 -21492
rect 19120 -23080 19178 -23068
rect 19578 -21492 19636 -21480
rect 19578 -23068 19590 -21492
rect 19624 -23068 19636 -21492
rect 19578 -23080 19636 -23068
rect 20036 -21492 20094 -21480
rect 20036 -23068 20048 -21492
rect 20082 -23068 20094 -21492
rect 20036 -23080 20094 -23068
rect 11233 -24157 11291 -24145
rect 11233 -25333 11245 -24157
rect 11279 -25333 11291 -24157
rect 11233 -25345 11291 -25333
rect 11691 -24157 11749 -24145
rect 11691 -25333 11703 -24157
rect 11737 -25333 11749 -24157
rect 11691 -25345 11749 -25333
rect 12149 -24157 12207 -24145
rect 12149 -25333 12161 -24157
rect 12195 -25333 12207 -24157
rect 12149 -25345 12207 -25333
rect 12607 -24157 12665 -24145
rect 12607 -25333 12619 -24157
rect 12653 -25333 12665 -24157
rect 12607 -25345 12665 -25333
rect 13065 -24157 13123 -24145
rect 13065 -25333 13077 -24157
rect 13111 -25333 13123 -24157
rect 13065 -25345 13123 -25333
rect 13523 -24157 13581 -24145
rect 13523 -25333 13535 -24157
rect 13569 -25333 13581 -24157
rect 13523 -25345 13581 -25333
rect 13981 -24157 14039 -24145
rect 13981 -25333 13993 -24157
rect 14027 -25333 14039 -24157
rect 13981 -25345 14039 -25333
rect 14439 -24157 14497 -24145
rect 14439 -25333 14451 -24157
rect 14485 -25333 14497 -24157
rect 14439 -25345 14497 -25333
rect 14897 -24157 14955 -24145
rect 14897 -25333 14909 -24157
rect 14943 -25333 14955 -24157
rect 14897 -25345 14955 -25333
rect 15355 -24157 15413 -24145
rect 15355 -25333 15367 -24157
rect 15401 -25333 15413 -24157
rect 15355 -25345 15413 -25333
rect 15813 -24157 15871 -24145
rect 15813 -25333 15825 -24157
rect 15859 -25333 15871 -24157
rect 15813 -25345 15871 -25333
rect 16233 -24157 16291 -24145
rect 16233 -25333 16245 -24157
rect 16279 -25333 16291 -24157
rect 16233 -25345 16291 -25333
rect 16691 -24157 16749 -24145
rect 16691 -25333 16703 -24157
rect 16737 -25333 16749 -24157
rect 16691 -25345 16749 -25333
rect 17149 -24157 17207 -24145
rect 17149 -25333 17161 -24157
rect 17195 -25333 17207 -24157
rect 17149 -25345 17207 -25333
rect 17607 -24157 17665 -24145
rect 17607 -25333 17619 -24157
rect 17653 -25333 17665 -24157
rect 17607 -25345 17665 -25333
rect 18065 -24157 18123 -24145
rect 18065 -25333 18077 -24157
rect 18111 -25333 18123 -24157
rect 18065 -25345 18123 -25333
rect 18523 -24157 18581 -24145
rect 18523 -25333 18535 -24157
rect 18569 -25333 18581 -24157
rect 18523 -25345 18581 -25333
rect 18981 -24157 19039 -24145
rect 18981 -25333 18993 -24157
rect 19027 -25333 19039 -24157
rect 18981 -25345 19039 -25333
rect 19439 -24157 19497 -24145
rect 19439 -25333 19451 -24157
rect 19485 -25333 19497 -24157
rect 19439 -25345 19497 -25333
rect 19897 -24157 19955 -24145
rect 19897 -25333 19909 -24157
rect 19943 -25333 19955 -24157
rect 19897 -25345 19955 -25333
rect 20355 -24157 20413 -24145
rect 20355 -25333 20367 -24157
rect 20401 -25333 20413 -24157
rect 20355 -25345 20413 -25333
rect 20813 -24157 20871 -24145
rect 20813 -25333 20825 -24157
rect 20859 -25333 20871 -24157
rect 20813 -25345 20871 -25333
rect 26792 -21492 26850 -21480
rect 26792 -23068 26804 -21492
rect 26838 -23068 26850 -21492
rect 26792 -23080 26850 -23068
rect 27250 -21492 27308 -21480
rect 27250 -23068 27262 -21492
rect 27296 -23068 27308 -21492
rect 27250 -23080 27308 -23068
rect 27708 -21492 27766 -21480
rect 27708 -23068 27720 -21492
rect 27754 -23068 27766 -21492
rect 27708 -23080 27766 -23068
rect 28166 -21492 28224 -21480
rect 28166 -23068 28178 -21492
rect 28212 -23068 28224 -21492
rect 28166 -23080 28224 -23068
rect 28624 -21492 28682 -21480
rect 28624 -23068 28636 -21492
rect 28670 -23068 28682 -21492
rect 28624 -23080 28682 -23068
rect 29082 -21492 29140 -21480
rect 29082 -23068 29094 -21492
rect 29128 -23068 29140 -21492
rect 29082 -23080 29140 -23068
rect 29540 -21492 29598 -21480
rect 29540 -23068 29552 -21492
rect 29586 -23068 29598 -21492
rect 29540 -23080 29598 -23068
rect 29998 -21492 30056 -21480
rect 29998 -23068 30010 -21492
rect 30044 -23068 30056 -21492
rect 29998 -23080 30056 -23068
rect 30456 -21492 30514 -21480
rect 30456 -23068 30468 -21492
rect 30502 -23068 30514 -21492
rect 30456 -23080 30514 -23068
rect 30914 -21492 30972 -21480
rect 30914 -23068 30926 -21492
rect 30960 -23068 30972 -21492
rect 30914 -23080 30972 -23068
rect 31372 -21492 31430 -21480
rect 31372 -23068 31384 -21492
rect 31418 -23068 31430 -21492
rect 31372 -23080 31430 -23068
rect 31830 -21492 31888 -21480
rect 31830 -23068 31842 -21492
rect 31876 -23068 31888 -21492
rect 31830 -23080 31888 -23068
rect 32288 -21492 32346 -21480
rect 32288 -23068 32300 -21492
rect 32334 -23068 32346 -21492
rect 32288 -23080 32346 -23068
rect 32746 -21492 32804 -21480
rect 32746 -23068 32758 -21492
rect 32792 -23068 32804 -21492
rect 32746 -23080 32804 -23068
rect 33204 -21492 33262 -21480
rect 33204 -23068 33216 -21492
rect 33250 -23068 33262 -21492
rect 33204 -23080 33262 -23068
rect 33662 -21492 33720 -21480
rect 33662 -23068 33674 -21492
rect 33708 -23068 33720 -21492
rect 33662 -23080 33720 -23068
rect 34120 -21492 34178 -21480
rect 34120 -23068 34132 -21492
rect 34166 -23068 34178 -21492
rect 34120 -23080 34178 -23068
rect 34578 -21492 34636 -21480
rect 34578 -23068 34590 -21492
rect 34624 -23068 34636 -21492
rect 34578 -23080 34636 -23068
rect 35036 -21492 35094 -21480
rect 35036 -23068 35048 -21492
rect 35082 -23068 35094 -21492
rect 35036 -23080 35094 -23068
rect 26233 -24157 26291 -24145
rect 26233 -25333 26245 -24157
rect 26279 -25333 26291 -24157
rect 26233 -25345 26291 -25333
rect 26691 -24157 26749 -24145
rect 26691 -25333 26703 -24157
rect 26737 -25333 26749 -24157
rect 26691 -25345 26749 -25333
rect 27149 -24157 27207 -24145
rect 27149 -25333 27161 -24157
rect 27195 -25333 27207 -24157
rect 27149 -25345 27207 -25333
rect 27607 -24157 27665 -24145
rect 27607 -25333 27619 -24157
rect 27653 -25333 27665 -24157
rect 27607 -25345 27665 -25333
rect 28065 -24157 28123 -24145
rect 28065 -25333 28077 -24157
rect 28111 -25333 28123 -24157
rect 28065 -25345 28123 -25333
rect 28523 -24157 28581 -24145
rect 28523 -25333 28535 -24157
rect 28569 -25333 28581 -24157
rect 28523 -25345 28581 -25333
rect 28981 -24157 29039 -24145
rect 28981 -25333 28993 -24157
rect 29027 -25333 29039 -24157
rect 28981 -25345 29039 -25333
rect 29439 -24157 29497 -24145
rect 29439 -25333 29451 -24157
rect 29485 -25333 29497 -24157
rect 29439 -25345 29497 -25333
rect 29897 -24157 29955 -24145
rect 29897 -25333 29909 -24157
rect 29943 -25333 29955 -24157
rect 29897 -25345 29955 -25333
rect 30355 -24157 30413 -24145
rect 30355 -25333 30367 -24157
rect 30401 -25333 30413 -24157
rect 30355 -25345 30413 -25333
rect 30813 -24157 30871 -24145
rect 30813 -25333 30825 -24157
rect 30859 -25333 30871 -24157
rect 30813 -25345 30871 -25333
rect 31233 -24157 31291 -24145
rect 31233 -25333 31245 -24157
rect 31279 -25333 31291 -24157
rect 31233 -25345 31291 -25333
rect 31691 -24157 31749 -24145
rect 31691 -25333 31703 -24157
rect 31737 -25333 31749 -24157
rect 31691 -25345 31749 -25333
rect 32149 -24157 32207 -24145
rect 32149 -25333 32161 -24157
rect 32195 -25333 32207 -24157
rect 32149 -25345 32207 -25333
rect 32607 -24157 32665 -24145
rect 32607 -25333 32619 -24157
rect 32653 -25333 32665 -24157
rect 32607 -25345 32665 -25333
rect 33065 -24157 33123 -24145
rect 33065 -25333 33077 -24157
rect 33111 -25333 33123 -24157
rect 33065 -25345 33123 -25333
rect 33523 -24157 33581 -24145
rect 33523 -25333 33535 -24157
rect 33569 -25333 33581 -24157
rect 33523 -25345 33581 -25333
rect 33981 -24157 34039 -24145
rect 33981 -25333 33993 -24157
rect 34027 -25333 34039 -24157
rect 33981 -25345 34039 -25333
rect 34439 -24157 34497 -24145
rect 34439 -25333 34451 -24157
rect 34485 -25333 34497 -24157
rect 34439 -25345 34497 -25333
rect 34897 -24157 34955 -24145
rect 34897 -25333 34909 -24157
rect 34943 -25333 34955 -24157
rect 34897 -25345 34955 -25333
rect 35355 -24157 35413 -24145
rect 35355 -25333 35367 -24157
rect 35401 -25333 35413 -24157
rect 35355 -25345 35413 -25333
rect 35813 -24157 35871 -24145
rect 35813 -25333 35825 -24157
rect 35859 -25333 35871 -24157
rect 35813 -25345 35871 -25333
<< ndiffc >>
rect 17634 3056 17668 3232
rect 18092 3056 18126 3232
rect 18550 3056 18584 3232
rect 19008 3056 19042 3232
rect 19466 3056 19500 3232
rect 19924 3056 19958 3232
rect 20382 3056 20416 3232
rect 20840 3056 20874 3232
rect 21298 3056 21332 3232
rect 21756 3056 21790 3232
rect 22214 3056 22248 3232
rect 26396 3056 26430 3232
rect 26854 3056 26888 3232
rect 27312 3056 27346 3232
rect 27770 3056 27804 3232
rect 28228 3056 28262 3232
rect 28686 3056 28720 3232
rect 29144 3056 29178 3232
rect 29602 3056 29636 3232
rect 30060 3056 30094 3232
rect 30518 3056 30552 3232
rect 30976 3056 31010 3232
rect 31618 2393 31652 2427
rect 31618 2325 31652 2359
rect 31702 2393 31736 2427
rect 31702 2325 31736 2359
rect 31863 2397 31897 2431
rect 31947 2389 31981 2423
rect 32031 2397 32065 2431
rect 32115 2389 32149 2423
rect 32199 2396 32233 2430
rect 11244 -8826 11278 -8650
rect 11702 -8826 11736 -8650
rect 12160 -8826 12194 -8650
rect 12618 -8826 12652 -8650
rect 13076 -8826 13110 -8650
rect 13534 -8826 13568 -8650
rect 13992 -8826 14026 -8650
rect 14450 -8826 14484 -8650
rect 14908 -8826 14942 -8650
rect 15366 -8826 15400 -8650
rect 15824 -8826 15858 -8650
rect 16244 -8826 16278 -8650
rect 16702 -8826 16736 -8650
rect 17160 -8826 17194 -8650
rect 17618 -8826 17652 -8650
rect 18076 -8826 18110 -8650
rect 18534 -8826 18568 -8650
rect 18992 -8826 19026 -8650
rect 19450 -8826 19484 -8650
rect 19908 -8826 19942 -8650
rect 20366 -8826 20400 -8650
rect 20824 -8826 20858 -8650
rect 11244 -9494 11278 -9318
rect 11702 -9494 11736 -9318
rect 12160 -9494 12194 -9318
rect 12618 -9494 12652 -9318
rect 13076 -9494 13110 -9318
rect 13534 -9494 13568 -9318
rect 13992 -9494 14026 -9318
rect 14450 -9494 14484 -9318
rect 14908 -9494 14942 -9318
rect 15366 -9494 15400 -9318
rect 15824 -9494 15858 -9318
rect 26244 -8826 26278 -8650
rect 26702 -8826 26736 -8650
rect 27160 -8826 27194 -8650
rect 27618 -8826 27652 -8650
rect 28076 -8826 28110 -8650
rect 28534 -8826 28568 -8650
rect 28992 -8826 29026 -8650
rect 29450 -8826 29484 -8650
rect 29908 -8826 29942 -8650
rect 30366 -8826 30400 -8650
rect 30824 -8826 30858 -8650
rect 31244 -8826 31278 -8650
rect 31702 -8826 31736 -8650
rect 32160 -8826 32194 -8650
rect 32618 -8826 32652 -8650
rect 33076 -8826 33110 -8650
rect 33534 -8826 33568 -8650
rect 33992 -8826 34026 -8650
rect 34450 -8826 34484 -8650
rect 34908 -8826 34942 -8650
rect 35366 -8826 35400 -8650
rect 35824 -8826 35858 -8650
rect 26244 -9494 26278 -9318
rect 26702 -9494 26736 -9318
rect 27160 -9494 27194 -9318
rect 27618 -9494 27652 -9318
rect 28076 -9494 28110 -9318
rect 28534 -9494 28568 -9318
rect 28992 -9494 29026 -9318
rect 29450 -9494 29484 -9318
rect 29908 -9494 29942 -9318
rect 30366 -9494 30400 -9318
rect 30824 -9494 30858 -9318
rect 20176 -12286 20210 -12110
rect 20634 -12286 20668 -12110
rect 21092 -12286 21126 -12110
rect 21550 -12286 21584 -12110
rect 22008 -12286 22042 -12110
rect 22466 -12286 22500 -12110
rect 22924 -12286 22958 -12110
rect 23382 -12286 23416 -12110
rect 23840 -12286 23874 -12110
rect 24298 -12286 24332 -12110
rect 24756 -12286 24790 -12110
rect 15176 -12954 15210 -12778
rect 15634 -12954 15668 -12778
rect 16092 -12954 16126 -12778
rect 16550 -12954 16584 -12778
rect 17008 -12954 17042 -12778
rect 17466 -12954 17500 -12778
rect 17924 -12954 17958 -12778
rect 18382 -12954 18416 -12778
rect 18840 -12954 18874 -12778
rect 19298 -12954 19332 -12778
rect 19756 -12954 19790 -12778
rect 20176 -12954 20210 -12778
rect 20634 -12954 20668 -12778
rect 21092 -12954 21126 -12778
rect 21550 -12954 21584 -12778
rect 22008 -12954 22042 -12778
rect 22466 -12954 22500 -12778
rect 22924 -12954 22958 -12778
rect 23382 -12954 23416 -12778
rect 23840 -12954 23874 -12778
rect 24298 -12954 24332 -12778
rect 24756 -12954 24790 -12778
rect 35176 -12286 35210 -12110
rect 35634 -12286 35668 -12110
rect 36092 -12286 36126 -12110
rect 36550 -12286 36584 -12110
rect 37008 -12286 37042 -12110
rect 37466 -12286 37500 -12110
rect 37924 -12286 37958 -12110
rect 38382 -12286 38416 -12110
rect 38840 -12286 38874 -12110
rect 39298 -12286 39332 -12110
rect 39756 -12286 39790 -12110
rect 30176 -12954 30210 -12778
rect 30634 -12954 30668 -12778
rect 31092 -12954 31126 -12778
rect 31550 -12954 31584 -12778
rect 32008 -12954 32042 -12778
rect 32466 -12954 32500 -12778
rect 32924 -12954 32958 -12778
rect 33382 -12954 33416 -12778
rect 33840 -12954 33874 -12778
rect 34298 -12954 34332 -12778
rect 34756 -12954 34790 -12778
rect 35176 -12954 35210 -12778
rect 35634 -12954 35668 -12778
rect 36092 -12954 36126 -12778
rect 36550 -12954 36584 -12778
rect 37008 -12954 37042 -12778
rect 37466 -12954 37500 -12778
rect 37924 -12954 37958 -12778
rect 38382 -12954 38416 -12778
rect 38840 -12954 38874 -12778
rect 39298 -12954 39332 -12778
rect 39756 -12954 39790 -12778
rect 11244 -26826 11278 -26650
rect 11702 -26826 11736 -26650
rect 12160 -26826 12194 -26650
rect 12618 -26826 12652 -26650
rect 13076 -26826 13110 -26650
rect 13534 -26826 13568 -26650
rect 13992 -26826 14026 -26650
rect 14450 -26826 14484 -26650
rect 14908 -26826 14942 -26650
rect 15366 -26826 15400 -26650
rect 15824 -26826 15858 -26650
rect 16244 -26826 16278 -26650
rect 16702 -26826 16736 -26650
rect 17160 -26826 17194 -26650
rect 17618 -26826 17652 -26650
rect 18076 -26826 18110 -26650
rect 18534 -26826 18568 -26650
rect 18992 -26826 19026 -26650
rect 19450 -26826 19484 -26650
rect 19908 -26826 19942 -26650
rect 20366 -26826 20400 -26650
rect 20824 -26826 20858 -26650
rect 11244 -27494 11278 -27318
rect 11702 -27494 11736 -27318
rect 12160 -27494 12194 -27318
rect 12618 -27494 12652 -27318
rect 13076 -27494 13110 -27318
rect 13534 -27494 13568 -27318
rect 13992 -27494 14026 -27318
rect 14450 -27494 14484 -27318
rect 14908 -27494 14942 -27318
rect 15366 -27494 15400 -27318
rect 15824 -27494 15858 -27318
rect 26244 -26826 26278 -26650
rect 26702 -26826 26736 -26650
rect 27160 -26826 27194 -26650
rect 27618 -26826 27652 -26650
rect 28076 -26826 28110 -26650
rect 28534 -26826 28568 -26650
rect 28992 -26826 29026 -26650
rect 29450 -26826 29484 -26650
rect 29908 -26826 29942 -26650
rect 30366 -26826 30400 -26650
rect 30824 -26826 30858 -26650
rect 31244 -26826 31278 -26650
rect 31702 -26826 31736 -26650
rect 32160 -26826 32194 -26650
rect 32618 -26826 32652 -26650
rect 33076 -26826 33110 -26650
rect 33534 -26826 33568 -26650
rect 33992 -26826 34026 -26650
rect 34450 -26826 34484 -26650
rect 34908 -26826 34942 -26650
rect 35366 -26826 35400 -26650
rect 35824 -26826 35858 -26650
rect 26244 -27494 26278 -27318
rect 26702 -27494 26736 -27318
rect 27160 -27494 27194 -27318
rect 27618 -27494 27652 -27318
rect 28076 -27494 28110 -27318
rect 28534 -27494 28568 -27318
rect 28992 -27494 29026 -27318
rect 29450 -27494 29484 -27318
rect 29908 -27494 29942 -27318
rect 30366 -27494 30400 -27318
rect 30824 -27494 30858 -27318
<< pdiffc >>
rect 15802 -195 15836 1381
rect 16260 -195 16294 1381
rect 16718 -195 16752 1381
rect 17176 -195 17210 1381
rect 17634 -195 17668 1381
rect 18092 -195 18126 1381
rect 18550 -195 18584 1381
rect 19008 -195 19042 1381
rect 19466 -195 19500 1381
rect 19924 -195 19958 1381
rect 20382 -195 20416 1381
rect 20840 -195 20874 1381
rect 21298 -195 21332 1381
rect 21756 -195 21790 1381
rect 22214 -195 22248 1381
rect 22672 -195 22706 1381
rect 23130 -195 23164 1381
rect 23588 -195 23622 1381
rect 24046 -195 24080 1381
rect 26397 625 26431 1801
rect 26855 625 26889 1801
rect 27313 625 27347 1801
rect 27771 625 27805 1801
rect 28229 625 28263 1801
rect 28687 625 28721 1801
rect 29145 625 29179 1801
rect 29603 625 29637 1801
rect 30061 625 30095 1801
rect 30519 625 30553 1801
rect 30977 625 31011 1801
rect 31618 2141 31652 2175
rect 31618 2073 31652 2107
rect 31618 2005 31652 2039
rect 31702 2141 31736 2175
rect 31702 2073 31736 2107
rect 31702 2005 31736 2039
rect 31863 2141 31897 2175
rect 31863 2073 31897 2107
rect 31863 2005 31897 2039
rect 31947 2141 31981 2175
rect 31947 2073 31981 2107
rect 31947 2005 31981 2039
rect 32031 2073 32065 2107
rect 32031 2005 32065 2039
rect 32115 2141 32149 2175
rect 32115 2073 32149 2107
rect 32115 2005 32149 2039
rect 32199 2005 32233 2039
rect 11804 -5068 11838 -3492
rect 12262 -5068 12296 -3492
rect 12720 -5068 12754 -3492
rect 13178 -5068 13212 -3492
rect 13636 -5068 13670 -3492
rect 14094 -5068 14128 -3492
rect 14552 -5068 14586 -3492
rect 15010 -5068 15044 -3492
rect 15468 -5068 15502 -3492
rect 15926 -5068 15960 -3492
rect 16384 -5068 16418 -3492
rect 16842 -5068 16876 -3492
rect 17300 -5068 17334 -3492
rect 17758 -5068 17792 -3492
rect 18216 -5068 18250 -3492
rect 18674 -5068 18708 -3492
rect 19132 -5068 19166 -3492
rect 19590 -5068 19624 -3492
rect 20048 -5068 20082 -3492
rect 11245 -7333 11279 -6157
rect 11703 -7333 11737 -6157
rect 12161 -7333 12195 -6157
rect 12619 -7333 12653 -6157
rect 13077 -7333 13111 -6157
rect 13535 -7333 13569 -6157
rect 13993 -7333 14027 -6157
rect 14451 -7333 14485 -6157
rect 14909 -7333 14943 -6157
rect 15367 -7333 15401 -6157
rect 15825 -7333 15859 -6157
rect 16245 -7333 16279 -6157
rect 16703 -7333 16737 -6157
rect 17161 -7333 17195 -6157
rect 17619 -7333 17653 -6157
rect 18077 -7333 18111 -6157
rect 18535 -7333 18569 -6157
rect 18993 -7333 19027 -6157
rect 19451 -7333 19485 -6157
rect 19909 -7333 19943 -6157
rect 20367 -7333 20401 -6157
rect 20825 -7333 20859 -6157
rect 26804 -5068 26838 -3492
rect 27262 -5068 27296 -3492
rect 27720 -5068 27754 -3492
rect 28178 -5068 28212 -3492
rect 28636 -5068 28670 -3492
rect 29094 -5068 29128 -3492
rect 29552 -5068 29586 -3492
rect 30010 -5068 30044 -3492
rect 30468 -5068 30502 -3492
rect 30926 -5068 30960 -3492
rect 31384 -5068 31418 -3492
rect 31842 -5068 31876 -3492
rect 32300 -5068 32334 -3492
rect 32758 -5068 32792 -3492
rect 33216 -5068 33250 -3492
rect 33674 -5068 33708 -3492
rect 34132 -5068 34166 -3492
rect 34590 -5068 34624 -3492
rect 35048 -5068 35082 -3492
rect 26245 -7333 26279 -6157
rect 26703 -7333 26737 -6157
rect 27161 -7333 27195 -6157
rect 27619 -7333 27653 -6157
rect 28077 -7333 28111 -6157
rect 28535 -7333 28569 -6157
rect 28993 -7333 29027 -6157
rect 29451 -7333 29485 -6157
rect 29909 -7333 29943 -6157
rect 30367 -7333 30401 -6157
rect 30825 -7333 30859 -6157
rect 31245 -7333 31279 -6157
rect 31703 -7333 31737 -6157
rect 32161 -7333 32195 -6157
rect 32619 -7333 32653 -6157
rect 33077 -7333 33111 -6157
rect 33535 -7333 33569 -6157
rect 33993 -7333 34027 -6157
rect 34451 -7333 34485 -6157
rect 34909 -7333 34943 -6157
rect 35367 -7333 35401 -6157
rect 35825 -7333 35859 -6157
rect 15175 -15447 15209 -14271
rect 15633 -15447 15667 -14271
rect 16091 -15447 16125 -14271
rect 16549 -15447 16583 -14271
rect 17007 -15447 17041 -14271
rect 17465 -15447 17499 -14271
rect 17923 -15447 17957 -14271
rect 18381 -15447 18415 -14271
rect 18839 -15447 18873 -14271
rect 19297 -15447 19331 -14271
rect 19755 -15447 19789 -14271
rect 20175 -15447 20209 -14271
rect 20633 -15447 20667 -14271
rect 21091 -15447 21125 -14271
rect 21549 -15447 21583 -14271
rect 22007 -15447 22041 -14271
rect 22465 -15447 22499 -14271
rect 22923 -15447 22957 -14271
rect 23381 -15447 23415 -14271
rect 23839 -15447 23873 -14271
rect 24297 -15447 24331 -14271
rect 24755 -15447 24789 -14271
rect 15952 -18112 15986 -16536
rect 16410 -18112 16444 -16536
rect 16868 -18112 16902 -16536
rect 17326 -18112 17360 -16536
rect 17784 -18112 17818 -16536
rect 18242 -18112 18276 -16536
rect 18700 -18112 18734 -16536
rect 19158 -18112 19192 -16536
rect 19616 -18112 19650 -16536
rect 20074 -18112 20108 -16536
rect 20532 -18112 20566 -16536
rect 20990 -18112 21024 -16536
rect 21448 -18112 21482 -16536
rect 21906 -18112 21940 -16536
rect 22364 -18112 22398 -16536
rect 22822 -18112 22856 -16536
rect 23280 -18112 23314 -16536
rect 23738 -18112 23772 -16536
rect 24196 -18112 24230 -16536
rect 30175 -15447 30209 -14271
rect 30633 -15447 30667 -14271
rect 31091 -15447 31125 -14271
rect 31549 -15447 31583 -14271
rect 32007 -15447 32041 -14271
rect 32465 -15447 32499 -14271
rect 32923 -15447 32957 -14271
rect 33381 -15447 33415 -14271
rect 33839 -15447 33873 -14271
rect 34297 -15447 34331 -14271
rect 34755 -15447 34789 -14271
rect 35175 -15447 35209 -14271
rect 35633 -15447 35667 -14271
rect 36091 -15447 36125 -14271
rect 36549 -15447 36583 -14271
rect 37007 -15447 37041 -14271
rect 37465 -15447 37499 -14271
rect 37923 -15447 37957 -14271
rect 38381 -15447 38415 -14271
rect 38839 -15447 38873 -14271
rect 39297 -15447 39331 -14271
rect 39755 -15447 39789 -14271
rect 30952 -18112 30986 -16536
rect 31410 -18112 31444 -16536
rect 31868 -18112 31902 -16536
rect 32326 -18112 32360 -16536
rect 32784 -18112 32818 -16536
rect 33242 -18112 33276 -16536
rect 33700 -18112 33734 -16536
rect 34158 -18112 34192 -16536
rect 34616 -18112 34650 -16536
rect 35074 -18112 35108 -16536
rect 35532 -18112 35566 -16536
rect 35990 -18112 36024 -16536
rect 36448 -18112 36482 -16536
rect 36906 -18112 36940 -16536
rect 37364 -18112 37398 -16536
rect 37822 -18112 37856 -16536
rect 38280 -18112 38314 -16536
rect 38738 -18112 38772 -16536
rect 39196 -18112 39230 -16536
rect 11804 -23068 11838 -21492
rect 12262 -23068 12296 -21492
rect 12720 -23068 12754 -21492
rect 13178 -23068 13212 -21492
rect 13636 -23068 13670 -21492
rect 14094 -23068 14128 -21492
rect 14552 -23068 14586 -21492
rect 15010 -23068 15044 -21492
rect 15468 -23068 15502 -21492
rect 15926 -23068 15960 -21492
rect 16384 -23068 16418 -21492
rect 16842 -23068 16876 -21492
rect 17300 -23068 17334 -21492
rect 17758 -23068 17792 -21492
rect 18216 -23068 18250 -21492
rect 18674 -23068 18708 -21492
rect 19132 -23068 19166 -21492
rect 19590 -23068 19624 -21492
rect 20048 -23068 20082 -21492
rect 11245 -25333 11279 -24157
rect 11703 -25333 11737 -24157
rect 12161 -25333 12195 -24157
rect 12619 -25333 12653 -24157
rect 13077 -25333 13111 -24157
rect 13535 -25333 13569 -24157
rect 13993 -25333 14027 -24157
rect 14451 -25333 14485 -24157
rect 14909 -25333 14943 -24157
rect 15367 -25333 15401 -24157
rect 15825 -25333 15859 -24157
rect 16245 -25333 16279 -24157
rect 16703 -25333 16737 -24157
rect 17161 -25333 17195 -24157
rect 17619 -25333 17653 -24157
rect 18077 -25333 18111 -24157
rect 18535 -25333 18569 -24157
rect 18993 -25333 19027 -24157
rect 19451 -25333 19485 -24157
rect 19909 -25333 19943 -24157
rect 20367 -25333 20401 -24157
rect 20825 -25333 20859 -24157
rect 26804 -23068 26838 -21492
rect 27262 -23068 27296 -21492
rect 27720 -23068 27754 -21492
rect 28178 -23068 28212 -21492
rect 28636 -23068 28670 -21492
rect 29094 -23068 29128 -21492
rect 29552 -23068 29586 -21492
rect 30010 -23068 30044 -21492
rect 30468 -23068 30502 -21492
rect 30926 -23068 30960 -21492
rect 31384 -23068 31418 -21492
rect 31842 -23068 31876 -21492
rect 32300 -23068 32334 -21492
rect 32758 -23068 32792 -21492
rect 33216 -23068 33250 -21492
rect 33674 -23068 33708 -21492
rect 34132 -23068 34166 -21492
rect 34590 -23068 34624 -21492
rect 35048 -23068 35082 -21492
rect 26245 -25333 26279 -24157
rect 26703 -25333 26737 -24157
rect 27161 -25333 27195 -24157
rect 27619 -25333 27653 -24157
rect 28077 -25333 28111 -24157
rect 28535 -25333 28569 -24157
rect 28993 -25333 29027 -24157
rect 29451 -25333 29485 -24157
rect 29909 -25333 29943 -24157
rect 30367 -25333 30401 -24157
rect 30825 -25333 30859 -24157
rect 31245 -25333 31279 -24157
rect 31703 -25333 31737 -24157
rect 32161 -25333 32195 -24157
rect 32619 -25333 32653 -24157
rect 33077 -25333 33111 -24157
rect 33535 -25333 33569 -24157
rect 33993 -25333 34027 -24157
rect 34451 -25333 34485 -24157
rect 34909 -25333 34943 -24157
rect 35367 -25333 35401 -24157
rect 35825 -25333 35859 -24157
<< psubdiff >>
rect 15426 4210 15588 4310
rect 24288 4210 24450 4310
rect 15426 4148 15526 4210
rect 24350 4148 24450 4210
rect 15426 2610 15526 2672
rect 24350 2610 24450 2672
rect 15426 2510 15588 2610
rect 24288 2510 24450 2610
rect 26008 4210 26170 4310
rect 31290 4210 31452 4310
rect 26008 4148 26108 4210
rect 31352 4148 31452 4210
rect 26008 2530 26108 2592
rect 31352 2530 31452 2592
rect 26008 2430 26170 2530
rect 31290 2430 31452 2530
rect 10818 -8208 10980 -8108
rect 21100 -8208 21262 -8108
rect 10818 -8270 10918 -8208
rect 21162 -8270 21262 -8208
rect 10818 -10472 10918 -10410
rect 21162 -10472 21262 -10410
rect 10818 -10572 10980 -10472
rect 21100 -10572 21262 -10472
rect 25818 -8208 25980 -8108
rect 36100 -8208 36262 -8108
rect 25818 -8270 25918 -8208
rect 36162 -8270 36262 -8208
rect 25818 -10472 25918 -10410
rect 36162 -10472 36262 -10410
rect 25818 -10572 25980 -10472
rect 36100 -10572 36262 -10472
rect 14772 -11132 14934 -11032
rect 25054 -11132 25216 -11032
rect 14772 -11194 14872 -11132
rect 25116 -11194 25216 -11132
rect 14772 -13396 14872 -13334
rect 25116 -13396 25216 -13334
rect 14772 -13496 14934 -13396
rect 25054 -13496 25216 -13396
rect 29772 -11132 29934 -11032
rect 40054 -11132 40216 -11032
rect 29772 -11194 29872 -11132
rect 40116 -11194 40216 -11132
rect 29772 -13396 29872 -13334
rect 40116 -13396 40216 -13334
rect 29772 -13496 29934 -13396
rect 40054 -13496 40216 -13396
rect 10818 -26208 10980 -26108
rect 21100 -26208 21262 -26108
rect 10818 -26270 10918 -26208
rect 21162 -26270 21262 -26208
rect 10818 -28472 10918 -28410
rect 21162 -28472 21262 -28410
rect 10818 -28572 10980 -28472
rect 21100 -28572 21262 -28472
rect 25818 -26208 25980 -26108
rect 36100 -26208 36262 -26108
rect 25818 -26270 25918 -26208
rect 36162 -26270 36262 -26208
rect 25818 -28472 25918 -28410
rect 36162 -28472 36262 -28410
rect 25818 -28572 25980 -28472
rect 36100 -28572 36262 -28472
<< nsubdiff >>
rect 15426 2174 15588 2274
rect 24288 2174 24450 2274
rect 15426 2112 15526 2174
rect 24350 2112 24450 2174
rect 15426 -1558 15526 -1496
rect 24350 -1558 24450 -1496
rect 15426 -1658 15588 -1558
rect 24288 -1658 24450 -1558
rect 26008 2094 26170 2194
rect 31290 2094 31452 2194
rect 26008 2032 26108 2094
rect 31352 2032 31452 2094
rect 26008 -1558 26108 -1496
rect 31352 -1558 31452 -1496
rect 26008 -1658 26170 -1558
rect 31290 -1658 31452 -1558
rect 10818 -2128 10980 -2028
rect 21100 -2128 21262 -2028
rect 10818 -2190 10918 -2128
rect 21162 -2190 21262 -2128
rect 10818 -7772 10918 -7710
rect 21162 -7772 21262 -7710
rect 10818 -7872 10980 -7772
rect 21100 -7872 21262 -7772
rect 25818 -2128 25980 -2028
rect 36100 -2128 36262 -2028
rect 25818 -2190 25918 -2128
rect 36162 -2190 36262 -2128
rect 25818 -7772 25918 -7710
rect 36162 -7772 36262 -7710
rect 25818 -7872 25980 -7772
rect 36100 -7872 36262 -7772
rect 14772 -13832 14934 -13732
rect 25054 -13832 25216 -13732
rect 14772 -13894 14872 -13832
rect 25116 -13894 25216 -13832
rect 14772 -19476 14872 -19414
rect 25116 -19476 25216 -19414
rect 14772 -19576 14934 -19476
rect 25054 -19576 25216 -19476
rect 29772 -13832 29934 -13732
rect 40054 -13832 40216 -13732
rect 29772 -13894 29872 -13832
rect 40116 -13894 40216 -13832
rect 29772 -19476 29872 -19414
rect 40116 -19476 40216 -19414
rect 29772 -19576 29934 -19476
rect 40054 -19576 40216 -19476
rect 10818 -20128 10980 -20028
rect 21100 -20128 21262 -20028
rect 10818 -20190 10918 -20128
rect 21162 -20190 21262 -20128
rect 10818 -25772 10918 -25710
rect 21162 -25772 21262 -25710
rect 10818 -25872 10980 -25772
rect 21100 -25872 21262 -25772
rect 25818 -20128 25980 -20028
rect 36100 -20128 36262 -20028
rect 25818 -20190 25918 -20128
rect 36162 -20190 36262 -20128
rect 25818 -25772 25918 -25710
rect 36162 -25772 36262 -25710
rect 25818 -25872 25980 -25772
rect 36100 -25872 36262 -25772
<< psubdiffcont >>
rect 15588 4210 24288 4310
rect 15426 2672 15526 4148
rect 24350 2672 24450 4148
rect 15588 2510 24288 2610
rect 26170 4210 31290 4310
rect 26008 2592 26108 4148
rect 31352 2592 31452 4148
rect 26170 2430 31290 2530
rect 10980 -8208 21100 -8108
rect 10818 -10410 10918 -8270
rect 21162 -10410 21262 -8270
rect 10980 -10572 21100 -10472
rect 25980 -8208 36100 -8108
rect 25818 -10410 25918 -8270
rect 36162 -10410 36262 -8270
rect 25980 -10572 36100 -10472
rect 14934 -11132 25054 -11032
rect 14772 -13334 14872 -11194
rect 25116 -13334 25216 -11194
rect 14934 -13496 25054 -13396
rect 29934 -11132 40054 -11032
rect 29772 -13334 29872 -11194
rect 40116 -13334 40216 -11194
rect 29934 -13496 40054 -13396
rect 10980 -26208 21100 -26108
rect 10818 -28410 10918 -26270
rect 21162 -28410 21262 -26270
rect 10980 -28572 21100 -28472
rect 25980 -26208 36100 -26108
rect 25818 -28410 25918 -26270
rect 36162 -28410 36262 -26270
rect 25980 -28572 36100 -28472
<< nsubdiffcont >>
rect 15588 2174 24288 2274
rect 15426 -1496 15526 2112
rect 24350 -1496 24450 2112
rect 15588 -1658 24288 -1558
rect 26170 2094 31290 2194
rect 26008 -1496 26108 2032
rect 31352 -1496 31452 2032
rect 26170 -1658 31290 -1558
rect 10980 -2128 21100 -2028
rect 10818 -7710 10918 -2190
rect 21162 -7710 21262 -2190
rect 10980 -7872 21100 -7772
rect 25980 -2128 36100 -2028
rect 25818 -7710 25918 -2190
rect 36162 -7710 36262 -2190
rect 25980 -7872 36100 -7772
rect 14934 -13832 25054 -13732
rect 14772 -19414 14872 -13894
rect 25116 -19414 25216 -13894
rect 14934 -19576 25054 -19476
rect 29934 -13832 40054 -13732
rect 29772 -19414 29872 -13894
rect 40116 -19414 40216 -13894
rect 29934 -19576 40054 -19476
rect 10980 -20128 21100 -20028
rect 10818 -25710 10918 -20190
rect 21162 -25710 21262 -20190
rect 10980 -25872 21100 -25772
rect 25980 -20128 36100 -20028
rect 25818 -25710 25918 -20190
rect 36162 -25710 36262 -20190
rect 25980 -25872 36100 -25772
<< poly >>
rect 17754 3316 18006 3332
rect 17754 3299 17770 3316
rect 17680 3282 17770 3299
rect 17990 3299 18006 3316
rect 18212 3316 18464 3332
rect 18212 3299 18228 3316
rect 17990 3282 18080 3299
rect 17680 3244 18080 3282
rect 18138 3282 18228 3299
rect 18448 3299 18464 3316
rect 18670 3316 18922 3332
rect 18670 3299 18686 3316
rect 18448 3282 18538 3299
rect 18138 3244 18538 3282
rect 18596 3282 18686 3299
rect 18906 3299 18922 3316
rect 19128 3316 19380 3332
rect 19128 3299 19144 3316
rect 18906 3282 18996 3299
rect 18596 3244 18996 3282
rect 19054 3282 19144 3299
rect 19364 3299 19380 3316
rect 19586 3316 19838 3332
rect 19586 3299 19602 3316
rect 19364 3282 19454 3299
rect 19054 3244 19454 3282
rect 19512 3282 19602 3299
rect 19822 3299 19838 3316
rect 20044 3316 20296 3332
rect 20044 3299 20060 3316
rect 19822 3282 19912 3299
rect 19512 3244 19912 3282
rect 19970 3282 20060 3299
rect 20280 3299 20296 3316
rect 20502 3316 20754 3332
rect 20502 3299 20518 3316
rect 20280 3282 20370 3299
rect 19970 3244 20370 3282
rect 20428 3282 20518 3299
rect 20738 3299 20754 3316
rect 20960 3316 21212 3332
rect 20960 3299 20976 3316
rect 20738 3282 20828 3299
rect 20428 3244 20828 3282
rect 20886 3282 20976 3299
rect 21196 3299 21212 3316
rect 21418 3316 21670 3332
rect 21418 3299 21434 3316
rect 21196 3282 21286 3299
rect 20886 3244 21286 3282
rect 21344 3282 21434 3299
rect 21654 3299 21670 3316
rect 21876 3316 22128 3332
rect 21876 3299 21892 3316
rect 21654 3282 21744 3299
rect 21344 3244 21744 3282
rect 21802 3282 21892 3299
rect 22112 3299 22128 3316
rect 22112 3282 22202 3299
rect 21802 3244 22202 3282
rect 17680 3006 18080 3044
rect 17680 2989 17770 3006
rect 17754 2972 17770 2989
rect 17990 2989 18080 3006
rect 18138 3006 18538 3044
rect 18138 2989 18228 3006
rect 17990 2972 18006 2989
rect 17754 2956 18006 2972
rect 18212 2972 18228 2989
rect 18448 2989 18538 3006
rect 18596 3006 18996 3044
rect 18596 2989 18686 3006
rect 18448 2972 18464 2989
rect 18212 2956 18464 2972
rect 18670 2972 18686 2989
rect 18906 2989 18996 3006
rect 19054 3006 19454 3044
rect 19054 2989 19144 3006
rect 18906 2972 18922 2989
rect 18670 2956 18922 2972
rect 19128 2972 19144 2989
rect 19364 2989 19454 3006
rect 19512 3006 19912 3044
rect 19512 2989 19602 3006
rect 19364 2972 19380 2989
rect 19128 2956 19380 2972
rect 19586 2972 19602 2989
rect 19822 2989 19912 3006
rect 19970 3006 20370 3044
rect 19970 2989 20060 3006
rect 19822 2972 19838 2989
rect 19586 2956 19838 2972
rect 20044 2972 20060 2989
rect 20280 2989 20370 3006
rect 20428 3006 20828 3044
rect 20428 2989 20518 3006
rect 20280 2972 20296 2989
rect 20044 2956 20296 2972
rect 20502 2972 20518 2989
rect 20738 2989 20828 3006
rect 20886 3006 21286 3044
rect 20886 2989 20976 3006
rect 20738 2972 20754 2989
rect 20502 2956 20754 2972
rect 20960 2972 20976 2989
rect 21196 2989 21286 3006
rect 21344 3006 21744 3044
rect 21344 2989 21434 3006
rect 21196 2972 21212 2989
rect 20960 2956 21212 2972
rect 21418 2972 21434 2989
rect 21654 2989 21744 3006
rect 21802 3006 22202 3044
rect 21802 2989 21892 3006
rect 21654 2972 21670 2989
rect 21418 2956 21670 2972
rect 21876 2972 21892 2989
rect 22112 2989 22202 3006
rect 22112 2972 22128 2989
rect 21876 2956 22128 2972
rect 26516 3316 26768 3332
rect 26516 3299 26532 3316
rect 26442 3282 26532 3299
rect 26752 3299 26768 3316
rect 26974 3316 27226 3332
rect 26974 3299 26990 3316
rect 26752 3282 26842 3299
rect 26442 3244 26842 3282
rect 26900 3282 26990 3299
rect 27210 3299 27226 3316
rect 27432 3316 27684 3332
rect 27432 3299 27448 3316
rect 27210 3282 27300 3299
rect 26900 3244 27300 3282
rect 27358 3282 27448 3299
rect 27668 3299 27684 3316
rect 27890 3316 28142 3332
rect 27890 3299 27906 3316
rect 27668 3282 27758 3299
rect 27358 3244 27758 3282
rect 27816 3282 27906 3299
rect 28126 3299 28142 3316
rect 28348 3316 28600 3332
rect 28348 3299 28364 3316
rect 28126 3282 28216 3299
rect 27816 3244 28216 3282
rect 28274 3282 28364 3299
rect 28584 3299 28600 3316
rect 28806 3316 29058 3332
rect 28806 3299 28822 3316
rect 28584 3282 28674 3299
rect 28274 3244 28674 3282
rect 28732 3282 28822 3299
rect 29042 3299 29058 3316
rect 29264 3316 29516 3332
rect 29264 3299 29280 3316
rect 29042 3282 29132 3299
rect 28732 3244 29132 3282
rect 29190 3282 29280 3299
rect 29500 3299 29516 3316
rect 29722 3316 29974 3332
rect 29722 3299 29738 3316
rect 29500 3282 29590 3299
rect 29190 3244 29590 3282
rect 29648 3282 29738 3299
rect 29958 3299 29974 3316
rect 30180 3316 30432 3332
rect 30180 3299 30196 3316
rect 29958 3282 30048 3299
rect 29648 3244 30048 3282
rect 30106 3282 30196 3299
rect 30416 3299 30432 3316
rect 30638 3316 30890 3332
rect 30638 3299 30654 3316
rect 30416 3282 30506 3299
rect 30106 3244 30506 3282
rect 30564 3282 30654 3299
rect 30874 3299 30890 3316
rect 30874 3282 30964 3299
rect 30564 3244 30964 3282
rect 26442 3006 26842 3044
rect 26442 2989 26532 3006
rect 26516 2972 26532 2989
rect 26752 2989 26842 3006
rect 26900 3006 27300 3044
rect 26900 2989 26990 3006
rect 26752 2972 26768 2989
rect 26516 2956 26768 2972
rect 26974 2972 26990 2989
rect 27210 2989 27300 3006
rect 27358 3006 27758 3044
rect 27358 2989 27448 3006
rect 27210 2972 27226 2989
rect 26974 2956 27226 2972
rect 27432 2972 27448 2989
rect 27668 2989 27758 3006
rect 27816 3006 28216 3044
rect 27816 2989 27906 3006
rect 27668 2972 27684 2989
rect 27432 2956 27684 2972
rect 27890 2972 27906 2989
rect 28126 2989 28216 3006
rect 28274 3006 28674 3044
rect 28274 2989 28364 3006
rect 28126 2972 28142 2989
rect 27890 2956 28142 2972
rect 28348 2972 28364 2989
rect 28584 2989 28674 3006
rect 28732 3006 29132 3044
rect 28732 2989 28822 3006
rect 28584 2972 28600 2989
rect 28348 2956 28600 2972
rect 28806 2972 28822 2989
rect 29042 2989 29132 3006
rect 29190 3006 29590 3044
rect 29190 2989 29280 3006
rect 29042 2972 29058 2989
rect 28806 2956 29058 2972
rect 29264 2972 29280 2989
rect 29500 2989 29590 3006
rect 29648 3006 30048 3044
rect 29648 2989 29738 3006
rect 29500 2972 29516 2989
rect 29264 2956 29516 2972
rect 29722 2972 29738 2989
rect 29958 2989 30048 3006
rect 30106 3006 30506 3044
rect 30106 2989 30196 3006
rect 29958 2972 29974 2989
rect 29722 2956 29974 2972
rect 30180 2972 30196 2989
rect 30416 2989 30506 3006
rect 30564 3006 30964 3044
rect 30564 2989 30654 3006
rect 30416 2972 30432 2989
rect 30180 2956 30432 2972
rect 30638 2972 30654 2989
rect 30874 2989 30964 3006
rect 30874 2972 30890 2989
rect 30638 2956 30890 2972
rect 31662 2443 31692 2469
rect 31907 2443 31937 2469
rect 31991 2443 32021 2469
rect 32075 2443 32105 2469
rect 32159 2443 32189 2469
rect 31662 2291 31692 2313
rect 31907 2291 31937 2313
rect 31991 2291 32021 2313
rect 32075 2291 32105 2313
rect 32159 2291 32189 2313
rect 31606 2275 31692 2291
rect 31606 2241 31622 2275
rect 31656 2241 31692 2275
rect 31606 2225 31692 2241
rect 31839 2275 32189 2291
rect 31839 2241 31855 2275
rect 31889 2241 31947 2275
rect 31981 2241 32031 2275
rect 32065 2241 32115 2275
rect 32149 2241 32189 2275
rect 31839 2225 32189 2241
rect 15922 1474 16174 1490
rect 15922 1457 15938 1474
rect 15848 1440 15938 1457
rect 16158 1457 16174 1474
rect 16380 1474 16632 1490
rect 16380 1457 16396 1474
rect 16158 1440 16248 1457
rect 15848 1393 16248 1440
rect 16306 1440 16396 1457
rect 16616 1457 16632 1474
rect 16838 1474 17090 1490
rect 16838 1457 16854 1474
rect 16616 1440 16706 1457
rect 16306 1393 16706 1440
rect 16764 1440 16854 1457
rect 17074 1457 17090 1474
rect 17296 1474 17548 1490
rect 17296 1457 17312 1474
rect 17074 1440 17164 1457
rect 16764 1393 17164 1440
rect 17222 1440 17312 1457
rect 17532 1457 17548 1474
rect 17754 1474 18006 1490
rect 17754 1457 17770 1474
rect 17532 1440 17622 1457
rect 17222 1393 17622 1440
rect 17680 1440 17770 1457
rect 17990 1457 18006 1474
rect 18212 1474 18464 1490
rect 18212 1457 18228 1474
rect 17990 1440 18080 1457
rect 17680 1393 18080 1440
rect 18138 1440 18228 1457
rect 18448 1457 18464 1474
rect 18670 1474 18922 1490
rect 18670 1457 18686 1474
rect 18448 1440 18538 1457
rect 18138 1393 18538 1440
rect 18596 1440 18686 1457
rect 18906 1457 18922 1474
rect 19128 1474 19380 1490
rect 19128 1457 19144 1474
rect 18906 1440 18996 1457
rect 18596 1393 18996 1440
rect 19054 1440 19144 1457
rect 19364 1457 19380 1474
rect 19586 1474 19838 1490
rect 19586 1457 19602 1474
rect 19364 1440 19454 1457
rect 19054 1393 19454 1440
rect 19512 1440 19602 1457
rect 19822 1457 19838 1474
rect 20044 1474 20296 1490
rect 20044 1457 20060 1474
rect 19822 1440 19912 1457
rect 19512 1393 19912 1440
rect 19970 1440 20060 1457
rect 20280 1457 20296 1474
rect 20502 1474 20754 1490
rect 20502 1457 20518 1474
rect 20280 1440 20370 1457
rect 19970 1393 20370 1440
rect 20428 1440 20518 1457
rect 20738 1457 20754 1474
rect 20960 1474 21212 1490
rect 20960 1457 20976 1474
rect 20738 1440 20828 1457
rect 20428 1393 20828 1440
rect 20886 1440 20976 1457
rect 21196 1457 21212 1474
rect 21418 1474 21670 1490
rect 21418 1457 21434 1474
rect 21196 1440 21286 1457
rect 20886 1393 21286 1440
rect 21344 1440 21434 1457
rect 21654 1457 21670 1474
rect 21876 1474 22128 1490
rect 21876 1457 21892 1474
rect 21654 1440 21744 1457
rect 21344 1393 21744 1440
rect 21802 1440 21892 1457
rect 22112 1457 22128 1474
rect 22334 1474 22586 1490
rect 22334 1457 22350 1474
rect 22112 1440 22202 1457
rect 21802 1393 22202 1440
rect 22260 1440 22350 1457
rect 22570 1457 22586 1474
rect 22792 1474 23044 1490
rect 22792 1457 22808 1474
rect 22570 1440 22660 1457
rect 22260 1393 22660 1440
rect 22718 1440 22808 1457
rect 23028 1457 23044 1474
rect 23250 1474 23502 1490
rect 23250 1457 23266 1474
rect 23028 1440 23118 1457
rect 22718 1393 23118 1440
rect 23176 1440 23266 1457
rect 23486 1457 23502 1474
rect 23708 1474 23960 1490
rect 23708 1457 23724 1474
rect 23486 1440 23576 1457
rect 23176 1393 23576 1440
rect 23634 1440 23724 1457
rect 23944 1457 23960 1474
rect 23944 1440 24034 1457
rect 23634 1393 24034 1440
rect 15848 -254 16248 -207
rect 15848 -271 15938 -254
rect 15922 -288 15938 -271
rect 16158 -271 16248 -254
rect 16306 -254 16706 -207
rect 16306 -271 16396 -254
rect 16158 -288 16174 -271
rect 15922 -304 16174 -288
rect 16380 -288 16396 -271
rect 16616 -271 16706 -254
rect 16764 -254 17164 -207
rect 16764 -271 16854 -254
rect 16616 -288 16632 -271
rect 16380 -304 16632 -288
rect 16838 -288 16854 -271
rect 17074 -271 17164 -254
rect 17222 -254 17622 -207
rect 17222 -271 17312 -254
rect 17074 -288 17090 -271
rect 16838 -304 17090 -288
rect 17296 -288 17312 -271
rect 17532 -271 17622 -254
rect 17680 -254 18080 -207
rect 17680 -271 17770 -254
rect 17532 -288 17548 -271
rect 17296 -304 17548 -288
rect 17754 -288 17770 -271
rect 17990 -271 18080 -254
rect 18138 -254 18538 -207
rect 18138 -271 18228 -254
rect 17990 -288 18006 -271
rect 17754 -304 18006 -288
rect 18212 -288 18228 -271
rect 18448 -271 18538 -254
rect 18596 -254 18996 -207
rect 18596 -271 18686 -254
rect 18448 -288 18464 -271
rect 18212 -304 18464 -288
rect 18670 -288 18686 -271
rect 18906 -271 18996 -254
rect 19054 -254 19454 -207
rect 19054 -271 19144 -254
rect 18906 -288 18922 -271
rect 18670 -304 18922 -288
rect 19128 -288 19144 -271
rect 19364 -271 19454 -254
rect 19512 -254 19912 -207
rect 19512 -271 19602 -254
rect 19364 -288 19380 -271
rect 19128 -304 19380 -288
rect 19586 -288 19602 -271
rect 19822 -271 19912 -254
rect 19970 -254 20370 -207
rect 19970 -271 20060 -254
rect 19822 -288 19838 -271
rect 19586 -304 19838 -288
rect 20044 -288 20060 -271
rect 20280 -271 20370 -254
rect 20428 -254 20828 -207
rect 20428 -271 20518 -254
rect 20280 -288 20296 -271
rect 20044 -304 20296 -288
rect 20502 -288 20518 -271
rect 20738 -271 20828 -254
rect 20886 -254 21286 -207
rect 20886 -271 20976 -254
rect 20738 -288 20754 -271
rect 20502 -304 20754 -288
rect 20960 -288 20976 -271
rect 21196 -271 21286 -254
rect 21344 -254 21744 -207
rect 21344 -271 21434 -254
rect 21196 -288 21212 -271
rect 20960 -304 21212 -288
rect 21418 -288 21434 -271
rect 21654 -271 21744 -254
rect 21802 -254 22202 -207
rect 21802 -271 21892 -254
rect 21654 -288 21670 -271
rect 21418 -304 21670 -288
rect 21876 -288 21892 -271
rect 22112 -271 22202 -254
rect 22260 -254 22660 -207
rect 22260 -271 22350 -254
rect 22112 -288 22128 -271
rect 21876 -304 22128 -288
rect 22334 -288 22350 -271
rect 22570 -271 22660 -254
rect 22718 -254 23118 -207
rect 22718 -271 22808 -254
rect 22570 -288 22586 -271
rect 22334 -304 22586 -288
rect 22792 -288 22808 -271
rect 23028 -271 23118 -254
rect 23176 -254 23576 -207
rect 23176 -271 23266 -254
rect 23028 -288 23044 -271
rect 22792 -304 23044 -288
rect 23250 -288 23266 -271
rect 23486 -271 23576 -254
rect 23634 -254 24034 -207
rect 23634 -271 23724 -254
rect 23486 -288 23502 -271
rect 23250 -304 23502 -288
rect 23708 -288 23724 -271
rect 23944 -271 24034 -254
rect 23944 -288 23960 -271
rect 23708 -304 23960 -288
rect 31662 2193 31692 2225
rect 31907 2193 31937 2225
rect 31991 2193 32021 2225
rect 32075 2193 32105 2225
rect 32159 2193 32189 2225
rect 26517 1894 26769 1910
rect 26517 1877 26533 1894
rect 26443 1860 26533 1877
rect 26753 1877 26769 1894
rect 26975 1894 27227 1910
rect 26975 1877 26991 1894
rect 26753 1860 26843 1877
rect 26443 1813 26843 1860
rect 26901 1860 26991 1877
rect 27211 1877 27227 1894
rect 27433 1894 27685 1910
rect 27433 1877 27449 1894
rect 27211 1860 27301 1877
rect 26901 1813 27301 1860
rect 27359 1860 27449 1877
rect 27669 1877 27685 1894
rect 27891 1894 28143 1910
rect 27891 1877 27907 1894
rect 27669 1860 27759 1877
rect 27359 1813 27759 1860
rect 27817 1860 27907 1877
rect 28127 1877 28143 1894
rect 28349 1894 28601 1910
rect 28349 1877 28365 1894
rect 28127 1860 28217 1877
rect 27817 1813 28217 1860
rect 28275 1860 28365 1877
rect 28585 1877 28601 1894
rect 28807 1894 29059 1910
rect 28807 1877 28823 1894
rect 28585 1860 28675 1877
rect 28275 1813 28675 1860
rect 28733 1860 28823 1877
rect 29043 1877 29059 1894
rect 29265 1894 29517 1910
rect 29265 1877 29281 1894
rect 29043 1860 29133 1877
rect 28733 1813 29133 1860
rect 29191 1860 29281 1877
rect 29501 1877 29517 1894
rect 29723 1894 29975 1910
rect 29723 1877 29739 1894
rect 29501 1860 29591 1877
rect 29191 1813 29591 1860
rect 29649 1860 29739 1877
rect 29959 1877 29975 1894
rect 30181 1894 30433 1910
rect 30181 1877 30197 1894
rect 29959 1860 30049 1877
rect 29649 1813 30049 1860
rect 30107 1860 30197 1877
rect 30417 1877 30433 1894
rect 30639 1894 30891 1910
rect 30639 1877 30655 1894
rect 30417 1860 30507 1877
rect 30107 1813 30507 1860
rect 30565 1860 30655 1877
rect 30875 1877 30891 1894
rect 30875 1860 30965 1877
rect 30565 1813 30965 1860
rect 26443 566 26843 613
rect 26443 549 26533 566
rect 26517 532 26533 549
rect 26753 549 26843 566
rect 26901 566 27301 613
rect 26901 549 26991 566
rect 26753 532 26769 549
rect 26517 516 26769 532
rect 26975 532 26991 549
rect 27211 549 27301 566
rect 27359 566 27759 613
rect 27359 549 27449 566
rect 27211 532 27227 549
rect 26975 516 27227 532
rect 27433 532 27449 549
rect 27669 549 27759 566
rect 27817 566 28217 613
rect 27817 549 27907 566
rect 27669 532 27685 549
rect 27433 516 27685 532
rect 27891 532 27907 549
rect 28127 549 28217 566
rect 28275 566 28675 613
rect 28275 549 28365 566
rect 28127 532 28143 549
rect 27891 516 28143 532
rect 28349 532 28365 549
rect 28585 549 28675 566
rect 28733 566 29133 613
rect 28733 549 28823 566
rect 28585 532 28601 549
rect 28349 516 28601 532
rect 28807 532 28823 549
rect 29043 549 29133 566
rect 29191 566 29591 613
rect 29191 549 29281 566
rect 29043 532 29059 549
rect 28807 516 29059 532
rect 29265 532 29281 549
rect 29501 549 29591 566
rect 29649 566 30049 613
rect 29649 549 29739 566
rect 29501 532 29517 549
rect 29265 516 29517 532
rect 29723 532 29739 549
rect 29959 549 30049 566
rect 30107 566 30507 613
rect 30107 549 30197 566
rect 29959 532 29975 549
rect 29723 516 29975 532
rect 30181 532 30197 549
rect 30417 549 30507 566
rect 30565 566 30965 613
rect 30565 549 30655 566
rect 30417 532 30433 549
rect 30181 516 30433 532
rect 30639 532 30655 549
rect 30875 549 30965 566
rect 30875 532 30891 549
rect 30639 516 30891 532
rect 31662 1967 31692 1993
rect 31907 1967 31937 1993
rect 31991 1967 32021 1993
rect 32075 1967 32105 1993
rect 32159 1967 32189 1993
rect 11924 -3399 12176 -3383
rect 11924 -3416 11940 -3399
rect 11850 -3433 11940 -3416
rect 12160 -3416 12176 -3399
rect 12382 -3399 12634 -3383
rect 12382 -3416 12398 -3399
rect 12160 -3433 12250 -3416
rect 11850 -3480 12250 -3433
rect 12308 -3433 12398 -3416
rect 12618 -3416 12634 -3399
rect 12840 -3399 13092 -3383
rect 12840 -3416 12856 -3399
rect 12618 -3433 12708 -3416
rect 12308 -3480 12708 -3433
rect 12766 -3433 12856 -3416
rect 13076 -3416 13092 -3399
rect 13298 -3399 13550 -3383
rect 13298 -3416 13314 -3399
rect 13076 -3433 13166 -3416
rect 12766 -3480 13166 -3433
rect 13224 -3433 13314 -3416
rect 13534 -3416 13550 -3399
rect 13756 -3399 14008 -3383
rect 13756 -3416 13772 -3399
rect 13534 -3433 13624 -3416
rect 13224 -3480 13624 -3433
rect 13682 -3433 13772 -3416
rect 13992 -3416 14008 -3399
rect 14214 -3399 14466 -3383
rect 14214 -3416 14230 -3399
rect 13992 -3433 14082 -3416
rect 13682 -3480 14082 -3433
rect 14140 -3433 14230 -3416
rect 14450 -3416 14466 -3399
rect 14672 -3399 14924 -3383
rect 14672 -3416 14688 -3399
rect 14450 -3433 14540 -3416
rect 14140 -3480 14540 -3433
rect 14598 -3433 14688 -3416
rect 14908 -3416 14924 -3399
rect 15130 -3399 15382 -3383
rect 15130 -3416 15146 -3399
rect 14908 -3433 14998 -3416
rect 14598 -3480 14998 -3433
rect 15056 -3433 15146 -3416
rect 15366 -3416 15382 -3399
rect 15588 -3399 15840 -3383
rect 15588 -3416 15604 -3399
rect 15366 -3433 15456 -3416
rect 15056 -3480 15456 -3433
rect 15514 -3433 15604 -3416
rect 15824 -3416 15840 -3399
rect 16046 -3399 16298 -3383
rect 16046 -3416 16062 -3399
rect 15824 -3433 15914 -3416
rect 15514 -3480 15914 -3433
rect 15972 -3433 16062 -3416
rect 16282 -3416 16298 -3399
rect 16504 -3399 16756 -3383
rect 16504 -3416 16520 -3399
rect 16282 -3433 16372 -3416
rect 15972 -3480 16372 -3433
rect 16430 -3433 16520 -3416
rect 16740 -3416 16756 -3399
rect 16962 -3399 17214 -3383
rect 16962 -3416 16978 -3399
rect 16740 -3433 16830 -3416
rect 16430 -3480 16830 -3433
rect 16888 -3433 16978 -3416
rect 17198 -3416 17214 -3399
rect 17420 -3399 17672 -3383
rect 17420 -3416 17436 -3399
rect 17198 -3433 17288 -3416
rect 16888 -3480 17288 -3433
rect 17346 -3433 17436 -3416
rect 17656 -3416 17672 -3399
rect 17878 -3399 18130 -3383
rect 17878 -3416 17894 -3399
rect 17656 -3433 17746 -3416
rect 17346 -3480 17746 -3433
rect 17804 -3433 17894 -3416
rect 18114 -3416 18130 -3399
rect 18336 -3399 18588 -3383
rect 18336 -3416 18352 -3399
rect 18114 -3433 18204 -3416
rect 17804 -3480 18204 -3433
rect 18262 -3433 18352 -3416
rect 18572 -3416 18588 -3399
rect 18794 -3399 19046 -3383
rect 18794 -3416 18810 -3399
rect 18572 -3433 18662 -3416
rect 18262 -3480 18662 -3433
rect 18720 -3433 18810 -3416
rect 19030 -3416 19046 -3399
rect 19252 -3399 19504 -3383
rect 19252 -3416 19268 -3399
rect 19030 -3433 19120 -3416
rect 18720 -3480 19120 -3433
rect 19178 -3433 19268 -3416
rect 19488 -3416 19504 -3399
rect 19710 -3399 19962 -3383
rect 19710 -3416 19726 -3399
rect 19488 -3433 19578 -3416
rect 19178 -3480 19578 -3433
rect 19636 -3433 19726 -3416
rect 19946 -3416 19962 -3399
rect 19946 -3433 20036 -3416
rect 19636 -3480 20036 -3433
rect 11850 -5127 12250 -5080
rect 11850 -5144 11940 -5127
rect 11924 -5161 11940 -5144
rect 12160 -5144 12250 -5127
rect 12308 -5127 12708 -5080
rect 12308 -5144 12398 -5127
rect 12160 -5161 12176 -5144
rect 11924 -5177 12176 -5161
rect 12382 -5161 12398 -5144
rect 12618 -5144 12708 -5127
rect 12766 -5127 13166 -5080
rect 12766 -5144 12856 -5127
rect 12618 -5161 12634 -5144
rect 12382 -5177 12634 -5161
rect 12840 -5161 12856 -5144
rect 13076 -5144 13166 -5127
rect 13224 -5127 13624 -5080
rect 13224 -5144 13314 -5127
rect 13076 -5161 13092 -5144
rect 12840 -5177 13092 -5161
rect 13298 -5161 13314 -5144
rect 13534 -5144 13624 -5127
rect 13682 -5127 14082 -5080
rect 13682 -5144 13772 -5127
rect 13534 -5161 13550 -5144
rect 13298 -5177 13550 -5161
rect 13756 -5161 13772 -5144
rect 13992 -5144 14082 -5127
rect 14140 -5127 14540 -5080
rect 14140 -5144 14230 -5127
rect 13992 -5161 14008 -5144
rect 13756 -5177 14008 -5161
rect 14214 -5161 14230 -5144
rect 14450 -5144 14540 -5127
rect 14598 -5127 14998 -5080
rect 14598 -5144 14688 -5127
rect 14450 -5161 14466 -5144
rect 14214 -5177 14466 -5161
rect 14672 -5161 14688 -5144
rect 14908 -5144 14998 -5127
rect 15056 -5127 15456 -5080
rect 15056 -5144 15146 -5127
rect 14908 -5161 14924 -5144
rect 14672 -5177 14924 -5161
rect 15130 -5161 15146 -5144
rect 15366 -5144 15456 -5127
rect 15514 -5127 15914 -5080
rect 15514 -5144 15604 -5127
rect 15366 -5161 15382 -5144
rect 15130 -5177 15382 -5161
rect 15588 -5161 15604 -5144
rect 15824 -5144 15914 -5127
rect 15972 -5127 16372 -5080
rect 15972 -5144 16062 -5127
rect 15824 -5161 15840 -5144
rect 15588 -5177 15840 -5161
rect 16046 -5161 16062 -5144
rect 16282 -5144 16372 -5127
rect 16430 -5127 16830 -5080
rect 16430 -5144 16520 -5127
rect 16282 -5161 16298 -5144
rect 16046 -5177 16298 -5161
rect 16504 -5161 16520 -5144
rect 16740 -5144 16830 -5127
rect 16888 -5127 17288 -5080
rect 16888 -5144 16978 -5127
rect 16740 -5161 16756 -5144
rect 16504 -5177 16756 -5161
rect 16962 -5161 16978 -5144
rect 17198 -5144 17288 -5127
rect 17346 -5127 17746 -5080
rect 17346 -5144 17436 -5127
rect 17198 -5161 17214 -5144
rect 16962 -5177 17214 -5161
rect 17420 -5161 17436 -5144
rect 17656 -5144 17746 -5127
rect 17804 -5127 18204 -5080
rect 17804 -5144 17894 -5127
rect 17656 -5161 17672 -5144
rect 17420 -5177 17672 -5161
rect 17878 -5161 17894 -5144
rect 18114 -5144 18204 -5127
rect 18262 -5127 18662 -5080
rect 18262 -5144 18352 -5127
rect 18114 -5161 18130 -5144
rect 17878 -5177 18130 -5161
rect 18336 -5161 18352 -5144
rect 18572 -5144 18662 -5127
rect 18720 -5127 19120 -5080
rect 18720 -5144 18810 -5127
rect 18572 -5161 18588 -5144
rect 18336 -5177 18588 -5161
rect 18794 -5161 18810 -5144
rect 19030 -5144 19120 -5127
rect 19178 -5127 19578 -5080
rect 19178 -5144 19268 -5127
rect 19030 -5161 19046 -5144
rect 18794 -5177 19046 -5161
rect 19252 -5161 19268 -5144
rect 19488 -5144 19578 -5127
rect 19636 -5127 20036 -5080
rect 19636 -5144 19726 -5127
rect 19488 -5161 19504 -5144
rect 19252 -5177 19504 -5161
rect 19710 -5161 19726 -5144
rect 19946 -5144 20036 -5127
rect 19946 -5161 19962 -5144
rect 19710 -5177 19962 -5161
rect 11365 -6064 11617 -6048
rect 11365 -6081 11381 -6064
rect 11291 -6098 11381 -6081
rect 11601 -6081 11617 -6064
rect 11823 -6064 12075 -6048
rect 11823 -6081 11839 -6064
rect 11601 -6098 11691 -6081
rect 11291 -6145 11691 -6098
rect 11749 -6098 11839 -6081
rect 12059 -6081 12075 -6064
rect 12281 -6064 12533 -6048
rect 12281 -6081 12297 -6064
rect 12059 -6098 12149 -6081
rect 11749 -6145 12149 -6098
rect 12207 -6098 12297 -6081
rect 12517 -6081 12533 -6064
rect 12739 -6064 12991 -6048
rect 12739 -6081 12755 -6064
rect 12517 -6098 12607 -6081
rect 12207 -6145 12607 -6098
rect 12665 -6098 12755 -6081
rect 12975 -6081 12991 -6064
rect 13197 -6064 13449 -6048
rect 13197 -6081 13213 -6064
rect 12975 -6098 13065 -6081
rect 12665 -6145 13065 -6098
rect 13123 -6098 13213 -6081
rect 13433 -6081 13449 -6064
rect 13655 -6064 13907 -6048
rect 13655 -6081 13671 -6064
rect 13433 -6098 13523 -6081
rect 13123 -6145 13523 -6098
rect 13581 -6098 13671 -6081
rect 13891 -6081 13907 -6064
rect 14113 -6064 14365 -6048
rect 14113 -6081 14129 -6064
rect 13891 -6098 13981 -6081
rect 13581 -6145 13981 -6098
rect 14039 -6098 14129 -6081
rect 14349 -6081 14365 -6064
rect 14571 -6064 14823 -6048
rect 14571 -6081 14587 -6064
rect 14349 -6098 14439 -6081
rect 14039 -6145 14439 -6098
rect 14497 -6098 14587 -6081
rect 14807 -6081 14823 -6064
rect 15029 -6064 15281 -6048
rect 15029 -6081 15045 -6064
rect 14807 -6098 14897 -6081
rect 14497 -6145 14897 -6098
rect 14955 -6098 15045 -6081
rect 15265 -6081 15281 -6064
rect 15487 -6064 15739 -6048
rect 15487 -6081 15503 -6064
rect 15265 -6098 15355 -6081
rect 14955 -6145 15355 -6098
rect 15413 -6098 15503 -6081
rect 15723 -6081 15739 -6064
rect 16365 -6064 16617 -6048
rect 16365 -6081 16381 -6064
rect 15723 -6098 15813 -6081
rect 15413 -6145 15813 -6098
rect 16291 -6098 16381 -6081
rect 16601 -6081 16617 -6064
rect 16823 -6064 17075 -6048
rect 16823 -6081 16839 -6064
rect 16601 -6098 16691 -6081
rect 16291 -6145 16691 -6098
rect 16749 -6098 16839 -6081
rect 17059 -6081 17075 -6064
rect 17281 -6064 17533 -6048
rect 17281 -6081 17297 -6064
rect 17059 -6098 17149 -6081
rect 16749 -6145 17149 -6098
rect 17207 -6098 17297 -6081
rect 17517 -6081 17533 -6064
rect 17739 -6064 17991 -6048
rect 17739 -6081 17755 -6064
rect 17517 -6098 17607 -6081
rect 17207 -6145 17607 -6098
rect 17665 -6098 17755 -6081
rect 17975 -6081 17991 -6064
rect 18197 -6064 18449 -6048
rect 18197 -6081 18213 -6064
rect 17975 -6098 18065 -6081
rect 17665 -6145 18065 -6098
rect 18123 -6098 18213 -6081
rect 18433 -6081 18449 -6064
rect 18655 -6064 18907 -6048
rect 18655 -6081 18671 -6064
rect 18433 -6098 18523 -6081
rect 18123 -6145 18523 -6098
rect 18581 -6098 18671 -6081
rect 18891 -6081 18907 -6064
rect 19113 -6064 19365 -6048
rect 19113 -6081 19129 -6064
rect 18891 -6098 18981 -6081
rect 18581 -6145 18981 -6098
rect 19039 -6098 19129 -6081
rect 19349 -6081 19365 -6064
rect 19571 -6064 19823 -6048
rect 19571 -6081 19587 -6064
rect 19349 -6098 19439 -6081
rect 19039 -6145 19439 -6098
rect 19497 -6098 19587 -6081
rect 19807 -6081 19823 -6064
rect 20029 -6064 20281 -6048
rect 20029 -6081 20045 -6064
rect 19807 -6098 19897 -6081
rect 19497 -6145 19897 -6098
rect 19955 -6098 20045 -6081
rect 20265 -6081 20281 -6064
rect 20487 -6064 20739 -6048
rect 20487 -6081 20503 -6064
rect 20265 -6098 20355 -6081
rect 19955 -6145 20355 -6098
rect 20413 -6098 20503 -6081
rect 20723 -6081 20739 -6064
rect 20723 -6098 20813 -6081
rect 20413 -6145 20813 -6098
rect 11291 -7392 11691 -7345
rect 11291 -7409 11381 -7392
rect 11365 -7426 11381 -7409
rect 11601 -7409 11691 -7392
rect 11749 -7392 12149 -7345
rect 11749 -7409 11839 -7392
rect 11601 -7426 11617 -7409
rect 11365 -7442 11617 -7426
rect 11823 -7426 11839 -7409
rect 12059 -7409 12149 -7392
rect 12207 -7392 12607 -7345
rect 12207 -7409 12297 -7392
rect 12059 -7426 12075 -7409
rect 11823 -7442 12075 -7426
rect 12281 -7426 12297 -7409
rect 12517 -7409 12607 -7392
rect 12665 -7392 13065 -7345
rect 12665 -7409 12755 -7392
rect 12517 -7426 12533 -7409
rect 12281 -7442 12533 -7426
rect 12739 -7426 12755 -7409
rect 12975 -7409 13065 -7392
rect 13123 -7392 13523 -7345
rect 13123 -7409 13213 -7392
rect 12975 -7426 12991 -7409
rect 12739 -7442 12991 -7426
rect 13197 -7426 13213 -7409
rect 13433 -7409 13523 -7392
rect 13581 -7392 13981 -7345
rect 13581 -7409 13671 -7392
rect 13433 -7426 13449 -7409
rect 13197 -7442 13449 -7426
rect 13655 -7426 13671 -7409
rect 13891 -7409 13981 -7392
rect 14039 -7392 14439 -7345
rect 14039 -7409 14129 -7392
rect 13891 -7426 13907 -7409
rect 13655 -7442 13907 -7426
rect 14113 -7426 14129 -7409
rect 14349 -7409 14439 -7392
rect 14497 -7392 14897 -7345
rect 14497 -7409 14587 -7392
rect 14349 -7426 14365 -7409
rect 14113 -7442 14365 -7426
rect 14571 -7426 14587 -7409
rect 14807 -7409 14897 -7392
rect 14955 -7392 15355 -7345
rect 14955 -7409 15045 -7392
rect 14807 -7426 14823 -7409
rect 14571 -7442 14823 -7426
rect 15029 -7426 15045 -7409
rect 15265 -7409 15355 -7392
rect 15413 -7392 15813 -7345
rect 15413 -7409 15503 -7392
rect 15265 -7426 15281 -7409
rect 15029 -7442 15281 -7426
rect 15487 -7426 15503 -7409
rect 15723 -7409 15813 -7392
rect 16291 -7392 16691 -7345
rect 16291 -7409 16381 -7392
rect 15723 -7426 15739 -7409
rect 15487 -7442 15739 -7426
rect 16365 -7426 16381 -7409
rect 16601 -7409 16691 -7392
rect 16749 -7392 17149 -7345
rect 16749 -7409 16839 -7392
rect 16601 -7426 16617 -7409
rect 16365 -7442 16617 -7426
rect 16823 -7426 16839 -7409
rect 17059 -7409 17149 -7392
rect 17207 -7392 17607 -7345
rect 17207 -7409 17297 -7392
rect 17059 -7426 17075 -7409
rect 16823 -7442 17075 -7426
rect 17281 -7426 17297 -7409
rect 17517 -7409 17607 -7392
rect 17665 -7392 18065 -7345
rect 17665 -7409 17755 -7392
rect 17517 -7426 17533 -7409
rect 17281 -7442 17533 -7426
rect 17739 -7426 17755 -7409
rect 17975 -7409 18065 -7392
rect 18123 -7392 18523 -7345
rect 18123 -7409 18213 -7392
rect 17975 -7426 17991 -7409
rect 17739 -7442 17991 -7426
rect 18197 -7426 18213 -7409
rect 18433 -7409 18523 -7392
rect 18581 -7392 18981 -7345
rect 18581 -7409 18671 -7392
rect 18433 -7426 18449 -7409
rect 18197 -7442 18449 -7426
rect 18655 -7426 18671 -7409
rect 18891 -7409 18981 -7392
rect 19039 -7392 19439 -7345
rect 19039 -7409 19129 -7392
rect 18891 -7426 18907 -7409
rect 18655 -7442 18907 -7426
rect 19113 -7426 19129 -7409
rect 19349 -7409 19439 -7392
rect 19497 -7392 19897 -7345
rect 19497 -7409 19587 -7392
rect 19349 -7426 19365 -7409
rect 19113 -7442 19365 -7426
rect 19571 -7426 19587 -7409
rect 19807 -7409 19897 -7392
rect 19955 -7392 20355 -7345
rect 19955 -7409 20045 -7392
rect 19807 -7426 19823 -7409
rect 19571 -7442 19823 -7426
rect 20029 -7426 20045 -7409
rect 20265 -7409 20355 -7392
rect 20413 -7392 20813 -7345
rect 20413 -7409 20503 -7392
rect 20265 -7426 20281 -7409
rect 20029 -7442 20281 -7426
rect 20487 -7426 20503 -7409
rect 20723 -7409 20813 -7392
rect 20723 -7426 20739 -7409
rect 20487 -7442 20739 -7426
rect 26924 -3399 27176 -3383
rect 26924 -3416 26940 -3399
rect 26850 -3433 26940 -3416
rect 27160 -3416 27176 -3399
rect 27382 -3399 27634 -3383
rect 27382 -3416 27398 -3399
rect 27160 -3433 27250 -3416
rect 26850 -3480 27250 -3433
rect 27308 -3433 27398 -3416
rect 27618 -3416 27634 -3399
rect 27840 -3399 28092 -3383
rect 27840 -3416 27856 -3399
rect 27618 -3433 27708 -3416
rect 27308 -3480 27708 -3433
rect 27766 -3433 27856 -3416
rect 28076 -3416 28092 -3399
rect 28298 -3399 28550 -3383
rect 28298 -3416 28314 -3399
rect 28076 -3433 28166 -3416
rect 27766 -3480 28166 -3433
rect 28224 -3433 28314 -3416
rect 28534 -3416 28550 -3399
rect 28756 -3399 29008 -3383
rect 28756 -3416 28772 -3399
rect 28534 -3433 28624 -3416
rect 28224 -3480 28624 -3433
rect 28682 -3433 28772 -3416
rect 28992 -3416 29008 -3399
rect 29214 -3399 29466 -3383
rect 29214 -3416 29230 -3399
rect 28992 -3433 29082 -3416
rect 28682 -3480 29082 -3433
rect 29140 -3433 29230 -3416
rect 29450 -3416 29466 -3399
rect 29672 -3399 29924 -3383
rect 29672 -3416 29688 -3399
rect 29450 -3433 29540 -3416
rect 29140 -3480 29540 -3433
rect 29598 -3433 29688 -3416
rect 29908 -3416 29924 -3399
rect 30130 -3399 30382 -3383
rect 30130 -3416 30146 -3399
rect 29908 -3433 29998 -3416
rect 29598 -3480 29998 -3433
rect 30056 -3433 30146 -3416
rect 30366 -3416 30382 -3399
rect 30588 -3399 30840 -3383
rect 30588 -3416 30604 -3399
rect 30366 -3433 30456 -3416
rect 30056 -3480 30456 -3433
rect 30514 -3433 30604 -3416
rect 30824 -3416 30840 -3399
rect 31046 -3399 31298 -3383
rect 31046 -3416 31062 -3399
rect 30824 -3433 30914 -3416
rect 30514 -3480 30914 -3433
rect 30972 -3433 31062 -3416
rect 31282 -3416 31298 -3399
rect 31504 -3399 31756 -3383
rect 31504 -3416 31520 -3399
rect 31282 -3433 31372 -3416
rect 30972 -3480 31372 -3433
rect 31430 -3433 31520 -3416
rect 31740 -3416 31756 -3399
rect 31962 -3399 32214 -3383
rect 31962 -3416 31978 -3399
rect 31740 -3433 31830 -3416
rect 31430 -3480 31830 -3433
rect 31888 -3433 31978 -3416
rect 32198 -3416 32214 -3399
rect 32420 -3399 32672 -3383
rect 32420 -3416 32436 -3399
rect 32198 -3433 32288 -3416
rect 31888 -3480 32288 -3433
rect 32346 -3433 32436 -3416
rect 32656 -3416 32672 -3399
rect 32878 -3399 33130 -3383
rect 32878 -3416 32894 -3399
rect 32656 -3433 32746 -3416
rect 32346 -3480 32746 -3433
rect 32804 -3433 32894 -3416
rect 33114 -3416 33130 -3399
rect 33336 -3399 33588 -3383
rect 33336 -3416 33352 -3399
rect 33114 -3433 33204 -3416
rect 32804 -3480 33204 -3433
rect 33262 -3433 33352 -3416
rect 33572 -3416 33588 -3399
rect 33794 -3399 34046 -3383
rect 33794 -3416 33810 -3399
rect 33572 -3433 33662 -3416
rect 33262 -3480 33662 -3433
rect 33720 -3433 33810 -3416
rect 34030 -3416 34046 -3399
rect 34252 -3399 34504 -3383
rect 34252 -3416 34268 -3399
rect 34030 -3433 34120 -3416
rect 33720 -3480 34120 -3433
rect 34178 -3433 34268 -3416
rect 34488 -3416 34504 -3399
rect 34710 -3399 34962 -3383
rect 34710 -3416 34726 -3399
rect 34488 -3433 34578 -3416
rect 34178 -3480 34578 -3433
rect 34636 -3433 34726 -3416
rect 34946 -3416 34962 -3399
rect 34946 -3433 35036 -3416
rect 34636 -3480 35036 -3433
rect 26850 -5127 27250 -5080
rect 26850 -5144 26940 -5127
rect 26924 -5161 26940 -5144
rect 27160 -5144 27250 -5127
rect 27308 -5127 27708 -5080
rect 27308 -5144 27398 -5127
rect 27160 -5161 27176 -5144
rect 26924 -5177 27176 -5161
rect 27382 -5161 27398 -5144
rect 27618 -5144 27708 -5127
rect 27766 -5127 28166 -5080
rect 27766 -5144 27856 -5127
rect 27618 -5161 27634 -5144
rect 27382 -5177 27634 -5161
rect 27840 -5161 27856 -5144
rect 28076 -5144 28166 -5127
rect 28224 -5127 28624 -5080
rect 28224 -5144 28314 -5127
rect 28076 -5161 28092 -5144
rect 27840 -5177 28092 -5161
rect 28298 -5161 28314 -5144
rect 28534 -5144 28624 -5127
rect 28682 -5127 29082 -5080
rect 28682 -5144 28772 -5127
rect 28534 -5161 28550 -5144
rect 28298 -5177 28550 -5161
rect 28756 -5161 28772 -5144
rect 28992 -5144 29082 -5127
rect 29140 -5127 29540 -5080
rect 29140 -5144 29230 -5127
rect 28992 -5161 29008 -5144
rect 28756 -5177 29008 -5161
rect 29214 -5161 29230 -5144
rect 29450 -5144 29540 -5127
rect 29598 -5127 29998 -5080
rect 29598 -5144 29688 -5127
rect 29450 -5161 29466 -5144
rect 29214 -5177 29466 -5161
rect 29672 -5161 29688 -5144
rect 29908 -5144 29998 -5127
rect 30056 -5127 30456 -5080
rect 30056 -5144 30146 -5127
rect 29908 -5161 29924 -5144
rect 29672 -5177 29924 -5161
rect 30130 -5161 30146 -5144
rect 30366 -5144 30456 -5127
rect 30514 -5127 30914 -5080
rect 30514 -5144 30604 -5127
rect 30366 -5161 30382 -5144
rect 30130 -5177 30382 -5161
rect 30588 -5161 30604 -5144
rect 30824 -5144 30914 -5127
rect 30972 -5127 31372 -5080
rect 30972 -5144 31062 -5127
rect 30824 -5161 30840 -5144
rect 30588 -5177 30840 -5161
rect 31046 -5161 31062 -5144
rect 31282 -5144 31372 -5127
rect 31430 -5127 31830 -5080
rect 31430 -5144 31520 -5127
rect 31282 -5161 31298 -5144
rect 31046 -5177 31298 -5161
rect 31504 -5161 31520 -5144
rect 31740 -5144 31830 -5127
rect 31888 -5127 32288 -5080
rect 31888 -5144 31978 -5127
rect 31740 -5161 31756 -5144
rect 31504 -5177 31756 -5161
rect 31962 -5161 31978 -5144
rect 32198 -5144 32288 -5127
rect 32346 -5127 32746 -5080
rect 32346 -5144 32436 -5127
rect 32198 -5161 32214 -5144
rect 31962 -5177 32214 -5161
rect 32420 -5161 32436 -5144
rect 32656 -5144 32746 -5127
rect 32804 -5127 33204 -5080
rect 32804 -5144 32894 -5127
rect 32656 -5161 32672 -5144
rect 32420 -5177 32672 -5161
rect 32878 -5161 32894 -5144
rect 33114 -5144 33204 -5127
rect 33262 -5127 33662 -5080
rect 33262 -5144 33352 -5127
rect 33114 -5161 33130 -5144
rect 32878 -5177 33130 -5161
rect 33336 -5161 33352 -5144
rect 33572 -5144 33662 -5127
rect 33720 -5127 34120 -5080
rect 33720 -5144 33810 -5127
rect 33572 -5161 33588 -5144
rect 33336 -5177 33588 -5161
rect 33794 -5161 33810 -5144
rect 34030 -5144 34120 -5127
rect 34178 -5127 34578 -5080
rect 34178 -5144 34268 -5127
rect 34030 -5161 34046 -5144
rect 33794 -5177 34046 -5161
rect 34252 -5161 34268 -5144
rect 34488 -5144 34578 -5127
rect 34636 -5127 35036 -5080
rect 34636 -5144 34726 -5127
rect 34488 -5161 34504 -5144
rect 34252 -5177 34504 -5161
rect 34710 -5161 34726 -5144
rect 34946 -5144 35036 -5127
rect 34946 -5161 34962 -5144
rect 34710 -5177 34962 -5161
rect 26365 -6064 26617 -6048
rect 26365 -6081 26381 -6064
rect 26291 -6098 26381 -6081
rect 26601 -6081 26617 -6064
rect 26823 -6064 27075 -6048
rect 26823 -6081 26839 -6064
rect 26601 -6098 26691 -6081
rect 26291 -6145 26691 -6098
rect 26749 -6098 26839 -6081
rect 27059 -6081 27075 -6064
rect 27281 -6064 27533 -6048
rect 27281 -6081 27297 -6064
rect 27059 -6098 27149 -6081
rect 26749 -6145 27149 -6098
rect 27207 -6098 27297 -6081
rect 27517 -6081 27533 -6064
rect 27739 -6064 27991 -6048
rect 27739 -6081 27755 -6064
rect 27517 -6098 27607 -6081
rect 27207 -6145 27607 -6098
rect 27665 -6098 27755 -6081
rect 27975 -6081 27991 -6064
rect 28197 -6064 28449 -6048
rect 28197 -6081 28213 -6064
rect 27975 -6098 28065 -6081
rect 27665 -6145 28065 -6098
rect 28123 -6098 28213 -6081
rect 28433 -6081 28449 -6064
rect 28655 -6064 28907 -6048
rect 28655 -6081 28671 -6064
rect 28433 -6098 28523 -6081
rect 28123 -6145 28523 -6098
rect 28581 -6098 28671 -6081
rect 28891 -6081 28907 -6064
rect 29113 -6064 29365 -6048
rect 29113 -6081 29129 -6064
rect 28891 -6098 28981 -6081
rect 28581 -6145 28981 -6098
rect 29039 -6098 29129 -6081
rect 29349 -6081 29365 -6064
rect 29571 -6064 29823 -6048
rect 29571 -6081 29587 -6064
rect 29349 -6098 29439 -6081
rect 29039 -6145 29439 -6098
rect 29497 -6098 29587 -6081
rect 29807 -6081 29823 -6064
rect 30029 -6064 30281 -6048
rect 30029 -6081 30045 -6064
rect 29807 -6098 29897 -6081
rect 29497 -6145 29897 -6098
rect 29955 -6098 30045 -6081
rect 30265 -6081 30281 -6064
rect 30487 -6064 30739 -6048
rect 30487 -6081 30503 -6064
rect 30265 -6098 30355 -6081
rect 29955 -6145 30355 -6098
rect 30413 -6098 30503 -6081
rect 30723 -6081 30739 -6064
rect 31365 -6064 31617 -6048
rect 31365 -6081 31381 -6064
rect 30723 -6098 30813 -6081
rect 30413 -6145 30813 -6098
rect 31291 -6098 31381 -6081
rect 31601 -6081 31617 -6064
rect 31823 -6064 32075 -6048
rect 31823 -6081 31839 -6064
rect 31601 -6098 31691 -6081
rect 31291 -6145 31691 -6098
rect 31749 -6098 31839 -6081
rect 32059 -6081 32075 -6064
rect 32281 -6064 32533 -6048
rect 32281 -6081 32297 -6064
rect 32059 -6098 32149 -6081
rect 31749 -6145 32149 -6098
rect 32207 -6098 32297 -6081
rect 32517 -6081 32533 -6064
rect 32739 -6064 32991 -6048
rect 32739 -6081 32755 -6064
rect 32517 -6098 32607 -6081
rect 32207 -6145 32607 -6098
rect 32665 -6098 32755 -6081
rect 32975 -6081 32991 -6064
rect 33197 -6064 33449 -6048
rect 33197 -6081 33213 -6064
rect 32975 -6098 33065 -6081
rect 32665 -6145 33065 -6098
rect 33123 -6098 33213 -6081
rect 33433 -6081 33449 -6064
rect 33655 -6064 33907 -6048
rect 33655 -6081 33671 -6064
rect 33433 -6098 33523 -6081
rect 33123 -6145 33523 -6098
rect 33581 -6098 33671 -6081
rect 33891 -6081 33907 -6064
rect 34113 -6064 34365 -6048
rect 34113 -6081 34129 -6064
rect 33891 -6098 33981 -6081
rect 33581 -6145 33981 -6098
rect 34039 -6098 34129 -6081
rect 34349 -6081 34365 -6064
rect 34571 -6064 34823 -6048
rect 34571 -6081 34587 -6064
rect 34349 -6098 34439 -6081
rect 34039 -6145 34439 -6098
rect 34497 -6098 34587 -6081
rect 34807 -6081 34823 -6064
rect 35029 -6064 35281 -6048
rect 35029 -6081 35045 -6064
rect 34807 -6098 34897 -6081
rect 34497 -6145 34897 -6098
rect 34955 -6098 35045 -6081
rect 35265 -6081 35281 -6064
rect 35487 -6064 35739 -6048
rect 35487 -6081 35503 -6064
rect 35265 -6098 35355 -6081
rect 34955 -6145 35355 -6098
rect 35413 -6098 35503 -6081
rect 35723 -6081 35739 -6064
rect 35723 -6098 35813 -6081
rect 35413 -6145 35813 -6098
rect 26291 -7392 26691 -7345
rect 26291 -7409 26381 -7392
rect 26365 -7426 26381 -7409
rect 26601 -7409 26691 -7392
rect 26749 -7392 27149 -7345
rect 26749 -7409 26839 -7392
rect 26601 -7426 26617 -7409
rect 26365 -7442 26617 -7426
rect 26823 -7426 26839 -7409
rect 27059 -7409 27149 -7392
rect 27207 -7392 27607 -7345
rect 27207 -7409 27297 -7392
rect 27059 -7426 27075 -7409
rect 26823 -7442 27075 -7426
rect 27281 -7426 27297 -7409
rect 27517 -7409 27607 -7392
rect 27665 -7392 28065 -7345
rect 27665 -7409 27755 -7392
rect 27517 -7426 27533 -7409
rect 27281 -7442 27533 -7426
rect 27739 -7426 27755 -7409
rect 27975 -7409 28065 -7392
rect 28123 -7392 28523 -7345
rect 28123 -7409 28213 -7392
rect 27975 -7426 27991 -7409
rect 27739 -7442 27991 -7426
rect 28197 -7426 28213 -7409
rect 28433 -7409 28523 -7392
rect 28581 -7392 28981 -7345
rect 28581 -7409 28671 -7392
rect 28433 -7426 28449 -7409
rect 28197 -7442 28449 -7426
rect 28655 -7426 28671 -7409
rect 28891 -7409 28981 -7392
rect 29039 -7392 29439 -7345
rect 29039 -7409 29129 -7392
rect 28891 -7426 28907 -7409
rect 28655 -7442 28907 -7426
rect 29113 -7426 29129 -7409
rect 29349 -7409 29439 -7392
rect 29497 -7392 29897 -7345
rect 29497 -7409 29587 -7392
rect 29349 -7426 29365 -7409
rect 29113 -7442 29365 -7426
rect 29571 -7426 29587 -7409
rect 29807 -7409 29897 -7392
rect 29955 -7392 30355 -7345
rect 29955 -7409 30045 -7392
rect 29807 -7426 29823 -7409
rect 29571 -7442 29823 -7426
rect 30029 -7426 30045 -7409
rect 30265 -7409 30355 -7392
rect 30413 -7392 30813 -7345
rect 30413 -7409 30503 -7392
rect 30265 -7426 30281 -7409
rect 30029 -7442 30281 -7426
rect 30487 -7426 30503 -7409
rect 30723 -7409 30813 -7392
rect 31291 -7392 31691 -7345
rect 31291 -7409 31381 -7392
rect 30723 -7426 30739 -7409
rect 30487 -7442 30739 -7426
rect 31365 -7426 31381 -7409
rect 31601 -7409 31691 -7392
rect 31749 -7392 32149 -7345
rect 31749 -7409 31839 -7392
rect 31601 -7426 31617 -7409
rect 31365 -7442 31617 -7426
rect 31823 -7426 31839 -7409
rect 32059 -7409 32149 -7392
rect 32207 -7392 32607 -7345
rect 32207 -7409 32297 -7392
rect 32059 -7426 32075 -7409
rect 31823 -7442 32075 -7426
rect 32281 -7426 32297 -7409
rect 32517 -7409 32607 -7392
rect 32665 -7392 33065 -7345
rect 32665 -7409 32755 -7392
rect 32517 -7426 32533 -7409
rect 32281 -7442 32533 -7426
rect 32739 -7426 32755 -7409
rect 32975 -7409 33065 -7392
rect 33123 -7392 33523 -7345
rect 33123 -7409 33213 -7392
rect 32975 -7426 32991 -7409
rect 32739 -7442 32991 -7426
rect 33197 -7426 33213 -7409
rect 33433 -7409 33523 -7392
rect 33581 -7392 33981 -7345
rect 33581 -7409 33671 -7392
rect 33433 -7426 33449 -7409
rect 33197 -7442 33449 -7426
rect 33655 -7426 33671 -7409
rect 33891 -7409 33981 -7392
rect 34039 -7392 34439 -7345
rect 34039 -7409 34129 -7392
rect 33891 -7426 33907 -7409
rect 33655 -7442 33907 -7426
rect 34113 -7426 34129 -7409
rect 34349 -7409 34439 -7392
rect 34497 -7392 34897 -7345
rect 34497 -7409 34587 -7392
rect 34349 -7426 34365 -7409
rect 34113 -7442 34365 -7426
rect 34571 -7426 34587 -7409
rect 34807 -7409 34897 -7392
rect 34955 -7392 35355 -7345
rect 34955 -7409 35045 -7392
rect 34807 -7426 34823 -7409
rect 34571 -7442 34823 -7426
rect 35029 -7426 35045 -7409
rect 35265 -7409 35355 -7392
rect 35413 -7392 35813 -7345
rect 35413 -7409 35503 -7392
rect 35265 -7426 35281 -7409
rect 35029 -7442 35281 -7426
rect 35487 -7426 35503 -7409
rect 35723 -7409 35813 -7392
rect 35723 -7426 35739 -7409
rect 35487 -7442 35739 -7426
rect 11364 -8566 11616 -8550
rect 11364 -8583 11380 -8566
rect 11290 -8600 11380 -8583
rect 11600 -8583 11616 -8566
rect 11822 -8566 12074 -8550
rect 11822 -8583 11838 -8566
rect 11600 -8600 11690 -8583
rect 11290 -8638 11690 -8600
rect 11748 -8600 11838 -8583
rect 12058 -8583 12074 -8566
rect 12280 -8566 12532 -8550
rect 12280 -8583 12296 -8566
rect 12058 -8600 12148 -8583
rect 11748 -8638 12148 -8600
rect 12206 -8600 12296 -8583
rect 12516 -8583 12532 -8566
rect 12738 -8566 12990 -8550
rect 12738 -8583 12754 -8566
rect 12516 -8600 12606 -8583
rect 12206 -8638 12606 -8600
rect 12664 -8600 12754 -8583
rect 12974 -8583 12990 -8566
rect 13196 -8566 13448 -8550
rect 13196 -8583 13212 -8566
rect 12974 -8600 13064 -8583
rect 12664 -8638 13064 -8600
rect 13122 -8600 13212 -8583
rect 13432 -8583 13448 -8566
rect 13654 -8566 13906 -8550
rect 13654 -8583 13670 -8566
rect 13432 -8600 13522 -8583
rect 13122 -8638 13522 -8600
rect 13580 -8600 13670 -8583
rect 13890 -8583 13906 -8566
rect 14112 -8566 14364 -8550
rect 14112 -8583 14128 -8566
rect 13890 -8600 13980 -8583
rect 13580 -8638 13980 -8600
rect 14038 -8600 14128 -8583
rect 14348 -8583 14364 -8566
rect 14570 -8566 14822 -8550
rect 14570 -8583 14586 -8566
rect 14348 -8600 14438 -8583
rect 14038 -8638 14438 -8600
rect 14496 -8600 14586 -8583
rect 14806 -8583 14822 -8566
rect 15028 -8566 15280 -8550
rect 15028 -8583 15044 -8566
rect 14806 -8600 14896 -8583
rect 14496 -8638 14896 -8600
rect 14954 -8600 15044 -8583
rect 15264 -8583 15280 -8566
rect 15486 -8566 15738 -8550
rect 15486 -8583 15502 -8566
rect 15264 -8600 15354 -8583
rect 14954 -8638 15354 -8600
rect 15412 -8600 15502 -8583
rect 15722 -8583 15738 -8566
rect 16364 -8566 16616 -8550
rect 16364 -8583 16380 -8566
rect 15722 -8600 15812 -8583
rect 15412 -8638 15812 -8600
rect 16290 -8600 16380 -8583
rect 16600 -8583 16616 -8566
rect 16822 -8566 17074 -8550
rect 16822 -8583 16838 -8566
rect 16600 -8600 16690 -8583
rect 16290 -8638 16690 -8600
rect 16748 -8600 16838 -8583
rect 17058 -8583 17074 -8566
rect 17280 -8566 17532 -8550
rect 17280 -8583 17296 -8566
rect 17058 -8600 17148 -8583
rect 16748 -8638 17148 -8600
rect 17206 -8600 17296 -8583
rect 17516 -8583 17532 -8566
rect 17738 -8566 17990 -8550
rect 17738 -8583 17754 -8566
rect 17516 -8600 17606 -8583
rect 17206 -8638 17606 -8600
rect 17664 -8600 17754 -8583
rect 17974 -8583 17990 -8566
rect 18196 -8566 18448 -8550
rect 18196 -8583 18212 -8566
rect 17974 -8600 18064 -8583
rect 17664 -8638 18064 -8600
rect 18122 -8600 18212 -8583
rect 18432 -8583 18448 -8566
rect 18654 -8566 18906 -8550
rect 18654 -8583 18670 -8566
rect 18432 -8600 18522 -8583
rect 18122 -8638 18522 -8600
rect 18580 -8600 18670 -8583
rect 18890 -8583 18906 -8566
rect 19112 -8566 19364 -8550
rect 19112 -8583 19128 -8566
rect 18890 -8600 18980 -8583
rect 18580 -8638 18980 -8600
rect 19038 -8600 19128 -8583
rect 19348 -8583 19364 -8566
rect 19570 -8566 19822 -8550
rect 19570 -8583 19586 -8566
rect 19348 -8600 19438 -8583
rect 19038 -8638 19438 -8600
rect 19496 -8600 19586 -8583
rect 19806 -8583 19822 -8566
rect 20028 -8566 20280 -8550
rect 20028 -8583 20044 -8566
rect 19806 -8600 19896 -8583
rect 19496 -8638 19896 -8600
rect 19954 -8600 20044 -8583
rect 20264 -8583 20280 -8566
rect 20486 -8566 20738 -8550
rect 20486 -8583 20502 -8566
rect 20264 -8600 20354 -8583
rect 19954 -8638 20354 -8600
rect 20412 -8600 20502 -8583
rect 20722 -8583 20738 -8566
rect 20722 -8600 20812 -8583
rect 20412 -8638 20812 -8600
rect 11290 -8876 11690 -8838
rect 11290 -8893 11380 -8876
rect 11364 -8910 11380 -8893
rect 11600 -8893 11690 -8876
rect 11748 -8876 12148 -8838
rect 11748 -8893 11838 -8876
rect 11600 -8910 11616 -8893
rect 11364 -8926 11616 -8910
rect 11822 -8910 11838 -8893
rect 12058 -8893 12148 -8876
rect 12206 -8876 12606 -8838
rect 12206 -8893 12296 -8876
rect 12058 -8910 12074 -8893
rect 11822 -8926 12074 -8910
rect 12280 -8910 12296 -8893
rect 12516 -8893 12606 -8876
rect 12664 -8876 13064 -8838
rect 12664 -8893 12754 -8876
rect 12516 -8910 12532 -8893
rect 12280 -8926 12532 -8910
rect 12738 -8910 12754 -8893
rect 12974 -8893 13064 -8876
rect 13122 -8876 13522 -8838
rect 13122 -8893 13212 -8876
rect 12974 -8910 12990 -8893
rect 12738 -8926 12990 -8910
rect 13196 -8910 13212 -8893
rect 13432 -8893 13522 -8876
rect 13580 -8876 13980 -8838
rect 13580 -8893 13670 -8876
rect 13432 -8910 13448 -8893
rect 13196 -8926 13448 -8910
rect 13654 -8910 13670 -8893
rect 13890 -8893 13980 -8876
rect 14038 -8876 14438 -8838
rect 14038 -8893 14128 -8876
rect 13890 -8910 13906 -8893
rect 13654 -8926 13906 -8910
rect 14112 -8910 14128 -8893
rect 14348 -8893 14438 -8876
rect 14496 -8876 14896 -8838
rect 14496 -8893 14586 -8876
rect 14348 -8910 14364 -8893
rect 14112 -8926 14364 -8910
rect 14570 -8910 14586 -8893
rect 14806 -8893 14896 -8876
rect 14954 -8876 15354 -8838
rect 14954 -8893 15044 -8876
rect 14806 -8910 14822 -8893
rect 14570 -8926 14822 -8910
rect 15028 -8910 15044 -8893
rect 15264 -8893 15354 -8876
rect 15412 -8876 15812 -8838
rect 15412 -8893 15502 -8876
rect 15264 -8910 15280 -8893
rect 15028 -8926 15280 -8910
rect 15486 -8910 15502 -8893
rect 15722 -8893 15812 -8876
rect 16290 -8876 16690 -8838
rect 16290 -8893 16380 -8876
rect 15722 -8910 15738 -8893
rect 15486 -8926 15738 -8910
rect 16364 -8910 16380 -8893
rect 16600 -8893 16690 -8876
rect 16748 -8876 17148 -8838
rect 16748 -8893 16838 -8876
rect 16600 -8910 16616 -8893
rect 16364 -8926 16616 -8910
rect 16822 -8910 16838 -8893
rect 17058 -8893 17148 -8876
rect 17206 -8876 17606 -8838
rect 17206 -8893 17296 -8876
rect 17058 -8910 17074 -8893
rect 16822 -8926 17074 -8910
rect 17280 -8910 17296 -8893
rect 17516 -8893 17606 -8876
rect 17664 -8876 18064 -8838
rect 17664 -8893 17754 -8876
rect 17516 -8910 17532 -8893
rect 17280 -8926 17532 -8910
rect 17738 -8910 17754 -8893
rect 17974 -8893 18064 -8876
rect 18122 -8876 18522 -8838
rect 18122 -8893 18212 -8876
rect 17974 -8910 17990 -8893
rect 17738 -8926 17990 -8910
rect 18196 -8910 18212 -8893
rect 18432 -8893 18522 -8876
rect 18580 -8876 18980 -8838
rect 18580 -8893 18670 -8876
rect 18432 -8910 18448 -8893
rect 18196 -8926 18448 -8910
rect 18654 -8910 18670 -8893
rect 18890 -8893 18980 -8876
rect 19038 -8876 19438 -8838
rect 19038 -8893 19128 -8876
rect 18890 -8910 18906 -8893
rect 18654 -8926 18906 -8910
rect 19112 -8910 19128 -8893
rect 19348 -8893 19438 -8876
rect 19496 -8876 19896 -8838
rect 19496 -8893 19586 -8876
rect 19348 -8910 19364 -8893
rect 19112 -8926 19364 -8910
rect 19570 -8910 19586 -8893
rect 19806 -8893 19896 -8876
rect 19954 -8876 20354 -8838
rect 19954 -8893 20044 -8876
rect 19806 -8910 19822 -8893
rect 19570 -8926 19822 -8910
rect 20028 -8910 20044 -8893
rect 20264 -8893 20354 -8876
rect 20412 -8876 20812 -8838
rect 20412 -8893 20502 -8876
rect 20264 -8910 20280 -8893
rect 20028 -8926 20280 -8910
rect 20486 -8910 20502 -8893
rect 20722 -8893 20812 -8876
rect 20722 -8910 20738 -8893
rect 20486 -8926 20738 -8910
rect 11364 -9234 11616 -9218
rect 11364 -9251 11380 -9234
rect 11290 -9268 11380 -9251
rect 11600 -9251 11616 -9234
rect 11822 -9234 12074 -9218
rect 11822 -9251 11838 -9234
rect 11600 -9268 11690 -9251
rect 11290 -9306 11690 -9268
rect 11748 -9268 11838 -9251
rect 12058 -9251 12074 -9234
rect 12280 -9234 12532 -9218
rect 12280 -9251 12296 -9234
rect 12058 -9268 12148 -9251
rect 11748 -9306 12148 -9268
rect 12206 -9268 12296 -9251
rect 12516 -9251 12532 -9234
rect 12738 -9234 12990 -9218
rect 12738 -9251 12754 -9234
rect 12516 -9268 12606 -9251
rect 12206 -9306 12606 -9268
rect 12664 -9268 12754 -9251
rect 12974 -9251 12990 -9234
rect 13196 -9234 13448 -9218
rect 13196 -9251 13212 -9234
rect 12974 -9268 13064 -9251
rect 12664 -9306 13064 -9268
rect 13122 -9268 13212 -9251
rect 13432 -9251 13448 -9234
rect 13654 -9234 13906 -9218
rect 13654 -9251 13670 -9234
rect 13432 -9268 13522 -9251
rect 13122 -9306 13522 -9268
rect 13580 -9268 13670 -9251
rect 13890 -9251 13906 -9234
rect 14112 -9234 14364 -9218
rect 14112 -9251 14128 -9234
rect 13890 -9268 13980 -9251
rect 13580 -9306 13980 -9268
rect 14038 -9268 14128 -9251
rect 14348 -9251 14364 -9234
rect 14570 -9234 14822 -9218
rect 14570 -9251 14586 -9234
rect 14348 -9268 14438 -9251
rect 14038 -9306 14438 -9268
rect 14496 -9268 14586 -9251
rect 14806 -9251 14822 -9234
rect 15028 -9234 15280 -9218
rect 15028 -9251 15044 -9234
rect 14806 -9268 14896 -9251
rect 14496 -9306 14896 -9268
rect 14954 -9268 15044 -9251
rect 15264 -9251 15280 -9234
rect 15486 -9234 15738 -9218
rect 15486 -9251 15502 -9234
rect 15264 -9268 15354 -9251
rect 14954 -9306 15354 -9268
rect 15412 -9268 15502 -9251
rect 15722 -9251 15738 -9234
rect 15722 -9268 15812 -9251
rect 15412 -9306 15812 -9268
rect 11290 -9544 11690 -9506
rect 11290 -9561 11380 -9544
rect 11364 -9578 11380 -9561
rect 11600 -9561 11690 -9544
rect 11748 -9544 12148 -9506
rect 11748 -9561 11838 -9544
rect 11600 -9578 11616 -9561
rect 11364 -9594 11616 -9578
rect 11822 -9578 11838 -9561
rect 12058 -9561 12148 -9544
rect 12206 -9544 12606 -9506
rect 12206 -9561 12296 -9544
rect 12058 -9578 12074 -9561
rect 11822 -9594 12074 -9578
rect 12280 -9578 12296 -9561
rect 12516 -9561 12606 -9544
rect 12664 -9544 13064 -9506
rect 12664 -9561 12754 -9544
rect 12516 -9578 12532 -9561
rect 12280 -9594 12532 -9578
rect 12738 -9578 12754 -9561
rect 12974 -9561 13064 -9544
rect 13122 -9544 13522 -9506
rect 13122 -9561 13212 -9544
rect 12974 -9578 12990 -9561
rect 12738 -9594 12990 -9578
rect 13196 -9578 13212 -9561
rect 13432 -9561 13522 -9544
rect 13580 -9544 13980 -9506
rect 13580 -9561 13670 -9544
rect 13432 -9578 13448 -9561
rect 13196 -9594 13448 -9578
rect 13654 -9578 13670 -9561
rect 13890 -9561 13980 -9544
rect 14038 -9544 14438 -9506
rect 14038 -9561 14128 -9544
rect 13890 -9578 13906 -9561
rect 13654 -9594 13906 -9578
rect 14112 -9578 14128 -9561
rect 14348 -9561 14438 -9544
rect 14496 -9544 14896 -9506
rect 14496 -9561 14586 -9544
rect 14348 -9578 14364 -9561
rect 14112 -9594 14364 -9578
rect 14570 -9578 14586 -9561
rect 14806 -9561 14896 -9544
rect 14954 -9544 15354 -9506
rect 14954 -9561 15044 -9544
rect 14806 -9578 14822 -9561
rect 14570 -9594 14822 -9578
rect 15028 -9578 15044 -9561
rect 15264 -9561 15354 -9544
rect 15412 -9544 15812 -9506
rect 15412 -9561 15502 -9544
rect 15264 -9578 15280 -9561
rect 15028 -9594 15280 -9578
rect 15486 -9578 15502 -9561
rect 15722 -9561 15812 -9544
rect 15722 -9578 15738 -9561
rect 15486 -9594 15738 -9578
rect 26364 -8566 26616 -8550
rect 26364 -8583 26380 -8566
rect 26290 -8600 26380 -8583
rect 26600 -8583 26616 -8566
rect 26822 -8566 27074 -8550
rect 26822 -8583 26838 -8566
rect 26600 -8600 26690 -8583
rect 26290 -8638 26690 -8600
rect 26748 -8600 26838 -8583
rect 27058 -8583 27074 -8566
rect 27280 -8566 27532 -8550
rect 27280 -8583 27296 -8566
rect 27058 -8600 27148 -8583
rect 26748 -8638 27148 -8600
rect 27206 -8600 27296 -8583
rect 27516 -8583 27532 -8566
rect 27738 -8566 27990 -8550
rect 27738 -8583 27754 -8566
rect 27516 -8600 27606 -8583
rect 27206 -8638 27606 -8600
rect 27664 -8600 27754 -8583
rect 27974 -8583 27990 -8566
rect 28196 -8566 28448 -8550
rect 28196 -8583 28212 -8566
rect 27974 -8600 28064 -8583
rect 27664 -8638 28064 -8600
rect 28122 -8600 28212 -8583
rect 28432 -8583 28448 -8566
rect 28654 -8566 28906 -8550
rect 28654 -8583 28670 -8566
rect 28432 -8600 28522 -8583
rect 28122 -8638 28522 -8600
rect 28580 -8600 28670 -8583
rect 28890 -8583 28906 -8566
rect 29112 -8566 29364 -8550
rect 29112 -8583 29128 -8566
rect 28890 -8600 28980 -8583
rect 28580 -8638 28980 -8600
rect 29038 -8600 29128 -8583
rect 29348 -8583 29364 -8566
rect 29570 -8566 29822 -8550
rect 29570 -8583 29586 -8566
rect 29348 -8600 29438 -8583
rect 29038 -8638 29438 -8600
rect 29496 -8600 29586 -8583
rect 29806 -8583 29822 -8566
rect 30028 -8566 30280 -8550
rect 30028 -8583 30044 -8566
rect 29806 -8600 29896 -8583
rect 29496 -8638 29896 -8600
rect 29954 -8600 30044 -8583
rect 30264 -8583 30280 -8566
rect 30486 -8566 30738 -8550
rect 30486 -8583 30502 -8566
rect 30264 -8600 30354 -8583
rect 29954 -8638 30354 -8600
rect 30412 -8600 30502 -8583
rect 30722 -8583 30738 -8566
rect 31364 -8566 31616 -8550
rect 31364 -8583 31380 -8566
rect 30722 -8600 30812 -8583
rect 30412 -8638 30812 -8600
rect 31290 -8600 31380 -8583
rect 31600 -8583 31616 -8566
rect 31822 -8566 32074 -8550
rect 31822 -8583 31838 -8566
rect 31600 -8600 31690 -8583
rect 31290 -8638 31690 -8600
rect 31748 -8600 31838 -8583
rect 32058 -8583 32074 -8566
rect 32280 -8566 32532 -8550
rect 32280 -8583 32296 -8566
rect 32058 -8600 32148 -8583
rect 31748 -8638 32148 -8600
rect 32206 -8600 32296 -8583
rect 32516 -8583 32532 -8566
rect 32738 -8566 32990 -8550
rect 32738 -8583 32754 -8566
rect 32516 -8600 32606 -8583
rect 32206 -8638 32606 -8600
rect 32664 -8600 32754 -8583
rect 32974 -8583 32990 -8566
rect 33196 -8566 33448 -8550
rect 33196 -8583 33212 -8566
rect 32974 -8600 33064 -8583
rect 32664 -8638 33064 -8600
rect 33122 -8600 33212 -8583
rect 33432 -8583 33448 -8566
rect 33654 -8566 33906 -8550
rect 33654 -8583 33670 -8566
rect 33432 -8600 33522 -8583
rect 33122 -8638 33522 -8600
rect 33580 -8600 33670 -8583
rect 33890 -8583 33906 -8566
rect 34112 -8566 34364 -8550
rect 34112 -8583 34128 -8566
rect 33890 -8600 33980 -8583
rect 33580 -8638 33980 -8600
rect 34038 -8600 34128 -8583
rect 34348 -8583 34364 -8566
rect 34570 -8566 34822 -8550
rect 34570 -8583 34586 -8566
rect 34348 -8600 34438 -8583
rect 34038 -8638 34438 -8600
rect 34496 -8600 34586 -8583
rect 34806 -8583 34822 -8566
rect 35028 -8566 35280 -8550
rect 35028 -8583 35044 -8566
rect 34806 -8600 34896 -8583
rect 34496 -8638 34896 -8600
rect 34954 -8600 35044 -8583
rect 35264 -8583 35280 -8566
rect 35486 -8566 35738 -8550
rect 35486 -8583 35502 -8566
rect 35264 -8600 35354 -8583
rect 34954 -8638 35354 -8600
rect 35412 -8600 35502 -8583
rect 35722 -8583 35738 -8566
rect 35722 -8600 35812 -8583
rect 35412 -8638 35812 -8600
rect 26290 -8876 26690 -8838
rect 26290 -8893 26380 -8876
rect 26364 -8910 26380 -8893
rect 26600 -8893 26690 -8876
rect 26748 -8876 27148 -8838
rect 26748 -8893 26838 -8876
rect 26600 -8910 26616 -8893
rect 26364 -8926 26616 -8910
rect 26822 -8910 26838 -8893
rect 27058 -8893 27148 -8876
rect 27206 -8876 27606 -8838
rect 27206 -8893 27296 -8876
rect 27058 -8910 27074 -8893
rect 26822 -8926 27074 -8910
rect 27280 -8910 27296 -8893
rect 27516 -8893 27606 -8876
rect 27664 -8876 28064 -8838
rect 27664 -8893 27754 -8876
rect 27516 -8910 27532 -8893
rect 27280 -8926 27532 -8910
rect 27738 -8910 27754 -8893
rect 27974 -8893 28064 -8876
rect 28122 -8876 28522 -8838
rect 28122 -8893 28212 -8876
rect 27974 -8910 27990 -8893
rect 27738 -8926 27990 -8910
rect 28196 -8910 28212 -8893
rect 28432 -8893 28522 -8876
rect 28580 -8876 28980 -8838
rect 28580 -8893 28670 -8876
rect 28432 -8910 28448 -8893
rect 28196 -8926 28448 -8910
rect 28654 -8910 28670 -8893
rect 28890 -8893 28980 -8876
rect 29038 -8876 29438 -8838
rect 29038 -8893 29128 -8876
rect 28890 -8910 28906 -8893
rect 28654 -8926 28906 -8910
rect 29112 -8910 29128 -8893
rect 29348 -8893 29438 -8876
rect 29496 -8876 29896 -8838
rect 29496 -8893 29586 -8876
rect 29348 -8910 29364 -8893
rect 29112 -8926 29364 -8910
rect 29570 -8910 29586 -8893
rect 29806 -8893 29896 -8876
rect 29954 -8876 30354 -8838
rect 29954 -8893 30044 -8876
rect 29806 -8910 29822 -8893
rect 29570 -8926 29822 -8910
rect 30028 -8910 30044 -8893
rect 30264 -8893 30354 -8876
rect 30412 -8876 30812 -8838
rect 30412 -8893 30502 -8876
rect 30264 -8910 30280 -8893
rect 30028 -8926 30280 -8910
rect 30486 -8910 30502 -8893
rect 30722 -8893 30812 -8876
rect 31290 -8876 31690 -8838
rect 31290 -8893 31380 -8876
rect 30722 -8910 30738 -8893
rect 30486 -8926 30738 -8910
rect 31364 -8910 31380 -8893
rect 31600 -8893 31690 -8876
rect 31748 -8876 32148 -8838
rect 31748 -8893 31838 -8876
rect 31600 -8910 31616 -8893
rect 31364 -8926 31616 -8910
rect 31822 -8910 31838 -8893
rect 32058 -8893 32148 -8876
rect 32206 -8876 32606 -8838
rect 32206 -8893 32296 -8876
rect 32058 -8910 32074 -8893
rect 31822 -8926 32074 -8910
rect 32280 -8910 32296 -8893
rect 32516 -8893 32606 -8876
rect 32664 -8876 33064 -8838
rect 32664 -8893 32754 -8876
rect 32516 -8910 32532 -8893
rect 32280 -8926 32532 -8910
rect 32738 -8910 32754 -8893
rect 32974 -8893 33064 -8876
rect 33122 -8876 33522 -8838
rect 33122 -8893 33212 -8876
rect 32974 -8910 32990 -8893
rect 32738 -8926 32990 -8910
rect 33196 -8910 33212 -8893
rect 33432 -8893 33522 -8876
rect 33580 -8876 33980 -8838
rect 33580 -8893 33670 -8876
rect 33432 -8910 33448 -8893
rect 33196 -8926 33448 -8910
rect 33654 -8910 33670 -8893
rect 33890 -8893 33980 -8876
rect 34038 -8876 34438 -8838
rect 34038 -8893 34128 -8876
rect 33890 -8910 33906 -8893
rect 33654 -8926 33906 -8910
rect 34112 -8910 34128 -8893
rect 34348 -8893 34438 -8876
rect 34496 -8876 34896 -8838
rect 34496 -8893 34586 -8876
rect 34348 -8910 34364 -8893
rect 34112 -8926 34364 -8910
rect 34570 -8910 34586 -8893
rect 34806 -8893 34896 -8876
rect 34954 -8876 35354 -8838
rect 34954 -8893 35044 -8876
rect 34806 -8910 34822 -8893
rect 34570 -8926 34822 -8910
rect 35028 -8910 35044 -8893
rect 35264 -8893 35354 -8876
rect 35412 -8876 35812 -8838
rect 35412 -8893 35502 -8876
rect 35264 -8910 35280 -8893
rect 35028 -8926 35280 -8910
rect 35486 -8910 35502 -8893
rect 35722 -8893 35812 -8876
rect 35722 -8910 35738 -8893
rect 35486 -8926 35738 -8910
rect 26364 -9234 26616 -9218
rect 26364 -9251 26380 -9234
rect 26290 -9268 26380 -9251
rect 26600 -9251 26616 -9234
rect 26822 -9234 27074 -9218
rect 26822 -9251 26838 -9234
rect 26600 -9268 26690 -9251
rect 26290 -9306 26690 -9268
rect 26748 -9268 26838 -9251
rect 27058 -9251 27074 -9234
rect 27280 -9234 27532 -9218
rect 27280 -9251 27296 -9234
rect 27058 -9268 27148 -9251
rect 26748 -9306 27148 -9268
rect 27206 -9268 27296 -9251
rect 27516 -9251 27532 -9234
rect 27738 -9234 27990 -9218
rect 27738 -9251 27754 -9234
rect 27516 -9268 27606 -9251
rect 27206 -9306 27606 -9268
rect 27664 -9268 27754 -9251
rect 27974 -9251 27990 -9234
rect 28196 -9234 28448 -9218
rect 28196 -9251 28212 -9234
rect 27974 -9268 28064 -9251
rect 27664 -9306 28064 -9268
rect 28122 -9268 28212 -9251
rect 28432 -9251 28448 -9234
rect 28654 -9234 28906 -9218
rect 28654 -9251 28670 -9234
rect 28432 -9268 28522 -9251
rect 28122 -9306 28522 -9268
rect 28580 -9268 28670 -9251
rect 28890 -9251 28906 -9234
rect 29112 -9234 29364 -9218
rect 29112 -9251 29128 -9234
rect 28890 -9268 28980 -9251
rect 28580 -9306 28980 -9268
rect 29038 -9268 29128 -9251
rect 29348 -9251 29364 -9234
rect 29570 -9234 29822 -9218
rect 29570 -9251 29586 -9234
rect 29348 -9268 29438 -9251
rect 29038 -9306 29438 -9268
rect 29496 -9268 29586 -9251
rect 29806 -9251 29822 -9234
rect 30028 -9234 30280 -9218
rect 30028 -9251 30044 -9234
rect 29806 -9268 29896 -9251
rect 29496 -9306 29896 -9268
rect 29954 -9268 30044 -9251
rect 30264 -9251 30280 -9234
rect 30486 -9234 30738 -9218
rect 30486 -9251 30502 -9234
rect 30264 -9268 30354 -9251
rect 29954 -9306 30354 -9268
rect 30412 -9268 30502 -9251
rect 30722 -9251 30738 -9234
rect 30722 -9268 30812 -9251
rect 30412 -9306 30812 -9268
rect 26290 -9544 26690 -9506
rect 26290 -9561 26380 -9544
rect 26364 -9578 26380 -9561
rect 26600 -9561 26690 -9544
rect 26748 -9544 27148 -9506
rect 26748 -9561 26838 -9544
rect 26600 -9578 26616 -9561
rect 26364 -9594 26616 -9578
rect 26822 -9578 26838 -9561
rect 27058 -9561 27148 -9544
rect 27206 -9544 27606 -9506
rect 27206 -9561 27296 -9544
rect 27058 -9578 27074 -9561
rect 26822 -9594 27074 -9578
rect 27280 -9578 27296 -9561
rect 27516 -9561 27606 -9544
rect 27664 -9544 28064 -9506
rect 27664 -9561 27754 -9544
rect 27516 -9578 27532 -9561
rect 27280 -9594 27532 -9578
rect 27738 -9578 27754 -9561
rect 27974 -9561 28064 -9544
rect 28122 -9544 28522 -9506
rect 28122 -9561 28212 -9544
rect 27974 -9578 27990 -9561
rect 27738 -9594 27990 -9578
rect 28196 -9578 28212 -9561
rect 28432 -9561 28522 -9544
rect 28580 -9544 28980 -9506
rect 28580 -9561 28670 -9544
rect 28432 -9578 28448 -9561
rect 28196 -9594 28448 -9578
rect 28654 -9578 28670 -9561
rect 28890 -9561 28980 -9544
rect 29038 -9544 29438 -9506
rect 29038 -9561 29128 -9544
rect 28890 -9578 28906 -9561
rect 28654 -9594 28906 -9578
rect 29112 -9578 29128 -9561
rect 29348 -9561 29438 -9544
rect 29496 -9544 29896 -9506
rect 29496 -9561 29586 -9544
rect 29348 -9578 29364 -9561
rect 29112 -9594 29364 -9578
rect 29570 -9578 29586 -9561
rect 29806 -9561 29896 -9544
rect 29954 -9544 30354 -9506
rect 29954 -9561 30044 -9544
rect 29806 -9578 29822 -9561
rect 29570 -9594 29822 -9578
rect 30028 -9578 30044 -9561
rect 30264 -9561 30354 -9544
rect 30412 -9544 30812 -9506
rect 30412 -9561 30502 -9544
rect 30264 -9578 30280 -9561
rect 30028 -9594 30280 -9578
rect 30486 -9578 30502 -9561
rect 30722 -9561 30812 -9544
rect 30722 -9578 30738 -9561
rect 30486 -9594 30738 -9578
rect 20296 -12026 20548 -12010
rect 20296 -12043 20312 -12026
rect 20222 -12060 20312 -12043
rect 20532 -12043 20548 -12026
rect 20754 -12026 21006 -12010
rect 20754 -12043 20770 -12026
rect 20532 -12060 20622 -12043
rect 20222 -12098 20622 -12060
rect 20680 -12060 20770 -12043
rect 20990 -12043 21006 -12026
rect 21212 -12026 21464 -12010
rect 21212 -12043 21228 -12026
rect 20990 -12060 21080 -12043
rect 20680 -12098 21080 -12060
rect 21138 -12060 21228 -12043
rect 21448 -12043 21464 -12026
rect 21670 -12026 21922 -12010
rect 21670 -12043 21686 -12026
rect 21448 -12060 21538 -12043
rect 21138 -12098 21538 -12060
rect 21596 -12060 21686 -12043
rect 21906 -12043 21922 -12026
rect 22128 -12026 22380 -12010
rect 22128 -12043 22144 -12026
rect 21906 -12060 21996 -12043
rect 21596 -12098 21996 -12060
rect 22054 -12060 22144 -12043
rect 22364 -12043 22380 -12026
rect 22586 -12026 22838 -12010
rect 22586 -12043 22602 -12026
rect 22364 -12060 22454 -12043
rect 22054 -12098 22454 -12060
rect 22512 -12060 22602 -12043
rect 22822 -12043 22838 -12026
rect 23044 -12026 23296 -12010
rect 23044 -12043 23060 -12026
rect 22822 -12060 22912 -12043
rect 22512 -12098 22912 -12060
rect 22970 -12060 23060 -12043
rect 23280 -12043 23296 -12026
rect 23502 -12026 23754 -12010
rect 23502 -12043 23518 -12026
rect 23280 -12060 23370 -12043
rect 22970 -12098 23370 -12060
rect 23428 -12060 23518 -12043
rect 23738 -12043 23754 -12026
rect 23960 -12026 24212 -12010
rect 23960 -12043 23976 -12026
rect 23738 -12060 23828 -12043
rect 23428 -12098 23828 -12060
rect 23886 -12060 23976 -12043
rect 24196 -12043 24212 -12026
rect 24418 -12026 24670 -12010
rect 24418 -12043 24434 -12026
rect 24196 -12060 24286 -12043
rect 23886 -12098 24286 -12060
rect 24344 -12060 24434 -12043
rect 24654 -12043 24670 -12026
rect 24654 -12060 24744 -12043
rect 24344 -12098 24744 -12060
rect 20222 -12336 20622 -12298
rect 20222 -12353 20312 -12336
rect 20296 -12370 20312 -12353
rect 20532 -12353 20622 -12336
rect 20680 -12336 21080 -12298
rect 20680 -12353 20770 -12336
rect 20532 -12370 20548 -12353
rect 20296 -12386 20548 -12370
rect 20754 -12370 20770 -12353
rect 20990 -12353 21080 -12336
rect 21138 -12336 21538 -12298
rect 21138 -12353 21228 -12336
rect 20990 -12370 21006 -12353
rect 20754 -12386 21006 -12370
rect 21212 -12370 21228 -12353
rect 21448 -12353 21538 -12336
rect 21596 -12336 21996 -12298
rect 21596 -12353 21686 -12336
rect 21448 -12370 21464 -12353
rect 21212 -12386 21464 -12370
rect 21670 -12370 21686 -12353
rect 21906 -12353 21996 -12336
rect 22054 -12336 22454 -12298
rect 22054 -12353 22144 -12336
rect 21906 -12370 21922 -12353
rect 21670 -12386 21922 -12370
rect 22128 -12370 22144 -12353
rect 22364 -12353 22454 -12336
rect 22512 -12336 22912 -12298
rect 22512 -12353 22602 -12336
rect 22364 -12370 22380 -12353
rect 22128 -12386 22380 -12370
rect 22586 -12370 22602 -12353
rect 22822 -12353 22912 -12336
rect 22970 -12336 23370 -12298
rect 22970 -12353 23060 -12336
rect 22822 -12370 22838 -12353
rect 22586 -12386 22838 -12370
rect 23044 -12370 23060 -12353
rect 23280 -12353 23370 -12336
rect 23428 -12336 23828 -12298
rect 23428 -12353 23518 -12336
rect 23280 -12370 23296 -12353
rect 23044 -12386 23296 -12370
rect 23502 -12370 23518 -12353
rect 23738 -12353 23828 -12336
rect 23886 -12336 24286 -12298
rect 23886 -12353 23976 -12336
rect 23738 -12370 23754 -12353
rect 23502 -12386 23754 -12370
rect 23960 -12370 23976 -12353
rect 24196 -12353 24286 -12336
rect 24344 -12336 24744 -12298
rect 24344 -12353 24434 -12336
rect 24196 -12370 24212 -12353
rect 23960 -12386 24212 -12370
rect 24418 -12370 24434 -12353
rect 24654 -12353 24744 -12336
rect 24654 -12370 24670 -12353
rect 24418 -12386 24670 -12370
rect 15296 -12694 15548 -12678
rect 15296 -12711 15312 -12694
rect 15222 -12728 15312 -12711
rect 15532 -12711 15548 -12694
rect 15754 -12694 16006 -12678
rect 15754 -12711 15770 -12694
rect 15532 -12728 15622 -12711
rect 15222 -12766 15622 -12728
rect 15680 -12728 15770 -12711
rect 15990 -12711 16006 -12694
rect 16212 -12694 16464 -12678
rect 16212 -12711 16228 -12694
rect 15990 -12728 16080 -12711
rect 15680 -12766 16080 -12728
rect 16138 -12728 16228 -12711
rect 16448 -12711 16464 -12694
rect 16670 -12694 16922 -12678
rect 16670 -12711 16686 -12694
rect 16448 -12728 16538 -12711
rect 16138 -12766 16538 -12728
rect 16596 -12728 16686 -12711
rect 16906 -12711 16922 -12694
rect 17128 -12694 17380 -12678
rect 17128 -12711 17144 -12694
rect 16906 -12728 16996 -12711
rect 16596 -12766 16996 -12728
rect 17054 -12728 17144 -12711
rect 17364 -12711 17380 -12694
rect 17586 -12694 17838 -12678
rect 17586 -12711 17602 -12694
rect 17364 -12728 17454 -12711
rect 17054 -12766 17454 -12728
rect 17512 -12728 17602 -12711
rect 17822 -12711 17838 -12694
rect 18044 -12694 18296 -12678
rect 18044 -12711 18060 -12694
rect 17822 -12728 17912 -12711
rect 17512 -12766 17912 -12728
rect 17970 -12728 18060 -12711
rect 18280 -12711 18296 -12694
rect 18502 -12694 18754 -12678
rect 18502 -12711 18518 -12694
rect 18280 -12728 18370 -12711
rect 17970 -12766 18370 -12728
rect 18428 -12728 18518 -12711
rect 18738 -12711 18754 -12694
rect 18960 -12694 19212 -12678
rect 18960 -12711 18976 -12694
rect 18738 -12728 18828 -12711
rect 18428 -12766 18828 -12728
rect 18886 -12728 18976 -12711
rect 19196 -12711 19212 -12694
rect 19418 -12694 19670 -12678
rect 19418 -12711 19434 -12694
rect 19196 -12728 19286 -12711
rect 18886 -12766 19286 -12728
rect 19344 -12728 19434 -12711
rect 19654 -12711 19670 -12694
rect 20296 -12694 20548 -12678
rect 20296 -12711 20312 -12694
rect 19654 -12728 19744 -12711
rect 19344 -12766 19744 -12728
rect 20222 -12728 20312 -12711
rect 20532 -12711 20548 -12694
rect 20754 -12694 21006 -12678
rect 20754 -12711 20770 -12694
rect 20532 -12728 20622 -12711
rect 20222 -12766 20622 -12728
rect 20680 -12728 20770 -12711
rect 20990 -12711 21006 -12694
rect 21212 -12694 21464 -12678
rect 21212 -12711 21228 -12694
rect 20990 -12728 21080 -12711
rect 20680 -12766 21080 -12728
rect 21138 -12728 21228 -12711
rect 21448 -12711 21464 -12694
rect 21670 -12694 21922 -12678
rect 21670 -12711 21686 -12694
rect 21448 -12728 21538 -12711
rect 21138 -12766 21538 -12728
rect 21596 -12728 21686 -12711
rect 21906 -12711 21922 -12694
rect 22128 -12694 22380 -12678
rect 22128 -12711 22144 -12694
rect 21906 -12728 21996 -12711
rect 21596 -12766 21996 -12728
rect 22054 -12728 22144 -12711
rect 22364 -12711 22380 -12694
rect 22586 -12694 22838 -12678
rect 22586 -12711 22602 -12694
rect 22364 -12728 22454 -12711
rect 22054 -12766 22454 -12728
rect 22512 -12728 22602 -12711
rect 22822 -12711 22838 -12694
rect 23044 -12694 23296 -12678
rect 23044 -12711 23060 -12694
rect 22822 -12728 22912 -12711
rect 22512 -12766 22912 -12728
rect 22970 -12728 23060 -12711
rect 23280 -12711 23296 -12694
rect 23502 -12694 23754 -12678
rect 23502 -12711 23518 -12694
rect 23280 -12728 23370 -12711
rect 22970 -12766 23370 -12728
rect 23428 -12728 23518 -12711
rect 23738 -12711 23754 -12694
rect 23960 -12694 24212 -12678
rect 23960 -12711 23976 -12694
rect 23738 -12728 23828 -12711
rect 23428 -12766 23828 -12728
rect 23886 -12728 23976 -12711
rect 24196 -12711 24212 -12694
rect 24418 -12694 24670 -12678
rect 24418 -12711 24434 -12694
rect 24196 -12728 24286 -12711
rect 23886 -12766 24286 -12728
rect 24344 -12728 24434 -12711
rect 24654 -12711 24670 -12694
rect 24654 -12728 24744 -12711
rect 24344 -12766 24744 -12728
rect 15222 -13004 15622 -12966
rect 15222 -13021 15312 -13004
rect 15296 -13038 15312 -13021
rect 15532 -13021 15622 -13004
rect 15680 -13004 16080 -12966
rect 15680 -13021 15770 -13004
rect 15532 -13038 15548 -13021
rect 15296 -13054 15548 -13038
rect 15754 -13038 15770 -13021
rect 15990 -13021 16080 -13004
rect 16138 -13004 16538 -12966
rect 16138 -13021 16228 -13004
rect 15990 -13038 16006 -13021
rect 15754 -13054 16006 -13038
rect 16212 -13038 16228 -13021
rect 16448 -13021 16538 -13004
rect 16596 -13004 16996 -12966
rect 16596 -13021 16686 -13004
rect 16448 -13038 16464 -13021
rect 16212 -13054 16464 -13038
rect 16670 -13038 16686 -13021
rect 16906 -13021 16996 -13004
rect 17054 -13004 17454 -12966
rect 17054 -13021 17144 -13004
rect 16906 -13038 16922 -13021
rect 16670 -13054 16922 -13038
rect 17128 -13038 17144 -13021
rect 17364 -13021 17454 -13004
rect 17512 -13004 17912 -12966
rect 17512 -13021 17602 -13004
rect 17364 -13038 17380 -13021
rect 17128 -13054 17380 -13038
rect 17586 -13038 17602 -13021
rect 17822 -13021 17912 -13004
rect 17970 -13004 18370 -12966
rect 17970 -13021 18060 -13004
rect 17822 -13038 17838 -13021
rect 17586 -13054 17838 -13038
rect 18044 -13038 18060 -13021
rect 18280 -13021 18370 -13004
rect 18428 -13004 18828 -12966
rect 18428 -13021 18518 -13004
rect 18280 -13038 18296 -13021
rect 18044 -13054 18296 -13038
rect 18502 -13038 18518 -13021
rect 18738 -13021 18828 -13004
rect 18886 -13004 19286 -12966
rect 18886 -13021 18976 -13004
rect 18738 -13038 18754 -13021
rect 18502 -13054 18754 -13038
rect 18960 -13038 18976 -13021
rect 19196 -13021 19286 -13004
rect 19344 -13004 19744 -12966
rect 19344 -13021 19434 -13004
rect 19196 -13038 19212 -13021
rect 18960 -13054 19212 -13038
rect 19418 -13038 19434 -13021
rect 19654 -13021 19744 -13004
rect 20222 -13004 20622 -12966
rect 20222 -13021 20312 -13004
rect 19654 -13038 19670 -13021
rect 19418 -13054 19670 -13038
rect 20296 -13038 20312 -13021
rect 20532 -13021 20622 -13004
rect 20680 -13004 21080 -12966
rect 20680 -13021 20770 -13004
rect 20532 -13038 20548 -13021
rect 20296 -13054 20548 -13038
rect 20754 -13038 20770 -13021
rect 20990 -13021 21080 -13004
rect 21138 -13004 21538 -12966
rect 21138 -13021 21228 -13004
rect 20990 -13038 21006 -13021
rect 20754 -13054 21006 -13038
rect 21212 -13038 21228 -13021
rect 21448 -13021 21538 -13004
rect 21596 -13004 21996 -12966
rect 21596 -13021 21686 -13004
rect 21448 -13038 21464 -13021
rect 21212 -13054 21464 -13038
rect 21670 -13038 21686 -13021
rect 21906 -13021 21996 -13004
rect 22054 -13004 22454 -12966
rect 22054 -13021 22144 -13004
rect 21906 -13038 21922 -13021
rect 21670 -13054 21922 -13038
rect 22128 -13038 22144 -13021
rect 22364 -13021 22454 -13004
rect 22512 -13004 22912 -12966
rect 22512 -13021 22602 -13004
rect 22364 -13038 22380 -13021
rect 22128 -13054 22380 -13038
rect 22586 -13038 22602 -13021
rect 22822 -13021 22912 -13004
rect 22970 -13004 23370 -12966
rect 22970 -13021 23060 -13004
rect 22822 -13038 22838 -13021
rect 22586 -13054 22838 -13038
rect 23044 -13038 23060 -13021
rect 23280 -13021 23370 -13004
rect 23428 -13004 23828 -12966
rect 23428 -13021 23518 -13004
rect 23280 -13038 23296 -13021
rect 23044 -13054 23296 -13038
rect 23502 -13038 23518 -13021
rect 23738 -13021 23828 -13004
rect 23886 -13004 24286 -12966
rect 23886 -13021 23976 -13004
rect 23738 -13038 23754 -13021
rect 23502 -13054 23754 -13038
rect 23960 -13038 23976 -13021
rect 24196 -13021 24286 -13004
rect 24344 -13004 24744 -12966
rect 24344 -13021 24434 -13004
rect 24196 -13038 24212 -13021
rect 23960 -13054 24212 -13038
rect 24418 -13038 24434 -13021
rect 24654 -13021 24744 -13004
rect 24654 -13038 24670 -13021
rect 24418 -13054 24670 -13038
rect 35296 -12026 35548 -12010
rect 35296 -12043 35312 -12026
rect 35222 -12060 35312 -12043
rect 35532 -12043 35548 -12026
rect 35754 -12026 36006 -12010
rect 35754 -12043 35770 -12026
rect 35532 -12060 35622 -12043
rect 35222 -12098 35622 -12060
rect 35680 -12060 35770 -12043
rect 35990 -12043 36006 -12026
rect 36212 -12026 36464 -12010
rect 36212 -12043 36228 -12026
rect 35990 -12060 36080 -12043
rect 35680 -12098 36080 -12060
rect 36138 -12060 36228 -12043
rect 36448 -12043 36464 -12026
rect 36670 -12026 36922 -12010
rect 36670 -12043 36686 -12026
rect 36448 -12060 36538 -12043
rect 36138 -12098 36538 -12060
rect 36596 -12060 36686 -12043
rect 36906 -12043 36922 -12026
rect 37128 -12026 37380 -12010
rect 37128 -12043 37144 -12026
rect 36906 -12060 36996 -12043
rect 36596 -12098 36996 -12060
rect 37054 -12060 37144 -12043
rect 37364 -12043 37380 -12026
rect 37586 -12026 37838 -12010
rect 37586 -12043 37602 -12026
rect 37364 -12060 37454 -12043
rect 37054 -12098 37454 -12060
rect 37512 -12060 37602 -12043
rect 37822 -12043 37838 -12026
rect 38044 -12026 38296 -12010
rect 38044 -12043 38060 -12026
rect 37822 -12060 37912 -12043
rect 37512 -12098 37912 -12060
rect 37970 -12060 38060 -12043
rect 38280 -12043 38296 -12026
rect 38502 -12026 38754 -12010
rect 38502 -12043 38518 -12026
rect 38280 -12060 38370 -12043
rect 37970 -12098 38370 -12060
rect 38428 -12060 38518 -12043
rect 38738 -12043 38754 -12026
rect 38960 -12026 39212 -12010
rect 38960 -12043 38976 -12026
rect 38738 -12060 38828 -12043
rect 38428 -12098 38828 -12060
rect 38886 -12060 38976 -12043
rect 39196 -12043 39212 -12026
rect 39418 -12026 39670 -12010
rect 39418 -12043 39434 -12026
rect 39196 -12060 39286 -12043
rect 38886 -12098 39286 -12060
rect 39344 -12060 39434 -12043
rect 39654 -12043 39670 -12026
rect 39654 -12060 39744 -12043
rect 39344 -12098 39744 -12060
rect 35222 -12336 35622 -12298
rect 35222 -12353 35312 -12336
rect 35296 -12370 35312 -12353
rect 35532 -12353 35622 -12336
rect 35680 -12336 36080 -12298
rect 35680 -12353 35770 -12336
rect 35532 -12370 35548 -12353
rect 35296 -12386 35548 -12370
rect 35754 -12370 35770 -12353
rect 35990 -12353 36080 -12336
rect 36138 -12336 36538 -12298
rect 36138 -12353 36228 -12336
rect 35990 -12370 36006 -12353
rect 35754 -12386 36006 -12370
rect 36212 -12370 36228 -12353
rect 36448 -12353 36538 -12336
rect 36596 -12336 36996 -12298
rect 36596 -12353 36686 -12336
rect 36448 -12370 36464 -12353
rect 36212 -12386 36464 -12370
rect 36670 -12370 36686 -12353
rect 36906 -12353 36996 -12336
rect 37054 -12336 37454 -12298
rect 37054 -12353 37144 -12336
rect 36906 -12370 36922 -12353
rect 36670 -12386 36922 -12370
rect 37128 -12370 37144 -12353
rect 37364 -12353 37454 -12336
rect 37512 -12336 37912 -12298
rect 37512 -12353 37602 -12336
rect 37364 -12370 37380 -12353
rect 37128 -12386 37380 -12370
rect 37586 -12370 37602 -12353
rect 37822 -12353 37912 -12336
rect 37970 -12336 38370 -12298
rect 37970 -12353 38060 -12336
rect 37822 -12370 37838 -12353
rect 37586 -12386 37838 -12370
rect 38044 -12370 38060 -12353
rect 38280 -12353 38370 -12336
rect 38428 -12336 38828 -12298
rect 38428 -12353 38518 -12336
rect 38280 -12370 38296 -12353
rect 38044 -12386 38296 -12370
rect 38502 -12370 38518 -12353
rect 38738 -12353 38828 -12336
rect 38886 -12336 39286 -12298
rect 38886 -12353 38976 -12336
rect 38738 -12370 38754 -12353
rect 38502 -12386 38754 -12370
rect 38960 -12370 38976 -12353
rect 39196 -12353 39286 -12336
rect 39344 -12336 39744 -12298
rect 39344 -12353 39434 -12336
rect 39196 -12370 39212 -12353
rect 38960 -12386 39212 -12370
rect 39418 -12370 39434 -12353
rect 39654 -12353 39744 -12336
rect 39654 -12370 39670 -12353
rect 39418 -12386 39670 -12370
rect 30296 -12694 30548 -12678
rect 30296 -12711 30312 -12694
rect 30222 -12728 30312 -12711
rect 30532 -12711 30548 -12694
rect 30754 -12694 31006 -12678
rect 30754 -12711 30770 -12694
rect 30532 -12728 30622 -12711
rect 30222 -12766 30622 -12728
rect 30680 -12728 30770 -12711
rect 30990 -12711 31006 -12694
rect 31212 -12694 31464 -12678
rect 31212 -12711 31228 -12694
rect 30990 -12728 31080 -12711
rect 30680 -12766 31080 -12728
rect 31138 -12728 31228 -12711
rect 31448 -12711 31464 -12694
rect 31670 -12694 31922 -12678
rect 31670 -12711 31686 -12694
rect 31448 -12728 31538 -12711
rect 31138 -12766 31538 -12728
rect 31596 -12728 31686 -12711
rect 31906 -12711 31922 -12694
rect 32128 -12694 32380 -12678
rect 32128 -12711 32144 -12694
rect 31906 -12728 31996 -12711
rect 31596 -12766 31996 -12728
rect 32054 -12728 32144 -12711
rect 32364 -12711 32380 -12694
rect 32586 -12694 32838 -12678
rect 32586 -12711 32602 -12694
rect 32364 -12728 32454 -12711
rect 32054 -12766 32454 -12728
rect 32512 -12728 32602 -12711
rect 32822 -12711 32838 -12694
rect 33044 -12694 33296 -12678
rect 33044 -12711 33060 -12694
rect 32822 -12728 32912 -12711
rect 32512 -12766 32912 -12728
rect 32970 -12728 33060 -12711
rect 33280 -12711 33296 -12694
rect 33502 -12694 33754 -12678
rect 33502 -12711 33518 -12694
rect 33280 -12728 33370 -12711
rect 32970 -12766 33370 -12728
rect 33428 -12728 33518 -12711
rect 33738 -12711 33754 -12694
rect 33960 -12694 34212 -12678
rect 33960 -12711 33976 -12694
rect 33738 -12728 33828 -12711
rect 33428 -12766 33828 -12728
rect 33886 -12728 33976 -12711
rect 34196 -12711 34212 -12694
rect 34418 -12694 34670 -12678
rect 34418 -12711 34434 -12694
rect 34196 -12728 34286 -12711
rect 33886 -12766 34286 -12728
rect 34344 -12728 34434 -12711
rect 34654 -12711 34670 -12694
rect 35296 -12694 35548 -12678
rect 35296 -12711 35312 -12694
rect 34654 -12728 34744 -12711
rect 34344 -12766 34744 -12728
rect 35222 -12728 35312 -12711
rect 35532 -12711 35548 -12694
rect 35754 -12694 36006 -12678
rect 35754 -12711 35770 -12694
rect 35532 -12728 35622 -12711
rect 35222 -12766 35622 -12728
rect 35680 -12728 35770 -12711
rect 35990 -12711 36006 -12694
rect 36212 -12694 36464 -12678
rect 36212 -12711 36228 -12694
rect 35990 -12728 36080 -12711
rect 35680 -12766 36080 -12728
rect 36138 -12728 36228 -12711
rect 36448 -12711 36464 -12694
rect 36670 -12694 36922 -12678
rect 36670 -12711 36686 -12694
rect 36448 -12728 36538 -12711
rect 36138 -12766 36538 -12728
rect 36596 -12728 36686 -12711
rect 36906 -12711 36922 -12694
rect 37128 -12694 37380 -12678
rect 37128 -12711 37144 -12694
rect 36906 -12728 36996 -12711
rect 36596 -12766 36996 -12728
rect 37054 -12728 37144 -12711
rect 37364 -12711 37380 -12694
rect 37586 -12694 37838 -12678
rect 37586 -12711 37602 -12694
rect 37364 -12728 37454 -12711
rect 37054 -12766 37454 -12728
rect 37512 -12728 37602 -12711
rect 37822 -12711 37838 -12694
rect 38044 -12694 38296 -12678
rect 38044 -12711 38060 -12694
rect 37822 -12728 37912 -12711
rect 37512 -12766 37912 -12728
rect 37970 -12728 38060 -12711
rect 38280 -12711 38296 -12694
rect 38502 -12694 38754 -12678
rect 38502 -12711 38518 -12694
rect 38280 -12728 38370 -12711
rect 37970 -12766 38370 -12728
rect 38428 -12728 38518 -12711
rect 38738 -12711 38754 -12694
rect 38960 -12694 39212 -12678
rect 38960 -12711 38976 -12694
rect 38738 -12728 38828 -12711
rect 38428 -12766 38828 -12728
rect 38886 -12728 38976 -12711
rect 39196 -12711 39212 -12694
rect 39418 -12694 39670 -12678
rect 39418 -12711 39434 -12694
rect 39196 -12728 39286 -12711
rect 38886 -12766 39286 -12728
rect 39344 -12728 39434 -12711
rect 39654 -12711 39670 -12694
rect 39654 -12728 39744 -12711
rect 39344 -12766 39744 -12728
rect 30222 -13004 30622 -12966
rect 30222 -13021 30312 -13004
rect 30296 -13038 30312 -13021
rect 30532 -13021 30622 -13004
rect 30680 -13004 31080 -12966
rect 30680 -13021 30770 -13004
rect 30532 -13038 30548 -13021
rect 30296 -13054 30548 -13038
rect 30754 -13038 30770 -13021
rect 30990 -13021 31080 -13004
rect 31138 -13004 31538 -12966
rect 31138 -13021 31228 -13004
rect 30990 -13038 31006 -13021
rect 30754 -13054 31006 -13038
rect 31212 -13038 31228 -13021
rect 31448 -13021 31538 -13004
rect 31596 -13004 31996 -12966
rect 31596 -13021 31686 -13004
rect 31448 -13038 31464 -13021
rect 31212 -13054 31464 -13038
rect 31670 -13038 31686 -13021
rect 31906 -13021 31996 -13004
rect 32054 -13004 32454 -12966
rect 32054 -13021 32144 -13004
rect 31906 -13038 31922 -13021
rect 31670 -13054 31922 -13038
rect 32128 -13038 32144 -13021
rect 32364 -13021 32454 -13004
rect 32512 -13004 32912 -12966
rect 32512 -13021 32602 -13004
rect 32364 -13038 32380 -13021
rect 32128 -13054 32380 -13038
rect 32586 -13038 32602 -13021
rect 32822 -13021 32912 -13004
rect 32970 -13004 33370 -12966
rect 32970 -13021 33060 -13004
rect 32822 -13038 32838 -13021
rect 32586 -13054 32838 -13038
rect 33044 -13038 33060 -13021
rect 33280 -13021 33370 -13004
rect 33428 -13004 33828 -12966
rect 33428 -13021 33518 -13004
rect 33280 -13038 33296 -13021
rect 33044 -13054 33296 -13038
rect 33502 -13038 33518 -13021
rect 33738 -13021 33828 -13004
rect 33886 -13004 34286 -12966
rect 33886 -13021 33976 -13004
rect 33738 -13038 33754 -13021
rect 33502 -13054 33754 -13038
rect 33960 -13038 33976 -13021
rect 34196 -13021 34286 -13004
rect 34344 -13004 34744 -12966
rect 34344 -13021 34434 -13004
rect 34196 -13038 34212 -13021
rect 33960 -13054 34212 -13038
rect 34418 -13038 34434 -13021
rect 34654 -13021 34744 -13004
rect 35222 -13004 35622 -12966
rect 35222 -13021 35312 -13004
rect 34654 -13038 34670 -13021
rect 34418 -13054 34670 -13038
rect 35296 -13038 35312 -13021
rect 35532 -13021 35622 -13004
rect 35680 -13004 36080 -12966
rect 35680 -13021 35770 -13004
rect 35532 -13038 35548 -13021
rect 35296 -13054 35548 -13038
rect 35754 -13038 35770 -13021
rect 35990 -13021 36080 -13004
rect 36138 -13004 36538 -12966
rect 36138 -13021 36228 -13004
rect 35990 -13038 36006 -13021
rect 35754 -13054 36006 -13038
rect 36212 -13038 36228 -13021
rect 36448 -13021 36538 -13004
rect 36596 -13004 36996 -12966
rect 36596 -13021 36686 -13004
rect 36448 -13038 36464 -13021
rect 36212 -13054 36464 -13038
rect 36670 -13038 36686 -13021
rect 36906 -13021 36996 -13004
rect 37054 -13004 37454 -12966
rect 37054 -13021 37144 -13004
rect 36906 -13038 36922 -13021
rect 36670 -13054 36922 -13038
rect 37128 -13038 37144 -13021
rect 37364 -13021 37454 -13004
rect 37512 -13004 37912 -12966
rect 37512 -13021 37602 -13004
rect 37364 -13038 37380 -13021
rect 37128 -13054 37380 -13038
rect 37586 -13038 37602 -13021
rect 37822 -13021 37912 -13004
rect 37970 -13004 38370 -12966
rect 37970 -13021 38060 -13004
rect 37822 -13038 37838 -13021
rect 37586 -13054 37838 -13038
rect 38044 -13038 38060 -13021
rect 38280 -13021 38370 -13004
rect 38428 -13004 38828 -12966
rect 38428 -13021 38518 -13004
rect 38280 -13038 38296 -13021
rect 38044 -13054 38296 -13038
rect 38502 -13038 38518 -13021
rect 38738 -13021 38828 -13004
rect 38886 -13004 39286 -12966
rect 38886 -13021 38976 -13004
rect 38738 -13038 38754 -13021
rect 38502 -13054 38754 -13038
rect 38960 -13038 38976 -13021
rect 39196 -13021 39286 -13004
rect 39344 -13004 39744 -12966
rect 39344 -13021 39434 -13004
rect 39196 -13038 39212 -13021
rect 38960 -13054 39212 -13038
rect 39418 -13038 39434 -13021
rect 39654 -13021 39744 -13004
rect 39654 -13038 39670 -13021
rect 39418 -13054 39670 -13038
rect 15295 -14178 15547 -14162
rect 15295 -14195 15311 -14178
rect 15221 -14212 15311 -14195
rect 15531 -14195 15547 -14178
rect 15753 -14178 16005 -14162
rect 15753 -14195 15769 -14178
rect 15531 -14212 15621 -14195
rect 15221 -14259 15621 -14212
rect 15679 -14212 15769 -14195
rect 15989 -14195 16005 -14178
rect 16211 -14178 16463 -14162
rect 16211 -14195 16227 -14178
rect 15989 -14212 16079 -14195
rect 15679 -14259 16079 -14212
rect 16137 -14212 16227 -14195
rect 16447 -14195 16463 -14178
rect 16669 -14178 16921 -14162
rect 16669 -14195 16685 -14178
rect 16447 -14212 16537 -14195
rect 16137 -14259 16537 -14212
rect 16595 -14212 16685 -14195
rect 16905 -14195 16921 -14178
rect 17127 -14178 17379 -14162
rect 17127 -14195 17143 -14178
rect 16905 -14212 16995 -14195
rect 16595 -14259 16995 -14212
rect 17053 -14212 17143 -14195
rect 17363 -14195 17379 -14178
rect 17585 -14178 17837 -14162
rect 17585 -14195 17601 -14178
rect 17363 -14212 17453 -14195
rect 17053 -14259 17453 -14212
rect 17511 -14212 17601 -14195
rect 17821 -14195 17837 -14178
rect 18043 -14178 18295 -14162
rect 18043 -14195 18059 -14178
rect 17821 -14212 17911 -14195
rect 17511 -14259 17911 -14212
rect 17969 -14212 18059 -14195
rect 18279 -14195 18295 -14178
rect 18501 -14178 18753 -14162
rect 18501 -14195 18517 -14178
rect 18279 -14212 18369 -14195
rect 17969 -14259 18369 -14212
rect 18427 -14212 18517 -14195
rect 18737 -14195 18753 -14178
rect 18959 -14178 19211 -14162
rect 18959 -14195 18975 -14178
rect 18737 -14212 18827 -14195
rect 18427 -14259 18827 -14212
rect 18885 -14212 18975 -14195
rect 19195 -14195 19211 -14178
rect 19417 -14178 19669 -14162
rect 19417 -14195 19433 -14178
rect 19195 -14212 19285 -14195
rect 18885 -14259 19285 -14212
rect 19343 -14212 19433 -14195
rect 19653 -14195 19669 -14178
rect 20295 -14178 20547 -14162
rect 20295 -14195 20311 -14178
rect 19653 -14212 19743 -14195
rect 19343 -14259 19743 -14212
rect 20221 -14212 20311 -14195
rect 20531 -14195 20547 -14178
rect 20753 -14178 21005 -14162
rect 20753 -14195 20769 -14178
rect 20531 -14212 20621 -14195
rect 20221 -14259 20621 -14212
rect 20679 -14212 20769 -14195
rect 20989 -14195 21005 -14178
rect 21211 -14178 21463 -14162
rect 21211 -14195 21227 -14178
rect 20989 -14212 21079 -14195
rect 20679 -14259 21079 -14212
rect 21137 -14212 21227 -14195
rect 21447 -14195 21463 -14178
rect 21669 -14178 21921 -14162
rect 21669 -14195 21685 -14178
rect 21447 -14212 21537 -14195
rect 21137 -14259 21537 -14212
rect 21595 -14212 21685 -14195
rect 21905 -14195 21921 -14178
rect 22127 -14178 22379 -14162
rect 22127 -14195 22143 -14178
rect 21905 -14212 21995 -14195
rect 21595 -14259 21995 -14212
rect 22053 -14212 22143 -14195
rect 22363 -14195 22379 -14178
rect 22585 -14178 22837 -14162
rect 22585 -14195 22601 -14178
rect 22363 -14212 22453 -14195
rect 22053 -14259 22453 -14212
rect 22511 -14212 22601 -14195
rect 22821 -14195 22837 -14178
rect 23043 -14178 23295 -14162
rect 23043 -14195 23059 -14178
rect 22821 -14212 22911 -14195
rect 22511 -14259 22911 -14212
rect 22969 -14212 23059 -14195
rect 23279 -14195 23295 -14178
rect 23501 -14178 23753 -14162
rect 23501 -14195 23517 -14178
rect 23279 -14212 23369 -14195
rect 22969 -14259 23369 -14212
rect 23427 -14212 23517 -14195
rect 23737 -14195 23753 -14178
rect 23959 -14178 24211 -14162
rect 23959 -14195 23975 -14178
rect 23737 -14212 23827 -14195
rect 23427 -14259 23827 -14212
rect 23885 -14212 23975 -14195
rect 24195 -14195 24211 -14178
rect 24417 -14178 24669 -14162
rect 24417 -14195 24433 -14178
rect 24195 -14212 24285 -14195
rect 23885 -14259 24285 -14212
rect 24343 -14212 24433 -14195
rect 24653 -14195 24669 -14178
rect 24653 -14212 24743 -14195
rect 24343 -14259 24743 -14212
rect 15221 -15506 15621 -15459
rect 15221 -15523 15311 -15506
rect 15295 -15540 15311 -15523
rect 15531 -15523 15621 -15506
rect 15679 -15506 16079 -15459
rect 15679 -15523 15769 -15506
rect 15531 -15540 15547 -15523
rect 15295 -15556 15547 -15540
rect 15753 -15540 15769 -15523
rect 15989 -15523 16079 -15506
rect 16137 -15506 16537 -15459
rect 16137 -15523 16227 -15506
rect 15989 -15540 16005 -15523
rect 15753 -15556 16005 -15540
rect 16211 -15540 16227 -15523
rect 16447 -15523 16537 -15506
rect 16595 -15506 16995 -15459
rect 16595 -15523 16685 -15506
rect 16447 -15540 16463 -15523
rect 16211 -15556 16463 -15540
rect 16669 -15540 16685 -15523
rect 16905 -15523 16995 -15506
rect 17053 -15506 17453 -15459
rect 17053 -15523 17143 -15506
rect 16905 -15540 16921 -15523
rect 16669 -15556 16921 -15540
rect 17127 -15540 17143 -15523
rect 17363 -15523 17453 -15506
rect 17511 -15506 17911 -15459
rect 17511 -15523 17601 -15506
rect 17363 -15540 17379 -15523
rect 17127 -15556 17379 -15540
rect 17585 -15540 17601 -15523
rect 17821 -15523 17911 -15506
rect 17969 -15506 18369 -15459
rect 17969 -15523 18059 -15506
rect 17821 -15540 17837 -15523
rect 17585 -15556 17837 -15540
rect 18043 -15540 18059 -15523
rect 18279 -15523 18369 -15506
rect 18427 -15506 18827 -15459
rect 18427 -15523 18517 -15506
rect 18279 -15540 18295 -15523
rect 18043 -15556 18295 -15540
rect 18501 -15540 18517 -15523
rect 18737 -15523 18827 -15506
rect 18885 -15506 19285 -15459
rect 18885 -15523 18975 -15506
rect 18737 -15540 18753 -15523
rect 18501 -15556 18753 -15540
rect 18959 -15540 18975 -15523
rect 19195 -15523 19285 -15506
rect 19343 -15506 19743 -15459
rect 19343 -15523 19433 -15506
rect 19195 -15540 19211 -15523
rect 18959 -15556 19211 -15540
rect 19417 -15540 19433 -15523
rect 19653 -15523 19743 -15506
rect 20221 -15506 20621 -15459
rect 20221 -15523 20311 -15506
rect 19653 -15540 19669 -15523
rect 19417 -15556 19669 -15540
rect 20295 -15540 20311 -15523
rect 20531 -15523 20621 -15506
rect 20679 -15506 21079 -15459
rect 20679 -15523 20769 -15506
rect 20531 -15540 20547 -15523
rect 20295 -15556 20547 -15540
rect 20753 -15540 20769 -15523
rect 20989 -15523 21079 -15506
rect 21137 -15506 21537 -15459
rect 21137 -15523 21227 -15506
rect 20989 -15540 21005 -15523
rect 20753 -15556 21005 -15540
rect 21211 -15540 21227 -15523
rect 21447 -15523 21537 -15506
rect 21595 -15506 21995 -15459
rect 21595 -15523 21685 -15506
rect 21447 -15540 21463 -15523
rect 21211 -15556 21463 -15540
rect 21669 -15540 21685 -15523
rect 21905 -15523 21995 -15506
rect 22053 -15506 22453 -15459
rect 22053 -15523 22143 -15506
rect 21905 -15540 21921 -15523
rect 21669 -15556 21921 -15540
rect 22127 -15540 22143 -15523
rect 22363 -15523 22453 -15506
rect 22511 -15506 22911 -15459
rect 22511 -15523 22601 -15506
rect 22363 -15540 22379 -15523
rect 22127 -15556 22379 -15540
rect 22585 -15540 22601 -15523
rect 22821 -15523 22911 -15506
rect 22969 -15506 23369 -15459
rect 22969 -15523 23059 -15506
rect 22821 -15540 22837 -15523
rect 22585 -15556 22837 -15540
rect 23043 -15540 23059 -15523
rect 23279 -15523 23369 -15506
rect 23427 -15506 23827 -15459
rect 23427 -15523 23517 -15506
rect 23279 -15540 23295 -15523
rect 23043 -15556 23295 -15540
rect 23501 -15540 23517 -15523
rect 23737 -15523 23827 -15506
rect 23885 -15506 24285 -15459
rect 23885 -15523 23975 -15506
rect 23737 -15540 23753 -15523
rect 23501 -15556 23753 -15540
rect 23959 -15540 23975 -15523
rect 24195 -15523 24285 -15506
rect 24343 -15506 24743 -15459
rect 24343 -15523 24433 -15506
rect 24195 -15540 24211 -15523
rect 23959 -15556 24211 -15540
rect 24417 -15540 24433 -15523
rect 24653 -15523 24743 -15506
rect 24653 -15540 24669 -15523
rect 24417 -15556 24669 -15540
rect 16072 -16443 16324 -16427
rect 16072 -16460 16088 -16443
rect 15998 -16477 16088 -16460
rect 16308 -16460 16324 -16443
rect 16530 -16443 16782 -16427
rect 16530 -16460 16546 -16443
rect 16308 -16477 16398 -16460
rect 15998 -16524 16398 -16477
rect 16456 -16477 16546 -16460
rect 16766 -16460 16782 -16443
rect 16988 -16443 17240 -16427
rect 16988 -16460 17004 -16443
rect 16766 -16477 16856 -16460
rect 16456 -16524 16856 -16477
rect 16914 -16477 17004 -16460
rect 17224 -16460 17240 -16443
rect 17446 -16443 17698 -16427
rect 17446 -16460 17462 -16443
rect 17224 -16477 17314 -16460
rect 16914 -16524 17314 -16477
rect 17372 -16477 17462 -16460
rect 17682 -16460 17698 -16443
rect 17904 -16443 18156 -16427
rect 17904 -16460 17920 -16443
rect 17682 -16477 17772 -16460
rect 17372 -16524 17772 -16477
rect 17830 -16477 17920 -16460
rect 18140 -16460 18156 -16443
rect 18362 -16443 18614 -16427
rect 18362 -16460 18378 -16443
rect 18140 -16477 18230 -16460
rect 17830 -16524 18230 -16477
rect 18288 -16477 18378 -16460
rect 18598 -16460 18614 -16443
rect 18820 -16443 19072 -16427
rect 18820 -16460 18836 -16443
rect 18598 -16477 18688 -16460
rect 18288 -16524 18688 -16477
rect 18746 -16477 18836 -16460
rect 19056 -16460 19072 -16443
rect 19278 -16443 19530 -16427
rect 19278 -16460 19294 -16443
rect 19056 -16477 19146 -16460
rect 18746 -16524 19146 -16477
rect 19204 -16477 19294 -16460
rect 19514 -16460 19530 -16443
rect 19736 -16443 19988 -16427
rect 19736 -16460 19752 -16443
rect 19514 -16477 19604 -16460
rect 19204 -16524 19604 -16477
rect 19662 -16477 19752 -16460
rect 19972 -16460 19988 -16443
rect 20194 -16443 20446 -16427
rect 20194 -16460 20210 -16443
rect 19972 -16477 20062 -16460
rect 19662 -16524 20062 -16477
rect 20120 -16477 20210 -16460
rect 20430 -16460 20446 -16443
rect 20652 -16443 20904 -16427
rect 20652 -16460 20668 -16443
rect 20430 -16477 20520 -16460
rect 20120 -16524 20520 -16477
rect 20578 -16477 20668 -16460
rect 20888 -16460 20904 -16443
rect 21110 -16443 21362 -16427
rect 21110 -16460 21126 -16443
rect 20888 -16477 20978 -16460
rect 20578 -16524 20978 -16477
rect 21036 -16477 21126 -16460
rect 21346 -16460 21362 -16443
rect 21568 -16443 21820 -16427
rect 21568 -16460 21584 -16443
rect 21346 -16477 21436 -16460
rect 21036 -16524 21436 -16477
rect 21494 -16477 21584 -16460
rect 21804 -16460 21820 -16443
rect 22026 -16443 22278 -16427
rect 22026 -16460 22042 -16443
rect 21804 -16477 21894 -16460
rect 21494 -16524 21894 -16477
rect 21952 -16477 22042 -16460
rect 22262 -16460 22278 -16443
rect 22484 -16443 22736 -16427
rect 22484 -16460 22500 -16443
rect 22262 -16477 22352 -16460
rect 21952 -16524 22352 -16477
rect 22410 -16477 22500 -16460
rect 22720 -16460 22736 -16443
rect 22942 -16443 23194 -16427
rect 22942 -16460 22958 -16443
rect 22720 -16477 22810 -16460
rect 22410 -16524 22810 -16477
rect 22868 -16477 22958 -16460
rect 23178 -16460 23194 -16443
rect 23400 -16443 23652 -16427
rect 23400 -16460 23416 -16443
rect 23178 -16477 23268 -16460
rect 22868 -16524 23268 -16477
rect 23326 -16477 23416 -16460
rect 23636 -16460 23652 -16443
rect 23858 -16443 24110 -16427
rect 23858 -16460 23874 -16443
rect 23636 -16477 23726 -16460
rect 23326 -16524 23726 -16477
rect 23784 -16477 23874 -16460
rect 24094 -16460 24110 -16443
rect 24094 -16477 24184 -16460
rect 23784 -16524 24184 -16477
rect 15998 -18171 16398 -18124
rect 15998 -18188 16088 -18171
rect 16072 -18205 16088 -18188
rect 16308 -18188 16398 -18171
rect 16456 -18171 16856 -18124
rect 16456 -18188 16546 -18171
rect 16308 -18205 16324 -18188
rect 16072 -18221 16324 -18205
rect 16530 -18205 16546 -18188
rect 16766 -18188 16856 -18171
rect 16914 -18171 17314 -18124
rect 16914 -18188 17004 -18171
rect 16766 -18205 16782 -18188
rect 16530 -18221 16782 -18205
rect 16988 -18205 17004 -18188
rect 17224 -18188 17314 -18171
rect 17372 -18171 17772 -18124
rect 17372 -18188 17462 -18171
rect 17224 -18205 17240 -18188
rect 16988 -18221 17240 -18205
rect 17446 -18205 17462 -18188
rect 17682 -18188 17772 -18171
rect 17830 -18171 18230 -18124
rect 17830 -18188 17920 -18171
rect 17682 -18205 17698 -18188
rect 17446 -18221 17698 -18205
rect 17904 -18205 17920 -18188
rect 18140 -18188 18230 -18171
rect 18288 -18171 18688 -18124
rect 18288 -18188 18378 -18171
rect 18140 -18205 18156 -18188
rect 17904 -18221 18156 -18205
rect 18362 -18205 18378 -18188
rect 18598 -18188 18688 -18171
rect 18746 -18171 19146 -18124
rect 18746 -18188 18836 -18171
rect 18598 -18205 18614 -18188
rect 18362 -18221 18614 -18205
rect 18820 -18205 18836 -18188
rect 19056 -18188 19146 -18171
rect 19204 -18171 19604 -18124
rect 19204 -18188 19294 -18171
rect 19056 -18205 19072 -18188
rect 18820 -18221 19072 -18205
rect 19278 -18205 19294 -18188
rect 19514 -18188 19604 -18171
rect 19662 -18171 20062 -18124
rect 19662 -18188 19752 -18171
rect 19514 -18205 19530 -18188
rect 19278 -18221 19530 -18205
rect 19736 -18205 19752 -18188
rect 19972 -18188 20062 -18171
rect 20120 -18171 20520 -18124
rect 20120 -18188 20210 -18171
rect 19972 -18205 19988 -18188
rect 19736 -18221 19988 -18205
rect 20194 -18205 20210 -18188
rect 20430 -18188 20520 -18171
rect 20578 -18171 20978 -18124
rect 20578 -18188 20668 -18171
rect 20430 -18205 20446 -18188
rect 20194 -18221 20446 -18205
rect 20652 -18205 20668 -18188
rect 20888 -18188 20978 -18171
rect 21036 -18171 21436 -18124
rect 21036 -18188 21126 -18171
rect 20888 -18205 20904 -18188
rect 20652 -18221 20904 -18205
rect 21110 -18205 21126 -18188
rect 21346 -18188 21436 -18171
rect 21494 -18171 21894 -18124
rect 21494 -18188 21584 -18171
rect 21346 -18205 21362 -18188
rect 21110 -18221 21362 -18205
rect 21568 -18205 21584 -18188
rect 21804 -18188 21894 -18171
rect 21952 -18171 22352 -18124
rect 21952 -18188 22042 -18171
rect 21804 -18205 21820 -18188
rect 21568 -18221 21820 -18205
rect 22026 -18205 22042 -18188
rect 22262 -18188 22352 -18171
rect 22410 -18171 22810 -18124
rect 22410 -18188 22500 -18171
rect 22262 -18205 22278 -18188
rect 22026 -18221 22278 -18205
rect 22484 -18205 22500 -18188
rect 22720 -18188 22810 -18171
rect 22868 -18171 23268 -18124
rect 22868 -18188 22958 -18171
rect 22720 -18205 22736 -18188
rect 22484 -18221 22736 -18205
rect 22942 -18205 22958 -18188
rect 23178 -18188 23268 -18171
rect 23326 -18171 23726 -18124
rect 23326 -18188 23416 -18171
rect 23178 -18205 23194 -18188
rect 22942 -18221 23194 -18205
rect 23400 -18205 23416 -18188
rect 23636 -18188 23726 -18171
rect 23784 -18171 24184 -18124
rect 23784 -18188 23874 -18171
rect 23636 -18205 23652 -18188
rect 23400 -18221 23652 -18205
rect 23858 -18205 23874 -18188
rect 24094 -18188 24184 -18171
rect 24094 -18205 24110 -18188
rect 23858 -18221 24110 -18205
rect 30295 -14178 30547 -14162
rect 30295 -14195 30311 -14178
rect 30221 -14212 30311 -14195
rect 30531 -14195 30547 -14178
rect 30753 -14178 31005 -14162
rect 30753 -14195 30769 -14178
rect 30531 -14212 30621 -14195
rect 30221 -14259 30621 -14212
rect 30679 -14212 30769 -14195
rect 30989 -14195 31005 -14178
rect 31211 -14178 31463 -14162
rect 31211 -14195 31227 -14178
rect 30989 -14212 31079 -14195
rect 30679 -14259 31079 -14212
rect 31137 -14212 31227 -14195
rect 31447 -14195 31463 -14178
rect 31669 -14178 31921 -14162
rect 31669 -14195 31685 -14178
rect 31447 -14212 31537 -14195
rect 31137 -14259 31537 -14212
rect 31595 -14212 31685 -14195
rect 31905 -14195 31921 -14178
rect 32127 -14178 32379 -14162
rect 32127 -14195 32143 -14178
rect 31905 -14212 31995 -14195
rect 31595 -14259 31995 -14212
rect 32053 -14212 32143 -14195
rect 32363 -14195 32379 -14178
rect 32585 -14178 32837 -14162
rect 32585 -14195 32601 -14178
rect 32363 -14212 32453 -14195
rect 32053 -14259 32453 -14212
rect 32511 -14212 32601 -14195
rect 32821 -14195 32837 -14178
rect 33043 -14178 33295 -14162
rect 33043 -14195 33059 -14178
rect 32821 -14212 32911 -14195
rect 32511 -14259 32911 -14212
rect 32969 -14212 33059 -14195
rect 33279 -14195 33295 -14178
rect 33501 -14178 33753 -14162
rect 33501 -14195 33517 -14178
rect 33279 -14212 33369 -14195
rect 32969 -14259 33369 -14212
rect 33427 -14212 33517 -14195
rect 33737 -14195 33753 -14178
rect 33959 -14178 34211 -14162
rect 33959 -14195 33975 -14178
rect 33737 -14212 33827 -14195
rect 33427 -14259 33827 -14212
rect 33885 -14212 33975 -14195
rect 34195 -14195 34211 -14178
rect 34417 -14178 34669 -14162
rect 34417 -14195 34433 -14178
rect 34195 -14212 34285 -14195
rect 33885 -14259 34285 -14212
rect 34343 -14212 34433 -14195
rect 34653 -14195 34669 -14178
rect 35295 -14178 35547 -14162
rect 35295 -14195 35311 -14178
rect 34653 -14212 34743 -14195
rect 34343 -14259 34743 -14212
rect 35221 -14212 35311 -14195
rect 35531 -14195 35547 -14178
rect 35753 -14178 36005 -14162
rect 35753 -14195 35769 -14178
rect 35531 -14212 35621 -14195
rect 35221 -14259 35621 -14212
rect 35679 -14212 35769 -14195
rect 35989 -14195 36005 -14178
rect 36211 -14178 36463 -14162
rect 36211 -14195 36227 -14178
rect 35989 -14212 36079 -14195
rect 35679 -14259 36079 -14212
rect 36137 -14212 36227 -14195
rect 36447 -14195 36463 -14178
rect 36669 -14178 36921 -14162
rect 36669 -14195 36685 -14178
rect 36447 -14212 36537 -14195
rect 36137 -14259 36537 -14212
rect 36595 -14212 36685 -14195
rect 36905 -14195 36921 -14178
rect 37127 -14178 37379 -14162
rect 37127 -14195 37143 -14178
rect 36905 -14212 36995 -14195
rect 36595 -14259 36995 -14212
rect 37053 -14212 37143 -14195
rect 37363 -14195 37379 -14178
rect 37585 -14178 37837 -14162
rect 37585 -14195 37601 -14178
rect 37363 -14212 37453 -14195
rect 37053 -14259 37453 -14212
rect 37511 -14212 37601 -14195
rect 37821 -14195 37837 -14178
rect 38043 -14178 38295 -14162
rect 38043 -14195 38059 -14178
rect 37821 -14212 37911 -14195
rect 37511 -14259 37911 -14212
rect 37969 -14212 38059 -14195
rect 38279 -14195 38295 -14178
rect 38501 -14178 38753 -14162
rect 38501 -14195 38517 -14178
rect 38279 -14212 38369 -14195
rect 37969 -14259 38369 -14212
rect 38427 -14212 38517 -14195
rect 38737 -14195 38753 -14178
rect 38959 -14178 39211 -14162
rect 38959 -14195 38975 -14178
rect 38737 -14212 38827 -14195
rect 38427 -14259 38827 -14212
rect 38885 -14212 38975 -14195
rect 39195 -14195 39211 -14178
rect 39417 -14178 39669 -14162
rect 39417 -14195 39433 -14178
rect 39195 -14212 39285 -14195
rect 38885 -14259 39285 -14212
rect 39343 -14212 39433 -14195
rect 39653 -14195 39669 -14178
rect 39653 -14212 39743 -14195
rect 39343 -14259 39743 -14212
rect 30221 -15506 30621 -15459
rect 30221 -15523 30311 -15506
rect 30295 -15540 30311 -15523
rect 30531 -15523 30621 -15506
rect 30679 -15506 31079 -15459
rect 30679 -15523 30769 -15506
rect 30531 -15540 30547 -15523
rect 30295 -15556 30547 -15540
rect 30753 -15540 30769 -15523
rect 30989 -15523 31079 -15506
rect 31137 -15506 31537 -15459
rect 31137 -15523 31227 -15506
rect 30989 -15540 31005 -15523
rect 30753 -15556 31005 -15540
rect 31211 -15540 31227 -15523
rect 31447 -15523 31537 -15506
rect 31595 -15506 31995 -15459
rect 31595 -15523 31685 -15506
rect 31447 -15540 31463 -15523
rect 31211 -15556 31463 -15540
rect 31669 -15540 31685 -15523
rect 31905 -15523 31995 -15506
rect 32053 -15506 32453 -15459
rect 32053 -15523 32143 -15506
rect 31905 -15540 31921 -15523
rect 31669 -15556 31921 -15540
rect 32127 -15540 32143 -15523
rect 32363 -15523 32453 -15506
rect 32511 -15506 32911 -15459
rect 32511 -15523 32601 -15506
rect 32363 -15540 32379 -15523
rect 32127 -15556 32379 -15540
rect 32585 -15540 32601 -15523
rect 32821 -15523 32911 -15506
rect 32969 -15506 33369 -15459
rect 32969 -15523 33059 -15506
rect 32821 -15540 32837 -15523
rect 32585 -15556 32837 -15540
rect 33043 -15540 33059 -15523
rect 33279 -15523 33369 -15506
rect 33427 -15506 33827 -15459
rect 33427 -15523 33517 -15506
rect 33279 -15540 33295 -15523
rect 33043 -15556 33295 -15540
rect 33501 -15540 33517 -15523
rect 33737 -15523 33827 -15506
rect 33885 -15506 34285 -15459
rect 33885 -15523 33975 -15506
rect 33737 -15540 33753 -15523
rect 33501 -15556 33753 -15540
rect 33959 -15540 33975 -15523
rect 34195 -15523 34285 -15506
rect 34343 -15506 34743 -15459
rect 34343 -15523 34433 -15506
rect 34195 -15540 34211 -15523
rect 33959 -15556 34211 -15540
rect 34417 -15540 34433 -15523
rect 34653 -15523 34743 -15506
rect 35221 -15506 35621 -15459
rect 35221 -15523 35311 -15506
rect 34653 -15540 34669 -15523
rect 34417 -15556 34669 -15540
rect 35295 -15540 35311 -15523
rect 35531 -15523 35621 -15506
rect 35679 -15506 36079 -15459
rect 35679 -15523 35769 -15506
rect 35531 -15540 35547 -15523
rect 35295 -15556 35547 -15540
rect 35753 -15540 35769 -15523
rect 35989 -15523 36079 -15506
rect 36137 -15506 36537 -15459
rect 36137 -15523 36227 -15506
rect 35989 -15540 36005 -15523
rect 35753 -15556 36005 -15540
rect 36211 -15540 36227 -15523
rect 36447 -15523 36537 -15506
rect 36595 -15506 36995 -15459
rect 36595 -15523 36685 -15506
rect 36447 -15540 36463 -15523
rect 36211 -15556 36463 -15540
rect 36669 -15540 36685 -15523
rect 36905 -15523 36995 -15506
rect 37053 -15506 37453 -15459
rect 37053 -15523 37143 -15506
rect 36905 -15540 36921 -15523
rect 36669 -15556 36921 -15540
rect 37127 -15540 37143 -15523
rect 37363 -15523 37453 -15506
rect 37511 -15506 37911 -15459
rect 37511 -15523 37601 -15506
rect 37363 -15540 37379 -15523
rect 37127 -15556 37379 -15540
rect 37585 -15540 37601 -15523
rect 37821 -15523 37911 -15506
rect 37969 -15506 38369 -15459
rect 37969 -15523 38059 -15506
rect 37821 -15540 37837 -15523
rect 37585 -15556 37837 -15540
rect 38043 -15540 38059 -15523
rect 38279 -15523 38369 -15506
rect 38427 -15506 38827 -15459
rect 38427 -15523 38517 -15506
rect 38279 -15540 38295 -15523
rect 38043 -15556 38295 -15540
rect 38501 -15540 38517 -15523
rect 38737 -15523 38827 -15506
rect 38885 -15506 39285 -15459
rect 38885 -15523 38975 -15506
rect 38737 -15540 38753 -15523
rect 38501 -15556 38753 -15540
rect 38959 -15540 38975 -15523
rect 39195 -15523 39285 -15506
rect 39343 -15506 39743 -15459
rect 39343 -15523 39433 -15506
rect 39195 -15540 39211 -15523
rect 38959 -15556 39211 -15540
rect 39417 -15540 39433 -15523
rect 39653 -15523 39743 -15506
rect 39653 -15540 39669 -15523
rect 39417 -15556 39669 -15540
rect 31072 -16443 31324 -16427
rect 31072 -16460 31088 -16443
rect 30998 -16477 31088 -16460
rect 31308 -16460 31324 -16443
rect 31530 -16443 31782 -16427
rect 31530 -16460 31546 -16443
rect 31308 -16477 31398 -16460
rect 30998 -16524 31398 -16477
rect 31456 -16477 31546 -16460
rect 31766 -16460 31782 -16443
rect 31988 -16443 32240 -16427
rect 31988 -16460 32004 -16443
rect 31766 -16477 31856 -16460
rect 31456 -16524 31856 -16477
rect 31914 -16477 32004 -16460
rect 32224 -16460 32240 -16443
rect 32446 -16443 32698 -16427
rect 32446 -16460 32462 -16443
rect 32224 -16477 32314 -16460
rect 31914 -16524 32314 -16477
rect 32372 -16477 32462 -16460
rect 32682 -16460 32698 -16443
rect 32904 -16443 33156 -16427
rect 32904 -16460 32920 -16443
rect 32682 -16477 32772 -16460
rect 32372 -16524 32772 -16477
rect 32830 -16477 32920 -16460
rect 33140 -16460 33156 -16443
rect 33362 -16443 33614 -16427
rect 33362 -16460 33378 -16443
rect 33140 -16477 33230 -16460
rect 32830 -16524 33230 -16477
rect 33288 -16477 33378 -16460
rect 33598 -16460 33614 -16443
rect 33820 -16443 34072 -16427
rect 33820 -16460 33836 -16443
rect 33598 -16477 33688 -16460
rect 33288 -16524 33688 -16477
rect 33746 -16477 33836 -16460
rect 34056 -16460 34072 -16443
rect 34278 -16443 34530 -16427
rect 34278 -16460 34294 -16443
rect 34056 -16477 34146 -16460
rect 33746 -16524 34146 -16477
rect 34204 -16477 34294 -16460
rect 34514 -16460 34530 -16443
rect 34736 -16443 34988 -16427
rect 34736 -16460 34752 -16443
rect 34514 -16477 34604 -16460
rect 34204 -16524 34604 -16477
rect 34662 -16477 34752 -16460
rect 34972 -16460 34988 -16443
rect 35194 -16443 35446 -16427
rect 35194 -16460 35210 -16443
rect 34972 -16477 35062 -16460
rect 34662 -16524 35062 -16477
rect 35120 -16477 35210 -16460
rect 35430 -16460 35446 -16443
rect 35652 -16443 35904 -16427
rect 35652 -16460 35668 -16443
rect 35430 -16477 35520 -16460
rect 35120 -16524 35520 -16477
rect 35578 -16477 35668 -16460
rect 35888 -16460 35904 -16443
rect 36110 -16443 36362 -16427
rect 36110 -16460 36126 -16443
rect 35888 -16477 35978 -16460
rect 35578 -16524 35978 -16477
rect 36036 -16477 36126 -16460
rect 36346 -16460 36362 -16443
rect 36568 -16443 36820 -16427
rect 36568 -16460 36584 -16443
rect 36346 -16477 36436 -16460
rect 36036 -16524 36436 -16477
rect 36494 -16477 36584 -16460
rect 36804 -16460 36820 -16443
rect 37026 -16443 37278 -16427
rect 37026 -16460 37042 -16443
rect 36804 -16477 36894 -16460
rect 36494 -16524 36894 -16477
rect 36952 -16477 37042 -16460
rect 37262 -16460 37278 -16443
rect 37484 -16443 37736 -16427
rect 37484 -16460 37500 -16443
rect 37262 -16477 37352 -16460
rect 36952 -16524 37352 -16477
rect 37410 -16477 37500 -16460
rect 37720 -16460 37736 -16443
rect 37942 -16443 38194 -16427
rect 37942 -16460 37958 -16443
rect 37720 -16477 37810 -16460
rect 37410 -16524 37810 -16477
rect 37868 -16477 37958 -16460
rect 38178 -16460 38194 -16443
rect 38400 -16443 38652 -16427
rect 38400 -16460 38416 -16443
rect 38178 -16477 38268 -16460
rect 37868 -16524 38268 -16477
rect 38326 -16477 38416 -16460
rect 38636 -16460 38652 -16443
rect 38858 -16443 39110 -16427
rect 38858 -16460 38874 -16443
rect 38636 -16477 38726 -16460
rect 38326 -16524 38726 -16477
rect 38784 -16477 38874 -16460
rect 39094 -16460 39110 -16443
rect 39094 -16477 39184 -16460
rect 38784 -16524 39184 -16477
rect 30998 -18171 31398 -18124
rect 30998 -18188 31088 -18171
rect 31072 -18205 31088 -18188
rect 31308 -18188 31398 -18171
rect 31456 -18171 31856 -18124
rect 31456 -18188 31546 -18171
rect 31308 -18205 31324 -18188
rect 31072 -18221 31324 -18205
rect 31530 -18205 31546 -18188
rect 31766 -18188 31856 -18171
rect 31914 -18171 32314 -18124
rect 31914 -18188 32004 -18171
rect 31766 -18205 31782 -18188
rect 31530 -18221 31782 -18205
rect 31988 -18205 32004 -18188
rect 32224 -18188 32314 -18171
rect 32372 -18171 32772 -18124
rect 32372 -18188 32462 -18171
rect 32224 -18205 32240 -18188
rect 31988 -18221 32240 -18205
rect 32446 -18205 32462 -18188
rect 32682 -18188 32772 -18171
rect 32830 -18171 33230 -18124
rect 32830 -18188 32920 -18171
rect 32682 -18205 32698 -18188
rect 32446 -18221 32698 -18205
rect 32904 -18205 32920 -18188
rect 33140 -18188 33230 -18171
rect 33288 -18171 33688 -18124
rect 33288 -18188 33378 -18171
rect 33140 -18205 33156 -18188
rect 32904 -18221 33156 -18205
rect 33362 -18205 33378 -18188
rect 33598 -18188 33688 -18171
rect 33746 -18171 34146 -18124
rect 33746 -18188 33836 -18171
rect 33598 -18205 33614 -18188
rect 33362 -18221 33614 -18205
rect 33820 -18205 33836 -18188
rect 34056 -18188 34146 -18171
rect 34204 -18171 34604 -18124
rect 34204 -18188 34294 -18171
rect 34056 -18205 34072 -18188
rect 33820 -18221 34072 -18205
rect 34278 -18205 34294 -18188
rect 34514 -18188 34604 -18171
rect 34662 -18171 35062 -18124
rect 34662 -18188 34752 -18171
rect 34514 -18205 34530 -18188
rect 34278 -18221 34530 -18205
rect 34736 -18205 34752 -18188
rect 34972 -18188 35062 -18171
rect 35120 -18171 35520 -18124
rect 35120 -18188 35210 -18171
rect 34972 -18205 34988 -18188
rect 34736 -18221 34988 -18205
rect 35194 -18205 35210 -18188
rect 35430 -18188 35520 -18171
rect 35578 -18171 35978 -18124
rect 35578 -18188 35668 -18171
rect 35430 -18205 35446 -18188
rect 35194 -18221 35446 -18205
rect 35652 -18205 35668 -18188
rect 35888 -18188 35978 -18171
rect 36036 -18171 36436 -18124
rect 36036 -18188 36126 -18171
rect 35888 -18205 35904 -18188
rect 35652 -18221 35904 -18205
rect 36110 -18205 36126 -18188
rect 36346 -18188 36436 -18171
rect 36494 -18171 36894 -18124
rect 36494 -18188 36584 -18171
rect 36346 -18205 36362 -18188
rect 36110 -18221 36362 -18205
rect 36568 -18205 36584 -18188
rect 36804 -18188 36894 -18171
rect 36952 -18171 37352 -18124
rect 36952 -18188 37042 -18171
rect 36804 -18205 36820 -18188
rect 36568 -18221 36820 -18205
rect 37026 -18205 37042 -18188
rect 37262 -18188 37352 -18171
rect 37410 -18171 37810 -18124
rect 37410 -18188 37500 -18171
rect 37262 -18205 37278 -18188
rect 37026 -18221 37278 -18205
rect 37484 -18205 37500 -18188
rect 37720 -18188 37810 -18171
rect 37868 -18171 38268 -18124
rect 37868 -18188 37958 -18171
rect 37720 -18205 37736 -18188
rect 37484 -18221 37736 -18205
rect 37942 -18205 37958 -18188
rect 38178 -18188 38268 -18171
rect 38326 -18171 38726 -18124
rect 38326 -18188 38416 -18171
rect 38178 -18205 38194 -18188
rect 37942 -18221 38194 -18205
rect 38400 -18205 38416 -18188
rect 38636 -18188 38726 -18171
rect 38784 -18171 39184 -18124
rect 38784 -18188 38874 -18171
rect 38636 -18205 38652 -18188
rect 38400 -18221 38652 -18205
rect 38858 -18205 38874 -18188
rect 39094 -18188 39184 -18171
rect 39094 -18205 39110 -18188
rect 38858 -18221 39110 -18205
rect 11924 -21399 12176 -21383
rect 11924 -21416 11940 -21399
rect 11850 -21433 11940 -21416
rect 12160 -21416 12176 -21399
rect 12382 -21399 12634 -21383
rect 12382 -21416 12398 -21399
rect 12160 -21433 12250 -21416
rect 11850 -21480 12250 -21433
rect 12308 -21433 12398 -21416
rect 12618 -21416 12634 -21399
rect 12840 -21399 13092 -21383
rect 12840 -21416 12856 -21399
rect 12618 -21433 12708 -21416
rect 12308 -21480 12708 -21433
rect 12766 -21433 12856 -21416
rect 13076 -21416 13092 -21399
rect 13298 -21399 13550 -21383
rect 13298 -21416 13314 -21399
rect 13076 -21433 13166 -21416
rect 12766 -21480 13166 -21433
rect 13224 -21433 13314 -21416
rect 13534 -21416 13550 -21399
rect 13756 -21399 14008 -21383
rect 13756 -21416 13772 -21399
rect 13534 -21433 13624 -21416
rect 13224 -21480 13624 -21433
rect 13682 -21433 13772 -21416
rect 13992 -21416 14008 -21399
rect 14214 -21399 14466 -21383
rect 14214 -21416 14230 -21399
rect 13992 -21433 14082 -21416
rect 13682 -21480 14082 -21433
rect 14140 -21433 14230 -21416
rect 14450 -21416 14466 -21399
rect 14672 -21399 14924 -21383
rect 14672 -21416 14688 -21399
rect 14450 -21433 14540 -21416
rect 14140 -21480 14540 -21433
rect 14598 -21433 14688 -21416
rect 14908 -21416 14924 -21399
rect 15130 -21399 15382 -21383
rect 15130 -21416 15146 -21399
rect 14908 -21433 14998 -21416
rect 14598 -21480 14998 -21433
rect 15056 -21433 15146 -21416
rect 15366 -21416 15382 -21399
rect 15588 -21399 15840 -21383
rect 15588 -21416 15604 -21399
rect 15366 -21433 15456 -21416
rect 15056 -21480 15456 -21433
rect 15514 -21433 15604 -21416
rect 15824 -21416 15840 -21399
rect 16046 -21399 16298 -21383
rect 16046 -21416 16062 -21399
rect 15824 -21433 15914 -21416
rect 15514 -21480 15914 -21433
rect 15972 -21433 16062 -21416
rect 16282 -21416 16298 -21399
rect 16504 -21399 16756 -21383
rect 16504 -21416 16520 -21399
rect 16282 -21433 16372 -21416
rect 15972 -21480 16372 -21433
rect 16430 -21433 16520 -21416
rect 16740 -21416 16756 -21399
rect 16962 -21399 17214 -21383
rect 16962 -21416 16978 -21399
rect 16740 -21433 16830 -21416
rect 16430 -21480 16830 -21433
rect 16888 -21433 16978 -21416
rect 17198 -21416 17214 -21399
rect 17420 -21399 17672 -21383
rect 17420 -21416 17436 -21399
rect 17198 -21433 17288 -21416
rect 16888 -21480 17288 -21433
rect 17346 -21433 17436 -21416
rect 17656 -21416 17672 -21399
rect 17878 -21399 18130 -21383
rect 17878 -21416 17894 -21399
rect 17656 -21433 17746 -21416
rect 17346 -21480 17746 -21433
rect 17804 -21433 17894 -21416
rect 18114 -21416 18130 -21399
rect 18336 -21399 18588 -21383
rect 18336 -21416 18352 -21399
rect 18114 -21433 18204 -21416
rect 17804 -21480 18204 -21433
rect 18262 -21433 18352 -21416
rect 18572 -21416 18588 -21399
rect 18794 -21399 19046 -21383
rect 18794 -21416 18810 -21399
rect 18572 -21433 18662 -21416
rect 18262 -21480 18662 -21433
rect 18720 -21433 18810 -21416
rect 19030 -21416 19046 -21399
rect 19252 -21399 19504 -21383
rect 19252 -21416 19268 -21399
rect 19030 -21433 19120 -21416
rect 18720 -21480 19120 -21433
rect 19178 -21433 19268 -21416
rect 19488 -21416 19504 -21399
rect 19710 -21399 19962 -21383
rect 19710 -21416 19726 -21399
rect 19488 -21433 19578 -21416
rect 19178 -21480 19578 -21433
rect 19636 -21433 19726 -21416
rect 19946 -21416 19962 -21399
rect 19946 -21433 20036 -21416
rect 19636 -21480 20036 -21433
rect 11850 -23127 12250 -23080
rect 11850 -23144 11940 -23127
rect 11924 -23161 11940 -23144
rect 12160 -23144 12250 -23127
rect 12308 -23127 12708 -23080
rect 12308 -23144 12398 -23127
rect 12160 -23161 12176 -23144
rect 11924 -23177 12176 -23161
rect 12382 -23161 12398 -23144
rect 12618 -23144 12708 -23127
rect 12766 -23127 13166 -23080
rect 12766 -23144 12856 -23127
rect 12618 -23161 12634 -23144
rect 12382 -23177 12634 -23161
rect 12840 -23161 12856 -23144
rect 13076 -23144 13166 -23127
rect 13224 -23127 13624 -23080
rect 13224 -23144 13314 -23127
rect 13076 -23161 13092 -23144
rect 12840 -23177 13092 -23161
rect 13298 -23161 13314 -23144
rect 13534 -23144 13624 -23127
rect 13682 -23127 14082 -23080
rect 13682 -23144 13772 -23127
rect 13534 -23161 13550 -23144
rect 13298 -23177 13550 -23161
rect 13756 -23161 13772 -23144
rect 13992 -23144 14082 -23127
rect 14140 -23127 14540 -23080
rect 14140 -23144 14230 -23127
rect 13992 -23161 14008 -23144
rect 13756 -23177 14008 -23161
rect 14214 -23161 14230 -23144
rect 14450 -23144 14540 -23127
rect 14598 -23127 14998 -23080
rect 14598 -23144 14688 -23127
rect 14450 -23161 14466 -23144
rect 14214 -23177 14466 -23161
rect 14672 -23161 14688 -23144
rect 14908 -23144 14998 -23127
rect 15056 -23127 15456 -23080
rect 15056 -23144 15146 -23127
rect 14908 -23161 14924 -23144
rect 14672 -23177 14924 -23161
rect 15130 -23161 15146 -23144
rect 15366 -23144 15456 -23127
rect 15514 -23127 15914 -23080
rect 15514 -23144 15604 -23127
rect 15366 -23161 15382 -23144
rect 15130 -23177 15382 -23161
rect 15588 -23161 15604 -23144
rect 15824 -23144 15914 -23127
rect 15972 -23127 16372 -23080
rect 15972 -23144 16062 -23127
rect 15824 -23161 15840 -23144
rect 15588 -23177 15840 -23161
rect 16046 -23161 16062 -23144
rect 16282 -23144 16372 -23127
rect 16430 -23127 16830 -23080
rect 16430 -23144 16520 -23127
rect 16282 -23161 16298 -23144
rect 16046 -23177 16298 -23161
rect 16504 -23161 16520 -23144
rect 16740 -23144 16830 -23127
rect 16888 -23127 17288 -23080
rect 16888 -23144 16978 -23127
rect 16740 -23161 16756 -23144
rect 16504 -23177 16756 -23161
rect 16962 -23161 16978 -23144
rect 17198 -23144 17288 -23127
rect 17346 -23127 17746 -23080
rect 17346 -23144 17436 -23127
rect 17198 -23161 17214 -23144
rect 16962 -23177 17214 -23161
rect 17420 -23161 17436 -23144
rect 17656 -23144 17746 -23127
rect 17804 -23127 18204 -23080
rect 17804 -23144 17894 -23127
rect 17656 -23161 17672 -23144
rect 17420 -23177 17672 -23161
rect 17878 -23161 17894 -23144
rect 18114 -23144 18204 -23127
rect 18262 -23127 18662 -23080
rect 18262 -23144 18352 -23127
rect 18114 -23161 18130 -23144
rect 17878 -23177 18130 -23161
rect 18336 -23161 18352 -23144
rect 18572 -23144 18662 -23127
rect 18720 -23127 19120 -23080
rect 18720 -23144 18810 -23127
rect 18572 -23161 18588 -23144
rect 18336 -23177 18588 -23161
rect 18794 -23161 18810 -23144
rect 19030 -23144 19120 -23127
rect 19178 -23127 19578 -23080
rect 19178 -23144 19268 -23127
rect 19030 -23161 19046 -23144
rect 18794 -23177 19046 -23161
rect 19252 -23161 19268 -23144
rect 19488 -23144 19578 -23127
rect 19636 -23127 20036 -23080
rect 19636 -23144 19726 -23127
rect 19488 -23161 19504 -23144
rect 19252 -23177 19504 -23161
rect 19710 -23161 19726 -23144
rect 19946 -23144 20036 -23127
rect 19946 -23161 19962 -23144
rect 19710 -23177 19962 -23161
rect 11365 -24064 11617 -24048
rect 11365 -24081 11381 -24064
rect 11291 -24098 11381 -24081
rect 11601 -24081 11617 -24064
rect 11823 -24064 12075 -24048
rect 11823 -24081 11839 -24064
rect 11601 -24098 11691 -24081
rect 11291 -24145 11691 -24098
rect 11749 -24098 11839 -24081
rect 12059 -24081 12075 -24064
rect 12281 -24064 12533 -24048
rect 12281 -24081 12297 -24064
rect 12059 -24098 12149 -24081
rect 11749 -24145 12149 -24098
rect 12207 -24098 12297 -24081
rect 12517 -24081 12533 -24064
rect 12739 -24064 12991 -24048
rect 12739 -24081 12755 -24064
rect 12517 -24098 12607 -24081
rect 12207 -24145 12607 -24098
rect 12665 -24098 12755 -24081
rect 12975 -24081 12991 -24064
rect 13197 -24064 13449 -24048
rect 13197 -24081 13213 -24064
rect 12975 -24098 13065 -24081
rect 12665 -24145 13065 -24098
rect 13123 -24098 13213 -24081
rect 13433 -24081 13449 -24064
rect 13655 -24064 13907 -24048
rect 13655 -24081 13671 -24064
rect 13433 -24098 13523 -24081
rect 13123 -24145 13523 -24098
rect 13581 -24098 13671 -24081
rect 13891 -24081 13907 -24064
rect 14113 -24064 14365 -24048
rect 14113 -24081 14129 -24064
rect 13891 -24098 13981 -24081
rect 13581 -24145 13981 -24098
rect 14039 -24098 14129 -24081
rect 14349 -24081 14365 -24064
rect 14571 -24064 14823 -24048
rect 14571 -24081 14587 -24064
rect 14349 -24098 14439 -24081
rect 14039 -24145 14439 -24098
rect 14497 -24098 14587 -24081
rect 14807 -24081 14823 -24064
rect 15029 -24064 15281 -24048
rect 15029 -24081 15045 -24064
rect 14807 -24098 14897 -24081
rect 14497 -24145 14897 -24098
rect 14955 -24098 15045 -24081
rect 15265 -24081 15281 -24064
rect 15487 -24064 15739 -24048
rect 15487 -24081 15503 -24064
rect 15265 -24098 15355 -24081
rect 14955 -24145 15355 -24098
rect 15413 -24098 15503 -24081
rect 15723 -24081 15739 -24064
rect 16365 -24064 16617 -24048
rect 16365 -24081 16381 -24064
rect 15723 -24098 15813 -24081
rect 15413 -24145 15813 -24098
rect 16291 -24098 16381 -24081
rect 16601 -24081 16617 -24064
rect 16823 -24064 17075 -24048
rect 16823 -24081 16839 -24064
rect 16601 -24098 16691 -24081
rect 16291 -24145 16691 -24098
rect 16749 -24098 16839 -24081
rect 17059 -24081 17075 -24064
rect 17281 -24064 17533 -24048
rect 17281 -24081 17297 -24064
rect 17059 -24098 17149 -24081
rect 16749 -24145 17149 -24098
rect 17207 -24098 17297 -24081
rect 17517 -24081 17533 -24064
rect 17739 -24064 17991 -24048
rect 17739 -24081 17755 -24064
rect 17517 -24098 17607 -24081
rect 17207 -24145 17607 -24098
rect 17665 -24098 17755 -24081
rect 17975 -24081 17991 -24064
rect 18197 -24064 18449 -24048
rect 18197 -24081 18213 -24064
rect 17975 -24098 18065 -24081
rect 17665 -24145 18065 -24098
rect 18123 -24098 18213 -24081
rect 18433 -24081 18449 -24064
rect 18655 -24064 18907 -24048
rect 18655 -24081 18671 -24064
rect 18433 -24098 18523 -24081
rect 18123 -24145 18523 -24098
rect 18581 -24098 18671 -24081
rect 18891 -24081 18907 -24064
rect 19113 -24064 19365 -24048
rect 19113 -24081 19129 -24064
rect 18891 -24098 18981 -24081
rect 18581 -24145 18981 -24098
rect 19039 -24098 19129 -24081
rect 19349 -24081 19365 -24064
rect 19571 -24064 19823 -24048
rect 19571 -24081 19587 -24064
rect 19349 -24098 19439 -24081
rect 19039 -24145 19439 -24098
rect 19497 -24098 19587 -24081
rect 19807 -24081 19823 -24064
rect 20029 -24064 20281 -24048
rect 20029 -24081 20045 -24064
rect 19807 -24098 19897 -24081
rect 19497 -24145 19897 -24098
rect 19955 -24098 20045 -24081
rect 20265 -24081 20281 -24064
rect 20487 -24064 20739 -24048
rect 20487 -24081 20503 -24064
rect 20265 -24098 20355 -24081
rect 19955 -24145 20355 -24098
rect 20413 -24098 20503 -24081
rect 20723 -24081 20739 -24064
rect 20723 -24098 20813 -24081
rect 20413 -24145 20813 -24098
rect 11291 -25392 11691 -25345
rect 11291 -25409 11381 -25392
rect 11365 -25426 11381 -25409
rect 11601 -25409 11691 -25392
rect 11749 -25392 12149 -25345
rect 11749 -25409 11839 -25392
rect 11601 -25426 11617 -25409
rect 11365 -25442 11617 -25426
rect 11823 -25426 11839 -25409
rect 12059 -25409 12149 -25392
rect 12207 -25392 12607 -25345
rect 12207 -25409 12297 -25392
rect 12059 -25426 12075 -25409
rect 11823 -25442 12075 -25426
rect 12281 -25426 12297 -25409
rect 12517 -25409 12607 -25392
rect 12665 -25392 13065 -25345
rect 12665 -25409 12755 -25392
rect 12517 -25426 12533 -25409
rect 12281 -25442 12533 -25426
rect 12739 -25426 12755 -25409
rect 12975 -25409 13065 -25392
rect 13123 -25392 13523 -25345
rect 13123 -25409 13213 -25392
rect 12975 -25426 12991 -25409
rect 12739 -25442 12991 -25426
rect 13197 -25426 13213 -25409
rect 13433 -25409 13523 -25392
rect 13581 -25392 13981 -25345
rect 13581 -25409 13671 -25392
rect 13433 -25426 13449 -25409
rect 13197 -25442 13449 -25426
rect 13655 -25426 13671 -25409
rect 13891 -25409 13981 -25392
rect 14039 -25392 14439 -25345
rect 14039 -25409 14129 -25392
rect 13891 -25426 13907 -25409
rect 13655 -25442 13907 -25426
rect 14113 -25426 14129 -25409
rect 14349 -25409 14439 -25392
rect 14497 -25392 14897 -25345
rect 14497 -25409 14587 -25392
rect 14349 -25426 14365 -25409
rect 14113 -25442 14365 -25426
rect 14571 -25426 14587 -25409
rect 14807 -25409 14897 -25392
rect 14955 -25392 15355 -25345
rect 14955 -25409 15045 -25392
rect 14807 -25426 14823 -25409
rect 14571 -25442 14823 -25426
rect 15029 -25426 15045 -25409
rect 15265 -25409 15355 -25392
rect 15413 -25392 15813 -25345
rect 15413 -25409 15503 -25392
rect 15265 -25426 15281 -25409
rect 15029 -25442 15281 -25426
rect 15487 -25426 15503 -25409
rect 15723 -25409 15813 -25392
rect 16291 -25392 16691 -25345
rect 16291 -25409 16381 -25392
rect 15723 -25426 15739 -25409
rect 15487 -25442 15739 -25426
rect 16365 -25426 16381 -25409
rect 16601 -25409 16691 -25392
rect 16749 -25392 17149 -25345
rect 16749 -25409 16839 -25392
rect 16601 -25426 16617 -25409
rect 16365 -25442 16617 -25426
rect 16823 -25426 16839 -25409
rect 17059 -25409 17149 -25392
rect 17207 -25392 17607 -25345
rect 17207 -25409 17297 -25392
rect 17059 -25426 17075 -25409
rect 16823 -25442 17075 -25426
rect 17281 -25426 17297 -25409
rect 17517 -25409 17607 -25392
rect 17665 -25392 18065 -25345
rect 17665 -25409 17755 -25392
rect 17517 -25426 17533 -25409
rect 17281 -25442 17533 -25426
rect 17739 -25426 17755 -25409
rect 17975 -25409 18065 -25392
rect 18123 -25392 18523 -25345
rect 18123 -25409 18213 -25392
rect 17975 -25426 17991 -25409
rect 17739 -25442 17991 -25426
rect 18197 -25426 18213 -25409
rect 18433 -25409 18523 -25392
rect 18581 -25392 18981 -25345
rect 18581 -25409 18671 -25392
rect 18433 -25426 18449 -25409
rect 18197 -25442 18449 -25426
rect 18655 -25426 18671 -25409
rect 18891 -25409 18981 -25392
rect 19039 -25392 19439 -25345
rect 19039 -25409 19129 -25392
rect 18891 -25426 18907 -25409
rect 18655 -25442 18907 -25426
rect 19113 -25426 19129 -25409
rect 19349 -25409 19439 -25392
rect 19497 -25392 19897 -25345
rect 19497 -25409 19587 -25392
rect 19349 -25426 19365 -25409
rect 19113 -25442 19365 -25426
rect 19571 -25426 19587 -25409
rect 19807 -25409 19897 -25392
rect 19955 -25392 20355 -25345
rect 19955 -25409 20045 -25392
rect 19807 -25426 19823 -25409
rect 19571 -25442 19823 -25426
rect 20029 -25426 20045 -25409
rect 20265 -25409 20355 -25392
rect 20413 -25392 20813 -25345
rect 20413 -25409 20503 -25392
rect 20265 -25426 20281 -25409
rect 20029 -25442 20281 -25426
rect 20487 -25426 20503 -25409
rect 20723 -25409 20813 -25392
rect 20723 -25426 20739 -25409
rect 20487 -25442 20739 -25426
rect 26924 -21399 27176 -21383
rect 26924 -21416 26940 -21399
rect 26850 -21433 26940 -21416
rect 27160 -21416 27176 -21399
rect 27382 -21399 27634 -21383
rect 27382 -21416 27398 -21399
rect 27160 -21433 27250 -21416
rect 26850 -21480 27250 -21433
rect 27308 -21433 27398 -21416
rect 27618 -21416 27634 -21399
rect 27840 -21399 28092 -21383
rect 27840 -21416 27856 -21399
rect 27618 -21433 27708 -21416
rect 27308 -21480 27708 -21433
rect 27766 -21433 27856 -21416
rect 28076 -21416 28092 -21399
rect 28298 -21399 28550 -21383
rect 28298 -21416 28314 -21399
rect 28076 -21433 28166 -21416
rect 27766 -21480 28166 -21433
rect 28224 -21433 28314 -21416
rect 28534 -21416 28550 -21399
rect 28756 -21399 29008 -21383
rect 28756 -21416 28772 -21399
rect 28534 -21433 28624 -21416
rect 28224 -21480 28624 -21433
rect 28682 -21433 28772 -21416
rect 28992 -21416 29008 -21399
rect 29214 -21399 29466 -21383
rect 29214 -21416 29230 -21399
rect 28992 -21433 29082 -21416
rect 28682 -21480 29082 -21433
rect 29140 -21433 29230 -21416
rect 29450 -21416 29466 -21399
rect 29672 -21399 29924 -21383
rect 29672 -21416 29688 -21399
rect 29450 -21433 29540 -21416
rect 29140 -21480 29540 -21433
rect 29598 -21433 29688 -21416
rect 29908 -21416 29924 -21399
rect 30130 -21399 30382 -21383
rect 30130 -21416 30146 -21399
rect 29908 -21433 29998 -21416
rect 29598 -21480 29998 -21433
rect 30056 -21433 30146 -21416
rect 30366 -21416 30382 -21399
rect 30588 -21399 30840 -21383
rect 30588 -21416 30604 -21399
rect 30366 -21433 30456 -21416
rect 30056 -21480 30456 -21433
rect 30514 -21433 30604 -21416
rect 30824 -21416 30840 -21399
rect 31046 -21399 31298 -21383
rect 31046 -21416 31062 -21399
rect 30824 -21433 30914 -21416
rect 30514 -21480 30914 -21433
rect 30972 -21433 31062 -21416
rect 31282 -21416 31298 -21399
rect 31504 -21399 31756 -21383
rect 31504 -21416 31520 -21399
rect 31282 -21433 31372 -21416
rect 30972 -21480 31372 -21433
rect 31430 -21433 31520 -21416
rect 31740 -21416 31756 -21399
rect 31962 -21399 32214 -21383
rect 31962 -21416 31978 -21399
rect 31740 -21433 31830 -21416
rect 31430 -21480 31830 -21433
rect 31888 -21433 31978 -21416
rect 32198 -21416 32214 -21399
rect 32420 -21399 32672 -21383
rect 32420 -21416 32436 -21399
rect 32198 -21433 32288 -21416
rect 31888 -21480 32288 -21433
rect 32346 -21433 32436 -21416
rect 32656 -21416 32672 -21399
rect 32878 -21399 33130 -21383
rect 32878 -21416 32894 -21399
rect 32656 -21433 32746 -21416
rect 32346 -21480 32746 -21433
rect 32804 -21433 32894 -21416
rect 33114 -21416 33130 -21399
rect 33336 -21399 33588 -21383
rect 33336 -21416 33352 -21399
rect 33114 -21433 33204 -21416
rect 32804 -21480 33204 -21433
rect 33262 -21433 33352 -21416
rect 33572 -21416 33588 -21399
rect 33794 -21399 34046 -21383
rect 33794 -21416 33810 -21399
rect 33572 -21433 33662 -21416
rect 33262 -21480 33662 -21433
rect 33720 -21433 33810 -21416
rect 34030 -21416 34046 -21399
rect 34252 -21399 34504 -21383
rect 34252 -21416 34268 -21399
rect 34030 -21433 34120 -21416
rect 33720 -21480 34120 -21433
rect 34178 -21433 34268 -21416
rect 34488 -21416 34504 -21399
rect 34710 -21399 34962 -21383
rect 34710 -21416 34726 -21399
rect 34488 -21433 34578 -21416
rect 34178 -21480 34578 -21433
rect 34636 -21433 34726 -21416
rect 34946 -21416 34962 -21399
rect 34946 -21433 35036 -21416
rect 34636 -21480 35036 -21433
rect 26850 -23127 27250 -23080
rect 26850 -23144 26940 -23127
rect 26924 -23161 26940 -23144
rect 27160 -23144 27250 -23127
rect 27308 -23127 27708 -23080
rect 27308 -23144 27398 -23127
rect 27160 -23161 27176 -23144
rect 26924 -23177 27176 -23161
rect 27382 -23161 27398 -23144
rect 27618 -23144 27708 -23127
rect 27766 -23127 28166 -23080
rect 27766 -23144 27856 -23127
rect 27618 -23161 27634 -23144
rect 27382 -23177 27634 -23161
rect 27840 -23161 27856 -23144
rect 28076 -23144 28166 -23127
rect 28224 -23127 28624 -23080
rect 28224 -23144 28314 -23127
rect 28076 -23161 28092 -23144
rect 27840 -23177 28092 -23161
rect 28298 -23161 28314 -23144
rect 28534 -23144 28624 -23127
rect 28682 -23127 29082 -23080
rect 28682 -23144 28772 -23127
rect 28534 -23161 28550 -23144
rect 28298 -23177 28550 -23161
rect 28756 -23161 28772 -23144
rect 28992 -23144 29082 -23127
rect 29140 -23127 29540 -23080
rect 29140 -23144 29230 -23127
rect 28992 -23161 29008 -23144
rect 28756 -23177 29008 -23161
rect 29214 -23161 29230 -23144
rect 29450 -23144 29540 -23127
rect 29598 -23127 29998 -23080
rect 29598 -23144 29688 -23127
rect 29450 -23161 29466 -23144
rect 29214 -23177 29466 -23161
rect 29672 -23161 29688 -23144
rect 29908 -23144 29998 -23127
rect 30056 -23127 30456 -23080
rect 30056 -23144 30146 -23127
rect 29908 -23161 29924 -23144
rect 29672 -23177 29924 -23161
rect 30130 -23161 30146 -23144
rect 30366 -23144 30456 -23127
rect 30514 -23127 30914 -23080
rect 30514 -23144 30604 -23127
rect 30366 -23161 30382 -23144
rect 30130 -23177 30382 -23161
rect 30588 -23161 30604 -23144
rect 30824 -23144 30914 -23127
rect 30972 -23127 31372 -23080
rect 30972 -23144 31062 -23127
rect 30824 -23161 30840 -23144
rect 30588 -23177 30840 -23161
rect 31046 -23161 31062 -23144
rect 31282 -23144 31372 -23127
rect 31430 -23127 31830 -23080
rect 31430 -23144 31520 -23127
rect 31282 -23161 31298 -23144
rect 31046 -23177 31298 -23161
rect 31504 -23161 31520 -23144
rect 31740 -23144 31830 -23127
rect 31888 -23127 32288 -23080
rect 31888 -23144 31978 -23127
rect 31740 -23161 31756 -23144
rect 31504 -23177 31756 -23161
rect 31962 -23161 31978 -23144
rect 32198 -23144 32288 -23127
rect 32346 -23127 32746 -23080
rect 32346 -23144 32436 -23127
rect 32198 -23161 32214 -23144
rect 31962 -23177 32214 -23161
rect 32420 -23161 32436 -23144
rect 32656 -23144 32746 -23127
rect 32804 -23127 33204 -23080
rect 32804 -23144 32894 -23127
rect 32656 -23161 32672 -23144
rect 32420 -23177 32672 -23161
rect 32878 -23161 32894 -23144
rect 33114 -23144 33204 -23127
rect 33262 -23127 33662 -23080
rect 33262 -23144 33352 -23127
rect 33114 -23161 33130 -23144
rect 32878 -23177 33130 -23161
rect 33336 -23161 33352 -23144
rect 33572 -23144 33662 -23127
rect 33720 -23127 34120 -23080
rect 33720 -23144 33810 -23127
rect 33572 -23161 33588 -23144
rect 33336 -23177 33588 -23161
rect 33794 -23161 33810 -23144
rect 34030 -23144 34120 -23127
rect 34178 -23127 34578 -23080
rect 34178 -23144 34268 -23127
rect 34030 -23161 34046 -23144
rect 33794 -23177 34046 -23161
rect 34252 -23161 34268 -23144
rect 34488 -23144 34578 -23127
rect 34636 -23127 35036 -23080
rect 34636 -23144 34726 -23127
rect 34488 -23161 34504 -23144
rect 34252 -23177 34504 -23161
rect 34710 -23161 34726 -23144
rect 34946 -23144 35036 -23127
rect 34946 -23161 34962 -23144
rect 34710 -23177 34962 -23161
rect 26365 -24064 26617 -24048
rect 26365 -24081 26381 -24064
rect 26291 -24098 26381 -24081
rect 26601 -24081 26617 -24064
rect 26823 -24064 27075 -24048
rect 26823 -24081 26839 -24064
rect 26601 -24098 26691 -24081
rect 26291 -24145 26691 -24098
rect 26749 -24098 26839 -24081
rect 27059 -24081 27075 -24064
rect 27281 -24064 27533 -24048
rect 27281 -24081 27297 -24064
rect 27059 -24098 27149 -24081
rect 26749 -24145 27149 -24098
rect 27207 -24098 27297 -24081
rect 27517 -24081 27533 -24064
rect 27739 -24064 27991 -24048
rect 27739 -24081 27755 -24064
rect 27517 -24098 27607 -24081
rect 27207 -24145 27607 -24098
rect 27665 -24098 27755 -24081
rect 27975 -24081 27991 -24064
rect 28197 -24064 28449 -24048
rect 28197 -24081 28213 -24064
rect 27975 -24098 28065 -24081
rect 27665 -24145 28065 -24098
rect 28123 -24098 28213 -24081
rect 28433 -24081 28449 -24064
rect 28655 -24064 28907 -24048
rect 28655 -24081 28671 -24064
rect 28433 -24098 28523 -24081
rect 28123 -24145 28523 -24098
rect 28581 -24098 28671 -24081
rect 28891 -24081 28907 -24064
rect 29113 -24064 29365 -24048
rect 29113 -24081 29129 -24064
rect 28891 -24098 28981 -24081
rect 28581 -24145 28981 -24098
rect 29039 -24098 29129 -24081
rect 29349 -24081 29365 -24064
rect 29571 -24064 29823 -24048
rect 29571 -24081 29587 -24064
rect 29349 -24098 29439 -24081
rect 29039 -24145 29439 -24098
rect 29497 -24098 29587 -24081
rect 29807 -24081 29823 -24064
rect 30029 -24064 30281 -24048
rect 30029 -24081 30045 -24064
rect 29807 -24098 29897 -24081
rect 29497 -24145 29897 -24098
rect 29955 -24098 30045 -24081
rect 30265 -24081 30281 -24064
rect 30487 -24064 30739 -24048
rect 30487 -24081 30503 -24064
rect 30265 -24098 30355 -24081
rect 29955 -24145 30355 -24098
rect 30413 -24098 30503 -24081
rect 30723 -24081 30739 -24064
rect 31365 -24064 31617 -24048
rect 31365 -24081 31381 -24064
rect 30723 -24098 30813 -24081
rect 30413 -24145 30813 -24098
rect 31291 -24098 31381 -24081
rect 31601 -24081 31617 -24064
rect 31823 -24064 32075 -24048
rect 31823 -24081 31839 -24064
rect 31601 -24098 31691 -24081
rect 31291 -24145 31691 -24098
rect 31749 -24098 31839 -24081
rect 32059 -24081 32075 -24064
rect 32281 -24064 32533 -24048
rect 32281 -24081 32297 -24064
rect 32059 -24098 32149 -24081
rect 31749 -24145 32149 -24098
rect 32207 -24098 32297 -24081
rect 32517 -24081 32533 -24064
rect 32739 -24064 32991 -24048
rect 32739 -24081 32755 -24064
rect 32517 -24098 32607 -24081
rect 32207 -24145 32607 -24098
rect 32665 -24098 32755 -24081
rect 32975 -24081 32991 -24064
rect 33197 -24064 33449 -24048
rect 33197 -24081 33213 -24064
rect 32975 -24098 33065 -24081
rect 32665 -24145 33065 -24098
rect 33123 -24098 33213 -24081
rect 33433 -24081 33449 -24064
rect 33655 -24064 33907 -24048
rect 33655 -24081 33671 -24064
rect 33433 -24098 33523 -24081
rect 33123 -24145 33523 -24098
rect 33581 -24098 33671 -24081
rect 33891 -24081 33907 -24064
rect 34113 -24064 34365 -24048
rect 34113 -24081 34129 -24064
rect 33891 -24098 33981 -24081
rect 33581 -24145 33981 -24098
rect 34039 -24098 34129 -24081
rect 34349 -24081 34365 -24064
rect 34571 -24064 34823 -24048
rect 34571 -24081 34587 -24064
rect 34349 -24098 34439 -24081
rect 34039 -24145 34439 -24098
rect 34497 -24098 34587 -24081
rect 34807 -24081 34823 -24064
rect 35029 -24064 35281 -24048
rect 35029 -24081 35045 -24064
rect 34807 -24098 34897 -24081
rect 34497 -24145 34897 -24098
rect 34955 -24098 35045 -24081
rect 35265 -24081 35281 -24064
rect 35487 -24064 35739 -24048
rect 35487 -24081 35503 -24064
rect 35265 -24098 35355 -24081
rect 34955 -24145 35355 -24098
rect 35413 -24098 35503 -24081
rect 35723 -24081 35739 -24064
rect 35723 -24098 35813 -24081
rect 35413 -24145 35813 -24098
rect 26291 -25392 26691 -25345
rect 26291 -25409 26381 -25392
rect 26365 -25426 26381 -25409
rect 26601 -25409 26691 -25392
rect 26749 -25392 27149 -25345
rect 26749 -25409 26839 -25392
rect 26601 -25426 26617 -25409
rect 26365 -25442 26617 -25426
rect 26823 -25426 26839 -25409
rect 27059 -25409 27149 -25392
rect 27207 -25392 27607 -25345
rect 27207 -25409 27297 -25392
rect 27059 -25426 27075 -25409
rect 26823 -25442 27075 -25426
rect 27281 -25426 27297 -25409
rect 27517 -25409 27607 -25392
rect 27665 -25392 28065 -25345
rect 27665 -25409 27755 -25392
rect 27517 -25426 27533 -25409
rect 27281 -25442 27533 -25426
rect 27739 -25426 27755 -25409
rect 27975 -25409 28065 -25392
rect 28123 -25392 28523 -25345
rect 28123 -25409 28213 -25392
rect 27975 -25426 27991 -25409
rect 27739 -25442 27991 -25426
rect 28197 -25426 28213 -25409
rect 28433 -25409 28523 -25392
rect 28581 -25392 28981 -25345
rect 28581 -25409 28671 -25392
rect 28433 -25426 28449 -25409
rect 28197 -25442 28449 -25426
rect 28655 -25426 28671 -25409
rect 28891 -25409 28981 -25392
rect 29039 -25392 29439 -25345
rect 29039 -25409 29129 -25392
rect 28891 -25426 28907 -25409
rect 28655 -25442 28907 -25426
rect 29113 -25426 29129 -25409
rect 29349 -25409 29439 -25392
rect 29497 -25392 29897 -25345
rect 29497 -25409 29587 -25392
rect 29349 -25426 29365 -25409
rect 29113 -25442 29365 -25426
rect 29571 -25426 29587 -25409
rect 29807 -25409 29897 -25392
rect 29955 -25392 30355 -25345
rect 29955 -25409 30045 -25392
rect 29807 -25426 29823 -25409
rect 29571 -25442 29823 -25426
rect 30029 -25426 30045 -25409
rect 30265 -25409 30355 -25392
rect 30413 -25392 30813 -25345
rect 30413 -25409 30503 -25392
rect 30265 -25426 30281 -25409
rect 30029 -25442 30281 -25426
rect 30487 -25426 30503 -25409
rect 30723 -25409 30813 -25392
rect 31291 -25392 31691 -25345
rect 31291 -25409 31381 -25392
rect 30723 -25426 30739 -25409
rect 30487 -25442 30739 -25426
rect 31365 -25426 31381 -25409
rect 31601 -25409 31691 -25392
rect 31749 -25392 32149 -25345
rect 31749 -25409 31839 -25392
rect 31601 -25426 31617 -25409
rect 31365 -25442 31617 -25426
rect 31823 -25426 31839 -25409
rect 32059 -25409 32149 -25392
rect 32207 -25392 32607 -25345
rect 32207 -25409 32297 -25392
rect 32059 -25426 32075 -25409
rect 31823 -25442 32075 -25426
rect 32281 -25426 32297 -25409
rect 32517 -25409 32607 -25392
rect 32665 -25392 33065 -25345
rect 32665 -25409 32755 -25392
rect 32517 -25426 32533 -25409
rect 32281 -25442 32533 -25426
rect 32739 -25426 32755 -25409
rect 32975 -25409 33065 -25392
rect 33123 -25392 33523 -25345
rect 33123 -25409 33213 -25392
rect 32975 -25426 32991 -25409
rect 32739 -25442 32991 -25426
rect 33197 -25426 33213 -25409
rect 33433 -25409 33523 -25392
rect 33581 -25392 33981 -25345
rect 33581 -25409 33671 -25392
rect 33433 -25426 33449 -25409
rect 33197 -25442 33449 -25426
rect 33655 -25426 33671 -25409
rect 33891 -25409 33981 -25392
rect 34039 -25392 34439 -25345
rect 34039 -25409 34129 -25392
rect 33891 -25426 33907 -25409
rect 33655 -25442 33907 -25426
rect 34113 -25426 34129 -25409
rect 34349 -25409 34439 -25392
rect 34497 -25392 34897 -25345
rect 34497 -25409 34587 -25392
rect 34349 -25426 34365 -25409
rect 34113 -25442 34365 -25426
rect 34571 -25426 34587 -25409
rect 34807 -25409 34897 -25392
rect 34955 -25392 35355 -25345
rect 34955 -25409 35045 -25392
rect 34807 -25426 34823 -25409
rect 34571 -25442 34823 -25426
rect 35029 -25426 35045 -25409
rect 35265 -25409 35355 -25392
rect 35413 -25392 35813 -25345
rect 35413 -25409 35503 -25392
rect 35265 -25426 35281 -25409
rect 35029 -25442 35281 -25426
rect 35487 -25426 35503 -25409
rect 35723 -25409 35813 -25392
rect 35723 -25426 35739 -25409
rect 35487 -25442 35739 -25426
rect 11364 -26566 11616 -26550
rect 11364 -26583 11380 -26566
rect 11290 -26600 11380 -26583
rect 11600 -26583 11616 -26566
rect 11822 -26566 12074 -26550
rect 11822 -26583 11838 -26566
rect 11600 -26600 11690 -26583
rect 11290 -26638 11690 -26600
rect 11748 -26600 11838 -26583
rect 12058 -26583 12074 -26566
rect 12280 -26566 12532 -26550
rect 12280 -26583 12296 -26566
rect 12058 -26600 12148 -26583
rect 11748 -26638 12148 -26600
rect 12206 -26600 12296 -26583
rect 12516 -26583 12532 -26566
rect 12738 -26566 12990 -26550
rect 12738 -26583 12754 -26566
rect 12516 -26600 12606 -26583
rect 12206 -26638 12606 -26600
rect 12664 -26600 12754 -26583
rect 12974 -26583 12990 -26566
rect 13196 -26566 13448 -26550
rect 13196 -26583 13212 -26566
rect 12974 -26600 13064 -26583
rect 12664 -26638 13064 -26600
rect 13122 -26600 13212 -26583
rect 13432 -26583 13448 -26566
rect 13654 -26566 13906 -26550
rect 13654 -26583 13670 -26566
rect 13432 -26600 13522 -26583
rect 13122 -26638 13522 -26600
rect 13580 -26600 13670 -26583
rect 13890 -26583 13906 -26566
rect 14112 -26566 14364 -26550
rect 14112 -26583 14128 -26566
rect 13890 -26600 13980 -26583
rect 13580 -26638 13980 -26600
rect 14038 -26600 14128 -26583
rect 14348 -26583 14364 -26566
rect 14570 -26566 14822 -26550
rect 14570 -26583 14586 -26566
rect 14348 -26600 14438 -26583
rect 14038 -26638 14438 -26600
rect 14496 -26600 14586 -26583
rect 14806 -26583 14822 -26566
rect 15028 -26566 15280 -26550
rect 15028 -26583 15044 -26566
rect 14806 -26600 14896 -26583
rect 14496 -26638 14896 -26600
rect 14954 -26600 15044 -26583
rect 15264 -26583 15280 -26566
rect 15486 -26566 15738 -26550
rect 15486 -26583 15502 -26566
rect 15264 -26600 15354 -26583
rect 14954 -26638 15354 -26600
rect 15412 -26600 15502 -26583
rect 15722 -26583 15738 -26566
rect 16364 -26566 16616 -26550
rect 16364 -26583 16380 -26566
rect 15722 -26600 15812 -26583
rect 15412 -26638 15812 -26600
rect 16290 -26600 16380 -26583
rect 16600 -26583 16616 -26566
rect 16822 -26566 17074 -26550
rect 16822 -26583 16838 -26566
rect 16600 -26600 16690 -26583
rect 16290 -26638 16690 -26600
rect 16748 -26600 16838 -26583
rect 17058 -26583 17074 -26566
rect 17280 -26566 17532 -26550
rect 17280 -26583 17296 -26566
rect 17058 -26600 17148 -26583
rect 16748 -26638 17148 -26600
rect 17206 -26600 17296 -26583
rect 17516 -26583 17532 -26566
rect 17738 -26566 17990 -26550
rect 17738 -26583 17754 -26566
rect 17516 -26600 17606 -26583
rect 17206 -26638 17606 -26600
rect 17664 -26600 17754 -26583
rect 17974 -26583 17990 -26566
rect 18196 -26566 18448 -26550
rect 18196 -26583 18212 -26566
rect 17974 -26600 18064 -26583
rect 17664 -26638 18064 -26600
rect 18122 -26600 18212 -26583
rect 18432 -26583 18448 -26566
rect 18654 -26566 18906 -26550
rect 18654 -26583 18670 -26566
rect 18432 -26600 18522 -26583
rect 18122 -26638 18522 -26600
rect 18580 -26600 18670 -26583
rect 18890 -26583 18906 -26566
rect 19112 -26566 19364 -26550
rect 19112 -26583 19128 -26566
rect 18890 -26600 18980 -26583
rect 18580 -26638 18980 -26600
rect 19038 -26600 19128 -26583
rect 19348 -26583 19364 -26566
rect 19570 -26566 19822 -26550
rect 19570 -26583 19586 -26566
rect 19348 -26600 19438 -26583
rect 19038 -26638 19438 -26600
rect 19496 -26600 19586 -26583
rect 19806 -26583 19822 -26566
rect 20028 -26566 20280 -26550
rect 20028 -26583 20044 -26566
rect 19806 -26600 19896 -26583
rect 19496 -26638 19896 -26600
rect 19954 -26600 20044 -26583
rect 20264 -26583 20280 -26566
rect 20486 -26566 20738 -26550
rect 20486 -26583 20502 -26566
rect 20264 -26600 20354 -26583
rect 19954 -26638 20354 -26600
rect 20412 -26600 20502 -26583
rect 20722 -26583 20738 -26566
rect 20722 -26600 20812 -26583
rect 20412 -26638 20812 -26600
rect 11290 -26876 11690 -26838
rect 11290 -26893 11380 -26876
rect 11364 -26910 11380 -26893
rect 11600 -26893 11690 -26876
rect 11748 -26876 12148 -26838
rect 11748 -26893 11838 -26876
rect 11600 -26910 11616 -26893
rect 11364 -26926 11616 -26910
rect 11822 -26910 11838 -26893
rect 12058 -26893 12148 -26876
rect 12206 -26876 12606 -26838
rect 12206 -26893 12296 -26876
rect 12058 -26910 12074 -26893
rect 11822 -26926 12074 -26910
rect 12280 -26910 12296 -26893
rect 12516 -26893 12606 -26876
rect 12664 -26876 13064 -26838
rect 12664 -26893 12754 -26876
rect 12516 -26910 12532 -26893
rect 12280 -26926 12532 -26910
rect 12738 -26910 12754 -26893
rect 12974 -26893 13064 -26876
rect 13122 -26876 13522 -26838
rect 13122 -26893 13212 -26876
rect 12974 -26910 12990 -26893
rect 12738 -26926 12990 -26910
rect 13196 -26910 13212 -26893
rect 13432 -26893 13522 -26876
rect 13580 -26876 13980 -26838
rect 13580 -26893 13670 -26876
rect 13432 -26910 13448 -26893
rect 13196 -26926 13448 -26910
rect 13654 -26910 13670 -26893
rect 13890 -26893 13980 -26876
rect 14038 -26876 14438 -26838
rect 14038 -26893 14128 -26876
rect 13890 -26910 13906 -26893
rect 13654 -26926 13906 -26910
rect 14112 -26910 14128 -26893
rect 14348 -26893 14438 -26876
rect 14496 -26876 14896 -26838
rect 14496 -26893 14586 -26876
rect 14348 -26910 14364 -26893
rect 14112 -26926 14364 -26910
rect 14570 -26910 14586 -26893
rect 14806 -26893 14896 -26876
rect 14954 -26876 15354 -26838
rect 14954 -26893 15044 -26876
rect 14806 -26910 14822 -26893
rect 14570 -26926 14822 -26910
rect 15028 -26910 15044 -26893
rect 15264 -26893 15354 -26876
rect 15412 -26876 15812 -26838
rect 15412 -26893 15502 -26876
rect 15264 -26910 15280 -26893
rect 15028 -26926 15280 -26910
rect 15486 -26910 15502 -26893
rect 15722 -26893 15812 -26876
rect 16290 -26876 16690 -26838
rect 16290 -26893 16380 -26876
rect 15722 -26910 15738 -26893
rect 15486 -26926 15738 -26910
rect 16364 -26910 16380 -26893
rect 16600 -26893 16690 -26876
rect 16748 -26876 17148 -26838
rect 16748 -26893 16838 -26876
rect 16600 -26910 16616 -26893
rect 16364 -26926 16616 -26910
rect 16822 -26910 16838 -26893
rect 17058 -26893 17148 -26876
rect 17206 -26876 17606 -26838
rect 17206 -26893 17296 -26876
rect 17058 -26910 17074 -26893
rect 16822 -26926 17074 -26910
rect 17280 -26910 17296 -26893
rect 17516 -26893 17606 -26876
rect 17664 -26876 18064 -26838
rect 17664 -26893 17754 -26876
rect 17516 -26910 17532 -26893
rect 17280 -26926 17532 -26910
rect 17738 -26910 17754 -26893
rect 17974 -26893 18064 -26876
rect 18122 -26876 18522 -26838
rect 18122 -26893 18212 -26876
rect 17974 -26910 17990 -26893
rect 17738 -26926 17990 -26910
rect 18196 -26910 18212 -26893
rect 18432 -26893 18522 -26876
rect 18580 -26876 18980 -26838
rect 18580 -26893 18670 -26876
rect 18432 -26910 18448 -26893
rect 18196 -26926 18448 -26910
rect 18654 -26910 18670 -26893
rect 18890 -26893 18980 -26876
rect 19038 -26876 19438 -26838
rect 19038 -26893 19128 -26876
rect 18890 -26910 18906 -26893
rect 18654 -26926 18906 -26910
rect 19112 -26910 19128 -26893
rect 19348 -26893 19438 -26876
rect 19496 -26876 19896 -26838
rect 19496 -26893 19586 -26876
rect 19348 -26910 19364 -26893
rect 19112 -26926 19364 -26910
rect 19570 -26910 19586 -26893
rect 19806 -26893 19896 -26876
rect 19954 -26876 20354 -26838
rect 19954 -26893 20044 -26876
rect 19806 -26910 19822 -26893
rect 19570 -26926 19822 -26910
rect 20028 -26910 20044 -26893
rect 20264 -26893 20354 -26876
rect 20412 -26876 20812 -26838
rect 20412 -26893 20502 -26876
rect 20264 -26910 20280 -26893
rect 20028 -26926 20280 -26910
rect 20486 -26910 20502 -26893
rect 20722 -26893 20812 -26876
rect 20722 -26910 20738 -26893
rect 20486 -26926 20738 -26910
rect 11364 -27234 11616 -27218
rect 11364 -27251 11380 -27234
rect 11290 -27268 11380 -27251
rect 11600 -27251 11616 -27234
rect 11822 -27234 12074 -27218
rect 11822 -27251 11838 -27234
rect 11600 -27268 11690 -27251
rect 11290 -27306 11690 -27268
rect 11748 -27268 11838 -27251
rect 12058 -27251 12074 -27234
rect 12280 -27234 12532 -27218
rect 12280 -27251 12296 -27234
rect 12058 -27268 12148 -27251
rect 11748 -27306 12148 -27268
rect 12206 -27268 12296 -27251
rect 12516 -27251 12532 -27234
rect 12738 -27234 12990 -27218
rect 12738 -27251 12754 -27234
rect 12516 -27268 12606 -27251
rect 12206 -27306 12606 -27268
rect 12664 -27268 12754 -27251
rect 12974 -27251 12990 -27234
rect 13196 -27234 13448 -27218
rect 13196 -27251 13212 -27234
rect 12974 -27268 13064 -27251
rect 12664 -27306 13064 -27268
rect 13122 -27268 13212 -27251
rect 13432 -27251 13448 -27234
rect 13654 -27234 13906 -27218
rect 13654 -27251 13670 -27234
rect 13432 -27268 13522 -27251
rect 13122 -27306 13522 -27268
rect 13580 -27268 13670 -27251
rect 13890 -27251 13906 -27234
rect 14112 -27234 14364 -27218
rect 14112 -27251 14128 -27234
rect 13890 -27268 13980 -27251
rect 13580 -27306 13980 -27268
rect 14038 -27268 14128 -27251
rect 14348 -27251 14364 -27234
rect 14570 -27234 14822 -27218
rect 14570 -27251 14586 -27234
rect 14348 -27268 14438 -27251
rect 14038 -27306 14438 -27268
rect 14496 -27268 14586 -27251
rect 14806 -27251 14822 -27234
rect 15028 -27234 15280 -27218
rect 15028 -27251 15044 -27234
rect 14806 -27268 14896 -27251
rect 14496 -27306 14896 -27268
rect 14954 -27268 15044 -27251
rect 15264 -27251 15280 -27234
rect 15486 -27234 15738 -27218
rect 15486 -27251 15502 -27234
rect 15264 -27268 15354 -27251
rect 14954 -27306 15354 -27268
rect 15412 -27268 15502 -27251
rect 15722 -27251 15738 -27234
rect 15722 -27268 15812 -27251
rect 15412 -27306 15812 -27268
rect 11290 -27544 11690 -27506
rect 11290 -27561 11380 -27544
rect 11364 -27578 11380 -27561
rect 11600 -27561 11690 -27544
rect 11748 -27544 12148 -27506
rect 11748 -27561 11838 -27544
rect 11600 -27578 11616 -27561
rect 11364 -27594 11616 -27578
rect 11822 -27578 11838 -27561
rect 12058 -27561 12148 -27544
rect 12206 -27544 12606 -27506
rect 12206 -27561 12296 -27544
rect 12058 -27578 12074 -27561
rect 11822 -27594 12074 -27578
rect 12280 -27578 12296 -27561
rect 12516 -27561 12606 -27544
rect 12664 -27544 13064 -27506
rect 12664 -27561 12754 -27544
rect 12516 -27578 12532 -27561
rect 12280 -27594 12532 -27578
rect 12738 -27578 12754 -27561
rect 12974 -27561 13064 -27544
rect 13122 -27544 13522 -27506
rect 13122 -27561 13212 -27544
rect 12974 -27578 12990 -27561
rect 12738 -27594 12990 -27578
rect 13196 -27578 13212 -27561
rect 13432 -27561 13522 -27544
rect 13580 -27544 13980 -27506
rect 13580 -27561 13670 -27544
rect 13432 -27578 13448 -27561
rect 13196 -27594 13448 -27578
rect 13654 -27578 13670 -27561
rect 13890 -27561 13980 -27544
rect 14038 -27544 14438 -27506
rect 14038 -27561 14128 -27544
rect 13890 -27578 13906 -27561
rect 13654 -27594 13906 -27578
rect 14112 -27578 14128 -27561
rect 14348 -27561 14438 -27544
rect 14496 -27544 14896 -27506
rect 14496 -27561 14586 -27544
rect 14348 -27578 14364 -27561
rect 14112 -27594 14364 -27578
rect 14570 -27578 14586 -27561
rect 14806 -27561 14896 -27544
rect 14954 -27544 15354 -27506
rect 14954 -27561 15044 -27544
rect 14806 -27578 14822 -27561
rect 14570 -27594 14822 -27578
rect 15028 -27578 15044 -27561
rect 15264 -27561 15354 -27544
rect 15412 -27544 15812 -27506
rect 15412 -27561 15502 -27544
rect 15264 -27578 15280 -27561
rect 15028 -27594 15280 -27578
rect 15486 -27578 15502 -27561
rect 15722 -27561 15812 -27544
rect 15722 -27578 15738 -27561
rect 15486 -27594 15738 -27578
rect 26364 -26566 26616 -26550
rect 26364 -26583 26380 -26566
rect 26290 -26600 26380 -26583
rect 26600 -26583 26616 -26566
rect 26822 -26566 27074 -26550
rect 26822 -26583 26838 -26566
rect 26600 -26600 26690 -26583
rect 26290 -26638 26690 -26600
rect 26748 -26600 26838 -26583
rect 27058 -26583 27074 -26566
rect 27280 -26566 27532 -26550
rect 27280 -26583 27296 -26566
rect 27058 -26600 27148 -26583
rect 26748 -26638 27148 -26600
rect 27206 -26600 27296 -26583
rect 27516 -26583 27532 -26566
rect 27738 -26566 27990 -26550
rect 27738 -26583 27754 -26566
rect 27516 -26600 27606 -26583
rect 27206 -26638 27606 -26600
rect 27664 -26600 27754 -26583
rect 27974 -26583 27990 -26566
rect 28196 -26566 28448 -26550
rect 28196 -26583 28212 -26566
rect 27974 -26600 28064 -26583
rect 27664 -26638 28064 -26600
rect 28122 -26600 28212 -26583
rect 28432 -26583 28448 -26566
rect 28654 -26566 28906 -26550
rect 28654 -26583 28670 -26566
rect 28432 -26600 28522 -26583
rect 28122 -26638 28522 -26600
rect 28580 -26600 28670 -26583
rect 28890 -26583 28906 -26566
rect 29112 -26566 29364 -26550
rect 29112 -26583 29128 -26566
rect 28890 -26600 28980 -26583
rect 28580 -26638 28980 -26600
rect 29038 -26600 29128 -26583
rect 29348 -26583 29364 -26566
rect 29570 -26566 29822 -26550
rect 29570 -26583 29586 -26566
rect 29348 -26600 29438 -26583
rect 29038 -26638 29438 -26600
rect 29496 -26600 29586 -26583
rect 29806 -26583 29822 -26566
rect 30028 -26566 30280 -26550
rect 30028 -26583 30044 -26566
rect 29806 -26600 29896 -26583
rect 29496 -26638 29896 -26600
rect 29954 -26600 30044 -26583
rect 30264 -26583 30280 -26566
rect 30486 -26566 30738 -26550
rect 30486 -26583 30502 -26566
rect 30264 -26600 30354 -26583
rect 29954 -26638 30354 -26600
rect 30412 -26600 30502 -26583
rect 30722 -26583 30738 -26566
rect 31364 -26566 31616 -26550
rect 31364 -26583 31380 -26566
rect 30722 -26600 30812 -26583
rect 30412 -26638 30812 -26600
rect 31290 -26600 31380 -26583
rect 31600 -26583 31616 -26566
rect 31822 -26566 32074 -26550
rect 31822 -26583 31838 -26566
rect 31600 -26600 31690 -26583
rect 31290 -26638 31690 -26600
rect 31748 -26600 31838 -26583
rect 32058 -26583 32074 -26566
rect 32280 -26566 32532 -26550
rect 32280 -26583 32296 -26566
rect 32058 -26600 32148 -26583
rect 31748 -26638 32148 -26600
rect 32206 -26600 32296 -26583
rect 32516 -26583 32532 -26566
rect 32738 -26566 32990 -26550
rect 32738 -26583 32754 -26566
rect 32516 -26600 32606 -26583
rect 32206 -26638 32606 -26600
rect 32664 -26600 32754 -26583
rect 32974 -26583 32990 -26566
rect 33196 -26566 33448 -26550
rect 33196 -26583 33212 -26566
rect 32974 -26600 33064 -26583
rect 32664 -26638 33064 -26600
rect 33122 -26600 33212 -26583
rect 33432 -26583 33448 -26566
rect 33654 -26566 33906 -26550
rect 33654 -26583 33670 -26566
rect 33432 -26600 33522 -26583
rect 33122 -26638 33522 -26600
rect 33580 -26600 33670 -26583
rect 33890 -26583 33906 -26566
rect 34112 -26566 34364 -26550
rect 34112 -26583 34128 -26566
rect 33890 -26600 33980 -26583
rect 33580 -26638 33980 -26600
rect 34038 -26600 34128 -26583
rect 34348 -26583 34364 -26566
rect 34570 -26566 34822 -26550
rect 34570 -26583 34586 -26566
rect 34348 -26600 34438 -26583
rect 34038 -26638 34438 -26600
rect 34496 -26600 34586 -26583
rect 34806 -26583 34822 -26566
rect 35028 -26566 35280 -26550
rect 35028 -26583 35044 -26566
rect 34806 -26600 34896 -26583
rect 34496 -26638 34896 -26600
rect 34954 -26600 35044 -26583
rect 35264 -26583 35280 -26566
rect 35486 -26566 35738 -26550
rect 35486 -26583 35502 -26566
rect 35264 -26600 35354 -26583
rect 34954 -26638 35354 -26600
rect 35412 -26600 35502 -26583
rect 35722 -26583 35738 -26566
rect 35722 -26600 35812 -26583
rect 35412 -26638 35812 -26600
rect 26290 -26876 26690 -26838
rect 26290 -26893 26380 -26876
rect 26364 -26910 26380 -26893
rect 26600 -26893 26690 -26876
rect 26748 -26876 27148 -26838
rect 26748 -26893 26838 -26876
rect 26600 -26910 26616 -26893
rect 26364 -26926 26616 -26910
rect 26822 -26910 26838 -26893
rect 27058 -26893 27148 -26876
rect 27206 -26876 27606 -26838
rect 27206 -26893 27296 -26876
rect 27058 -26910 27074 -26893
rect 26822 -26926 27074 -26910
rect 27280 -26910 27296 -26893
rect 27516 -26893 27606 -26876
rect 27664 -26876 28064 -26838
rect 27664 -26893 27754 -26876
rect 27516 -26910 27532 -26893
rect 27280 -26926 27532 -26910
rect 27738 -26910 27754 -26893
rect 27974 -26893 28064 -26876
rect 28122 -26876 28522 -26838
rect 28122 -26893 28212 -26876
rect 27974 -26910 27990 -26893
rect 27738 -26926 27990 -26910
rect 28196 -26910 28212 -26893
rect 28432 -26893 28522 -26876
rect 28580 -26876 28980 -26838
rect 28580 -26893 28670 -26876
rect 28432 -26910 28448 -26893
rect 28196 -26926 28448 -26910
rect 28654 -26910 28670 -26893
rect 28890 -26893 28980 -26876
rect 29038 -26876 29438 -26838
rect 29038 -26893 29128 -26876
rect 28890 -26910 28906 -26893
rect 28654 -26926 28906 -26910
rect 29112 -26910 29128 -26893
rect 29348 -26893 29438 -26876
rect 29496 -26876 29896 -26838
rect 29496 -26893 29586 -26876
rect 29348 -26910 29364 -26893
rect 29112 -26926 29364 -26910
rect 29570 -26910 29586 -26893
rect 29806 -26893 29896 -26876
rect 29954 -26876 30354 -26838
rect 29954 -26893 30044 -26876
rect 29806 -26910 29822 -26893
rect 29570 -26926 29822 -26910
rect 30028 -26910 30044 -26893
rect 30264 -26893 30354 -26876
rect 30412 -26876 30812 -26838
rect 30412 -26893 30502 -26876
rect 30264 -26910 30280 -26893
rect 30028 -26926 30280 -26910
rect 30486 -26910 30502 -26893
rect 30722 -26893 30812 -26876
rect 31290 -26876 31690 -26838
rect 31290 -26893 31380 -26876
rect 30722 -26910 30738 -26893
rect 30486 -26926 30738 -26910
rect 31364 -26910 31380 -26893
rect 31600 -26893 31690 -26876
rect 31748 -26876 32148 -26838
rect 31748 -26893 31838 -26876
rect 31600 -26910 31616 -26893
rect 31364 -26926 31616 -26910
rect 31822 -26910 31838 -26893
rect 32058 -26893 32148 -26876
rect 32206 -26876 32606 -26838
rect 32206 -26893 32296 -26876
rect 32058 -26910 32074 -26893
rect 31822 -26926 32074 -26910
rect 32280 -26910 32296 -26893
rect 32516 -26893 32606 -26876
rect 32664 -26876 33064 -26838
rect 32664 -26893 32754 -26876
rect 32516 -26910 32532 -26893
rect 32280 -26926 32532 -26910
rect 32738 -26910 32754 -26893
rect 32974 -26893 33064 -26876
rect 33122 -26876 33522 -26838
rect 33122 -26893 33212 -26876
rect 32974 -26910 32990 -26893
rect 32738 -26926 32990 -26910
rect 33196 -26910 33212 -26893
rect 33432 -26893 33522 -26876
rect 33580 -26876 33980 -26838
rect 33580 -26893 33670 -26876
rect 33432 -26910 33448 -26893
rect 33196 -26926 33448 -26910
rect 33654 -26910 33670 -26893
rect 33890 -26893 33980 -26876
rect 34038 -26876 34438 -26838
rect 34038 -26893 34128 -26876
rect 33890 -26910 33906 -26893
rect 33654 -26926 33906 -26910
rect 34112 -26910 34128 -26893
rect 34348 -26893 34438 -26876
rect 34496 -26876 34896 -26838
rect 34496 -26893 34586 -26876
rect 34348 -26910 34364 -26893
rect 34112 -26926 34364 -26910
rect 34570 -26910 34586 -26893
rect 34806 -26893 34896 -26876
rect 34954 -26876 35354 -26838
rect 34954 -26893 35044 -26876
rect 34806 -26910 34822 -26893
rect 34570 -26926 34822 -26910
rect 35028 -26910 35044 -26893
rect 35264 -26893 35354 -26876
rect 35412 -26876 35812 -26838
rect 35412 -26893 35502 -26876
rect 35264 -26910 35280 -26893
rect 35028 -26926 35280 -26910
rect 35486 -26910 35502 -26893
rect 35722 -26893 35812 -26876
rect 35722 -26910 35738 -26893
rect 35486 -26926 35738 -26910
rect 26364 -27234 26616 -27218
rect 26364 -27251 26380 -27234
rect 26290 -27268 26380 -27251
rect 26600 -27251 26616 -27234
rect 26822 -27234 27074 -27218
rect 26822 -27251 26838 -27234
rect 26600 -27268 26690 -27251
rect 26290 -27306 26690 -27268
rect 26748 -27268 26838 -27251
rect 27058 -27251 27074 -27234
rect 27280 -27234 27532 -27218
rect 27280 -27251 27296 -27234
rect 27058 -27268 27148 -27251
rect 26748 -27306 27148 -27268
rect 27206 -27268 27296 -27251
rect 27516 -27251 27532 -27234
rect 27738 -27234 27990 -27218
rect 27738 -27251 27754 -27234
rect 27516 -27268 27606 -27251
rect 27206 -27306 27606 -27268
rect 27664 -27268 27754 -27251
rect 27974 -27251 27990 -27234
rect 28196 -27234 28448 -27218
rect 28196 -27251 28212 -27234
rect 27974 -27268 28064 -27251
rect 27664 -27306 28064 -27268
rect 28122 -27268 28212 -27251
rect 28432 -27251 28448 -27234
rect 28654 -27234 28906 -27218
rect 28654 -27251 28670 -27234
rect 28432 -27268 28522 -27251
rect 28122 -27306 28522 -27268
rect 28580 -27268 28670 -27251
rect 28890 -27251 28906 -27234
rect 29112 -27234 29364 -27218
rect 29112 -27251 29128 -27234
rect 28890 -27268 28980 -27251
rect 28580 -27306 28980 -27268
rect 29038 -27268 29128 -27251
rect 29348 -27251 29364 -27234
rect 29570 -27234 29822 -27218
rect 29570 -27251 29586 -27234
rect 29348 -27268 29438 -27251
rect 29038 -27306 29438 -27268
rect 29496 -27268 29586 -27251
rect 29806 -27251 29822 -27234
rect 30028 -27234 30280 -27218
rect 30028 -27251 30044 -27234
rect 29806 -27268 29896 -27251
rect 29496 -27306 29896 -27268
rect 29954 -27268 30044 -27251
rect 30264 -27251 30280 -27234
rect 30486 -27234 30738 -27218
rect 30486 -27251 30502 -27234
rect 30264 -27268 30354 -27251
rect 29954 -27306 30354 -27268
rect 30412 -27268 30502 -27251
rect 30722 -27251 30738 -27234
rect 30722 -27268 30812 -27251
rect 30412 -27306 30812 -27268
rect 26290 -27544 26690 -27506
rect 26290 -27561 26380 -27544
rect 26364 -27578 26380 -27561
rect 26600 -27561 26690 -27544
rect 26748 -27544 27148 -27506
rect 26748 -27561 26838 -27544
rect 26600 -27578 26616 -27561
rect 26364 -27594 26616 -27578
rect 26822 -27578 26838 -27561
rect 27058 -27561 27148 -27544
rect 27206 -27544 27606 -27506
rect 27206 -27561 27296 -27544
rect 27058 -27578 27074 -27561
rect 26822 -27594 27074 -27578
rect 27280 -27578 27296 -27561
rect 27516 -27561 27606 -27544
rect 27664 -27544 28064 -27506
rect 27664 -27561 27754 -27544
rect 27516 -27578 27532 -27561
rect 27280 -27594 27532 -27578
rect 27738 -27578 27754 -27561
rect 27974 -27561 28064 -27544
rect 28122 -27544 28522 -27506
rect 28122 -27561 28212 -27544
rect 27974 -27578 27990 -27561
rect 27738 -27594 27990 -27578
rect 28196 -27578 28212 -27561
rect 28432 -27561 28522 -27544
rect 28580 -27544 28980 -27506
rect 28580 -27561 28670 -27544
rect 28432 -27578 28448 -27561
rect 28196 -27594 28448 -27578
rect 28654 -27578 28670 -27561
rect 28890 -27561 28980 -27544
rect 29038 -27544 29438 -27506
rect 29038 -27561 29128 -27544
rect 28890 -27578 28906 -27561
rect 28654 -27594 28906 -27578
rect 29112 -27578 29128 -27561
rect 29348 -27561 29438 -27544
rect 29496 -27544 29896 -27506
rect 29496 -27561 29586 -27544
rect 29348 -27578 29364 -27561
rect 29112 -27594 29364 -27578
rect 29570 -27578 29586 -27561
rect 29806 -27561 29896 -27544
rect 29954 -27544 30354 -27506
rect 29954 -27561 30044 -27544
rect 29806 -27578 29822 -27561
rect 29570 -27594 29822 -27578
rect 30028 -27578 30044 -27561
rect 30264 -27561 30354 -27544
rect 30412 -27544 30812 -27506
rect 30412 -27561 30502 -27544
rect 30264 -27578 30280 -27561
rect 30028 -27594 30280 -27578
rect 30486 -27578 30502 -27561
rect 30722 -27561 30812 -27544
rect 30722 -27578 30738 -27561
rect 30486 -27594 30738 -27578
<< polycont >>
rect 17770 3282 17990 3316
rect 18228 3282 18448 3316
rect 18686 3282 18906 3316
rect 19144 3282 19364 3316
rect 19602 3282 19822 3316
rect 20060 3282 20280 3316
rect 20518 3282 20738 3316
rect 20976 3282 21196 3316
rect 21434 3282 21654 3316
rect 21892 3282 22112 3316
rect 17770 2972 17990 3006
rect 18228 2972 18448 3006
rect 18686 2972 18906 3006
rect 19144 2972 19364 3006
rect 19602 2972 19822 3006
rect 20060 2972 20280 3006
rect 20518 2972 20738 3006
rect 20976 2972 21196 3006
rect 21434 2972 21654 3006
rect 21892 2972 22112 3006
rect 26532 3282 26752 3316
rect 26990 3282 27210 3316
rect 27448 3282 27668 3316
rect 27906 3282 28126 3316
rect 28364 3282 28584 3316
rect 28822 3282 29042 3316
rect 29280 3282 29500 3316
rect 29738 3282 29958 3316
rect 30196 3282 30416 3316
rect 30654 3282 30874 3316
rect 26532 2972 26752 3006
rect 26990 2972 27210 3006
rect 27448 2972 27668 3006
rect 27906 2972 28126 3006
rect 28364 2972 28584 3006
rect 28822 2972 29042 3006
rect 29280 2972 29500 3006
rect 29738 2972 29958 3006
rect 30196 2972 30416 3006
rect 30654 2972 30874 3006
rect 31622 2241 31656 2275
rect 31855 2241 31889 2275
rect 31947 2241 31981 2275
rect 32031 2241 32065 2275
rect 32115 2241 32149 2275
rect 15938 1440 16158 1474
rect 16396 1440 16616 1474
rect 16854 1440 17074 1474
rect 17312 1440 17532 1474
rect 17770 1440 17990 1474
rect 18228 1440 18448 1474
rect 18686 1440 18906 1474
rect 19144 1440 19364 1474
rect 19602 1440 19822 1474
rect 20060 1440 20280 1474
rect 20518 1440 20738 1474
rect 20976 1440 21196 1474
rect 21434 1440 21654 1474
rect 21892 1440 22112 1474
rect 22350 1440 22570 1474
rect 22808 1440 23028 1474
rect 23266 1440 23486 1474
rect 23724 1440 23944 1474
rect 15938 -288 16158 -254
rect 16396 -288 16616 -254
rect 16854 -288 17074 -254
rect 17312 -288 17532 -254
rect 17770 -288 17990 -254
rect 18228 -288 18448 -254
rect 18686 -288 18906 -254
rect 19144 -288 19364 -254
rect 19602 -288 19822 -254
rect 20060 -288 20280 -254
rect 20518 -288 20738 -254
rect 20976 -288 21196 -254
rect 21434 -288 21654 -254
rect 21892 -288 22112 -254
rect 22350 -288 22570 -254
rect 22808 -288 23028 -254
rect 23266 -288 23486 -254
rect 23724 -288 23944 -254
rect 26533 1860 26753 1894
rect 26991 1860 27211 1894
rect 27449 1860 27669 1894
rect 27907 1860 28127 1894
rect 28365 1860 28585 1894
rect 28823 1860 29043 1894
rect 29281 1860 29501 1894
rect 29739 1860 29959 1894
rect 30197 1860 30417 1894
rect 30655 1860 30875 1894
rect 26533 532 26753 566
rect 26991 532 27211 566
rect 27449 532 27669 566
rect 27907 532 28127 566
rect 28365 532 28585 566
rect 28823 532 29043 566
rect 29281 532 29501 566
rect 29739 532 29959 566
rect 30197 532 30417 566
rect 30655 532 30875 566
rect 11940 -3433 12160 -3399
rect 12398 -3433 12618 -3399
rect 12856 -3433 13076 -3399
rect 13314 -3433 13534 -3399
rect 13772 -3433 13992 -3399
rect 14230 -3433 14450 -3399
rect 14688 -3433 14908 -3399
rect 15146 -3433 15366 -3399
rect 15604 -3433 15824 -3399
rect 16062 -3433 16282 -3399
rect 16520 -3433 16740 -3399
rect 16978 -3433 17198 -3399
rect 17436 -3433 17656 -3399
rect 17894 -3433 18114 -3399
rect 18352 -3433 18572 -3399
rect 18810 -3433 19030 -3399
rect 19268 -3433 19488 -3399
rect 19726 -3433 19946 -3399
rect 11940 -5161 12160 -5127
rect 12398 -5161 12618 -5127
rect 12856 -5161 13076 -5127
rect 13314 -5161 13534 -5127
rect 13772 -5161 13992 -5127
rect 14230 -5161 14450 -5127
rect 14688 -5161 14908 -5127
rect 15146 -5161 15366 -5127
rect 15604 -5161 15824 -5127
rect 16062 -5161 16282 -5127
rect 16520 -5161 16740 -5127
rect 16978 -5161 17198 -5127
rect 17436 -5161 17656 -5127
rect 17894 -5161 18114 -5127
rect 18352 -5161 18572 -5127
rect 18810 -5161 19030 -5127
rect 19268 -5161 19488 -5127
rect 19726 -5161 19946 -5127
rect 11381 -6098 11601 -6064
rect 11839 -6098 12059 -6064
rect 12297 -6098 12517 -6064
rect 12755 -6098 12975 -6064
rect 13213 -6098 13433 -6064
rect 13671 -6098 13891 -6064
rect 14129 -6098 14349 -6064
rect 14587 -6098 14807 -6064
rect 15045 -6098 15265 -6064
rect 15503 -6098 15723 -6064
rect 16381 -6098 16601 -6064
rect 16839 -6098 17059 -6064
rect 17297 -6098 17517 -6064
rect 17755 -6098 17975 -6064
rect 18213 -6098 18433 -6064
rect 18671 -6098 18891 -6064
rect 19129 -6098 19349 -6064
rect 19587 -6098 19807 -6064
rect 20045 -6098 20265 -6064
rect 20503 -6098 20723 -6064
rect 11381 -7426 11601 -7392
rect 11839 -7426 12059 -7392
rect 12297 -7426 12517 -7392
rect 12755 -7426 12975 -7392
rect 13213 -7426 13433 -7392
rect 13671 -7426 13891 -7392
rect 14129 -7426 14349 -7392
rect 14587 -7426 14807 -7392
rect 15045 -7426 15265 -7392
rect 15503 -7426 15723 -7392
rect 16381 -7426 16601 -7392
rect 16839 -7426 17059 -7392
rect 17297 -7426 17517 -7392
rect 17755 -7426 17975 -7392
rect 18213 -7426 18433 -7392
rect 18671 -7426 18891 -7392
rect 19129 -7426 19349 -7392
rect 19587 -7426 19807 -7392
rect 20045 -7426 20265 -7392
rect 20503 -7426 20723 -7392
rect 26940 -3433 27160 -3399
rect 27398 -3433 27618 -3399
rect 27856 -3433 28076 -3399
rect 28314 -3433 28534 -3399
rect 28772 -3433 28992 -3399
rect 29230 -3433 29450 -3399
rect 29688 -3433 29908 -3399
rect 30146 -3433 30366 -3399
rect 30604 -3433 30824 -3399
rect 31062 -3433 31282 -3399
rect 31520 -3433 31740 -3399
rect 31978 -3433 32198 -3399
rect 32436 -3433 32656 -3399
rect 32894 -3433 33114 -3399
rect 33352 -3433 33572 -3399
rect 33810 -3433 34030 -3399
rect 34268 -3433 34488 -3399
rect 34726 -3433 34946 -3399
rect 26940 -5161 27160 -5127
rect 27398 -5161 27618 -5127
rect 27856 -5161 28076 -5127
rect 28314 -5161 28534 -5127
rect 28772 -5161 28992 -5127
rect 29230 -5161 29450 -5127
rect 29688 -5161 29908 -5127
rect 30146 -5161 30366 -5127
rect 30604 -5161 30824 -5127
rect 31062 -5161 31282 -5127
rect 31520 -5161 31740 -5127
rect 31978 -5161 32198 -5127
rect 32436 -5161 32656 -5127
rect 32894 -5161 33114 -5127
rect 33352 -5161 33572 -5127
rect 33810 -5161 34030 -5127
rect 34268 -5161 34488 -5127
rect 34726 -5161 34946 -5127
rect 26381 -6098 26601 -6064
rect 26839 -6098 27059 -6064
rect 27297 -6098 27517 -6064
rect 27755 -6098 27975 -6064
rect 28213 -6098 28433 -6064
rect 28671 -6098 28891 -6064
rect 29129 -6098 29349 -6064
rect 29587 -6098 29807 -6064
rect 30045 -6098 30265 -6064
rect 30503 -6098 30723 -6064
rect 31381 -6098 31601 -6064
rect 31839 -6098 32059 -6064
rect 32297 -6098 32517 -6064
rect 32755 -6098 32975 -6064
rect 33213 -6098 33433 -6064
rect 33671 -6098 33891 -6064
rect 34129 -6098 34349 -6064
rect 34587 -6098 34807 -6064
rect 35045 -6098 35265 -6064
rect 35503 -6098 35723 -6064
rect 26381 -7426 26601 -7392
rect 26839 -7426 27059 -7392
rect 27297 -7426 27517 -7392
rect 27755 -7426 27975 -7392
rect 28213 -7426 28433 -7392
rect 28671 -7426 28891 -7392
rect 29129 -7426 29349 -7392
rect 29587 -7426 29807 -7392
rect 30045 -7426 30265 -7392
rect 30503 -7426 30723 -7392
rect 31381 -7426 31601 -7392
rect 31839 -7426 32059 -7392
rect 32297 -7426 32517 -7392
rect 32755 -7426 32975 -7392
rect 33213 -7426 33433 -7392
rect 33671 -7426 33891 -7392
rect 34129 -7426 34349 -7392
rect 34587 -7426 34807 -7392
rect 35045 -7426 35265 -7392
rect 35503 -7426 35723 -7392
rect 11380 -8600 11600 -8566
rect 11838 -8600 12058 -8566
rect 12296 -8600 12516 -8566
rect 12754 -8600 12974 -8566
rect 13212 -8600 13432 -8566
rect 13670 -8600 13890 -8566
rect 14128 -8600 14348 -8566
rect 14586 -8600 14806 -8566
rect 15044 -8600 15264 -8566
rect 15502 -8600 15722 -8566
rect 16380 -8600 16600 -8566
rect 16838 -8600 17058 -8566
rect 17296 -8600 17516 -8566
rect 17754 -8600 17974 -8566
rect 18212 -8600 18432 -8566
rect 18670 -8600 18890 -8566
rect 19128 -8600 19348 -8566
rect 19586 -8600 19806 -8566
rect 20044 -8600 20264 -8566
rect 20502 -8600 20722 -8566
rect 11380 -8910 11600 -8876
rect 11838 -8910 12058 -8876
rect 12296 -8910 12516 -8876
rect 12754 -8910 12974 -8876
rect 13212 -8910 13432 -8876
rect 13670 -8910 13890 -8876
rect 14128 -8910 14348 -8876
rect 14586 -8910 14806 -8876
rect 15044 -8910 15264 -8876
rect 15502 -8910 15722 -8876
rect 16380 -8910 16600 -8876
rect 16838 -8910 17058 -8876
rect 17296 -8910 17516 -8876
rect 17754 -8910 17974 -8876
rect 18212 -8910 18432 -8876
rect 18670 -8910 18890 -8876
rect 19128 -8910 19348 -8876
rect 19586 -8910 19806 -8876
rect 20044 -8910 20264 -8876
rect 20502 -8910 20722 -8876
rect 11380 -9268 11600 -9234
rect 11838 -9268 12058 -9234
rect 12296 -9268 12516 -9234
rect 12754 -9268 12974 -9234
rect 13212 -9268 13432 -9234
rect 13670 -9268 13890 -9234
rect 14128 -9268 14348 -9234
rect 14586 -9268 14806 -9234
rect 15044 -9268 15264 -9234
rect 15502 -9268 15722 -9234
rect 11380 -9578 11600 -9544
rect 11838 -9578 12058 -9544
rect 12296 -9578 12516 -9544
rect 12754 -9578 12974 -9544
rect 13212 -9578 13432 -9544
rect 13670 -9578 13890 -9544
rect 14128 -9578 14348 -9544
rect 14586 -9578 14806 -9544
rect 15044 -9578 15264 -9544
rect 15502 -9578 15722 -9544
rect 26380 -8600 26600 -8566
rect 26838 -8600 27058 -8566
rect 27296 -8600 27516 -8566
rect 27754 -8600 27974 -8566
rect 28212 -8600 28432 -8566
rect 28670 -8600 28890 -8566
rect 29128 -8600 29348 -8566
rect 29586 -8600 29806 -8566
rect 30044 -8600 30264 -8566
rect 30502 -8600 30722 -8566
rect 31380 -8600 31600 -8566
rect 31838 -8600 32058 -8566
rect 32296 -8600 32516 -8566
rect 32754 -8600 32974 -8566
rect 33212 -8600 33432 -8566
rect 33670 -8600 33890 -8566
rect 34128 -8600 34348 -8566
rect 34586 -8600 34806 -8566
rect 35044 -8600 35264 -8566
rect 35502 -8600 35722 -8566
rect 26380 -8910 26600 -8876
rect 26838 -8910 27058 -8876
rect 27296 -8910 27516 -8876
rect 27754 -8910 27974 -8876
rect 28212 -8910 28432 -8876
rect 28670 -8910 28890 -8876
rect 29128 -8910 29348 -8876
rect 29586 -8910 29806 -8876
rect 30044 -8910 30264 -8876
rect 30502 -8910 30722 -8876
rect 31380 -8910 31600 -8876
rect 31838 -8910 32058 -8876
rect 32296 -8910 32516 -8876
rect 32754 -8910 32974 -8876
rect 33212 -8910 33432 -8876
rect 33670 -8910 33890 -8876
rect 34128 -8910 34348 -8876
rect 34586 -8910 34806 -8876
rect 35044 -8910 35264 -8876
rect 35502 -8910 35722 -8876
rect 26380 -9268 26600 -9234
rect 26838 -9268 27058 -9234
rect 27296 -9268 27516 -9234
rect 27754 -9268 27974 -9234
rect 28212 -9268 28432 -9234
rect 28670 -9268 28890 -9234
rect 29128 -9268 29348 -9234
rect 29586 -9268 29806 -9234
rect 30044 -9268 30264 -9234
rect 30502 -9268 30722 -9234
rect 26380 -9578 26600 -9544
rect 26838 -9578 27058 -9544
rect 27296 -9578 27516 -9544
rect 27754 -9578 27974 -9544
rect 28212 -9578 28432 -9544
rect 28670 -9578 28890 -9544
rect 29128 -9578 29348 -9544
rect 29586 -9578 29806 -9544
rect 30044 -9578 30264 -9544
rect 30502 -9578 30722 -9544
rect 20312 -12060 20532 -12026
rect 20770 -12060 20990 -12026
rect 21228 -12060 21448 -12026
rect 21686 -12060 21906 -12026
rect 22144 -12060 22364 -12026
rect 22602 -12060 22822 -12026
rect 23060 -12060 23280 -12026
rect 23518 -12060 23738 -12026
rect 23976 -12060 24196 -12026
rect 24434 -12060 24654 -12026
rect 20312 -12370 20532 -12336
rect 20770 -12370 20990 -12336
rect 21228 -12370 21448 -12336
rect 21686 -12370 21906 -12336
rect 22144 -12370 22364 -12336
rect 22602 -12370 22822 -12336
rect 23060 -12370 23280 -12336
rect 23518 -12370 23738 -12336
rect 23976 -12370 24196 -12336
rect 24434 -12370 24654 -12336
rect 15312 -12728 15532 -12694
rect 15770 -12728 15990 -12694
rect 16228 -12728 16448 -12694
rect 16686 -12728 16906 -12694
rect 17144 -12728 17364 -12694
rect 17602 -12728 17822 -12694
rect 18060 -12728 18280 -12694
rect 18518 -12728 18738 -12694
rect 18976 -12728 19196 -12694
rect 19434 -12728 19654 -12694
rect 20312 -12728 20532 -12694
rect 20770 -12728 20990 -12694
rect 21228 -12728 21448 -12694
rect 21686 -12728 21906 -12694
rect 22144 -12728 22364 -12694
rect 22602 -12728 22822 -12694
rect 23060 -12728 23280 -12694
rect 23518 -12728 23738 -12694
rect 23976 -12728 24196 -12694
rect 24434 -12728 24654 -12694
rect 15312 -13038 15532 -13004
rect 15770 -13038 15990 -13004
rect 16228 -13038 16448 -13004
rect 16686 -13038 16906 -13004
rect 17144 -13038 17364 -13004
rect 17602 -13038 17822 -13004
rect 18060 -13038 18280 -13004
rect 18518 -13038 18738 -13004
rect 18976 -13038 19196 -13004
rect 19434 -13038 19654 -13004
rect 20312 -13038 20532 -13004
rect 20770 -13038 20990 -13004
rect 21228 -13038 21448 -13004
rect 21686 -13038 21906 -13004
rect 22144 -13038 22364 -13004
rect 22602 -13038 22822 -13004
rect 23060 -13038 23280 -13004
rect 23518 -13038 23738 -13004
rect 23976 -13038 24196 -13004
rect 24434 -13038 24654 -13004
rect 35312 -12060 35532 -12026
rect 35770 -12060 35990 -12026
rect 36228 -12060 36448 -12026
rect 36686 -12060 36906 -12026
rect 37144 -12060 37364 -12026
rect 37602 -12060 37822 -12026
rect 38060 -12060 38280 -12026
rect 38518 -12060 38738 -12026
rect 38976 -12060 39196 -12026
rect 39434 -12060 39654 -12026
rect 35312 -12370 35532 -12336
rect 35770 -12370 35990 -12336
rect 36228 -12370 36448 -12336
rect 36686 -12370 36906 -12336
rect 37144 -12370 37364 -12336
rect 37602 -12370 37822 -12336
rect 38060 -12370 38280 -12336
rect 38518 -12370 38738 -12336
rect 38976 -12370 39196 -12336
rect 39434 -12370 39654 -12336
rect 30312 -12728 30532 -12694
rect 30770 -12728 30990 -12694
rect 31228 -12728 31448 -12694
rect 31686 -12728 31906 -12694
rect 32144 -12728 32364 -12694
rect 32602 -12728 32822 -12694
rect 33060 -12728 33280 -12694
rect 33518 -12728 33738 -12694
rect 33976 -12728 34196 -12694
rect 34434 -12728 34654 -12694
rect 35312 -12728 35532 -12694
rect 35770 -12728 35990 -12694
rect 36228 -12728 36448 -12694
rect 36686 -12728 36906 -12694
rect 37144 -12728 37364 -12694
rect 37602 -12728 37822 -12694
rect 38060 -12728 38280 -12694
rect 38518 -12728 38738 -12694
rect 38976 -12728 39196 -12694
rect 39434 -12728 39654 -12694
rect 30312 -13038 30532 -13004
rect 30770 -13038 30990 -13004
rect 31228 -13038 31448 -13004
rect 31686 -13038 31906 -13004
rect 32144 -13038 32364 -13004
rect 32602 -13038 32822 -13004
rect 33060 -13038 33280 -13004
rect 33518 -13038 33738 -13004
rect 33976 -13038 34196 -13004
rect 34434 -13038 34654 -13004
rect 35312 -13038 35532 -13004
rect 35770 -13038 35990 -13004
rect 36228 -13038 36448 -13004
rect 36686 -13038 36906 -13004
rect 37144 -13038 37364 -13004
rect 37602 -13038 37822 -13004
rect 38060 -13038 38280 -13004
rect 38518 -13038 38738 -13004
rect 38976 -13038 39196 -13004
rect 39434 -13038 39654 -13004
rect 15311 -14212 15531 -14178
rect 15769 -14212 15989 -14178
rect 16227 -14212 16447 -14178
rect 16685 -14212 16905 -14178
rect 17143 -14212 17363 -14178
rect 17601 -14212 17821 -14178
rect 18059 -14212 18279 -14178
rect 18517 -14212 18737 -14178
rect 18975 -14212 19195 -14178
rect 19433 -14212 19653 -14178
rect 20311 -14212 20531 -14178
rect 20769 -14212 20989 -14178
rect 21227 -14212 21447 -14178
rect 21685 -14212 21905 -14178
rect 22143 -14212 22363 -14178
rect 22601 -14212 22821 -14178
rect 23059 -14212 23279 -14178
rect 23517 -14212 23737 -14178
rect 23975 -14212 24195 -14178
rect 24433 -14212 24653 -14178
rect 15311 -15540 15531 -15506
rect 15769 -15540 15989 -15506
rect 16227 -15540 16447 -15506
rect 16685 -15540 16905 -15506
rect 17143 -15540 17363 -15506
rect 17601 -15540 17821 -15506
rect 18059 -15540 18279 -15506
rect 18517 -15540 18737 -15506
rect 18975 -15540 19195 -15506
rect 19433 -15540 19653 -15506
rect 20311 -15540 20531 -15506
rect 20769 -15540 20989 -15506
rect 21227 -15540 21447 -15506
rect 21685 -15540 21905 -15506
rect 22143 -15540 22363 -15506
rect 22601 -15540 22821 -15506
rect 23059 -15540 23279 -15506
rect 23517 -15540 23737 -15506
rect 23975 -15540 24195 -15506
rect 24433 -15540 24653 -15506
rect 16088 -16477 16308 -16443
rect 16546 -16477 16766 -16443
rect 17004 -16477 17224 -16443
rect 17462 -16477 17682 -16443
rect 17920 -16477 18140 -16443
rect 18378 -16477 18598 -16443
rect 18836 -16477 19056 -16443
rect 19294 -16477 19514 -16443
rect 19752 -16477 19972 -16443
rect 20210 -16477 20430 -16443
rect 20668 -16477 20888 -16443
rect 21126 -16477 21346 -16443
rect 21584 -16477 21804 -16443
rect 22042 -16477 22262 -16443
rect 22500 -16477 22720 -16443
rect 22958 -16477 23178 -16443
rect 23416 -16477 23636 -16443
rect 23874 -16477 24094 -16443
rect 16088 -18205 16308 -18171
rect 16546 -18205 16766 -18171
rect 17004 -18205 17224 -18171
rect 17462 -18205 17682 -18171
rect 17920 -18205 18140 -18171
rect 18378 -18205 18598 -18171
rect 18836 -18205 19056 -18171
rect 19294 -18205 19514 -18171
rect 19752 -18205 19972 -18171
rect 20210 -18205 20430 -18171
rect 20668 -18205 20888 -18171
rect 21126 -18205 21346 -18171
rect 21584 -18205 21804 -18171
rect 22042 -18205 22262 -18171
rect 22500 -18205 22720 -18171
rect 22958 -18205 23178 -18171
rect 23416 -18205 23636 -18171
rect 23874 -18205 24094 -18171
rect 30311 -14212 30531 -14178
rect 30769 -14212 30989 -14178
rect 31227 -14212 31447 -14178
rect 31685 -14212 31905 -14178
rect 32143 -14212 32363 -14178
rect 32601 -14212 32821 -14178
rect 33059 -14212 33279 -14178
rect 33517 -14212 33737 -14178
rect 33975 -14212 34195 -14178
rect 34433 -14212 34653 -14178
rect 35311 -14212 35531 -14178
rect 35769 -14212 35989 -14178
rect 36227 -14212 36447 -14178
rect 36685 -14212 36905 -14178
rect 37143 -14212 37363 -14178
rect 37601 -14212 37821 -14178
rect 38059 -14212 38279 -14178
rect 38517 -14212 38737 -14178
rect 38975 -14212 39195 -14178
rect 39433 -14212 39653 -14178
rect 30311 -15540 30531 -15506
rect 30769 -15540 30989 -15506
rect 31227 -15540 31447 -15506
rect 31685 -15540 31905 -15506
rect 32143 -15540 32363 -15506
rect 32601 -15540 32821 -15506
rect 33059 -15540 33279 -15506
rect 33517 -15540 33737 -15506
rect 33975 -15540 34195 -15506
rect 34433 -15540 34653 -15506
rect 35311 -15540 35531 -15506
rect 35769 -15540 35989 -15506
rect 36227 -15540 36447 -15506
rect 36685 -15540 36905 -15506
rect 37143 -15540 37363 -15506
rect 37601 -15540 37821 -15506
rect 38059 -15540 38279 -15506
rect 38517 -15540 38737 -15506
rect 38975 -15540 39195 -15506
rect 39433 -15540 39653 -15506
rect 31088 -16477 31308 -16443
rect 31546 -16477 31766 -16443
rect 32004 -16477 32224 -16443
rect 32462 -16477 32682 -16443
rect 32920 -16477 33140 -16443
rect 33378 -16477 33598 -16443
rect 33836 -16477 34056 -16443
rect 34294 -16477 34514 -16443
rect 34752 -16477 34972 -16443
rect 35210 -16477 35430 -16443
rect 35668 -16477 35888 -16443
rect 36126 -16477 36346 -16443
rect 36584 -16477 36804 -16443
rect 37042 -16477 37262 -16443
rect 37500 -16477 37720 -16443
rect 37958 -16477 38178 -16443
rect 38416 -16477 38636 -16443
rect 38874 -16477 39094 -16443
rect 31088 -18205 31308 -18171
rect 31546 -18205 31766 -18171
rect 32004 -18205 32224 -18171
rect 32462 -18205 32682 -18171
rect 32920 -18205 33140 -18171
rect 33378 -18205 33598 -18171
rect 33836 -18205 34056 -18171
rect 34294 -18205 34514 -18171
rect 34752 -18205 34972 -18171
rect 35210 -18205 35430 -18171
rect 35668 -18205 35888 -18171
rect 36126 -18205 36346 -18171
rect 36584 -18205 36804 -18171
rect 37042 -18205 37262 -18171
rect 37500 -18205 37720 -18171
rect 37958 -18205 38178 -18171
rect 38416 -18205 38636 -18171
rect 38874 -18205 39094 -18171
rect 11940 -21433 12160 -21399
rect 12398 -21433 12618 -21399
rect 12856 -21433 13076 -21399
rect 13314 -21433 13534 -21399
rect 13772 -21433 13992 -21399
rect 14230 -21433 14450 -21399
rect 14688 -21433 14908 -21399
rect 15146 -21433 15366 -21399
rect 15604 -21433 15824 -21399
rect 16062 -21433 16282 -21399
rect 16520 -21433 16740 -21399
rect 16978 -21433 17198 -21399
rect 17436 -21433 17656 -21399
rect 17894 -21433 18114 -21399
rect 18352 -21433 18572 -21399
rect 18810 -21433 19030 -21399
rect 19268 -21433 19488 -21399
rect 19726 -21433 19946 -21399
rect 11940 -23161 12160 -23127
rect 12398 -23161 12618 -23127
rect 12856 -23161 13076 -23127
rect 13314 -23161 13534 -23127
rect 13772 -23161 13992 -23127
rect 14230 -23161 14450 -23127
rect 14688 -23161 14908 -23127
rect 15146 -23161 15366 -23127
rect 15604 -23161 15824 -23127
rect 16062 -23161 16282 -23127
rect 16520 -23161 16740 -23127
rect 16978 -23161 17198 -23127
rect 17436 -23161 17656 -23127
rect 17894 -23161 18114 -23127
rect 18352 -23161 18572 -23127
rect 18810 -23161 19030 -23127
rect 19268 -23161 19488 -23127
rect 19726 -23161 19946 -23127
rect 11381 -24098 11601 -24064
rect 11839 -24098 12059 -24064
rect 12297 -24098 12517 -24064
rect 12755 -24098 12975 -24064
rect 13213 -24098 13433 -24064
rect 13671 -24098 13891 -24064
rect 14129 -24098 14349 -24064
rect 14587 -24098 14807 -24064
rect 15045 -24098 15265 -24064
rect 15503 -24098 15723 -24064
rect 16381 -24098 16601 -24064
rect 16839 -24098 17059 -24064
rect 17297 -24098 17517 -24064
rect 17755 -24098 17975 -24064
rect 18213 -24098 18433 -24064
rect 18671 -24098 18891 -24064
rect 19129 -24098 19349 -24064
rect 19587 -24098 19807 -24064
rect 20045 -24098 20265 -24064
rect 20503 -24098 20723 -24064
rect 11381 -25426 11601 -25392
rect 11839 -25426 12059 -25392
rect 12297 -25426 12517 -25392
rect 12755 -25426 12975 -25392
rect 13213 -25426 13433 -25392
rect 13671 -25426 13891 -25392
rect 14129 -25426 14349 -25392
rect 14587 -25426 14807 -25392
rect 15045 -25426 15265 -25392
rect 15503 -25426 15723 -25392
rect 16381 -25426 16601 -25392
rect 16839 -25426 17059 -25392
rect 17297 -25426 17517 -25392
rect 17755 -25426 17975 -25392
rect 18213 -25426 18433 -25392
rect 18671 -25426 18891 -25392
rect 19129 -25426 19349 -25392
rect 19587 -25426 19807 -25392
rect 20045 -25426 20265 -25392
rect 20503 -25426 20723 -25392
rect 26940 -21433 27160 -21399
rect 27398 -21433 27618 -21399
rect 27856 -21433 28076 -21399
rect 28314 -21433 28534 -21399
rect 28772 -21433 28992 -21399
rect 29230 -21433 29450 -21399
rect 29688 -21433 29908 -21399
rect 30146 -21433 30366 -21399
rect 30604 -21433 30824 -21399
rect 31062 -21433 31282 -21399
rect 31520 -21433 31740 -21399
rect 31978 -21433 32198 -21399
rect 32436 -21433 32656 -21399
rect 32894 -21433 33114 -21399
rect 33352 -21433 33572 -21399
rect 33810 -21433 34030 -21399
rect 34268 -21433 34488 -21399
rect 34726 -21433 34946 -21399
rect 26940 -23161 27160 -23127
rect 27398 -23161 27618 -23127
rect 27856 -23161 28076 -23127
rect 28314 -23161 28534 -23127
rect 28772 -23161 28992 -23127
rect 29230 -23161 29450 -23127
rect 29688 -23161 29908 -23127
rect 30146 -23161 30366 -23127
rect 30604 -23161 30824 -23127
rect 31062 -23161 31282 -23127
rect 31520 -23161 31740 -23127
rect 31978 -23161 32198 -23127
rect 32436 -23161 32656 -23127
rect 32894 -23161 33114 -23127
rect 33352 -23161 33572 -23127
rect 33810 -23161 34030 -23127
rect 34268 -23161 34488 -23127
rect 34726 -23161 34946 -23127
rect 26381 -24098 26601 -24064
rect 26839 -24098 27059 -24064
rect 27297 -24098 27517 -24064
rect 27755 -24098 27975 -24064
rect 28213 -24098 28433 -24064
rect 28671 -24098 28891 -24064
rect 29129 -24098 29349 -24064
rect 29587 -24098 29807 -24064
rect 30045 -24098 30265 -24064
rect 30503 -24098 30723 -24064
rect 31381 -24098 31601 -24064
rect 31839 -24098 32059 -24064
rect 32297 -24098 32517 -24064
rect 32755 -24098 32975 -24064
rect 33213 -24098 33433 -24064
rect 33671 -24098 33891 -24064
rect 34129 -24098 34349 -24064
rect 34587 -24098 34807 -24064
rect 35045 -24098 35265 -24064
rect 35503 -24098 35723 -24064
rect 26381 -25426 26601 -25392
rect 26839 -25426 27059 -25392
rect 27297 -25426 27517 -25392
rect 27755 -25426 27975 -25392
rect 28213 -25426 28433 -25392
rect 28671 -25426 28891 -25392
rect 29129 -25426 29349 -25392
rect 29587 -25426 29807 -25392
rect 30045 -25426 30265 -25392
rect 30503 -25426 30723 -25392
rect 31381 -25426 31601 -25392
rect 31839 -25426 32059 -25392
rect 32297 -25426 32517 -25392
rect 32755 -25426 32975 -25392
rect 33213 -25426 33433 -25392
rect 33671 -25426 33891 -25392
rect 34129 -25426 34349 -25392
rect 34587 -25426 34807 -25392
rect 35045 -25426 35265 -25392
rect 35503 -25426 35723 -25392
rect 11380 -26600 11600 -26566
rect 11838 -26600 12058 -26566
rect 12296 -26600 12516 -26566
rect 12754 -26600 12974 -26566
rect 13212 -26600 13432 -26566
rect 13670 -26600 13890 -26566
rect 14128 -26600 14348 -26566
rect 14586 -26600 14806 -26566
rect 15044 -26600 15264 -26566
rect 15502 -26600 15722 -26566
rect 16380 -26600 16600 -26566
rect 16838 -26600 17058 -26566
rect 17296 -26600 17516 -26566
rect 17754 -26600 17974 -26566
rect 18212 -26600 18432 -26566
rect 18670 -26600 18890 -26566
rect 19128 -26600 19348 -26566
rect 19586 -26600 19806 -26566
rect 20044 -26600 20264 -26566
rect 20502 -26600 20722 -26566
rect 11380 -26910 11600 -26876
rect 11838 -26910 12058 -26876
rect 12296 -26910 12516 -26876
rect 12754 -26910 12974 -26876
rect 13212 -26910 13432 -26876
rect 13670 -26910 13890 -26876
rect 14128 -26910 14348 -26876
rect 14586 -26910 14806 -26876
rect 15044 -26910 15264 -26876
rect 15502 -26910 15722 -26876
rect 16380 -26910 16600 -26876
rect 16838 -26910 17058 -26876
rect 17296 -26910 17516 -26876
rect 17754 -26910 17974 -26876
rect 18212 -26910 18432 -26876
rect 18670 -26910 18890 -26876
rect 19128 -26910 19348 -26876
rect 19586 -26910 19806 -26876
rect 20044 -26910 20264 -26876
rect 20502 -26910 20722 -26876
rect 11380 -27268 11600 -27234
rect 11838 -27268 12058 -27234
rect 12296 -27268 12516 -27234
rect 12754 -27268 12974 -27234
rect 13212 -27268 13432 -27234
rect 13670 -27268 13890 -27234
rect 14128 -27268 14348 -27234
rect 14586 -27268 14806 -27234
rect 15044 -27268 15264 -27234
rect 15502 -27268 15722 -27234
rect 11380 -27578 11600 -27544
rect 11838 -27578 12058 -27544
rect 12296 -27578 12516 -27544
rect 12754 -27578 12974 -27544
rect 13212 -27578 13432 -27544
rect 13670 -27578 13890 -27544
rect 14128 -27578 14348 -27544
rect 14586 -27578 14806 -27544
rect 15044 -27578 15264 -27544
rect 15502 -27578 15722 -27544
rect 26380 -26600 26600 -26566
rect 26838 -26600 27058 -26566
rect 27296 -26600 27516 -26566
rect 27754 -26600 27974 -26566
rect 28212 -26600 28432 -26566
rect 28670 -26600 28890 -26566
rect 29128 -26600 29348 -26566
rect 29586 -26600 29806 -26566
rect 30044 -26600 30264 -26566
rect 30502 -26600 30722 -26566
rect 31380 -26600 31600 -26566
rect 31838 -26600 32058 -26566
rect 32296 -26600 32516 -26566
rect 32754 -26600 32974 -26566
rect 33212 -26600 33432 -26566
rect 33670 -26600 33890 -26566
rect 34128 -26600 34348 -26566
rect 34586 -26600 34806 -26566
rect 35044 -26600 35264 -26566
rect 35502 -26600 35722 -26566
rect 26380 -26910 26600 -26876
rect 26838 -26910 27058 -26876
rect 27296 -26910 27516 -26876
rect 27754 -26910 27974 -26876
rect 28212 -26910 28432 -26876
rect 28670 -26910 28890 -26876
rect 29128 -26910 29348 -26876
rect 29586 -26910 29806 -26876
rect 30044 -26910 30264 -26876
rect 30502 -26910 30722 -26876
rect 31380 -26910 31600 -26876
rect 31838 -26910 32058 -26876
rect 32296 -26910 32516 -26876
rect 32754 -26910 32974 -26876
rect 33212 -26910 33432 -26876
rect 33670 -26910 33890 -26876
rect 34128 -26910 34348 -26876
rect 34586 -26910 34806 -26876
rect 35044 -26910 35264 -26876
rect 35502 -26910 35722 -26876
rect 26380 -27268 26600 -27234
rect 26838 -27268 27058 -27234
rect 27296 -27268 27516 -27234
rect 27754 -27268 27974 -27234
rect 28212 -27268 28432 -27234
rect 28670 -27268 28890 -27234
rect 29128 -27268 29348 -27234
rect 29586 -27268 29806 -27234
rect 30044 -27268 30264 -27234
rect 30502 -27268 30722 -27234
rect 26380 -27578 26600 -27544
rect 26838 -27578 27058 -27544
rect 27296 -27578 27516 -27544
rect 27754 -27578 27974 -27544
rect 28212 -27578 28432 -27544
rect 28670 -27578 28890 -27544
rect 29128 -27578 29348 -27544
rect 29586 -27578 29806 -27544
rect 30044 -27578 30264 -27544
rect 30502 -27578 30722 -27544
<< locali >>
rect 15426 4148 15526 4310
rect 24350 4148 24450 4310
rect 17754 3282 17770 3316
rect 17990 3282 18006 3316
rect 18212 3282 18228 3316
rect 18448 3282 18464 3316
rect 18670 3282 18686 3316
rect 18906 3282 18922 3316
rect 19128 3282 19144 3316
rect 19364 3282 19380 3316
rect 19586 3282 19602 3316
rect 19822 3282 19838 3316
rect 20044 3282 20060 3316
rect 20280 3282 20296 3316
rect 20502 3282 20518 3316
rect 20738 3282 20754 3316
rect 20960 3282 20976 3316
rect 21196 3282 21212 3316
rect 21418 3282 21434 3316
rect 21654 3282 21670 3316
rect 21876 3282 21892 3316
rect 22112 3282 22128 3316
rect 17634 3232 17668 3248
rect 17634 3040 17668 3056
rect 18092 3232 18126 3248
rect 18092 3040 18126 3056
rect 18550 3232 18584 3248
rect 18550 3040 18584 3056
rect 19008 3232 19042 3248
rect 19008 3040 19042 3056
rect 19466 3232 19500 3248
rect 19466 3040 19500 3056
rect 19924 3232 19958 3248
rect 19924 3040 19958 3056
rect 20382 3232 20416 3248
rect 20382 3040 20416 3056
rect 20840 3232 20874 3248
rect 20840 3040 20874 3056
rect 21298 3232 21332 3248
rect 21298 3040 21332 3056
rect 21756 3232 21790 3248
rect 21756 3040 21790 3056
rect 22214 3232 22248 3248
rect 22214 3040 22248 3056
rect 17754 2972 17770 3006
rect 17990 2972 18006 3006
rect 18212 2972 18228 3006
rect 18448 2972 18464 3006
rect 18670 2972 18686 3006
rect 18906 2972 18922 3006
rect 19128 2972 19144 3006
rect 19364 2972 19380 3006
rect 19586 2972 19602 3006
rect 19822 2972 19838 3006
rect 20044 2972 20060 3006
rect 20280 2972 20296 3006
rect 20502 2972 20518 3006
rect 20738 2972 20754 3006
rect 20960 2972 20976 3006
rect 21196 2972 21212 3006
rect 21418 2972 21434 3006
rect 21654 2972 21670 3006
rect 21876 2972 21892 3006
rect 22112 2972 22128 3006
rect 15426 2510 15526 2672
rect 24350 2510 24450 2672
rect 26008 4148 26108 4310
rect 31352 4148 31452 4310
rect 26516 3282 26532 3316
rect 26752 3282 26768 3316
rect 26974 3282 26990 3316
rect 27210 3282 27226 3316
rect 27432 3282 27448 3316
rect 27668 3282 27684 3316
rect 27890 3282 27906 3316
rect 28126 3282 28142 3316
rect 28348 3282 28364 3316
rect 28584 3282 28600 3316
rect 28806 3282 28822 3316
rect 29042 3282 29058 3316
rect 29264 3282 29280 3316
rect 29500 3282 29516 3316
rect 29722 3282 29738 3316
rect 29958 3282 29974 3316
rect 30180 3282 30196 3316
rect 30416 3282 30432 3316
rect 30638 3282 30654 3316
rect 30874 3282 30890 3316
rect 26396 3232 26430 3248
rect 26396 3040 26430 3056
rect 26854 3232 26888 3248
rect 26854 3040 26888 3056
rect 27312 3232 27346 3248
rect 27312 3040 27346 3056
rect 27770 3232 27804 3248
rect 27770 3040 27804 3056
rect 28228 3232 28262 3248
rect 28228 3040 28262 3056
rect 28686 3232 28720 3248
rect 28686 3040 28720 3056
rect 29144 3232 29178 3248
rect 29144 3040 29178 3056
rect 29602 3232 29636 3248
rect 29602 3040 29636 3056
rect 30060 3232 30094 3248
rect 30060 3040 30094 3056
rect 30518 3232 30552 3248
rect 30518 3040 30552 3056
rect 30976 3232 31010 3248
rect 30976 3040 31010 3056
rect 26516 2972 26532 3006
rect 26752 2972 26768 3006
rect 26974 2972 26990 3006
rect 27210 2972 27226 3006
rect 27432 2972 27448 3006
rect 27668 2972 27684 3006
rect 27890 2972 27906 3006
rect 28126 2972 28142 3006
rect 28348 2972 28364 3006
rect 28584 2972 28600 3006
rect 28806 2972 28822 3006
rect 29042 2972 29058 3006
rect 29264 2972 29280 3006
rect 29500 2972 29516 3006
rect 29722 2972 29738 3006
rect 29958 2972 29974 3006
rect 30180 2972 30196 3006
rect 30416 2972 30432 3006
rect 30638 2972 30654 3006
rect 30874 2972 30890 3006
rect 26008 2430 26108 2592
rect 31352 2430 31452 2592
rect 31542 2473 31571 2507
rect 31605 2473 31663 2507
rect 31697 2473 31755 2507
rect 31789 2473 31847 2507
rect 31881 2473 31939 2507
rect 31973 2473 32031 2507
rect 32065 2473 32123 2507
rect 32157 2473 32215 2507
rect 32249 2473 32278 2507
rect 31606 2427 31652 2473
rect 31606 2393 31618 2427
rect 31606 2359 31652 2393
rect 31606 2325 31618 2359
rect 31606 2309 31652 2325
rect 31686 2427 31752 2439
rect 31686 2393 31702 2427
rect 31736 2393 31752 2427
rect 31686 2359 31752 2393
rect 31844 2431 31897 2473
rect 31844 2397 31863 2431
rect 31844 2381 31897 2397
rect 31931 2423 31997 2439
rect 31931 2389 31947 2423
rect 31981 2389 31997 2423
rect 31686 2325 31702 2359
rect 31736 2325 31752 2359
rect 31686 2313 31752 2325
rect 31706 2276 31752 2313
rect 31931 2345 31997 2389
rect 32031 2431 32065 2473
rect 32031 2381 32065 2397
rect 32099 2423 32165 2439
rect 32099 2389 32115 2423
rect 32149 2389 32165 2423
rect 32099 2345 32165 2389
rect 32199 2430 32249 2473
rect 32233 2396 32249 2430
rect 32199 2380 32249 2396
rect 31931 2309 32252 2345
rect 32199 2276 32252 2309
rect 31606 2274 31622 2275
rect 15426 2112 15526 2274
rect 24350 2112 24450 2274
rect 31656 2241 31672 2275
rect 31654 2227 31672 2241
rect 31706 2228 31712 2276
rect 31839 2228 31848 2275
rect 31896 2241 31947 2275
rect 31981 2241 32031 2275
rect 32065 2241 32115 2275
rect 32149 2241 32165 2275
rect 31896 2228 32165 2241
rect 15922 1440 15938 1474
rect 16158 1440 16174 1474
rect 16380 1440 16396 1474
rect 16616 1440 16632 1474
rect 16838 1440 16854 1474
rect 17074 1440 17090 1474
rect 17296 1440 17312 1474
rect 17532 1440 17548 1474
rect 17754 1440 17770 1474
rect 17990 1440 18006 1474
rect 18212 1440 18228 1474
rect 18448 1440 18464 1474
rect 18670 1440 18686 1474
rect 18906 1440 18922 1474
rect 19128 1440 19144 1474
rect 19364 1440 19380 1474
rect 19586 1440 19602 1474
rect 19822 1440 19838 1474
rect 20044 1440 20060 1474
rect 20280 1440 20296 1474
rect 20502 1440 20518 1474
rect 20738 1440 20754 1474
rect 20960 1440 20976 1474
rect 21196 1440 21212 1474
rect 21418 1440 21434 1474
rect 21654 1440 21670 1474
rect 21876 1440 21892 1474
rect 22112 1440 22128 1474
rect 22334 1440 22350 1474
rect 22570 1440 22586 1474
rect 22792 1440 22808 1474
rect 23028 1440 23044 1474
rect 23250 1440 23266 1474
rect 23486 1440 23502 1474
rect 23708 1440 23724 1474
rect 23944 1440 23960 1474
rect 15802 1381 15836 1397
rect 15802 -211 15836 -195
rect 16260 1381 16294 1397
rect 16260 -211 16294 -195
rect 16718 1381 16752 1397
rect 16718 -211 16752 -195
rect 17176 1381 17210 1397
rect 17176 -211 17210 -195
rect 17634 1381 17668 1397
rect 17634 -211 17668 -195
rect 18092 1381 18126 1397
rect 18092 -211 18126 -195
rect 18550 1381 18584 1397
rect 18550 -211 18584 -195
rect 19008 1381 19042 1397
rect 19008 -211 19042 -195
rect 19466 1381 19500 1397
rect 19466 -211 19500 -195
rect 19924 1381 19958 1397
rect 19924 -211 19958 -195
rect 20382 1381 20416 1397
rect 20382 -211 20416 -195
rect 20840 1381 20874 1397
rect 20840 -211 20874 -195
rect 21298 1381 21332 1397
rect 21298 -211 21332 -195
rect 21756 1381 21790 1397
rect 21756 -211 21790 -195
rect 22214 1381 22248 1397
rect 22214 -211 22248 -195
rect 22672 1381 22706 1397
rect 22672 -211 22706 -195
rect 23130 1381 23164 1397
rect 23130 -211 23164 -195
rect 23588 1381 23622 1397
rect 23588 -211 23622 -195
rect 24046 1381 24080 1397
rect 24046 -211 24080 -195
rect 15922 -288 15938 -254
rect 16158 -288 16174 -254
rect 16380 -288 16396 -254
rect 16616 -288 16632 -254
rect 16838 -288 16854 -254
rect 17074 -288 17090 -254
rect 17296 -288 17312 -254
rect 17532 -288 17548 -254
rect 17754 -288 17770 -254
rect 17990 -288 18006 -254
rect 18212 -288 18228 -254
rect 18448 -288 18464 -254
rect 18670 -288 18686 -254
rect 18906 -288 18922 -254
rect 19128 -288 19144 -254
rect 19364 -288 19380 -254
rect 19586 -288 19602 -254
rect 19822 -288 19838 -254
rect 20044 -288 20060 -254
rect 20280 -288 20296 -254
rect 20502 -288 20518 -254
rect 20738 -288 20754 -254
rect 20960 -288 20976 -254
rect 21196 -288 21212 -254
rect 21418 -288 21434 -254
rect 21654 -288 21670 -254
rect 21876 -288 21892 -254
rect 22112 -288 22128 -254
rect 22334 -288 22350 -254
rect 22570 -288 22586 -254
rect 22792 -288 22808 -254
rect 23028 -288 23044 -254
rect 23250 -288 23266 -254
rect 23486 -288 23502 -254
rect 23708 -288 23724 -254
rect 23944 -288 23960 -254
rect 15426 -1658 15526 -1496
rect 24350 -1658 24450 -1496
rect 26008 2032 26108 2194
rect 31352 2032 31452 2194
rect 31706 2193 31752 2228
rect 31839 2225 32165 2228
rect 32199 2228 32204 2276
rect 31610 2175 31652 2191
rect 31610 2141 31618 2175
rect 31610 2107 31652 2141
rect 31610 2073 31618 2107
rect 31610 2039 31652 2073
rect 31610 2005 31618 2039
rect 31610 1963 31652 2005
rect 31686 2175 31752 2193
rect 32199 2191 32252 2228
rect 31686 2141 31702 2175
rect 31736 2141 31752 2175
rect 31686 2107 31752 2141
rect 31686 2073 31702 2107
rect 31736 2073 31752 2107
rect 31686 2039 31752 2073
rect 31686 2005 31702 2039
rect 31736 2005 31752 2039
rect 31686 1997 31752 2005
rect 31844 2175 31897 2191
rect 31844 2141 31863 2175
rect 31844 2107 31897 2141
rect 31844 2073 31863 2107
rect 31844 2039 31897 2073
rect 31844 2005 31863 2039
rect 31844 1963 31897 2005
rect 31931 2175 32252 2191
rect 31931 2141 31947 2175
rect 31981 2157 32115 2175
rect 31981 2141 31997 2157
rect 31931 2107 31997 2141
rect 32099 2141 32115 2157
rect 32149 2153 32252 2175
rect 32149 2141 32165 2153
rect 31931 2073 31947 2107
rect 31981 2073 31997 2107
rect 31931 2039 31997 2073
rect 31931 2005 31947 2039
rect 31981 2005 31997 2039
rect 31931 1997 31997 2005
rect 32031 2107 32065 2123
rect 32031 2039 32065 2073
rect 32031 1963 32065 2005
rect 32099 2107 32165 2141
rect 32099 2073 32115 2107
rect 32149 2073 32165 2107
rect 32099 2039 32165 2073
rect 32099 2005 32115 2039
rect 32149 2005 32165 2039
rect 32099 1997 32165 2005
rect 32199 2039 32241 2055
rect 32233 2005 32241 2039
rect 32199 1963 32241 2005
rect 31542 1929 31571 1963
rect 31605 1929 31663 1963
rect 31697 1929 31755 1963
rect 31789 1929 31847 1963
rect 31881 1929 31939 1963
rect 31973 1929 32031 1963
rect 32065 1929 32123 1963
rect 32157 1929 32215 1963
rect 32249 1929 32278 1963
rect 26517 1860 26533 1894
rect 26753 1860 26769 1894
rect 26975 1860 26991 1894
rect 27211 1860 27227 1894
rect 27433 1860 27449 1894
rect 27669 1860 27685 1894
rect 27891 1860 27907 1894
rect 28127 1860 28143 1894
rect 28349 1860 28365 1894
rect 28585 1860 28601 1894
rect 28807 1860 28823 1894
rect 29043 1860 29059 1894
rect 29265 1860 29281 1894
rect 29501 1860 29517 1894
rect 29723 1860 29739 1894
rect 29959 1860 29975 1894
rect 30181 1860 30197 1894
rect 30417 1860 30433 1894
rect 30639 1860 30655 1894
rect 30875 1860 30891 1894
rect 26397 1801 26431 1817
rect 26397 609 26431 625
rect 26855 1801 26889 1817
rect 26855 609 26889 625
rect 27313 1801 27347 1817
rect 27313 609 27347 625
rect 27771 1801 27805 1817
rect 27771 609 27805 625
rect 28229 1801 28263 1817
rect 28229 609 28263 625
rect 28687 1801 28721 1817
rect 28687 609 28721 625
rect 29145 1801 29179 1817
rect 29145 609 29179 625
rect 29603 1801 29637 1817
rect 29603 609 29637 625
rect 30061 1801 30095 1817
rect 30061 609 30095 625
rect 30519 1801 30553 1817
rect 30519 609 30553 625
rect 30977 1801 31011 1817
rect 30977 609 31011 625
rect 26517 532 26533 566
rect 26753 532 26769 566
rect 26975 532 26991 566
rect 27211 532 27227 566
rect 27433 532 27449 566
rect 27669 532 27685 566
rect 27891 532 27907 566
rect 28127 532 28143 566
rect 28349 532 28365 566
rect 28585 532 28601 566
rect 28807 532 28823 566
rect 29043 532 29059 566
rect 29265 532 29281 566
rect 29501 532 29517 566
rect 29723 532 29739 566
rect 29959 532 29975 566
rect 30181 532 30197 566
rect 30417 532 30433 566
rect 30639 532 30655 566
rect 30875 532 30891 566
rect 26008 -1658 26108 -1496
rect 31352 -1658 31452 -1496
rect 10818 -2190 10918 -2028
rect 21162 -2190 21262 -2028
rect 11924 -3433 11940 -3399
rect 12160 -3433 12176 -3399
rect 12382 -3433 12398 -3399
rect 12618 -3433 12634 -3399
rect 12840 -3433 12856 -3399
rect 13076 -3433 13092 -3399
rect 13298 -3433 13314 -3399
rect 13534 -3433 13550 -3399
rect 13756 -3433 13772 -3399
rect 13992 -3433 14008 -3399
rect 14214 -3433 14230 -3399
rect 14450 -3433 14466 -3399
rect 14672 -3433 14688 -3399
rect 14908 -3433 14924 -3399
rect 15130 -3433 15146 -3399
rect 15366 -3433 15382 -3399
rect 15588 -3433 15604 -3399
rect 15824 -3433 15840 -3399
rect 16046 -3433 16062 -3399
rect 16282 -3433 16298 -3399
rect 16504 -3433 16520 -3399
rect 16740 -3433 16756 -3399
rect 16962 -3433 16978 -3399
rect 17198 -3433 17214 -3399
rect 17420 -3433 17436 -3399
rect 17656 -3433 17672 -3399
rect 17878 -3433 17894 -3399
rect 18114 -3433 18130 -3399
rect 18336 -3433 18352 -3399
rect 18572 -3433 18588 -3399
rect 18794 -3433 18810 -3399
rect 19030 -3433 19046 -3399
rect 19252 -3433 19268 -3399
rect 19488 -3433 19504 -3399
rect 19710 -3433 19726 -3399
rect 19946 -3433 19962 -3399
rect 11804 -3492 11838 -3476
rect 11804 -5084 11838 -5068
rect 12262 -3492 12296 -3476
rect 12262 -5084 12296 -5068
rect 12720 -3492 12754 -3476
rect 12720 -5084 12754 -5068
rect 13178 -3492 13212 -3476
rect 13178 -5084 13212 -5068
rect 13636 -3492 13670 -3476
rect 13636 -5084 13670 -5068
rect 14094 -3492 14128 -3476
rect 14094 -5084 14128 -5068
rect 14552 -3492 14586 -3476
rect 14552 -5084 14586 -5068
rect 15010 -3492 15044 -3476
rect 15010 -5084 15044 -5068
rect 15468 -3492 15502 -3476
rect 15468 -5084 15502 -5068
rect 15926 -3492 15960 -3476
rect 15926 -5084 15960 -5068
rect 16384 -3492 16418 -3476
rect 16384 -5084 16418 -5068
rect 16842 -3492 16876 -3476
rect 16842 -5084 16876 -5068
rect 17300 -3492 17334 -3476
rect 17300 -5084 17334 -5068
rect 17758 -3492 17792 -3476
rect 17758 -5084 17792 -5068
rect 18216 -3492 18250 -3476
rect 18216 -5084 18250 -5068
rect 18674 -3492 18708 -3476
rect 18674 -5084 18708 -5068
rect 19132 -3492 19166 -3476
rect 19132 -5084 19166 -5068
rect 19590 -3492 19624 -3476
rect 19590 -5084 19624 -5068
rect 20048 -3492 20082 -3476
rect 20048 -5084 20082 -5068
rect 11924 -5161 11940 -5127
rect 12160 -5161 12176 -5127
rect 12382 -5161 12398 -5127
rect 12618 -5161 12634 -5127
rect 12840 -5161 12856 -5127
rect 13076 -5161 13092 -5127
rect 13298 -5161 13314 -5127
rect 13534 -5161 13550 -5127
rect 13756 -5161 13772 -5127
rect 13992 -5161 14008 -5127
rect 14214 -5161 14230 -5127
rect 14450 -5161 14466 -5127
rect 14672 -5161 14688 -5127
rect 14908 -5161 14924 -5127
rect 15130 -5161 15146 -5127
rect 15366 -5161 15382 -5127
rect 15588 -5161 15604 -5127
rect 15824 -5161 15840 -5127
rect 16046 -5161 16062 -5127
rect 16282 -5161 16298 -5127
rect 16504 -5161 16520 -5127
rect 16740 -5161 16756 -5127
rect 16962 -5161 16978 -5127
rect 17198 -5161 17214 -5127
rect 17420 -5161 17436 -5127
rect 17656 -5161 17672 -5127
rect 17878 -5161 17894 -5127
rect 18114 -5161 18130 -5127
rect 18336 -5161 18352 -5127
rect 18572 -5161 18588 -5127
rect 18794 -5161 18810 -5127
rect 19030 -5161 19046 -5127
rect 19252 -5161 19268 -5127
rect 19488 -5161 19504 -5127
rect 19710 -5161 19726 -5127
rect 19946 -5161 19962 -5127
rect 15682 -5244 16142 -5238
rect 15682 -5292 15688 -5244
rect 15736 -5292 16142 -5244
rect 15682 -5298 16142 -5292
rect 11365 -6098 11381 -6064
rect 11601 -6098 11617 -6064
rect 11823 -6098 11839 -6064
rect 12059 -6098 12075 -6064
rect 12281 -6098 12297 -6064
rect 12517 -6098 12533 -6064
rect 12739 -6098 12755 -6064
rect 12975 -6098 12991 -6064
rect 13197 -6098 13213 -6064
rect 13433 -6098 13449 -6064
rect 13655 -6098 13671 -6064
rect 13891 -6098 13907 -6064
rect 14113 -6098 14129 -6064
rect 14349 -6098 14365 -6064
rect 14571 -6098 14587 -6064
rect 14807 -6098 14823 -6064
rect 15029 -6098 15045 -6064
rect 15265 -6098 15281 -6064
rect 15487 -6098 15503 -6064
rect 15723 -6098 15739 -6064
rect 16365 -6098 16381 -6064
rect 16601 -6098 16617 -6064
rect 16823 -6098 16839 -6064
rect 17059 -6098 17075 -6064
rect 17281 -6098 17297 -6064
rect 17517 -6098 17533 -6064
rect 17739 -6098 17755 -6064
rect 17975 -6098 17991 -6064
rect 18197 -6098 18213 -6064
rect 18433 -6098 18449 -6064
rect 18655 -6098 18671 -6064
rect 18891 -6098 18907 -6064
rect 19113 -6098 19129 -6064
rect 19349 -6098 19365 -6064
rect 19571 -6098 19587 -6064
rect 19807 -6098 19823 -6064
rect 20029 -6098 20045 -6064
rect 20265 -6098 20281 -6064
rect 20487 -6098 20503 -6064
rect 20723 -6098 20739 -6064
rect 11245 -6157 11279 -6141
rect 11245 -7349 11279 -7333
rect 11703 -6157 11737 -6141
rect 11703 -7349 11737 -7333
rect 12161 -6157 12195 -6141
rect 12161 -7349 12195 -7333
rect 12619 -6157 12653 -6141
rect 12619 -7349 12653 -7333
rect 13077 -6157 13111 -6141
rect 13077 -7349 13111 -7333
rect 13535 -6157 13569 -6141
rect 13535 -7349 13569 -7333
rect 13993 -6157 14027 -6141
rect 13993 -7349 14027 -7333
rect 14451 -6157 14485 -6141
rect 14451 -7349 14485 -7333
rect 14909 -6157 14943 -6141
rect 14909 -7349 14943 -7333
rect 15367 -6157 15401 -6141
rect 15367 -7349 15401 -7333
rect 15825 -6157 15859 -6141
rect 15825 -7349 15859 -7333
rect 16245 -6157 16279 -6141
rect 16245 -7349 16279 -7333
rect 16703 -6157 16737 -6141
rect 16703 -7349 16737 -7333
rect 17161 -6157 17195 -6141
rect 17161 -7349 17195 -7333
rect 17619 -6157 17653 -6141
rect 17619 -7349 17653 -7333
rect 18077 -6157 18111 -6141
rect 18077 -7349 18111 -7333
rect 18535 -6157 18569 -6141
rect 18535 -7349 18569 -7333
rect 18993 -6157 19027 -6141
rect 18993 -7349 19027 -7333
rect 19451 -6157 19485 -6141
rect 19451 -7349 19485 -7333
rect 19909 -6157 19943 -6141
rect 19909 -7349 19943 -7333
rect 20367 -6157 20401 -6141
rect 20367 -7349 20401 -7333
rect 20825 -6157 20859 -6141
rect 20825 -7349 20859 -7333
rect 11365 -7426 11381 -7392
rect 11601 -7426 11617 -7392
rect 11823 -7426 11839 -7392
rect 12059 -7426 12075 -7392
rect 12281 -7426 12297 -7392
rect 12517 -7426 12533 -7392
rect 12739 -7426 12755 -7392
rect 12975 -7426 12991 -7392
rect 13197 -7426 13213 -7392
rect 13433 -7426 13449 -7392
rect 13655 -7426 13671 -7392
rect 13891 -7426 13907 -7392
rect 14113 -7426 14129 -7392
rect 14349 -7426 14365 -7392
rect 14571 -7426 14587 -7392
rect 14807 -7426 14823 -7392
rect 15029 -7426 15045 -7392
rect 15265 -7426 15281 -7392
rect 15487 -7426 15503 -7392
rect 15723 -7426 15739 -7392
rect 16365 -7426 16381 -7392
rect 16601 -7426 16617 -7392
rect 16823 -7426 16839 -7392
rect 17059 -7426 17075 -7392
rect 17281 -7426 17297 -7392
rect 17517 -7426 17533 -7392
rect 17739 -7426 17755 -7392
rect 17975 -7426 17991 -7392
rect 18197 -7426 18213 -7392
rect 18433 -7426 18449 -7392
rect 18655 -7426 18671 -7392
rect 18891 -7426 18907 -7392
rect 19113 -7426 19129 -7392
rect 19349 -7426 19365 -7392
rect 19571 -7426 19587 -7392
rect 19807 -7426 19823 -7392
rect 20029 -7426 20045 -7392
rect 20265 -7426 20281 -7392
rect 20487 -7426 20503 -7392
rect 20723 -7426 20739 -7392
rect 10818 -7872 10918 -7710
rect 21162 -7872 21262 -7710
rect 25818 -2190 25918 -2028
rect 36162 -2190 36262 -2028
rect 26924 -3433 26940 -3399
rect 27160 -3433 27176 -3399
rect 27382 -3433 27398 -3399
rect 27618 -3433 27634 -3399
rect 27840 -3433 27856 -3399
rect 28076 -3433 28092 -3399
rect 28298 -3433 28314 -3399
rect 28534 -3433 28550 -3399
rect 28756 -3433 28772 -3399
rect 28992 -3433 29008 -3399
rect 29214 -3433 29230 -3399
rect 29450 -3433 29466 -3399
rect 29672 -3433 29688 -3399
rect 29908 -3433 29924 -3399
rect 30130 -3433 30146 -3399
rect 30366 -3433 30382 -3399
rect 30588 -3433 30604 -3399
rect 30824 -3433 30840 -3399
rect 31046 -3433 31062 -3399
rect 31282 -3433 31298 -3399
rect 31504 -3433 31520 -3399
rect 31740 -3433 31756 -3399
rect 31962 -3433 31978 -3399
rect 32198 -3433 32214 -3399
rect 32420 -3433 32436 -3399
rect 32656 -3433 32672 -3399
rect 32878 -3433 32894 -3399
rect 33114 -3433 33130 -3399
rect 33336 -3433 33352 -3399
rect 33572 -3433 33588 -3399
rect 33794 -3433 33810 -3399
rect 34030 -3433 34046 -3399
rect 34252 -3433 34268 -3399
rect 34488 -3433 34504 -3399
rect 34710 -3433 34726 -3399
rect 34946 -3433 34962 -3399
rect 26804 -3492 26838 -3476
rect 26804 -5084 26838 -5068
rect 27262 -3492 27296 -3476
rect 27262 -5084 27296 -5068
rect 27720 -3492 27754 -3476
rect 27720 -5084 27754 -5068
rect 28178 -3492 28212 -3476
rect 28178 -5084 28212 -5068
rect 28636 -3492 28670 -3476
rect 28636 -5084 28670 -5068
rect 29094 -3492 29128 -3476
rect 29094 -5084 29128 -5068
rect 29552 -3492 29586 -3476
rect 29552 -5084 29586 -5068
rect 30010 -3492 30044 -3476
rect 30010 -5084 30044 -5068
rect 30468 -3492 30502 -3476
rect 30468 -5084 30502 -5068
rect 30926 -3492 30960 -3476
rect 30926 -5084 30960 -5068
rect 31384 -3492 31418 -3476
rect 31384 -5084 31418 -5068
rect 31842 -3492 31876 -3476
rect 31842 -5084 31876 -5068
rect 32300 -3492 32334 -3476
rect 32300 -5084 32334 -5068
rect 32758 -3492 32792 -3476
rect 32758 -5084 32792 -5068
rect 33216 -3492 33250 -3476
rect 33216 -5084 33250 -5068
rect 33674 -3492 33708 -3476
rect 33674 -5084 33708 -5068
rect 34132 -3492 34166 -3476
rect 34132 -5084 34166 -5068
rect 34590 -3492 34624 -3476
rect 34590 -5084 34624 -5068
rect 35048 -3492 35082 -3476
rect 35048 -5084 35082 -5068
rect 26924 -5161 26940 -5127
rect 27160 -5161 27176 -5127
rect 27382 -5161 27398 -5127
rect 27618 -5161 27634 -5127
rect 27840 -5161 27856 -5127
rect 28076 -5161 28092 -5127
rect 28298 -5161 28314 -5127
rect 28534 -5161 28550 -5127
rect 28756 -5161 28772 -5127
rect 28992 -5161 29008 -5127
rect 29214 -5161 29230 -5127
rect 29450 -5161 29466 -5127
rect 29672 -5161 29688 -5127
rect 29908 -5161 29924 -5127
rect 30130 -5161 30146 -5127
rect 30366 -5161 30382 -5127
rect 30588 -5161 30604 -5127
rect 30824 -5161 30840 -5127
rect 31046 -5161 31062 -5127
rect 31282 -5161 31298 -5127
rect 31504 -5161 31520 -5127
rect 31740 -5161 31756 -5127
rect 31962 -5161 31978 -5127
rect 32198 -5161 32214 -5127
rect 32420 -5161 32436 -5127
rect 32656 -5161 32672 -5127
rect 32878 -5161 32894 -5127
rect 33114 -5161 33130 -5127
rect 33336 -5161 33352 -5127
rect 33572 -5161 33588 -5127
rect 33794 -5161 33810 -5127
rect 34030 -5161 34046 -5127
rect 34252 -5161 34268 -5127
rect 34488 -5161 34504 -5127
rect 34710 -5161 34726 -5127
rect 34946 -5161 34962 -5127
rect 30682 -5244 31142 -5238
rect 30682 -5292 30688 -5244
rect 30736 -5292 31142 -5244
rect 30682 -5298 31142 -5292
rect 26365 -6098 26381 -6064
rect 26601 -6098 26617 -6064
rect 26823 -6098 26839 -6064
rect 27059 -6098 27075 -6064
rect 27281 -6098 27297 -6064
rect 27517 -6098 27533 -6064
rect 27739 -6098 27755 -6064
rect 27975 -6098 27991 -6064
rect 28197 -6098 28213 -6064
rect 28433 -6098 28449 -6064
rect 28655 -6098 28671 -6064
rect 28891 -6098 28907 -6064
rect 29113 -6098 29129 -6064
rect 29349 -6098 29365 -6064
rect 29571 -6098 29587 -6064
rect 29807 -6098 29823 -6064
rect 30029 -6098 30045 -6064
rect 30265 -6098 30281 -6064
rect 30487 -6098 30503 -6064
rect 30723 -6098 30739 -6064
rect 31365 -6098 31381 -6064
rect 31601 -6098 31617 -6064
rect 31823 -6098 31839 -6064
rect 32059 -6098 32075 -6064
rect 32281 -6098 32297 -6064
rect 32517 -6098 32533 -6064
rect 32739 -6098 32755 -6064
rect 32975 -6098 32991 -6064
rect 33197 -6098 33213 -6064
rect 33433 -6098 33449 -6064
rect 33655 -6098 33671 -6064
rect 33891 -6098 33907 -6064
rect 34113 -6098 34129 -6064
rect 34349 -6098 34365 -6064
rect 34571 -6098 34587 -6064
rect 34807 -6098 34823 -6064
rect 35029 -6098 35045 -6064
rect 35265 -6098 35281 -6064
rect 35487 -6098 35503 -6064
rect 35723 -6098 35739 -6064
rect 26245 -6157 26279 -6141
rect 26245 -7349 26279 -7333
rect 26703 -6157 26737 -6141
rect 26703 -7349 26737 -7333
rect 27161 -6157 27195 -6141
rect 27161 -7349 27195 -7333
rect 27619 -6157 27653 -6141
rect 27619 -7349 27653 -7333
rect 28077 -6157 28111 -6141
rect 28077 -7349 28111 -7333
rect 28535 -6157 28569 -6141
rect 28535 -7349 28569 -7333
rect 28993 -6157 29027 -6141
rect 28993 -7349 29027 -7333
rect 29451 -6157 29485 -6141
rect 29451 -7349 29485 -7333
rect 29909 -6157 29943 -6141
rect 29909 -7349 29943 -7333
rect 30367 -6157 30401 -6141
rect 30367 -7349 30401 -7333
rect 30825 -6157 30859 -6141
rect 30825 -7349 30859 -7333
rect 31245 -6157 31279 -6141
rect 31245 -7349 31279 -7333
rect 31703 -6157 31737 -6141
rect 31703 -7349 31737 -7333
rect 32161 -6157 32195 -6141
rect 32161 -7349 32195 -7333
rect 32619 -6157 32653 -6141
rect 32619 -7349 32653 -7333
rect 33077 -6157 33111 -6141
rect 33077 -7349 33111 -7333
rect 33535 -6157 33569 -6141
rect 33535 -7349 33569 -7333
rect 33993 -6157 34027 -6141
rect 33993 -7349 34027 -7333
rect 34451 -6157 34485 -6141
rect 34451 -7349 34485 -7333
rect 34909 -6157 34943 -6141
rect 34909 -7349 34943 -7333
rect 35367 -6157 35401 -6141
rect 35367 -7349 35401 -7333
rect 35825 -6157 35859 -6141
rect 35825 -7349 35859 -7333
rect 26365 -7426 26381 -7392
rect 26601 -7426 26617 -7392
rect 26823 -7426 26839 -7392
rect 27059 -7426 27075 -7392
rect 27281 -7426 27297 -7392
rect 27517 -7426 27533 -7392
rect 27739 -7426 27755 -7392
rect 27975 -7426 27991 -7392
rect 28197 -7426 28213 -7392
rect 28433 -7426 28449 -7392
rect 28655 -7426 28671 -7392
rect 28891 -7426 28907 -7392
rect 29113 -7426 29129 -7392
rect 29349 -7426 29365 -7392
rect 29571 -7426 29587 -7392
rect 29807 -7426 29823 -7392
rect 30029 -7426 30045 -7392
rect 30265 -7426 30281 -7392
rect 30487 -7426 30503 -7392
rect 30723 -7426 30739 -7392
rect 31365 -7426 31381 -7392
rect 31601 -7426 31617 -7392
rect 31823 -7426 31839 -7392
rect 32059 -7426 32075 -7392
rect 32281 -7426 32297 -7392
rect 32517 -7426 32533 -7392
rect 32739 -7426 32755 -7392
rect 32975 -7426 32991 -7392
rect 33197 -7426 33213 -7392
rect 33433 -7426 33449 -7392
rect 33655 -7426 33671 -7392
rect 33891 -7426 33907 -7392
rect 34113 -7426 34129 -7392
rect 34349 -7426 34365 -7392
rect 34571 -7426 34587 -7392
rect 34807 -7426 34823 -7392
rect 35029 -7426 35045 -7392
rect 35265 -7426 35281 -7392
rect 35487 -7426 35503 -7392
rect 35723 -7426 35739 -7392
rect 25818 -7872 25918 -7710
rect 36162 -7872 36262 -7710
rect 10818 -8270 10918 -8108
rect 21162 -8270 21262 -8108
rect 11364 -8600 11380 -8566
rect 11600 -8600 11616 -8566
rect 11822 -8600 11838 -8566
rect 12058 -8600 12074 -8566
rect 12280 -8600 12296 -8566
rect 12516 -8600 12532 -8566
rect 12738 -8600 12754 -8566
rect 12974 -8600 12990 -8566
rect 13196 -8600 13212 -8566
rect 13432 -8600 13448 -8566
rect 13654 -8600 13670 -8566
rect 13890 -8600 13906 -8566
rect 14112 -8600 14128 -8566
rect 14348 -8600 14364 -8566
rect 14570 -8600 14586 -8566
rect 14806 -8600 14822 -8566
rect 15028 -8600 15044 -8566
rect 15264 -8600 15280 -8566
rect 15486 -8600 15502 -8566
rect 15722 -8600 15738 -8566
rect 16364 -8600 16380 -8566
rect 16600 -8600 16616 -8566
rect 16822 -8600 16838 -8566
rect 17058 -8600 17074 -8566
rect 17280 -8600 17296 -8566
rect 17516 -8600 17532 -8566
rect 17738 -8600 17754 -8566
rect 17974 -8600 17990 -8566
rect 18196 -8600 18212 -8566
rect 18432 -8600 18448 -8566
rect 18654 -8600 18670 -8566
rect 18890 -8600 18906 -8566
rect 19112 -8600 19128 -8566
rect 19348 -8600 19364 -8566
rect 19570 -8600 19586 -8566
rect 19806 -8600 19822 -8566
rect 20028 -8600 20044 -8566
rect 20264 -8600 20280 -8566
rect 20486 -8600 20502 -8566
rect 20722 -8600 20738 -8566
rect 11244 -8650 11278 -8634
rect 11244 -8842 11278 -8826
rect 11702 -8650 11736 -8634
rect 11702 -8842 11736 -8826
rect 12160 -8650 12194 -8634
rect 12160 -8842 12194 -8826
rect 12618 -8650 12652 -8634
rect 12618 -8842 12652 -8826
rect 13076 -8650 13110 -8634
rect 13076 -8842 13110 -8826
rect 13534 -8650 13568 -8634
rect 13534 -8842 13568 -8826
rect 13992 -8650 14026 -8634
rect 13992 -8842 14026 -8826
rect 14450 -8650 14484 -8634
rect 14450 -8842 14484 -8826
rect 14908 -8650 14942 -8634
rect 14908 -8842 14942 -8826
rect 15366 -8650 15400 -8634
rect 15366 -8842 15400 -8826
rect 15824 -8650 15858 -8634
rect 15824 -8842 15858 -8826
rect 16244 -8650 16278 -8634
rect 16244 -8842 16278 -8826
rect 16702 -8650 16736 -8634
rect 16702 -8842 16736 -8826
rect 17160 -8650 17194 -8634
rect 17160 -8842 17194 -8826
rect 17618 -8650 17652 -8634
rect 17618 -8842 17652 -8826
rect 18076 -8650 18110 -8634
rect 18076 -8842 18110 -8826
rect 18534 -8650 18568 -8634
rect 18534 -8842 18568 -8826
rect 18992 -8650 19026 -8634
rect 18992 -8842 19026 -8826
rect 19450 -8650 19484 -8634
rect 19450 -8842 19484 -8826
rect 19908 -8650 19942 -8634
rect 19908 -8842 19942 -8826
rect 20366 -8650 20400 -8634
rect 20366 -8842 20400 -8826
rect 20824 -8650 20858 -8634
rect 20824 -8842 20858 -8826
rect 11364 -8910 11380 -8876
rect 11600 -8910 11616 -8876
rect 11822 -8910 11838 -8876
rect 12058 -8910 12074 -8876
rect 12280 -8910 12296 -8876
rect 12516 -8910 12532 -8876
rect 12738 -8910 12754 -8876
rect 12974 -8910 12990 -8876
rect 13196 -8910 13212 -8876
rect 13432 -8910 13448 -8876
rect 13654 -8910 13670 -8876
rect 13890 -8910 13906 -8876
rect 14112 -8910 14128 -8876
rect 14348 -8910 14364 -8876
rect 14570 -8910 14586 -8876
rect 14806 -8910 14822 -8876
rect 15028 -8910 15044 -8876
rect 15264 -8910 15280 -8876
rect 15486 -8910 15502 -8876
rect 15722 -8910 15738 -8876
rect 16364 -8910 16380 -8876
rect 16600 -8910 16616 -8876
rect 16822 -8910 16838 -8876
rect 17058 -8910 17074 -8876
rect 17280 -8910 17296 -8876
rect 17516 -8910 17532 -8876
rect 17738 -8910 17754 -8876
rect 17974 -8910 17990 -8876
rect 18196 -8910 18212 -8876
rect 18432 -8910 18448 -8876
rect 18654 -8910 18670 -8876
rect 18890 -8910 18906 -8876
rect 19112 -8910 19128 -8876
rect 19348 -8910 19364 -8876
rect 19570 -8910 19586 -8876
rect 19806 -8910 19822 -8876
rect 20028 -8910 20044 -8876
rect 20264 -8910 20280 -8876
rect 20486 -8910 20502 -8876
rect 20722 -8910 20738 -8876
rect 11364 -9268 11380 -9234
rect 11600 -9268 11616 -9234
rect 11822 -9268 11838 -9234
rect 12058 -9268 12074 -9234
rect 12280 -9268 12296 -9234
rect 12516 -9268 12532 -9234
rect 12738 -9268 12754 -9234
rect 12974 -9268 12990 -9234
rect 13196 -9268 13212 -9234
rect 13432 -9268 13448 -9234
rect 13654 -9268 13670 -9234
rect 13890 -9268 13906 -9234
rect 14112 -9268 14128 -9234
rect 14348 -9268 14364 -9234
rect 14570 -9268 14586 -9234
rect 14806 -9268 14822 -9234
rect 15028 -9268 15044 -9234
rect 15264 -9268 15280 -9234
rect 15486 -9268 15502 -9234
rect 15722 -9268 15738 -9234
rect 11244 -9318 11278 -9302
rect 11244 -9510 11278 -9494
rect 11702 -9318 11736 -9302
rect 11702 -9510 11736 -9494
rect 12160 -9318 12194 -9302
rect 12160 -9510 12194 -9494
rect 12618 -9318 12652 -9302
rect 12618 -9510 12652 -9494
rect 13076 -9318 13110 -9302
rect 13076 -9510 13110 -9494
rect 13534 -9318 13568 -9302
rect 13534 -9510 13568 -9494
rect 13992 -9318 14026 -9302
rect 13992 -9510 14026 -9494
rect 14450 -9318 14484 -9302
rect 14450 -9510 14484 -9494
rect 14908 -9318 14942 -9302
rect 14908 -9510 14942 -9494
rect 15366 -9318 15400 -9302
rect 15366 -9510 15400 -9494
rect 15824 -9318 15858 -9302
rect 15824 -9510 15858 -9494
rect 11364 -9578 11380 -9544
rect 11600 -9578 11616 -9544
rect 11822 -9578 11838 -9544
rect 12058 -9578 12074 -9544
rect 12280 -9578 12296 -9544
rect 12516 -9578 12532 -9544
rect 12738 -9578 12754 -9544
rect 12974 -9578 12990 -9544
rect 13196 -9578 13212 -9544
rect 13432 -9578 13448 -9544
rect 13654 -9578 13670 -9544
rect 13890 -9578 13906 -9544
rect 14112 -9578 14128 -9544
rect 14348 -9578 14364 -9544
rect 14570 -9578 14586 -9544
rect 14806 -9578 14822 -9544
rect 15028 -9578 15044 -9544
rect 15264 -9578 15280 -9544
rect 15486 -9578 15502 -9544
rect 15722 -9578 15738 -9544
rect 10818 -10572 10918 -10410
rect 21162 -10572 21262 -10410
rect 25818 -8270 25918 -8108
rect 36162 -8270 36262 -8108
rect 26364 -8600 26380 -8566
rect 26600 -8600 26616 -8566
rect 26822 -8600 26838 -8566
rect 27058 -8600 27074 -8566
rect 27280 -8600 27296 -8566
rect 27516 -8600 27532 -8566
rect 27738 -8600 27754 -8566
rect 27974 -8600 27990 -8566
rect 28196 -8600 28212 -8566
rect 28432 -8600 28448 -8566
rect 28654 -8600 28670 -8566
rect 28890 -8600 28906 -8566
rect 29112 -8600 29128 -8566
rect 29348 -8600 29364 -8566
rect 29570 -8600 29586 -8566
rect 29806 -8600 29822 -8566
rect 30028 -8600 30044 -8566
rect 30264 -8600 30280 -8566
rect 30486 -8600 30502 -8566
rect 30722 -8600 30738 -8566
rect 31364 -8600 31380 -8566
rect 31600 -8600 31616 -8566
rect 31822 -8600 31838 -8566
rect 32058 -8600 32074 -8566
rect 32280 -8600 32296 -8566
rect 32516 -8600 32532 -8566
rect 32738 -8600 32754 -8566
rect 32974 -8600 32990 -8566
rect 33196 -8600 33212 -8566
rect 33432 -8600 33448 -8566
rect 33654 -8600 33670 -8566
rect 33890 -8600 33906 -8566
rect 34112 -8600 34128 -8566
rect 34348 -8600 34364 -8566
rect 34570 -8600 34586 -8566
rect 34806 -8600 34822 -8566
rect 35028 -8600 35044 -8566
rect 35264 -8600 35280 -8566
rect 35486 -8600 35502 -8566
rect 35722 -8600 35738 -8566
rect 26244 -8650 26278 -8634
rect 26244 -8842 26278 -8826
rect 26702 -8650 26736 -8634
rect 26702 -8842 26736 -8826
rect 27160 -8650 27194 -8634
rect 27160 -8842 27194 -8826
rect 27618 -8650 27652 -8634
rect 27618 -8842 27652 -8826
rect 28076 -8650 28110 -8634
rect 28076 -8842 28110 -8826
rect 28534 -8650 28568 -8634
rect 28534 -8842 28568 -8826
rect 28992 -8650 29026 -8634
rect 28992 -8842 29026 -8826
rect 29450 -8650 29484 -8634
rect 29450 -8842 29484 -8826
rect 29908 -8650 29942 -8634
rect 29908 -8842 29942 -8826
rect 30366 -8650 30400 -8634
rect 30366 -8842 30400 -8826
rect 30824 -8650 30858 -8634
rect 30824 -8842 30858 -8826
rect 31244 -8650 31278 -8634
rect 31244 -8842 31278 -8826
rect 31702 -8650 31736 -8634
rect 31702 -8842 31736 -8826
rect 32160 -8650 32194 -8634
rect 32160 -8842 32194 -8826
rect 32618 -8650 32652 -8634
rect 32618 -8842 32652 -8826
rect 33076 -8650 33110 -8634
rect 33076 -8842 33110 -8826
rect 33534 -8650 33568 -8634
rect 33534 -8842 33568 -8826
rect 33992 -8650 34026 -8634
rect 33992 -8842 34026 -8826
rect 34450 -8650 34484 -8634
rect 34450 -8842 34484 -8826
rect 34908 -8650 34942 -8634
rect 34908 -8842 34942 -8826
rect 35366 -8650 35400 -8634
rect 35366 -8842 35400 -8826
rect 35824 -8650 35858 -8634
rect 35824 -8842 35858 -8826
rect 26364 -8910 26380 -8876
rect 26600 -8910 26616 -8876
rect 26822 -8910 26838 -8876
rect 27058 -8910 27074 -8876
rect 27280 -8910 27296 -8876
rect 27516 -8910 27532 -8876
rect 27738 -8910 27754 -8876
rect 27974 -8910 27990 -8876
rect 28196 -8910 28212 -8876
rect 28432 -8910 28448 -8876
rect 28654 -8910 28670 -8876
rect 28890 -8910 28906 -8876
rect 29112 -8910 29128 -8876
rect 29348 -8910 29364 -8876
rect 29570 -8910 29586 -8876
rect 29806 -8910 29822 -8876
rect 30028 -8910 30044 -8876
rect 30264 -8910 30280 -8876
rect 30486 -8910 30502 -8876
rect 30722 -8910 30738 -8876
rect 31364 -8910 31380 -8876
rect 31600 -8910 31616 -8876
rect 31822 -8910 31838 -8876
rect 32058 -8910 32074 -8876
rect 32280 -8910 32296 -8876
rect 32516 -8910 32532 -8876
rect 32738 -8910 32754 -8876
rect 32974 -8910 32990 -8876
rect 33196 -8910 33212 -8876
rect 33432 -8910 33448 -8876
rect 33654 -8910 33670 -8876
rect 33890 -8910 33906 -8876
rect 34112 -8910 34128 -8876
rect 34348 -8910 34364 -8876
rect 34570 -8910 34586 -8876
rect 34806 -8910 34822 -8876
rect 35028 -8910 35044 -8876
rect 35264 -8910 35280 -8876
rect 35486 -8910 35502 -8876
rect 35722 -8910 35738 -8876
rect 26364 -9268 26380 -9234
rect 26600 -9268 26616 -9234
rect 26822 -9268 26838 -9234
rect 27058 -9268 27074 -9234
rect 27280 -9268 27296 -9234
rect 27516 -9268 27532 -9234
rect 27738 -9268 27754 -9234
rect 27974 -9268 27990 -9234
rect 28196 -9268 28212 -9234
rect 28432 -9268 28448 -9234
rect 28654 -9268 28670 -9234
rect 28890 -9268 28906 -9234
rect 29112 -9268 29128 -9234
rect 29348 -9268 29364 -9234
rect 29570 -9268 29586 -9234
rect 29806 -9268 29822 -9234
rect 30028 -9268 30044 -9234
rect 30264 -9268 30280 -9234
rect 30486 -9268 30502 -9234
rect 30722 -9268 30738 -9234
rect 26244 -9318 26278 -9302
rect 26244 -9510 26278 -9494
rect 26702 -9318 26736 -9302
rect 26702 -9510 26736 -9494
rect 27160 -9318 27194 -9302
rect 27160 -9510 27194 -9494
rect 27618 -9318 27652 -9302
rect 27618 -9510 27652 -9494
rect 28076 -9318 28110 -9302
rect 28076 -9510 28110 -9494
rect 28534 -9318 28568 -9302
rect 28534 -9510 28568 -9494
rect 28992 -9318 29026 -9302
rect 28992 -9510 29026 -9494
rect 29450 -9318 29484 -9302
rect 29450 -9510 29484 -9494
rect 29908 -9318 29942 -9302
rect 29908 -9510 29942 -9494
rect 30366 -9318 30400 -9302
rect 30366 -9510 30400 -9494
rect 30824 -9318 30858 -9302
rect 30824 -9510 30858 -9494
rect 26364 -9578 26380 -9544
rect 26600 -9578 26616 -9544
rect 26822 -9578 26838 -9544
rect 27058 -9578 27074 -9544
rect 27280 -9578 27296 -9544
rect 27516 -9578 27532 -9544
rect 27738 -9578 27754 -9544
rect 27974 -9578 27990 -9544
rect 28196 -9578 28212 -9544
rect 28432 -9578 28448 -9544
rect 28654 -9578 28670 -9544
rect 28890 -9578 28906 -9544
rect 29112 -9578 29128 -9544
rect 29348 -9578 29364 -9544
rect 29570 -9578 29586 -9544
rect 29806 -9578 29822 -9544
rect 30028 -9578 30044 -9544
rect 30264 -9578 30280 -9544
rect 30486 -9578 30502 -9544
rect 30722 -9578 30738 -9544
rect 25818 -10572 25918 -10410
rect 36162 -10572 36262 -10410
rect 14772 -11194 14872 -11032
rect 25116 -11194 25216 -11032
rect 20296 -12060 20312 -12026
rect 20532 -12060 20548 -12026
rect 20754 -12060 20770 -12026
rect 20990 -12060 21006 -12026
rect 21212 -12060 21228 -12026
rect 21448 -12060 21464 -12026
rect 21670 -12060 21686 -12026
rect 21906 -12060 21922 -12026
rect 22128 -12060 22144 -12026
rect 22364 -12060 22380 -12026
rect 22586 -12060 22602 -12026
rect 22822 -12060 22838 -12026
rect 23044 -12060 23060 -12026
rect 23280 -12060 23296 -12026
rect 23502 -12060 23518 -12026
rect 23738 -12060 23754 -12026
rect 23960 -12060 23976 -12026
rect 24196 -12060 24212 -12026
rect 24418 -12060 24434 -12026
rect 24654 -12060 24670 -12026
rect 20176 -12110 20210 -12094
rect 20176 -12302 20210 -12286
rect 20634 -12110 20668 -12094
rect 20634 -12302 20668 -12286
rect 21092 -12110 21126 -12094
rect 21092 -12302 21126 -12286
rect 21550 -12110 21584 -12094
rect 21550 -12302 21584 -12286
rect 22008 -12110 22042 -12094
rect 22008 -12302 22042 -12286
rect 22466 -12110 22500 -12094
rect 22466 -12302 22500 -12286
rect 22924 -12110 22958 -12094
rect 22924 -12302 22958 -12286
rect 23382 -12110 23416 -12094
rect 23382 -12302 23416 -12286
rect 23840 -12110 23874 -12094
rect 23840 -12302 23874 -12286
rect 24298 -12110 24332 -12094
rect 24298 -12302 24332 -12286
rect 24756 -12110 24790 -12094
rect 24756 -12302 24790 -12286
rect 20296 -12370 20312 -12336
rect 20532 -12370 20548 -12336
rect 20754 -12370 20770 -12336
rect 20990 -12370 21006 -12336
rect 21212 -12370 21228 -12336
rect 21448 -12370 21464 -12336
rect 21670 -12370 21686 -12336
rect 21906 -12370 21922 -12336
rect 22128 -12370 22144 -12336
rect 22364 -12370 22380 -12336
rect 22586 -12370 22602 -12336
rect 22822 -12370 22838 -12336
rect 23044 -12370 23060 -12336
rect 23280 -12370 23296 -12336
rect 23502 -12370 23518 -12336
rect 23738 -12370 23754 -12336
rect 23960 -12370 23976 -12336
rect 24196 -12370 24212 -12336
rect 24418 -12370 24434 -12336
rect 24654 -12370 24670 -12336
rect 15296 -12728 15312 -12694
rect 15532 -12728 15548 -12694
rect 15754 -12728 15770 -12694
rect 15990 -12728 16006 -12694
rect 16212 -12728 16228 -12694
rect 16448 -12728 16464 -12694
rect 16670 -12728 16686 -12694
rect 16906 -12728 16922 -12694
rect 17128 -12728 17144 -12694
rect 17364 -12728 17380 -12694
rect 17586 -12728 17602 -12694
rect 17822 -12728 17838 -12694
rect 18044 -12728 18060 -12694
rect 18280 -12728 18296 -12694
rect 18502 -12728 18518 -12694
rect 18738 -12728 18754 -12694
rect 18960 -12728 18976 -12694
rect 19196 -12728 19212 -12694
rect 19418 -12728 19434 -12694
rect 19654 -12728 19670 -12694
rect 20296 -12728 20312 -12694
rect 20532 -12728 20548 -12694
rect 20754 -12728 20770 -12694
rect 20990 -12728 21006 -12694
rect 21212 -12728 21228 -12694
rect 21448 -12728 21464 -12694
rect 21670 -12728 21686 -12694
rect 21906 -12728 21922 -12694
rect 22128 -12728 22144 -12694
rect 22364 -12728 22380 -12694
rect 22586 -12728 22602 -12694
rect 22822 -12728 22838 -12694
rect 23044 -12728 23060 -12694
rect 23280 -12728 23296 -12694
rect 23502 -12728 23518 -12694
rect 23738 -12728 23754 -12694
rect 23960 -12728 23976 -12694
rect 24196 -12728 24212 -12694
rect 24418 -12728 24434 -12694
rect 24654 -12728 24670 -12694
rect 15176 -12778 15210 -12762
rect 15176 -12970 15210 -12954
rect 15634 -12778 15668 -12762
rect 15634 -12970 15668 -12954
rect 16092 -12778 16126 -12762
rect 16092 -12970 16126 -12954
rect 16550 -12778 16584 -12762
rect 16550 -12970 16584 -12954
rect 17008 -12778 17042 -12762
rect 17008 -12970 17042 -12954
rect 17466 -12778 17500 -12762
rect 17466 -12970 17500 -12954
rect 17924 -12778 17958 -12762
rect 17924 -12970 17958 -12954
rect 18382 -12778 18416 -12762
rect 18382 -12970 18416 -12954
rect 18840 -12778 18874 -12762
rect 18840 -12970 18874 -12954
rect 19298 -12778 19332 -12762
rect 19298 -12970 19332 -12954
rect 19756 -12778 19790 -12762
rect 19756 -12970 19790 -12954
rect 20176 -12778 20210 -12762
rect 20176 -12970 20210 -12954
rect 20634 -12778 20668 -12762
rect 20634 -12970 20668 -12954
rect 21092 -12778 21126 -12762
rect 21092 -12970 21126 -12954
rect 21550 -12778 21584 -12762
rect 21550 -12970 21584 -12954
rect 22008 -12778 22042 -12762
rect 22008 -12970 22042 -12954
rect 22466 -12778 22500 -12762
rect 22466 -12970 22500 -12954
rect 22924 -12778 22958 -12762
rect 22924 -12970 22958 -12954
rect 23382 -12778 23416 -12762
rect 23382 -12970 23416 -12954
rect 23840 -12778 23874 -12762
rect 23840 -12970 23874 -12954
rect 24298 -12778 24332 -12762
rect 24298 -12970 24332 -12954
rect 24756 -12778 24790 -12762
rect 24756 -12970 24790 -12954
rect 15296 -13038 15312 -13004
rect 15532 -13038 15548 -13004
rect 15754 -13038 15770 -13004
rect 15990 -13038 16006 -13004
rect 16212 -13038 16228 -13004
rect 16448 -13038 16464 -13004
rect 16670 -13038 16686 -13004
rect 16906 -13038 16922 -13004
rect 17128 -13038 17144 -13004
rect 17364 -13038 17380 -13004
rect 17586 -13038 17602 -13004
rect 17822 -13038 17838 -13004
rect 18044 -13038 18060 -13004
rect 18280 -13038 18296 -13004
rect 18502 -13038 18518 -13004
rect 18738 -13038 18754 -13004
rect 18960 -13038 18976 -13004
rect 19196 -13038 19212 -13004
rect 19418 -13038 19434 -13004
rect 19654 -13038 19670 -13004
rect 20296 -13038 20312 -13004
rect 20532 -13038 20548 -13004
rect 20754 -13038 20770 -13004
rect 20990 -13038 21006 -13004
rect 21212 -13038 21228 -13004
rect 21448 -13038 21464 -13004
rect 21670 -13038 21686 -13004
rect 21906 -13038 21922 -13004
rect 22128 -13038 22144 -13004
rect 22364 -13038 22380 -13004
rect 22586 -13038 22602 -13004
rect 22822 -13038 22838 -13004
rect 23044 -13038 23060 -13004
rect 23280 -13038 23296 -13004
rect 23502 -13038 23518 -13004
rect 23738 -13038 23754 -13004
rect 23960 -13038 23976 -13004
rect 24196 -13038 24212 -13004
rect 24418 -13038 24434 -13004
rect 24654 -13038 24670 -13004
rect 14772 -13496 14872 -13334
rect 25116 -13496 25216 -13334
rect 29772 -11194 29872 -11032
rect 40116 -11194 40216 -11032
rect 35296 -12060 35312 -12026
rect 35532 -12060 35548 -12026
rect 35754 -12060 35770 -12026
rect 35990 -12060 36006 -12026
rect 36212 -12060 36228 -12026
rect 36448 -12060 36464 -12026
rect 36670 -12060 36686 -12026
rect 36906 -12060 36922 -12026
rect 37128 -12060 37144 -12026
rect 37364 -12060 37380 -12026
rect 37586 -12060 37602 -12026
rect 37822 -12060 37838 -12026
rect 38044 -12060 38060 -12026
rect 38280 -12060 38296 -12026
rect 38502 -12060 38518 -12026
rect 38738 -12060 38754 -12026
rect 38960 -12060 38976 -12026
rect 39196 -12060 39212 -12026
rect 39418 -12060 39434 -12026
rect 39654 -12060 39670 -12026
rect 35176 -12110 35210 -12094
rect 35176 -12302 35210 -12286
rect 35634 -12110 35668 -12094
rect 35634 -12302 35668 -12286
rect 36092 -12110 36126 -12094
rect 36092 -12302 36126 -12286
rect 36550 -12110 36584 -12094
rect 36550 -12302 36584 -12286
rect 37008 -12110 37042 -12094
rect 37008 -12302 37042 -12286
rect 37466 -12110 37500 -12094
rect 37466 -12302 37500 -12286
rect 37924 -12110 37958 -12094
rect 37924 -12302 37958 -12286
rect 38382 -12110 38416 -12094
rect 38382 -12302 38416 -12286
rect 38840 -12110 38874 -12094
rect 38840 -12302 38874 -12286
rect 39298 -12110 39332 -12094
rect 39298 -12302 39332 -12286
rect 39756 -12110 39790 -12094
rect 39756 -12302 39790 -12286
rect 35296 -12370 35312 -12336
rect 35532 -12370 35548 -12336
rect 35754 -12370 35770 -12336
rect 35990 -12370 36006 -12336
rect 36212 -12370 36228 -12336
rect 36448 -12370 36464 -12336
rect 36670 -12370 36686 -12336
rect 36906 -12370 36922 -12336
rect 37128 -12370 37144 -12336
rect 37364 -12370 37380 -12336
rect 37586 -12370 37602 -12336
rect 37822 -12370 37838 -12336
rect 38044 -12370 38060 -12336
rect 38280 -12370 38296 -12336
rect 38502 -12370 38518 -12336
rect 38738 -12370 38754 -12336
rect 38960 -12370 38976 -12336
rect 39196 -12370 39212 -12336
rect 39418 -12370 39434 -12336
rect 39654 -12370 39670 -12336
rect 30296 -12728 30312 -12694
rect 30532 -12728 30548 -12694
rect 30754 -12728 30770 -12694
rect 30990 -12728 31006 -12694
rect 31212 -12728 31228 -12694
rect 31448 -12728 31464 -12694
rect 31670 -12728 31686 -12694
rect 31906 -12728 31922 -12694
rect 32128 -12728 32144 -12694
rect 32364 -12728 32380 -12694
rect 32586 -12728 32602 -12694
rect 32822 -12728 32838 -12694
rect 33044 -12728 33060 -12694
rect 33280 -12728 33296 -12694
rect 33502 -12728 33518 -12694
rect 33738 -12728 33754 -12694
rect 33960 -12728 33976 -12694
rect 34196 -12728 34212 -12694
rect 34418 -12728 34434 -12694
rect 34654 -12728 34670 -12694
rect 35296 -12728 35312 -12694
rect 35532 -12728 35548 -12694
rect 35754 -12728 35770 -12694
rect 35990 -12728 36006 -12694
rect 36212 -12728 36228 -12694
rect 36448 -12728 36464 -12694
rect 36670 -12728 36686 -12694
rect 36906 -12728 36922 -12694
rect 37128 -12728 37144 -12694
rect 37364 -12728 37380 -12694
rect 37586 -12728 37602 -12694
rect 37822 -12728 37838 -12694
rect 38044 -12728 38060 -12694
rect 38280 -12728 38296 -12694
rect 38502 -12728 38518 -12694
rect 38738 -12728 38754 -12694
rect 38960 -12728 38976 -12694
rect 39196 -12728 39212 -12694
rect 39418 -12728 39434 -12694
rect 39654 -12728 39670 -12694
rect 30176 -12778 30210 -12762
rect 30176 -12970 30210 -12954
rect 30634 -12778 30668 -12762
rect 30634 -12970 30668 -12954
rect 31092 -12778 31126 -12762
rect 31092 -12970 31126 -12954
rect 31550 -12778 31584 -12762
rect 31550 -12970 31584 -12954
rect 32008 -12778 32042 -12762
rect 32008 -12970 32042 -12954
rect 32466 -12778 32500 -12762
rect 32466 -12970 32500 -12954
rect 32924 -12778 32958 -12762
rect 32924 -12970 32958 -12954
rect 33382 -12778 33416 -12762
rect 33382 -12970 33416 -12954
rect 33840 -12778 33874 -12762
rect 33840 -12970 33874 -12954
rect 34298 -12778 34332 -12762
rect 34298 -12970 34332 -12954
rect 34756 -12778 34790 -12762
rect 34756 -12970 34790 -12954
rect 35176 -12778 35210 -12762
rect 35176 -12970 35210 -12954
rect 35634 -12778 35668 -12762
rect 35634 -12970 35668 -12954
rect 36092 -12778 36126 -12762
rect 36092 -12970 36126 -12954
rect 36550 -12778 36584 -12762
rect 36550 -12970 36584 -12954
rect 37008 -12778 37042 -12762
rect 37008 -12970 37042 -12954
rect 37466 -12778 37500 -12762
rect 37466 -12970 37500 -12954
rect 37924 -12778 37958 -12762
rect 37924 -12970 37958 -12954
rect 38382 -12778 38416 -12762
rect 38382 -12970 38416 -12954
rect 38840 -12778 38874 -12762
rect 38840 -12970 38874 -12954
rect 39298 -12778 39332 -12762
rect 39298 -12970 39332 -12954
rect 39756 -12778 39790 -12762
rect 39756 -12970 39790 -12954
rect 30296 -13038 30312 -13004
rect 30532 -13038 30548 -13004
rect 30754 -13038 30770 -13004
rect 30990 -13038 31006 -13004
rect 31212 -13038 31228 -13004
rect 31448 -13038 31464 -13004
rect 31670 -13038 31686 -13004
rect 31906 -13038 31922 -13004
rect 32128 -13038 32144 -13004
rect 32364 -13038 32380 -13004
rect 32586 -13038 32602 -13004
rect 32822 -13038 32838 -13004
rect 33044 -13038 33060 -13004
rect 33280 -13038 33296 -13004
rect 33502 -13038 33518 -13004
rect 33738 -13038 33754 -13004
rect 33960 -13038 33976 -13004
rect 34196 -13038 34212 -13004
rect 34418 -13038 34434 -13004
rect 34654 -13038 34670 -13004
rect 35296 -13038 35312 -13004
rect 35532 -13038 35548 -13004
rect 35754 -13038 35770 -13004
rect 35990 -13038 36006 -13004
rect 36212 -13038 36228 -13004
rect 36448 -13038 36464 -13004
rect 36670 -13038 36686 -13004
rect 36906 -13038 36922 -13004
rect 37128 -13038 37144 -13004
rect 37364 -13038 37380 -13004
rect 37586 -13038 37602 -13004
rect 37822 -13038 37838 -13004
rect 38044 -13038 38060 -13004
rect 38280 -13038 38296 -13004
rect 38502 -13038 38518 -13004
rect 38738 -13038 38754 -13004
rect 38960 -13038 38976 -13004
rect 39196 -13038 39212 -13004
rect 39418 -13038 39434 -13004
rect 39654 -13038 39670 -13004
rect 29772 -13496 29872 -13334
rect 40116 -13496 40216 -13334
rect 14772 -13894 14872 -13732
rect 25116 -13894 25216 -13732
rect 15295 -14212 15311 -14178
rect 15531 -14212 15547 -14178
rect 15753 -14212 15769 -14178
rect 15989 -14212 16005 -14178
rect 16211 -14212 16227 -14178
rect 16447 -14212 16463 -14178
rect 16669 -14212 16685 -14178
rect 16905 -14212 16921 -14178
rect 17127 -14212 17143 -14178
rect 17363 -14212 17379 -14178
rect 17585 -14212 17601 -14178
rect 17821 -14212 17837 -14178
rect 18043 -14212 18059 -14178
rect 18279 -14212 18295 -14178
rect 18501 -14212 18517 -14178
rect 18737 -14212 18753 -14178
rect 18959 -14212 18975 -14178
rect 19195 -14212 19211 -14178
rect 19417 -14212 19433 -14178
rect 19653 -14212 19669 -14178
rect 20295 -14212 20311 -14178
rect 20531 -14212 20547 -14178
rect 20753 -14212 20769 -14178
rect 20989 -14212 21005 -14178
rect 21211 -14212 21227 -14178
rect 21447 -14212 21463 -14178
rect 21669 -14212 21685 -14178
rect 21905 -14212 21921 -14178
rect 22127 -14212 22143 -14178
rect 22363 -14212 22379 -14178
rect 22585 -14212 22601 -14178
rect 22821 -14212 22837 -14178
rect 23043 -14212 23059 -14178
rect 23279 -14212 23295 -14178
rect 23501 -14212 23517 -14178
rect 23737 -14212 23753 -14178
rect 23959 -14212 23975 -14178
rect 24195 -14212 24211 -14178
rect 24417 -14212 24433 -14178
rect 24653 -14212 24669 -14178
rect 15175 -14271 15209 -14255
rect 15175 -15463 15209 -15447
rect 15633 -14271 15667 -14255
rect 15633 -15463 15667 -15447
rect 16091 -14271 16125 -14255
rect 16091 -15463 16125 -15447
rect 16549 -14271 16583 -14255
rect 16549 -15463 16583 -15447
rect 17007 -14271 17041 -14255
rect 17007 -15463 17041 -15447
rect 17465 -14271 17499 -14255
rect 17465 -15463 17499 -15447
rect 17923 -14271 17957 -14255
rect 17923 -15463 17957 -15447
rect 18381 -14271 18415 -14255
rect 18381 -15463 18415 -15447
rect 18839 -14271 18873 -14255
rect 18839 -15463 18873 -15447
rect 19297 -14271 19331 -14255
rect 19297 -15463 19331 -15447
rect 19755 -14271 19789 -14255
rect 19755 -15463 19789 -15447
rect 20175 -14271 20209 -14255
rect 20175 -15463 20209 -15447
rect 20633 -14271 20667 -14255
rect 20633 -15463 20667 -15447
rect 21091 -14271 21125 -14255
rect 21091 -15463 21125 -15447
rect 21549 -14271 21583 -14255
rect 21549 -15463 21583 -15447
rect 22007 -14271 22041 -14255
rect 22007 -15463 22041 -15447
rect 22465 -14271 22499 -14255
rect 22465 -15463 22499 -15447
rect 22923 -14271 22957 -14255
rect 22923 -15463 22957 -15447
rect 23381 -14271 23415 -14255
rect 23381 -15463 23415 -15447
rect 23839 -14271 23873 -14255
rect 23839 -15463 23873 -15447
rect 24297 -14271 24331 -14255
rect 24297 -15463 24331 -15447
rect 24755 -14271 24789 -14255
rect 24755 -15463 24789 -15447
rect 15295 -15540 15311 -15506
rect 15531 -15540 15547 -15506
rect 15753 -15540 15769 -15506
rect 15989 -15540 16005 -15506
rect 16211 -15540 16227 -15506
rect 16447 -15540 16463 -15506
rect 16669 -15540 16685 -15506
rect 16905 -15540 16921 -15506
rect 17127 -15540 17143 -15506
rect 17363 -15540 17379 -15506
rect 17585 -15540 17601 -15506
rect 17821 -15540 17837 -15506
rect 18043 -15540 18059 -15506
rect 18279 -15540 18295 -15506
rect 18501 -15540 18517 -15506
rect 18737 -15540 18753 -15506
rect 18959 -15540 18975 -15506
rect 19195 -15540 19211 -15506
rect 19417 -15540 19433 -15506
rect 19653 -15540 19669 -15506
rect 20295 -15540 20311 -15506
rect 20531 -15540 20547 -15506
rect 20753 -15540 20769 -15506
rect 20989 -15540 21005 -15506
rect 21211 -15540 21227 -15506
rect 21447 -15540 21463 -15506
rect 21669 -15540 21685 -15506
rect 21905 -15540 21921 -15506
rect 22127 -15540 22143 -15506
rect 22363 -15540 22379 -15506
rect 22585 -15540 22601 -15506
rect 22821 -15540 22837 -15506
rect 23043 -15540 23059 -15506
rect 23279 -15540 23295 -15506
rect 23501 -15540 23517 -15506
rect 23737 -15540 23753 -15506
rect 23959 -15540 23975 -15506
rect 24195 -15540 24211 -15506
rect 24417 -15540 24433 -15506
rect 24653 -15540 24669 -15506
rect 19892 -16312 20352 -16306
rect 19892 -16360 20298 -16312
rect 20346 -16360 20352 -16312
rect 19892 -16366 20352 -16360
rect 16072 -16477 16088 -16443
rect 16308 -16477 16324 -16443
rect 16530 -16477 16546 -16443
rect 16766 -16477 16782 -16443
rect 16988 -16477 17004 -16443
rect 17224 -16477 17240 -16443
rect 17446 -16477 17462 -16443
rect 17682 -16477 17698 -16443
rect 17904 -16477 17920 -16443
rect 18140 -16477 18156 -16443
rect 18362 -16477 18378 -16443
rect 18598 -16477 18614 -16443
rect 18820 -16477 18836 -16443
rect 19056 -16477 19072 -16443
rect 19278 -16477 19294 -16443
rect 19514 -16477 19530 -16443
rect 19736 -16477 19752 -16443
rect 19972 -16477 19988 -16443
rect 20194 -16477 20210 -16443
rect 20430 -16477 20446 -16443
rect 20652 -16477 20668 -16443
rect 20888 -16477 20904 -16443
rect 21110 -16477 21126 -16443
rect 21346 -16477 21362 -16443
rect 21568 -16477 21584 -16443
rect 21804 -16477 21820 -16443
rect 22026 -16477 22042 -16443
rect 22262 -16477 22278 -16443
rect 22484 -16477 22500 -16443
rect 22720 -16477 22736 -16443
rect 22942 -16477 22958 -16443
rect 23178 -16477 23194 -16443
rect 23400 -16477 23416 -16443
rect 23636 -16477 23652 -16443
rect 23858 -16477 23874 -16443
rect 24094 -16477 24110 -16443
rect 15952 -16536 15986 -16520
rect 15952 -18128 15986 -18112
rect 16410 -16536 16444 -16520
rect 16410 -18128 16444 -18112
rect 16868 -16536 16902 -16520
rect 16868 -18128 16902 -18112
rect 17326 -16536 17360 -16520
rect 17326 -18128 17360 -18112
rect 17784 -16536 17818 -16520
rect 17784 -18128 17818 -18112
rect 18242 -16536 18276 -16520
rect 18242 -18128 18276 -18112
rect 18700 -16536 18734 -16520
rect 18700 -18128 18734 -18112
rect 19158 -16536 19192 -16520
rect 19158 -18128 19192 -18112
rect 19616 -16536 19650 -16520
rect 19616 -18128 19650 -18112
rect 20074 -16536 20108 -16520
rect 20074 -18128 20108 -18112
rect 20532 -16536 20566 -16520
rect 20532 -18128 20566 -18112
rect 20990 -16536 21024 -16520
rect 20990 -18128 21024 -18112
rect 21448 -16536 21482 -16520
rect 21448 -18128 21482 -18112
rect 21906 -16536 21940 -16520
rect 21906 -18128 21940 -18112
rect 22364 -16536 22398 -16520
rect 22364 -18128 22398 -18112
rect 22822 -16536 22856 -16520
rect 22822 -18128 22856 -18112
rect 23280 -16536 23314 -16520
rect 23280 -18128 23314 -18112
rect 23738 -16536 23772 -16520
rect 23738 -18128 23772 -18112
rect 24196 -16536 24230 -16520
rect 24196 -18128 24230 -18112
rect 16072 -18205 16088 -18171
rect 16308 -18205 16324 -18171
rect 16530 -18205 16546 -18171
rect 16766 -18205 16782 -18171
rect 16988 -18205 17004 -18171
rect 17224 -18205 17240 -18171
rect 17446 -18205 17462 -18171
rect 17682 -18205 17698 -18171
rect 17904 -18205 17920 -18171
rect 18140 -18205 18156 -18171
rect 18362 -18205 18378 -18171
rect 18598 -18205 18614 -18171
rect 18820 -18205 18836 -18171
rect 19056 -18205 19072 -18171
rect 19278 -18205 19294 -18171
rect 19514 -18205 19530 -18171
rect 19736 -18205 19752 -18171
rect 19972 -18205 19988 -18171
rect 20194 -18205 20210 -18171
rect 20430 -18205 20446 -18171
rect 20652 -18205 20668 -18171
rect 20888 -18205 20904 -18171
rect 21110 -18205 21126 -18171
rect 21346 -18205 21362 -18171
rect 21568 -18205 21584 -18171
rect 21804 -18205 21820 -18171
rect 22026 -18205 22042 -18171
rect 22262 -18205 22278 -18171
rect 22484 -18205 22500 -18171
rect 22720 -18205 22736 -18171
rect 22942 -18205 22958 -18171
rect 23178 -18205 23194 -18171
rect 23400 -18205 23416 -18171
rect 23636 -18205 23652 -18171
rect 23858 -18205 23874 -18171
rect 24094 -18205 24110 -18171
rect 14772 -19576 14872 -19414
rect 25116 -19576 25216 -19414
rect 29772 -13894 29872 -13732
rect 40116 -13894 40216 -13732
rect 30295 -14212 30311 -14178
rect 30531 -14212 30547 -14178
rect 30753 -14212 30769 -14178
rect 30989 -14212 31005 -14178
rect 31211 -14212 31227 -14178
rect 31447 -14212 31463 -14178
rect 31669 -14212 31685 -14178
rect 31905 -14212 31921 -14178
rect 32127 -14212 32143 -14178
rect 32363 -14212 32379 -14178
rect 32585 -14212 32601 -14178
rect 32821 -14212 32837 -14178
rect 33043 -14212 33059 -14178
rect 33279 -14212 33295 -14178
rect 33501 -14212 33517 -14178
rect 33737 -14212 33753 -14178
rect 33959 -14212 33975 -14178
rect 34195 -14212 34211 -14178
rect 34417 -14212 34433 -14178
rect 34653 -14212 34669 -14178
rect 35295 -14212 35311 -14178
rect 35531 -14212 35547 -14178
rect 35753 -14212 35769 -14178
rect 35989 -14212 36005 -14178
rect 36211 -14212 36227 -14178
rect 36447 -14212 36463 -14178
rect 36669 -14212 36685 -14178
rect 36905 -14212 36921 -14178
rect 37127 -14212 37143 -14178
rect 37363 -14212 37379 -14178
rect 37585 -14212 37601 -14178
rect 37821 -14212 37837 -14178
rect 38043 -14212 38059 -14178
rect 38279 -14212 38295 -14178
rect 38501 -14212 38517 -14178
rect 38737 -14212 38753 -14178
rect 38959 -14212 38975 -14178
rect 39195 -14212 39211 -14178
rect 39417 -14212 39433 -14178
rect 39653 -14212 39669 -14178
rect 30175 -14271 30209 -14255
rect 30175 -15463 30209 -15447
rect 30633 -14271 30667 -14255
rect 30633 -15463 30667 -15447
rect 31091 -14271 31125 -14255
rect 31091 -15463 31125 -15447
rect 31549 -14271 31583 -14255
rect 31549 -15463 31583 -15447
rect 32007 -14271 32041 -14255
rect 32007 -15463 32041 -15447
rect 32465 -14271 32499 -14255
rect 32465 -15463 32499 -15447
rect 32923 -14271 32957 -14255
rect 32923 -15463 32957 -15447
rect 33381 -14271 33415 -14255
rect 33381 -15463 33415 -15447
rect 33839 -14271 33873 -14255
rect 33839 -15463 33873 -15447
rect 34297 -14271 34331 -14255
rect 34297 -15463 34331 -15447
rect 34755 -14271 34789 -14255
rect 34755 -15463 34789 -15447
rect 35175 -14271 35209 -14255
rect 35175 -15463 35209 -15447
rect 35633 -14271 35667 -14255
rect 35633 -15463 35667 -15447
rect 36091 -14271 36125 -14255
rect 36091 -15463 36125 -15447
rect 36549 -14271 36583 -14255
rect 36549 -15463 36583 -15447
rect 37007 -14271 37041 -14255
rect 37007 -15463 37041 -15447
rect 37465 -14271 37499 -14255
rect 37465 -15463 37499 -15447
rect 37923 -14271 37957 -14255
rect 37923 -15463 37957 -15447
rect 38381 -14271 38415 -14255
rect 38381 -15463 38415 -15447
rect 38839 -14271 38873 -14255
rect 38839 -15463 38873 -15447
rect 39297 -14271 39331 -14255
rect 39297 -15463 39331 -15447
rect 39755 -14271 39789 -14255
rect 39755 -15463 39789 -15447
rect 30295 -15540 30311 -15506
rect 30531 -15540 30547 -15506
rect 30753 -15540 30769 -15506
rect 30989 -15540 31005 -15506
rect 31211 -15540 31227 -15506
rect 31447 -15540 31463 -15506
rect 31669 -15540 31685 -15506
rect 31905 -15540 31921 -15506
rect 32127 -15540 32143 -15506
rect 32363 -15540 32379 -15506
rect 32585 -15540 32601 -15506
rect 32821 -15540 32837 -15506
rect 33043 -15540 33059 -15506
rect 33279 -15540 33295 -15506
rect 33501 -15540 33517 -15506
rect 33737 -15540 33753 -15506
rect 33959 -15540 33975 -15506
rect 34195 -15540 34211 -15506
rect 34417 -15540 34433 -15506
rect 34653 -15540 34669 -15506
rect 35295 -15540 35311 -15506
rect 35531 -15540 35547 -15506
rect 35753 -15540 35769 -15506
rect 35989 -15540 36005 -15506
rect 36211 -15540 36227 -15506
rect 36447 -15540 36463 -15506
rect 36669 -15540 36685 -15506
rect 36905 -15540 36921 -15506
rect 37127 -15540 37143 -15506
rect 37363 -15540 37379 -15506
rect 37585 -15540 37601 -15506
rect 37821 -15540 37837 -15506
rect 38043 -15540 38059 -15506
rect 38279 -15540 38295 -15506
rect 38501 -15540 38517 -15506
rect 38737 -15540 38753 -15506
rect 38959 -15540 38975 -15506
rect 39195 -15540 39211 -15506
rect 39417 -15540 39433 -15506
rect 39653 -15540 39669 -15506
rect 34892 -16312 35352 -16306
rect 34892 -16360 35298 -16312
rect 35346 -16360 35352 -16312
rect 34892 -16366 35352 -16360
rect 31072 -16477 31088 -16443
rect 31308 -16477 31324 -16443
rect 31530 -16477 31546 -16443
rect 31766 -16477 31782 -16443
rect 31988 -16477 32004 -16443
rect 32224 -16477 32240 -16443
rect 32446 -16477 32462 -16443
rect 32682 -16477 32698 -16443
rect 32904 -16477 32920 -16443
rect 33140 -16477 33156 -16443
rect 33362 -16477 33378 -16443
rect 33598 -16477 33614 -16443
rect 33820 -16477 33836 -16443
rect 34056 -16477 34072 -16443
rect 34278 -16477 34294 -16443
rect 34514 -16477 34530 -16443
rect 34736 -16477 34752 -16443
rect 34972 -16477 34988 -16443
rect 35194 -16477 35210 -16443
rect 35430 -16477 35446 -16443
rect 35652 -16477 35668 -16443
rect 35888 -16477 35904 -16443
rect 36110 -16477 36126 -16443
rect 36346 -16477 36362 -16443
rect 36568 -16477 36584 -16443
rect 36804 -16477 36820 -16443
rect 37026 -16477 37042 -16443
rect 37262 -16477 37278 -16443
rect 37484 -16477 37500 -16443
rect 37720 -16477 37736 -16443
rect 37942 -16477 37958 -16443
rect 38178 -16477 38194 -16443
rect 38400 -16477 38416 -16443
rect 38636 -16477 38652 -16443
rect 38858 -16477 38874 -16443
rect 39094 -16477 39110 -16443
rect 30952 -16536 30986 -16520
rect 30952 -18128 30986 -18112
rect 31410 -16536 31444 -16520
rect 31410 -18128 31444 -18112
rect 31868 -16536 31902 -16520
rect 31868 -18128 31902 -18112
rect 32326 -16536 32360 -16520
rect 32326 -18128 32360 -18112
rect 32784 -16536 32818 -16520
rect 32784 -18128 32818 -18112
rect 33242 -16536 33276 -16520
rect 33242 -18128 33276 -18112
rect 33700 -16536 33734 -16520
rect 33700 -18128 33734 -18112
rect 34158 -16536 34192 -16520
rect 34158 -18128 34192 -18112
rect 34616 -16536 34650 -16520
rect 34616 -18128 34650 -18112
rect 35074 -16536 35108 -16520
rect 35074 -18128 35108 -18112
rect 35532 -16536 35566 -16520
rect 35532 -18128 35566 -18112
rect 35990 -16536 36024 -16520
rect 35990 -18128 36024 -18112
rect 36448 -16536 36482 -16520
rect 36448 -18128 36482 -18112
rect 36906 -16536 36940 -16520
rect 36906 -18128 36940 -18112
rect 37364 -16536 37398 -16520
rect 37364 -18128 37398 -18112
rect 37822 -16536 37856 -16520
rect 37822 -18128 37856 -18112
rect 38280 -16536 38314 -16520
rect 38280 -18128 38314 -18112
rect 38738 -16536 38772 -16520
rect 38738 -18128 38772 -18112
rect 39196 -16536 39230 -16520
rect 39196 -18128 39230 -18112
rect 31072 -18205 31088 -18171
rect 31308 -18205 31324 -18171
rect 31530 -18205 31546 -18171
rect 31766 -18205 31782 -18171
rect 31988 -18205 32004 -18171
rect 32224 -18205 32240 -18171
rect 32446 -18205 32462 -18171
rect 32682 -18205 32698 -18171
rect 32904 -18205 32920 -18171
rect 33140 -18205 33156 -18171
rect 33362 -18205 33378 -18171
rect 33598 -18205 33614 -18171
rect 33820 -18205 33836 -18171
rect 34056 -18205 34072 -18171
rect 34278 -18205 34294 -18171
rect 34514 -18205 34530 -18171
rect 34736 -18205 34752 -18171
rect 34972 -18205 34988 -18171
rect 35194 -18205 35210 -18171
rect 35430 -18205 35446 -18171
rect 35652 -18205 35668 -18171
rect 35888 -18205 35904 -18171
rect 36110 -18205 36126 -18171
rect 36346 -18205 36362 -18171
rect 36568 -18205 36584 -18171
rect 36804 -18205 36820 -18171
rect 37026 -18205 37042 -18171
rect 37262 -18205 37278 -18171
rect 37484 -18205 37500 -18171
rect 37720 -18205 37736 -18171
rect 37942 -18205 37958 -18171
rect 38178 -18205 38194 -18171
rect 38400 -18205 38416 -18171
rect 38636 -18205 38652 -18171
rect 38858 -18205 38874 -18171
rect 39094 -18205 39110 -18171
rect 29772 -19576 29872 -19414
rect 40116 -19576 40216 -19414
rect 10818 -20190 10918 -20028
rect 21162 -20190 21262 -20028
rect 11924 -21433 11940 -21399
rect 12160 -21433 12176 -21399
rect 12382 -21433 12398 -21399
rect 12618 -21433 12634 -21399
rect 12840 -21433 12856 -21399
rect 13076 -21433 13092 -21399
rect 13298 -21433 13314 -21399
rect 13534 -21433 13550 -21399
rect 13756 -21433 13772 -21399
rect 13992 -21433 14008 -21399
rect 14214 -21433 14230 -21399
rect 14450 -21433 14466 -21399
rect 14672 -21433 14688 -21399
rect 14908 -21433 14924 -21399
rect 15130 -21433 15146 -21399
rect 15366 -21433 15382 -21399
rect 15588 -21433 15604 -21399
rect 15824 -21433 15840 -21399
rect 16046 -21433 16062 -21399
rect 16282 -21433 16298 -21399
rect 16504 -21433 16520 -21399
rect 16740 -21433 16756 -21399
rect 16962 -21433 16978 -21399
rect 17198 -21433 17214 -21399
rect 17420 -21433 17436 -21399
rect 17656 -21433 17672 -21399
rect 17878 -21433 17894 -21399
rect 18114 -21433 18130 -21399
rect 18336 -21433 18352 -21399
rect 18572 -21433 18588 -21399
rect 18794 -21433 18810 -21399
rect 19030 -21433 19046 -21399
rect 19252 -21433 19268 -21399
rect 19488 -21433 19504 -21399
rect 19710 -21433 19726 -21399
rect 19946 -21433 19962 -21399
rect 11804 -21492 11838 -21476
rect 11804 -23084 11838 -23068
rect 12262 -21492 12296 -21476
rect 12262 -23084 12296 -23068
rect 12720 -21492 12754 -21476
rect 12720 -23084 12754 -23068
rect 13178 -21492 13212 -21476
rect 13178 -23084 13212 -23068
rect 13636 -21492 13670 -21476
rect 13636 -23084 13670 -23068
rect 14094 -21492 14128 -21476
rect 14094 -23084 14128 -23068
rect 14552 -21492 14586 -21476
rect 14552 -23084 14586 -23068
rect 15010 -21492 15044 -21476
rect 15010 -23084 15044 -23068
rect 15468 -21492 15502 -21476
rect 15468 -23084 15502 -23068
rect 15926 -21492 15960 -21476
rect 15926 -23084 15960 -23068
rect 16384 -21492 16418 -21476
rect 16384 -23084 16418 -23068
rect 16842 -21492 16876 -21476
rect 16842 -23084 16876 -23068
rect 17300 -21492 17334 -21476
rect 17300 -23084 17334 -23068
rect 17758 -21492 17792 -21476
rect 17758 -23084 17792 -23068
rect 18216 -21492 18250 -21476
rect 18216 -23084 18250 -23068
rect 18674 -21492 18708 -21476
rect 18674 -23084 18708 -23068
rect 19132 -21492 19166 -21476
rect 19132 -23084 19166 -23068
rect 19590 -21492 19624 -21476
rect 19590 -23084 19624 -23068
rect 20048 -21492 20082 -21476
rect 20048 -23084 20082 -23068
rect 11924 -23161 11940 -23127
rect 12160 -23161 12176 -23127
rect 12382 -23161 12398 -23127
rect 12618 -23161 12634 -23127
rect 12840 -23161 12856 -23127
rect 13076 -23161 13092 -23127
rect 13298 -23161 13314 -23127
rect 13534 -23161 13550 -23127
rect 13756 -23161 13772 -23127
rect 13992 -23161 14008 -23127
rect 14214 -23161 14230 -23127
rect 14450 -23161 14466 -23127
rect 14672 -23161 14688 -23127
rect 14908 -23161 14924 -23127
rect 15130 -23161 15146 -23127
rect 15366 -23161 15382 -23127
rect 15588 -23161 15604 -23127
rect 15824 -23161 15840 -23127
rect 16046 -23161 16062 -23127
rect 16282 -23161 16298 -23127
rect 16504 -23161 16520 -23127
rect 16740 -23161 16756 -23127
rect 16962 -23161 16978 -23127
rect 17198 -23161 17214 -23127
rect 17420 -23161 17436 -23127
rect 17656 -23161 17672 -23127
rect 17878 -23161 17894 -23127
rect 18114 -23161 18130 -23127
rect 18336 -23161 18352 -23127
rect 18572 -23161 18588 -23127
rect 18794 -23161 18810 -23127
rect 19030 -23161 19046 -23127
rect 19252 -23161 19268 -23127
rect 19488 -23161 19504 -23127
rect 19710 -23161 19726 -23127
rect 19946 -23161 19962 -23127
rect 15682 -23244 16142 -23238
rect 15682 -23292 15688 -23244
rect 15736 -23292 16142 -23244
rect 15682 -23298 16142 -23292
rect 11365 -24098 11381 -24064
rect 11601 -24098 11617 -24064
rect 11823 -24098 11839 -24064
rect 12059 -24098 12075 -24064
rect 12281 -24098 12297 -24064
rect 12517 -24098 12533 -24064
rect 12739 -24098 12755 -24064
rect 12975 -24098 12991 -24064
rect 13197 -24098 13213 -24064
rect 13433 -24098 13449 -24064
rect 13655 -24098 13671 -24064
rect 13891 -24098 13907 -24064
rect 14113 -24098 14129 -24064
rect 14349 -24098 14365 -24064
rect 14571 -24098 14587 -24064
rect 14807 -24098 14823 -24064
rect 15029 -24098 15045 -24064
rect 15265 -24098 15281 -24064
rect 15487 -24098 15503 -24064
rect 15723 -24098 15739 -24064
rect 16365 -24098 16381 -24064
rect 16601 -24098 16617 -24064
rect 16823 -24098 16839 -24064
rect 17059 -24098 17075 -24064
rect 17281 -24098 17297 -24064
rect 17517 -24098 17533 -24064
rect 17739 -24098 17755 -24064
rect 17975 -24098 17991 -24064
rect 18197 -24098 18213 -24064
rect 18433 -24098 18449 -24064
rect 18655 -24098 18671 -24064
rect 18891 -24098 18907 -24064
rect 19113 -24098 19129 -24064
rect 19349 -24098 19365 -24064
rect 19571 -24098 19587 -24064
rect 19807 -24098 19823 -24064
rect 20029 -24098 20045 -24064
rect 20265 -24098 20281 -24064
rect 20487 -24098 20503 -24064
rect 20723 -24098 20739 -24064
rect 11245 -24157 11279 -24141
rect 11245 -25349 11279 -25333
rect 11703 -24157 11737 -24141
rect 11703 -25349 11737 -25333
rect 12161 -24157 12195 -24141
rect 12161 -25349 12195 -25333
rect 12619 -24157 12653 -24141
rect 12619 -25349 12653 -25333
rect 13077 -24157 13111 -24141
rect 13077 -25349 13111 -25333
rect 13535 -24157 13569 -24141
rect 13535 -25349 13569 -25333
rect 13993 -24157 14027 -24141
rect 13993 -25349 14027 -25333
rect 14451 -24157 14485 -24141
rect 14451 -25349 14485 -25333
rect 14909 -24157 14943 -24141
rect 14909 -25349 14943 -25333
rect 15367 -24157 15401 -24141
rect 15367 -25349 15401 -25333
rect 15825 -24157 15859 -24141
rect 15825 -25349 15859 -25333
rect 16245 -24157 16279 -24141
rect 16245 -25349 16279 -25333
rect 16703 -24157 16737 -24141
rect 16703 -25349 16737 -25333
rect 17161 -24157 17195 -24141
rect 17161 -25349 17195 -25333
rect 17619 -24157 17653 -24141
rect 17619 -25349 17653 -25333
rect 18077 -24157 18111 -24141
rect 18077 -25349 18111 -25333
rect 18535 -24157 18569 -24141
rect 18535 -25349 18569 -25333
rect 18993 -24157 19027 -24141
rect 18993 -25349 19027 -25333
rect 19451 -24157 19485 -24141
rect 19451 -25349 19485 -25333
rect 19909 -24157 19943 -24141
rect 19909 -25349 19943 -25333
rect 20367 -24157 20401 -24141
rect 20367 -25349 20401 -25333
rect 20825 -24157 20859 -24141
rect 20825 -25349 20859 -25333
rect 11365 -25426 11381 -25392
rect 11601 -25426 11617 -25392
rect 11823 -25426 11839 -25392
rect 12059 -25426 12075 -25392
rect 12281 -25426 12297 -25392
rect 12517 -25426 12533 -25392
rect 12739 -25426 12755 -25392
rect 12975 -25426 12991 -25392
rect 13197 -25426 13213 -25392
rect 13433 -25426 13449 -25392
rect 13655 -25426 13671 -25392
rect 13891 -25426 13907 -25392
rect 14113 -25426 14129 -25392
rect 14349 -25426 14365 -25392
rect 14571 -25426 14587 -25392
rect 14807 -25426 14823 -25392
rect 15029 -25426 15045 -25392
rect 15265 -25426 15281 -25392
rect 15487 -25426 15503 -25392
rect 15723 -25426 15739 -25392
rect 16365 -25426 16381 -25392
rect 16601 -25426 16617 -25392
rect 16823 -25426 16839 -25392
rect 17059 -25426 17075 -25392
rect 17281 -25426 17297 -25392
rect 17517 -25426 17533 -25392
rect 17739 -25426 17755 -25392
rect 17975 -25426 17991 -25392
rect 18197 -25426 18213 -25392
rect 18433 -25426 18449 -25392
rect 18655 -25426 18671 -25392
rect 18891 -25426 18907 -25392
rect 19113 -25426 19129 -25392
rect 19349 -25426 19365 -25392
rect 19571 -25426 19587 -25392
rect 19807 -25426 19823 -25392
rect 20029 -25426 20045 -25392
rect 20265 -25426 20281 -25392
rect 20487 -25426 20503 -25392
rect 20723 -25426 20739 -25392
rect 10818 -25872 10918 -25710
rect 21162 -25872 21262 -25710
rect 25818 -20190 25918 -20028
rect 36162 -20190 36262 -20028
rect 26924 -21433 26940 -21399
rect 27160 -21433 27176 -21399
rect 27382 -21433 27398 -21399
rect 27618 -21433 27634 -21399
rect 27840 -21433 27856 -21399
rect 28076 -21433 28092 -21399
rect 28298 -21433 28314 -21399
rect 28534 -21433 28550 -21399
rect 28756 -21433 28772 -21399
rect 28992 -21433 29008 -21399
rect 29214 -21433 29230 -21399
rect 29450 -21433 29466 -21399
rect 29672 -21433 29688 -21399
rect 29908 -21433 29924 -21399
rect 30130 -21433 30146 -21399
rect 30366 -21433 30382 -21399
rect 30588 -21433 30604 -21399
rect 30824 -21433 30840 -21399
rect 31046 -21433 31062 -21399
rect 31282 -21433 31298 -21399
rect 31504 -21433 31520 -21399
rect 31740 -21433 31756 -21399
rect 31962 -21433 31978 -21399
rect 32198 -21433 32214 -21399
rect 32420 -21433 32436 -21399
rect 32656 -21433 32672 -21399
rect 32878 -21433 32894 -21399
rect 33114 -21433 33130 -21399
rect 33336 -21433 33352 -21399
rect 33572 -21433 33588 -21399
rect 33794 -21433 33810 -21399
rect 34030 -21433 34046 -21399
rect 34252 -21433 34268 -21399
rect 34488 -21433 34504 -21399
rect 34710 -21433 34726 -21399
rect 34946 -21433 34962 -21399
rect 26804 -21492 26838 -21476
rect 26804 -23084 26838 -23068
rect 27262 -21492 27296 -21476
rect 27262 -23084 27296 -23068
rect 27720 -21492 27754 -21476
rect 27720 -23084 27754 -23068
rect 28178 -21492 28212 -21476
rect 28178 -23084 28212 -23068
rect 28636 -21492 28670 -21476
rect 28636 -23084 28670 -23068
rect 29094 -21492 29128 -21476
rect 29094 -23084 29128 -23068
rect 29552 -21492 29586 -21476
rect 29552 -23084 29586 -23068
rect 30010 -21492 30044 -21476
rect 30010 -23084 30044 -23068
rect 30468 -21492 30502 -21476
rect 30468 -23084 30502 -23068
rect 30926 -21492 30960 -21476
rect 30926 -23084 30960 -23068
rect 31384 -21492 31418 -21476
rect 31384 -23084 31418 -23068
rect 31842 -21492 31876 -21476
rect 31842 -23084 31876 -23068
rect 32300 -21492 32334 -21476
rect 32300 -23084 32334 -23068
rect 32758 -21492 32792 -21476
rect 32758 -23084 32792 -23068
rect 33216 -21492 33250 -21476
rect 33216 -23084 33250 -23068
rect 33674 -21492 33708 -21476
rect 33674 -23084 33708 -23068
rect 34132 -21492 34166 -21476
rect 34132 -23084 34166 -23068
rect 34590 -21492 34624 -21476
rect 34590 -23084 34624 -23068
rect 35048 -21492 35082 -21476
rect 35048 -23084 35082 -23068
rect 26924 -23161 26940 -23127
rect 27160 -23161 27176 -23127
rect 27382 -23161 27398 -23127
rect 27618 -23161 27634 -23127
rect 27840 -23161 27856 -23127
rect 28076 -23161 28092 -23127
rect 28298 -23161 28314 -23127
rect 28534 -23161 28550 -23127
rect 28756 -23161 28772 -23127
rect 28992 -23161 29008 -23127
rect 29214 -23161 29230 -23127
rect 29450 -23161 29466 -23127
rect 29672 -23161 29688 -23127
rect 29908 -23161 29924 -23127
rect 30130 -23161 30146 -23127
rect 30366 -23161 30382 -23127
rect 30588 -23161 30604 -23127
rect 30824 -23161 30840 -23127
rect 31046 -23161 31062 -23127
rect 31282 -23161 31298 -23127
rect 31504 -23161 31520 -23127
rect 31740 -23161 31756 -23127
rect 31962 -23161 31978 -23127
rect 32198 -23161 32214 -23127
rect 32420 -23161 32436 -23127
rect 32656 -23161 32672 -23127
rect 32878 -23161 32894 -23127
rect 33114 -23161 33130 -23127
rect 33336 -23161 33352 -23127
rect 33572 -23161 33588 -23127
rect 33794 -23161 33810 -23127
rect 34030 -23161 34046 -23127
rect 34252 -23161 34268 -23127
rect 34488 -23161 34504 -23127
rect 34710 -23161 34726 -23127
rect 34946 -23161 34962 -23127
rect 30682 -23244 31142 -23238
rect 30682 -23292 30688 -23244
rect 30736 -23292 31142 -23244
rect 30682 -23298 31142 -23292
rect 26365 -24098 26381 -24064
rect 26601 -24098 26617 -24064
rect 26823 -24098 26839 -24064
rect 27059 -24098 27075 -24064
rect 27281 -24098 27297 -24064
rect 27517 -24098 27533 -24064
rect 27739 -24098 27755 -24064
rect 27975 -24098 27991 -24064
rect 28197 -24098 28213 -24064
rect 28433 -24098 28449 -24064
rect 28655 -24098 28671 -24064
rect 28891 -24098 28907 -24064
rect 29113 -24098 29129 -24064
rect 29349 -24098 29365 -24064
rect 29571 -24098 29587 -24064
rect 29807 -24098 29823 -24064
rect 30029 -24098 30045 -24064
rect 30265 -24098 30281 -24064
rect 30487 -24098 30503 -24064
rect 30723 -24098 30739 -24064
rect 31365 -24098 31381 -24064
rect 31601 -24098 31617 -24064
rect 31823 -24098 31839 -24064
rect 32059 -24098 32075 -24064
rect 32281 -24098 32297 -24064
rect 32517 -24098 32533 -24064
rect 32739 -24098 32755 -24064
rect 32975 -24098 32991 -24064
rect 33197 -24098 33213 -24064
rect 33433 -24098 33449 -24064
rect 33655 -24098 33671 -24064
rect 33891 -24098 33907 -24064
rect 34113 -24098 34129 -24064
rect 34349 -24098 34365 -24064
rect 34571 -24098 34587 -24064
rect 34807 -24098 34823 -24064
rect 35029 -24098 35045 -24064
rect 35265 -24098 35281 -24064
rect 35487 -24098 35503 -24064
rect 35723 -24098 35739 -24064
rect 26245 -24157 26279 -24141
rect 26245 -25349 26279 -25333
rect 26703 -24157 26737 -24141
rect 26703 -25349 26737 -25333
rect 27161 -24157 27195 -24141
rect 27161 -25349 27195 -25333
rect 27619 -24157 27653 -24141
rect 27619 -25349 27653 -25333
rect 28077 -24157 28111 -24141
rect 28077 -25349 28111 -25333
rect 28535 -24157 28569 -24141
rect 28535 -25349 28569 -25333
rect 28993 -24157 29027 -24141
rect 28993 -25349 29027 -25333
rect 29451 -24157 29485 -24141
rect 29451 -25349 29485 -25333
rect 29909 -24157 29943 -24141
rect 29909 -25349 29943 -25333
rect 30367 -24157 30401 -24141
rect 30367 -25349 30401 -25333
rect 30825 -24157 30859 -24141
rect 30825 -25349 30859 -25333
rect 31245 -24157 31279 -24141
rect 31245 -25349 31279 -25333
rect 31703 -24157 31737 -24141
rect 31703 -25349 31737 -25333
rect 32161 -24157 32195 -24141
rect 32161 -25349 32195 -25333
rect 32619 -24157 32653 -24141
rect 32619 -25349 32653 -25333
rect 33077 -24157 33111 -24141
rect 33077 -25349 33111 -25333
rect 33535 -24157 33569 -24141
rect 33535 -25349 33569 -25333
rect 33993 -24157 34027 -24141
rect 33993 -25349 34027 -25333
rect 34451 -24157 34485 -24141
rect 34451 -25349 34485 -25333
rect 34909 -24157 34943 -24141
rect 34909 -25349 34943 -25333
rect 35367 -24157 35401 -24141
rect 35367 -25349 35401 -25333
rect 35825 -24157 35859 -24141
rect 35825 -25349 35859 -25333
rect 26365 -25426 26381 -25392
rect 26601 -25426 26617 -25392
rect 26823 -25426 26839 -25392
rect 27059 -25426 27075 -25392
rect 27281 -25426 27297 -25392
rect 27517 -25426 27533 -25392
rect 27739 -25426 27755 -25392
rect 27975 -25426 27991 -25392
rect 28197 -25426 28213 -25392
rect 28433 -25426 28449 -25392
rect 28655 -25426 28671 -25392
rect 28891 -25426 28907 -25392
rect 29113 -25426 29129 -25392
rect 29349 -25426 29365 -25392
rect 29571 -25426 29587 -25392
rect 29807 -25426 29823 -25392
rect 30029 -25426 30045 -25392
rect 30265 -25426 30281 -25392
rect 30487 -25426 30503 -25392
rect 30723 -25426 30739 -25392
rect 31365 -25426 31381 -25392
rect 31601 -25426 31617 -25392
rect 31823 -25426 31839 -25392
rect 32059 -25426 32075 -25392
rect 32281 -25426 32297 -25392
rect 32517 -25426 32533 -25392
rect 32739 -25426 32755 -25392
rect 32975 -25426 32991 -25392
rect 33197 -25426 33213 -25392
rect 33433 -25426 33449 -25392
rect 33655 -25426 33671 -25392
rect 33891 -25426 33907 -25392
rect 34113 -25426 34129 -25392
rect 34349 -25426 34365 -25392
rect 34571 -25426 34587 -25392
rect 34807 -25426 34823 -25392
rect 35029 -25426 35045 -25392
rect 35265 -25426 35281 -25392
rect 35487 -25426 35503 -25392
rect 35723 -25426 35739 -25392
rect 25818 -25872 25918 -25710
rect 36162 -25872 36262 -25710
rect 10818 -26270 10918 -26108
rect 21162 -26270 21262 -26108
rect 11364 -26600 11380 -26566
rect 11600 -26600 11616 -26566
rect 11822 -26600 11838 -26566
rect 12058 -26600 12074 -26566
rect 12280 -26600 12296 -26566
rect 12516 -26600 12532 -26566
rect 12738 -26600 12754 -26566
rect 12974 -26600 12990 -26566
rect 13196 -26600 13212 -26566
rect 13432 -26600 13448 -26566
rect 13654 -26600 13670 -26566
rect 13890 -26600 13906 -26566
rect 14112 -26600 14128 -26566
rect 14348 -26600 14364 -26566
rect 14570 -26600 14586 -26566
rect 14806 -26600 14822 -26566
rect 15028 -26600 15044 -26566
rect 15264 -26600 15280 -26566
rect 15486 -26600 15502 -26566
rect 15722 -26600 15738 -26566
rect 16364 -26600 16380 -26566
rect 16600 -26600 16616 -26566
rect 16822 -26600 16838 -26566
rect 17058 -26600 17074 -26566
rect 17280 -26600 17296 -26566
rect 17516 -26600 17532 -26566
rect 17738 -26600 17754 -26566
rect 17974 -26600 17990 -26566
rect 18196 -26600 18212 -26566
rect 18432 -26600 18448 -26566
rect 18654 -26600 18670 -26566
rect 18890 -26600 18906 -26566
rect 19112 -26600 19128 -26566
rect 19348 -26600 19364 -26566
rect 19570 -26600 19586 -26566
rect 19806 -26600 19822 -26566
rect 20028 -26600 20044 -26566
rect 20264 -26600 20280 -26566
rect 20486 -26600 20502 -26566
rect 20722 -26600 20738 -26566
rect 11244 -26650 11278 -26634
rect 11244 -26842 11278 -26826
rect 11702 -26650 11736 -26634
rect 11702 -26842 11736 -26826
rect 12160 -26650 12194 -26634
rect 12160 -26842 12194 -26826
rect 12618 -26650 12652 -26634
rect 12618 -26842 12652 -26826
rect 13076 -26650 13110 -26634
rect 13076 -26842 13110 -26826
rect 13534 -26650 13568 -26634
rect 13534 -26842 13568 -26826
rect 13992 -26650 14026 -26634
rect 13992 -26842 14026 -26826
rect 14450 -26650 14484 -26634
rect 14450 -26842 14484 -26826
rect 14908 -26650 14942 -26634
rect 14908 -26842 14942 -26826
rect 15366 -26650 15400 -26634
rect 15366 -26842 15400 -26826
rect 15824 -26650 15858 -26634
rect 15824 -26842 15858 -26826
rect 16244 -26650 16278 -26634
rect 16244 -26842 16278 -26826
rect 16702 -26650 16736 -26634
rect 16702 -26842 16736 -26826
rect 17160 -26650 17194 -26634
rect 17160 -26842 17194 -26826
rect 17618 -26650 17652 -26634
rect 17618 -26842 17652 -26826
rect 18076 -26650 18110 -26634
rect 18076 -26842 18110 -26826
rect 18534 -26650 18568 -26634
rect 18534 -26842 18568 -26826
rect 18992 -26650 19026 -26634
rect 18992 -26842 19026 -26826
rect 19450 -26650 19484 -26634
rect 19450 -26842 19484 -26826
rect 19908 -26650 19942 -26634
rect 19908 -26842 19942 -26826
rect 20366 -26650 20400 -26634
rect 20366 -26842 20400 -26826
rect 20824 -26650 20858 -26634
rect 20824 -26842 20858 -26826
rect 11364 -26910 11380 -26876
rect 11600 -26910 11616 -26876
rect 11822 -26910 11838 -26876
rect 12058 -26910 12074 -26876
rect 12280 -26910 12296 -26876
rect 12516 -26910 12532 -26876
rect 12738 -26910 12754 -26876
rect 12974 -26910 12990 -26876
rect 13196 -26910 13212 -26876
rect 13432 -26910 13448 -26876
rect 13654 -26910 13670 -26876
rect 13890 -26910 13906 -26876
rect 14112 -26910 14128 -26876
rect 14348 -26910 14364 -26876
rect 14570 -26910 14586 -26876
rect 14806 -26910 14822 -26876
rect 15028 -26910 15044 -26876
rect 15264 -26910 15280 -26876
rect 15486 -26910 15502 -26876
rect 15722 -26910 15738 -26876
rect 16364 -26910 16380 -26876
rect 16600 -26910 16616 -26876
rect 16822 -26910 16838 -26876
rect 17058 -26910 17074 -26876
rect 17280 -26910 17296 -26876
rect 17516 -26910 17532 -26876
rect 17738 -26910 17754 -26876
rect 17974 -26910 17990 -26876
rect 18196 -26910 18212 -26876
rect 18432 -26910 18448 -26876
rect 18654 -26910 18670 -26876
rect 18890 -26910 18906 -26876
rect 19112 -26910 19128 -26876
rect 19348 -26910 19364 -26876
rect 19570 -26910 19586 -26876
rect 19806 -26910 19822 -26876
rect 20028 -26910 20044 -26876
rect 20264 -26910 20280 -26876
rect 20486 -26910 20502 -26876
rect 20722 -26910 20738 -26876
rect 11364 -27268 11380 -27234
rect 11600 -27268 11616 -27234
rect 11822 -27268 11838 -27234
rect 12058 -27268 12074 -27234
rect 12280 -27268 12296 -27234
rect 12516 -27268 12532 -27234
rect 12738 -27268 12754 -27234
rect 12974 -27268 12990 -27234
rect 13196 -27268 13212 -27234
rect 13432 -27268 13448 -27234
rect 13654 -27268 13670 -27234
rect 13890 -27268 13906 -27234
rect 14112 -27268 14128 -27234
rect 14348 -27268 14364 -27234
rect 14570 -27268 14586 -27234
rect 14806 -27268 14822 -27234
rect 15028 -27268 15044 -27234
rect 15264 -27268 15280 -27234
rect 15486 -27268 15502 -27234
rect 15722 -27268 15738 -27234
rect 11244 -27318 11278 -27302
rect 11244 -27510 11278 -27494
rect 11702 -27318 11736 -27302
rect 11702 -27510 11736 -27494
rect 12160 -27318 12194 -27302
rect 12160 -27510 12194 -27494
rect 12618 -27318 12652 -27302
rect 12618 -27510 12652 -27494
rect 13076 -27318 13110 -27302
rect 13076 -27510 13110 -27494
rect 13534 -27318 13568 -27302
rect 13534 -27510 13568 -27494
rect 13992 -27318 14026 -27302
rect 13992 -27510 14026 -27494
rect 14450 -27318 14484 -27302
rect 14450 -27510 14484 -27494
rect 14908 -27318 14942 -27302
rect 14908 -27510 14942 -27494
rect 15366 -27318 15400 -27302
rect 15366 -27510 15400 -27494
rect 15824 -27318 15858 -27302
rect 15824 -27510 15858 -27494
rect 11364 -27578 11380 -27544
rect 11600 -27578 11616 -27544
rect 11822 -27578 11838 -27544
rect 12058 -27578 12074 -27544
rect 12280 -27578 12296 -27544
rect 12516 -27578 12532 -27544
rect 12738 -27578 12754 -27544
rect 12974 -27578 12990 -27544
rect 13196 -27578 13212 -27544
rect 13432 -27578 13448 -27544
rect 13654 -27578 13670 -27544
rect 13890 -27578 13906 -27544
rect 14112 -27578 14128 -27544
rect 14348 -27578 14364 -27544
rect 14570 -27578 14586 -27544
rect 14806 -27578 14822 -27544
rect 15028 -27578 15044 -27544
rect 15264 -27578 15280 -27544
rect 15486 -27578 15502 -27544
rect 15722 -27578 15738 -27544
rect 10818 -28572 10918 -28410
rect 21162 -28572 21262 -28410
rect 25818 -26270 25918 -26108
rect 36162 -26270 36262 -26108
rect 26364 -26600 26380 -26566
rect 26600 -26600 26616 -26566
rect 26822 -26600 26838 -26566
rect 27058 -26600 27074 -26566
rect 27280 -26600 27296 -26566
rect 27516 -26600 27532 -26566
rect 27738 -26600 27754 -26566
rect 27974 -26600 27990 -26566
rect 28196 -26600 28212 -26566
rect 28432 -26600 28448 -26566
rect 28654 -26600 28670 -26566
rect 28890 -26600 28906 -26566
rect 29112 -26600 29128 -26566
rect 29348 -26600 29364 -26566
rect 29570 -26600 29586 -26566
rect 29806 -26600 29822 -26566
rect 30028 -26600 30044 -26566
rect 30264 -26600 30280 -26566
rect 30486 -26600 30502 -26566
rect 30722 -26600 30738 -26566
rect 31364 -26600 31380 -26566
rect 31600 -26600 31616 -26566
rect 31822 -26600 31838 -26566
rect 32058 -26600 32074 -26566
rect 32280 -26600 32296 -26566
rect 32516 -26600 32532 -26566
rect 32738 -26600 32754 -26566
rect 32974 -26600 32990 -26566
rect 33196 -26600 33212 -26566
rect 33432 -26600 33448 -26566
rect 33654 -26600 33670 -26566
rect 33890 -26600 33906 -26566
rect 34112 -26600 34128 -26566
rect 34348 -26600 34364 -26566
rect 34570 -26600 34586 -26566
rect 34806 -26600 34822 -26566
rect 35028 -26600 35044 -26566
rect 35264 -26600 35280 -26566
rect 35486 -26600 35502 -26566
rect 35722 -26600 35738 -26566
rect 26244 -26650 26278 -26634
rect 26244 -26842 26278 -26826
rect 26702 -26650 26736 -26634
rect 26702 -26842 26736 -26826
rect 27160 -26650 27194 -26634
rect 27160 -26842 27194 -26826
rect 27618 -26650 27652 -26634
rect 27618 -26842 27652 -26826
rect 28076 -26650 28110 -26634
rect 28076 -26842 28110 -26826
rect 28534 -26650 28568 -26634
rect 28534 -26842 28568 -26826
rect 28992 -26650 29026 -26634
rect 28992 -26842 29026 -26826
rect 29450 -26650 29484 -26634
rect 29450 -26842 29484 -26826
rect 29908 -26650 29942 -26634
rect 29908 -26842 29942 -26826
rect 30366 -26650 30400 -26634
rect 30366 -26842 30400 -26826
rect 30824 -26650 30858 -26634
rect 30824 -26842 30858 -26826
rect 31244 -26650 31278 -26634
rect 31244 -26842 31278 -26826
rect 31702 -26650 31736 -26634
rect 31702 -26842 31736 -26826
rect 32160 -26650 32194 -26634
rect 32160 -26842 32194 -26826
rect 32618 -26650 32652 -26634
rect 32618 -26842 32652 -26826
rect 33076 -26650 33110 -26634
rect 33076 -26842 33110 -26826
rect 33534 -26650 33568 -26634
rect 33534 -26842 33568 -26826
rect 33992 -26650 34026 -26634
rect 33992 -26842 34026 -26826
rect 34450 -26650 34484 -26634
rect 34450 -26842 34484 -26826
rect 34908 -26650 34942 -26634
rect 34908 -26842 34942 -26826
rect 35366 -26650 35400 -26634
rect 35366 -26842 35400 -26826
rect 35824 -26650 35858 -26634
rect 35824 -26842 35858 -26826
rect 26364 -26910 26380 -26876
rect 26600 -26910 26616 -26876
rect 26822 -26910 26838 -26876
rect 27058 -26910 27074 -26876
rect 27280 -26910 27296 -26876
rect 27516 -26910 27532 -26876
rect 27738 -26910 27754 -26876
rect 27974 -26910 27990 -26876
rect 28196 -26910 28212 -26876
rect 28432 -26910 28448 -26876
rect 28654 -26910 28670 -26876
rect 28890 -26910 28906 -26876
rect 29112 -26910 29128 -26876
rect 29348 -26910 29364 -26876
rect 29570 -26910 29586 -26876
rect 29806 -26910 29822 -26876
rect 30028 -26910 30044 -26876
rect 30264 -26910 30280 -26876
rect 30486 -26910 30502 -26876
rect 30722 -26910 30738 -26876
rect 31364 -26910 31380 -26876
rect 31600 -26910 31616 -26876
rect 31822 -26910 31838 -26876
rect 32058 -26910 32074 -26876
rect 32280 -26910 32296 -26876
rect 32516 -26910 32532 -26876
rect 32738 -26910 32754 -26876
rect 32974 -26910 32990 -26876
rect 33196 -26910 33212 -26876
rect 33432 -26910 33448 -26876
rect 33654 -26910 33670 -26876
rect 33890 -26910 33906 -26876
rect 34112 -26910 34128 -26876
rect 34348 -26910 34364 -26876
rect 34570 -26910 34586 -26876
rect 34806 -26910 34822 -26876
rect 35028 -26910 35044 -26876
rect 35264 -26910 35280 -26876
rect 35486 -26910 35502 -26876
rect 35722 -26910 35738 -26876
rect 26364 -27268 26380 -27234
rect 26600 -27268 26616 -27234
rect 26822 -27268 26838 -27234
rect 27058 -27268 27074 -27234
rect 27280 -27268 27296 -27234
rect 27516 -27268 27532 -27234
rect 27738 -27268 27754 -27234
rect 27974 -27268 27990 -27234
rect 28196 -27268 28212 -27234
rect 28432 -27268 28448 -27234
rect 28654 -27268 28670 -27234
rect 28890 -27268 28906 -27234
rect 29112 -27268 29128 -27234
rect 29348 -27268 29364 -27234
rect 29570 -27268 29586 -27234
rect 29806 -27268 29822 -27234
rect 30028 -27268 30044 -27234
rect 30264 -27268 30280 -27234
rect 30486 -27268 30502 -27234
rect 30722 -27268 30738 -27234
rect 26244 -27318 26278 -27302
rect 26244 -27510 26278 -27494
rect 26702 -27318 26736 -27302
rect 26702 -27510 26736 -27494
rect 27160 -27318 27194 -27302
rect 27160 -27510 27194 -27494
rect 27618 -27318 27652 -27302
rect 27618 -27510 27652 -27494
rect 28076 -27318 28110 -27302
rect 28076 -27510 28110 -27494
rect 28534 -27318 28568 -27302
rect 28534 -27510 28568 -27494
rect 28992 -27318 29026 -27302
rect 28992 -27510 29026 -27494
rect 29450 -27318 29484 -27302
rect 29450 -27510 29484 -27494
rect 29908 -27318 29942 -27302
rect 29908 -27510 29942 -27494
rect 30366 -27318 30400 -27302
rect 30366 -27510 30400 -27494
rect 30824 -27318 30858 -27302
rect 30824 -27510 30858 -27494
rect 26364 -27578 26380 -27544
rect 26600 -27578 26616 -27544
rect 26822 -27578 26838 -27544
rect 27058 -27578 27074 -27544
rect 27280 -27578 27296 -27544
rect 27516 -27578 27532 -27544
rect 27738 -27578 27754 -27544
rect 27974 -27578 27990 -27544
rect 28196 -27578 28212 -27544
rect 28432 -27578 28448 -27544
rect 28654 -27578 28670 -27544
rect 28890 -27578 28906 -27544
rect 29112 -27578 29128 -27544
rect 29348 -27578 29364 -27544
rect 29570 -27578 29586 -27544
rect 29806 -27578 29822 -27544
rect 30028 -27578 30044 -27544
rect 30264 -27578 30280 -27544
rect 30486 -27578 30502 -27544
rect 30722 -27578 30738 -27544
rect 25818 -28572 25918 -28410
rect 36162 -28572 36262 -28410
<< viali >>
rect 15526 4210 15588 4310
rect 15588 4210 24288 4310
rect 24288 4210 24350 4310
rect 15426 2698 15526 4122
rect 17788 3282 17972 3316
rect 18246 3282 18430 3316
rect 18704 3282 18888 3316
rect 19162 3282 19346 3316
rect 19620 3282 19804 3316
rect 20078 3282 20262 3316
rect 20536 3282 20720 3316
rect 20994 3282 21178 3316
rect 21452 3282 21636 3316
rect 21910 3282 22094 3316
rect 17634 3056 17668 3232
rect 18092 3056 18126 3232
rect 18550 3056 18584 3232
rect 19008 3056 19042 3232
rect 19466 3056 19500 3232
rect 19924 3056 19958 3232
rect 20382 3056 20416 3232
rect 20840 3056 20874 3232
rect 21298 3056 21332 3232
rect 21756 3056 21790 3232
rect 22214 3056 22248 3232
rect 17788 2972 17972 3006
rect 18246 2972 18430 3006
rect 18704 2972 18888 3006
rect 19162 2972 19346 3006
rect 19620 2972 19804 3006
rect 20078 2972 20262 3006
rect 20536 2972 20720 3006
rect 20994 2972 21178 3006
rect 21452 2972 21636 3006
rect 21910 2972 22094 3006
rect 24350 2698 24450 4122
rect 15526 2510 15588 2610
rect 15588 2510 24288 2610
rect 24288 2510 24350 2610
rect 26108 4210 26170 4310
rect 26170 4210 31290 4310
rect 31290 4210 31352 4310
rect 26008 2614 26108 4126
rect 26550 3282 26734 3316
rect 27008 3282 27192 3316
rect 27466 3282 27650 3316
rect 27924 3282 28108 3316
rect 28382 3282 28566 3316
rect 28840 3282 29024 3316
rect 29298 3282 29482 3316
rect 29756 3282 29940 3316
rect 30214 3282 30398 3316
rect 30672 3282 30856 3316
rect 26396 3056 26430 3232
rect 26854 3056 26888 3232
rect 27312 3056 27346 3232
rect 27770 3056 27804 3232
rect 28228 3056 28262 3232
rect 28686 3056 28720 3232
rect 29144 3056 29178 3232
rect 29602 3056 29636 3232
rect 30060 3056 30094 3232
rect 30518 3056 30552 3232
rect 30976 3056 31010 3232
rect 26550 2972 26734 3006
rect 27008 2972 27192 3006
rect 27466 2972 27650 3006
rect 27924 2972 28108 3006
rect 28382 2972 28566 3006
rect 28840 2972 29024 3006
rect 29298 2972 29482 3006
rect 29756 2972 29940 3006
rect 30214 2972 30398 3006
rect 30672 2972 30856 3006
rect 31352 2614 31452 4126
rect 26108 2430 26170 2530
rect 26170 2430 31290 2530
rect 31290 2430 31352 2530
rect 31571 2473 31605 2507
rect 31663 2473 31697 2507
rect 31755 2473 31789 2507
rect 31847 2473 31881 2507
rect 31939 2473 31973 2507
rect 32031 2473 32065 2507
rect 32123 2473 32157 2507
rect 32215 2473 32249 2507
rect 15526 2174 15588 2274
rect 15588 2174 24288 2274
rect 24288 2174 24350 2274
rect 15426 -1360 15526 1976
rect 31606 2241 31622 2274
rect 31622 2241 31654 2274
rect 31606 2226 31654 2241
rect 31712 2228 31760 2276
rect 31848 2275 31896 2276
rect 31848 2241 31855 2275
rect 31855 2241 31889 2275
rect 31889 2241 31896 2275
rect 31848 2228 31896 2241
rect 15956 1440 16140 1474
rect 16414 1440 16598 1474
rect 16872 1440 17056 1474
rect 17330 1440 17514 1474
rect 17788 1440 17972 1474
rect 18246 1440 18430 1474
rect 18704 1440 18888 1474
rect 19162 1440 19346 1474
rect 19620 1440 19804 1474
rect 20078 1440 20262 1474
rect 20536 1440 20720 1474
rect 20994 1440 21178 1474
rect 21452 1440 21636 1474
rect 21910 1440 22094 1474
rect 22368 1440 22552 1474
rect 22826 1440 23010 1474
rect 23284 1440 23468 1474
rect 23742 1440 23926 1474
rect 15802 -195 15836 1381
rect 16260 -195 16294 1381
rect 16718 -195 16752 1381
rect 17176 -195 17210 1381
rect 17634 -195 17668 1381
rect 18092 -195 18126 1381
rect 18550 -195 18584 1381
rect 19008 -195 19042 1381
rect 19466 -195 19500 1381
rect 19924 -195 19958 1381
rect 20382 -195 20416 1381
rect 20840 -195 20874 1381
rect 21298 -195 21332 1381
rect 21756 -195 21790 1381
rect 22214 -195 22248 1381
rect 22672 -195 22706 1381
rect 23130 -195 23164 1381
rect 23588 -195 23622 1381
rect 24046 -195 24080 1381
rect 15956 -288 16140 -254
rect 16414 -288 16598 -254
rect 16872 -288 17056 -254
rect 17330 -288 17514 -254
rect 17788 -288 17972 -254
rect 18246 -288 18430 -254
rect 18704 -288 18888 -254
rect 19162 -288 19346 -254
rect 19620 -288 19804 -254
rect 20078 -288 20262 -254
rect 20536 -288 20720 -254
rect 20994 -288 21178 -254
rect 21452 -288 21636 -254
rect 21910 -288 22094 -254
rect 22368 -288 22552 -254
rect 22826 -288 23010 -254
rect 23284 -288 23468 -254
rect 23742 -288 23926 -254
rect 24350 -1360 24450 1976
rect 15526 -1658 15588 -1558
rect 15588 -1658 24288 -1558
rect 24288 -1658 24350 -1558
rect 26108 2094 26170 2194
rect 26170 2094 31290 2194
rect 31290 2094 31352 2194
rect 26008 -1375 26108 1911
rect 32204 2228 32252 2276
rect 31571 1929 31605 1963
rect 31663 1929 31697 1963
rect 31755 1929 31789 1963
rect 31847 1929 31881 1963
rect 31939 1929 31973 1963
rect 32031 1929 32065 1963
rect 32123 1929 32157 1963
rect 32215 1929 32249 1963
rect 26551 1860 26735 1894
rect 27009 1860 27193 1894
rect 27467 1860 27651 1894
rect 27925 1860 28109 1894
rect 28383 1860 28567 1894
rect 28841 1860 29025 1894
rect 29299 1860 29483 1894
rect 29757 1860 29941 1894
rect 30215 1860 30399 1894
rect 30673 1860 30857 1894
rect 26397 625 26431 1801
rect 26855 625 26889 1801
rect 27313 625 27347 1801
rect 27771 625 27805 1801
rect 28229 625 28263 1801
rect 28687 625 28721 1801
rect 29145 625 29179 1801
rect 29603 625 29637 1801
rect 30061 625 30095 1801
rect 30519 625 30553 1801
rect 30977 625 31011 1801
rect 26551 532 26735 566
rect 27009 532 27193 566
rect 27467 532 27651 566
rect 27925 532 28109 566
rect 28383 532 28567 566
rect 28841 532 29025 566
rect 29299 532 29483 566
rect 29757 532 29941 566
rect 30215 532 30399 566
rect 30673 532 30857 566
rect 31352 -1375 31452 1911
rect 26108 -1658 26170 -1558
rect 26170 -1658 31290 -1558
rect 31290 -1658 31352 -1558
rect 10918 -2128 10980 -2028
rect 10980 -2128 21100 -2028
rect 21100 -2128 21162 -2028
rect 10818 -7590 10918 -2418
rect 11958 -3433 12142 -3399
rect 12416 -3433 12600 -3399
rect 12874 -3433 13058 -3399
rect 13332 -3433 13516 -3399
rect 13790 -3433 13974 -3399
rect 14248 -3433 14432 -3399
rect 14706 -3433 14890 -3399
rect 15164 -3433 15348 -3399
rect 15622 -3433 15806 -3399
rect 16080 -3433 16264 -3399
rect 16538 -3433 16722 -3399
rect 16996 -3433 17180 -3399
rect 17454 -3433 17638 -3399
rect 17912 -3433 18096 -3399
rect 18370 -3433 18554 -3399
rect 18828 -3433 19012 -3399
rect 19286 -3433 19470 -3399
rect 19744 -3433 19928 -3399
rect 11804 -5068 11838 -3492
rect 12262 -5068 12296 -3492
rect 12720 -5068 12754 -3492
rect 13178 -5068 13212 -3492
rect 13636 -5068 13670 -3492
rect 14094 -5068 14128 -3492
rect 14552 -5068 14586 -3492
rect 15010 -5068 15044 -3492
rect 15468 -5068 15502 -3492
rect 15926 -5068 15960 -3492
rect 16384 -5068 16418 -3492
rect 16842 -5068 16876 -3492
rect 17300 -5068 17334 -3492
rect 17758 -5068 17792 -3492
rect 18216 -5068 18250 -3492
rect 18674 -5068 18708 -3492
rect 19132 -5068 19166 -3492
rect 19590 -5068 19624 -3492
rect 20048 -5068 20082 -3492
rect 11958 -5161 12142 -5127
rect 12416 -5161 12600 -5127
rect 12874 -5161 13058 -5127
rect 13332 -5161 13516 -5127
rect 13790 -5161 13974 -5127
rect 14248 -5161 14432 -5127
rect 14706 -5161 14890 -5127
rect 15164 -5161 15348 -5127
rect 15622 -5161 15806 -5127
rect 16080 -5161 16264 -5127
rect 16538 -5161 16722 -5127
rect 16996 -5161 17180 -5127
rect 17454 -5161 17638 -5127
rect 17912 -5161 18096 -5127
rect 18370 -5161 18554 -5127
rect 18828 -5161 19012 -5127
rect 19286 -5161 19470 -5127
rect 19744 -5161 19928 -5127
rect 15688 -5292 15736 -5244
rect 16142 -5298 16202 -5238
rect 11399 -6098 11583 -6064
rect 11857 -6098 12041 -6064
rect 12315 -6098 12499 -6064
rect 12773 -6098 12957 -6064
rect 13231 -6098 13415 -6064
rect 13689 -6098 13873 -6064
rect 14147 -6098 14331 -6064
rect 14605 -6098 14789 -6064
rect 15063 -6098 15247 -6064
rect 15521 -6098 15705 -6064
rect 16399 -6098 16583 -6064
rect 16857 -6098 17041 -6064
rect 17315 -6098 17499 -6064
rect 17773 -6098 17957 -6064
rect 18231 -6098 18415 -6064
rect 18689 -6098 18873 -6064
rect 19147 -6098 19331 -6064
rect 19605 -6098 19789 -6064
rect 20063 -6098 20247 -6064
rect 20521 -6098 20705 -6064
rect 11245 -7333 11279 -6157
rect 11703 -7333 11737 -6157
rect 12161 -7333 12195 -6157
rect 12619 -7333 12653 -6157
rect 13077 -7333 13111 -6157
rect 13535 -7333 13569 -6157
rect 13993 -7333 14027 -6157
rect 14451 -7333 14485 -6157
rect 14909 -7333 14943 -6157
rect 15367 -7333 15401 -6157
rect 15825 -7333 15859 -6157
rect 16245 -7333 16279 -6157
rect 16703 -7333 16737 -6157
rect 17161 -7333 17195 -6157
rect 17619 -7333 17653 -6157
rect 18077 -7333 18111 -6157
rect 18535 -7333 18569 -6157
rect 18993 -7333 19027 -6157
rect 19451 -7333 19485 -6157
rect 19909 -7333 19943 -6157
rect 20367 -7333 20401 -6157
rect 20825 -7333 20859 -6157
rect 11399 -7426 11583 -7392
rect 11857 -7426 12041 -7392
rect 12315 -7426 12499 -7392
rect 12773 -7426 12957 -7392
rect 13231 -7426 13415 -7392
rect 13689 -7426 13873 -7392
rect 14147 -7426 14331 -7392
rect 14605 -7426 14789 -7392
rect 15063 -7426 15247 -7392
rect 15521 -7426 15705 -7392
rect 16399 -7426 16583 -7392
rect 16857 -7426 17041 -7392
rect 17315 -7426 17499 -7392
rect 17773 -7426 17957 -7392
rect 18231 -7426 18415 -7392
rect 18689 -7426 18873 -7392
rect 19147 -7426 19331 -7392
rect 19605 -7426 19789 -7392
rect 20063 -7426 20247 -7392
rect 20521 -7426 20705 -7392
rect 21162 -7590 21262 -2418
rect 10918 -7872 10980 -7772
rect 10980 -7872 21100 -7772
rect 21100 -7872 21162 -7772
rect 25918 -2128 25980 -2028
rect 25980 -2128 36100 -2028
rect 36100 -2128 36162 -2028
rect 25818 -7590 25918 -2418
rect 26958 -3433 27142 -3399
rect 27416 -3433 27600 -3399
rect 27874 -3433 28058 -3399
rect 28332 -3433 28516 -3399
rect 28790 -3433 28974 -3399
rect 29248 -3433 29432 -3399
rect 29706 -3433 29890 -3399
rect 30164 -3433 30348 -3399
rect 30622 -3433 30806 -3399
rect 31080 -3433 31264 -3399
rect 31538 -3433 31722 -3399
rect 31996 -3433 32180 -3399
rect 32454 -3433 32638 -3399
rect 32912 -3433 33096 -3399
rect 33370 -3433 33554 -3399
rect 33828 -3433 34012 -3399
rect 34286 -3433 34470 -3399
rect 34744 -3433 34928 -3399
rect 26804 -5068 26838 -3492
rect 27262 -5068 27296 -3492
rect 27720 -5068 27754 -3492
rect 28178 -5068 28212 -3492
rect 28636 -5068 28670 -3492
rect 29094 -5068 29128 -3492
rect 29552 -5068 29586 -3492
rect 30010 -5068 30044 -3492
rect 30468 -5068 30502 -3492
rect 30926 -5068 30960 -3492
rect 31384 -5068 31418 -3492
rect 31842 -5068 31876 -3492
rect 32300 -5068 32334 -3492
rect 32758 -5068 32792 -3492
rect 33216 -5068 33250 -3492
rect 33674 -5068 33708 -3492
rect 34132 -5068 34166 -3492
rect 34590 -5068 34624 -3492
rect 35048 -5068 35082 -3492
rect 26958 -5161 27142 -5127
rect 27416 -5161 27600 -5127
rect 27874 -5161 28058 -5127
rect 28332 -5161 28516 -5127
rect 28790 -5161 28974 -5127
rect 29248 -5161 29432 -5127
rect 29706 -5161 29890 -5127
rect 30164 -5161 30348 -5127
rect 30622 -5161 30806 -5127
rect 31080 -5161 31264 -5127
rect 31538 -5161 31722 -5127
rect 31996 -5161 32180 -5127
rect 32454 -5161 32638 -5127
rect 32912 -5161 33096 -5127
rect 33370 -5161 33554 -5127
rect 33828 -5161 34012 -5127
rect 34286 -5161 34470 -5127
rect 34744 -5161 34928 -5127
rect 30688 -5292 30736 -5244
rect 31142 -5298 31202 -5238
rect 26399 -6098 26583 -6064
rect 26857 -6098 27041 -6064
rect 27315 -6098 27499 -6064
rect 27773 -6098 27957 -6064
rect 28231 -6098 28415 -6064
rect 28689 -6098 28873 -6064
rect 29147 -6098 29331 -6064
rect 29605 -6098 29789 -6064
rect 30063 -6098 30247 -6064
rect 30521 -6098 30705 -6064
rect 31399 -6098 31583 -6064
rect 31857 -6098 32041 -6064
rect 32315 -6098 32499 -6064
rect 32773 -6098 32957 -6064
rect 33231 -6098 33415 -6064
rect 33689 -6098 33873 -6064
rect 34147 -6098 34331 -6064
rect 34605 -6098 34789 -6064
rect 35063 -6098 35247 -6064
rect 35521 -6098 35705 -6064
rect 26245 -7333 26279 -6157
rect 26703 -7333 26737 -6157
rect 27161 -7333 27195 -6157
rect 27619 -7333 27653 -6157
rect 28077 -7333 28111 -6157
rect 28535 -7333 28569 -6157
rect 28993 -7333 29027 -6157
rect 29451 -7333 29485 -6157
rect 29909 -7333 29943 -6157
rect 30367 -7333 30401 -6157
rect 30825 -7333 30859 -6157
rect 31245 -7333 31279 -6157
rect 31703 -7333 31737 -6157
rect 32161 -7333 32195 -6157
rect 32619 -7333 32653 -6157
rect 33077 -7333 33111 -6157
rect 33535 -7333 33569 -6157
rect 33993 -7333 34027 -6157
rect 34451 -7333 34485 -6157
rect 34909 -7333 34943 -6157
rect 35367 -7333 35401 -6157
rect 35825 -7333 35859 -6157
rect 26399 -7426 26583 -7392
rect 26857 -7426 27041 -7392
rect 27315 -7426 27499 -7392
rect 27773 -7426 27957 -7392
rect 28231 -7426 28415 -7392
rect 28689 -7426 28873 -7392
rect 29147 -7426 29331 -7392
rect 29605 -7426 29789 -7392
rect 30063 -7426 30247 -7392
rect 30521 -7426 30705 -7392
rect 31399 -7426 31583 -7392
rect 31857 -7426 32041 -7392
rect 32315 -7426 32499 -7392
rect 32773 -7426 32957 -7392
rect 33231 -7426 33415 -7392
rect 33689 -7426 33873 -7392
rect 34147 -7426 34331 -7392
rect 34605 -7426 34789 -7392
rect 35063 -7426 35247 -7392
rect 35521 -7426 35705 -7392
rect 36162 -7590 36262 -2418
rect 25918 -7872 25980 -7772
rect 25980 -7872 36100 -7772
rect 36100 -7872 36162 -7772
rect 10918 -8208 10980 -8108
rect 10980 -8208 21100 -8108
rect 21100 -8208 21162 -8108
rect 10818 -10342 10918 -8338
rect 11398 -8600 11582 -8566
rect 11856 -8600 12040 -8566
rect 12314 -8600 12498 -8566
rect 12772 -8600 12956 -8566
rect 13230 -8600 13414 -8566
rect 13688 -8600 13872 -8566
rect 14146 -8600 14330 -8566
rect 14604 -8600 14788 -8566
rect 15062 -8600 15246 -8566
rect 15520 -8600 15704 -8566
rect 16398 -8600 16582 -8566
rect 16856 -8600 17040 -8566
rect 17314 -8600 17498 -8566
rect 17772 -8600 17956 -8566
rect 18230 -8600 18414 -8566
rect 18688 -8600 18872 -8566
rect 19146 -8600 19330 -8566
rect 19604 -8600 19788 -8566
rect 20062 -8600 20246 -8566
rect 20520 -8600 20704 -8566
rect 11244 -8826 11278 -8650
rect 11702 -8826 11736 -8650
rect 12160 -8826 12194 -8650
rect 12618 -8826 12652 -8650
rect 13076 -8826 13110 -8650
rect 13534 -8826 13568 -8650
rect 13992 -8826 14026 -8650
rect 14450 -8826 14484 -8650
rect 14908 -8826 14942 -8650
rect 15366 -8826 15400 -8650
rect 15824 -8826 15858 -8650
rect 16244 -8826 16278 -8650
rect 16702 -8826 16736 -8650
rect 17160 -8826 17194 -8650
rect 17618 -8826 17652 -8650
rect 18076 -8826 18110 -8650
rect 18534 -8826 18568 -8650
rect 18992 -8826 19026 -8650
rect 19450 -8826 19484 -8650
rect 19908 -8826 19942 -8650
rect 20366 -8826 20400 -8650
rect 20824 -8826 20858 -8650
rect 11398 -8910 11582 -8876
rect 11856 -8910 12040 -8876
rect 12314 -8910 12498 -8876
rect 12772 -8910 12956 -8876
rect 13230 -8910 13414 -8876
rect 13688 -8910 13872 -8876
rect 14146 -8910 14330 -8876
rect 14604 -8910 14788 -8876
rect 15062 -8910 15246 -8876
rect 15520 -8910 15704 -8876
rect 16398 -8910 16582 -8876
rect 16856 -8910 17040 -8876
rect 17314 -8910 17498 -8876
rect 17772 -8910 17956 -8876
rect 18230 -8910 18414 -8876
rect 18688 -8910 18872 -8876
rect 19146 -8910 19330 -8876
rect 19604 -8910 19788 -8876
rect 20062 -8910 20246 -8876
rect 20520 -8910 20704 -8876
rect 11398 -9268 11582 -9234
rect 11856 -9268 12040 -9234
rect 12314 -9268 12498 -9234
rect 12772 -9268 12956 -9234
rect 13230 -9268 13414 -9234
rect 13688 -9268 13872 -9234
rect 14146 -9268 14330 -9234
rect 14604 -9268 14788 -9234
rect 15062 -9268 15246 -9234
rect 15520 -9268 15704 -9234
rect 11244 -9494 11278 -9318
rect 11702 -9494 11736 -9318
rect 12160 -9494 12194 -9318
rect 12618 -9494 12652 -9318
rect 13076 -9494 13110 -9318
rect 13534 -9494 13568 -9318
rect 13992 -9494 14026 -9318
rect 14450 -9494 14484 -9318
rect 14908 -9494 14942 -9318
rect 15366 -9494 15400 -9318
rect 15824 -9494 15858 -9318
rect 11398 -9578 11582 -9544
rect 11856 -9578 12040 -9544
rect 12314 -9578 12498 -9544
rect 12772 -9578 12956 -9544
rect 13230 -9578 13414 -9544
rect 13688 -9578 13872 -9544
rect 14146 -9578 14330 -9544
rect 14604 -9578 14788 -9544
rect 15062 -9578 15246 -9544
rect 15520 -9578 15704 -9544
rect 21162 -10342 21262 -8338
rect 10918 -10572 10980 -10472
rect 10980 -10572 21100 -10472
rect 21100 -10572 21162 -10472
rect 25918 -8208 25980 -8108
rect 25980 -8208 36100 -8108
rect 36100 -8208 36162 -8108
rect 25818 -10342 25918 -8338
rect 26398 -8600 26582 -8566
rect 26856 -8600 27040 -8566
rect 27314 -8600 27498 -8566
rect 27772 -8600 27956 -8566
rect 28230 -8600 28414 -8566
rect 28688 -8600 28872 -8566
rect 29146 -8600 29330 -8566
rect 29604 -8600 29788 -8566
rect 30062 -8600 30246 -8566
rect 30520 -8600 30704 -8566
rect 31398 -8600 31582 -8566
rect 31856 -8600 32040 -8566
rect 32314 -8600 32498 -8566
rect 32772 -8600 32956 -8566
rect 33230 -8600 33414 -8566
rect 33688 -8600 33872 -8566
rect 34146 -8600 34330 -8566
rect 34604 -8600 34788 -8566
rect 35062 -8600 35246 -8566
rect 35520 -8600 35704 -8566
rect 26244 -8826 26278 -8650
rect 26702 -8826 26736 -8650
rect 27160 -8826 27194 -8650
rect 27618 -8826 27652 -8650
rect 28076 -8826 28110 -8650
rect 28534 -8826 28568 -8650
rect 28992 -8826 29026 -8650
rect 29450 -8826 29484 -8650
rect 29908 -8826 29942 -8650
rect 30366 -8826 30400 -8650
rect 30824 -8826 30858 -8650
rect 31244 -8826 31278 -8650
rect 31702 -8826 31736 -8650
rect 32160 -8826 32194 -8650
rect 32618 -8826 32652 -8650
rect 33076 -8826 33110 -8650
rect 33534 -8826 33568 -8650
rect 33992 -8826 34026 -8650
rect 34450 -8826 34484 -8650
rect 34908 -8826 34942 -8650
rect 35366 -8826 35400 -8650
rect 35824 -8826 35858 -8650
rect 26398 -8910 26582 -8876
rect 26856 -8910 27040 -8876
rect 27314 -8910 27498 -8876
rect 27772 -8910 27956 -8876
rect 28230 -8910 28414 -8876
rect 28688 -8910 28872 -8876
rect 29146 -8910 29330 -8876
rect 29604 -8910 29788 -8876
rect 30062 -8910 30246 -8876
rect 30520 -8910 30704 -8876
rect 31398 -8910 31582 -8876
rect 31856 -8910 32040 -8876
rect 32314 -8910 32498 -8876
rect 32772 -8910 32956 -8876
rect 33230 -8910 33414 -8876
rect 33688 -8910 33872 -8876
rect 34146 -8910 34330 -8876
rect 34604 -8910 34788 -8876
rect 35062 -8910 35246 -8876
rect 35520 -8910 35704 -8876
rect 26398 -9268 26582 -9234
rect 26856 -9268 27040 -9234
rect 27314 -9268 27498 -9234
rect 27772 -9268 27956 -9234
rect 28230 -9268 28414 -9234
rect 28688 -9268 28872 -9234
rect 29146 -9268 29330 -9234
rect 29604 -9268 29788 -9234
rect 30062 -9268 30246 -9234
rect 30520 -9268 30704 -9234
rect 26244 -9494 26278 -9318
rect 26702 -9494 26736 -9318
rect 27160 -9494 27194 -9318
rect 27618 -9494 27652 -9318
rect 28076 -9494 28110 -9318
rect 28534 -9494 28568 -9318
rect 28992 -9494 29026 -9318
rect 29450 -9494 29484 -9318
rect 29908 -9494 29942 -9318
rect 30366 -9494 30400 -9318
rect 30824 -9494 30858 -9318
rect 26398 -9578 26582 -9544
rect 26856 -9578 27040 -9544
rect 27314 -9578 27498 -9544
rect 27772 -9578 27956 -9544
rect 28230 -9578 28414 -9544
rect 28688 -9578 28872 -9544
rect 29146 -9578 29330 -9544
rect 29604 -9578 29788 -9544
rect 30062 -9578 30246 -9544
rect 30520 -9578 30704 -9544
rect 36162 -10342 36262 -8338
rect 25918 -10572 25980 -10472
rect 25980 -10572 36100 -10472
rect 36100 -10572 36162 -10472
rect 14872 -11132 14934 -11032
rect 14934 -11132 25054 -11032
rect 25054 -11132 25116 -11032
rect 14772 -13266 14872 -11262
rect 20330 -12060 20514 -12026
rect 20788 -12060 20972 -12026
rect 21246 -12060 21430 -12026
rect 21704 -12060 21888 -12026
rect 22162 -12060 22346 -12026
rect 22620 -12060 22804 -12026
rect 23078 -12060 23262 -12026
rect 23536 -12060 23720 -12026
rect 23994 -12060 24178 -12026
rect 24452 -12060 24636 -12026
rect 20176 -12286 20210 -12110
rect 20634 -12286 20668 -12110
rect 21092 -12286 21126 -12110
rect 21550 -12286 21584 -12110
rect 22008 -12286 22042 -12110
rect 22466 -12286 22500 -12110
rect 22924 -12286 22958 -12110
rect 23382 -12286 23416 -12110
rect 23840 -12286 23874 -12110
rect 24298 -12286 24332 -12110
rect 24756 -12286 24790 -12110
rect 20330 -12370 20514 -12336
rect 20788 -12370 20972 -12336
rect 21246 -12370 21430 -12336
rect 21704 -12370 21888 -12336
rect 22162 -12370 22346 -12336
rect 22620 -12370 22804 -12336
rect 23078 -12370 23262 -12336
rect 23536 -12370 23720 -12336
rect 23994 -12370 24178 -12336
rect 24452 -12370 24636 -12336
rect 15330 -12728 15514 -12694
rect 15788 -12728 15972 -12694
rect 16246 -12728 16430 -12694
rect 16704 -12728 16888 -12694
rect 17162 -12728 17346 -12694
rect 17620 -12728 17804 -12694
rect 18078 -12728 18262 -12694
rect 18536 -12728 18720 -12694
rect 18994 -12728 19178 -12694
rect 19452 -12728 19636 -12694
rect 20330 -12728 20514 -12694
rect 20788 -12728 20972 -12694
rect 21246 -12728 21430 -12694
rect 21704 -12728 21888 -12694
rect 22162 -12728 22346 -12694
rect 22620 -12728 22804 -12694
rect 23078 -12728 23262 -12694
rect 23536 -12728 23720 -12694
rect 23994 -12728 24178 -12694
rect 24452 -12728 24636 -12694
rect 15176 -12954 15210 -12778
rect 15634 -12954 15668 -12778
rect 16092 -12954 16126 -12778
rect 16550 -12954 16584 -12778
rect 17008 -12954 17042 -12778
rect 17466 -12954 17500 -12778
rect 17924 -12954 17958 -12778
rect 18382 -12954 18416 -12778
rect 18840 -12954 18874 -12778
rect 19298 -12954 19332 -12778
rect 19756 -12954 19790 -12778
rect 20176 -12954 20210 -12778
rect 20634 -12954 20668 -12778
rect 21092 -12954 21126 -12778
rect 21550 -12954 21584 -12778
rect 22008 -12954 22042 -12778
rect 22466 -12954 22500 -12778
rect 22924 -12954 22958 -12778
rect 23382 -12954 23416 -12778
rect 23840 -12954 23874 -12778
rect 24298 -12954 24332 -12778
rect 24756 -12954 24790 -12778
rect 15330 -13038 15514 -13004
rect 15788 -13038 15972 -13004
rect 16246 -13038 16430 -13004
rect 16704 -13038 16888 -13004
rect 17162 -13038 17346 -13004
rect 17620 -13038 17804 -13004
rect 18078 -13038 18262 -13004
rect 18536 -13038 18720 -13004
rect 18994 -13038 19178 -13004
rect 19452 -13038 19636 -13004
rect 20330 -13038 20514 -13004
rect 20788 -13038 20972 -13004
rect 21246 -13038 21430 -13004
rect 21704 -13038 21888 -13004
rect 22162 -13038 22346 -13004
rect 22620 -13038 22804 -13004
rect 23078 -13038 23262 -13004
rect 23536 -13038 23720 -13004
rect 23994 -13038 24178 -13004
rect 24452 -13038 24636 -13004
rect 25116 -13266 25216 -11262
rect 14872 -13496 14934 -13396
rect 14934 -13496 25054 -13396
rect 25054 -13496 25116 -13396
rect 29872 -11132 29934 -11032
rect 29934 -11132 40054 -11032
rect 40054 -11132 40116 -11032
rect 29772 -13266 29872 -11262
rect 35330 -12060 35514 -12026
rect 35788 -12060 35972 -12026
rect 36246 -12060 36430 -12026
rect 36704 -12060 36888 -12026
rect 37162 -12060 37346 -12026
rect 37620 -12060 37804 -12026
rect 38078 -12060 38262 -12026
rect 38536 -12060 38720 -12026
rect 38994 -12060 39178 -12026
rect 39452 -12060 39636 -12026
rect 35176 -12286 35210 -12110
rect 35634 -12286 35668 -12110
rect 36092 -12286 36126 -12110
rect 36550 -12286 36584 -12110
rect 37008 -12286 37042 -12110
rect 37466 -12286 37500 -12110
rect 37924 -12286 37958 -12110
rect 38382 -12286 38416 -12110
rect 38840 -12286 38874 -12110
rect 39298 -12286 39332 -12110
rect 39756 -12286 39790 -12110
rect 35330 -12370 35514 -12336
rect 35788 -12370 35972 -12336
rect 36246 -12370 36430 -12336
rect 36704 -12370 36888 -12336
rect 37162 -12370 37346 -12336
rect 37620 -12370 37804 -12336
rect 38078 -12370 38262 -12336
rect 38536 -12370 38720 -12336
rect 38994 -12370 39178 -12336
rect 39452 -12370 39636 -12336
rect 30330 -12728 30514 -12694
rect 30788 -12728 30972 -12694
rect 31246 -12728 31430 -12694
rect 31704 -12728 31888 -12694
rect 32162 -12728 32346 -12694
rect 32620 -12728 32804 -12694
rect 33078 -12728 33262 -12694
rect 33536 -12728 33720 -12694
rect 33994 -12728 34178 -12694
rect 34452 -12728 34636 -12694
rect 35330 -12728 35514 -12694
rect 35788 -12728 35972 -12694
rect 36246 -12728 36430 -12694
rect 36704 -12728 36888 -12694
rect 37162 -12728 37346 -12694
rect 37620 -12728 37804 -12694
rect 38078 -12728 38262 -12694
rect 38536 -12728 38720 -12694
rect 38994 -12728 39178 -12694
rect 39452 -12728 39636 -12694
rect 30176 -12954 30210 -12778
rect 30634 -12954 30668 -12778
rect 31092 -12954 31126 -12778
rect 31550 -12954 31584 -12778
rect 32008 -12954 32042 -12778
rect 32466 -12954 32500 -12778
rect 32924 -12954 32958 -12778
rect 33382 -12954 33416 -12778
rect 33840 -12954 33874 -12778
rect 34298 -12954 34332 -12778
rect 34756 -12954 34790 -12778
rect 35176 -12954 35210 -12778
rect 35634 -12954 35668 -12778
rect 36092 -12954 36126 -12778
rect 36550 -12954 36584 -12778
rect 37008 -12954 37042 -12778
rect 37466 -12954 37500 -12778
rect 37924 -12954 37958 -12778
rect 38382 -12954 38416 -12778
rect 38840 -12954 38874 -12778
rect 39298 -12954 39332 -12778
rect 39756 -12954 39790 -12778
rect 30330 -13038 30514 -13004
rect 30788 -13038 30972 -13004
rect 31246 -13038 31430 -13004
rect 31704 -13038 31888 -13004
rect 32162 -13038 32346 -13004
rect 32620 -13038 32804 -13004
rect 33078 -13038 33262 -13004
rect 33536 -13038 33720 -13004
rect 33994 -13038 34178 -13004
rect 34452 -13038 34636 -13004
rect 35330 -13038 35514 -13004
rect 35788 -13038 35972 -13004
rect 36246 -13038 36430 -13004
rect 36704 -13038 36888 -13004
rect 37162 -13038 37346 -13004
rect 37620 -13038 37804 -13004
rect 38078 -13038 38262 -13004
rect 38536 -13038 38720 -13004
rect 38994 -13038 39178 -13004
rect 39452 -13038 39636 -13004
rect 40116 -13266 40216 -11262
rect 29872 -13496 29934 -13396
rect 29934 -13496 40054 -13396
rect 40054 -13496 40116 -13396
rect 14872 -13832 14934 -13732
rect 14934 -13832 25054 -13732
rect 25054 -13832 25116 -13732
rect 14772 -19186 14872 -14014
rect 15329 -14212 15513 -14178
rect 15787 -14212 15971 -14178
rect 16245 -14212 16429 -14178
rect 16703 -14212 16887 -14178
rect 17161 -14212 17345 -14178
rect 17619 -14212 17803 -14178
rect 18077 -14212 18261 -14178
rect 18535 -14212 18719 -14178
rect 18993 -14212 19177 -14178
rect 19451 -14212 19635 -14178
rect 20329 -14212 20513 -14178
rect 20787 -14212 20971 -14178
rect 21245 -14212 21429 -14178
rect 21703 -14212 21887 -14178
rect 22161 -14212 22345 -14178
rect 22619 -14212 22803 -14178
rect 23077 -14212 23261 -14178
rect 23535 -14212 23719 -14178
rect 23993 -14212 24177 -14178
rect 24451 -14212 24635 -14178
rect 15175 -15447 15209 -14271
rect 15633 -15447 15667 -14271
rect 16091 -15447 16125 -14271
rect 16549 -15447 16583 -14271
rect 17007 -15447 17041 -14271
rect 17465 -15447 17499 -14271
rect 17923 -15447 17957 -14271
rect 18381 -15447 18415 -14271
rect 18839 -15447 18873 -14271
rect 19297 -15447 19331 -14271
rect 19755 -15447 19789 -14271
rect 20175 -15447 20209 -14271
rect 20633 -15447 20667 -14271
rect 21091 -15447 21125 -14271
rect 21549 -15447 21583 -14271
rect 22007 -15447 22041 -14271
rect 22465 -15447 22499 -14271
rect 22923 -15447 22957 -14271
rect 23381 -15447 23415 -14271
rect 23839 -15447 23873 -14271
rect 24297 -15447 24331 -14271
rect 24755 -15447 24789 -14271
rect 15329 -15540 15513 -15506
rect 15787 -15540 15971 -15506
rect 16245 -15540 16429 -15506
rect 16703 -15540 16887 -15506
rect 17161 -15540 17345 -15506
rect 17619 -15540 17803 -15506
rect 18077 -15540 18261 -15506
rect 18535 -15540 18719 -15506
rect 18993 -15540 19177 -15506
rect 19451 -15540 19635 -15506
rect 20329 -15540 20513 -15506
rect 20787 -15540 20971 -15506
rect 21245 -15540 21429 -15506
rect 21703 -15540 21887 -15506
rect 22161 -15540 22345 -15506
rect 22619 -15540 22803 -15506
rect 23077 -15540 23261 -15506
rect 23535 -15540 23719 -15506
rect 23993 -15540 24177 -15506
rect 24451 -15540 24635 -15506
rect 19832 -16366 19892 -16306
rect 20298 -16360 20346 -16312
rect 16106 -16477 16290 -16443
rect 16564 -16477 16748 -16443
rect 17022 -16477 17206 -16443
rect 17480 -16477 17664 -16443
rect 17938 -16477 18122 -16443
rect 18396 -16477 18580 -16443
rect 18854 -16477 19038 -16443
rect 19312 -16477 19496 -16443
rect 19770 -16477 19954 -16443
rect 20228 -16477 20412 -16443
rect 20686 -16477 20870 -16443
rect 21144 -16477 21328 -16443
rect 21602 -16477 21786 -16443
rect 22060 -16477 22244 -16443
rect 22518 -16477 22702 -16443
rect 22976 -16477 23160 -16443
rect 23434 -16477 23618 -16443
rect 23892 -16477 24076 -16443
rect 15952 -18112 15986 -16536
rect 16410 -18112 16444 -16536
rect 16868 -18112 16902 -16536
rect 17326 -18112 17360 -16536
rect 17784 -18112 17818 -16536
rect 18242 -18112 18276 -16536
rect 18700 -18112 18734 -16536
rect 19158 -18112 19192 -16536
rect 19616 -18112 19650 -16536
rect 20074 -18112 20108 -16536
rect 20532 -18112 20566 -16536
rect 20990 -18112 21024 -16536
rect 21448 -18112 21482 -16536
rect 21906 -18112 21940 -16536
rect 22364 -18112 22398 -16536
rect 22822 -18112 22856 -16536
rect 23280 -18112 23314 -16536
rect 23738 -18112 23772 -16536
rect 24196 -18112 24230 -16536
rect 16106 -18205 16290 -18171
rect 16564 -18205 16748 -18171
rect 17022 -18205 17206 -18171
rect 17480 -18205 17664 -18171
rect 17938 -18205 18122 -18171
rect 18396 -18205 18580 -18171
rect 18854 -18205 19038 -18171
rect 19312 -18205 19496 -18171
rect 19770 -18205 19954 -18171
rect 20228 -18205 20412 -18171
rect 20686 -18205 20870 -18171
rect 21144 -18205 21328 -18171
rect 21602 -18205 21786 -18171
rect 22060 -18205 22244 -18171
rect 22518 -18205 22702 -18171
rect 22976 -18205 23160 -18171
rect 23434 -18205 23618 -18171
rect 23892 -18205 24076 -18171
rect 25116 -19186 25216 -14014
rect 14872 -19576 14934 -19476
rect 14934 -19576 25054 -19476
rect 25054 -19576 25116 -19476
rect 29872 -13832 29934 -13732
rect 29934 -13832 40054 -13732
rect 40054 -13832 40116 -13732
rect 29772 -19186 29872 -14014
rect 30329 -14212 30513 -14178
rect 30787 -14212 30971 -14178
rect 31245 -14212 31429 -14178
rect 31703 -14212 31887 -14178
rect 32161 -14212 32345 -14178
rect 32619 -14212 32803 -14178
rect 33077 -14212 33261 -14178
rect 33535 -14212 33719 -14178
rect 33993 -14212 34177 -14178
rect 34451 -14212 34635 -14178
rect 35329 -14212 35513 -14178
rect 35787 -14212 35971 -14178
rect 36245 -14212 36429 -14178
rect 36703 -14212 36887 -14178
rect 37161 -14212 37345 -14178
rect 37619 -14212 37803 -14178
rect 38077 -14212 38261 -14178
rect 38535 -14212 38719 -14178
rect 38993 -14212 39177 -14178
rect 39451 -14212 39635 -14178
rect 30175 -15447 30209 -14271
rect 30633 -15447 30667 -14271
rect 31091 -15447 31125 -14271
rect 31549 -15447 31583 -14271
rect 32007 -15447 32041 -14271
rect 32465 -15447 32499 -14271
rect 32923 -15447 32957 -14271
rect 33381 -15447 33415 -14271
rect 33839 -15447 33873 -14271
rect 34297 -15447 34331 -14271
rect 34755 -15447 34789 -14271
rect 35175 -15447 35209 -14271
rect 35633 -15447 35667 -14271
rect 36091 -15447 36125 -14271
rect 36549 -15447 36583 -14271
rect 37007 -15447 37041 -14271
rect 37465 -15447 37499 -14271
rect 37923 -15447 37957 -14271
rect 38381 -15447 38415 -14271
rect 38839 -15447 38873 -14271
rect 39297 -15447 39331 -14271
rect 39755 -15447 39789 -14271
rect 30329 -15540 30513 -15506
rect 30787 -15540 30971 -15506
rect 31245 -15540 31429 -15506
rect 31703 -15540 31887 -15506
rect 32161 -15540 32345 -15506
rect 32619 -15540 32803 -15506
rect 33077 -15540 33261 -15506
rect 33535 -15540 33719 -15506
rect 33993 -15540 34177 -15506
rect 34451 -15540 34635 -15506
rect 35329 -15540 35513 -15506
rect 35787 -15540 35971 -15506
rect 36245 -15540 36429 -15506
rect 36703 -15540 36887 -15506
rect 37161 -15540 37345 -15506
rect 37619 -15540 37803 -15506
rect 38077 -15540 38261 -15506
rect 38535 -15540 38719 -15506
rect 38993 -15540 39177 -15506
rect 39451 -15540 39635 -15506
rect 34832 -16366 34892 -16306
rect 35298 -16360 35346 -16312
rect 31106 -16477 31290 -16443
rect 31564 -16477 31748 -16443
rect 32022 -16477 32206 -16443
rect 32480 -16477 32664 -16443
rect 32938 -16477 33122 -16443
rect 33396 -16477 33580 -16443
rect 33854 -16477 34038 -16443
rect 34312 -16477 34496 -16443
rect 34770 -16477 34954 -16443
rect 35228 -16477 35412 -16443
rect 35686 -16477 35870 -16443
rect 36144 -16477 36328 -16443
rect 36602 -16477 36786 -16443
rect 37060 -16477 37244 -16443
rect 37518 -16477 37702 -16443
rect 37976 -16477 38160 -16443
rect 38434 -16477 38618 -16443
rect 38892 -16477 39076 -16443
rect 30952 -18112 30986 -16536
rect 31410 -18112 31444 -16536
rect 31868 -18112 31902 -16536
rect 32326 -18112 32360 -16536
rect 32784 -18112 32818 -16536
rect 33242 -18112 33276 -16536
rect 33700 -18112 33734 -16536
rect 34158 -18112 34192 -16536
rect 34616 -18112 34650 -16536
rect 35074 -18112 35108 -16536
rect 35532 -18112 35566 -16536
rect 35990 -18112 36024 -16536
rect 36448 -18112 36482 -16536
rect 36906 -18112 36940 -16536
rect 37364 -18112 37398 -16536
rect 37822 -18112 37856 -16536
rect 38280 -18112 38314 -16536
rect 38738 -18112 38772 -16536
rect 39196 -18112 39230 -16536
rect 31106 -18205 31290 -18171
rect 31564 -18205 31748 -18171
rect 32022 -18205 32206 -18171
rect 32480 -18205 32664 -18171
rect 32938 -18205 33122 -18171
rect 33396 -18205 33580 -18171
rect 33854 -18205 34038 -18171
rect 34312 -18205 34496 -18171
rect 34770 -18205 34954 -18171
rect 35228 -18205 35412 -18171
rect 35686 -18205 35870 -18171
rect 36144 -18205 36328 -18171
rect 36602 -18205 36786 -18171
rect 37060 -18205 37244 -18171
rect 37518 -18205 37702 -18171
rect 37976 -18205 38160 -18171
rect 38434 -18205 38618 -18171
rect 38892 -18205 39076 -18171
rect 40116 -19186 40216 -14014
rect 29872 -19576 29934 -19476
rect 29934 -19576 40054 -19476
rect 40054 -19576 40116 -19476
rect 10918 -20128 10980 -20028
rect 10980 -20128 21100 -20028
rect 21100 -20128 21162 -20028
rect 10818 -25590 10918 -20418
rect 11958 -21433 12142 -21399
rect 12416 -21433 12600 -21399
rect 12874 -21433 13058 -21399
rect 13332 -21433 13516 -21399
rect 13790 -21433 13974 -21399
rect 14248 -21433 14432 -21399
rect 14706 -21433 14890 -21399
rect 15164 -21433 15348 -21399
rect 15622 -21433 15806 -21399
rect 16080 -21433 16264 -21399
rect 16538 -21433 16722 -21399
rect 16996 -21433 17180 -21399
rect 17454 -21433 17638 -21399
rect 17912 -21433 18096 -21399
rect 18370 -21433 18554 -21399
rect 18828 -21433 19012 -21399
rect 19286 -21433 19470 -21399
rect 19744 -21433 19928 -21399
rect 11804 -23068 11838 -21492
rect 12262 -23068 12296 -21492
rect 12720 -23068 12754 -21492
rect 13178 -23068 13212 -21492
rect 13636 -23068 13670 -21492
rect 14094 -23068 14128 -21492
rect 14552 -23068 14586 -21492
rect 15010 -23068 15044 -21492
rect 15468 -23068 15502 -21492
rect 15926 -23068 15960 -21492
rect 16384 -23068 16418 -21492
rect 16842 -23068 16876 -21492
rect 17300 -23068 17334 -21492
rect 17758 -23068 17792 -21492
rect 18216 -23068 18250 -21492
rect 18674 -23068 18708 -21492
rect 19132 -23068 19166 -21492
rect 19590 -23068 19624 -21492
rect 20048 -23068 20082 -21492
rect 11958 -23161 12142 -23127
rect 12416 -23161 12600 -23127
rect 12874 -23161 13058 -23127
rect 13332 -23161 13516 -23127
rect 13790 -23161 13974 -23127
rect 14248 -23161 14432 -23127
rect 14706 -23161 14890 -23127
rect 15164 -23161 15348 -23127
rect 15622 -23161 15806 -23127
rect 16080 -23161 16264 -23127
rect 16538 -23161 16722 -23127
rect 16996 -23161 17180 -23127
rect 17454 -23161 17638 -23127
rect 17912 -23161 18096 -23127
rect 18370 -23161 18554 -23127
rect 18828 -23161 19012 -23127
rect 19286 -23161 19470 -23127
rect 19744 -23161 19928 -23127
rect 15688 -23292 15736 -23244
rect 16142 -23298 16202 -23238
rect 11399 -24098 11583 -24064
rect 11857 -24098 12041 -24064
rect 12315 -24098 12499 -24064
rect 12773 -24098 12957 -24064
rect 13231 -24098 13415 -24064
rect 13689 -24098 13873 -24064
rect 14147 -24098 14331 -24064
rect 14605 -24098 14789 -24064
rect 15063 -24098 15247 -24064
rect 15521 -24098 15705 -24064
rect 16399 -24098 16583 -24064
rect 16857 -24098 17041 -24064
rect 17315 -24098 17499 -24064
rect 17773 -24098 17957 -24064
rect 18231 -24098 18415 -24064
rect 18689 -24098 18873 -24064
rect 19147 -24098 19331 -24064
rect 19605 -24098 19789 -24064
rect 20063 -24098 20247 -24064
rect 20521 -24098 20705 -24064
rect 11245 -25333 11279 -24157
rect 11703 -25333 11737 -24157
rect 12161 -25333 12195 -24157
rect 12619 -25333 12653 -24157
rect 13077 -25333 13111 -24157
rect 13535 -25333 13569 -24157
rect 13993 -25333 14027 -24157
rect 14451 -25333 14485 -24157
rect 14909 -25333 14943 -24157
rect 15367 -25333 15401 -24157
rect 15825 -25333 15859 -24157
rect 16245 -25333 16279 -24157
rect 16703 -25333 16737 -24157
rect 17161 -25333 17195 -24157
rect 17619 -25333 17653 -24157
rect 18077 -25333 18111 -24157
rect 18535 -25333 18569 -24157
rect 18993 -25333 19027 -24157
rect 19451 -25333 19485 -24157
rect 19909 -25333 19943 -24157
rect 20367 -25333 20401 -24157
rect 20825 -25333 20859 -24157
rect 11399 -25426 11583 -25392
rect 11857 -25426 12041 -25392
rect 12315 -25426 12499 -25392
rect 12773 -25426 12957 -25392
rect 13231 -25426 13415 -25392
rect 13689 -25426 13873 -25392
rect 14147 -25426 14331 -25392
rect 14605 -25426 14789 -25392
rect 15063 -25426 15247 -25392
rect 15521 -25426 15705 -25392
rect 16399 -25426 16583 -25392
rect 16857 -25426 17041 -25392
rect 17315 -25426 17499 -25392
rect 17773 -25426 17957 -25392
rect 18231 -25426 18415 -25392
rect 18689 -25426 18873 -25392
rect 19147 -25426 19331 -25392
rect 19605 -25426 19789 -25392
rect 20063 -25426 20247 -25392
rect 20521 -25426 20705 -25392
rect 21162 -25590 21262 -20418
rect 10918 -25872 10980 -25772
rect 10980 -25872 21100 -25772
rect 21100 -25872 21162 -25772
rect 25918 -20128 25980 -20028
rect 25980 -20128 36100 -20028
rect 36100 -20128 36162 -20028
rect 25818 -25590 25918 -20418
rect 26958 -21433 27142 -21399
rect 27416 -21433 27600 -21399
rect 27874 -21433 28058 -21399
rect 28332 -21433 28516 -21399
rect 28790 -21433 28974 -21399
rect 29248 -21433 29432 -21399
rect 29706 -21433 29890 -21399
rect 30164 -21433 30348 -21399
rect 30622 -21433 30806 -21399
rect 31080 -21433 31264 -21399
rect 31538 -21433 31722 -21399
rect 31996 -21433 32180 -21399
rect 32454 -21433 32638 -21399
rect 32912 -21433 33096 -21399
rect 33370 -21433 33554 -21399
rect 33828 -21433 34012 -21399
rect 34286 -21433 34470 -21399
rect 34744 -21433 34928 -21399
rect 26804 -23068 26838 -21492
rect 27262 -23068 27296 -21492
rect 27720 -23068 27754 -21492
rect 28178 -23068 28212 -21492
rect 28636 -23068 28670 -21492
rect 29094 -23068 29128 -21492
rect 29552 -23068 29586 -21492
rect 30010 -23068 30044 -21492
rect 30468 -23068 30502 -21492
rect 30926 -23068 30960 -21492
rect 31384 -23068 31418 -21492
rect 31842 -23068 31876 -21492
rect 32300 -23068 32334 -21492
rect 32758 -23068 32792 -21492
rect 33216 -23068 33250 -21492
rect 33674 -23068 33708 -21492
rect 34132 -23068 34166 -21492
rect 34590 -23068 34624 -21492
rect 35048 -23068 35082 -21492
rect 26958 -23161 27142 -23127
rect 27416 -23161 27600 -23127
rect 27874 -23161 28058 -23127
rect 28332 -23161 28516 -23127
rect 28790 -23161 28974 -23127
rect 29248 -23161 29432 -23127
rect 29706 -23161 29890 -23127
rect 30164 -23161 30348 -23127
rect 30622 -23161 30806 -23127
rect 31080 -23161 31264 -23127
rect 31538 -23161 31722 -23127
rect 31996 -23161 32180 -23127
rect 32454 -23161 32638 -23127
rect 32912 -23161 33096 -23127
rect 33370 -23161 33554 -23127
rect 33828 -23161 34012 -23127
rect 34286 -23161 34470 -23127
rect 34744 -23161 34928 -23127
rect 30688 -23292 30736 -23244
rect 31142 -23298 31202 -23238
rect 26399 -24098 26583 -24064
rect 26857 -24098 27041 -24064
rect 27315 -24098 27499 -24064
rect 27773 -24098 27957 -24064
rect 28231 -24098 28415 -24064
rect 28689 -24098 28873 -24064
rect 29147 -24098 29331 -24064
rect 29605 -24098 29789 -24064
rect 30063 -24098 30247 -24064
rect 30521 -24098 30705 -24064
rect 31399 -24098 31583 -24064
rect 31857 -24098 32041 -24064
rect 32315 -24098 32499 -24064
rect 32773 -24098 32957 -24064
rect 33231 -24098 33415 -24064
rect 33689 -24098 33873 -24064
rect 34147 -24098 34331 -24064
rect 34605 -24098 34789 -24064
rect 35063 -24098 35247 -24064
rect 35521 -24098 35705 -24064
rect 26245 -25333 26279 -24157
rect 26703 -25333 26737 -24157
rect 27161 -25333 27195 -24157
rect 27619 -25333 27653 -24157
rect 28077 -25333 28111 -24157
rect 28535 -25333 28569 -24157
rect 28993 -25333 29027 -24157
rect 29451 -25333 29485 -24157
rect 29909 -25333 29943 -24157
rect 30367 -25333 30401 -24157
rect 30825 -25333 30859 -24157
rect 31245 -25333 31279 -24157
rect 31703 -25333 31737 -24157
rect 32161 -25333 32195 -24157
rect 32619 -25333 32653 -24157
rect 33077 -25333 33111 -24157
rect 33535 -25333 33569 -24157
rect 33993 -25333 34027 -24157
rect 34451 -25333 34485 -24157
rect 34909 -25333 34943 -24157
rect 35367 -25333 35401 -24157
rect 35825 -25333 35859 -24157
rect 26399 -25426 26583 -25392
rect 26857 -25426 27041 -25392
rect 27315 -25426 27499 -25392
rect 27773 -25426 27957 -25392
rect 28231 -25426 28415 -25392
rect 28689 -25426 28873 -25392
rect 29147 -25426 29331 -25392
rect 29605 -25426 29789 -25392
rect 30063 -25426 30247 -25392
rect 30521 -25426 30705 -25392
rect 31399 -25426 31583 -25392
rect 31857 -25426 32041 -25392
rect 32315 -25426 32499 -25392
rect 32773 -25426 32957 -25392
rect 33231 -25426 33415 -25392
rect 33689 -25426 33873 -25392
rect 34147 -25426 34331 -25392
rect 34605 -25426 34789 -25392
rect 35063 -25426 35247 -25392
rect 35521 -25426 35705 -25392
rect 36162 -25590 36262 -20418
rect 25918 -25872 25980 -25772
rect 25980 -25872 36100 -25772
rect 36100 -25872 36162 -25772
rect 10918 -26208 10980 -26108
rect 10980 -26208 21100 -26108
rect 21100 -26208 21162 -26108
rect 10818 -28342 10918 -26338
rect 11398 -26600 11582 -26566
rect 11856 -26600 12040 -26566
rect 12314 -26600 12498 -26566
rect 12772 -26600 12956 -26566
rect 13230 -26600 13414 -26566
rect 13688 -26600 13872 -26566
rect 14146 -26600 14330 -26566
rect 14604 -26600 14788 -26566
rect 15062 -26600 15246 -26566
rect 15520 -26600 15704 -26566
rect 16398 -26600 16582 -26566
rect 16856 -26600 17040 -26566
rect 17314 -26600 17498 -26566
rect 17772 -26600 17956 -26566
rect 18230 -26600 18414 -26566
rect 18688 -26600 18872 -26566
rect 19146 -26600 19330 -26566
rect 19604 -26600 19788 -26566
rect 20062 -26600 20246 -26566
rect 20520 -26600 20704 -26566
rect 11244 -26826 11278 -26650
rect 11702 -26826 11736 -26650
rect 12160 -26826 12194 -26650
rect 12618 -26826 12652 -26650
rect 13076 -26826 13110 -26650
rect 13534 -26826 13568 -26650
rect 13992 -26826 14026 -26650
rect 14450 -26826 14484 -26650
rect 14908 -26826 14942 -26650
rect 15366 -26826 15400 -26650
rect 15824 -26826 15858 -26650
rect 16244 -26826 16278 -26650
rect 16702 -26826 16736 -26650
rect 17160 -26826 17194 -26650
rect 17618 -26826 17652 -26650
rect 18076 -26826 18110 -26650
rect 18534 -26826 18568 -26650
rect 18992 -26826 19026 -26650
rect 19450 -26826 19484 -26650
rect 19908 -26826 19942 -26650
rect 20366 -26826 20400 -26650
rect 20824 -26826 20858 -26650
rect 11398 -26910 11582 -26876
rect 11856 -26910 12040 -26876
rect 12314 -26910 12498 -26876
rect 12772 -26910 12956 -26876
rect 13230 -26910 13414 -26876
rect 13688 -26910 13872 -26876
rect 14146 -26910 14330 -26876
rect 14604 -26910 14788 -26876
rect 15062 -26910 15246 -26876
rect 15520 -26910 15704 -26876
rect 16398 -26910 16582 -26876
rect 16856 -26910 17040 -26876
rect 17314 -26910 17498 -26876
rect 17772 -26910 17956 -26876
rect 18230 -26910 18414 -26876
rect 18688 -26910 18872 -26876
rect 19146 -26910 19330 -26876
rect 19604 -26910 19788 -26876
rect 20062 -26910 20246 -26876
rect 20520 -26910 20704 -26876
rect 11398 -27268 11582 -27234
rect 11856 -27268 12040 -27234
rect 12314 -27268 12498 -27234
rect 12772 -27268 12956 -27234
rect 13230 -27268 13414 -27234
rect 13688 -27268 13872 -27234
rect 14146 -27268 14330 -27234
rect 14604 -27268 14788 -27234
rect 15062 -27268 15246 -27234
rect 15520 -27268 15704 -27234
rect 11244 -27494 11278 -27318
rect 11702 -27494 11736 -27318
rect 12160 -27494 12194 -27318
rect 12618 -27494 12652 -27318
rect 13076 -27494 13110 -27318
rect 13534 -27494 13568 -27318
rect 13992 -27494 14026 -27318
rect 14450 -27494 14484 -27318
rect 14908 -27494 14942 -27318
rect 15366 -27494 15400 -27318
rect 15824 -27494 15858 -27318
rect 11398 -27578 11582 -27544
rect 11856 -27578 12040 -27544
rect 12314 -27578 12498 -27544
rect 12772 -27578 12956 -27544
rect 13230 -27578 13414 -27544
rect 13688 -27578 13872 -27544
rect 14146 -27578 14330 -27544
rect 14604 -27578 14788 -27544
rect 15062 -27578 15246 -27544
rect 15520 -27578 15704 -27544
rect 21162 -28342 21262 -26338
rect 10918 -28572 10980 -28472
rect 10980 -28572 21100 -28472
rect 21100 -28572 21162 -28472
rect 25918 -26208 25980 -26108
rect 25980 -26208 36100 -26108
rect 36100 -26208 36162 -26108
rect 25818 -28342 25918 -26338
rect 26398 -26600 26582 -26566
rect 26856 -26600 27040 -26566
rect 27314 -26600 27498 -26566
rect 27772 -26600 27956 -26566
rect 28230 -26600 28414 -26566
rect 28688 -26600 28872 -26566
rect 29146 -26600 29330 -26566
rect 29604 -26600 29788 -26566
rect 30062 -26600 30246 -26566
rect 30520 -26600 30704 -26566
rect 31398 -26600 31582 -26566
rect 31856 -26600 32040 -26566
rect 32314 -26600 32498 -26566
rect 32772 -26600 32956 -26566
rect 33230 -26600 33414 -26566
rect 33688 -26600 33872 -26566
rect 34146 -26600 34330 -26566
rect 34604 -26600 34788 -26566
rect 35062 -26600 35246 -26566
rect 35520 -26600 35704 -26566
rect 26244 -26826 26278 -26650
rect 26702 -26826 26736 -26650
rect 27160 -26826 27194 -26650
rect 27618 -26826 27652 -26650
rect 28076 -26826 28110 -26650
rect 28534 -26826 28568 -26650
rect 28992 -26826 29026 -26650
rect 29450 -26826 29484 -26650
rect 29908 -26826 29942 -26650
rect 30366 -26826 30400 -26650
rect 30824 -26826 30858 -26650
rect 31244 -26826 31278 -26650
rect 31702 -26826 31736 -26650
rect 32160 -26826 32194 -26650
rect 32618 -26826 32652 -26650
rect 33076 -26826 33110 -26650
rect 33534 -26826 33568 -26650
rect 33992 -26826 34026 -26650
rect 34450 -26826 34484 -26650
rect 34908 -26826 34942 -26650
rect 35366 -26826 35400 -26650
rect 35824 -26826 35858 -26650
rect 26398 -26910 26582 -26876
rect 26856 -26910 27040 -26876
rect 27314 -26910 27498 -26876
rect 27772 -26910 27956 -26876
rect 28230 -26910 28414 -26876
rect 28688 -26910 28872 -26876
rect 29146 -26910 29330 -26876
rect 29604 -26910 29788 -26876
rect 30062 -26910 30246 -26876
rect 30520 -26910 30704 -26876
rect 31398 -26910 31582 -26876
rect 31856 -26910 32040 -26876
rect 32314 -26910 32498 -26876
rect 32772 -26910 32956 -26876
rect 33230 -26910 33414 -26876
rect 33688 -26910 33872 -26876
rect 34146 -26910 34330 -26876
rect 34604 -26910 34788 -26876
rect 35062 -26910 35246 -26876
rect 35520 -26910 35704 -26876
rect 26398 -27268 26582 -27234
rect 26856 -27268 27040 -27234
rect 27314 -27268 27498 -27234
rect 27772 -27268 27956 -27234
rect 28230 -27268 28414 -27234
rect 28688 -27268 28872 -27234
rect 29146 -27268 29330 -27234
rect 29604 -27268 29788 -27234
rect 30062 -27268 30246 -27234
rect 30520 -27268 30704 -27234
rect 26244 -27494 26278 -27318
rect 26702 -27494 26736 -27318
rect 27160 -27494 27194 -27318
rect 27618 -27494 27652 -27318
rect 28076 -27494 28110 -27318
rect 28534 -27494 28568 -27318
rect 28992 -27494 29026 -27318
rect 29450 -27494 29484 -27318
rect 29908 -27494 29942 -27318
rect 30366 -27494 30400 -27318
rect 30824 -27494 30858 -27318
rect 26398 -27578 26582 -27544
rect 26856 -27578 27040 -27544
rect 27314 -27578 27498 -27544
rect 27772 -27578 27956 -27544
rect 28230 -27578 28414 -27544
rect 28688 -27578 28872 -27544
rect 29146 -27578 29330 -27544
rect 29604 -27578 29788 -27544
rect 30062 -27578 30246 -27544
rect 30520 -27578 30704 -27544
rect 36162 -28342 36262 -26338
rect 25918 -28572 25980 -28472
rect 25980 -28572 36100 -28472
rect 36100 -28572 36162 -28472
<< metal1 >>
rect 15420 4310 24456 4316
rect 15420 4210 15526 4310
rect 24350 4210 24456 4310
rect 15420 4204 24456 4210
rect 15420 4122 15532 4204
rect 15420 2698 15426 4122
rect 15526 2698 15532 4122
rect 15914 3904 15924 4204
rect 23656 3904 23666 4204
rect 24344 4122 24456 4204
rect 17550 3726 22522 3756
rect 17550 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 22522 3726
rect 17550 3612 22522 3640
rect 17614 3232 17674 3612
rect 17854 3322 17914 3612
rect 18304 3388 21514 3448
rect 21574 3388 21580 3448
rect 18304 3322 18364 3388
rect 18766 3322 18826 3388
rect 19220 3322 19280 3388
rect 19682 3322 19742 3388
rect 20136 3322 20196 3388
rect 20586 3322 20646 3388
rect 21052 3322 21112 3388
rect 21508 3322 21568 3388
rect 17776 3316 17984 3322
rect 17776 3282 17788 3316
rect 17972 3282 17984 3316
rect 17776 3276 17984 3282
rect 18234 3316 18442 3322
rect 18234 3282 18246 3316
rect 18430 3282 18442 3316
rect 18234 3276 18442 3282
rect 18692 3316 18900 3322
rect 18692 3282 18704 3316
rect 18888 3282 18900 3316
rect 18692 3276 18900 3282
rect 19150 3316 19358 3322
rect 19150 3282 19162 3316
rect 19346 3282 19358 3316
rect 19150 3276 19358 3282
rect 19608 3316 19816 3322
rect 19608 3282 19620 3316
rect 19804 3282 19816 3316
rect 19608 3276 19816 3282
rect 20066 3316 20274 3322
rect 20066 3282 20078 3316
rect 20262 3282 20274 3316
rect 20066 3276 20274 3282
rect 20524 3316 20732 3322
rect 20524 3282 20536 3316
rect 20720 3282 20732 3316
rect 20524 3276 20732 3282
rect 20982 3316 21190 3322
rect 20982 3282 20994 3316
rect 21178 3282 21190 3316
rect 20982 3276 21190 3282
rect 21440 3316 21648 3322
rect 21440 3282 21452 3316
rect 21636 3282 21648 3316
rect 21440 3276 21648 3282
rect 17614 3202 17634 3232
rect 17628 3076 17634 3202
rect 15420 2616 15532 2698
rect 17622 3056 17634 3076
rect 17668 3076 17674 3232
rect 18086 3232 18132 3244
rect 18086 3084 18092 3232
rect 17668 3056 17682 3076
rect 17622 2616 17682 3056
rect 18078 3056 18092 3084
rect 18126 3084 18132 3232
rect 18544 3232 18590 3244
rect 18126 3056 18138 3084
rect 17776 3006 17984 3012
rect 17776 2972 17788 3006
rect 17972 2972 17984 3006
rect 17776 2966 17984 2972
rect 17850 2616 17910 2966
rect 18078 2768 18138 3056
rect 18544 3056 18550 3232
rect 18584 3056 18590 3232
rect 18544 3044 18590 3056
rect 19002 3232 19048 3244
rect 19002 3056 19008 3232
rect 19042 3056 19048 3232
rect 19002 3044 19048 3056
rect 19460 3232 19506 3244
rect 19460 3056 19466 3232
rect 19500 3056 19506 3232
rect 19460 3044 19506 3056
rect 19918 3232 19964 3244
rect 19918 3056 19924 3232
rect 19958 3056 19964 3232
rect 19918 3044 19964 3056
rect 20376 3232 20422 3244
rect 20376 3056 20382 3232
rect 20416 3056 20422 3232
rect 20376 3044 20422 3056
rect 20834 3232 20880 3244
rect 20834 3056 20840 3232
rect 20874 3056 20880 3232
rect 20834 3044 20880 3056
rect 21292 3232 21338 3244
rect 21292 3056 21298 3232
rect 21332 3056 21338 3232
rect 21742 3232 21802 3612
rect 21968 3322 22028 3612
rect 21898 3316 22106 3322
rect 21898 3282 21910 3316
rect 22094 3282 22106 3316
rect 21898 3276 22106 3282
rect 21742 3204 21756 3232
rect 21750 3076 21756 3204
rect 21292 3044 21338 3056
rect 21748 3056 21756 3076
rect 21790 3204 21802 3232
rect 22208 3232 22268 3612
rect 21790 3076 21796 3204
rect 21790 3056 21808 3076
rect 18234 3006 18442 3012
rect 18234 2972 18246 3006
rect 18430 2972 18442 3006
rect 18234 2966 18442 2972
rect 18692 3006 18900 3012
rect 18692 2972 18704 3006
rect 18888 2972 18900 3006
rect 18692 2966 18900 2972
rect 19150 3006 19358 3012
rect 19150 2972 19162 3006
rect 19346 2972 19358 3006
rect 19150 2966 19358 2972
rect 19608 3006 19816 3012
rect 19608 2972 19620 3006
rect 19804 2972 19816 3006
rect 19608 2966 19816 2972
rect 20066 3006 20274 3012
rect 20066 2972 20078 3006
rect 20262 2972 20274 3006
rect 20066 2966 20274 2972
rect 20524 3006 20732 3012
rect 20524 2972 20536 3006
rect 20720 2972 20732 3006
rect 20524 2966 20732 2972
rect 20982 3006 21190 3012
rect 20982 2972 20994 3006
rect 21178 2972 21190 3006
rect 20982 2966 21190 2972
rect 21440 3006 21648 3012
rect 21440 2972 21452 3006
rect 21636 2972 21648 3006
rect 21440 2966 21648 2972
rect 18310 2894 18376 2966
rect 18772 2894 18838 2966
rect 19226 2894 19292 2966
rect 19688 2894 19754 2966
rect 20142 2894 20208 2966
rect 20592 2894 20658 2966
rect 21058 2894 21124 2966
rect 21514 2894 21580 2966
rect 18310 2828 21580 2894
rect 18078 2702 18138 2708
rect 21748 2616 21808 3056
rect 22208 3056 22214 3232
rect 22248 3056 22268 3232
rect 21898 3006 22106 3012
rect 21898 2972 21910 3006
rect 22094 2972 22106 3006
rect 21898 2966 22106 2972
rect 21976 2616 22036 2966
rect 22208 2616 22268 3056
rect 24344 2698 24350 4122
rect 24450 2698 24456 4122
rect 24344 2616 24456 2698
rect 15420 2610 24456 2616
rect 15420 2510 15526 2610
rect 24350 2510 24456 2610
rect 15420 2504 24456 2510
rect 26002 4310 31458 4316
rect 26002 4210 26108 4310
rect 31352 4210 31458 4310
rect 26002 4204 31458 4210
rect 26002 4126 26114 4204
rect 26002 2614 26008 4126
rect 26108 2614 26114 4126
rect 26714 3904 26724 4204
rect 30736 3904 30746 4204
rect 31346 4126 31458 4204
rect 26312 3726 31284 3756
rect 26312 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 31284 3726
rect 26312 3612 31284 3640
rect 26376 3232 26436 3612
rect 26616 3322 26676 3612
rect 26538 3316 26746 3322
rect 26538 3282 26550 3316
rect 26734 3282 26746 3316
rect 26538 3276 26746 3282
rect 26376 3202 26396 3232
rect 26390 3076 26396 3202
rect 26002 2536 26114 2614
rect 26384 3056 26396 3076
rect 26430 3076 26436 3232
rect 26840 3232 26900 3612
rect 27066 3388 30330 3448
rect 27066 3322 27126 3388
rect 27528 3322 27588 3388
rect 27982 3322 28042 3388
rect 28444 3322 28504 3388
rect 28898 3322 28958 3388
rect 29348 3322 29408 3388
rect 29814 3322 29874 3388
rect 30270 3322 30330 3388
rect 30730 3322 30790 3612
rect 26996 3316 27204 3322
rect 26996 3282 27008 3316
rect 27192 3282 27204 3316
rect 26996 3276 27204 3282
rect 27454 3316 27662 3322
rect 27454 3282 27466 3316
rect 27650 3282 27662 3316
rect 27454 3276 27662 3282
rect 27912 3316 28120 3322
rect 27912 3282 27924 3316
rect 28108 3282 28120 3316
rect 27912 3276 28120 3282
rect 28370 3316 28578 3322
rect 28370 3282 28382 3316
rect 28566 3282 28578 3316
rect 28370 3276 28578 3282
rect 28828 3316 29036 3322
rect 28828 3282 28840 3316
rect 29024 3282 29036 3316
rect 28828 3276 29036 3282
rect 29286 3316 29494 3322
rect 29286 3282 29298 3316
rect 29482 3282 29494 3316
rect 29286 3276 29494 3282
rect 29744 3316 29952 3322
rect 29744 3282 29756 3316
rect 29940 3282 29952 3316
rect 29744 3276 29952 3282
rect 30202 3316 30410 3322
rect 30202 3282 30214 3316
rect 30398 3282 30410 3316
rect 30202 3276 30410 3282
rect 30660 3316 30868 3322
rect 30660 3282 30672 3316
rect 30856 3282 30868 3316
rect 30660 3276 30868 3282
rect 26430 3056 26444 3076
rect 26384 2536 26444 3056
rect 26840 3056 26854 3232
rect 26888 3056 26900 3232
rect 26538 3006 26746 3012
rect 26538 2972 26550 3006
rect 26734 2972 26746 3006
rect 26538 2966 26746 2972
rect 26612 2536 26672 2966
rect 26840 2536 26900 3056
rect 27306 3232 27352 3244
rect 27306 3056 27312 3232
rect 27346 3056 27352 3232
rect 27306 3044 27352 3056
rect 27764 3232 27810 3244
rect 27764 3056 27770 3232
rect 27804 3056 27810 3232
rect 27764 3044 27810 3056
rect 28222 3232 28268 3244
rect 28222 3056 28228 3232
rect 28262 3056 28268 3232
rect 28222 3044 28268 3056
rect 28680 3232 28726 3244
rect 28680 3056 28686 3232
rect 28720 3056 28726 3232
rect 28680 3044 28726 3056
rect 29138 3232 29184 3244
rect 29138 3056 29144 3232
rect 29178 3056 29184 3232
rect 29138 3044 29184 3056
rect 29596 3232 29642 3244
rect 29596 3056 29602 3232
rect 29636 3056 29642 3232
rect 29596 3044 29642 3056
rect 30054 3232 30100 3244
rect 30054 3056 30060 3232
rect 30094 3056 30100 3232
rect 30512 3232 30558 3244
rect 30512 3110 30518 3232
rect 30054 3044 30100 3056
rect 30504 3056 30518 3110
rect 30552 3110 30558 3232
rect 30970 3232 31030 3612
rect 30552 3056 30564 3110
rect 26996 3006 27204 3012
rect 26996 2972 27008 3006
rect 27192 2972 27204 3006
rect 26996 2966 27204 2972
rect 27454 3006 27662 3012
rect 27454 2972 27466 3006
rect 27650 2972 27662 3006
rect 27454 2966 27662 2972
rect 27912 3006 28120 3012
rect 27912 2972 27924 3006
rect 28108 2972 28120 3006
rect 27912 2966 28120 2972
rect 28370 3006 28578 3012
rect 28370 2972 28382 3006
rect 28566 2972 28578 3006
rect 28370 2966 28578 2972
rect 28828 3006 29036 3012
rect 28828 2972 28840 3006
rect 29024 2972 29036 3006
rect 28828 2966 29036 2972
rect 29286 3006 29494 3012
rect 29286 2972 29298 3006
rect 29482 2972 29494 3006
rect 29286 2966 29494 2972
rect 29744 3006 29952 3012
rect 29744 2972 29756 3006
rect 29940 2972 29952 3006
rect 29744 2966 29952 2972
rect 30202 3006 30410 3012
rect 30202 2972 30214 3006
rect 30398 2972 30410 3006
rect 30202 2966 30410 2972
rect 27066 2894 27126 2966
rect 27528 2894 27588 2966
rect 27982 2896 28042 2966
rect 27976 2894 27982 2896
rect 27059 2834 27066 2894
rect 27126 2834 27528 2894
rect 27588 2836 27982 2894
rect 28042 2894 28048 2896
rect 28444 2894 28504 2966
rect 28898 2894 28958 2966
rect 29348 2894 29408 2966
rect 29814 2894 29874 2966
rect 30270 2894 30330 2966
rect 28042 2836 28444 2894
rect 27588 2834 28444 2836
rect 28504 2834 28898 2894
rect 28958 2834 29348 2894
rect 29408 2834 29814 2894
rect 29874 2834 30270 2894
rect 30330 2834 30337 2894
rect 27059 2828 30337 2834
rect 30504 2686 30564 3056
rect 30970 3056 30976 3232
rect 31010 3056 31030 3232
rect 30660 3006 30868 3012
rect 30660 2972 30672 3006
rect 30856 2972 30868 3006
rect 30660 2966 30868 2972
rect 30498 2626 30504 2686
rect 30564 2626 30570 2686
rect 30738 2536 30798 2966
rect 30970 2536 31030 3056
rect 31346 2614 31352 4126
rect 31452 2614 31458 4126
rect 31346 2538 31458 2614
rect 31346 2536 32278 2538
rect 26002 2530 32278 2536
rect 26002 2430 26108 2530
rect 31352 2507 32278 2530
rect 31352 2473 31571 2507
rect 31605 2473 31663 2507
rect 31697 2473 31755 2507
rect 31789 2473 31847 2507
rect 31881 2473 31939 2507
rect 31973 2473 32031 2507
rect 32065 2473 32123 2507
rect 32157 2473 32215 2507
rect 32249 2473 32278 2507
rect 31352 2442 32278 2473
rect 31352 2430 31458 2442
rect 26002 2424 31458 2430
rect 30504 2344 30564 2350
rect 25234 2284 30504 2344
rect 30564 2284 31566 2344
rect 15420 2274 24456 2280
rect 15420 2174 15526 2274
rect 24350 2174 24456 2274
rect 15420 2168 24456 2174
rect 15420 1976 15532 2168
rect 15420 -996 15426 1976
rect 15036 -1056 15426 -996
rect 15420 -1360 15426 -1056
rect 15526 1614 15532 1976
rect 15790 1614 15850 2168
rect 16018 1614 16078 2168
rect 16244 1614 16304 2168
rect 16702 2026 23178 2086
rect 15526 1554 16304 1614
rect 16468 1554 16474 1614
rect 16534 1554 16540 1614
rect 15526 -996 15532 1554
rect 15790 1381 15850 1554
rect 16018 1480 16078 1554
rect 15944 1474 16152 1480
rect 15944 1440 15956 1474
rect 16140 1440 16152 1474
rect 15944 1434 16152 1440
rect 15790 1322 15802 1381
rect 15796 -162 15802 1322
rect 15788 -195 15802 -162
rect 15836 1322 15850 1381
rect 16244 1381 16304 1554
rect 16474 1480 16534 1554
rect 16402 1474 16610 1480
rect 16402 1440 16414 1474
rect 16598 1440 16610 1474
rect 16402 1434 16610 1440
rect 16244 1338 16260 1381
rect 15836 -162 15842 1322
rect 16254 -130 16260 1338
rect 15836 -195 15848 -162
rect 15788 -982 15848 -195
rect 16246 -195 16260 -130
rect 16294 1338 16304 1381
rect 16702 1381 16762 2026
rect 17620 1902 22264 1962
rect 16924 1554 16930 1614
rect 16990 1554 16996 1614
rect 17384 1554 17390 1614
rect 17450 1554 17456 1614
rect 16930 1480 16990 1554
rect 17390 1480 17450 1554
rect 16860 1474 17068 1480
rect 16860 1440 16872 1474
rect 17056 1440 17068 1474
rect 16860 1434 17068 1440
rect 17318 1474 17526 1480
rect 17318 1440 17330 1474
rect 17514 1440 17526 1474
rect 17318 1434 17526 1440
rect 16294 -130 16300 1338
rect 16702 1298 16718 1381
rect 16294 -195 16306 -130
rect 15944 -254 16152 -248
rect 15944 -288 15956 -254
rect 16140 -288 16152 -254
rect 15944 -294 16152 -288
rect 16020 -982 16080 -294
rect 16246 -982 16306 -195
rect 16712 -195 16718 1298
rect 16752 1298 16762 1381
rect 17170 1381 17216 1393
rect 16752 -195 16758 1298
rect 17170 -136 17176 1381
rect 16712 -207 16758 -195
rect 17162 -195 17176 -136
rect 17210 -136 17216 1381
rect 17620 1381 17680 1902
rect 18528 1778 21344 1838
rect 17840 1554 17846 1614
rect 17906 1554 17912 1614
rect 18298 1554 18304 1614
rect 18364 1554 18370 1614
rect 17846 1480 17906 1554
rect 18304 1480 18364 1554
rect 17776 1474 17984 1480
rect 17776 1440 17788 1474
rect 17972 1440 17984 1474
rect 17776 1434 17984 1440
rect 18234 1474 18442 1480
rect 18234 1440 18246 1474
rect 18430 1440 18442 1474
rect 18234 1434 18442 1440
rect 18528 1393 18588 1778
rect 19452 1662 20430 1722
rect 18762 1554 18768 1614
rect 18828 1554 18834 1614
rect 19216 1554 19222 1614
rect 19282 1554 19288 1614
rect 18768 1480 18828 1554
rect 19222 1480 19282 1554
rect 18692 1474 18900 1480
rect 18692 1440 18704 1474
rect 18888 1440 18900 1474
rect 18692 1434 18900 1440
rect 19150 1474 19358 1480
rect 19150 1440 19162 1474
rect 19346 1440 19358 1474
rect 19150 1434 19358 1440
rect 17620 1304 17634 1381
rect 17210 -195 17222 -136
rect 16402 -254 16610 -248
rect 16402 -288 16414 -254
rect 16598 -288 16610 -254
rect 16402 -294 16610 -288
rect 16860 -254 17068 -248
rect 16860 -288 16872 -254
rect 17056 -288 17068 -254
rect 16860 -294 17068 -288
rect 16478 -360 16538 -294
rect 16934 -360 16994 -294
rect 16472 -420 16478 -360
rect 16538 -420 16544 -360
rect 16928 -420 16934 -360
rect 16994 -420 17000 -360
rect 17162 -728 17222 -195
rect 17628 -195 17634 1304
rect 17668 1304 17680 1381
rect 18086 1381 18132 1393
rect 17668 -195 17674 1304
rect 18086 -134 18092 1381
rect 17628 -207 17674 -195
rect 18078 -195 18092 -134
rect 18126 -134 18132 1381
rect 18528 1381 18590 1393
rect 18528 1310 18550 1381
rect 18126 -195 18138 -134
rect 17318 -254 17526 -248
rect 17318 -288 17330 -254
rect 17514 -288 17526 -254
rect 17318 -294 17526 -288
rect 17776 -254 17984 -248
rect 17776 -288 17788 -254
rect 17972 -288 17984 -254
rect 17776 -294 17984 -288
rect 17394 -360 17454 -294
rect 17850 -360 17910 -294
rect 17388 -420 17394 -360
rect 17454 -420 17460 -360
rect 17844 -420 17850 -360
rect 17910 -420 17916 -360
rect 18078 -594 18138 -195
rect 18544 -195 18550 1310
rect 18584 -195 18590 1381
rect 19002 1381 19048 1393
rect 19002 -116 19008 1381
rect 18544 -207 18590 -195
rect 18994 -195 19008 -116
rect 19042 -116 19048 1381
rect 19452 1381 19512 1662
rect 19676 1554 19682 1614
rect 19742 1554 19748 1614
rect 19906 1554 19912 1614
rect 19972 1554 19978 1614
rect 20134 1554 20140 1614
rect 20200 1554 20206 1614
rect 19682 1480 19742 1554
rect 19608 1474 19816 1480
rect 19608 1440 19620 1474
rect 19804 1440 19816 1474
rect 19608 1434 19816 1440
rect 19452 1302 19466 1381
rect 19042 -195 19054 -116
rect 18234 -254 18442 -248
rect 18234 -288 18246 -254
rect 18430 -288 18442 -254
rect 18234 -294 18442 -288
rect 18692 -254 18900 -248
rect 18692 -288 18704 -254
rect 18888 -288 18900 -254
rect 18692 -294 18900 -288
rect 18308 -360 18368 -294
rect 18772 -360 18832 -294
rect 18302 -420 18308 -360
rect 18368 -420 18374 -360
rect 18766 -420 18772 -360
rect 18832 -420 18838 -360
rect 18994 -470 19054 -195
rect 19460 -195 19466 1302
rect 19500 1302 19512 1381
rect 19912 1381 19972 1554
rect 20140 1480 20200 1554
rect 20066 1474 20274 1480
rect 20066 1440 20078 1474
rect 20262 1440 20274 1474
rect 20066 1434 20274 1440
rect 19912 1332 19924 1381
rect 19500 -195 19506 1302
rect 19460 -207 19506 -195
rect 19918 -195 19924 1332
rect 19958 1332 19972 1381
rect 20370 1381 20430 1662
rect 20590 1554 20596 1614
rect 20656 1554 20662 1614
rect 21050 1554 21056 1614
rect 21116 1554 21122 1614
rect 20596 1480 20656 1554
rect 21056 1480 21116 1554
rect 20524 1474 20732 1480
rect 20524 1440 20536 1474
rect 20720 1440 20732 1474
rect 20524 1434 20732 1440
rect 20982 1474 21190 1480
rect 20982 1440 20994 1474
rect 21178 1440 21190 1474
rect 20982 1434 21190 1440
rect 20370 1354 20382 1381
rect 19958 -195 19964 1332
rect 19918 -207 19964 -195
rect 20376 -195 20382 1354
rect 20416 1354 20430 1381
rect 20834 1381 20880 1393
rect 20416 -195 20422 1354
rect 20834 -150 20840 1381
rect 20376 -207 20422 -195
rect 20824 -195 20840 -150
rect 20874 -150 20880 1381
rect 21284 1381 21344 1778
rect 21506 1554 21512 1614
rect 21572 1554 21578 1614
rect 21962 1554 21968 1614
rect 22028 1554 22034 1614
rect 21512 1480 21572 1554
rect 21968 1480 22028 1554
rect 21440 1474 21648 1480
rect 21440 1440 21452 1474
rect 21636 1440 21648 1474
rect 21440 1434 21648 1440
rect 21898 1474 22106 1480
rect 21898 1440 21910 1474
rect 22094 1440 22106 1474
rect 21898 1434 22106 1440
rect 21284 1350 21298 1381
rect 20874 -195 20884 -150
rect 19150 -254 19358 -248
rect 19150 -288 19162 -254
rect 19346 -288 19358 -254
rect 19150 -294 19358 -288
rect 19608 -254 19816 -248
rect 19608 -288 19620 -254
rect 19804 -288 19816 -254
rect 19608 -294 19816 -288
rect 20066 -254 20274 -248
rect 20066 -288 20078 -254
rect 20262 -288 20274 -254
rect 20066 -294 20274 -288
rect 20524 -254 20732 -248
rect 20524 -288 20536 -254
rect 20720 -288 20732 -254
rect 20524 -294 20732 -288
rect 19222 -360 19282 -294
rect 19678 -360 19738 -294
rect 20146 -360 20206 -294
rect 20604 -360 20664 -294
rect 19216 -420 19222 -360
rect 19282 -420 19288 -360
rect 19672 -420 19678 -360
rect 19738 -420 19744 -360
rect 20140 -420 20146 -360
rect 20206 -420 20212 -360
rect 20598 -420 20604 -360
rect 20664 -420 20670 -360
rect 20824 -470 20884 -195
rect 21292 -195 21298 1350
rect 21332 1350 21344 1381
rect 21750 1381 21796 1393
rect 21332 -195 21338 1350
rect 21750 -136 21756 1381
rect 21292 -207 21338 -195
rect 21740 -195 21756 -136
rect 21790 -136 21796 1381
rect 22204 1381 22264 1902
rect 22418 1554 22424 1614
rect 22484 1554 22490 1614
rect 22876 1554 22882 1614
rect 22942 1554 22948 1614
rect 22424 1480 22484 1554
rect 22882 1480 22942 1554
rect 22356 1474 22564 1480
rect 22356 1440 22368 1474
rect 22552 1440 22564 1474
rect 22356 1434 22564 1440
rect 22814 1474 23022 1480
rect 22814 1440 22826 1474
rect 23010 1440 23022 1474
rect 22814 1434 23022 1440
rect 22204 1314 22214 1381
rect 21790 -195 21800 -136
rect 20982 -254 21190 -248
rect 20982 -288 20994 -254
rect 21178 -288 21190 -254
rect 20982 -294 21190 -288
rect 21440 -254 21648 -248
rect 21440 -288 21452 -254
rect 21636 -288 21648 -254
rect 21440 -294 21648 -288
rect 21060 -360 21120 -294
rect 21516 -360 21576 -294
rect 21054 -420 21060 -360
rect 21120 -420 21126 -360
rect 21510 -420 21516 -360
rect 21576 -420 21582 -360
rect 18994 -530 20884 -470
rect 21740 -594 21800 -195
rect 22208 -195 22214 1314
rect 22248 1314 22264 1381
rect 22666 1381 22712 1393
rect 22248 -195 22254 1314
rect 22666 -138 22672 1381
rect 22208 -207 22254 -195
rect 22660 -195 22672 -138
rect 22706 -138 22712 1381
rect 23118 1381 23178 2026
rect 23572 1614 23632 2168
rect 23804 1614 23864 2168
rect 24030 1614 24090 2168
rect 24344 1976 24456 2168
rect 24344 1614 24350 1976
rect 23336 1554 23342 1614
rect 23402 1554 23408 1614
rect 23572 1554 24350 1614
rect 23342 1480 23402 1554
rect 23272 1474 23480 1480
rect 23272 1440 23284 1474
rect 23468 1440 23480 1474
rect 23272 1434 23480 1440
rect 23118 1322 23130 1381
rect 22706 -195 22720 -138
rect 21898 -254 22106 -248
rect 21898 -288 21910 -254
rect 22094 -288 22106 -254
rect 21898 -294 22106 -288
rect 22356 -254 22564 -248
rect 22356 -288 22368 -254
rect 22552 -288 22564 -254
rect 22356 -294 22564 -288
rect 21972 -360 22032 -294
rect 22428 -360 22488 -294
rect 21966 -420 21972 -360
rect 22032 -420 22038 -360
rect 22422 -420 22428 -360
rect 22488 -420 22494 -360
rect 18078 -654 21800 -594
rect 22660 -728 22720 -195
rect 23124 -195 23130 1322
rect 23164 1322 23178 1381
rect 23572 1381 23632 1554
rect 23804 1480 23864 1554
rect 23730 1474 23938 1480
rect 23730 1440 23742 1474
rect 23926 1440 23938 1474
rect 23730 1434 23938 1440
rect 23164 -195 23170 1322
rect 23572 1320 23588 1381
rect 23582 -118 23588 1320
rect 23124 -207 23170 -195
rect 23576 -195 23588 -118
rect 23622 1320 23632 1381
rect 24030 1381 24090 1554
rect 24030 1338 24046 1381
rect 23622 -118 23628 1320
rect 23622 -195 23636 -118
rect 24040 -124 24046 1338
rect 22814 -254 23022 -248
rect 22814 -288 22826 -254
rect 23010 -288 23022 -254
rect 22814 -294 23022 -288
rect 23272 -254 23480 -248
rect 23272 -288 23284 -254
rect 23468 -288 23480 -254
rect 23272 -294 23480 -288
rect 22886 -360 22946 -294
rect 23346 -360 23406 -294
rect 22880 -420 22886 -360
rect 22946 -420 22952 -360
rect 23340 -420 23346 -360
rect 23406 -420 23412 -360
rect 17162 -788 22720 -728
rect 23576 -982 23636 -195
rect 24034 -195 24046 -124
rect 24080 1338 24090 1381
rect 24080 -124 24086 1338
rect 24080 -195 24094 -124
rect 23730 -254 23938 -248
rect 23730 -288 23742 -254
rect 23926 -288 23938 -254
rect 23730 -294 23938 -288
rect 23806 -982 23866 -294
rect 24034 -982 24094 -195
rect 24344 -982 24350 1554
rect 15760 -992 24350 -982
rect 15760 -996 15774 -992
rect 15526 -1056 15774 -996
rect 15526 -1360 15532 -1056
rect 15760 -1078 15774 -1056
rect 15870 -1078 16374 -992
rect 16470 -1078 16974 -992
rect 17070 -1078 17574 -992
rect 17670 -1078 18174 -992
rect 18270 -1078 18774 -992
rect 18870 -1078 19374 -992
rect 19470 -1078 19974 -992
rect 20070 -1078 20574 -992
rect 20670 -1078 21174 -992
rect 21270 -1078 21774 -992
rect 21870 -1078 22374 -992
rect 22470 -1078 22974 -992
rect 23070 -1078 23574 -992
rect 23670 -1078 23994 -992
rect 24090 -1078 24350 -992
rect 15760 -1092 24350 -1078
rect 15420 -1552 15532 -1360
rect 15914 -1552 15924 -1252
rect 23656 -1552 23666 -1252
rect 24344 -1360 24350 -1092
rect 24450 -982 24456 1976
rect 24450 -1092 24458 -982
rect 24450 -1360 24456 -1092
rect 24344 -1552 24456 -1360
rect 15420 -1558 24456 -1552
rect 15420 -1658 15526 -1558
rect 24350 -1658 24456 -1558
rect 15420 -1664 24456 -1658
rect 10812 -2028 21268 -2022
rect 10812 -2128 10918 -2028
rect 21162 -2128 21268 -2028
rect 10812 -2134 21268 -2128
rect 10812 -2418 10924 -2134
rect 10812 -7590 10818 -2418
rect 10918 -5240 10924 -2418
rect 11524 -2434 11534 -2134
rect 20546 -2434 20556 -2134
rect 21156 -2418 21268 -2134
rect 11762 -2608 20118 -2594
rect 11762 -2694 11776 -2608
rect 11872 -2694 12376 -2608
rect 12472 -2694 12976 -2608
rect 13072 -2694 13576 -2608
rect 13672 -2694 14176 -2608
rect 14272 -2694 14776 -2608
rect 14872 -2694 15376 -2608
rect 15472 -2694 15976 -2608
rect 16072 -2694 16576 -2608
rect 16672 -2694 17176 -2608
rect 17272 -2694 17776 -2608
rect 17872 -2694 18376 -2608
rect 18472 -2694 18976 -2608
rect 19072 -2694 19576 -2608
rect 19672 -2694 19996 -2608
rect 20092 -2694 20118 -2608
rect 11762 -2704 20118 -2694
rect 11790 -3492 11850 -2704
rect 12022 -3393 12082 -2704
rect 11946 -3399 12154 -3393
rect 11946 -3433 11958 -3399
rect 12142 -3433 12154 -3399
rect 11946 -3439 12154 -3433
rect 11790 -3524 11804 -3492
rect 11798 -5008 11804 -3524
rect 11792 -5068 11804 -5008
rect 11838 -3524 11850 -3492
rect 12248 -3492 12308 -2704
rect 13164 -2958 18722 -2898
rect 12474 -3326 12480 -3266
rect 12540 -3326 12546 -3266
rect 12930 -3326 12936 -3266
rect 12996 -3326 13002 -3266
rect 12480 -3393 12540 -3326
rect 12936 -3393 12996 -3326
rect 12404 -3399 12612 -3393
rect 12404 -3433 12416 -3399
rect 12600 -3433 12612 -3399
rect 12404 -3439 12612 -3433
rect 12862 -3399 13070 -3393
rect 12862 -3433 12874 -3399
rect 13058 -3433 13070 -3399
rect 12862 -3439 13070 -3433
rect 11838 -5008 11844 -3524
rect 12248 -3556 12262 -3492
rect 11838 -5068 11852 -5008
rect 12256 -5024 12262 -3556
rect 11792 -5240 11852 -5068
rect 12246 -5068 12262 -5024
rect 12296 -3556 12308 -3492
rect 12714 -3492 12760 -3480
rect 12296 -5024 12302 -3556
rect 12714 -4984 12720 -3492
rect 12296 -5068 12306 -5024
rect 11946 -5127 12154 -5121
rect 11946 -5161 11958 -5127
rect 12142 -5161 12154 -5127
rect 11946 -5167 12154 -5161
rect 12020 -5240 12080 -5167
rect 12246 -5240 12306 -5068
rect 12704 -5068 12720 -4984
rect 12754 -4984 12760 -3492
rect 13164 -3492 13224 -2958
rect 14080 -3092 17802 -3032
rect 13390 -3326 13396 -3266
rect 13456 -3326 13462 -3266
rect 13846 -3326 13852 -3266
rect 13912 -3326 13918 -3266
rect 13396 -3393 13456 -3326
rect 13852 -3393 13912 -3326
rect 13320 -3399 13528 -3393
rect 13320 -3433 13332 -3399
rect 13516 -3433 13528 -3399
rect 13320 -3439 13528 -3433
rect 13778 -3399 13986 -3393
rect 13778 -3433 13790 -3399
rect 13974 -3433 13986 -3399
rect 13778 -3439 13986 -3433
rect 13164 -3550 13178 -3492
rect 12754 -5068 12764 -4984
rect 12404 -5127 12612 -5121
rect 12404 -5161 12416 -5127
rect 12600 -5161 12612 -5127
rect 12404 -5167 12612 -5161
rect 12476 -5240 12536 -5167
rect 10918 -5300 12306 -5240
rect 12470 -5300 12476 -5240
rect 12536 -5300 12542 -5240
rect 10918 -5672 10924 -5300
rect 11792 -5672 11852 -5300
rect 10918 -5732 11852 -5672
rect 12704 -5720 12764 -5068
rect 13172 -5068 13178 -3550
rect 13212 -3550 13224 -3492
rect 13630 -3492 13676 -3480
rect 13212 -5068 13218 -3550
rect 13630 -4990 13636 -3492
rect 13172 -5080 13218 -5068
rect 13622 -5068 13636 -4990
rect 13670 -4990 13676 -3492
rect 14080 -3492 14140 -3092
rect 14996 -3216 16886 -3156
rect 14304 -3326 14310 -3266
rect 14370 -3326 14376 -3266
rect 14768 -3326 14774 -3266
rect 14834 -3326 14840 -3266
rect 14310 -3393 14370 -3326
rect 14774 -3393 14834 -3326
rect 14236 -3399 14444 -3393
rect 14236 -3433 14248 -3399
rect 14432 -3433 14444 -3399
rect 14236 -3439 14444 -3433
rect 14694 -3399 14902 -3393
rect 14694 -3433 14706 -3399
rect 14890 -3433 14902 -3399
rect 14694 -3439 14902 -3433
rect 14080 -3552 14094 -3492
rect 13670 -5068 13682 -4990
rect 12862 -5127 13070 -5121
rect 12862 -5161 12874 -5127
rect 13058 -5161 13070 -5127
rect 12862 -5167 13070 -5161
rect 13320 -5127 13528 -5121
rect 13320 -5161 13332 -5127
rect 13516 -5161 13528 -5127
rect 13320 -5167 13528 -5161
rect 12932 -5240 12992 -5167
rect 13392 -5240 13452 -5167
rect 12926 -5300 12932 -5240
rect 12992 -5300 12998 -5240
rect 13386 -5300 13392 -5240
rect 13452 -5300 13458 -5240
rect 13622 -5590 13682 -5068
rect 14088 -5068 14094 -3552
rect 14128 -3552 14140 -3492
rect 14546 -3492 14592 -3480
rect 14128 -5068 14134 -3552
rect 14546 -4996 14552 -3492
rect 14088 -5080 14134 -5068
rect 14530 -5068 14552 -4996
rect 14586 -5068 14592 -3492
rect 14996 -3492 15056 -3216
rect 15218 -3326 15224 -3266
rect 15284 -3326 15290 -3266
rect 15674 -3326 15680 -3266
rect 15740 -3326 15746 -3266
rect 16142 -3326 16148 -3266
rect 16208 -3326 16214 -3266
rect 16600 -3326 16606 -3266
rect 16666 -3326 16672 -3266
rect 15224 -3393 15284 -3326
rect 15680 -3393 15740 -3326
rect 16148 -3393 16208 -3326
rect 16606 -3393 16666 -3326
rect 15152 -3399 15360 -3393
rect 15152 -3433 15164 -3399
rect 15348 -3433 15360 -3399
rect 15152 -3439 15360 -3433
rect 15610 -3399 15818 -3393
rect 15610 -3433 15622 -3399
rect 15806 -3433 15818 -3399
rect 15610 -3439 15818 -3433
rect 16068 -3399 16276 -3393
rect 16068 -3433 16080 -3399
rect 16264 -3433 16276 -3399
rect 16068 -3439 16276 -3433
rect 16526 -3399 16734 -3393
rect 16526 -3433 16538 -3399
rect 16722 -3433 16734 -3399
rect 16526 -3439 16734 -3433
rect 14996 -3570 15010 -3492
rect 14530 -5080 14592 -5068
rect 15004 -5068 15010 -3570
rect 15044 -3570 15056 -3492
rect 15462 -3492 15508 -3480
rect 15044 -5068 15050 -3570
rect 15462 -4988 15468 -3492
rect 15004 -5080 15050 -5068
rect 15454 -5068 15468 -4988
rect 15502 -4988 15508 -3492
rect 15920 -3492 15966 -3480
rect 15502 -5068 15514 -4988
rect 15920 -5046 15926 -3492
rect 13778 -5127 13986 -5121
rect 13778 -5161 13790 -5127
rect 13974 -5161 13986 -5127
rect 13778 -5167 13986 -5161
rect 14236 -5127 14444 -5121
rect 14236 -5161 14248 -5127
rect 14432 -5161 14444 -5127
rect 14236 -5167 14444 -5161
rect 13848 -5240 13908 -5167
rect 14306 -5240 14366 -5167
rect 13842 -5300 13848 -5240
rect 13908 -5300 13914 -5240
rect 14300 -5300 14306 -5240
rect 14366 -5300 14372 -5240
rect 14530 -5464 14590 -5080
rect 14694 -5127 14902 -5121
rect 14694 -5161 14706 -5127
rect 14890 -5161 14902 -5127
rect 14694 -5167 14902 -5161
rect 15152 -5127 15360 -5121
rect 15152 -5161 15164 -5127
rect 15348 -5161 15360 -5127
rect 15152 -5167 15360 -5161
rect 14770 -5240 14830 -5167
rect 15224 -5240 15284 -5167
rect 14764 -5300 14770 -5240
rect 14830 -5300 14836 -5240
rect 15218 -5300 15224 -5240
rect 15284 -5300 15290 -5240
rect 15454 -5348 15514 -5068
rect 15916 -5068 15926 -5046
rect 15960 -5046 15966 -3492
rect 16378 -3492 16424 -3480
rect 16378 -5040 16384 -3492
rect 15960 -5068 15976 -5046
rect 15610 -5127 15818 -5121
rect 15610 -5161 15622 -5127
rect 15806 -5161 15818 -5127
rect 15610 -5167 15818 -5161
rect 15682 -5238 15742 -5167
rect 15916 -5228 15976 -5068
rect 16372 -5068 16384 -5040
rect 16418 -5040 16424 -3492
rect 16826 -3492 16886 -3216
rect 17056 -3326 17062 -3266
rect 17122 -3326 17128 -3266
rect 17512 -3326 17518 -3266
rect 17578 -3326 17584 -3266
rect 17062 -3393 17122 -3326
rect 17518 -3393 17578 -3326
rect 16984 -3399 17192 -3393
rect 16984 -3433 16996 -3399
rect 17180 -3433 17192 -3399
rect 16984 -3439 17192 -3433
rect 17442 -3399 17650 -3393
rect 17442 -3433 17454 -3399
rect 17638 -3433 17650 -3399
rect 17442 -3439 17650 -3433
rect 16826 -3536 16842 -3492
rect 16418 -5068 16432 -5040
rect 16068 -5127 16276 -5121
rect 16068 -5161 16080 -5127
rect 16264 -5161 16276 -5127
rect 16068 -5167 16276 -5161
rect 15676 -5240 15748 -5238
rect 15676 -5300 15682 -5240
rect 15742 -5300 15748 -5240
rect 16142 -5232 16202 -5167
rect 15916 -5294 15976 -5288
rect 16130 -5238 16214 -5232
rect 16130 -5300 16142 -5238
rect 16202 -5300 16214 -5238
rect 16130 -5304 16214 -5300
rect 16372 -5348 16432 -5068
rect 16836 -5068 16842 -3536
rect 16876 -3536 16886 -3492
rect 17294 -3492 17340 -3480
rect 16876 -5068 16882 -3536
rect 17294 -5036 17300 -3492
rect 16836 -5080 16882 -5068
rect 17286 -5068 17300 -5036
rect 17334 -5036 17340 -3492
rect 17742 -3492 17802 -3092
rect 17968 -3326 17974 -3266
rect 18034 -3326 18040 -3266
rect 18424 -3326 18430 -3266
rect 18490 -3326 18496 -3266
rect 17974 -3393 18034 -3326
rect 18430 -3393 18490 -3326
rect 17900 -3399 18108 -3393
rect 17900 -3433 17912 -3399
rect 18096 -3433 18108 -3399
rect 17900 -3439 18108 -3433
rect 18358 -3399 18566 -3393
rect 18358 -3433 18370 -3399
rect 18554 -3433 18566 -3399
rect 18358 -3439 18566 -3433
rect 17742 -3550 17758 -3492
rect 17334 -5068 17346 -5036
rect 16526 -5127 16734 -5121
rect 16526 -5161 16538 -5127
rect 16722 -5161 16734 -5127
rect 16526 -5167 16734 -5161
rect 16984 -5127 17192 -5121
rect 16984 -5161 16996 -5127
rect 17180 -5161 17192 -5127
rect 16984 -5167 17192 -5161
rect 16598 -5240 16658 -5167
rect 17058 -5240 17118 -5167
rect 16592 -5300 16598 -5240
rect 16658 -5300 16664 -5240
rect 17052 -5300 17058 -5240
rect 17118 -5300 17124 -5240
rect 15454 -5408 16432 -5348
rect 17286 -5464 17346 -5068
rect 17752 -5068 17758 -3550
rect 17792 -3550 17802 -3492
rect 18210 -3492 18256 -3480
rect 17792 -5068 17798 -3550
rect 18210 -5000 18216 -3492
rect 17752 -5080 17798 -5068
rect 18206 -5068 18216 -5000
rect 18250 -5000 18256 -3492
rect 18662 -3492 18722 -2958
rect 18882 -3326 18888 -3266
rect 18948 -3326 18954 -3266
rect 19342 -3326 19348 -3266
rect 19408 -3326 19414 -3266
rect 18888 -3393 18948 -3326
rect 19348 -3393 19408 -3326
rect 18816 -3399 19024 -3393
rect 18816 -3433 18828 -3399
rect 19012 -3433 19024 -3399
rect 18816 -3439 19024 -3433
rect 19274 -3399 19482 -3393
rect 19274 -3433 19286 -3399
rect 19470 -3433 19482 -3399
rect 19274 -3439 19482 -3433
rect 18662 -3548 18674 -3492
rect 18250 -5068 18266 -5000
rect 17442 -5127 17650 -5121
rect 17442 -5161 17454 -5127
rect 17638 -5161 17650 -5127
rect 17442 -5167 17650 -5161
rect 17900 -5127 18108 -5121
rect 17900 -5161 17912 -5127
rect 18096 -5161 18108 -5127
rect 17900 -5167 18108 -5161
rect 17514 -5240 17574 -5167
rect 17970 -5240 18030 -5167
rect 17508 -5300 17514 -5240
rect 17574 -5300 17580 -5240
rect 17964 -5300 17970 -5240
rect 18030 -5300 18036 -5240
rect 14530 -5524 17346 -5464
rect 18206 -5590 18266 -5068
rect 18668 -5068 18674 -3548
rect 18708 -3548 18722 -3492
rect 19126 -3492 19172 -3480
rect 18708 -5068 18714 -3548
rect 19126 -5008 19132 -3492
rect 18668 -5080 18714 -5068
rect 19120 -5068 19132 -5008
rect 19166 -5008 19172 -3492
rect 19578 -3492 19638 -2704
rect 19808 -3393 19868 -2704
rect 19732 -3399 19940 -3393
rect 19732 -3433 19744 -3399
rect 19928 -3433 19940 -3399
rect 19732 -3439 19940 -3433
rect 19578 -3568 19590 -3492
rect 19584 -5006 19590 -3568
rect 19166 -5068 19180 -5008
rect 18358 -5127 18566 -5121
rect 18358 -5161 18370 -5127
rect 18554 -5161 18566 -5127
rect 18358 -5167 18566 -5161
rect 18816 -5127 19024 -5121
rect 18816 -5161 18828 -5127
rect 19012 -5161 19024 -5127
rect 18816 -5167 19024 -5161
rect 18426 -5240 18486 -5167
rect 18884 -5240 18944 -5167
rect 18420 -5300 18426 -5240
rect 18486 -5300 18492 -5240
rect 18878 -5300 18884 -5240
rect 18944 -5300 18950 -5240
rect 13622 -5650 18266 -5590
rect 19120 -5720 19180 -5068
rect 19574 -5068 19590 -5006
rect 19624 -3568 19638 -3492
rect 20036 -3492 20096 -2704
rect 20036 -3562 20048 -3492
rect 19624 -5006 19630 -3568
rect 19624 -5068 19634 -5006
rect 20042 -5024 20048 -3562
rect 19274 -5127 19482 -5121
rect 19274 -5161 19286 -5127
rect 19470 -5161 19482 -5127
rect 19274 -5167 19482 -5161
rect 19344 -5240 19404 -5167
rect 19338 -5300 19344 -5240
rect 19404 -5300 19410 -5240
rect 19574 -5242 19634 -5068
rect 20032 -5068 20048 -5024
rect 20082 -3562 20096 -3492
rect 20082 -5024 20088 -3562
rect 20082 -5068 20092 -5024
rect 19732 -5127 19940 -5121
rect 19732 -5161 19744 -5127
rect 19928 -5161 19940 -5127
rect 19732 -5167 19940 -5161
rect 19806 -5242 19866 -5167
rect 20032 -5242 20092 -5068
rect 21156 -5242 21162 -2418
rect 19574 -5302 21162 -5242
rect 10918 -7590 10924 -5732
rect 11232 -6157 11292 -5732
rect 11460 -6058 11520 -5732
rect 12704 -5780 19180 -5720
rect 20032 -5736 20092 -5302
rect 21156 -5736 21162 -5302
rect 20032 -5796 21162 -5736
rect 11684 -5886 11690 -5826
rect 11750 -5886 11756 -5826
rect 11387 -6064 11595 -6058
rect 11387 -6098 11399 -6064
rect 11583 -6098 11595 -6064
rect 11387 -6104 11595 -6098
rect 11232 -6204 11245 -6157
rect 11239 -7312 11245 -6204
rect 10812 -7766 10924 -7590
rect 11232 -7333 11245 -7312
rect 11279 -6204 11292 -6157
rect 11690 -6157 11750 -5886
rect 11922 -5988 15124 -5928
rect 15184 -5988 15190 -5928
rect 11922 -6058 11982 -5988
rect 12384 -6058 12444 -5988
rect 12838 -6058 12898 -5988
rect 13300 -6058 13360 -5988
rect 13754 -6058 13814 -5988
rect 14204 -6058 14264 -5988
rect 14670 -6058 14730 -5988
rect 15126 -6058 15186 -5988
rect 15582 -6006 16750 -5946
rect 15582 -6058 15642 -6006
rect 11845 -6064 12053 -6058
rect 11845 -6098 11857 -6064
rect 12041 -6098 12053 -6064
rect 11845 -6104 12053 -6098
rect 12303 -6064 12511 -6058
rect 12303 -6098 12315 -6064
rect 12499 -6098 12511 -6064
rect 12303 -6104 12511 -6098
rect 12761 -6064 12969 -6058
rect 12761 -6098 12773 -6064
rect 12957 -6098 12969 -6064
rect 12761 -6104 12969 -6098
rect 13219 -6064 13427 -6058
rect 13219 -6098 13231 -6064
rect 13415 -6098 13427 -6064
rect 13219 -6104 13427 -6098
rect 13677 -6064 13885 -6058
rect 13677 -6098 13689 -6064
rect 13873 -6098 13885 -6064
rect 13677 -6104 13885 -6098
rect 14135 -6064 14343 -6058
rect 14135 -6098 14147 -6064
rect 14331 -6098 14343 -6064
rect 14135 -6104 14343 -6098
rect 14593 -6064 14801 -6058
rect 14593 -6098 14605 -6064
rect 14789 -6098 14801 -6064
rect 14593 -6104 14801 -6098
rect 15051 -6064 15259 -6058
rect 15051 -6098 15063 -6064
rect 15247 -6098 15259 -6064
rect 15051 -6104 15259 -6098
rect 15509 -6064 15717 -6058
rect 15509 -6098 15521 -6064
rect 15705 -6098 15717 -6064
rect 15509 -6104 15717 -6098
rect 11279 -7312 11285 -6204
rect 11690 -6224 11703 -6157
rect 11279 -7333 11292 -7312
rect 11232 -7766 11292 -7333
rect 11697 -7333 11703 -6224
rect 11737 -6224 11750 -6157
rect 12155 -6157 12201 -6145
rect 11737 -7333 11743 -6224
rect 11697 -7345 11743 -7333
rect 12155 -7333 12161 -6157
rect 12195 -7333 12201 -6157
rect 12155 -7345 12201 -7333
rect 12613 -6157 12659 -6145
rect 12613 -7333 12619 -6157
rect 12653 -7333 12659 -6157
rect 12613 -7345 12659 -7333
rect 13071 -6157 13117 -6145
rect 13071 -7333 13077 -6157
rect 13111 -7333 13117 -6157
rect 13071 -7345 13117 -7333
rect 13529 -6157 13575 -6145
rect 13529 -7333 13535 -6157
rect 13569 -7333 13575 -6157
rect 13529 -7345 13575 -7333
rect 13987 -6157 14033 -6145
rect 13987 -7333 13993 -6157
rect 14027 -7333 14033 -6157
rect 13987 -7345 14033 -7333
rect 14445 -6157 14491 -6145
rect 14445 -7333 14451 -6157
rect 14485 -7333 14491 -6157
rect 14445 -7345 14491 -7333
rect 14903 -6157 14949 -6145
rect 14903 -7333 14909 -6157
rect 14943 -7333 14949 -6157
rect 15361 -6157 15407 -6145
rect 15361 -7266 15367 -6157
rect 14903 -7345 14949 -7333
rect 15352 -7333 15367 -7266
rect 15401 -7266 15407 -6157
rect 15812 -6157 15872 -6006
rect 15812 -6172 15825 -6157
rect 15401 -7333 15412 -7266
rect 15819 -7298 15825 -6172
rect 11387 -7392 11595 -7386
rect 11387 -7426 11399 -7392
rect 11583 -7426 11595 -7392
rect 11387 -7432 11595 -7426
rect 11845 -7392 12053 -7386
rect 11845 -7426 11857 -7392
rect 12041 -7426 12053 -7392
rect 11845 -7432 12053 -7426
rect 12303 -7392 12511 -7386
rect 12303 -7426 12315 -7392
rect 12499 -7426 12511 -7392
rect 12303 -7432 12511 -7426
rect 12761 -7392 12969 -7386
rect 12761 -7426 12773 -7392
rect 12957 -7426 12969 -7392
rect 12761 -7432 12969 -7426
rect 13219 -7392 13427 -7386
rect 13219 -7426 13231 -7392
rect 13415 -7426 13427 -7392
rect 13219 -7432 13427 -7426
rect 13677 -7392 13885 -7386
rect 13677 -7426 13689 -7392
rect 13873 -7426 13885 -7392
rect 13677 -7432 13885 -7426
rect 14135 -7392 14343 -7386
rect 14135 -7426 14147 -7392
rect 14331 -7426 14343 -7392
rect 14135 -7432 14343 -7426
rect 14593 -7392 14801 -7386
rect 14593 -7426 14605 -7392
rect 14789 -7426 14801 -7392
rect 14593 -7432 14801 -7426
rect 15051 -7392 15259 -7386
rect 15051 -7426 15063 -7392
rect 15247 -7426 15259 -7392
rect 15051 -7432 15259 -7426
rect 11460 -7766 11520 -7432
rect 11914 -7500 11974 -7432
rect 12376 -7500 12436 -7432
rect 12830 -7500 12890 -7432
rect 13292 -7500 13352 -7432
rect 13746 -7500 13806 -7432
rect 14196 -7500 14256 -7432
rect 14662 -7500 14722 -7432
rect 15118 -7500 15178 -7432
rect 11914 -7504 12830 -7500
rect 11974 -7560 12376 -7504
rect 11914 -7570 11974 -7564
rect 12436 -7560 12830 -7504
rect 12890 -7560 13292 -7500
rect 13352 -7506 14196 -7500
rect 13352 -7560 13746 -7506
rect 12376 -7570 12436 -7564
rect 12830 -7566 12890 -7560
rect 13292 -7566 13352 -7560
rect 13806 -7560 14196 -7506
rect 14256 -7560 14662 -7500
rect 14722 -7504 15178 -7500
rect 14722 -7560 15118 -7504
rect 14196 -7566 14256 -7560
rect 14662 -7566 14722 -7560
rect 13746 -7572 13806 -7566
rect 15118 -7570 15178 -7564
rect 15352 -7626 15412 -7333
rect 15810 -7333 15825 -7298
rect 15859 -6172 15872 -6157
rect 16232 -6157 16292 -6006
rect 16464 -6058 16524 -6006
rect 16387 -6064 16595 -6058
rect 16387 -6098 16399 -6064
rect 16583 -6098 16595 -6064
rect 16387 -6104 16595 -6098
rect 15859 -7298 15865 -6172
rect 16232 -6178 16245 -6157
rect 16239 -7298 16245 -6178
rect 15859 -7333 15870 -7298
rect 15509 -7392 15717 -7386
rect 15509 -7426 15521 -7392
rect 15705 -7426 15717 -7392
rect 15509 -7432 15717 -7426
rect 15346 -7686 15352 -7626
rect 15412 -7686 15418 -7626
rect 15582 -7766 15642 -7432
rect 15810 -7766 15870 -7333
rect 16230 -7333 16245 -7298
rect 16279 -6178 16292 -6157
rect 16690 -6157 16750 -6006
rect 16916 -5988 20180 -5928
rect 16916 -6058 16976 -5988
rect 17378 -6058 17438 -5988
rect 17832 -6058 17892 -5988
rect 18294 -6058 18354 -5988
rect 18748 -6058 18808 -5988
rect 19198 -6058 19258 -5988
rect 19664 -6058 19724 -5988
rect 20120 -6058 20180 -5988
rect 20582 -6058 20642 -5796
rect 16845 -6064 17053 -6058
rect 16845 -6098 16857 -6064
rect 17041 -6098 17053 -6064
rect 16845 -6104 17053 -6098
rect 17303 -6064 17511 -6058
rect 17303 -6098 17315 -6064
rect 17499 -6098 17511 -6064
rect 17303 -6104 17511 -6098
rect 17761 -6064 17969 -6058
rect 17761 -6098 17773 -6064
rect 17957 -6098 17969 -6064
rect 17761 -6104 17969 -6098
rect 18219 -6064 18427 -6058
rect 18219 -6098 18231 -6064
rect 18415 -6098 18427 -6064
rect 18219 -6104 18427 -6098
rect 18677 -6064 18885 -6058
rect 18677 -6098 18689 -6064
rect 18873 -6098 18885 -6064
rect 18677 -6104 18885 -6098
rect 19135 -6064 19343 -6058
rect 19135 -6098 19147 -6064
rect 19331 -6098 19343 -6064
rect 19135 -6104 19343 -6098
rect 19593 -6064 19801 -6058
rect 19593 -6098 19605 -6064
rect 19789 -6098 19801 -6064
rect 19593 -6104 19801 -6098
rect 20051 -6064 20259 -6058
rect 20051 -6098 20063 -6064
rect 20247 -6098 20259 -6064
rect 20051 -6104 20259 -6098
rect 20509 -6064 20717 -6058
rect 20509 -6098 20521 -6064
rect 20705 -6098 20717 -6064
rect 20509 -6104 20717 -6098
rect 16279 -7298 16285 -6178
rect 16690 -6200 16703 -6157
rect 16697 -7292 16703 -6200
rect 16279 -7333 16290 -7298
rect 16230 -7766 16290 -7333
rect 16688 -7333 16703 -7292
rect 16737 -6200 16750 -6157
rect 17155 -6157 17201 -6145
rect 16737 -7292 16743 -6200
rect 16737 -7333 16748 -7292
rect 16387 -7392 16595 -7386
rect 16387 -7426 16399 -7392
rect 16583 -7426 16595 -7392
rect 16387 -7432 16595 -7426
rect 16458 -7766 16518 -7432
rect 16688 -7766 16748 -7333
rect 17155 -7333 17161 -6157
rect 17195 -7333 17201 -6157
rect 17155 -7345 17201 -7333
rect 17613 -6157 17659 -6145
rect 17613 -7333 17619 -6157
rect 17653 -7333 17659 -6157
rect 17613 -7345 17659 -7333
rect 18071 -6157 18117 -6145
rect 18071 -7333 18077 -6157
rect 18111 -7333 18117 -6157
rect 18071 -7345 18117 -7333
rect 18529 -6157 18575 -6145
rect 18529 -7333 18535 -6157
rect 18569 -7333 18575 -6157
rect 18529 -7345 18575 -7333
rect 18987 -6157 19033 -6145
rect 18987 -7333 18993 -6157
rect 19027 -7333 19033 -6157
rect 18987 -7345 19033 -7333
rect 19445 -6157 19491 -6145
rect 19445 -7333 19451 -6157
rect 19485 -7333 19491 -6157
rect 19445 -7345 19491 -7333
rect 19903 -6157 19949 -6145
rect 19903 -7333 19909 -6157
rect 19943 -7333 19949 -6157
rect 20361 -6157 20407 -6145
rect 20361 -7326 20367 -6157
rect 19903 -7345 19949 -7333
rect 20352 -7333 20367 -7326
rect 20401 -7326 20407 -6157
rect 20808 -6157 20868 -5796
rect 20808 -6210 20825 -6157
rect 20819 -7300 20825 -6210
rect 20401 -7333 20412 -7326
rect 16845 -7392 17053 -7386
rect 16845 -7426 16857 -7392
rect 17041 -7426 17053 -7392
rect 16845 -7432 17053 -7426
rect 17303 -7392 17511 -7386
rect 17303 -7426 17315 -7392
rect 17499 -7426 17511 -7392
rect 17303 -7432 17511 -7426
rect 17761 -7392 17969 -7386
rect 17761 -7426 17773 -7392
rect 17957 -7426 17969 -7392
rect 17761 -7432 17969 -7426
rect 18219 -7392 18427 -7386
rect 18219 -7426 18231 -7392
rect 18415 -7426 18427 -7392
rect 18219 -7432 18427 -7426
rect 18677 -7392 18885 -7386
rect 18677 -7426 18689 -7392
rect 18873 -7426 18885 -7392
rect 18677 -7432 18885 -7426
rect 19135 -7392 19343 -7386
rect 19135 -7426 19147 -7392
rect 19331 -7426 19343 -7392
rect 19135 -7432 19343 -7426
rect 19593 -7392 19801 -7386
rect 19593 -7426 19605 -7392
rect 19789 -7426 19801 -7392
rect 19593 -7432 19801 -7426
rect 20051 -7392 20259 -7386
rect 20051 -7426 20063 -7392
rect 20247 -7426 20259 -7392
rect 20051 -7432 20259 -7426
rect 16916 -7500 16976 -7432
rect 17378 -7496 17438 -7432
rect 16916 -7504 17378 -7500
rect 16976 -7556 17378 -7504
rect 17832 -7500 17892 -7432
rect 18294 -7500 18354 -7432
rect 18748 -7500 18808 -7432
rect 19198 -7496 19258 -7432
rect 17438 -7502 19198 -7500
rect 17438 -7556 17832 -7502
rect 16976 -7560 17832 -7556
rect 17378 -7562 17438 -7560
rect 17892 -7560 18294 -7502
rect 16916 -7570 16976 -7564
rect 17832 -7568 17892 -7562
rect 18354 -7560 18748 -7502
rect 18294 -7568 18354 -7562
rect 18808 -7556 19198 -7502
rect 19664 -7500 19724 -7432
rect 20120 -7500 20180 -7432
rect 19258 -7502 20180 -7500
rect 19258 -7556 19664 -7502
rect 18808 -7560 19664 -7556
rect 19198 -7562 19258 -7560
rect 19724 -7560 20120 -7502
rect 18748 -7568 18808 -7562
rect 19664 -7568 19724 -7562
rect 20120 -7568 20180 -7562
rect 20352 -7632 20412 -7333
rect 20810 -7333 20825 -7300
rect 20859 -6210 20868 -6157
rect 20859 -7300 20865 -6210
rect 20859 -7333 20870 -7300
rect 20509 -7392 20717 -7386
rect 20509 -7426 20521 -7392
rect 20705 -7426 20717 -7392
rect 20509 -7432 20717 -7426
rect 20352 -7698 20412 -7692
rect 20582 -7766 20642 -7432
rect 20810 -7766 20870 -7333
rect 21156 -7590 21162 -5796
rect 21262 -7590 21268 -2418
rect 25234 -5664 25294 2284
rect 30504 2278 30564 2284
rect 31506 2280 31566 2284
rect 31506 2274 31666 2280
rect 31506 2226 31606 2274
rect 31654 2226 31666 2274
rect 31506 2220 31666 2226
rect 31700 2276 31908 2282
rect 31700 2228 31712 2276
rect 31760 2228 31848 2276
rect 31896 2228 31908 2276
rect 31700 2222 31908 2228
rect 32192 2276 32478 2282
rect 32192 2228 32204 2276
rect 32252 2228 32478 2276
rect 32192 2222 32478 2228
rect 25546 2200 25606 2206
rect 25400 -420 25406 -360
rect 25466 -420 25472 -360
rect 25406 -3260 25466 -420
rect 25406 -3266 25468 -3260
rect 25406 -3326 25408 -3266
rect 25406 -3332 25468 -3326
rect 25228 -5724 25234 -5664
rect 25294 -5724 25300 -5664
rect 21156 -7766 21268 -7590
rect 10812 -7772 21268 -7766
rect 10812 -7872 10918 -7772
rect 21162 -7872 21268 -7772
rect 10812 -7878 21268 -7872
rect 10812 -8108 21268 -8102
rect 10812 -8208 10918 -8108
rect 21162 -8208 21268 -8108
rect 10812 -8214 21268 -8208
rect 10812 -8338 10924 -8214
rect 10812 -10342 10818 -8338
rect 10918 -10342 10924 -8338
rect 11232 -8650 11292 -8214
rect 11462 -8560 11522 -8214
rect 15352 -8306 15412 -8300
rect 11920 -8440 12376 -8434
rect 11908 -8500 11914 -8440
rect 11974 -8494 12376 -8440
rect 12436 -8440 13292 -8434
rect 12436 -8494 12830 -8440
rect 11974 -8500 11980 -8494
rect 11914 -8560 11980 -8500
rect 12376 -8560 12442 -8494
rect 12824 -8500 12830 -8494
rect 12890 -8494 13292 -8440
rect 13352 -8494 13746 -8434
rect 13806 -8494 14196 -8434
rect 14256 -8440 15118 -8434
rect 14256 -8494 14662 -8440
rect 12890 -8500 12896 -8494
rect 12830 -8560 12896 -8500
rect 13292 -8560 13358 -8494
rect 13746 -8560 13812 -8494
rect 14196 -8560 14262 -8494
rect 14656 -8500 14662 -8494
rect 14722 -8494 15118 -8440
rect 15178 -8494 15184 -8434
rect 14722 -8500 14728 -8494
rect 14662 -8560 14728 -8500
rect 15118 -8560 15184 -8494
rect 11386 -8566 11594 -8560
rect 11386 -8600 11398 -8566
rect 11582 -8600 11594 -8566
rect 11386 -8606 11594 -8600
rect 11844 -8566 12052 -8560
rect 11844 -8600 11856 -8566
rect 12040 -8600 12052 -8566
rect 11844 -8606 12052 -8600
rect 12302 -8566 12510 -8560
rect 12302 -8600 12314 -8566
rect 12498 -8600 12510 -8566
rect 12302 -8606 12510 -8600
rect 12760 -8566 12968 -8560
rect 12760 -8600 12772 -8566
rect 12956 -8600 12968 -8566
rect 12760 -8606 12968 -8600
rect 13218 -8566 13426 -8560
rect 13218 -8600 13230 -8566
rect 13414 -8600 13426 -8566
rect 13218 -8606 13426 -8600
rect 13676 -8566 13884 -8560
rect 13676 -8600 13688 -8566
rect 13872 -8600 13884 -8566
rect 13676 -8606 13884 -8600
rect 14134 -8566 14342 -8560
rect 14134 -8600 14146 -8566
rect 14330 -8600 14342 -8566
rect 14134 -8606 14342 -8600
rect 14592 -8566 14800 -8560
rect 14592 -8600 14604 -8566
rect 14788 -8600 14800 -8566
rect 14592 -8606 14800 -8600
rect 15050 -8566 15258 -8560
rect 15050 -8600 15062 -8566
rect 15246 -8600 15258 -8566
rect 15050 -8606 15258 -8600
rect 11232 -8690 11244 -8650
rect 11238 -8786 11244 -8690
rect 11232 -8826 11244 -8786
rect 11278 -8690 11292 -8650
rect 11696 -8650 11742 -8638
rect 11278 -8786 11284 -8690
rect 11696 -8784 11702 -8650
rect 11278 -8826 11292 -8786
rect 11232 -9042 11292 -8826
rect 11688 -8826 11702 -8784
rect 11736 -8784 11742 -8650
rect 12154 -8650 12200 -8638
rect 11736 -8826 11748 -8784
rect 11386 -8876 11594 -8870
rect 11386 -8910 11398 -8876
rect 11582 -8910 11594 -8876
rect 11386 -8916 11594 -8910
rect 11460 -9042 11520 -8916
rect 11232 -9102 11520 -9042
rect 11232 -9318 11292 -9102
rect 11460 -9228 11520 -9102
rect 11386 -9234 11594 -9228
rect 11386 -9268 11398 -9234
rect 11582 -9268 11594 -9234
rect 11386 -9274 11594 -9268
rect 11232 -9338 11244 -9318
rect 11238 -9464 11244 -9338
rect 11224 -9494 11244 -9464
rect 11278 -9338 11292 -9318
rect 11688 -9318 11748 -8826
rect 12154 -8826 12160 -8650
rect 12194 -8826 12200 -8650
rect 12154 -8838 12200 -8826
rect 12612 -8650 12658 -8638
rect 12612 -8826 12618 -8650
rect 12652 -8826 12658 -8650
rect 12612 -8838 12658 -8826
rect 13070 -8650 13116 -8638
rect 13070 -8826 13076 -8650
rect 13110 -8826 13116 -8650
rect 13070 -8838 13116 -8826
rect 13528 -8650 13574 -8638
rect 13528 -8826 13534 -8650
rect 13568 -8826 13574 -8650
rect 13528 -8838 13574 -8826
rect 13986 -8650 14032 -8638
rect 13986 -8826 13992 -8650
rect 14026 -8826 14032 -8650
rect 13986 -8838 14032 -8826
rect 14444 -8650 14490 -8638
rect 14444 -8826 14450 -8650
rect 14484 -8826 14490 -8650
rect 14444 -8838 14490 -8826
rect 14902 -8650 14948 -8638
rect 14902 -8826 14908 -8650
rect 14942 -8826 14948 -8650
rect 15352 -8650 15412 -8366
rect 15580 -8560 15640 -8214
rect 15508 -8566 15716 -8560
rect 15508 -8600 15520 -8566
rect 15704 -8600 15716 -8566
rect 15508 -8606 15716 -8600
rect 15352 -8680 15366 -8650
rect 14902 -8838 14948 -8826
rect 15360 -8826 15366 -8680
rect 15400 -8680 15412 -8650
rect 15812 -8650 15872 -8214
rect 15812 -8678 15824 -8650
rect 15400 -8826 15406 -8680
rect 15818 -8770 15824 -8678
rect 15360 -8838 15406 -8826
rect 15812 -8826 15824 -8770
rect 15858 -8678 15872 -8650
rect 16232 -8650 16292 -8214
rect 16466 -8560 16526 -8214
rect 16386 -8566 16594 -8560
rect 16386 -8600 16398 -8566
rect 16582 -8600 16594 -8566
rect 16386 -8606 16594 -8600
rect 15858 -8770 15864 -8678
rect 16232 -8686 16244 -8650
rect 15858 -8826 15872 -8770
rect 16238 -8790 16244 -8686
rect 11844 -8876 12052 -8870
rect 11844 -8910 11856 -8876
rect 12040 -8910 12052 -8876
rect 11844 -8916 12052 -8910
rect 12302 -8876 12510 -8870
rect 12302 -8910 12314 -8876
rect 12498 -8910 12510 -8876
rect 12302 -8916 12510 -8910
rect 12760 -8876 12968 -8870
rect 12760 -8910 12772 -8876
rect 12956 -8910 12968 -8876
rect 12760 -8916 12968 -8910
rect 13218 -8876 13426 -8870
rect 13218 -8910 13230 -8876
rect 13414 -8910 13426 -8876
rect 13218 -8916 13426 -8910
rect 13676 -8876 13884 -8870
rect 13676 -8910 13688 -8876
rect 13872 -8910 13884 -8876
rect 13676 -8916 13884 -8910
rect 14134 -8876 14342 -8870
rect 14134 -8910 14146 -8876
rect 14330 -8910 14342 -8876
rect 14134 -8916 14342 -8910
rect 14592 -8876 14800 -8870
rect 14592 -8910 14604 -8876
rect 14788 -8910 14800 -8876
rect 14592 -8916 14800 -8910
rect 15050 -8876 15258 -8870
rect 15050 -8910 15062 -8876
rect 15246 -8910 15258 -8876
rect 15050 -8916 15258 -8910
rect 15508 -8876 15716 -8870
rect 15508 -8910 15520 -8876
rect 15704 -8910 15716 -8876
rect 15508 -8916 15716 -8910
rect 11914 -8982 11974 -8916
rect 12376 -8982 12436 -8916
rect 12830 -8982 12890 -8916
rect 13292 -8982 13352 -8916
rect 13746 -8982 13806 -8916
rect 14196 -8982 14256 -8916
rect 14662 -8982 14722 -8916
rect 15118 -8982 15178 -8916
rect 11914 -9042 15178 -8982
rect 11920 -9162 15184 -9102
rect 11920 -9228 11980 -9162
rect 12382 -9228 12442 -9162
rect 12836 -9228 12896 -9162
rect 13298 -9228 13358 -9162
rect 13752 -9228 13812 -9162
rect 14202 -9228 14262 -9162
rect 14668 -9228 14728 -9162
rect 15124 -9228 15184 -9162
rect 15580 -9228 15640 -8916
rect 11844 -9234 12052 -9228
rect 11844 -9268 11856 -9234
rect 12040 -9268 12052 -9234
rect 11844 -9274 12052 -9268
rect 12302 -9234 12510 -9228
rect 12302 -9268 12314 -9234
rect 12498 -9268 12510 -9234
rect 12302 -9274 12510 -9268
rect 12760 -9234 12968 -9228
rect 12760 -9268 12772 -9234
rect 12956 -9268 12968 -9234
rect 12760 -9274 12968 -9268
rect 13218 -9234 13426 -9228
rect 13218 -9268 13230 -9234
rect 13414 -9268 13426 -9234
rect 13218 -9274 13426 -9268
rect 13676 -9234 13884 -9228
rect 13676 -9268 13688 -9234
rect 13872 -9268 13884 -9234
rect 13676 -9274 13884 -9268
rect 14134 -9234 14342 -9228
rect 14134 -9268 14146 -9234
rect 14330 -9268 14342 -9234
rect 14134 -9274 14342 -9268
rect 14592 -9234 14800 -9228
rect 14592 -9268 14604 -9234
rect 14788 -9268 14800 -9234
rect 14592 -9274 14800 -9268
rect 15050 -9234 15258 -9228
rect 15050 -9268 15062 -9234
rect 15246 -9268 15258 -9234
rect 15050 -9274 15258 -9268
rect 15508 -9234 15716 -9228
rect 15508 -9268 15520 -9234
rect 15704 -9268 15716 -9234
rect 15508 -9274 15716 -9268
rect 11278 -9494 11284 -9338
rect 11688 -9346 11702 -9318
rect 11224 -9874 11284 -9494
rect 11696 -9494 11702 -9346
rect 11736 -9346 11748 -9318
rect 12154 -9318 12200 -9306
rect 11736 -9494 11742 -9346
rect 11696 -9506 11742 -9494
rect 12154 -9494 12160 -9318
rect 12194 -9494 12200 -9318
rect 12154 -9506 12200 -9494
rect 12612 -9318 12658 -9306
rect 12612 -9494 12618 -9318
rect 12652 -9494 12658 -9318
rect 12612 -9506 12658 -9494
rect 13070 -9318 13116 -9306
rect 13070 -9494 13076 -9318
rect 13110 -9494 13116 -9318
rect 13070 -9506 13116 -9494
rect 13528 -9318 13574 -9306
rect 13528 -9494 13534 -9318
rect 13568 -9494 13574 -9318
rect 13528 -9506 13574 -9494
rect 13986 -9318 14032 -9306
rect 13986 -9494 13992 -9318
rect 14026 -9494 14032 -9318
rect 13986 -9506 14032 -9494
rect 14444 -9318 14490 -9306
rect 14444 -9494 14450 -9318
rect 14484 -9494 14490 -9318
rect 14444 -9506 14490 -9494
rect 14902 -9318 14948 -9306
rect 14902 -9494 14908 -9318
rect 14942 -9494 14948 -9318
rect 15360 -9318 15406 -9306
rect 15360 -9466 15366 -9318
rect 14902 -9506 14948 -9494
rect 15352 -9494 15366 -9466
rect 15400 -9466 15406 -9318
rect 15812 -9318 15872 -8826
rect 15400 -9494 15412 -9466
rect 11386 -9544 11594 -9538
rect 11386 -9578 11398 -9544
rect 11582 -9578 11594 -9544
rect 11386 -9584 11594 -9578
rect 11844 -9544 12052 -9538
rect 11844 -9578 11856 -9544
rect 12040 -9578 12052 -9544
rect 11844 -9584 12052 -9578
rect 12302 -9544 12510 -9538
rect 12302 -9578 12314 -9544
rect 12498 -9578 12510 -9544
rect 12302 -9584 12510 -9578
rect 12760 -9544 12968 -9538
rect 12760 -9578 12772 -9544
rect 12956 -9578 12968 -9544
rect 12760 -9584 12968 -9578
rect 13218 -9544 13426 -9538
rect 13218 -9578 13230 -9544
rect 13414 -9578 13426 -9544
rect 13218 -9584 13426 -9578
rect 13676 -9544 13884 -9538
rect 13676 -9578 13688 -9544
rect 13872 -9578 13884 -9544
rect 13676 -9584 13884 -9578
rect 14134 -9544 14342 -9538
rect 14134 -9578 14146 -9544
rect 14330 -9578 14342 -9544
rect 14134 -9584 14342 -9578
rect 14592 -9544 14800 -9538
rect 14592 -9578 14604 -9544
rect 14788 -9578 14800 -9544
rect 14592 -9584 14800 -9578
rect 15050 -9544 15258 -9538
rect 15050 -9578 15062 -9544
rect 15246 -9578 15258 -9544
rect 15050 -9584 15258 -9578
rect 11464 -9874 11524 -9584
rect 11914 -9650 11974 -9584
rect 12376 -9650 12436 -9584
rect 12830 -9650 12890 -9584
rect 13292 -9650 13352 -9584
rect 13746 -9650 13806 -9584
rect 14196 -9650 14256 -9584
rect 14662 -9650 14722 -9584
rect 15118 -9650 15178 -9584
rect 11914 -9710 15116 -9650
rect 15176 -9710 15182 -9650
rect 15352 -9874 15412 -9494
rect 15812 -9494 15824 -9318
rect 15858 -9494 15872 -9318
rect 15508 -9544 15716 -9538
rect 15508 -9578 15520 -9544
rect 15704 -9578 15716 -9544
rect 15508 -9584 15716 -9578
rect 15578 -9874 15638 -9584
rect 15812 -9874 15872 -9494
rect 16228 -8826 16244 -8790
rect 16278 -8686 16292 -8650
rect 16688 -8650 16748 -8214
rect 20346 -8354 20352 -8294
rect 20412 -8354 20418 -8294
rect 19192 -8434 19198 -8430
rect 16910 -8494 16916 -8434
rect 16976 -8436 19198 -8434
rect 16976 -8494 17378 -8436
rect 16916 -8560 16980 -8494
rect 17372 -8496 17378 -8494
rect 17438 -8494 17832 -8436
rect 17438 -8496 17444 -8494
rect 17826 -8496 17832 -8494
rect 17892 -8494 18294 -8436
rect 17892 -8496 17898 -8494
rect 18288 -8496 18294 -8494
rect 18354 -8494 18748 -8436
rect 18354 -8496 18360 -8494
rect 18742 -8496 18748 -8494
rect 18808 -8490 19198 -8436
rect 19258 -8434 19264 -8430
rect 19258 -8490 19664 -8434
rect 18808 -8494 19664 -8490
rect 19724 -8494 20120 -8434
rect 20180 -8494 20186 -8434
rect 18808 -8496 18814 -8494
rect 17378 -8560 17442 -8496
rect 17832 -8560 17896 -8496
rect 18294 -8560 18358 -8496
rect 18748 -8560 18812 -8496
rect 19198 -8560 19262 -8494
rect 19664 -8560 19728 -8494
rect 20120 -8560 20184 -8494
rect 16844 -8566 17052 -8560
rect 16844 -8600 16856 -8566
rect 17040 -8600 17052 -8566
rect 16844 -8606 17052 -8600
rect 17302 -8566 17510 -8560
rect 17302 -8600 17314 -8566
rect 17498 -8600 17510 -8566
rect 17302 -8606 17510 -8600
rect 17760 -8566 17968 -8560
rect 17760 -8600 17772 -8566
rect 17956 -8600 17968 -8566
rect 17760 -8606 17968 -8600
rect 18218 -8566 18426 -8560
rect 18218 -8600 18230 -8566
rect 18414 -8600 18426 -8566
rect 18218 -8606 18426 -8600
rect 18676 -8566 18884 -8560
rect 18676 -8600 18688 -8566
rect 18872 -8600 18884 -8566
rect 18676 -8606 18884 -8600
rect 19134 -8566 19342 -8560
rect 19134 -8600 19146 -8566
rect 19330 -8600 19342 -8566
rect 19134 -8606 19342 -8600
rect 19592 -8566 19800 -8560
rect 19592 -8600 19604 -8566
rect 19788 -8600 19800 -8566
rect 19592 -8606 19800 -8600
rect 20050 -8566 20258 -8560
rect 20050 -8600 20062 -8566
rect 20246 -8600 20258 -8566
rect 20050 -8606 20258 -8600
rect 16278 -8790 16284 -8686
rect 16688 -8714 16702 -8650
rect 16696 -8782 16702 -8714
rect 16278 -8826 16288 -8790
rect 16228 -8980 16288 -8826
rect 16688 -8826 16702 -8782
rect 16736 -8714 16748 -8650
rect 17154 -8650 17200 -8638
rect 16736 -8782 16742 -8714
rect 16736 -8826 16748 -8782
rect 16386 -8876 16594 -8870
rect 16386 -8910 16398 -8876
rect 16582 -8910 16594 -8876
rect 16386 -8916 16594 -8910
rect 16456 -8980 16516 -8916
rect 16688 -8980 16748 -8826
rect 17154 -8826 17160 -8650
rect 17194 -8826 17200 -8650
rect 17154 -8838 17200 -8826
rect 17612 -8650 17658 -8638
rect 17612 -8826 17618 -8650
rect 17652 -8826 17658 -8650
rect 17612 -8838 17658 -8826
rect 18070 -8650 18116 -8638
rect 18070 -8826 18076 -8650
rect 18110 -8826 18116 -8650
rect 18070 -8838 18116 -8826
rect 18528 -8650 18574 -8638
rect 18528 -8826 18534 -8650
rect 18568 -8826 18574 -8650
rect 18528 -8838 18574 -8826
rect 18986 -8650 19032 -8638
rect 18986 -8826 18992 -8650
rect 19026 -8826 19032 -8650
rect 18986 -8838 19032 -8826
rect 19444 -8650 19490 -8638
rect 19444 -8826 19450 -8650
rect 19484 -8826 19490 -8650
rect 19444 -8838 19490 -8826
rect 19902 -8650 19948 -8638
rect 19902 -8826 19908 -8650
rect 19942 -8826 19948 -8650
rect 20352 -8650 20412 -8354
rect 20592 -8560 20652 -8214
rect 20508 -8566 20716 -8560
rect 20508 -8600 20520 -8566
rect 20704 -8600 20716 -8566
rect 20508 -8606 20716 -8600
rect 20352 -8692 20366 -8650
rect 19902 -8838 19948 -8826
rect 20360 -8826 20366 -8692
rect 20400 -8692 20412 -8650
rect 20810 -8650 20870 -8214
rect 20810 -8690 20824 -8650
rect 20400 -8826 20406 -8692
rect 20818 -8780 20824 -8690
rect 20360 -8838 20406 -8826
rect 20808 -8826 20824 -8780
rect 20858 -8690 20870 -8650
rect 21156 -8338 21268 -8214
rect 20858 -8780 20864 -8690
rect 20858 -8826 20868 -8780
rect 16844 -8876 17052 -8870
rect 16844 -8910 16856 -8876
rect 17040 -8910 17052 -8876
rect 16844 -8916 17052 -8910
rect 17302 -8876 17510 -8870
rect 17302 -8910 17314 -8876
rect 17498 -8910 17510 -8876
rect 17302 -8916 17510 -8910
rect 17760 -8876 17968 -8870
rect 17760 -8910 17772 -8876
rect 17956 -8910 17968 -8876
rect 17760 -8916 17968 -8910
rect 18218 -8876 18426 -8870
rect 18218 -8910 18230 -8876
rect 18414 -8910 18426 -8876
rect 18218 -8916 18426 -8910
rect 18676 -8876 18884 -8870
rect 18676 -8910 18688 -8876
rect 18872 -8910 18884 -8876
rect 18676 -8916 18884 -8910
rect 19134 -8876 19342 -8870
rect 19134 -8910 19146 -8876
rect 19330 -8910 19342 -8876
rect 19134 -8916 19342 -8910
rect 19592 -8876 19800 -8870
rect 19592 -8910 19604 -8876
rect 19788 -8910 19800 -8876
rect 19592 -8916 19800 -8910
rect 20050 -8876 20258 -8870
rect 20050 -8910 20062 -8876
rect 20246 -8910 20258 -8876
rect 20050 -8916 20258 -8910
rect 20508 -8876 20716 -8870
rect 20508 -8910 20520 -8876
rect 20704 -8910 20716 -8876
rect 20508 -8916 20716 -8910
rect 16228 -9040 16748 -8980
rect 16228 -9874 16288 -9040
rect 16456 -9874 16516 -9040
rect 16688 -9874 16748 -9040
rect 16914 -8982 16974 -8916
rect 17376 -8982 17436 -8916
rect 17830 -8982 17890 -8916
rect 18292 -8982 18352 -8916
rect 18746 -8982 18806 -8916
rect 19196 -8982 19256 -8916
rect 19662 -8982 19722 -8916
rect 20118 -8982 20178 -8916
rect 16914 -9042 20178 -8982
rect 20582 -9874 20642 -8916
rect 20808 -9874 20868 -8826
rect 11160 -9902 20930 -9874
rect 11160 -9988 11210 -9902
rect 11306 -9988 11790 -9902
rect 11886 -9988 12390 -9902
rect 12486 -9988 12990 -9902
rect 13086 -9988 13590 -9902
rect 13686 -9988 14190 -9902
rect 14286 -9988 14790 -9902
rect 14886 -9988 15390 -9902
rect 15486 -9988 15990 -9902
rect 16086 -9988 16590 -9902
rect 16686 -9988 17190 -9902
rect 17286 -9988 17790 -9902
rect 17886 -9988 18390 -9902
rect 18486 -9988 18990 -9902
rect 19086 -9988 19590 -9902
rect 19686 -9988 20190 -9902
rect 20286 -9988 20790 -9902
rect 20886 -9988 20930 -9902
rect 11160 -10018 20930 -9988
rect 10812 -10466 10924 -10342
rect 11524 -10466 11534 -10166
rect 20546 -10466 20556 -10166
rect 21156 -10342 21162 -8338
rect 21262 -10342 21268 -8338
rect 21156 -10466 21268 -10342
rect 10812 -10472 21268 -10466
rect 10812 -10572 10918 -10472
rect 21162 -10572 21268 -10472
rect 10812 -10578 21268 -10572
rect 14766 -11032 25222 -11026
rect 14766 -11132 14872 -11032
rect 25116 -11132 25222 -11032
rect 14766 -11138 25222 -11132
rect 14766 -11262 14878 -11138
rect 14766 -13266 14772 -11262
rect 14872 -13266 14878 -11262
rect 15478 -11438 15488 -11138
rect 24500 -11438 24510 -11138
rect 25110 -11262 25222 -11138
rect 15104 -11616 24874 -11586
rect 15104 -11702 15148 -11616
rect 15244 -11702 15748 -11616
rect 15844 -11702 16348 -11616
rect 16444 -11702 16948 -11616
rect 17044 -11702 17548 -11616
rect 17644 -11702 18148 -11616
rect 18244 -11702 18748 -11616
rect 18844 -11702 19348 -11616
rect 19444 -11702 19948 -11616
rect 20044 -11702 20548 -11616
rect 20644 -11702 21148 -11616
rect 21244 -11702 21748 -11616
rect 21844 -11702 22348 -11616
rect 22444 -11702 22948 -11616
rect 23044 -11702 23548 -11616
rect 23644 -11702 24148 -11616
rect 24244 -11702 24728 -11616
rect 24824 -11702 24874 -11616
rect 15104 -11730 24874 -11702
rect 15166 -12778 15226 -11730
rect 15392 -12688 15452 -11730
rect 15856 -12622 19120 -12562
rect 15856 -12688 15916 -12622
rect 16312 -12688 16372 -12622
rect 16778 -12688 16838 -12622
rect 17228 -12688 17288 -12622
rect 17682 -12688 17742 -12622
rect 18144 -12688 18204 -12622
rect 18598 -12688 18658 -12622
rect 19060 -12688 19120 -12622
rect 19286 -12564 19346 -11730
rect 19518 -12564 19578 -11730
rect 19746 -12564 19806 -11730
rect 19286 -12624 19806 -12564
rect 15318 -12694 15526 -12688
rect 15318 -12728 15330 -12694
rect 15514 -12728 15526 -12694
rect 15318 -12734 15526 -12728
rect 15776 -12694 15984 -12688
rect 15776 -12728 15788 -12694
rect 15972 -12728 15984 -12694
rect 15776 -12734 15984 -12728
rect 16234 -12694 16442 -12688
rect 16234 -12728 16246 -12694
rect 16430 -12728 16442 -12694
rect 16234 -12734 16442 -12728
rect 16692 -12694 16900 -12688
rect 16692 -12728 16704 -12694
rect 16888 -12728 16900 -12694
rect 16692 -12734 16900 -12728
rect 17150 -12694 17358 -12688
rect 17150 -12728 17162 -12694
rect 17346 -12728 17358 -12694
rect 17150 -12734 17358 -12728
rect 17608 -12694 17816 -12688
rect 17608 -12728 17620 -12694
rect 17804 -12728 17816 -12694
rect 17608 -12734 17816 -12728
rect 18066 -12694 18274 -12688
rect 18066 -12728 18078 -12694
rect 18262 -12728 18274 -12694
rect 18066 -12734 18274 -12728
rect 18524 -12694 18732 -12688
rect 18524 -12728 18536 -12694
rect 18720 -12728 18732 -12694
rect 18524 -12734 18732 -12728
rect 18982 -12694 19190 -12688
rect 18982 -12728 18994 -12694
rect 19178 -12728 19190 -12694
rect 18982 -12734 19190 -12728
rect 15166 -12824 15176 -12778
rect 15170 -12914 15176 -12824
rect 14766 -13390 14878 -13266
rect 15164 -12954 15176 -12914
rect 15210 -12824 15226 -12778
rect 15628 -12778 15674 -12766
rect 15210 -12914 15216 -12824
rect 15628 -12912 15634 -12778
rect 15210 -12954 15224 -12914
rect 15164 -13390 15224 -12954
rect 15622 -12954 15634 -12912
rect 15668 -12912 15674 -12778
rect 16086 -12778 16132 -12766
rect 15668 -12954 15682 -12912
rect 15318 -13004 15526 -12998
rect 15318 -13038 15330 -13004
rect 15514 -13038 15526 -13004
rect 15318 -13044 15526 -13038
rect 15382 -13390 15442 -13044
rect 15622 -13250 15682 -12954
rect 16086 -12954 16092 -12778
rect 16126 -12954 16132 -12778
rect 16086 -12966 16132 -12954
rect 16544 -12778 16590 -12766
rect 16544 -12954 16550 -12778
rect 16584 -12954 16590 -12778
rect 16544 -12966 16590 -12954
rect 17002 -12778 17048 -12766
rect 17002 -12954 17008 -12778
rect 17042 -12954 17048 -12778
rect 17002 -12966 17048 -12954
rect 17460 -12778 17506 -12766
rect 17460 -12954 17466 -12778
rect 17500 -12954 17506 -12778
rect 17460 -12966 17506 -12954
rect 17918 -12778 17964 -12766
rect 17918 -12954 17924 -12778
rect 17958 -12954 17964 -12778
rect 17918 -12966 17964 -12954
rect 18376 -12778 18422 -12766
rect 18376 -12954 18382 -12778
rect 18416 -12954 18422 -12778
rect 18376 -12966 18422 -12954
rect 18834 -12778 18880 -12766
rect 18834 -12954 18840 -12778
rect 18874 -12954 18880 -12778
rect 19286 -12778 19346 -12624
rect 19518 -12688 19578 -12624
rect 19440 -12694 19648 -12688
rect 19440 -12728 19452 -12694
rect 19636 -12728 19648 -12694
rect 19440 -12734 19648 -12728
rect 19286 -12822 19298 -12778
rect 19292 -12890 19298 -12822
rect 18834 -12966 18880 -12954
rect 19286 -12954 19298 -12890
rect 19332 -12822 19346 -12778
rect 19746 -12778 19806 -12624
rect 19746 -12814 19756 -12778
rect 19332 -12890 19338 -12822
rect 19332 -12954 19346 -12890
rect 19750 -12918 19756 -12814
rect 15776 -13004 15984 -12998
rect 15776 -13038 15788 -13004
rect 15972 -13038 15984 -13004
rect 15776 -13044 15984 -13038
rect 16234 -13004 16442 -12998
rect 16234 -13038 16246 -13004
rect 16430 -13038 16442 -13004
rect 16234 -13044 16442 -13038
rect 16692 -13004 16900 -12998
rect 16692 -13038 16704 -13004
rect 16888 -13038 16900 -13004
rect 16692 -13044 16900 -13038
rect 17150 -13004 17358 -12998
rect 17150 -13038 17162 -13004
rect 17346 -13038 17358 -13004
rect 17150 -13044 17358 -13038
rect 17608 -13004 17816 -12998
rect 17608 -13038 17620 -13004
rect 17804 -13038 17816 -13004
rect 17608 -13044 17816 -13038
rect 18066 -13004 18274 -12998
rect 18066 -13038 18078 -13004
rect 18262 -13038 18274 -13004
rect 18066 -13044 18274 -13038
rect 18524 -13004 18732 -12998
rect 18524 -13038 18536 -13004
rect 18720 -13038 18732 -13004
rect 18524 -13044 18732 -13038
rect 18982 -13004 19190 -12998
rect 18982 -13038 18994 -13004
rect 19178 -13038 19190 -13004
rect 18982 -13044 19190 -13038
rect 15850 -13110 15914 -13044
rect 16306 -13110 16370 -13044
rect 16772 -13110 16836 -13044
rect 17222 -13108 17286 -13044
rect 17676 -13108 17740 -13044
rect 18138 -13108 18202 -13044
rect 18592 -13108 18656 -13044
rect 17220 -13110 17226 -13108
rect 15848 -13170 15854 -13110
rect 15914 -13170 16310 -13110
rect 16370 -13114 17226 -13110
rect 16370 -13170 16776 -13114
rect 16770 -13174 16776 -13170
rect 16836 -13168 17226 -13114
rect 17286 -13110 17292 -13108
rect 17674 -13110 17680 -13108
rect 17286 -13168 17680 -13110
rect 17740 -13110 17746 -13108
rect 18136 -13110 18142 -13108
rect 17740 -13168 18142 -13110
rect 18202 -13110 18208 -13108
rect 18590 -13110 18596 -13108
rect 18202 -13168 18596 -13110
rect 18656 -13110 18662 -13108
rect 19054 -13110 19118 -13044
rect 18656 -13168 19058 -13110
rect 16836 -13170 19058 -13168
rect 19118 -13170 19124 -13110
rect 16836 -13174 16842 -13170
rect 15616 -13310 15622 -13250
rect 15682 -13310 15688 -13250
rect 19286 -13390 19346 -12954
rect 19742 -12954 19756 -12918
rect 19790 -12814 19806 -12778
rect 20162 -12110 20222 -11730
rect 20396 -12020 20456 -11730
rect 20318 -12026 20526 -12020
rect 20318 -12060 20330 -12026
rect 20514 -12060 20526 -12026
rect 20318 -12066 20526 -12060
rect 20162 -12286 20176 -12110
rect 20210 -12286 20222 -12110
rect 20622 -12110 20682 -11730
rect 20856 -11954 24062 -11894
rect 24122 -11954 24128 -11894
rect 20856 -12020 20916 -11954
rect 21312 -12020 21372 -11954
rect 21778 -12020 21838 -11954
rect 22228 -12020 22288 -11954
rect 22682 -12020 22742 -11954
rect 23144 -12020 23204 -11954
rect 23598 -12020 23658 -11954
rect 24060 -12020 24120 -11954
rect 24510 -12020 24570 -11730
rect 20776 -12026 20984 -12020
rect 20776 -12060 20788 -12026
rect 20972 -12060 20984 -12026
rect 20776 -12066 20984 -12060
rect 21234 -12026 21442 -12020
rect 21234 -12060 21246 -12026
rect 21430 -12060 21442 -12026
rect 21234 -12066 21442 -12060
rect 21692 -12026 21900 -12020
rect 21692 -12060 21704 -12026
rect 21888 -12060 21900 -12026
rect 21692 -12066 21900 -12060
rect 22150 -12026 22358 -12020
rect 22150 -12060 22162 -12026
rect 22346 -12060 22358 -12026
rect 22150 -12066 22358 -12060
rect 22608 -12026 22816 -12020
rect 22608 -12060 22620 -12026
rect 22804 -12060 22816 -12026
rect 22608 -12066 22816 -12060
rect 23066 -12026 23274 -12020
rect 23066 -12060 23078 -12026
rect 23262 -12060 23274 -12026
rect 23066 -12066 23274 -12060
rect 23524 -12026 23732 -12020
rect 23524 -12060 23536 -12026
rect 23720 -12060 23732 -12026
rect 23524 -12066 23732 -12060
rect 23982 -12026 24190 -12020
rect 23982 -12060 23994 -12026
rect 24178 -12060 24190 -12026
rect 23982 -12066 24190 -12060
rect 24440 -12026 24648 -12020
rect 24440 -12060 24452 -12026
rect 24636 -12060 24648 -12026
rect 24440 -12066 24648 -12060
rect 20622 -12138 20634 -12110
rect 20162 -12778 20222 -12286
rect 20628 -12286 20634 -12138
rect 20668 -12138 20682 -12110
rect 21086 -12110 21132 -12098
rect 20668 -12286 20674 -12138
rect 20628 -12298 20674 -12286
rect 21086 -12286 21092 -12110
rect 21126 -12286 21132 -12110
rect 21086 -12298 21132 -12286
rect 21544 -12110 21590 -12098
rect 21544 -12286 21550 -12110
rect 21584 -12286 21590 -12110
rect 21544 -12298 21590 -12286
rect 22002 -12110 22048 -12098
rect 22002 -12286 22008 -12110
rect 22042 -12286 22048 -12110
rect 22002 -12298 22048 -12286
rect 22460 -12110 22506 -12098
rect 22460 -12286 22466 -12110
rect 22500 -12286 22506 -12110
rect 22460 -12298 22506 -12286
rect 22918 -12110 22964 -12098
rect 22918 -12286 22924 -12110
rect 22958 -12286 22964 -12110
rect 22918 -12298 22964 -12286
rect 23376 -12110 23422 -12098
rect 23376 -12286 23382 -12110
rect 23416 -12286 23422 -12110
rect 23376 -12298 23422 -12286
rect 23834 -12110 23880 -12098
rect 23834 -12286 23840 -12110
rect 23874 -12286 23880 -12110
rect 24292 -12110 24338 -12098
rect 24292 -12258 24298 -12110
rect 23834 -12298 23880 -12286
rect 24286 -12286 24298 -12258
rect 24332 -12258 24338 -12110
rect 24750 -12110 24810 -11730
rect 24332 -12286 24346 -12258
rect 24750 -12266 24756 -12110
rect 20318 -12336 20526 -12330
rect 20318 -12370 20330 -12336
rect 20514 -12370 20526 -12336
rect 20318 -12376 20526 -12370
rect 20776 -12336 20984 -12330
rect 20776 -12370 20788 -12336
rect 20972 -12370 20984 -12336
rect 20776 -12376 20984 -12370
rect 21234 -12336 21442 -12330
rect 21234 -12370 21246 -12336
rect 21430 -12370 21442 -12336
rect 21234 -12376 21442 -12370
rect 21692 -12336 21900 -12330
rect 21692 -12370 21704 -12336
rect 21888 -12370 21900 -12336
rect 21692 -12376 21900 -12370
rect 22150 -12336 22358 -12330
rect 22150 -12370 22162 -12336
rect 22346 -12370 22358 -12336
rect 22150 -12376 22358 -12370
rect 22608 -12336 22816 -12330
rect 22608 -12370 22620 -12336
rect 22804 -12370 22816 -12336
rect 22608 -12376 22816 -12370
rect 23066 -12336 23274 -12330
rect 23066 -12370 23078 -12336
rect 23262 -12370 23274 -12336
rect 23066 -12376 23274 -12370
rect 23524 -12336 23732 -12330
rect 23524 -12370 23536 -12336
rect 23720 -12370 23732 -12336
rect 23524 -12376 23732 -12370
rect 23982 -12336 24190 -12330
rect 23982 -12370 23994 -12336
rect 24178 -12370 24190 -12336
rect 23982 -12376 24190 -12370
rect 20394 -12688 20454 -12376
rect 20850 -12442 20910 -12376
rect 21306 -12442 21366 -12376
rect 21772 -12442 21832 -12376
rect 22222 -12442 22282 -12376
rect 22676 -12442 22736 -12376
rect 23138 -12442 23198 -12376
rect 23592 -12442 23652 -12376
rect 24054 -12442 24114 -12376
rect 20850 -12502 24114 -12442
rect 20856 -12622 24120 -12562
rect 20856 -12688 20916 -12622
rect 21312 -12688 21372 -12622
rect 21778 -12688 21838 -12622
rect 22228 -12688 22288 -12622
rect 22682 -12688 22742 -12622
rect 23144 -12688 23204 -12622
rect 23598 -12688 23658 -12622
rect 24060 -12688 24120 -12622
rect 20318 -12694 20526 -12688
rect 20318 -12728 20330 -12694
rect 20514 -12728 20526 -12694
rect 20318 -12734 20526 -12728
rect 20776 -12694 20984 -12688
rect 20776 -12728 20788 -12694
rect 20972 -12728 20984 -12694
rect 20776 -12734 20984 -12728
rect 21234 -12694 21442 -12688
rect 21234 -12728 21246 -12694
rect 21430 -12728 21442 -12694
rect 21234 -12734 21442 -12728
rect 21692 -12694 21900 -12688
rect 21692 -12728 21704 -12694
rect 21888 -12728 21900 -12694
rect 21692 -12734 21900 -12728
rect 22150 -12694 22358 -12688
rect 22150 -12728 22162 -12694
rect 22346 -12728 22358 -12694
rect 22150 -12734 22358 -12728
rect 22608 -12694 22816 -12688
rect 22608 -12728 22620 -12694
rect 22804 -12728 22816 -12694
rect 22608 -12734 22816 -12728
rect 23066 -12694 23274 -12688
rect 23066 -12728 23078 -12694
rect 23262 -12728 23274 -12694
rect 23066 -12734 23274 -12728
rect 23524 -12694 23732 -12688
rect 23524 -12728 23536 -12694
rect 23720 -12728 23732 -12694
rect 23524 -12734 23732 -12728
rect 23982 -12694 24190 -12688
rect 23982 -12728 23994 -12694
rect 24178 -12728 24190 -12694
rect 23982 -12734 24190 -12728
rect 19790 -12918 19796 -12814
rect 20162 -12834 20176 -12778
rect 19790 -12954 19802 -12918
rect 20170 -12926 20176 -12834
rect 19440 -13004 19648 -12998
rect 19440 -13038 19452 -13004
rect 19636 -13038 19648 -13004
rect 19440 -13044 19648 -13038
rect 19508 -13390 19568 -13044
rect 19742 -13390 19802 -12954
rect 20162 -12954 20176 -12926
rect 20210 -12834 20222 -12778
rect 20628 -12778 20674 -12766
rect 20210 -12926 20216 -12834
rect 20628 -12924 20634 -12778
rect 20210 -12954 20222 -12926
rect 20162 -13390 20222 -12954
rect 20622 -12954 20634 -12924
rect 20668 -12924 20674 -12778
rect 21086 -12778 21132 -12766
rect 20668 -12954 20682 -12924
rect 20318 -13004 20526 -12998
rect 20318 -13038 20330 -13004
rect 20514 -13038 20526 -13004
rect 20318 -13044 20526 -13038
rect 20394 -13390 20454 -13044
rect 20622 -13238 20682 -12954
rect 21086 -12954 21092 -12778
rect 21126 -12954 21132 -12778
rect 21086 -12966 21132 -12954
rect 21544 -12778 21590 -12766
rect 21544 -12954 21550 -12778
rect 21584 -12954 21590 -12778
rect 21544 -12966 21590 -12954
rect 22002 -12778 22048 -12766
rect 22002 -12954 22008 -12778
rect 22042 -12954 22048 -12778
rect 22002 -12966 22048 -12954
rect 22460 -12778 22506 -12766
rect 22460 -12954 22466 -12778
rect 22500 -12954 22506 -12778
rect 22460 -12966 22506 -12954
rect 22918 -12778 22964 -12766
rect 22918 -12954 22924 -12778
rect 22958 -12954 22964 -12778
rect 22918 -12966 22964 -12954
rect 23376 -12778 23422 -12766
rect 23376 -12954 23382 -12778
rect 23416 -12954 23422 -12778
rect 23376 -12966 23422 -12954
rect 23834 -12778 23880 -12766
rect 23834 -12954 23840 -12778
rect 23874 -12954 23880 -12778
rect 24286 -12778 24346 -12286
rect 24742 -12286 24756 -12266
rect 24790 -12140 24810 -12110
rect 24790 -12266 24796 -12140
rect 24790 -12286 24802 -12266
rect 24440 -12336 24648 -12330
rect 24440 -12370 24452 -12336
rect 24636 -12370 24648 -12336
rect 24440 -12376 24648 -12370
rect 24514 -12502 24574 -12376
rect 24742 -12502 24802 -12286
rect 24514 -12562 24802 -12502
rect 24514 -12688 24574 -12562
rect 24440 -12694 24648 -12688
rect 24440 -12728 24452 -12694
rect 24636 -12728 24648 -12694
rect 24440 -12734 24648 -12728
rect 24286 -12820 24298 -12778
rect 23834 -12966 23880 -12954
rect 24292 -12954 24298 -12820
rect 24332 -12820 24346 -12778
rect 24742 -12778 24802 -12562
rect 24742 -12818 24756 -12778
rect 24332 -12954 24338 -12820
rect 24750 -12914 24756 -12818
rect 24292 -12966 24338 -12954
rect 24742 -12954 24756 -12914
rect 24790 -12818 24802 -12778
rect 24790 -12914 24796 -12818
rect 24790 -12954 24802 -12914
rect 20776 -13004 20984 -12998
rect 20776 -13038 20788 -13004
rect 20972 -13038 20984 -13004
rect 20776 -13044 20984 -13038
rect 21234 -13004 21442 -12998
rect 21234 -13038 21246 -13004
rect 21430 -13038 21442 -13004
rect 21234 -13044 21442 -13038
rect 21692 -13004 21900 -12998
rect 21692 -13038 21704 -13004
rect 21888 -13038 21900 -13004
rect 21692 -13044 21900 -13038
rect 22150 -13004 22358 -12998
rect 22150 -13038 22162 -13004
rect 22346 -13038 22358 -13004
rect 22150 -13044 22358 -13038
rect 22608 -13004 22816 -12998
rect 22608 -13038 22620 -13004
rect 22804 -13038 22816 -13004
rect 22608 -13044 22816 -13038
rect 23066 -13004 23274 -12998
rect 23066 -13038 23078 -13004
rect 23262 -13038 23274 -13004
rect 23066 -13044 23274 -13038
rect 23524 -13004 23732 -12998
rect 23524 -13038 23536 -13004
rect 23720 -13038 23732 -13004
rect 23524 -13044 23732 -13038
rect 23982 -13004 24190 -12998
rect 23982 -13038 23994 -13004
rect 24178 -13038 24190 -13004
rect 23982 -13044 24190 -13038
rect 24440 -13004 24648 -12998
rect 24440 -13038 24452 -13004
rect 24636 -13038 24648 -13004
rect 24440 -13044 24648 -13038
rect 20850 -13110 20916 -13044
rect 21306 -13104 21372 -13044
rect 21306 -13110 21312 -13104
rect 20850 -13170 20856 -13110
rect 20916 -13164 21312 -13110
rect 21372 -13110 21378 -13104
rect 21772 -13110 21838 -13044
rect 22222 -13110 22288 -13044
rect 22676 -13110 22742 -13044
rect 23138 -13104 23204 -13044
rect 23138 -13110 23144 -13104
rect 21372 -13164 21778 -13110
rect 20916 -13170 21778 -13164
rect 21838 -13170 22228 -13110
rect 22288 -13170 22682 -13110
rect 22742 -13164 23144 -13110
rect 23204 -13110 23210 -13104
rect 23592 -13110 23658 -13044
rect 24054 -13104 24120 -13044
rect 24054 -13110 24060 -13104
rect 23204 -13164 23598 -13110
rect 22742 -13170 23598 -13164
rect 23658 -13164 24060 -13110
rect 24120 -13164 24126 -13104
rect 23658 -13170 24114 -13164
rect 20622 -13304 20682 -13298
rect 24512 -13390 24572 -13044
rect 24742 -13390 24802 -12954
rect 25110 -13266 25116 -11262
rect 25216 -13266 25222 -11262
rect 25110 -13390 25222 -13266
rect 14766 -13396 25222 -13390
rect 14766 -13496 14872 -13396
rect 25116 -13496 25222 -13396
rect 14766 -13502 25222 -13496
rect 14766 -13732 25222 -13726
rect 14766 -13832 14872 -13732
rect 25116 -13832 25222 -13732
rect 14766 -13838 25222 -13832
rect 14766 -14014 14878 -13838
rect 14766 -19186 14772 -14014
rect 14872 -15808 14878 -14014
rect 15164 -14271 15224 -13838
rect 15392 -14172 15452 -13838
rect 15622 -13912 15682 -13906
rect 15317 -14178 15525 -14172
rect 15317 -14212 15329 -14178
rect 15513 -14212 15525 -14178
rect 15317 -14218 15525 -14212
rect 15164 -14304 15175 -14271
rect 15169 -15394 15175 -14304
rect 15166 -15447 15175 -15394
rect 15209 -14304 15224 -14271
rect 15622 -14271 15682 -13972
rect 15854 -14042 15914 -14036
rect 16310 -14042 16370 -14036
rect 17226 -14042 17286 -14036
rect 15914 -14102 16310 -14044
rect 16776 -14044 16836 -14042
rect 16370 -14048 17226 -14044
rect 16370 -14102 16776 -14048
rect 15854 -14104 16776 -14102
rect 15854 -14172 15914 -14104
rect 16310 -14172 16370 -14104
rect 16836 -14102 17226 -14048
rect 17680 -14042 17740 -14036
rect 17286 -14102 17680 -14044
rect 18142 -14042 18202 -14036
rect 19058 -14040 19118 -14034
rect 17740 -14102 18142 -14044
rect 18596 -14044 18656 -14042
rect 18202 -14048 19058 -14044
rect 18202 -14102 18596 -14048
rect 16836 -14104 18596 -14102
rect 16776 -14172 16836 -14108
rect 17226 -14172 17286 -14104
rect 17680 -14172 17740 -14104
rect 18142 -14172 18202 -14104
rect 18656 -14100 19058 -14048
rect 18656 -14104 19118 -14100
rect 18596 -14172 18656 -14108
rect 19058 -14172 19118 -14104
rect 15775 -14178 15983 -14172
rect 15775 -14212 15787 -14178
rect 15971 -14212 15983 -14178
rect 15775 -14218 15983 -14212
rect 16233 -14178 16441 -14172
rect 16233 -14212 16245 -14178
rect 16429 -14212 16441 -14178
rect 16233 -14218 16441 -14212
rect 16691 -14178 16899 -14172
rect 16691 -14212 16703 -14178
rect 16887 -14212 16899 -14178
rect 16691 -14218 16899 -14212
rect 17149 -14178 17357 -14172
rect 17149 -14212 17161 -14178
rect 17345 -14212 17357 -14178
rect 17149 -14218 17357 -14212
rect 17607 -14178 17815 -14172
rect 17607 -14212 17619 -14178
rect 17803 -14212 17815 -14178
rect 17607 -14218 17815 -14212
rect 18065 -14178 18273 -14172
rect 18065 -14212 18077 -14178
rect 18261 -14212 18273 -14178
rect 18065 -14218 18273 -14212
rect 18523 -14178 18731 -14172
rect 18523 -14212 18535 -14178
rect 18719 -14212 18731 -14178
rect 18523 -14218 18731 -14212
rect 18981 -14178 19189 -14172
rect 18981 -14212 18993 -14178
rect 19177 -14212 19189 -14178
rect 18981 -14218 19189 -14212
rect 15622 -14278 15633 -14271
rect 15209 -15394 15215 -14304
rect 15209 -15447 15226 -15394
rect 15166 -15808 15226 -15447
rect 15627 -15447 15633 -14278
rect 15667 -14278 15682 -14271
rect 16085 -14271 16131 -14259
rect 15667 -15447 15673 -14278
rect 15627 -15459 15673 -15447
rect 16085 -15447 16091 -14271
rect 16125 -15447 16131 -14271
rect 16085 -15459 16131 -15447
rect 16543 -14271 16589 -14259
rect 16543 -15447 16549 -14271
rect 16583 -15447 16589 -14271
rect 16543 -15459 16589 -15447
rect 17001 -14271 17047 -14259
rect 17001 -15447 17007 -14271
rect 17041 -15447 17047 -14271
rect 17001 -15459 17047 -15447
rect 17459 -14271 17505 -14259
rect 17459 -15447 17465 -14271
rect 17499 -15447 17505 -14271
rect 17459 -15459 17505 -15447
rect 17917 -14271 17963 -14259
rect 17917 -15447 17923 -14271
rect 17957 -15447 17963 -14271
rect 17917 -15459 17963 -15447
rect 18375 -14271 18421 -14259
rect 18375 -15447 18381 -14271
rect 18415 -15447 18421 -14271
rect 18375 -15459 18421 -15447
rect 18833 -14271 18879 -14259
rect 18833 -15447 18839 -14271
rect 18873 -15447 18879 -14271
rect 19286 -14271 19346 -13838
rect 19516 -14172 19576 -13838
rect 19439 -14178 19647 -14172
rect 19439 -14212 19451 -14178
rect 19635 -14212 19647 -14178
rect 19439 -14218 19647 -14212
rect 19286 -14312 19297 -14271
rect 19291 -15404 19297 -14312
rect 18833 -15459 18879 -15447
rect 19284 -15447 19297 -15404
rect 19331 -14312 19346 -14271
rect 19744 -14271 19804 -13838
rect 19744 -14306 19755 -14271
rect 19331 -15404 19337 -14312
rect 19331 -15447 19344 -15404
rect 19749 -15426 19755 -14306
rect 15317 -15506 15525 -15500
rect 15317 -15540 15329 -15506
rect 15513 -15540 15525 -15506
rect 15317 -15546 15525 -15540
rect 15775 -15506 15983 -15500
rect 15775 -15540 15787 -15506
rect 15971 -15540 15983 -15506
rect 15775 -15546 15983 -15540
rect 16233 -15506 16441 -15500
rect 16233 -15540 16245 -15506
rect 16429 -15540 16441 -15506
rect 16233 -15546 16441 -15540
rect 16691 -15506 16899 -15500
rect 16691 -15540 16703 -15506
rect 16887 -15540 16899 -15506
rect 16691 -15546 16899 -15540
rect 17149 -15506 17357 -15500
rect 17149 -15540 17161 -15506
rect 17345 -15540 17357 -15506
rect 17149 -15546 17357 -15540
rect 17607 -15506 17815 -15500
rect 17607 -15540 17619 -15506
rect 17803 -15540 17815 -15506
rect 17607 -15546 17815 -15540
rect 18065 -15506 18273 -15500
rect 18065 -15540 18077 -15506
rect 18261 -15540 18273 -15506
rect 18065 -15546 18273 -15540
rect 18523 -15506 18731 -15500
rect 18523 -15540 18535 -15506
rect 18719 -15540 18731 -15506
rect 18523 -15546 18731 -15540
rect 18981 -15506 19189 -15500
rect 18981 -15540 18993 -15506
rect 19177 -15540 19189 -15506
rect 18981 -15546 19189 -15540
rect 15392 -15808 15452 -15546
rect 15854 -15616 15914 -15546
rect 16310 -15616 16370 -15546
rect 16776 -15616 16836 -15546
rect 17226 -15616 17286 -15546
rect 17680 -15616 17740 -15546
rect 18142 -15616 18202 -15546
rect 18596 -15616 18656 -15546
rect 19058 -15616 19118 -15546
rect 15854 -15676 19118 -15616
rect 19284 -15598 19344 -15447
rect 19742 -15447 19755 -15426
rect 19789 -14306 19804 -14271
rect 20164 -14271 20224 -13838
rect 20392 -14172 20452 -13838
rect 20616 -13978 20622 -13918
rect 20682 -13978 20688 -13918
rect 20317 -14178 20525 -14172
rect 20317 -14212 20329 -14178
rect 20513 -14212 20525 -14178
rect 20317 -14218 20525 -14212
rect 20164 -14306 20175 -14271
rect 19789 -15426 19795 -14306
rect 19789 -15447 19802 -15426
rect 20169 -15432 20175 -14306
rect 19439 -15506 19647 -15500
rect 19439 -15540 19451 -15506
rect 19635 -15540 19647 -15506
rect 19439 -15546 19647 -15540
rect 19510 -15598 19570 -15546
rect 19742 -15598 19802 -15447
rect 20162 -15447 20175 -15432
rect 20209 -14306 20224 -14271
rect 20622 -14271 20682 -13978
rect 20856 -14040 20916 -14034
rect 22228 -14038 22288 -14032
rect 21312 -14044 21372 -14038
rect 21778 -14044 21838 -14038
rect 20916 -14100 21312 -14044
rect 20856 -14104 21312 -14100
rect 21372 -14104 21778 -14044
rect 21838 -14098 22228 -14044
rect 22682 -14044 22742 -14038
rect 23144 -14044 23204 -14038
rect 23598 -14040 23658 -14034
rect 22288 -14098 22682 -14044
rect 21838 -14104 22682 -14098
rect 22742 -14104 23144 -14044
rect 23204 -14100 23598 -14044
rect 24060 -14040 24120 -14034
rect 23658 -14100 24060 -14044
rect 23204 -14104 24120 -14100
rect 20856 -14172 20916 -14104
rect 21312 -14172 21372 -14104
rect 21778 -14172 21838 -14104
rect 22228 -14172 22288 -14104
rect 22682 -14172 22742 -14104
rect 23144 -14172 23204 -14104
rect 23598 -14172 23658 -14104
rect 24060 -14172 24120 -14104
rect 24514 -14172 24574 -13838
rect 20775 -14178 20983 -14172
rect 20775 -14212 20787 -14178
rect 20971 -14212 20983 -14178
rect 20775 -14218 20983 -14212
rect 21233 -14178 21441 -14172
rect 21233 -14212 21245 -14178
rect 21429 -14212 21441 -14178
rect 21233 -14218 21441 -14212
rect 21691 -14178 21899 -14172
rect 21691 -14212 21703 -14178
rect 21887 -14212 21899 -14178
rect 21691 -14218 21899 -14212
rect 22149 -14178 22357 -14172
rect 22149 -14212 22161 -14178
rect 22345 -14212 22357 -14178
rect 22149 -14218 22357 -14212
rect 22607 -14178 22815 -14172
rect 22607 -14212 22619 -14178
rect 22803 -14212 22815 -14178
rect 22607 -14218 22815 -14212
rect 23065 -14178 23273 -14172
rect 23065 -14212 23077 -14178
rect 23261 -14212 23273 -14178
rect 23065 -14218 23273 -14212
rect 23523 -14178 23731 -14172
rect 23523 -14212 23535 -14178
rect 23719 -14212 23731 -14178
rect 23523 -14218 23731 -14212
rect 23981 -14178 24189 -14172
rect 23981 -14212 23993 -14178
rect 24177 -14212 24189 -14178
rect 23981 -14218 24189 -14212
rect 24439 -14178 24647 -14172
rect 24439 -14212 24451 -14178
rect 24635 -14212 24647 -14178
rect 24439 -14218 24647 -14212
rect 20209 -15432 20215 -14306
rect 20622 -14338 20633 -14271
rect 20209 -15447 20222 -15432
rect 20162 -15598 20222 -15447
rect 20627 -15447 20633 -14338
rect 20667 -14338 20682 -14271
rect 21085 -14271 21131 -14259
rect 20667 -15447 20673 -14338
rect 20627 -15459 20673 -15447
rect 21085 -15447 21091 -14271
rect 21125 -15447 21131 -14271
rect 21085 -15459 21131 -15447
rect 21543 -14271 21589 -14259
rect 21543 -15447 21549 -14271
rect 21583 -15447 21589 -14271
rect 21543 -15459 21589 -15447
rect 22001 -14271 22047 -14259
rect 22001 -15447 22007 -14271
rect 22041 -15447 22047 -14271
rect 22001 -15459 22047 -15447
rect 22459 -14271 22505 -14259
rect 22459 -15447 22465 -14271
rect 22499 -15447 22505 -14271
rect 22459 -15459 22505 -15447
rect 22917 -14271 22963 -14259
rect 22917 -15447 22923 -14271
rect 22957 -15447 22963 -14271
rect 22917 -15459 22963 -15447
rect 23375 -14271 23421 -14259
rect 23375 -15447 23381 -14271
rect 23415 -15447 23421 -14271
rect 23375 -15459 23421 -15447
rect 23833 -14271 23879 -14259
rect 23833 -15447 23839 -14271
rect 23873 -15447 23879 -14271
rect 24291 -14271 24337 -14259
rect 24291 -15380 24297 -14271
rect 23833 -15459 23879 -15447
rect 24284 -15447 24297 -15380
rect 24331 -15380 24337 -14271
rect 24742 -14271 24802 -13838
rect 24742 -14292 24755 -14271
rect 24331 -15447 24344 -15380
rect 24749 -15400 24755 -14292
rect 20317 -15506 20525 -15500
rect 20317 -15540 20329 -15506
rect 20513 -15540 20525 -15506
rect 20317 -15546 20525 -15540
rect 20775 -15506 20983 -15500
rect 20775 -15540 20787 -15506
rect 20971 -15540 20983 -15506
rect 20775 -15546 20983 -15540
rect 21233 -15506 21441 -15500
rect 21233 -15540 21245 -15506
rect 21429 -15540 21441 -15506
rect 21233 -15546 21441 -15540
rect 21691 -15506 21899 -15500
rect 21691 -15540 21703 -15506
rect 21887 -15540 21899 -15506
rect 21691 -15546 21899 -15540
rect 22149 -15506 22357 -15500
rect 22149 -15540 22161 -15506
rect 22345 -15540 22357 -15506
rect 22149 -15546 22357 -15540
rect 22607 -15506 22815 -15500
rect 22607 -15540 22619 -15506
rect 22803 -15540 22815 -15506
rect 22607 -15546 22815 -15540
rect 23065 -15506 23273 -15500
rect 23065 -15540 23077 -15506
rect 23261 -15540 23273 -15506
rect 23065 -15546 23273 -15540
rect 23523 -15506 23731 -15500
rect 23523 -15540 23535 -15506
rect 23719 -15540 23731 -15506
rect 23523 -15546 23731 -15540
rect 23981 -15506 24189 -15500
rect 23981 -15540 23993 -15506
rect 24177 -15540 24189 -15506
rect 23981 -15546 24189 -15540
rect 20392 -15598 20452 -15546
rect 19284 -15658 20452 -15598
rect 20848 -15616 20908 -15546
rect 21304 -15616 21364 -15546
rect 21770 -15616 21830 -15546
rect 22220 -15616 22280 -15546
rect 22674 -15616 22734 -15546
rect 23136 -15616 23196 -15546
rect 23590 -15616 23650 -15546
rect 24052 -15616 24112 -15546
rect 20848 -15676 24112 -15616
rect 24284 -15718 24344 -15447
rect 24742 -15447 24755 -15400
rect 24789 -14292 24802 -14271
rect 25110 -14014 25222 -13838
rect 24789 -15400 24795 -14292
rect 24789 -15447 24802 -15400
rect 24439 -15506 24647 -15500
rect 24439 -15540 24451 -15506
rect 24635 -15540 24647 -15506
rect 24439 -15546 24647 -15540
rect 24278 -15778 24284 -15718
rect 24344 -15778 24350 -15718
rect 14872 -15868 16002 -15808
rect 14872 -16302 14878 -15868
rect 15942 -16302 16002 -15868
rect 16854 -15884 23330 -15824
rect 24514 -15872 24574 -15546
rect 24742 -15872 24802 -15447
rect 25110 -15872 25116 -14014
rect 14872 -16362 16460 -16302
rect 14872 -19186 14878 -16362
rect 15942 -16536 16002 -16362
rect 16168 -16437 16228 -16362
rect 16094 -16443 16302 -16437
rect 16094 -16477 16106 -16443
rect 16290 -16477 16302 -16443
rect 16094 -16483 16302 -16477
rect 15942 -16580 15952 -16536
rect 15946 -18042 15952 -16580
rect 15938 -18112 15952 -18042
rect 15986 -16580 16002 -16536
rect 16400 -16536 16460 -16362
rect 16624 -16364 16630 -16304
rect 16690 -16364 16696 -16304
rect 16630 -16437 16690 -16364
rect 16552 -16443 16760 -16437
rect 16552 -16477 16564 -16443
rect 16748 -16477 16760 -16443
rect 16552 -16483 16760 -16477
rect 15986 -18042 15992 -16580
rect 16400 -16598 16410 -16536
rect 16404 -18036 16410 -16598
rect 15986 -18112 15998 -18042
rect 15938 -18900 15998 -18112
rect 16396 -18112 16410 -18036
rect 16444 -16598 16460 -16536
rect 16854 -16536 16914 -15884
rect 17768 -16014 22412 -15954
rect 17084 -16364 17090 -16304
rect 17150 -16364 17156 -16304
rect 17542 -16364 17548 -16304
rect 17608 -16364 17614 -16304
rect 17090 -16437 17150 -16364
rect 17548 -16437 17608 -16364
rect 17010 -16443 17218 -16437
rect 17010 -16477 17022 -16443
rect 17206 -16477 17218 -16443
rect 17010 -16483 17218 -16477
rect 17468 -16443 17676 -16437
rect 17468 -16477 17480 -16443
rect 17664 -16477 17676 -16443
rect 17468 -16483 17676 -16477
rect 16854 -16596 16868 -16536
rect 16444 -18036 16450 -16598
rect 16444 -18112 16456 -18036
rect 16094 -18171 16302 -18165
rect 16094 -18205 16106 -18171
rect 16290 -18205 16302 -18171
rect 16094 -18211 16302 -18205
rect 16166 -18900 16226 -18211
rect 16396 -18900 16456 -18112
rect 16862 -18112 16868 -16596
rect 16902 -16596 16914 -16536
rect 17320 -16536 17366 -16524
rect 16902 -18112 16908 -16596
rect 17320 -18056 17326 -16536
rect 16862 -18124 16908 -18112
rect 17312 -18112 17326 -18056
rect 17360 -18056 17366 -16536
rect 17768 -16536 17828 -16014
rect 18688 -16140 21504 -16080
rect 17998 -16364 18004 -16304
rect 18064 -16364 18070 -16304
rect 18454 -16364 18460 -16304
rect 18520 -16364 18526 -16304
rect 18004 -16437 18064 -16364
rect 18460 -16437 18520 -16364
rect 17926 -16443 18134 -16437
rect 17926 -16477 17938 -16443
rect 18122 -16477 18134 -16443
rect 17926 -16483 18134 -16477
rect 18384 -16443 18592 -16437
rect 18384 -16477 18396 -16443
rect 18580 -16477 18592 -16443
rect 18384 -16483 18592 -16477
rect 17768 -16604 17784 -16536
rect 17360 -18112 17372 -18056
rect 16552 -18171 16760 -18165
rect 16552 -18205 16564 -18171
rect 16748 -18205 16760 -18171
rect 16552 -18211 16760 -18205
rect 17010 -18171 17218 -18165
rect 17010 -18205 17022 -18171
rect 17206 -18205 17218 -18171
rect 17010 -18211 17218 -18205
rect 16626 -18278 16686 -18211
rect 17086 -18278 17146 -18211
rect 16620 -18338 16626 -18278
rect 16686 -18338 16692 -18278
rect 17080 -18338 17086 -18278
rect 17146 -18338 17152 -18278
rect 17312 -18646 17372 -18112
rect 17778 -18112 17784 -16604
rect 17818 -16604 17828 -16536
rect 18236 -16536 18282 -16524
rect 17818 -18112 17824 -16604
rect 18236 -18054 18242 -16536
rect 17778 -18124 17824 -18112
rect 18232 -18112 18242 -18054
rect 18276 -18054 18282 -16536
rect 18688 -16536 18748 -16140
rect 19602 -16256 20580 -16196
rect 18910 -16364 18916 -16304
rect 18976 -16364 18982 -16304
rect 19370 -16364 19376 -16304
rect 19436 -16364 19442 -16304
rect 18916 -16437 18976 -16364
rect 19376 -16437 19436 -16364
rect 18842 -16443 19050 -16437
rect 18842 -16477 18854 -16443
rect 19038 -16477 19050 -16443
rect 18842 -16483 19050 -16477
rect 19300 -16443 19508 -16437
rect 19300 -16477 19312 -16443
rect 19496 -16477 19508 -16443
rect 19300 -16483 19508 -16477
rect 18688 -16568 18700 -16536
rect 18276 -18112 18292 -18054
rect 17468 -18171 17676 -18165
rect 17468 -18205 17480 -18171
rect 17664 -18205 17676 -18171
rect 17468 -18211 17676 -18205
rect 17926 -18171 18134 -18165
rect 17926 -18205 17938 -18171
rect 18122 -18205 18134 -18171
rect 17926 -18211 18134 -18205
rect 17544 -18278 17604 -18211
rect 18000 -18278 18060 -18211
rect 17538 -18338 17544 -18278
rect 17604 -18338 17610 -18278
rect 17994 -18338 18000 -18278
rect 18060 -18338 18066 -18278
rect 18232 -18512 18292 -18112
rect 18694 -18112 18700 -16568
rect 18734 -16568 18748 -16536
rect 19152 -16536 19198 -16524
rect 18734 -18112 18740 -16568
rect 19152 -18068 19158 -16536
rect 18694 -18124 18740 -18112
rect 19148 -18112 19158 -18068
rect 19192 -18068 19198 -16536
rect 19602 -16536 19662 -16256
rect 19820 -16304 19904 -16300
rect 19820 -16366 19832 -16304
rect 19892 -16366 19904 -16304
rect 19820 -16372 19904 -16366
rect 20058 -16316 20118 -16310
rect 19832 -16437 19892 -16372
rect 20286 -16364 20292 -16304
rect 20352 -16364 20358 -16304
rect 20286 -16366 20358 -16364
rect 19758 -16443 19966 -16437
rect 19758 -16477 19770 -16443
rect 19954 -16477 19966 -16443
rect 19758 -16483 19966 -16477
rect 19602 -16564 19616 -16536
rect 19192 -18112 19208 -18068
rect 18384 -18171 18592 -18165
rect 18384 -18205 18396 -18171
rect 18580 -18205 18592 -18171
rect 18384 -18211 18592 -18205
rect 18842 -18171 19050 -18165
rect 18842 -18205 18854 -18171
rect 19038 -18205 19050 -18171
rect 18842 -18211 19050 -18205
rect 18456 -18278 18516 -18211
rect 18912 -18278 18972 -18211
rect 18450 -18338 18456 -18278
rect 18516 -18338 18522 -18278
rect 18906 -18338 18912 -18278
rect 18972 -18338 18978 -18278
rect 19148 -18388 19208 -18112
rect 19610 -18112 19616 -16564
rect 19650 -16564 19662 -16536
rect 20058 -16536 20118 -16376
rect 20292 -16437 20352 -16366
rect 20216 -16443 20424 -16437
rect 20216 -16477 20228 -16443
rect 20412 -16477 20424 -16443
rect 20216 -16483 20424 -16477
rect 20058 -16558 20074 -16536
rect 19650 -18112 19656 -16564
rect 19610 -18124 19656 -18112
rect 20068 -18112 20074 -16558
rect 20108 -16558 20118 -16536
rect 20520 -16536 20580 -16256
rect 20744 -16364 20750 -16304
rect 20810 -16364 20816 -16304
rect 21198 -16364 21204 -16304
rect 21264 -16364 21270 -16304
rect 20750 -16437 20810 -16364
rect 21204 -16437 21264 -16364
rect 20674 -16443 20882 -16437
rect 20674 -16477 20686 -16443
rect 20870 -16477 20882 -16443
rect 20674 -16483 20882 -16477
rect 21132 -16443 21340 -16437
rect 21132 -16477 21144 -16443
rect 21328 -16477 21340 -16443
rect 21132 -16483 21340 -16477
rect 21444 -16524 21504 -16140
rect 21662 -16364 21668 -16304
rect 21728 -16364 21734 -16304
rect 22120 -16364 22126 -16304
rect 22186 -16364 22192 -16304
rect 21668 -16437 21728 -16364
rect 22126 -16437 22186 -16364
rect 21590 -16443 21798 -16437
rect 21590 -16477 21602 -16443
rect 21786 -16477 21798 -16443
rect 21590 -16483 21798 -16477
rect 22048 -16443 22256 -16437
rect 22048 -16477 22060 -16443
rect 22244 -16477 22256 -16443
rect 22048 -16483 22256 -16477
rect 20108 -18112 20114 -16558
rect 20520 -16616 20532 -16536
rect 20068 -18124 20114 -18112
rect 20526 -18112 20532 -16616
rect 20566 -16616 20580 -16536
rect 20984 -16536 21030 -16524
rect 20566 -18112 20572 -16616
rect 20984 -18034 20990 -16536
rect 20526 -18124 20572 -18112
rect 20978 -18112 20990 -18034
rect 21024 -18034 21030 -16536
rect 21442 -16536 21504 -16524
rect 21024 -18112 21038 -18034
rect 19300 -18171 19508 -18165
rect 19300 -18205 19312 -18171
rect 19496 -18205 19508 -18171
rect 19300 -18211 19508 -18205
rect 19758 -18171 19966 -18165
rect 19758 -18205 19770 -18171
rect 19954 -18205 19966 -18171
rect 19758 -18211 19966 -18205
rect 20216 -18171 20424 -18165
rect 20216 -18205 20228 -18171
rect 20412 -18205 20424 -18171
rect 20216 -18211 20424 -18205
rect 20674 -18171 20882 -18165
rect 20674 -18205 20686 -18171
rect 20870 -18205 20882 -18171
rect 20674 -18211 20882 -18205
rect 19368 -18278 19428 -18211
rect 19826 -18278 19886 -18211
rect 20294 -18278 20354 -18211
rect 20750 -18278 20810 -18211
rect 19362 -18338 19368 -18278
rect 19428 -18338 19434 -18278
rect 19820 -18338 19826 -18278
rect 19886 -18338 19892 -18278
rect 20288 -18338 20294 -18278
rect 20354 -18338 20360 -18278
rect 20744 -18338 20750 -18278
rect 20810 -18338 20816 -18278
rect 20978 -18388 21038 -18112
rect 21442 -18112 21448 -16536
rect 21482 -16608 21504 -16536
rect 21900 -16536 21946 -16524
rect 21482 -18112 21488 -16608
rect 21900 -18052 21906 -16536
rect 21442 -18124 21488 -18112
rect 21894 -18112 21906 -18052
rect 21940 -18052 21946 -16536
rect 22352 -16536 22412 -16014
rect 22576 -16364 22582 -16304
rect 22642 -16364 22648 -16304
rect 23036 -16364 23042 -16304
rect 23102 -16364 23108 -16304
rect 22582 -16437 22642 -16364
rect 23042 -16437 23102 -16364
rect 22506 -16443 22714 -16437
rect 22506 -16477 22518 -16443
rect 22702 -16477 22714 -16443
rect 22506 -16483 22714 -16477
rect 22964 -16443 23172 -16437
rect 22964 -16477 22976 -16443
rect 23160 -16477 23172 -16443
rect 22964 -16483 23172 -16477
rect 22352 -16614 22364 -16536
rect 21940 -18112 21954 -18052
rect 21132 -18171 21340 -18165
rect 21132 -18205 21144 -18171
rect 21328 -18205 21340 -18171
rect 21132 -18211 21340 -18205
rect 21590 -18171 21798 -18165
rect 21590 -18205 21602 -18171
rect 21786 -18205 21798 -18171
rect 21590 -18211 21798 -18205
rect 21200 -18278 21260 -18211
rect 21664 -18278 21724 -18211
rect 21194 -18338 21200 -18278
rect 21260 -18338 21266 -18278
rect 21658 -18338 21664 -18278
rect 21724 -18338 21730 -18278
rect 19148 -18448 21038 -18388
rect 21894 -18512 21954 -18112
rect 22358 -18112 22364 -16614
rect 22398 -16614 22412 -16536
rect 22816 -16536 22862 -16524
rect 22398 -18112 22404 -16614
rect 22816 -18054 22822 -16536
rect 22358 -18124 22404 -18112
rect 22810 -18112 22822 -18054
rect 22856 -18054 22862 -16536
rect 23270 -16536 23330 -15884
rect 24182 -15932 25116 -15872
rect 24182 -16304 24242 -15932
rect 25110 -16304 25116 -15932
rect 23492 -16364 23498 -16304
rect 23558 -16364 23564 -16304
rect 23728 -16364 25116 -16304
rect 23498 -16437 23558 -16364
rect 23422 -16443 23630 -16437
rect 23422 -16477 23434 -16443
rect 23618 -16477 23630 -16443
rect 23422 -16483 23630 -16477
rect 23270 -16620 23280 -16536
rect 22856 -18112 22870 -18054
rect 22048 -18171 22256 -18165
rect 22048 -18205 22060 -18171
rect 22244 -18205 22256 -18171
rect 22048 -18211 22256 -18205
rect 22506 -18171 22714 -18165
rect 22506 -18205 22518 -18171
rect 22702 -18205 22714 -18171
rect 22506 -18211 22714 -18205
rect 22122 -18278 22182 -18211
rect 22578 -18278 22638 -18211
rect 22116 -18338 22122 -18278
rect 22182 -18338 22188 -18278
rect 22572 -18338 22578 -18278
rect 22638 -18338 22644 -18278
rect 18232 -18572 21954 -18512
rect 22810 -18646 22870 -18112
rect 23274 -18112 23280 -16620
rect 23314 -16620 23330 -16536
rect 23728 -16536 23788 -16364
rect 23954 -16437 24014 -16364
rect 23880 -16443 24088 -16437
rect 23880 -16477 23892 -16443
rect 24076 -16477 24088 -16443
rect 23880 -16483 24088 -16477
rect 23728 -16580 23738 -16536
rect 23314 -18112 23320 -16620
rect 23732 -18048 23738 -16580
rect 23274 -18124 23320 -18112
rect 23726 -18112 23738 -18048
rect 23772 -16580 23788 -16536
rect 24182 -16536 24242 -16364
rect 23772 -18048 23778 -16580
rect 24182 -16596 24196 -16536
rect 23772 -18112 23786 -18048
rect 24190 -18080 24196 -16596
rect 22964 -18171 23172 -18165
rect 22964 -18205 22976 -18171
rect 23160 -18205 23172 -18171
rect 22964 -18211 23172 -18205
rect 23422 -18171 23630 -18165
rect 23422 -18205 23434 -18171
rect 23618 -18205 23630 -18171
rect 23422 -18211 23630 -18205
rect 23038 -18278 23098 -18211
rect 23494 -18278 23554 -18211
rect 23032 -18338 23038 -18278
rect 23098 -18338 23104 -18278
rect 23488 -18338 23494 -18278
rect 23554 -18338 23560 -18278
rect 17312 -18706 22870 -18646
rect 23726 -18900 23786 -18112
rect 24184 -18112 24196 -18080
rect 24230 -16596 24242 -16536
rect 24230 -18080 24236 -16596
rect 24230 -18112 24244 -18080
rect 23880 -18171 24088 -18165
rect 23880 -18205 23892 -18171
rect 24076 -18205 24088 -18171
rect 23880 -18211 24088 -18205
rect 23952 -18900 24012 -18211
rect 24184 -18900 24244 -18112
rect 15916 -18910 24272 -18900
rect 15916 -18996 15942 -18910
rect 16038 -18996 16362 -18910
rect 16458 -18996 16962 -18910
rect 17058 -18996 17562 -18910
rect 17658 -18996 18162 -18910
rect 18258 -18996 18762 -18910
rect 18858 -18996 19362 -18910
rect 19458 -18996 19962 -18910
rect 20058 -18996 20562 -18910
rect 20658 -18996 21162 -18910
rect 21258 -18996 21762 -18910
rect 21858 -18996 22362 -18910
rect 22458 -18996 22962 -18910
rect 23058 -18996 23562 -18910
rect 23658 -18996 24162 -18910
rect 24258 -18996 24272 -18910
rect 15916 -19010 24272 -18996
rect 14766 -19470 14878 -19186
rect 15478 -19470 15488 -19170
rect 24500 -19470 24510 -19170
rect 25110 -19186 25116 -16364
rect 25216 -19186 25222 -14014
rect 25110 -19470 25222 -19186
rect 14766 -19476 25222 -19470
rect 14766 -19576 14872 -19476
rect 25116 -19576 25222 -19476
rect 14766 -19582 25222 -19576
rect 25406 -16304 25466 -3332
rect 25546 -9650 25606 2140
rect 26002 2194 31458 2200
rect 26002 2094 26108 2194
rect 31352 2094 31458 2194
rect 26002 2088 31458 2094
rect 26002 1911 26114 2088
rect 26002 -982 26008 1911
rect 26000 -1092 26008 -982
rect 26002 -1375 26008 -1092
rect 26108 420 26114 1911
rect 26384 1801 26444 2088
rect 26612 1900 26672 2088
rect 26539 1894 26747 1900
rect 26539 1860 26551 1894
rect 26735 1860 26747 1894
rect 26539 1854 26747 1860
rect 26384 1778 26397 1801
rect 26391 670 26397 1778
rect 26384 625 26397 670
rect 26431 1778 26444 1801
rect 26842 1801 26902 2088
rect 30504 2032 30564 2038
rect 27066 2026 27126 2032
rect 27528 2026 27588 2032
rect 27982 2026 28042 2032
rect 28444 2026 28504 2032
rect 28898 2026 28958 2032
rect 29348 2026 29408 2032
rect 29814 2026 29874 2032
rect 30270 2026 30330 2032
rect 27060 1966 27066 2026
rect 27126 1966 27528 2026
rect 27588 1966 27982 2026
rect 28042 1966 28444 2026
rect 28504 1966 28898 2026
rect 28958 1966 29348 2026
rect 29408 1966 29814 2026
rect 29874 1966 30270 2026
rect 30330 1966 30336 2026
rect 27066 1900 27126 1966
rect 27528 1900 27588 1966
rect 27982 1900 28042 1966
rect 28444 1900 28504 1966
rect 28898 1900 28958 1966
rect 29348 1900 29408 1966
rect 29814 1900 29874 1966
rect 30270 1900 30330 1966
rect 26997 1894 27205 1900
rect 26997 1860 27009 1894
rect 27193 1860 27205 1894
rect 26997 1854 27205 1860
rect 27455 1894 27663 1900
rect 27455 1860 27467 1894
rect 27651 1860 27663 1894
rect 27455 1854 27663 1860
rect 27913 1894 28121 1900
rect 27913 1860 27925 1894
rect 28109 1860 28121 1894
rect 27913 1854 28121 1860
rect 28371 1894 28579 1900
rect 28371 1860 28383 1894
rect 28567 1860 28579 1894
rect 28371 1854 28579 1860
rect 28829 1894 29037 1900
rect 28829 1860 28841 1894
rect 29025 1860 29037 1894
rect 28829 1854 29037 1860
rect 29287 1894 29495 1900
rect 29287 1860 29299 1894
rect 29483 1860 29495 1894
rect 29287 1854 29495 1860
rect 29745 1894 29953 1900
rect 29745 1860 29757 1894
rect 29941 1860 29953 1894
rect 29745 1854 29953 1860
rect 30203 1894 30411 1900
rect 30203 1860 30215 1894
rect 30399 1860 30411 1894
rect 30203 1854 30411 1860
rect 26431 670 26437 1778
rect 26431 625 26444 670
rect 26384 420 26444 625
rect 26842 625 26855 1801
rect 26889 625 26902 1801
rect 26539 566 26747 572
rect 26539 532 26551 566
rect 26735 532 26747 566
rect 26539 526 26747 532
rect 26612 420 26672 526
rect 26842 420 26902 625
rect 27307 1801 27353 1813
rect 27307 625 27313 1801
rect 27347 625 27353 1801
rect 27307 613 27353 625
rect 27765 1801 27811 1813
rect 27765 625 27771 1801
rect 27805 625 27811 1801
rect 27765 613 27811 625
rect 28223 1801 28269 1813
rect 28223 625 28229 1801
rect 28263 625 28269 1801
rect 28223 613 28269 625
rect 28681 1801 28727 1813
rect 28681 625 28687 1801
rect 28721 625 28727 1801
rect 28681 613 28727 625
rect 29139 1801 29185 1813
rect 29139 625 29145 1801
rect 29179 625 29185 1801
rect 29139 613 29185 625
rect 29597 1801 29643 1813
rect 29597 625 29603 1801
rect 29637 625 29643 1801
rect 29597 613 29643 625
rect 30055 1801 30101 1813
rect 30055 625 30061 1801
rect 30095 625 30101 1801
rect 30504 1801 30564 1972
rect 30734 1900 30794 2088
rect 30661 1894 30869 1900
rect 30661 1860 30673 1894
rect 30857 1860 30869 1894
rect 30661 1854 30869 1860
rect 30504 1732 30519 1801
rect 30055 613 30101 625
rect 30513 625 30519 1732
rect 30553 1732 30564 1801
rect 30962 1801 31022 2088
rect 30962 1764 30977 1801
rect 30553 625 30559 1732
rect 30971 638 30977 1764
rect 30513 613 30559 625
rect 30964 625 30977 638
rect 31011 1764 31022 1801
rect 31346 1994 31458 2088
rect 31346 1963 32278 1994
rect 31346 1929 31571 1963
rect 31605 1929 31663 1963
rect 31697 1929 31755 1963
rect 31789 1929 31847 1963
rect 31881 1929 31939 1963
rect 31973 1929 32031 1963
rect 32065 1929 32123 1963
rect 32157 1929 32215 1963
rect 32249 1929 32278 1963
rect 31346 1911 32278 1929
rect 31011 638 31017 1764
rect 31011 625 31024 638
rect 26997 566 27205 572
rect 26997 532 27009 566
rect 27193 532 27205 566
rect 26997 526 27205 532
rect 27455 566 27663 572
rect 27455 532 27467 566
rect 27651 532 27663 566
rect 27455 526 27663 532
rect 27913 566 28121 572
rect 27913 532 27925 566
rect 28109 532 28121 566
rect 27913 526 28121 532
rect 28371 566 28579 572
rect 28371 532 28383 566
rect 28567 532 28579 566
rect 28371 526 28579 532
rect 28829 566 29037 572
rect 28829 532 28841 566
rect 29025 532 29037 566
rect 28829 526 29037 532
rect 29287 566 29495 572
rect 29287 532 29299 566
rect 29483 532 29495 566
rect 29287 526 29495 532
rect 29745 566 29953 572
rect 29745 532 29757 566
rect 29941 532 29953 566
rect 29745 526 29953 532
rect 30203 566 30411 572
rect 30203 532 30215 566
rect 30399 532 30411 566
rect 30203 526 30411 532
rect 30661 566 30869 572
rect 30661 532 30673 566
rect 30857 532 30869 566
rect 30661 526 30869 532
rect 26108 360 26902 420
rect 27074 454 27134 526
rect 27536 454 27596 526
rect 27990 454 28050 526
rect 28452 454 28512 526
rect 28906 454 28966 526
rect 29356 454 29416 526
rect 29822 454 29882 526
rect 30278 454 30338 526
rect 30734 472 30794 526
rect 30964 472 31024 625
rect 31346 472 31352 1911
rect 27074 394 30278 454
rect 30338 394 30344 454
rect 30734 412 31352 472
rect 26108 -982 26114 360
rect 26384 -982 26444 360
rect 26612 -982 26672 360
rect 26842 -982 26902 360
rect 30734 -982 30794 412
rect 30964 -982 31024 412
rect 26108 -992 31274 -982
rect 26108 -1078 26290 -992
rect 26386 -1078 26890 -992
rect 26986 -1078 27490 -992
rect 27586 -1078 28090 -992
rect 28186 -1078 28690 -992
rect 28786 -1078 29290 -992
rect 29386 -1078 29890 -992
rect 29986 -1078 30490 -992
rect 30586 -1078 31090 -992
rect 31186 -1078 31274 -992
rect 26108 -1092 31274 -1078
rect 26108 -1375 26114 -1092
rect 26002 -1552 26114 -1375
rect 26714 -1552 26724 -1252
rect 30736 -1552 30746 -1252
rect 31346 -1375 31352 412
rect 31452 1898 32278 1911
rect 31452 -1375 31458 1898
rect 31346 -1552 31458 -1375
rect 26002 -1558 31458 -1552
rect 26002 -1658 26108 -1558
rect 31352 -1658 31458 -1558
rect 26002 -1664 31458 -1658
rect 25812 -2028 36268 -2022
rect 25812 -2128 25918 -2028
rect 36162 -2128 36268 -2028
rect 25812 -2134 36268 -2128
rect 25812 -2418 25924 -2134
rect 25812 -7590 25818 -2418
rect 25918 -5240 25924 -2418
rect 26524 -2434 26534 -2134
rect 35546 -2434 35556 -2134
rect 36156 -2418 36268 -2134
rect 26762 -2608 35118 -2594
rect 26762 -2694 26776 -2608
rect 26872 -2694 27376 -2608
rect 27472 -2694 27976 -2608
rect 28072 -2694 28576 -2608
rect 28672 -2694 29176 -2608
rect 29272 -2694 29776 -2608
rect 29872 -2694 30376 -2608
rect 30472 -2694 30976 -2608
rect 31072 -2694 31576 -2608
rect 31672 -2694 32176 -2608
rect 32272 -2694 32776 -2608
rect 32872 -2694 33376 -2608
rect 33472 -2694 33976 -2608
rect 34072 -2694 34576 -2608
rect 34672 -2694 34996 -2608
rect 35092 -2694 35118 -2608
rect 26762 -2704 35118 -2694
rect 26790 -3492 26850 -2704
rect 27022 -3393 27082 -2704
rect 26946 -3399 27154 -3393
rect 26946 -3433 26958 -3399
rect 27142 -3433 27154 -3399
rect 26946 -3439 27154 -3433
rect 26790 -3524 26804 -3492
rect 26798 -5008 26804 -3524
rect 26792 -5068 26804 -5008
rect 26838 -3524 26850 -3492
rect 27248 -3492 27308 -2704
rect 28164 -2958 33722 -2898
rect 27474 -3326 27480 -3266
rect 27540 -3326 27546 -3266
rect 27930 -3326 27936 -3266
rect 27996 -3326 28002 -3266
rect 27480 -3393 27540 -3326
rect 27936 -3393 27996 -3326
rect 27404 -3399 27612 -3393
rect 27404 -3433 27416 -3399
rect 27600 -3433 27612 -3399
rect 27404 -3439 27612 -3433
rect 27862 -3399 28070 -3393
rect 27862 -3433 27874 -3399
rect 28058 -3433 28070 -3399
rect 27862 -3439 28070 -3433
rect 26838 -5008 26844 -3524
rect 27248 -3556 27262 -3492
rect 26838 -5068 26852 -5008
rect 27256 -5024 27262 -3556
rect 26792 -5240 26852 -5068
rect 27246 -5068 27262 -5024
rect 27296 -3556 27308 -3492
rect 27714 -3492 27760 -3480
rect 27296 -5024 27302 -3556
rect 27714 -4984 27720 -3492
rect 27296 -5068 27306 -5024
rect 26946 -5127 27154 -5121
rect 26946 -5161 26958 -5127
rect 27142 -5161 27154 -5127
rect 26946 -5167 27154 -5161
rect 27020 -5240 27080 -5167
rect 27246 -5240 27306 -5068
rect 27704 -5068 27720 -4984
rect 27754 -4984 27760 -3492
rect 28164 -3492 28224 -2958
rect 29080 -3092 32802 -3032
rect 28390 -3326 28396 -3266
rect 28456 -3326 28462 -3266
rect 28846 -3326 28852 -3266
rect 28912 -3326 28918 -3266
rect 28396 -3393 28456 -3326
rect 28852 -3393 28912 -3326
rect 28320 -3399 28528 -3393
rect 28320 -3433 28332 -3399
rect 28516 -3433 28528 -3399
rect 28320 -3439 28528 -3433
rect 28778 -3399 28986 -3393
rect 28778 -3433 28790 -3399
rect 28974 -3433 28986 -3399
rect 28778 -3439 28986 -3433
rect 28164 -3550 28178 -3492
rect 27754 -5068 27764 -4984
rect 27404 -5127 27612 -5121
rect 27404 -5161 27416 -5127
rect 27600 -5161 27612 -5127
rect 27404 -5167 27612 -5161
rect 27476 -5240 27536 -5167
rect 25918 -5300 27306 -5240
rect 27470 -5300 27476 -5240
rect 27536 -5300 27542 -5240
rect 25918 -5672 25924 -5300
rect 26792 -5672 26852 -5300
rect 25918 -5732 26852 -5672
rect 27704 -5720 27764 -5068
rect 28172 -5068 28178 -3550
rect 28212 -3550 28224 -3492
rect 28630 -3492 28676 -3480
rect 28212 -5068 28218 -3550
rect 28630 -4990 28636 -3492
rect 28172 -5080 28218 -5068
rect 28622 -5068 28636 -4990
rect 28670 -4990 28676 -3492
rect 29080 -3492 29140 -3092
rect 29996 -3216 31886 -3156
rect 29304 -3326 29310 -3266
rect 29370 -3326 29376 -3266
rect 29768 -3326 29774 -3266
rect 29834 -3326 29840 -3266
rect 29310 -3393 29370 -3326
rect 29774 -3393 29834 -3326
rect 29236 -3399 29444 -3393
rect 29236 -3433 29248 -3399
rect 29432 -3433 29444 -3399
rect 29236 -3439 29444 -3433
rect 29694 -3399 29902 -3393
rect 29694 -3433 29706 -3399
rect 29890 -3433 29902 -3399
rect 29694 -3439 29902 -3433
rect 29080 -3552 29094 -3492
rect 28670 -5068 28682 -4990
rect 27862 -5127 28070 -5121
rect 27862 -5161 27874 -5127
rect 28058 -5161 28070 -5127
rect 27862 -5167 28070 -5161
rect 28320 -5127 28528 -5121
rect 28320 -5161 28332 -5127
rect 28516 -5161 28528 -5127
rect 28320 -5167 28528 -5161
rect 27932 -5240 27992 -5167
rect 28392 -5240 28452 -5167
rect 27926 -5300 27932 -5240
rect 27992 -5300 27998 -5240
rect 28386 -5300 28392 -5240
rect 28452 -5300 28458 -5240
rect 28622 -5590 28682 -5068
rect 29088 -5068 29094 -3552
rect 29128 -3552 29140 -3492
rect 29546 -3492 29592 -3480
rect 29128 -5068 29134 -3552
rect 29546 -4996 29552 -3492
rect 29088 -5080 29134 -5068
rect 29530 -5068 29552 -4996
rect 29586 -5068 29592 -3492
rect 29996 -3492 30056 -3216
rect 30218 -3326 30224 -3266
rect 30284 -3326 30290 -3266
rect 30674 -3326 30680 -3266
rect 30740 -3326 30746 -3266
rect 31142 -3326 31148 -3266
rect 31208 -3326 31214 -3266
rect 31600 -3326 31606 -3266
rect 31666 -3326 31672 -3266
rect 30224 -3393 30284 -3326
rect 30680 -3393 30740 -3326
rect 31148 -3393 31208 -3326
rect 31606 -3393 31666 -3326
rect 30152 -3399 30360 -3393
rect 30152 -3433 30164 -3399
rect 30348 -3433 30360 -3399
rect 30152 -3439 30360 -3433
rect 30610 -3399 30818 -3393
rect 30610 -3433 30622 -3399
rect 30806 -3433 30818 -3399
rect 30610 -3439 30818 -3433
rect 31068 -3399 31276 -3393
rect 31068 -3433 31080 -3399
rect 31264 -3433 31276 -3399
rect 31068 -3439 31276 -3433
rect 31526 -3399 31734 -3393
rect 31526 -3433 31538 -3399
rect 31722 -3433 31734 -3399
rect 31526 -3439 31734 -3433
rect 29996 -3570 30010 -3492
rect 29530 -5080 29592 -5068
rect 30004 -5068 30010 -3570
rect 30044 -3570 30056 -3492
rect 30462 -3492 30508 -3480
rect 30044 -5068 30050 -3570
rect 30462 -4988 30468 -3492
rect 30004 -5080 30050 -5068
rect 30454 -5068 30468 -4988
rect 30502 -4988 30508 -3492
rect 30920 -3492 30966 -3480
rect 30502 -5068 30514 -4988
rect 30920 -5046 30926 -3492
rect 28778 -5127 28986 -5121
rect 28778 -5161 28790 -5127
rect 28974 -5161 28986 -5127
rect 28778 -5167 28986 -5161
rect 29236 -5127 29444 -5121
rect 29236 -5161 29248 -5127
rect 29432 -5161 29444 -5127
rect 29236 -5167 29444 -5161
rect 28848 -5240 28908 -5167
rect 29306 -5240 29366 -5167
rect 28842 -5300 28848 -5240
rect 28908 -5300 28914 -5240
rect 29300 -5300 29306 -5240
rect 29366 -5300 29372 -5240
rect 29530 -5464 29590 -5080
rect 29694 -5127 29902 -5121
rect 29694 -5161 29706 -5127
rect 29890 -5161 29902 -5127
rect 29694 -5167 29902 -5161
rect 30152 -5127 30360 -5121
rect 30152 -5161 30164 -5127
rect 30348 -5161 30360 -5127
rect 30152 -5167 30360 -5161
rect 29770 -5240 29830 -5167
rect 30224 -5240 30284 -5167
rect 29764 -5300 29770 -5240
rect 29830 -5300 29836 -5240
rect 30218 -5300 30224 -5240
rect 30284 -5300 30290 -5240
rect 30454 -5348 30514 -5068
rect 30916 -5068 30926 -5046
rect 30960 -5046 30966 -3492
rect 31378 -3492 31424 -3480
rect 31378 -5040 31384 -3492
rect 30960 -5068 30976 -5046
rect 30610 -5127 30818 -5121
rect 30610 -5161 30622 -5127
rect 30806 -5161 30818 -5127
rect 30610 -5167 30818 -5161
rect 30682 -5238 30742 -5167
rect 30916 -5228 30976 -5068
rect 31372 -5068 31384 -5040
rect 31418 -5040 31424 -3492
rect 31826 -3492 31886 -3216
rect 32056 -3326 32062 -3266
rect 32122 -3326 32128 -3266
rect 32512 -3326 32518 -3266
rect 32578 -3326 32584 -3266
rect 32062 -3393 32122 -3326
rect 32518 -3393 32578 -3326
rect 31984 -3399 32192 -3393
rect 31984 -3433 31996 -3399
rect 32180 -3433 32192 -3399
rect 31984 -3439 32192 -3433
rect 32442 -3399 32650 -3393
rect 32442 -3433 32454 -3399
rect 32638 -3433 32650 -3399
rect 32442 -3439 32650 -3433
rect 31826 -3536 31842 -3492
rect 31418 -5068 31432 -5040
rect 31068 -5127 31276 -5121
rect 31068 -5161 31080 -5127
rect 31264 -5161 31276 -5127
rect 31068 -5167 31276 -5161
rect 30676 -5240 30748 -5238
rect 30676 -5300 30682 -5240
rect 30742 -5300 30748 -5240
rect 31142 -5232 31202 -5167
rect 30916 -5294 30976 -5288
rect 31130 -5238 31214 -5232
rect 31130 -5300 31142 -5238
rect 31202 -5300 31214 -5238
rect 31130 -5304 31214 -5300
rect 31372 -5348 31432 -5068
rect 31836 -5068 31842 -3536
rect 31876 -3536 31886 -3492
rect 32294 -3492 32340 -3480
rect 31876 -5068 31882 -3536
rect 32294 -5036 32300 -3492
rect 31836 -5080 31882 -5068
rect 32286 -5068 32300 -5036
rect 32334 -5036 32340 -3492
rect 32742 -3492 32802 -3092
rect 32968 -3326 32974 -3266
rect 33034 -3326 33040 -3266
rect 33424 -3326 33430 -3266
rect 33490 -3326 33496 -3266
rect 32974 -3393 33034 -3326
rect 33430 -3393 33490 -3326
rect 32900 -3399 33108 -3393
rect 32900 -3433 32912 -3399
rect 33096 -3433 33108 -3399
rect 32900 -3439 33108 -3433
rect 33358 -3399 33566 -3393
rect 33358 -3433 33370 -3399
rect 33554 -3433 33566 -3399
rect 33358 -3439 33566 -3433
rect 32742 -3550 32758 -3492
rect 32334 -5068 32346 -5036
rect 31526 -5127 31734 -5121
rect 31526 -5161 31538 -5127
rect 31722 -5161 31734 -5127
rect 31526 -5167 31734 -5161
rect 31984 -5127 32192 -5121
rect 31984 -5161 31996 -5127
rect 32180 -5161 32192 -5127
rect 31984 -5167 32192 -5161
rect 31598 -5240 31658 -5167
rect 32058 -5240 32118 -5167
rect 31592 -5300 31598 -5240
rect 31658 -5300 31664 -5240
rect 32052 -5300 32058 -5240
rect 32118 -5300 32124 -5240
rect 30454 -5408 31432 -5348
rect 32286 -5464 32346 -5068
rect 32752 -5068 32758 -3550
rect 32792 -3550 32802 -3492
rect 33210 -3492 33256 -3480
rect 32792 -5068 32798 -3550
rect 33210 -5000 33216 -3492
rect 32752 -5080 32798 -5068
rect 33206 -5068 33216 -5000
rect 33250 -5000 33256 -3492
rect 33662 -3492 33722 -2958
rect 33882 -3326 33888 -3266
rect 33948 -3326 33954 -3266
rect 34342 -3326 34348 -3266
rect 34408 -3326 34414 -3266
rect 33888 -3393 33948 -3326
rect 34348 -3393 34408 -3326
rect 33816 -3399 34024 -3393
rect 33816 -3433 33828 -3399
rect 34012 -3433 34024 -3399
rect 33816 -3439 34024 -3433
rect 34274 -3399 34482 -3393
rect 34274 -3433 34286 -3399
rect 34470 -3433 34482 -3399
rect 34274 -3439 34482 -3433
rect 33662 -3548 33674 -3492
rect 33250 -5068 33266 -5000
rect 32442 -5127 32650 -5121
rect 32442 -5161 32454 -5127
rect 32638 -5161 32650 -5127
rect 32442 -5167 32650 -5161
rect 32900 -5127 33108 -5121
rect 32900 -5161 32912 -5127
rect 33096 -5161 33108 -5127
rect 32900 -5167 33108 -5161
rect 32514 -5240 32574 -5167
rect 32970 -5240 33030 -5167
rect 32508 -5300 32514 -5240
rect 32574 -5300 32580 -5240
rect 32964 -5300 32970 -5240
rect 33030 -5300 33036 -5240
rect 29530 -5524 32346 -5464
rect 33206 -5590 33266 -5068
rect 33668 -5068 33674 -3548
rect 33708 -3548 33722 -3492
rect 34126 -3492 34172 -3480
rect 33708 -5068 33714 -3548
rect 34126 -5008 34132 -3492
rect 33668 -5080 33714 -5068
rect 34120 -5068 34132 -5008
rect 34166 -5008 34172 -3492
rect 34578 -3492 34638 -2704
rect 34808 -3393 34868 -2704
rect 34732 -3399 34940 -3393
rect 34732 -3433 34744 -3399
rect 34928 -3433 34940 -3399
rect 34732 -3439 34940 -3433
rect 34578 -3568 34590 -3492
rect 34584 -5006 34590 -3568
rect 34166 -5068 34180 -5008
rect 33358 -5127 33566 -5121
rect 33358 -5161 33370 -5127
rect 33554 -5161 33566 -5127
rect 33358 -5167 33566 -5161
rect 33816 -5127 34024 -5121
rect 33816 -5161 33828 -5127
rect 34012 -5161 34024 -5127
rect 33816 -5167 34024 -5161
rect 33426 -5240 33486 -5167
rect 33884 -5240 33944 -5167
rect 33420 -5300 33426 -5240
rect 33486 -5300 33492 -5240
rect 33878 -5300 33884 -5240
rect 33944 -5300 33950 -5240
rect 28622 -5650 33266 -5590
rect 34120 -5720 34180 -5068
rect 34574 -5068 34590 -5006
rect 34624 -3568 34638 -3492
rect 35036 -3492 35096 -2704
rect 35036 -3562 35048 -3492
rect 34624 -5006 34630 -3568
rect 34624 -5068 34634 -5006
rect 35042 -5024 35048 -3562
rect 34274 -5127 34482 -5121
rect 34274 -5161 34286 -5127
rect 34470 -5161 34482 -5127
rect 34274 -5167 34482 -5161
rect 34344 -5240 34404 -5167
rect 34338 -5300 34344 -5240
rect 34404 -5300 34410 -5240
rect 34574 -5242 34634 -5068
rect 35032 -5068 35048 -5024
rect 35082 -3562 35096 -3492
rect 35082 -5024 35088 -3562
rect 35082 -5068 35092 -5024
rect 34732 -5127 34940 -5121
rect 34732 -5161 34744 -5127
rect 34928 -5161 34940 -5127
rect 34732 -5167 34940 -5161
rect 34806 -5242 34866 -5167
rect 35032 -5242 35092 -5068
rect 36156 -5242 36162 -2418
rect 34574 -5302 36162 -5242
rect 25918 -7590 25924 -5732
rect 26232 -6157 26292 -5732
rect 26460 -6058 26520 -5732
rect 27704 -5780 34180 -5720
rect 35032 -5736 35092 -5302
rect 36156 -5736 36162 -5302
rect 35032 -5796 36162 -5736
rect 26684 -5886 26690 -5826
rect 26750 -5886 26756 -5826
rect 26387 -6064 26595 -6058
rect 26387 -6098 26399 -6064
rect 26583 -6098 26595 -6064
rect 26387 -6104 26595 -6098
rect 26232 -6204 26245 -6157
rect 26239 -7312 26245 -6204
rect 25812 -7766 25924 -7590
rect 26232 -7333 26245 -7312
rect 26279 -6204 26292 -6157
rect 26690 -6157 26750 -5886
rect 26922 -5988 30186 -5928
rect 26922 -6058 26982 -5988
rect 27384 -6058 27444 -5988
rect 27838 -6058 27898 -5988
rect 28300 -6058 28360 -5988
rect 28754 -6058 28814 -5988
rect 29204 -6058 29264 -5988
rect 29670 -6058 29730 -5988
rect 30126 -6058 30186 -5988
rect 30582 -6006 31750 -5946
rect 30582 -6058 30642 -6006
rect 26845 -6064 27053 -6058
rect 26845 -6098 26857 -6064
rect 27041 -6098 27053 -6064
rect 26845 -6104 27053 -6098
rect 27303 -6064 27511 -6058
rect 27303 -6098 27315 -6064
rect 27499 -6098 27511 -6064
rect 27303 -6104 27511 -6098
rect 27761 -6064 27969 -6058
rect 27761 -6098 27773 -6064
rect 27957 -6098 27969 -6064
rect 27761 -6104 27969 -6098
rect 28219 -6064 28427 -6058
rect 28219 -6098 28231 -6064
rect 28415 -6098 28427 -6064
rect 28219 -6104 28427 -6098
rect 28677 -6064 28885 -6058
rect 28677 -6098 28689 -6064
rect 28873 -6098 28885 -6064
rect 28677 -6104 28885 -6098
rect 29135 -6064 29343 -6058
rect 29135 -6098 29147 -6064
rect 29331 -6098 29343 -6064
rect 29135 -6104 29343 -6098
rect 29593 -6064 29801 -6058
rect 29593 -6098 29605 -6064
rect 29789 -6098 29801 -6064
rect 29593 -6104 29801 -6098
rect 30051 -6064 30259 -6058
rect 30051 -6098 30063 -6064
rect 30247 -6098 30259 -6064
rect 30051 -6104 30259 -6098
rect 30509 -6064 30717 -6058
rect 30509 -6098 30521 -6064
rect 30705 -6098 30717 -6064
rect 30509 -6104 30717 -6098
rect 26279 -7312 26285 -6204
rect 26690 -6224 26703 -6157
rect 26279 -7333 26292 -7312
rect 26232 -7766 26292 -7333
rect 26697 -7333 26703 -6224
rect 26737 -6224 26750 -6157
rect 27155 -6157 27201 -6145
rect 26737 -7333 26743 -6224
rect 26697 -7345 26743 -7333
rect 27155 -7333 27161 -6157
rect 27195 -7333 27201 -6157
rect 27155 -7345 27201 -7333
rect 27613 -6157 27659 -6145
rect 27613 -7333 27619 -6157
rect 27653 -7333 27659 -6157
rect 27613 -7345 27659 -7333
rect 28071 -6157 28117 -6145
rect 28071 -7333 28077 -6157
rect 28111 -7333 28117 -6157
rect 28071 -7345 28117 -7333
rect 28529 -6157 28575 -6145
rect 28529 -7333 28535 -6157
rect 28569 -7333 28575 -6157
rect 28529 -7345 28575 -7333
rect 28987 -6157 29033 -6145
rect 28987 -7333 28993 -6157
rect 29027 -7333 29033 -6157
rect 28987 -7345 29033 -7333
rect 29445 -6157 29491 -6145
rect 29445 -7333 29451 -6157
rect 29485 -7333 29491 -6157
rect 29445 -7345 29491 -7333
rect 29903 -6157 29949 -6145
rect 29903 -7333 29909 -6157
rect 29943 -7333 29949 -6157
rect 30361 -6157 30407 -6145
rect 30361 -7266 30367 -6157
rect 29903 -7345 29949 -7333
rect 30352 -7333 30367 -7266
rect 30401 -7266 30407 -6157
rect 30812 -6157 30872 -6006
rect 30812 -6172 30825 -6157
rect 30401 -7333 30412 -7266
rect 30819 -7298 30825 -6172
rect 26387 -7392 26595 -7386
rect 26387 -7426 26399 -7392
rect 26583 -7426 26595 -7392
rect 26387 -7432 26595 -7426
rect 26845 -7392 27053 -7386
rect 26845 -7426 26857 -7392
rect 27041 -7426 27053 -7392
rect 26845 -7432 27053 -7426
rect 27303 -7392 27511 -7386
rect 27303 -7426 27315 -7392
rect 27499 -7426 27511 -7392
rect 27303 -7432 27511 -7426
rect 27761 -7392 27969 -7386
rect 27761 -7426 27773 -7392
rect 27957 -7426 27969 -7392
rect 27761 -7432 27969 -7426
rect 28219 -7392 28427 -7386
rect 28219 -7426 28231 -7392
rect 28415 -7426 28427 -7392
rect 28219 -7432 28427 -7426
rect 28677 -7392 28885 -7386
rect 28677 -7426 28689 -7392
rect 28873 -7426 28885 -7392
rect 28677 -7432 28885 -7426
rect 29135 -7392 29343 -7386
rect 29135 -7426 29147 -7392
rect 29331 -7426 29343 -7392
rect 29135 -7432 29343 -7426
rect 29593 -7392 29801 -7386
rect 29593 -7426 29605 -7392
rect 29789 -7426 29801 -7392
rect 29593 -7432 29801 -7426
rect 30051 -7392 30259 -7386
rect 30051 -7426 30063 -7392
rect 30247 -7426 30259 -7392
rect 30051 -7432 30259 -7426
rect 26460 -7766 26520 -7432
rect 26914 -7500 26974 -7432
rect 27376 -7500 27436 -7432
rect 27830 -7500 27890 -7432
rect 28292 -7500 28352 -7432
rect 28746 -7500 28806 -7432
rect 29196 -7500 29256 -7432
rect 29662 -7500 29722 -7432
rect 30118 -7500 30178 -7432
rect 26914 -7504 27830 -7500
rect 26974 -7560 27376 -7504
rect 26914 -7570 26974 -7564
rect 27436 -7560 27830 -7504
rect 27890 -7560 28292 -7500
rect 28352 -7506 29196 -7500
rect 28352 -7560 28746 -7506
rect 27376 -7570 27436 -7564
rect 27830 -7566 27890 -7560
rect 28292 -7566 28352 -7560
rect 28806 -7560 29196 -7506
rect 29256 -7560 29662 -7500
rect 29722 -7504 30178 -7500
rect 29722 -7560 30118 -7504
rect 29196 -7566 29256 -7560
rect 29662 -7566 29722 -7560
rect 28746 -7572 28806 -7566
rect 30118 -7570 30178 -7564
rect 30352 -7626 30412 -7333
rect 30810 -7333 30825 -7298
rect 30859 -6172 30872 -6157
rect 31232 -6157 31292 -6006
rect 31464 -6058 31524 -6006
rect 31387 -6064 31595 -6058
rect 31387 -6098 31399 -6064
rect 31583 -6098 31595 -6064
rect 31387 -6104 31595 -6098
rect 30859 -7298 30865 -6172
rect 31232 -6178 31245 -6157
rect 31239 -7298 31245 -6178
rect 30859 -7333 30870 -7298
rect 30509 -7392 30717 -7386
rect 30509 -7426 30521 -7392
rect 30705 -7426 30717 -7392
rect 30509 -7432 30717 -7426
rect 30346 -7686 30352 -7626
rect 30412 -7686 30418 -7626
rect 30582 -7766 30642 -7432
rect 30810 -7766 30870 -7333
rect 31230 -7333 31245 -7298
rect 31279 -6178 31292 -6157
rect 31690 -6157 31750 -6006
rect 31916 -5988 35180 -5928
rect 31916 -6058 31976 -5988
rect 32378 -6058 32438 -5988
rect 32832 -6058 32892 -5988
rect 33294 -6058 33354 -5988
rect 33748 -6058 33808 -5988
rect 34198 -6058 34258 -5988
rect 34664 -6058 34724 -5988
rect 35120 -6058 35180 -5988
rect 35582 -6058 35642 -5796
rect 31845 -6064 32053 -6058
rect 31845 -6098 31857 -6064
rect 32041 -6098 32053 -6064
rect 31845 -6104 32053 -6098
rect 32303 -6064 32511 -6058
rect 32303 -6098 32315 -6064
rect 32499 -6098 32511 -6064
rect 32303 -6104 32511 -6098
rect 32761 -6064 32969 -6058
rect 32761 -6098 32773 -6064
rect 32957 -6098 32969 -6064
rect 32761 -6104 32969 -6098
rect 33219 -6064 33427 -6058
rect 33219 -6098 33231 -6064
rect 33415 -6098 33427 -6064
rect 33219 -6104 33427 -6098
rect 33677 -6064 33885 -6058
rect 33677 -6098 33689 -6064
rect 33873 -6098 33885 -6064
rect 33677 -6104 33885 -6098
rect 34135 -6064 34343 -6058
rect 34135 -6098 34147 -6064
rect 34331 -6098 34343 -6064
rect 34135 -6104 34343 -6098
rect 34593 -6064 34801 -6058
rect 34593 -6098 34605 -6064
rect 34789 -6098 34801 -6064
rect 34593 -6104 34801 -6098
rect 35051 -6064 35259 -6058
rect 35051 -6098 35063 -6064
rect 35247 -6098 35259 -6064
rect 35051 -6104 35259 -6098
rect 35509 -6064 35717 -6058
rect 35509 -6098 35521 -6064
rect 35705 -6098 35717 -6064
rect 35509 -6104 35717 -6098
rect 31279 -7298 31285 -6178
rect 31690 -6200 31703 -6157
rect 31697 -7292 31703 -6200
rect 31279 -7333 31290 -7298
rect 31230 -7766 31290 -7333
rect 31688 -7333 31703 -7292
rect 31737 -6200 31750 -6157
rect 32155 -6157 32201 -6145
rect 31737 -7292 31743 -6200
rect 31737 -7333 31748 -7292
rect 31387 -7392 31595 -7386
rect 31387 -7426 31399 -7392
rect 31583 -7426 31595 -7392
rect 31387 -7432 31595 -7426
rect 31458 -7766 31518 -7432
rect 31688 -7766 31748 -7333
rect 32155 -7333 32161 -6157
rect 32195 -7333 32201 -6157
rect 32155 -7345 32201 -7333
rect 32613 -6157 32659 -6145
rect 32613 -7333 32619 -6157
rect 32653 -7333 32659 -6157
rect 32613 -7345 32659 -7333
rect 33071 -6157 33117 -6145
rect 33071 -7333 33077 -6157
rect 33111 -7333 33117 -6157
rect 33071 -7345 33117 -7333
rect 33529 -6157 33575 -6145
rect 33529 -7333 33535 -6157
rect 33569 -7333 33575 -6157
rect 33529 -7345 33575 -7333
rect 33987 -6157 34033 -6145
rect 33987 -7333 33993 -6157
rect 34027 -7333 34033 -6157
rect 33987 -7345 34033 -7333
rect 34445 -6157 34491 -6145
rect 34445 -7333 34451 -6157
rect 34485 -7333 34491 -6157
rect 34445 -7345 34491 -7333
rect 34903 -6157 34949 -6145
rect 34903 -7333 34909 -6157
rect 34943 -7333 34949 -6157
rect 35361 -6157 35407 -6145
rect 35361 -7326 35367 -6157
rect 34903 -7345 34949 -7333
rect 35352 -7333 35367 -7326
rect 35401 -7326 35407 -6157
rect 35808 -6157 35868 -5796
rect 35808 -6210 35825 -6157
rect 35819 -7300 35825 -6210
rect 35401 -7333 35412 -7326
rect 31845 -7392 32053 -7386
rect 31845 -7426 31857 -7392
rect 32041 -7426 32053 -7392
rect 31845 -7432 32053 -7426
rect 32303 -7392 32511 -7386
rect 32303 -7426 32315 -7392
rect 32499 -7426 32511 -7392
rect 32303 -7432 32511 -7426
rect 32761 -7392 32969 -7386
rect 32761 -7426 32773 -7392
rect 32957 -7426 32969 -7392
rect 32761 -7432 32969 -7426
rect 33219 -7392 33427 -7386
rect 33219 -7426 33231 -7392
rect 33415 -7426 33427 -7392
rect 33219 -7432 33427 -7426
rect 33677 -7392 33885 -7386
rect 33677 -7426 33689 -7392
rect 33873 -7426 33885 -7392
rect 33677 -7432 33885 -7426
rect 34135 -7392 34343 -7386
rect 34135 -7426 34147 -7392
rect 34331 -7426 34343 -7392
rect 34135 -7432 34343 -7426
rect 34593 -7392 34801 -7386
rect 34593 -7426 34605 -7392
rect 34789 -7426 34801 -7392
rect 34593 -7432 34801 -7426
rect 35051 -7392 35259 -7386
rect 35051 -7426 35063 -7392
rect 35247 -7426 35259 -7392
rect 35051 -7432 35259 -7426
rect 31916 -7500 31976 -7432
rect 32378 -7496 32438 -7432
rect 31916 -7504 32378 -7500
rect 31976 -7556 32378 -7504
rect 32832 -7500 32892 -7432
rect 33294 -7500 33354 -7432
rect 33748 -7500 33808 -7432
rect 34198 -7496 34258 -7432
rect 32438 -7502 34198 -7500
rect 32438 -7556 32832 -7502
rect 31976 -7560 32832 -7556
rect 32378 -7562 32438 -7560
rect 32892 -7560 33294 -7502
rect 31916 -7570 31976 -7564
rect 32832 -7568 32892 -7562
rect 33354 -7560 33748 -7502
rect 33294 -7568 33354 -7562
rect 33808 -7556 34198 -7502
rect 34664 -7500 34724 -7432
rect 35120 -7500 35180 -7432
rect 34258 -7502 35180 -7500
rect 34258 -7556 34664 -7502
rect 33808 -7560 34664 -7556
rect 34198 -7562 34258 -7560
rect 34724 -7560 35120 -7502
rect 33748 -7568 33808 -7562
rect 34664 -7568 34724 -7562
rect 35120 -7568 35180 -7562
rect 35352 -7632 35412 -7333
rect 35810 -7333 35825 -7300
rect 35859 -6210 35868 -6157
rect 35859 -7300 35865 -6210
rect 35859 -7333 35870 -7300
rect 35509 -7392 35717 -7386
rect 35509 -7426 35521 -7392
rect 35705 -7426 35717 -7392
rect 35509 -7432 35717 -7426
rect 35352 -7698 35412 -7692
rect 35582 -7766 35642 -7432
rect 35810 -7766 35870 -7333
rect 36156 -7590 36162 -5796
rect 36262 -7590 36268 -2418
rect 36156 -7766 36268 -7590
rect 25812 -7772 36268 -7766
rect 25812 -7872 25918 -7772
rect 36162 -7872 36268 -7772
rect 25812 -7878 36268 -7872
rect 25812 -8108 36268 -8102
rect 25812 -8208 25918 -8108
rect 36162 -8208 36268 -8108
rect 25812 -8214 36268 -8208
rect 25812 -8338 25924 -8214
rect 25540 -9710 25546 -9650
rect 25606 -9710 25612 -9650
rect 10812 -20028 21268 -20022
rect 10812 -20128 10918 -20028
rect 21162 -20128 21268 -20028
rect 10812 -20134 21268 -20128
rect 10812 -20418 10924 -20134
rect 10812 -25590 10818 -20418
rect 10918 -23240 10924 -20418
rect 11524 -20434 11534 -20134
rect 20546 -20434 20556 -20134
rect 21156 -20418 21268 -20134
rect 11762 -20608 20118 -20594
rect 11762 -20694 11776 -20608
rect 11872 -20694 12376 -20608
rect 12472 -20694 12976 -20608
rect 13072 -20694 13576 -20608
rect 13672 -20694 14176 -20608
rect 14272 -20694 14776 -20608
rect 14872 -20694 15376 -20608
rect 15472 -20694 15976 -20608
rect 16072 -20694 16576 -20608
rect 16672 -20694 17176 -20608
rect 17272 -20694 17776 -20608
rect 17872 -20694 18376 -20608
rect 18472 -20694 18976 -20608
rect 19072 -20694 19576 -20608
rect 19672 -20694 19996 -20608
rect 20092 -20694 20118 -20608
rect 11762 -20704 20118 -20694
rect 11790 -21492 11850 -20704
rect 12022 -21393 12082 -20704
rect 11946 -21399 12154 -21393
rect 11946 -21433 11958 -21399
rect 12142 -21433 12154 -21399
rect 11946 -21439 12154 -21433
rect 11790 -21524 11804 -21492
rect 11798 -23008 11804 -21524
rect 11792 -23068 11804 -23008
rect 11838 -21524 11850 -21492
rect 12248 -21492 12308 -20704
rect 13164 -20958 18722 -20898
rect 12474 -21326 12480 -21266
rect 12540 -21326 12546 -21266
rect 12930 -21326 12936 -21266
rect 12996 -21326 13002 -21266
rect 12480 -21393 12540 -21326
rect 12936 -21393 12996 -21326
rect 12404 -21399 12612 -21393
rect 12404 -21433 12416 -21399
rect 12600 -21433 12612 -21399
rect 12404 -21439 12612 -21433
rect 12862 -21399 13070 -21393
rect 12862 -21433 12874 -21399
rect 13058 -21433 13070 -21399
rect 12862 -21439 13070 -21433
rect 11838 -23008 11844 -21524
rect 12248 -21556 12262 -21492
rect 11838 -23068 11852 -23008
rect 12256 -23024 12262 -21556
rect 11792 -23240 11852 -23068
rect 12246 -23068 12262 -23024
rect 12296 -21556 12308 -21492
rect 12714 -21492 12760 -21480
rect 12296 -23024 12302 -21556
rect 12714 -22984 12720 -21492
rect 12296 -23068 12306 -23024
rect 11946 -23127 12154 -23121
rect 11946 -23161 11958 -23127
rect 12142 -23161 12154 -23127
rect 11946 -23167 12154 -23161
rect 12020 -23240 12080 -23167
rect 12246 -23240 12306 -23068
rect 12704 -23068 12720 -22984
rect 12754 -22984 12760 -21492
rect 13164 -21492 13224 -20958
rect 14080 -21092 17802 -21032
rect 13390 -21326 13396 -21266
rect 13456 -21326 13462 -21266
rect 13846 -21326 13852 -21266
rect 13912 -21326 13918 -21266
rect 13396 -21393 13456 -21326
rect 13852 -21393 13912 -21326
rect 13320 -21399 13528 -21393
rect 13320 -21433 13332 -21399
rect 13516 -21433 13528 -21399
rect 13320 -21439 13528 -21433
rect 13778 -21399 13986 -21393
rect 13778 -21433 13790 -21399
rect 13974 -21433 13986 -21399
rect 13778 -21439 13986 -21433
rect 13164 -21550 13178 -21492
rect 12754 -23068 12764 -22984
rect 12404 -23127 12612 -23121
rect 12404 -23161 12416 -23127
rect 12600 -23161 12612 -23127
rect 12404 -23167 12612 -23161
rect 12476 -23240 12536 -23167
rect 10918 -23300 12306 -23240
rect 12470 -23300 12476 -23240
rect 12536 -23300 12542 -23240
rect 10918 -23672 10924 -23300
rect 11792 -23672 11852 -23300
rect 10918 -23732 11852 -23672
rect 12704 -23720 12764 -23068
rect 13172 -23068 13178 -21550
rect 13212 -21550 13224 -21492
rect 13630 -21492 13676 -21480
rect 13212 -23068 13218 -21550
rect 13630 -22990 13636 -21492
rect 13172 -23080 13218 -23068
rect 13622 -23068 13636 -22990
rect 13670 -22990 13676 -21492
rect 14080 -21492 14140 -21092
rect 14996 -21216 16886 -21156
rect 14304 -21326 14310 -21266
rect 14370 -21326 14376 -21266
rect 14768 -21326 14774 -21266
rect 14834 -21326 14840 -21266
rect 14310 -21393 14370 -21326
rect 14774 -21393 14834 -21326
rect 14236 -21399 14444 -21393
rect 14236 -21433 14248 -21399
rect 14432 -21433 14444 -21399
rect 14236 -21439 14444 -21433
rect 14694 -21399 14902 -21393
rect 14694 -21433 14706 -21399
rect 14890 -21433 14902 -21399
rect 14694 -21439 14902 -21433
rect 14080 -21552 14094 -21492
rect 13670 -23068 13682 -22990
rect 12862 -23127 13070 -23121
rect 12862 -23161 12874 -23127
rect 13058 -23161 13070 -23127
rect 12862 -23167 13070 -23161
rect 13320 -23127 13528 -23121
rect 13320 -23161 13332 -23127
rect 13516 -23161 13528 -23127
rect 13320 -23167 13528 -23161
rect 12932 -23240 12992 -23167
rect 13392 -23240 13452 -23167
rect 12926 -23300 12932 -23240
rect 12992 -23300 12998 -23240
rect 13386 -23300 13392 -23240
rect 13452 -23300 13458 -23240
rect 13622 -23590 13682 -23068
rect 14088 -23068 14094 -21552
rect 14128 -21552 14140 -21492
rect 14546 -21492 14592 -21480
rect 14128 -23068 14134 -21552
rect 14546 -22996 14552 -21492
rect 14088 -23080 14134 -23068
rect 14530 -23068 14552 -22996
rect 14586 -23068 14592 -21492
rect 14996 -21492 15056 -21216
rect 15218 -21326 15224 -21266
rect 15284 -21326 15290 -21266
rect 15674 -21326 15680 -21266
rect 15740 -21326 15746 -21266
rect 16142 -21326 16148 -21266
rect 16208 -21326 16214 -21266
rect 16600 -21326 16606 -21266
rect 16666 -21326 16672 -21266
rect 15224 -21393 15284 -21326
rect 15680 -21393 15740 -21326
rect 16148 -21393 16208 -21326
rect 16606 -21393 16666 -21326
rect 15152 -21399 15360 -21393
rect 15152 -21433 15164 -21399
rect 15348 -21433 15360 -21399
rect 15152 -21439 15360 -21433
rect 15610 -21399 15818 -21393
rect 15610 -21433 15622 -21399
rect 15806 -21433 15818 -21399
rect 15610 -21439 15818 -21433
rect 16068 -21399 16276 -21393
rect 16068 -21433 16080 -21399
rect 16264 -21433 16276 -21399
rect 16068 -21439 16276 -21433
rect 16526 -21399 16734 -21393
rect 16526 -21433 16538 -21399
rect 16722 -21433 16734 -21399
rect 16526 -21439 16734 -21433
rect 14996 -21570 15010 -21492
rect 14530 -23080 14592 -23068
rect 15004 -23068 15010 -21570
rect 15044 -21570 15056 -21492
rect 15462 -21492 15508 -21480
rect 15044 -23068 15050 -21570
rect 15462 -22988 15468 -21492
rect 15004 -23080 15050 -23068
rect 15454 -23068 15468 -22988
rect 15502 -22988 15508 -21492
rect 15920 -21492 15966 -21480
rect 15502 -23068 15514 -22988
rect 15920 -23046 15926 -21492
rect 13778 -23127 13986 -23121
rect 13778 -23161 13790 -23127
rect 13974 -23161 13986 -23127
rect 13778 -23167 13986 -23161
rect 14236 -23127 14444 -23121
rect 14236 -23161 14248 -23127
rect 14432 -23161 14444 -23127
rect 14236 -23167 14444 -23161
rect 13848 -23240 13908 -23167
rect 14306 -23240 14366 -23167
rect 13842 -23300 13848 -23240
rect 13908 -23300 13914 -23240
rect 14300 -23300 14306 -23240
rect 14366 -23300 14372 -23240
rect 14530 -23464 14590 -23080
rect 14694 -23127 14902 -23121
rect 14694 -23161 14706 -23127
rect 14890 -23161 14902 -23127
rect 14694 -23167 14902 -23161
rect 15152 -23127 15360 -23121
rect 15152 -23161 15164 -23127
rect 15348 -23161 15360 -23127
rect 15152 -23167 15360 -23161
rect 14770 -23240 14830 -23167
rect 15224 -23240 15284 -23167
rect 14764 -23300 14770 -23240
rect 14830 -23300 14836 -23240
rect 15218 -23300 15224 -23240
rect 15284 -23300 15290 -23240
rect 15454 -23348 15514 -23068
rect 15916 -23068 15926 -23046
rect 15960 -23046 15966 -21492
rect 16378 -21492 16424 -21480
rect 16378 -23040 16384 -21492
rect 15960 -23068 15976 -23046
rect 15610 -23127 15818 -23121
rect 15610 -23161 15622 -23127
rect 15806 -23161 15818 -23127
rect 15610 -23167 15818 -23161
rect 15682 -23238 15742 -23167
rect 15916 -23228 15976 -23068
rect 16372 -23068 16384 -23040
rect 16418 -23040 16424 -21492
rect 16826 -21492 16886 -21216
rect 17056 -21326 17062 -21266
rect 17122 -21326 17128 -21266
rect 17512 -21326 17518 -21266
rect 17578 -21326 17584 -21266
rect 17062 -21393 17122 -21326
rect 17518 -21393 17578 -21326
rect 16984 -21399 17192 -21393
rect 16984 -21433 16996 -21399
rect 17180 -21433 17192 -21399
rect 16984 -21439 17192 -21433
rect 17442 -21399 17650 -21393
rect 17442 -21433 17454 -21399
rect 17638 -21433 17650 -21399
rect 17442 -21439 17650 -21433
rect 16826 -21536 16842 -21492
rect 16418 -23068 16432 -23040
rect 16068 -23127 16276 -23121
rect 16068 -23161 16080 -23127
rect 16264 -23161 16276 -23127
rect 16068 -23167 16276 -23161
rect 15676 -23240 15748 -23238
rect 15676 -23300 15682 -23240
rect 15742 -23300 15748 -23240
rect 16142 -23232 16202 -23167
rect 15916 -23294 15976 -23288
rect 16130 -23238 16214 -23232
rect 16130 -23300 16142 -23238
rect 16202 -23300 16214 -23238
rect 16130 -23304 16214 -23300
rect 16372 -23348 16432 -23068
rect 16836 -23068 16842 -21536
rect 16876 -21536 16886 -21492
rect 17294 -21492 17340 -21480
rect 16876 -23068 16882 -21536
rect 17294 -23036 17300 -21492
rect 16836 -23080 16882 -23068
rect 17286 -23068 17300 -23036
rect 17334 -23036 17340 -21492
rect 17742 -21492 17802 -21092
rect 17968 -21326 17974 -21266
rect 18034 -21326 18040 -21266
rect 18424 -21326 18430 -21266
rect 18490 -21326 18496 -21266
rect 17974 -21393 18034 -21326
rect 18430 -21393 18490 -21326
rect 17900 -21399 18108 -21393
rect 17900 -21433 17912 -21399
rect 18096 -21433 18108 -21399
rect 17900 -21439 18108 -21433
rect 18358 -21399 18566 -21393
rect 18358 -21433 18370 -21399
rect 18554 -21433 18566 -21399
rect 18358 -21439 18566 -21433
rect 17742 -21550 17758 -21492
rect 17334 -23068 17346 -23036
rect 16526 -23127 16734 -23121
rect 16526 -23161 16538 -23127
rect 16722 -23161 16734 -23127
rect 16526 -23167 16734 -23161
rect 16984 -23127 17192 -23121
rect 16984 -23161 16996 -23127
rect 17180 -23161 17192 -23127
rect 16984 -23167 17192 -23161
rect 16598 -23240 16658 -23167
rect 17058 -23240 17118 -23167
rect 16592 -23300 16598 -23240
rect 16658 -23300 16664 -23240
rect 17052 -23300 17058 -23240
rect 17118 -23300 17124 -23240
rect 15454 -23408 16432 -23348
rect 17286 -23464 17346 -23068
rect 17752 -23068 17758 -21550
rect 17792 -21550 17802 -21492
rect 18210 -21492 18256 -21480
rect 17792 -23068 17798 -21550
rect 18210 -23000 18216 -21492
rect 17752 -23080 17798 -23068
rect 18206 -23068 18216 -23000
rect 18250 -23000 18256 -21492
rect 18662 -21492 18722 -20958
rect 18882 -21326 18888 -21266
rect 18948 -21326 18954 -21266
rect 19342 -21326 19348 -21266
rect 19408 -21326 19414 -21266
rect 18888 -21393 18948 -21326
rect 19348 -21393 19408 -21326
rect 18816 -21399 19024 -21393
rect 18816 -21433 18828 -21399
rect 19012 -21433 19024 -21399
rect 18816 -21439 19024 -21433
rect 19274 -21399 19482 -21393
rect 19274 -21433 19286 -21399
rect 19470 -21433 19482 -21399
rect 19274 -21439 19482 -21433
rect 18662 -21548 18674 -21492
rect 18250 -23068 18266 -23000
rect 17442 -23127 17650 -23121
rect 17442 -23161 17454 -23127
rect 17638 -23161 17650 -23127
rect 17442 -23167 17650 -23161
rect 17900 -23127 18108 -23121
rect 17900 -23161 17912 -23127
rect 18096 -23161 18108 -23127
rect 17900 -23167 18108 -23161
rect 17514 -23240 17574 -23167
rect 17970 -23240 18030 -23167
rect 17508 -23300 17514 -23240
rect 17574 -23300 17580 -23240
rect 17964 -23300 17970 -23240
rect 18030 -23300 18036 -23240
rect 14530 -23524 17346 -23464
rect 18206 -23590 18266 -23068
rect 18668 -23068 18674 -21548
rect 18708 -21548 18722 -21492
rect 19126 -21492 19172 -21480
rect 18708 -23068 18714 -21548
rect 19126 -23008 19132 -21492
rect 18668 -23080 18714 -23068
rect 19120 -23068 19132 -23008
rect 19166 -23008 19172 -21492
rect 19578 -21492 19638 -20704
rect 19808 -21393 19868 -20704
rect 19732 -21399 19940 -21393
rect 19732 -21433 19744 -21399
rect 19928 -21433 19940 -21399
rect 19732 -21439 19940 -21433
rect 19578 -21568 19590 -21492
rect 19584 -23006 19590 -21568
rect 19166 -23068 19180 -23008
rect 18358 -23127 18566 -23121
rect 18358 -23161 18370 -23127
rect 18554 -23161 18566 -23127
rect 18358 -23167 18566 -23161
rect 18816 -23127 19024 -23121
rect 18816 -23161 18828 -23127
rect 19012 -23161 19024 -23127
rect 18816 -23167 19024 -23161
rect 18426 -23240 18486 -23167
rect 18884 -23240 18944 -23167
rect 18420 -23300 18426 -23240
rect 18486 -23300 18492 -23240
rect 18878 -23300 18884 -23240
rect 18944 -23300 18950 -23240
rect 13622 -23650 18266 -23590
rect 19120 -23720 19180 -23068
rect 19574 -23068 19590 -23006
rect 19624 -21568 19638 -21492
rect 20036 -21492 20096 -20704
rect 20036 -21562 20048 -21492
rect 19624 -23006 19630 -21568
rect 19624 -23068 19634 -23006
rect 20042 -23024 20048 -21562
rect 19274 -23127 19482 -23121
rect 19274 -23161 19286 -23127
rect 19470 -23161 19482 -23127
rect 19274 -23167 19482 -23161
rect 19344 -23240 19404 -23167
rect 19338 -23300 19344 -23240
rect 19404 -23300 19410 -23240
rect 19574 -23242 19634 -23068
rect 20032 -23068 20048 -23024
rect 20082 -21562 20096 -21492
rect 20082 -23024 20088 -21562
rect 20082 -23068 20092 -23024
rect 19732 -23127 19940 -23121
rect 19732 -23161 19744 -23127
rect 19928 -23161 19940 -23127
rect 19732 -23167 19940 -23161
rect 19806 -23242 19866 -23167
rect 20032 -23242 20092 -23068
rect 21156 -23242 21162 -20418
rect 19574 -23302 21162 -23242
rect 10918 -25590 10924 -23732
rect 11232 -24157 11292 -23732
rect 11460 -24058 11520 -23732
rect 12704 -23780 19180 -23720
rect 20032 -23736 20092 -23302
rect 21156 -23736 21162 -23302
rect 20032 -23796 21162 -23736
rect 11684 -23886 11690 -23826
rect 11750 -23886 11756 -23826
rect 11387 -24064 11595 -24058
rect 11387 -24098 11399 -24064
rect 11583 -24098 11595 -24064
rect 11387 -24104 11595 -24098
rect 11232 -24204 11245 -24157
rect 11239 -25312 11245 -24204
rect 10812 -25766 10924 -25590
rect 11232 -25333 11245 -25312
rect 11279 -24204 11292 -24157
rect 11690 -24157 11750 -23886
rect 11922 -23988 15186 -23928
rect 11922 -24058 11982 -23988
rect 12384 -24058 12444 -23988
rect 12838 -24058 12898 -23988
rect 13300 -24058 13360 -23988
rect 13754 -24058 13814 -23988
rect 14204 -24058 14264 -23988
rect 14670 -24058 14730 -23988
rect 15126 -24058 15186 -23988
rect 15582 -24006 16750 -23946
rect 15582 -24058 15642 -24006
rect 11845 -24064 12053 -24058
rect 11845 -24098 11857 -24064
rect 12041 -24098 12053 -24064
rect 11845 -24104 12053 -24098
rect 12303 -24064 12511 -24058
rect 12303 -24098 12315 -24064
rect 12499 -24098 12511 -24064
rect 12303 -24104 12511 -24098
rect 12761 -24064 12969 -24058
rect 12761 -24098 12773 -24064
rect 12957 -24098 12969 -24064
rect 12761 -24104 12969 -24098
rect 13219 -24064 13427 -24058
rect 13219 -24098 13231 -24064
rect 13415 -24098 13427 -24064
rect 13219 -24104 13427 -24098
rect 13677 -24064 13885 -24058
rect 13677 -24098 13689 -24064
rect 13873 -24098 13885 -24064
rect 13677 -24104 13885 -24098
rect 14135 -24064 14343 -24058
rect 14135 -24098 14147 -24064
rect 14331 -24098 14343 -24064
rect 14135 -24104 14343 -24098
rect 14593 -24064 14801 -24058
rect 14593 -24098 14605 -24064
rect 14789 -24098 14801 -24064
rect 14593 -24104 14801 -24098
rect 15051 -24064 15259 -24058
rect 15051 -24098 15063 -24064
rect 15247 -24098 15259 -24064
rect 15051 -24104 15259 -24098
rect 15509 -24064 15717 -24058
rect 15509 -24098 15521 -24064
rect 15705 -24098 15717 -24064
rect 15509 -24104 15717 -24098
rect 11279 -25312 11285 -24204
rect 11690 -24224 11703 -24157
rect 11279 -25333 11292 -25312
rect 11232 -25766 11292 -25333
rect 11697 -25333 11703 -24224
rect 11737 -24224 11750 -24157
rect 12155 -24157 12201 -24145
rect 11737 -25333 11743 -24224
rect 11697 -25345 11743 -25333
rect 12155 -25333 12161 -24157
rect 12195 -25333 12201 -24157
rect 12155 -25345 12201 -25333
rect 12613 -24157 12659 -24145
rect 12613 -25333 12619 -24157
rect 12653 -25333 12659 -24157
rect 12613 -25345 12659 -25333
rect 13071 -24157 13117 -24145
rect 13071 -25333 13077 -24157
rect 13111 -25333 13117 -24157
rect 13071 -25345 13117 -25333
rect 13529 -24157 13575 -24145
rect 13529 -25333 13535 -24157
rect 13569 -25333 13575 -24157
rect 13529 -25345 13575 -25333
rect 13987 -24157 14033 -24145
rect 13987 -25333 13993 -24157
rect 14027 -25333 14033 -24157
rect 13987 -25345 14033 -25333
rect 14445 -24157 14491 -24145
rect 14445 -25333 14451 -24157
rect 14485 -25333 14491 -24157
rect 14445 -25345 14491 -25333
rect 14903 -24157 14949 -24145
rect 14903 -25333 14909 -24157
rect 14943 -25333 14949 -24157
rect 15361 -24157 15407 -24145
rect 15361 -25266 15367 -24157
rect 14903 -25345 14949 -25333
rect 15352 -25333 15367 -25266
rect 15401 -25266 15407 -24157
rect 15812 -24157 15872 -24006
rect 15812 -24172 15825 -24157
rect 15401 -25333 15412 -25266
rect 15819 -25298 15825 -24172
rect 11387 -25392 11595 -25386
rect 11387 -25426 11399 -25392
rect 11583 -25426 11595 -25392
rect 11387 -25432 11595 -25426
rect 11845 -25392 12053 -25386
rect 11845 -25426 11857 -25392
rect 12041 -25426 12053 -25392
rect 11845 -25432 12053 -25426
rect 12303 -25392 12511 -25386
rect 12303 -25426 12315 -25392
rect 12499 -25426 12511 -25392
rect 12303 -25432 12511 -25426
rect 12761 -25392 12969 -25386
rect 12761 -25426 12773 -25392
rect 12957 -25426 12969 -25392
rect 12761 -25432 12969 -25426
rect 13219 -25392 13427 -25386
rect 13219 -25426 13231 -25392
rect 13415 -25426 13427 -25392
rect 13219 -25432 13427 -25426
rect 13677 -25392 13885 -25386
rect 13677 -25426 13689 -25392
rect 13873 -25426 13885 -25392
rect 13677 -25432 13885 -25426
rect 14135 -25392 14343 -25386
rect 14135 -25426 14147 -25392
rect 14331 -25426 14343 -25392
rect 14135 -25432 14343 -25426
rect 14593 -25392 14801 -25386
rect 14593 -25426 14605 -25392
rect 14789 -25426 14801 -25392
rect 14593 -25432 14801 -25426
rect 15051 -25392 15259 -25386
rect 15051 -25426 15063 -25392
rect 15247 -25426 15259 -25392
rect 15051 -25432 15259 -25426
rect 11460 -25766 11520 -25432
rect 11914 -25500 11974 -25432
rect 12376 -25500 12436 -25432
rect 12830 -25500 12890 -25432
rect 13292 -25500 13352 -25432
rect 13746 -25500 13806 -25432
rect 14196 -25500 14256 -25432
rect 14662 -25500 14722 -25432
rect 15118 -25500 15178 -25432
rect 11914 -25504 12830 -25500
rect 11974 -25560 12376 -25504
rect 11914 -25570 11974 -25564
rect 12436 -25560 12830 -25504
rect 12890 -25560 13292 -25500
rect 13352 -25506 14196 -25500
rect 13352 -25560 13746 -25506
rect 12376 -25570 12436 -25564
rect 12830 -25566 12890 -25560
rect 13292 -25566 13352 -25560
rect 13806 -25560 14196 -25506
rect 14256 -25560 14662 -25500
rect 14722 -25504 15178 -25500
rect 14722 -25560 15118 -25504
rect 14196 -25566 14256 -25560
rect 14662 -25566 14722 -25560
rect 13746 -25572 13806 -25566
rect 15118 -25570 15178 -25564
rect 15352 -25626 15412 -25333
rect 15810 -25333 15825 -25298
rect 15859 -24172 15872 -24157
rect 16232 -24157 16292 -24006
rect 16464 -24058 16524 -24006
rect 16387 -24064 16595 -24058
rect 16387 -24098 16399 -24064
rect 16583 -24098 16595 -24064
rect 16387 -24104 16595 -24098
rect 15859 -25298 15865 -24172
rect 16232 -24178 16245 -24157
rect 16239 -25298 16245 -24178
rect 15859 -25333 15870 -25298
rect 15509 -25392 15717 -25386
rect 15509 -25426 15521 -25392
rect 15705 -25426 15717 -25392
rect 15509 -25432 15717 -25426
rect 15346 -25686 15352 -25626
rect 15412 -25686 15418 -25626
rect 15582 -25766 15642 -25432
rect 15810 -25766 15870 -25333
rect 16230 -25333 16245 -25298
rect 16279 -24178 16292 -24157
rect 16690 -24157 16750 -24006
rect 16916 -23988 20180 -23928
rect 16916 -24058 16976 -23988
rect 17378 -24058 17438 -23988
rect 17832 -24058 17892 -23988
rect 18294 -24058 18354 -23988
rect 18748 -24058 18808 -23988
rect 19198 -24058 19258 -23988
rect 19664 -24058 19724 -23988
rect 20120 -24058 20180 -23988
rect 20582 -24058 20642 -23796
rect 16845 -24064 17053 -24058
rect 16845 -24098 16857 -24064
rect 17041 -24098 17053 -24064
rect 16845 -24104 17053 -24098
rect 17303 -24064 17511 -24058
rect 17303 -24098 17315 -24064
rect 17499 -24098 17511 -24064
rect 17303 -24104 17511 -24098
rect 17761 -24064 17969 -24058
rect 17761 -24098 17773 -24064
rect 17957 -24098 17969 -24064
rect 17761 -24104 17969 -24098
rect 18219 -24064 18427 -24058
rect 18219 -24098 18231 -24064
rect 18415 -24098 18427 -24064
rect 18219 -24104 18427 -24098
rect 18677 -24064 18885 -24058
rect 18677 -24098 18689 -24064
rect 18873 -24098 18885 -24064
rect 18677 -24104 18885 -24098
rect 19135 -24064 19343 -24058
rect 19135 -24098 19147 -24064
rect 19331 -24098 19343 -24064
rect 19135 -24104 19343 -24098
rect 19593 -24064 19801 -24058
rect 19593 -24098 19605 -24064
rect 19789 -24098 19801 -24064
rect 19593 -24104 19801 -24098
rect 20051 -24064 20259 -24058
rect 20051 -24098 20063 -24064
rect 20247 -24098 20259 -24064
rect 20051 -24104 20259 -24098
rect 20509 -24064 20717 -24058
rect 20509 -24098 20521 -24064
rect 20705 -24098 20717 -24064
rect 20509 -24104 20717 -24098
rect 16279 -25298 16285 -24178
rect 16690 -24200 16703 -24157
rect 16697 -25292 16703 -24200
rect 16279 -25333 16290 -25298
rect 16230 -25766 16290 -25333
rect 16688 -25333 16703 -25292
rect 16737 -24200 16750 -24157
rect 17155 -24157 17201 -24145
rect 16737 -25292 16743 -24200
rect 16737 -25333 16748 -25292
rect 16387 -25392 16595 -25386
rect 16387 -25426 16399 -25392
rect 16583 -25426 16595 -25392
rect 16387 -25432 16595 -25426
rect 16458 -25766 16518 -25432
rect 16688 -25766 16748 -25333
rect 17155 -25333 17161 -24157
rect 17195 -25333 17201 -24157
rect 17155 -25345 17201 -25333
rect 17613 -24157 17659 -24145
rect 17613 -25333 17619 -24157
rect 17653 -25333 17659 -24157
rect 17613 -25345 17659 -25333
rect 18071 -24157 18117 -24145
rect 18071 -25333 18077 -24157
rect 18111 -25333 18117 -24157
rect 18071 -25345 18117 -25333
rect 18529 -24157 18575 -24145
rect 18529 -25333 18535 -24157
rect 18569 -25333 18575 -24157
rect 18529 -25345 18575 -25333
rect 18987 -24157 19033 -24145
rect 18987 -25333 18993 -24157
rect 19027 -25333 19033 -24157
rect 18987 -25345 19033 -25333
rect 19445 -24157 19491 -24145
rect 19445 -25333 19451 -24157
rect 19485 -25333 19491 -24157
rect 19445 -25345 19491 -25333
rect 19903 -24157 19949 -24145
rect 19903 -25333 19909 -24157
rect 19943 -25333 19949 -24157
rect 20361 -24157 20407 -24145
rect 20361 -25326 20367 -24157
rect 19903 -25345 19949 -25333
rect 20352 -25333 20367 -25326
rect 20401 -25326 20407 -24157
rect 20808 -24157 20868 -23796
rect 20808 -24210 20825 -24157
rect 20819 -25300 20825 -24210
rect 20401 -25333 20412 -25326
rect 16845 -25392 17053 -25386
rect 16845 -25426 16857 -25392
rect 17041 -25426 17053 -25392
rect 16845 -25432 17053 -25426
rect 17303 -25392 17511 -25386
rect 17303 -25426 17315 -25392
rect 17499 -25426 17511 -25392
rect 17303 -25432 17511 -25426
rect 17761 -25392 17969 -25386
rect 17761 -25426 17773 -25392
rect 17957 -25426 17969 -25392
rect 17761 -25432 17969 -25426
rect 18219 -25392 18427 -25386
rect 18219 -25426 18231 -25392
rect 18415 -25426 18427 -25392
rect 18219 -25432 18427 -25426
rect 18677 -25392 18885 -25386
rect 18677 -25426 18689 -25392
rect 18873 -25426 18885 -25392
rect 18677 -25432 18885 -25426
rect 19135 -25392 19343 -25386
rect 19135 -25426 19147 -25392
rect 19331 -25426 19343 -25392
rect 19135 -25432 19343 -25426
rect 19593 -25392 19801 -25386
rect 19593 -25426 19605 -25392
rect 19789 -25426 19801 -25392
rect 19593 -25432 19801 -25426
rect 20051 -25392 20259 -25386
rect 20051 -25426 20063 -25392
rect 20247 -25426 20259 -25392
rect 20051 -25432 20259 -25426
rect 16916 -25500 16976 -25432
rect 17378 -25496 17438 -25432
rect 16916 -25504 17378 -25500
rect 16976 -25556 17378 -25504
rect 17832 -25500 17892 -25432
rect 18294 -25500 18354 -25432
rect 18748 -25500 18808 -25432
rect 19198 -25496 19258 -25432
rect 17438 -25502 19198 -25500
rect 17438 -25556 17832 -25502
rect 16976 -25560 17832 -25556
rect 17378 -25562 17438 -25560
rect 17892 -25560 18294 -25502
rect 16916 -25570 16976 -25564
rect 17832 -25568 17892 -25562
rect 18354 -25560 18748 -25502
rect 18294 -25568 18354 -25562
rect 18808 -25556 19198 -25502
rect 19664 -25500 19724 -25432
rect 20120 -25500 20180 -25432
rect 19258 -25502 20180 -25500
rect 19258 -25556 19664 -25502
rect 18808 -25560 19664 -25556
rect 19198 -25562 19258 -25560
rect 19724 -25560 20120 -25502
rect 18748 -25568 18808 -25562
rect 19664 -25568 19724 -25562
rect 20120 -25568 20180 -25562
rect 20352 -25632 20412 -25333
rect 20810 -25333 20825 -25300
rect 20859 -24210 20868 -24157
rect 20859 -25300 20865 -24210
rect 20859 -25333 20870 -25300
rect 20509 -25392 20717 -25386
rect 20509 -25426 20521 -25392
rect 20705 -25426 20717 -25392
rect 20509 -25432 20717 -25426
rect 20352 -25698 20412 -25692
rect 20582 -25766 20642 -25432
rect 20810 -25766 20870 -25333
rect 21156 -25590 21162 -23796
rect 21262 -25590 21268 -20418
rect 25406 -23240 25466 -16364
rect 25546 -11894 25606 -9710
rect 25812 -10342 25818 -8338
rect 25918 -10342 25924 -8338
rect 26232 -8650 26292 -8214
rect 26462 -8560 26522 -8214
rect 30352 -8306 30412 -8300
rect 26920 -8440 27376 -8434
rect 26908 -8500 26914 -8440
rect 26974 -8494 27376 -8440
rect 27436 -8440 28292 -8434
rect 27436 -8494 27830 -8440
rect 26974 -8500 26980 -8494
rect 26914 -8560 26980 -8500
rect 27376 -8560 27442 -8494
rect 27824 -8500 27830 -8494
rect 27890 -8494 28292 -8440
rect 28352 -8494 28746 -8434
rect 28806 -8494 29196 -8434
rect 29256 -8440 30118 -8434
rect 29256 -8494 29662 -8440
rect 27890 -8500 27896 -8494
rect 27830 -8560 27896 -8500
rect 28292 -8560 28358 -8494
rect 28746 -8560 28812 -8494
rect 29196 -8560 29262 -8494
rect 29656 -8500 29662 -8494
rect 29722 -8494 30118 -8440
rect 30178 -8494 30184 -8434
rect 29722 -8500 29728 -8494
rect 29662 -8560 29728 -8500
rect 30118 -8560 30184 -8494
rect 26386 -8566 26594 -8560
rect 26386 -8600 26398 -8566
rect 26582 -8600 26594 -8566
rect 26386 -8606 26594 -8600
rect 26844 -8566 27052 -8560
rect 26844 -8600 26856 -8566
rect 27040 -8600 27052 -8566
rect 26844 -8606 27052 -8600
rect 27302 -8566 27510 -8560
rect 27302 -8600 27314 -8566
rect 27498 -8600 27510 -8566
rect 27302 -8606 27510 -8600
rect 27760 -8566 27968 -8560
rect 27760 -8600 27772 -8566
rect 27956 -8600 27968 -8566
rect 27760 -8606 27968 -8600
rect 28218 -8566 28426 -8560
rect 28218 -8600 28230 -8566
rect 28414 -8600 28426 -8566
rect 28218 -8606 28426 -8600
rect 28676 -8566 28884 -8560
rect 28676 -8600 28688 -8566
rect 28872 -8600 28884 -8566
rect 28676 -8606 28884 -8600
rect 29134 -8566 29342 -8560
rect 29134 -8600 29146 -8566
rect 29330 -8600 29342 -8566
rect 29134 -8606 29342 -8600
rect 29592 -8566 29800 -8560
rect 29592 -8600 29604 -8566
rect 29788 -8600 29800 -8566
rect 29592 -8606 29800 -8600
rect 30050 -8566 30258 -8560
rect 30050 -8600 30062 -8566
rect 30246 -8600 30258 -8566
rect 30050 -8606 30258 -8600
rect 26232 -8690 26244 -8650
rect 26238 -8786 26244 -8690
rect 26232 -8826 26244 -8786
rect 26278 -8690 26292 -8650
rect 26696 -8650 26742 -8638
rect 26278 -8786 26284 -8690
rect 26696 -8784 26702 -8650
rect 26278 -8826 26292 -8786
rect 26232 -9042 26292 -8826
rect 26688 -8826 26702 -8784
rect 26736 -8784 26742 -8650
rect 27154 -8650 27200 -8638
rect 26736 -8826 26748 -8784
rect 26386 -8876 26594 -8870
rect 26386 -8910 26398 -8876
rect 26582 -8910 26594 -8876
rect 26386 -8916 26594 -8910
rect 26460 -9042 26520 -8916
rect 26232 -9102 26520 -9042
rect 26232 -9318 26292 -9102
rect 26460 -9228 26520 -9102
rect 26386 -9234 26594 -9228
rect 26386 -9268 26398 -9234
rect 26582 -9268 26594 -9234
rect 26386 -9274 26594 -9268
rect 26232 -9338 26244 -9318
rect 26238 -9464 26244 -9338
rect 26224 -9494 26244 -9464
rect 26278 -9338 26292 -9318
rect 26688 -9318 26748 -8826
rect 27154 -8826 27160 -8650
rect 27194 -8826 27200 -8650
rect 27154 -8838 27200 -8826
rect 27612 -8650 27658 -8638
rect 27612 -8826 27618 -8650
rect 27652 -8826 27658 -8650
rect 27612 -8838 27658 -8826
rect 28070 -8650 28116 -8638
rect 28070 -8826 28076 -8650
rect 28110 -8826 28116 -8650
rect 28070 -8838 28116 -8826
rect 28528 -8650 28574 -8638
rect 28528 -8826 28534 -8650
rect 28568 -8826 28574 -8650
rect 28528 -8838 28574 -8826
rect 28986 -8650 29032 -8638
rect 28986 -8826 28992 -8650
rect 29026 -8826 29032 -8650
rect 28986 -8838 29032 -8826
rect 29444 -8650 29490 -8638
rect 29444 -8826 29450 -8650
rect 29484 -8826 29490 -8650
rect 29444 -8838 29490 -8826
rect 29902 -8650 29948 -8638
rect 29902 -8826 29908 -8650
rect 29942 -8826 29948 -8650
rect 30352 -8650 30412 -8366
rect 30580 -8560 30640 -8214
rect 30508 -8566 30716 -8560
rect 30508 -8600 30520 -8566
rect 30704 -8600 30716 -8566
rect 30508 -8606 30716 -8600
rect 30352 -8680 30366 -8650
rect 29902 -8838 29948 -8826
rect 30360 -8826 30366 -8680
rect 30400 -8680 30412 -8650
rect 30812 -8650 30872 -8214
rect 30812 -8678 30824 -8650
rect 30400 -8826 30406 -8680
rect 30818 -8770 30824 -8678
rect 30360 -8838 30406 -8826
rect 30812 -8826 30824 -8770
rect 30858 -8678 30872 -8650
rect 31232 -8650 31292 -8214
rect 31466 -8560 31526 -8214
rect 31386 -8566 31594 -8560
rect 31386 -8600 31398 -8566
rect 31582 -8600 31594 -8566
rect 31386 -8606 31594 -8600
rect 30858 -8770 30864 -8678
rect 31232 -8686 31244 -8650
rect 30858 -8826 30872 -8770
rect 31238 -8790 31244 -8686
rect 26844 -8876 27052 -8870
rect 26844 -8910 26856 -8876
rect 27040 -8910 27052 -8876
rect 26844 -8916 27052 -8910
rect 27302 -8876 27510 -8870
rect 27302 -8910 27314 -8876
rect 27498 -8910 27510 -8876
rect 27302 -8916 27510 -8910
rect 27760 -8876 27968 -8870
rect 27760 -8910 27772 -8876
rect 27956 -8910 27968 -8876
rect 27760 -8916 27968 -8910
rect 28218 -8876 28426 -8870
rect 28218 -8910 28230 -8876
rect 28414 -8910 28426 -8876
rect 28218 -8916 28426 -8910
rect 28676 -8876 28884 -8870
rect 28676 -8910 28688 -8876
rect 28872 -8910 28884 -8876
rect 28676 -8916 28884 -8910
rect 29134 -8876 29342 -8870
rect 29134 -8910 29146 -8876
rect 29330 -8910 29342 -8876
rect 29134 -8916 29342 -8910
rect 29592 -8876 29800 -8870
rect 29592 -8910 29604 -8876
rect 29788 -8910 29800 -8876
rect 29592 -8916 29800 -8910
rect 30050 -8876 30258 -8870
rect 30050 -8910 30062 -8876
rect 30246 -8910 30258 -8876
rect 30050 -8916 30258 -8910
rect 30508 -8876 30716 -8870
rect 30508 -8910 30520 -8876
rect 30704 -8910 30716 -8876
rect 30508 -8916 30716 -8910
rect 26914 -8982 26974 -8916
rect 27376 -8982 27436 -8916
rect 27830 -8982 27890 -8916
rect 28292 -8982 28352 -8916
rect 28746 -8982 28806 -8916
rect 29196 -8982 29256 -8916
rect 29662 -8982 29722 -8916
rect 30118 -8982 30178 -8916
rect 26914 -9042 30178 -8982
rect 26920 -9162 30184 -9102
rect 26920 -9228 26980 -9162
rect 27382 -9228 27442 -9162
rect 27836 -9228 27896 -9162
rect 28298 -9228 28358 -9162
rect 28752 -9228 28812 -9162
rect 29202 -9228 29262 -9162
rect 29668 -9228 29728 -9162
rect 30124 -9228 30184 -9162
rect 30580 -9228 30640 -8916
rect 26844 -9234 27052 -9228
rect 26844 -9268 26856 -9234
rect 27040 -9268 27052 -9234
rect 26844 -9274 27052 -9268
rect 27302 -9234 27510 -9228
rect 27302 -9268 27314 -9234
rect 27498 -9268 27510 -9234
rect 27302 -9274 27510 -9268
rect 27760 -9234 27968 -9228
rect 27760 -9268 27772 -9234
rect 27956 -9268 27968 -9234
rect 27760 -9274 27968 -9268
rect 28218 -9234 28426 -9228
rect 28218 -9268 28230 -9234
rect 28414 -9268 28426 -9234
rect 28218 -9274 28426 -9268
rect 28676 -9234 28884 -9228
rect 28676 -9268 28688 -9234
rect 28872 -9268 28884 -9234
rect 28676 -9274 28884 -9268
rect 29134 -9234 29342 -9228
rect 29134 -9268 29146 -9234
rect 29330 -9268 29342 -9234
rect 29134 -9274 29342 -9268
rect 29592 -9234 29800 -9228
rect 29592 -9268 29604 -9234
rect 29788 -9268 29800 -9234
rect 29592 -9274 29800 -9268
rect 30050 -9234 30258 -9228
rect 30050 -9268 30062 -9234
rect 30246 -9268 30258 -9234
rect 30050 -9274 30258 -9268
rect 30508 -9234 30716 -9228
rect 30508 -9268 30520 -9234
rect 30704 -9268 30716 -9234
rect 30508 -9274 30716 -9268
rect 26278 -9494 26284 -9338
rect 26688 -9346 26702 -9318
rect 26224 -9874 26284 -9494
rect 26696 -9494 26702 -9346
rect 26736 -9346 26748 -9318
rect 27154 -9318 27200 -9306
rect 26736 -9494 26742 -9346
rect 26696 -9506 26742 -9494
rect 27154 -9494 27160 -9318
rect 27194 -9494 27200 -9318
rect 27154 -9506 27200 -9494
rect 27612 -9318 27658 -9306
rect 27612 -9494 27618 -9318
rect 27652 -9494 27658 -9318
rect 27612 -9506 27658 -9494
rect 28070 -9318 28116 -9306
rect 28070 -9494 28076 -9318
rect 28110 -9494 28116 -9318
rect 28070 -9506 28116 -9494
rect 28528 -9318 28574 -9306
rect 28528 -9494 28534 -9318
rect 28568 -9494 28574 -9318
rect 28528 -9506 28574 -9494
rect 28986 -9318 29032 -9306
rect 28986 -9494 28992 -9318
rect 29026 -9494 29032 -9318
rect 28986 -9506 29032 -9494
rect 29444 -9318 29490 -9306
rect 29444 -9494 29450 -9318
rect 29484 -9494 29490 -9318
rect 29444 -9506 29490 -9494
rect 29902 -9318 29948 -9306
rect 29902 -9494 29908 -9318
rect 29942 -9494 29948 -9318
rect 30360 -9318 30406 -9306
rect 30360 -9466 30366 -9318
rect 29902 -9506 29948 -9494
rect 30352 -9494 30366 -9466
rect 30400 -9466 30406 -9318
rect 30812 -9318 30872 -8826
rect 30400 -9494 30412 -9466
rect 26386 -9544 26594 -9538
rect 26386 -9578 26398 -9544
rect 26582 -9578 26594 -9544
rect 26386 -9584 26594 -9578
rect 26844 -9544 27052 -9538
rect 26844 -9578 26856 -9544
rect 27040 -9578 27052 -9544
rect 26844 -9584 27052 -9578
rect 27302 -9544 27510 -9538
rect 27302 -9578 27314 -9544
rect 27498 -9578 27510 -9544
rect 27302 -9584 27510 -9578
rect 27760 -9544 27968 -9538
rect 27760 -9578 27772 -9544
rect 27956 -9578 27968 -9544
rect 27760 -9584 27968 -9578
rect 28218 -9544 28426 -9538
rect 28218 -9578 28230 -9544
rect 28414 -9578 28426 -9544
rect 28218 -9584 28426 -9578
rect 28676 -9544 28884 -9538
rect 28676 -9578 28688 -9544
rect 28872 -9578 28884 -9544
rect 28676 -9584 28884 -9578
rect 29134 -9544 29342 -9538
rect 29134 -9578 29146 -9544
rect 29330 -9578 29342 -9544
rect 29134 -9584 29342 -9578
rect 29592 -9544 29800 -9538
rect 29592 -9578 29604 -9544
rect 29788 -9578 29800 -9544
rect 29592 -9584 29800 -9578
rect 30050 -9544 30258 -9538
rect 30050 -9578 30062 -9544
rect 30246 -9578 30258 -9544
rect 30050 -9584 30258 -9578
rect 26464 -9874 26524 -9584
rect 26914 -9650 26974 -9584
rect 27376 -9650 27436 -9584
rect 27830 -9650 27890 -9584
rect 28292 -9650 28352 -9584
rect 28746 -9650 28806 -9584
rect 29196 -9650 29256 -9584
rect 29662 -9650 29722 -9584
rect 30118 -9650 30178 -9584
rect 26974 -9710 30178 -9650
rect 26914 -9716 26974 -9710
rect 30352 -9874 30412 -9494
rect 30812 -9494 30824 -9318
rect 30858 -9494 30872 -9318
rect 30508 -9544 30716 -9538
rect 30508 -9578 30520 -9544
rect 30704 -9578 30716 -9544
rect 30508 -9584 30716 -9578
rect 30578 -9874 30638 -9584
rect 30812 -9874 30872 -9494
rect 31228 -8826 31244 -8790
rect 31278 -8686 31292 -8650
rect 31688 -8650 31748 -8214
rect 35346 -8354 35352 -8294
rect 35412 -8354 35418 -8294
rect 34192 -8434 34198 -8430
rect 31910 -8494 31916 -8434
rect 31976 -8436 34198 -8434
rect 31976 -8494 32378 -8436
rect 31916 -8560 31980 -8494
rect 32372 -8496 32378 -8494
rect 32438 -8494 32832 -8436
rect 32438 -8496 32444 -8494
rect 32826 -8496 32832 -8494
rect 32892 -8494 33294 -8436
rect 32892 -8496 32898 -8494
rect 33288 -8496 33294 -8494
rect 33354 -8494 33748 -8436
rect 33354 -8496 33360 -8494
rect 33742 -8496 33748 -8494
rect 33808 -8490 34198 -8436
rect 34258 -8434 34264 -8430
rect 34258 -8490 34664 -8434
rect 33808 -8494 34664 -8490
rect 34724 -8494 35120 -8434
rect 35180 -8494 35186 -8434
rect 33808 -8496 33814 -8494
rect 32378 -8560 32442 -8496
rect 32832 -8560 32896 -8496
rect 33294 -8560 33358 -8496
rect 33748 -8560 33812 -8496
rect 34198 -8560 34262 -8494
rect 34664 -8560 34728 -8494
rect 35120 -8560 35184 -8494
rect 31844 -8566 32052 -8560
rect 31844 -8600 31856 -8566
rect 32040 -8600 32052 -8566
rect 31844 -8606 32052 -8600
rect 32302 -8566 32510 -8560
rect 32302 -8600 32314 -8566
rect 32498 -8600 32510 -8566
rect 32302 -8606 32510 -8600
rect 32760 -8566 32968 -8560
rect 32760 -8600 32772 -8566
rect 32956 -8600 32968 -8566
rect 32760 -8606 32968 -8600
rect 33218 -8566 33426 -8560
rect 33218 -8600 33230 -8566
rect 33414 -8600 33426 -8566
rect 33218 -8606 33426 -8600
rect 33676 -8566 33884 -8560
rect 33676 -8600 33688 -8566
rect 33872 -8600 33884 -8566
rect 33676 -8606 33884 -8600
rect 34134 -8566 34342 -8560
rect 34134 -8600 34146 -8566
rect 34330 -8600 34342 -8566
rect 34134 -8606 34342 -8600
rect 34592 -8566 34800 -8560
rect 34592 -8600 34604 -8566
rect 34788 -8600 34800 -8566
rect 34592 -8606 34800 -8600
rect 35050 -8566 35258 -8560
rect 35050 -8600 35062 -8566
rect 35246 -8600 35258 -8566
rect 35050 -8606 35258 -8600
rect 31278 -8790 31284 -8686
rect 31688 -8714 31702 -8650
rect 31696 -8782 31702 -8714
rect 31278 -8826 31288 -8790
rect 31228 -8980 31288 -8826
rect 31688 -8826 31702 -8782
rect 31736 -8714 31748 -8650
rect 32154 -8650 32200 -8638
rect 31736 -8782 31742 -8714
rect 31736 -8826 31748 -8782
rect 31386 -8876 31594 -8870
rect 31386 -8910 31398 -8876
rect 31582 -8910 31594 -8876
rect 31386 -8916 31594 -8910
rect 31456 -8980 31516 -8916
rect 31688 -8980 31748 -8826
rect 32154 -8826 32160 -8650
rect 32194 -8826 32200 -8650
rect 32154 -8838 32200 -8826
rect 32612 -8650 32658 -8638
rect 32612 -8826 32618 -8650
rect 32652 -8826 32658 -8650
rect 32612 -8838 32658 -8826
rect 33070 -8650 33116 -8638
rect 33070 -8826 33076 -8650
rect 33110 -8826 33116 -8650
rect 33070 -8838 33116 -8826
rect 33528 -8650 33574 -8638
rect 33528 -8826 33534 -8650
rect 33568 -8826 33574 -8650
rect 33528 -8838 33574 -8826
rect 33986 -8650 34032 -8638
rect 33986 -8826 33992 -8650
rect 34026 -8826 34032 -8650
rect 33986 -8838 34032 -8826
rect 34444 -8650 34490 -8638
rect 34444 -8826 34450 -8650
rect 34484 -8826 34490 -8650
rect 34444 -8838 34490 -8826
rect 34902 -8650 34948 -8638
rect 34902 -8826 34908 -8650
rect 34942 -8826 34948 -8650
rect 35352 -8650 35412 -8354
rect 35592 -8560 35652 -8214
rect 35508 -8566 35716 -8560
rect 35508 -8600 35520 -8566
rect 35704 -8600 35716 -8566
rect 35508 -8606 35716 -8600
rect 35352 -8692 35366 -8650
rect 34902 -8838 34948 -8826
rect 35360 -8826 35366 -8692
rect 35400 -8692 35412 -8650
rect 35810 -8650 35870 -8214
rect 35810 -8690 35824 -8650
rect 35400 -8826 35406 -8692
rect 35818 -8780 35824 -8690
rect 35360 -8838 35406 -8826
rect 35808 -8826 35824 -8780
rect 35858 -8690 35870 -8650
rect 36156 -8338 36268 -8214
rect 35858 -8780 35864 -8690
rect 35858 -8826 35868 -8780
rect 31844 -8876 32052 -8870
rect 31844 -8910 31856 -8876
rect 32040 -8910 32052 -8876
rect 31844 -8916 32052 -8910
rect 32302 -8876 32510 -8870
rect 32302 -8910 32314 -8876
rect 32498 -8910 32510 -8876
rect 32302 -8916 32510 -8910
rect 32760 -8876 32968 -8870
rect 32760 -8910 32772 -8876
rect 32956 -8910 32968 -8876
rect 32760 -8916 32968 -8910
rect 33218 -8876 33426 -8870
rect 33218 -8910 33230 -8876
rect 33414 -8910 33426 -8876
rect 33218 -8916 33426 -8910
rect 33676 -8876 33884 -8870
rect 33676 -8910 33688 -8876
rect 33872 -8910 33884 -8876
rect 33676 -8916 33884 -8910
rect 34134 -8876 34342 -8870
rect 34134 -8910 34146 -8876
rect 34330 -8910 34342 -8876
rect 34134 -8916 34342 -8910
rect 34592 -8876 34800 -8870
rect 34592 -8910 34604 -8876
rect 34788 -8910 34800 -8876
rect 34592 -8916 34800 -8910
rect 35050 -8876 35258 -8870
rect 35050 -8910 35062 -8876
rect 35246 -8910 35258 -8876
rect 35050 -8916 35258 -8910
rect 35508 -8876 35716 -8870
rect 35508 -8910 35520 -8876
rect 35704 -8910 35716 -8876
rect 35508 -8916 35716 -8910
rect 31228 -9040 31748 -8980
rect 31228 -9874 31288 -9040
rect 31456 -9874 31516 -9040
rect 31688 -9874 31748 -9040
rect 31914 -8982 31974 -8916
rect 32376 -8982 32436 -8916
rect 32830 -8982 32890 -8916
rect 33292 -8982 33352 -8916
rect 33746 -8982 33806 -8916
rect 34196 -8982 34256 -8916
rect 34662 -8982 34722 -8916
rect 35118 -8982 35178 -8916
rect 31914 -9042 35178 -8982
rect 35582 -9874 35642 -8916
rect 35808 -9874 35868 -8826
rect 26160 -9902 35930 -9874
rect 26160 -9988 26210 -9902
rect 26306 -9988 26790 -9902
rect 26886 -9988 27390 -9902
rect 27486 -9988 27990 -9902
rect 28086 -9988 28590 -9902
rect 28686 -9988 29190 -9902
rect 29286 -9988 29790 -9902
rect 29886 -9988 30390 -9902
rect 30486 -9988 30990 -9902
rect 31086 -9988 31590 -9902
rect 31686 -9988 32190 -9902
rect 32286 -9988 32790 -9902
rect 32886 -9988 33390 -9902
rect 33486 -9988 33990 -9902
rect 34086 -9988 34590 -9902
rect 34686 -9988 35190 -9902
rect 35286 -9988 35790 -9902
rect 35886 -9988 35930 -9902
rect 26160 -10018 35930 -9988
rect 25812 -10466 25924 -10342
rect 26524 -10466 26534 -10166
rect 35546 -10466 35556 -10166
rect 36156 -10342 36162 -8338
rect 36262 -10342 36268 -8338
rect 36156 -10466 36268 -10342
rect 25812 -10472 36268 -10466
rect 25812 -10572 25918 -10472
rect 36162 -10572 36268 -10472
rect 25812 -10578 36268 -10572
rect 25400 -23300 25406 -23240
rect 25466 -23300 25472 -23240
rect 21156 -25766 21268 -25590
rect 10812 -25772 21268 -25766
rect 10812 -25872 10918 -25772
rect 21162 -25872 21268 -25772
rect 10812 -25878 21268 -25872
rect 10812 -26108 21268 -26102
rect 10812 -26208 10918 -26108
rect 21162 -26208 21268 -26108
rect 10812 -26214 21268 -26208
rect 10812 -26338 10924 -26214
rect 10812 -28342 10818 -26338
rect 10918 -28342 10924 -26338
rect 11232 -26650 11292 -26214
rect 11462 -26560 11522 -26214
rect 15352 -26306 15412 -26300
rect 11920 -26440 12376 -26434
rect 11908 -26500 11914 -26440
rect 11974 -26494 12376 -26440
rect 12436 -26440 13292 -26434
rect 12436 -26494 12830 -26440
rect 11974 -26500 11980 -26494
rect 11914 -26560 11980 -26500
rect 12376 -26560 12442 -26494
rect 12824 -26500 12830 -26494
rect 12890 -26494 13292 -26440
rect 13352 -26494 13746 -26434
rect 13806 -26494 14196 -26434
rect 14256 -26440 15118 -26434
rect 14256 -26494 14662 -26440
rect 12890 -26500 12896 -26494
rect 12830 -26560 12896 -26500
rect 13292 -26560 13358 -26494
rect 13746 -26560 13812 -26494
rect 14196 -26560 14262 -26494
rect 14656 -26500 14662 -26494
rect 14722 -26494 15118 -26440
rect 15178 -26494 15184 -26434
rect 14722 -26500 14728 -26494
rect 14662 -26560 14728 -26500
rect 15118 -26560 15184 -26494
rect 11386 -26566 11594 -26560
rect 11386 -26600 11398 -26566
rect 11582 -26600 11594 -26566
rect 11386 -26606 11594 -26600
rect 11844 -26566 12052 -26560
rect 11844 -26600 11856 -26566
rect 12040 -26600 12052 -26566
rect 11844 -26606 12052 -26600
rect 12302 -26566 12510 -26560
rect 12302 -26600 12314 -26566
rect 12498 -26600 12510 -26566
rect 12302 -26606 12510 -26600
rect 12760 -26566 12968 -26560
rect 12760 -26600 12772 -26566
rect 12956 -26600 12968 -26566
rect 12760 -26606 12968 -26600
rect 13218 -26566 13426 -26560
rect 13218 -26600 13230 -26566
rect 13414 -26600 13426 -26566
rect 13218 -26606 13426 -26600
rect 13676 -26566 13884 -26560
rect 13676 -26600 13688 -26566
rect 13872 -26600 13884 -26566
rect 13676 -26606 13884 -26600
rect 14134 -26566 14342 -26560
rect 14134 -26600 14146 -26566
rect 14330 -26600 14342 -26566
rect 14134 -26606 14342 -26600
rect 14592 -26566 14800 -26560
rect 14592 -26600 14604 -26566
rect 14788 -26600 14800 -26566
rect 14592 -26606 14800 -26600
rect 15050 -26566 15258 -26560
rect 15050 -26600 15062 -26566
rect 15246 -26600 15258 -26566
rect 15050 -26606 15258 -26600
rect 11232 -26690 11244 -26650
rect 11238 -26786 11244 -26690
rect 11232 -26826 11244 -26786
rect 11278 -26690 11292 -26650
rect 11696 -26650 11742 -26638
rect 11278 -26786 11284 -26690
rect 11696 -26784 11702 -26650
rect 11278 -26826 11292 -26786
rect 11232 -27042 11292 -26826
rect 11688 -26826 11702 -26784
rect 11736 -26784 11742 -26650
rect 12154 -26650 12200 -26638
rect 11736 -26826 11748 -26784
rect 11386 -26876 11594 -26870
rect 11386 -26910 11398 -26876
rect 11582 -26910 11594 -26876
rect 11386 -26916 11594 -26910
rect 11460 -27042 11520 -26916
rect 11232 -27102 11520 -27042
rect 11232 -27318 11292 -27102
rect 11460 -27228 11520 -27102
rect 11386 -27234 11594 -27228
rect 11386 -27268 11398 -27234
rect 11582 -27268 11594 -27234
rect 11386 -27274 11594 -27268
rect 11232 -27338 11244 -27318
rect 11238 -27464 11244 -27338
rect 11224 -27494 11244 -27464
rect 11278 -27338 11292 -27318
rect 11688 -27318 11748 -26826
rect 12154 -26826 12160 -26650
rect 12194 -26826 12200 -26650
rect 12154 -26838 12200 -26826
rect 12612 -26650 12658 -26638
rect 12612 -26826 12618 -26650
rect 12652 -26826 12658 -26650
rect 12612 -26838 12658 -26826
rect 13070 -26650 13116 -26638
rect 13070 -26826 13076 -26650
rect 13110 -26826 13116 -26650
rect 13070 -26838 13116 -26826
rect 13528 -26650 13574 -26638
rect 13528 -26826 13534 -26650
rect 13568 -26826 13574 -26650
rect 13528 -26838 13574 -26826
rect 13986 -26650 14032 -26638
rect 13986 -26826 13992 -26650
rect 14026 -26826 14032 -26650
rect 13986 -26838 14032 -26826
rect 14444 -26650 14490 -26638
rect 14444 -26826 14450 -26650
rect 14484 -26826 14490 -26650
rect 14444 -26838 14490 -26826
rect 14902 -26650 14948 -26638
rect 14902 -26826 14908 -26650
rect 14942 -26826 14948 -26650
rect 15352 -26650 15412 -26366
rect 15580 -26560 15640 -26214
rect 15508 -26566 15716 -26560
rect 15508 -26600 15520 -26566
rect 15704 -26600 15716 -26566
rect 15508 -26606 15716 -26600
rect 15352 -26680 15366 -26650
rect 14902 -26838 14948 -26826
rect 15360 -26826 15366 -26680
rect 15400 -26680 15412 -26650
rect 15812 -26650 15872 -26214
rect 15812 -26678 15824 -26650
rect 15400 -26826 15406 -26680
rect 15818 -26770 15824 -26678
rect 15360 -26838 15406 -26826
rect 15812 -26826 15824 -26770
rect 15858 -26678 15872 -26650
rect 16232 -26650 16292 -26214
rect 16466 -26560 16526 -26214
rect 16386 -26566 16594 -26560
rect 16386 -26600 16398 -26566
rect 16582 -26600 16594 -26566
rect 16386 -26606 16594 -26600
rect 15858 -26770 15864 -26678
rect 16232 -26686 16244 -26650
rect 15858 -26826 15872 -26770
rect 16238 -26790 16244 -26686
rect 11844 -26876 12052 -26870
rect 11844 -26910 11856 -26876
rect 12040 -26910 12052 -26876
rect 11844 -26916 12052 -26910
rect 12302 -26876 12510 -26870
rect 12302 -26910 12314 -26876
rect 12498 -26910 12510 -26876
rect 12302 -26916 12510 -26910
rect 12760 -26876 12968 -26870
rect 12760 -26910 12772 -26876
rect 12956 -26910 12968 -26876
rect 12760 -26916 12968 -26910
rect 13218 -26876 13426 -26870
rect 13218 -26910 13230 -26876
rect 13414 -26910 13426 -26876
rect 13218 -26916 13426 -26910
rect 13676 -26876 13884 -26870
rect 13676 -26910 13688 -26876
rect 13872 -26910 13884 -26876
rect 13676 -26916 13884 -26910
rect 14134 -26876 14342 -26870
rect 14134 -26910 14146 -26876
rect 14330 -26910 14342 -26876
rect 14134 -26916 14342 -26910
rect 14592 -26876 14800 -26870
rect 14592 -26910 14604 -26876
rect 14788 -26910 14800 -26876
rect 14592 -26916 14800 -26910
rect 15050 -26876 15258 -26870
rect 15050 -26910 15062 -26876
rect 15246 -26910 15258 -26876
rect 15050 -26916 15258 -26910
rect 15508 -26876 15716 -26870
rect 15508 -26910 15520 -26876
rect 15704 -26910 15716 -26876
rect 15508 -26916 15716 -26910
rect 11914 -26982 11974 -26916
rect 12376 -26982 12436 -26916
rect 12830 -26982 12890 -26916
rect 13292 -26982 13352 -26916
rect 13746 -26982 13806 -26916
rect 14196 -26982 14256 -26916
rect 14662 -26982 14722 -26916
rect 15118 -26982 15178 -26916
rect 11914 -27042 15178 -26982
rect 11920 -27162 15184 -27102
rect 11920 -27228 11980 -27162
rect 12382 -27228 12442 -27162
rect 12836 -27228 12896 -27162
rect 13298 -27228 13358 -27162
rect 13752 -27228 13812 -27162
rect 14202 -27228 14262 -27162
rect 14668 -27228 14728 -27162
rect 15124 -27228 15184 -27162
rect 15580 -27228 15640 -26916
rect 11844 -27234 12052 -27228
rect 11844 -27268 11856 -27234
rect 12040 -27268 12052 -27234
rect 11844 -27274 12052 -27268
rect 12302 -27234 12510 -27228
rect 12302 -27268 12314 -27234
rect 12498 -27268 12510 -27234
rect 12302 -27274 12510 -27268
rect 12760 -27234 12968 -27228
rect 12760 -27268 12772 -27234
rect 12956 -27268 12968 -27234
rect 12760 -27274 12968 -27268
rect 13218 -27234 13426 -27228
rect 13218 -27268 13230 -27234
rect 13414 -27268 13426 -27234
rect 13218 -27274 13426 -27268
rect 13676 -27234 13884 -27228
rect 13676 -27268 13688 -27234
rect 13872 -27268 13884 -27234
rect 13676 -27274 13884 -27268
rect 14134 -27234 14342 -27228
rect 14134 -27268 14146 -27234
rect 14330 -27268 14342 -27234
rect 14134 -27274 14342 -27268
rect 14592 -27234 14800 -27228
rect 14592 -27268 14604 -27234
rect 14788 -27268 14800 -27234
rect 14592 -27274 14800 -27268
rect 15050 -27234 15258 -27228
rect 15050 -27268 15062 -27234
rect 15246 -27268 15258 -27234
rect 15050 -27274 15258 -27268
rect 15508 -27234 15716 -27228
rect 15508 -27268 15520 -27234
rect 15704 -27268 15716 -27234
rect 15508 -27274 15716 -27268
rect 11278 -27494 11284 -27338
rect 11688 -27346 11702 -27318
rect 11224 -27874 11284 -27494
rect 11696 -27494 11702 -27346
rect 11736 -27346 11748 -27318
rect 12154 -27318 12200 -27306
rect 11736 -27494 11742 -27346
rect 11696 -27506 11742 -27494
rect 12154 -27494 12160 -27318
rect 12194 -27494 12200 -27318
rect 12154 -27506 12200 -27494
rect 12612 -27318 12658 -27306
rect 12612 -27494 12618 -27318
rect 12652 -27494 12658 -27318
rect 12612 -27506 12658 -27494
rect 13070 -27318 13116 -27306
rect 13070 -27494 13076 -27318
rect 13110 -27494 13116 -27318
rect 13070 -27506 13116 -27494
rect 13528 -27318 13574 -27306
rect 13528 -27494 13534 -27318
rect 13568 -27494 13574 -27318
rect 13528 -27506 13574 -27494
rect 13986 -27318 14032 -27306
rect 13986 -27494 13992 -27318
rect 14026 -27494 14032 -27318
rect 13986 -27506 14032 -27494
rect 14444 -27318 14490 -27306
rect 14444 -27494 14450 -27318
rect 14484 -27494 14490 -27318
rect 14444 -27506 14490 -27494
rect 14902 -27318 14948 -27306
rect 14902 -27494 14908 -27318
rect 14942 -27494 14948 -27318
rect 15360 -27318 15406 -27306
rect 15360 -27466 15366 -27318
rect 14902 -27506 14948 -27494
rect 15352 -27494 15366 -27466
rect 15400 -27466 15406 -27318
rect 15812 -27318 15872 -26826
rect 15400 -27494 15412 -27466
rect 11386 -27544 11594 -27538
rect 11386 -27578 11398 -27544
rect 11582 -27578 11594 -27544
rect 11386 -27584 11594 -27578
rect 11844 -27544 12052 -27538
rect 11844 -27578 11856 -27544
rect 12040 -27578 12052 -27544
rect 11844 -27584 12052 -27578
rect 12302 -27544 12510 -27538
rect 12302 -27578 12314 -27544
rect 12498 -27578 12510 -27544
rect 12302 -27584 12510 -27578
rect 12760 -27544 12968 -27538
rect 12760 -27578 12772 -27544
rect 12956 -27578 12968 -27544
rect 12760 -27584 12968 -27578
rect 13218 -27544 13426 -27538
rect 13218 -27578 13230 -27544
rect 13414 -27578 13426 -27544
rect 13218 -27584 13426 -27578
rect 13676 -27544 13884 -27538
rect 13676 -27578 13688 -27544
rect 13872 -27578 13884 -27544
rect 13676 -27584 13884 -27578
rect 14134 -27544 14342 -27538
rect 14134 -27578 14146 -27544
rect 14330 -27578 14342 -27544
rect 14134 -27584 14342 -27578
rect 14592 -27544 14800 -27538
rect 14592 -27578 14604 -27544
rect 14788 -27578 14800 -27544
rect 14592 -27584 14800 -27578
rect 15050 -27544 15258 -27538
rect 15050 -27578 15062 -27544
rect 15246 -27578 15258 -27544
rect 15050 -27584 15258 -27578
rect 11464 -27874 11524 -27584
rect 11914 -27650 11974 -27584
rect 12376 -27650 12436 -27584
rect 12830 -27650 12890 -27584
rect 13292 -27650 13352 -27584
rect 13746 -27650 13806 -27584
rect 14196 -27650 14256 -27584
rect 14662 -27650 14722 -27584
rect 15118 -27650 15178 -27584
rect 11914 -27710 15118 -27650
rect 15118 -27716 15178 -27710
rect 15352 -27874 15412 -27494
rect 15812 -27494 15824 -27318
rect 15858 -27494 15872 -27318
rect 15508 -27544 15716 -27538
rect 15508 -27578 15520 -27544
rect 15704 -27578 15716 -27544
rect 15508 -27584 15716 -27578
rect 15578 -27874 15638 -27584
rect 15812 -27874 15872 -27494
rect 16228 -26826 16244 -26790
rect 16278 -26686 16292 -26650
rect 16688 -26650 16748 -26214
rect 20346 -26354 20352 -26294
rect 20412 -26354 20418 -26294
rect 19192 -26434 19198 -26430
rect 16910 -26494 16916 -26434
rect 16976 -26436 19198 -26434
rect 16976 -26494 17378 -26436
rect 16916 -26560 16980 -26494
rect 17372 -26496 17378 -26494
rect 17438 -26494 17832 -26436
rect 17438 -26496 17444 -26494
rect 17826 -26496 17832 -26494
rect 17892 -26494 18294 -26436
rect 17892 -26496 17898 -26494
rect 18288 -26496 18294 -26494
rect 18354 -26494 18748 -26436
rect 18354 -26496 18360 -26494
rect 18742 -26496 18748 -26494
rect 18808 -26490 19198 -26436
rect 19258 -26434 19264 -26430
rect 19258 -26490 19664 -26434
rect 18808 -26494 19664 -26490
rect 19724 -26494 20120 -26434
rect 20180 -26494 20186 -26434
rect 18808 -26496 18814 -26494
rect 17378 -26560 17442 -26496
rect 17832 -26560 17896 -26496
rect 18294 -26560 18358 -26496
rect 18748 -26560 18812 -26496
rect 19198 -26560 19262 -26494
rect 19664 -26560 19728 -26494
rect 20120 -26560 20184 -26494
rect 16844 -26566 17052 -26560
rect 16844 -26600 16856 -26566
rect 17040 -26600 17052 -26566
rect 16844 -26606 17052 -26600
rect 17302 -26566 17510 -26560
rect 17302 -26600 17314 -26566
rect 17498 -26600 17510 -26566
rect 17302 -26606 17510 -26600
rect 17760 -26566 17968 -26560
rect 17760 -26600 17772 -26566
rect 17956 -26600 17968 -26566
rect 17760 -26606 17968 -26600
rect 18218 -26566 18426 -26560
rect 18218 -26600 18230 -26566
rect 18414 -26600 18426 -26566
rect 18218 -26606 18426 -26600
rect 18676 -26566 18884 -26560
rect 18676 -26600 18688 -26566
rect 18872 -26600 18884 -26566
rect 18676 -26606 18884 -26600
rect 19134 -26566 19342 -26560
rect 19134 -26600 19146 -26566
rect 19330 -26600 19342 -26566
rect 19134 -26606 19342 -26600
rect 19592 -26566 19800 -26560
rect 19592 -26600 19604 -26566
rect 19788 -26600 19800 -26566
rect 19592 -26606 19800 -26600
rect 20050 -26566 20258 -26560
rect 20050 -26600 20062 -26566
rect 20246 -26600 20258 -26566
rect 20050 -26606 20258 -26600
rect 16278 -26790 16284 -26686
rect 16688 -26714 16702 -26650
rect 16696 -26782 16702 -26714
rect 16278 -26826 16288 -26790
rect 16228 -26980 16288 -26826
rect 16688 -26826 16702 -26782
rect 16736 -26714 16748 -26650
rect 17154 -26650 17200 -26638
rect 16736 -26782 16742 -26714
rect 16736 -26826 16748 -26782
rect 16386 -26876 16594 -26870
rect 16386 -26910 16398 -26876
rect 16582 -26910 16594 -26876
rect 16386 -26916 16594 -26910
rect 16456 -26980 16516 -26916
rect 16688 -26980 16748 -26826
rect 17154 -26826 17160 -26650
rect 17194 -26826 17200 -26650
rect 17154 -26838 17200 -26826
rect 17612 -26650 17658 -26638
rect 17612 -26826 17618 -26650
rect 17652 -26826 17658 -26650
rect 17612 -26838 17658 -26826
rect 18070 -26650 18116 -26638
rect 18070 -26826 18076 -26650
rect 18110 -26826 18116 -26650
rect 18070 -26838 18116 -26826
rect 18528 -26650 18574 -26638
rect 18528 -26826 18534 -26650
rect 18568 -26826 18574 -26650
rect 18528 -26838 18574 -26826
rect 18986 -26650 19032 -26638
rect 18986 -26826 18992 -26650
rect 19026 -26826 19032 -26650
rect 18986 -26838 19032 -26826
rect 19444 -26650 19490 -26638
rect 19444 -26826 19450 -26650
rect 19484 -26826 19490 -26650
rect 19444 -26838 19490 -26826
rect 19902 -26650 19948 -26638
rect 19902 -26826 19908 -26650
rect 19942 -26826 19948 -26650
rect 20352 -26650 20412 -26354
rect 20592 -26560 20652 -26214
rect 20508 -26566 20716 -26560
rect 20508 -26600 20520 -26566
rect 20704 -26600 20716 -26566
rect 20508 -26606 20716 -26600
rect 20352 -26692 20366 -26650
rect 19902 -26838 19948 -26826
rect 20360 -26826 20366 -26692
rect 20400 -26692 20412 -26650
rect 20810 -26650 20870 -26214
rect 20810 -26690 20824 -26650
rect 20400 -26826 20406 -26692
rect 20818 -26780 20824 -26690
rect 20360 -26838 20406 -26826
rect 20808 -26826 20824 -26780
rect 20858 -26690 20870 -26650
rect 21156 -26338 21268 -26214
rect 20858 -26780 20864 -26690
rect 20858 -26826 20868 -26780
rect 16844 -26876 17052 -26870
rect 16844 -26910 16856 -26876
rect 17040 -26910 17052 -26876
rect 16844 -26916 17052 -26910
rect 17302 -26876 17510 -26870
rect 17302 -26910 17314 -26876
rect 17498 -26910 17510 -26876
rect 17302 -26916 17510 -26910
rect 17760 -26876 17968 -26870
rect 17760 -26910 17772 -26876
rect 17956 -26910 17968 -26876
rect 17760 -26916 17968 -26910
rect 18218 -26876 18426 -26870
rect 18218 -26910 18230 -26876
rect 18414 -26910 18426 -26876
rect 18218 -26916 18426 -26910
rect 18676 -26876 18884 -26870
rect 18676 -26910 18688 -26876
rect 18872 -26910 18884 -26876
rect 18676 -26916 18884 -26910
rect 19134 -26876 19342 -26870
rect 19134 -26910 19146 -26876
rect 19330 -26910 19342 -26876
rect 19134 -26916 19342 -26910
rect 19592 -26876 19800 -26870
rect 19592 -26910 19604 -26876
rect 19788 -26910 19800 -26876
rect 19592 -26916 19800 -26910
rect 20050 -26876 20258 -26870
rect 20050 -26910 20062 -26876
rect 20246 -26910 20258 -26876
rect 20050 -26916 20258 -26910
rect 20508 -26876 20716 -26870
rect 20508 -26910 20520 -26876
rect 20704 -26910 20716 -26876
rect 20508 -26916 20716 -26910
rect 16228 -27040 16748 -26980
rect 16228 -27874 16288 -27040
rect 16456 -27874 16516 -27040
rect 16688 -27874 16748 -27040
rect 16914 -26982 16974 -26916
rect 17376 -26982 17436 -26916
rect 17830 -26982 17890 -26916
rect 18292 -26982 18352 -26916
rect 18746 -26982 18806 -26916
rect 19196 -26982 19256 -26916
rect 19662 -26982 19722 -26916
rect 20118 -26982 20178 -26916
rect 16914 -27042 20178 -26982
rect 20582 -27874 20642 -26916
rect 20808 -27874 20868 -26826
rect 11160 -27902 20930 -27874
rect 11160 -27988 11210 -27902
rect 11306 -27988 11790 -27902
rect 11886 -27988 12390 -27902
rect 12486 -27988 12990 -27902
rect 13086 -27988 13590 -27902
rect 13686 -27988 14190 -27902
rect 14286 -27988 14790 -27902
rect 14886 -27988 15390 -27902
rect 15486 -27988 15990 -27902
rect 16086 -27988 16590 -27902
rect 16686 -27988 17190 -27902
rect 17286 -27988 17790 -27902
rect 17886 -27988 18390 -27902
rect 18486 -27988 18990 -27902
rect 19086 -27988 19590 -27902
rect 19686 -27988 20190 -27902
rect 20286 -27988 20790 -27902
rect 20886 -27988 20930 -27902
rect 11160 -28018 20930 -27988
rect 10812 -28466 10924 -28342
rect 11524 -28466 11534 -28166
rect 20546 -28466 20556 -28166
rect 21156 -28342 21162 -26338
rect 21262 -28342 21268 -26338
rect 25546 -27650 25606 -11954
rect 29766 -11032 40222 -11026
rect 29766 -11132 29872 -11032
rect 40116 -11132 40222 -11032
rect 29766 -11138 40222 -11132
rect 29766 -11262 29878 -11138
rect 29766 -13266 29772 -11262
rect 29872 -13266 29878 -11262
rect 30478 -11438 30488 -11138
rect 39500 -11438 39510 -11138
rect 40110 -11262 40222 -11138
rect 30104 -11616 39874 -11586
rect 30104 -11702 30148 -11616
rect 30244 -11702 30748 -11616
rect 30844 -11702 31348 -11616
rect 31444 -11702 31948 -11616
rect 32044 -11702 32548 -11616
rect 32644 -11702 33148 -11616
rect 33244 -11702 33748 -11616
rect 33844 -11702 34348 -11616
rect 34444 -11702 34948 -11616
rect 35044 -11702 35548 -11616
rect 35644 -11702 36148 -11616
rect 36244 -11702 36748 -11616
rect 36844 -11702 37348 -11616
rect 37444 -11702 37948 -11616
rect 38044 -11702 38548 -11616
rect 38644 -11702 39148 -11616
rect 39244 -11702 39728 -11616
rect 39824 -11702 39874 -11616
rect 30104 -11730 39874 -11702
rect 30166 -12778 30226 -11730
rect 30392 -12688 30452 -11730
rect 30856 -12622 34120 -12562
rect 30856 -12688 30916 -12622
rect 31312 -12688 31372 -12622
rect 31778 -12688 31838 -12622
rect 32228 -12688 32288 -12622
rect 32682 -12688 32742 -12622
rect 33144 -12688 33204 -12622
rect 33598 -12688 33658 -12622
rect 34060 -12688 34120 -12622
rect 34286 -12564 34346 -11730
rect 34518 -12564 34578 -11730
rect 34746 -12564 34806 -11730
rect 34286 -12624 34806 -12564
rect 30318 -12694 30526 -12688
rect 30318 -12728 30330 -12694
rect 30514 -12728 30526 -12694
rect 30318 -12734 30526 -12728
rect 30776 -12694 30984 -12688
rect 30776 -12728 30788 -12694
rect 30972 -12728 30984 -12694
rect 30776 -12734 30984 -12728
rect 31234 -12694 31442 -12688
rect 31234 -12728 31246 -12694
rect 31430 -12728 31442 -12694
rect 31234 -12734 31442 -12728
rect 31692 -12694 31900 -12688
rect 31692 -12728 31704 -12694
rect 31888 -12728 31900 -12694
rect 31692 -12734 31900 -12728
rect 32150 -12694 32358 -12688
rect 32150 -12728 32162 -12694
rect 32346 -12728 32358 -12694
rect 32150 -12734 32358 -12728
rect 32608 -12694 32816 -12688
rect 32608 -12728 32620 -12694
rect 32804 -12728 32816 -12694
rect 32608 -12734 32816 -12728
rect 33066 -12694 33274 -12688
rect 33066 -12728 33078 -12694
rect 33262 -12728 33274 -12694
rect 33066 -12734 33274 -12728
rect 33524 -12694 33732 -12688
rect 33524 -12728 33536 -12694
rect 33720 -12728 33732 -12694
rect 33524 -12734 33732 -12728
rect 33982 -12694 34190 -12688
rect 33982 -12728 33994 -12694
rect 34178 -12728 34190 -12694
rect 33982 -12734 34190 -12728
rect 30166 -12824 30176 -12778
rect 30170 -12914 30176 -12824
rect 29766 -13390 29878 -13266
rect 30164 -12954 30176 -12914
rect 30210 -12824 30226 -12778
rect 30628 -12778 30674 -12766
rect 30210 -12914 30216 -12824
rect 30628 -12912 30634 -12778
rect 30210 -12954 30224 -12914
rect 30164 -13390 30224 -12954
rect 30622 -12954 30634 -12912
rect 30668 -12912 30674 -12778
rect 31086 -12778 31132 -12766
rect 30668 -12954 30682 -12912
rect 30318 -13004 30526 -12998
rect 30318 -13038 30330 -13004
rect 30514 -13038 30526 -13004
rect 30318 -13044 30526 -13038
rect 30382 -13390 30442 -13044
rect 30622 -13250 30682 -12954
rect 31086 -12954 31092 -12778
rect 31126 -12954 31132 -12778
rect 31086 -12966 31132 -12954
rect 31544 -12778 31590 -12766
rect 31544 -12954 31550 -12778
rect 31584 -12954 31590 -12778
rect 31544 -12966 31590 -12954
rect 32002 -12778 32048 -12766
rect 32002 -12954 32008 -12778
rect 32042 -12954 32048 -12778
rect 32002 -12966 32048 -12954
rect 32460 -12778 32506 -12766
rect 32460 -12954 32466 -12778
rect 32500 -12954 32506 -12778
rect 32460 -12966 32506 -12954
rect 32918 -12778 32964 -12766
rect 32918 -12954 32924 -12778
rect 32958 -12954 32964 -12778
rect 32918 -12966 32964 -12954
rect 33376 -12778 33422 -12766
rect 33376 -12954 33382 -12778
rect 33416 -12954 33422 -12778
rect 33376 -12966 33422 -12954
rect 33834 -12778 33880 -12766
rect 33834 -12954 33840 -12778
rect 33874 -12954 33880 -12778
rect 34286 -12778 34346 -12624
rect 34518 -12688 34578 -12624
rect 34440 -12694 34648 -12688
rect 34440 -12728 34452 -12694
rect 34636 -12728 34648 -12694
rect 34440 -12734 34648 -12728
rect 34286 -12822 34298 -12778
rect 34292 -12890 34298 -12822
rect 33834 -12966 33880 -12954
rect 34286 -12954 34298 -12890
rect 34332 -12822 34346 -12778
rect 34746 -12778 34806 -12624
rect 34746 -12814 34756 -12778
rect 34332 -12890 34338 -12822
rect 34332 -12954 34346 -12890
rect 34750 -12918 34756 -12814
rect 30776 -13004 30984 -12998
rect 30776 -13038 30788 -13004
rect 30972 -13038 30984 -13004
rect 30776 -13044 30984 -13038
rect 31234 -13004 31442 -12998
rect 31234 -13038 31246 -13004
rect 31430 -13038 31442 -13004
rect 31234 -13044 31442 -13038
rect 31692 -13004 31900 -12998
rect 31692 -13038 31704 -13004
rect 31888 -13038 31900 -13004
rect 31692 -13044 31900 -13038
rect 32150 -13004 32358 -12998
rect 32150 -13038 32162 -13004
rect 32346 -13038 32358 -13004
rect 32150 -13044 32358 -13038
rect 32608 -13004 32816 -12998
rect 32608 -13038 32620 -13004
rect 32804 -13038 32816 -13004
rect 32608 -13044 32816 -13038
rect 33066 -13004 33274 -12998
rect 33066 -13038 33078 -13004
rect 33262 -13038 33274 -13004
rect 33066 -13044 33274 -13038
rect 33524 -13004 33732 -12998
rect 33524 -13038 33536 -13004
rect 33720 -13038 33732 -13004
rect 33524 -13044 33732 -13038
rect 33982 -13004 34190 -12998
rect 33982 -13038 33994 -13004
rect 34178 -13038 34190 -13004
rect 33982 -13044 34190 -13038
rect 30850 -13110 30914 -13044
rect 31306 -13110 31370 -13044
rect 31772 -13110 31836 -13044
rect 32222 -13108 32286 -13044
rect 32676 -13108 32740 -13044
rect 33138 -13108 33202 -13044
rect 33592 -13108 33656 -13044
rect 32220 -13110 32226 -13108
rect 30848 -13170 30854 -13110
rect 30914 -13170 31310 -13110
rect 31370 -13114 32226 -13110
rect 31370 -13170 31776 -13114
rect 31770 -13174 31776 -13170
rect 31836 -13168 32226 -13114
rect 32286 -13110 32292 -13108
rect 32674 -13110 32680 -13108
rect 32286 -13168 32680 -13110
rect 32740 -13110 32746 -13108
rect 33136 -13110 33142 -13108
rect 32740 -13168 33142 -13110
rect 33202 -13110 33208 -13108
rect 33590 -13110 33596 -13108
rect 33202 -13168 33596 -13110
rect 33656 -13110 33662 -13108
rect 34054 -13110 34118 -13044
rect 33656 -13168 34058 -13110
rect 31836 -13170 34058 -13168
rect 34118 -13170 34124 -13110
rect 31836 -13174 31842 -13170
rect 30616 -13310 30622 -13250
rect 30682 -13310 30688 -13250
rect 34286 -13390 34346 -12954
rect 34742 -12954 34756 -12918
rect 34790 -12814 34806 -12778
rect 35162 -12110 35222 -11730
rect 35396 -12020 35456 -11730
rect 35318 -12026 35526 -12020
rect 35318 -12060 35330 -12026
rect 35514 -12060 35526 -12026
rect 35318 -12066 35526 -12060
rect 35162 -12286 35176 -12110
rect 35210 -12286 35222 -12110
rect 35622 -12110 35682 -11730
rect 35856 -11894 35916 -11888
rect 35916 -11954 39120 -11894
rect 35856 -12020 35916 -11954
rect 36312 -12020 36372 -11954
rect 36778 -12020 36838 -11954
rect 37228 -12020 37288 -11954
rect 37682 -12020 37742 -11954
rect 38144 -12020 38204 -11954
rect 38598 -12020 38658 -11954
rect 39060 -12020 39120 -11954
rect 39510 -12020 39570 -11730
rect 35776 -12026 35984 -12020
rect 35776 -12060 35788 -12026
rect 35972 -12060 35984 -12026
rect 35776 -12066 35984 -12060
rect 36234 -12026 36442 -12020
rect 36234 -12060 36246 -12026
rect 36430 -12060 36442 -12026
rect 36234 -12066 36442 -12060
rect 36692 -12026 36900 -12020
rect 36692 -12060 36704 -12026
rect 36888 -12060 36900 -12026
rect 36692 -12066 36900 -12060
rect 37150 -12026 37358 -12020
rect 37150 -12060 37162 -12026
rect 37346 -12060 37358 -12026
rect 37150 -12066 37358 -12060
rect 37608 -12026 37816 -12020
rect 37608 -12060 37620 -12026
rect 37804 -12060 37816 -12026
rect 37608 -12066 37816 -12060
rect 38066 -12026 38274 -12020
rect 38066 -12060 38078 -12026
rect 38262 -12060 38274 -12026
rect 38066 -12066 38274 -12060
rect 38524 -12026 38732 -12020
rect 38524 -12060 38536 -12026
rect 38720 -12060 38732 -12026
rect 38524 -12066 38732 -12060
rect 38982 -12026 39190 -12020
rect 38982 -12060 38994 -12026
rect 39178 -12060 39190 -12026
rect 38982 -12066 39190 -12060
rect 39440 -12026 39648 -12020
rect 39440 -12060 39452 -12026
rect 39636 -12060 39648 -12026
rect 39440 -12066 39648 -12060
rect 35622 -12138 35634 -12110
rect 35162 -12778 35222 -12286
rect 35628 -12286 35634 -12138
rect 35668 -12138 35682 -12110
rect 36086 -12110 36132 -12098
rect 35668 -12286 35674 -12138
rect 35628 -12298 35674 -12286
rect 36086 -12286 36092 -12110
rect 36126 -12286 36132 -12110
rect 36086 -12298 36132 -12286
rect 36544 -12110 36590 -12098
rect 36544 -12286 36550 -12110
rect 36584 -12286 36590 -12110
rect 36544 -12298 36590 -12286
rect 37002 -12110 37048 -12098
rect 37002 -12286 37008 -12110
rect 37042 -12286 37048 -12110
rect 37002 -12298 37048 -12286
rect 37460 -12110 37506 -12098
rect 37460 -12286 37466 -12110
rect 37500 -12286 37506 -12110
rect 37460 -12298 37506 -12286
rect 37918 -12110 37964 -12098
rect 37918 -12286 37924 -12110
rect 37958 -12286 37964 -12110
rect 37918 -12298 37964 -12286
rect 38376 -12110 38422 -12098
rect 38376 -12286 38382 -12110
rect 38416 -12286 38422 -12110
rect 38376 -12298 38422 -12286
rect 38834 -12110 38880 -12098
rect 38834 -12286 38840 -12110
rect 38874 -12286 38880 -12110
rect 39292 -12110 39338 -12098
rect 39292 -12258 39298 -12110
rect 38834 -12298 38880 -12286
rect 39286 -12286 39298 -12258
rect 39332 -12258 39338 -12110
rect 39750 -12110 39810 -11730
rect 39332 -12286 39346 -12258
rect 39750 -12266 39756 -12110
rect 35318 -12336 35526 -12330
rect 35318 -12370 35330 -12336
rect 35514 -12370 35526 -12336
rect 35318 -12376 35526 -12370
rect 35776 -12336 35984 -12330
rect 35776 -12370 35788 -12336
rect 35972 -12370 35984 -12336
rect 35776 -12376 35984 -12370
rect 36234 -12336 36442 -12330
rect 36234 -12370 36246 -12336
rect 36430 -12370 36442 -12336
rect 36234 -12376 36442 -12370
rect 36692 -12336 36900 -12330
rect 36692 -12370 36704 -12336
rect 36888 -12370 36900 -12336
rect 36692 -12376 36900 -12370
rect 37150 -12336 37358 -12330
rect 37150 -12370 37162 -12336
rect 37346 -12370 37358 -12336
rect 37150 -12376 37358 -12370
rect 37608 -12336 37816 -12330
rect 37608 -12370 37620 -12336
rect 37804 -12370 37816 -12336
rect 37608 -12376 37816 -12370
rect 38066 -12336 38274 -12330
rect 38066 -12370 38078 -12336
rect 38262 -12370 38274 -12336
rect 38066 -12376 38274 -12370
rect 38524 -12336 38732 -12330
rect 38524 -12370 38536 -12336
rect 38720 -12370 38732 -12336
rect 38524 -12376 38732 -12370
rect 38982 -12336 39190 -12330
rect 38982 -12370 38994 -12336
rect 39178 -12370 39190 -12336
rect 38982 -12376 39190 -12370
rect 35394 -12688 35454 -12376
rect 35850 -12442 35910 -12376
rect 36306 -12442 36366 -12376
rect 36772 -12442 36832 -12376
rect 37222 -12442 37282 -12376
rect 37676 -12442 37736 -12376
rect 38138 -12442 38198 -12376
rect 38592 -12442 38652 -12376
rect 39054 -12442 39114 -12376
rect 35850 -12502 39114 -12442
rect 35856 -12622 39120 -12562
rect 35856 -12688 35916 -12622
rect 36312 -12688 36372 -12622
rect 36778 -12688 36838 -12622
rect 37228 -12688 37288 -12622
rect 37682 -12688 37742 -12622
rect 38144 -12688 38204 -12622
rect 38598 -12688 38658 -12622
rect 39060 -12688 39120 -12622
rect 35318 -12694 35526 -12688
rect 35318 -12728 35330 -12694
rect 35514 -12728 35526 -12694
rect 35318 -12734 35526 -12728
rect 35776 -12694 35984 -12688
rect 35776 -12728 35788 -12694
rect 35972 -12728 35984 -12694
rect 35776 -12734 35984 -12728
rect 36234 -12694 36442 -12688
rect 36234 -12728 36246 -12694
rect 36430 -12728 36442 -12694
rect 36234 -12734 36442 -12728
rect 36692 -12694 36900 -12688
rect 36692 -12728 36704 -12694
rect 36888 -12728 36900 -12694
rect 36692 -12734 36900 -12728
rect 37150 -12694 37358 -12688
rect 37150 -12728 37162 -12694
rect 37346 -12728 37358 -12694
rect 37150 -12734 37358 -12728
rect 37608 -12694 37816 -12688
rect 37608 -12728 37620 -12694
rect 37804 -12728 37816 -12694
rect 37608 -12734 37816 -12728
rect 38066 -12694 38274 -12688
rect 38066 -12728 38078 -12694
rect 38262 -12728 38274 -12694
rect 38066 -12734 38274 -12728
rect 38524 -12694 38732 -12688
rect 38524 -12728 38536 -12694
rect 38720 -12728 38732 -12694
rect 38524 -12734 38732 -12728
rect 38982 -12694 39190 -12688
rect 38982 -12728 38994 -12694
rect 39178 -12728 39190 -12694
rect 38982 -12734 39190 -12728
rect 34790 -12918 34796 -12814
rect 35162 -12834 35176 -12778
rect 34790 -12954 34802 -12918
rect 35170 -12926 35176 -12834
rect 34440 -13004 34648 -12998
rect 34440 -13038 34452 -13004
rect 34636 -13038 34648 -13004
rect 34440 -13044 34648 -13038
rect 34508 -13390 34568 -13044
rect 34742 -13390 34802 -12954
rect 35162 -12954 35176 -12926
rect 35210 -12834 35222 -12778
rect 35628 -12778 35674 -12766
rect 35210 -12926 35216 -12834
rect 35628 -12924 35634 -12778
rect 35210 -12954 35222 -12926
rect 35162 -13390 35222 -12954
rect 35622 -12954 35634 -12924
rect 35668 -12924 35674 -12778
rect 36086 -12778 36132 -12766
rect 35668 -12954 35682 -12924
rect 35318 -13004 35526 -12998
rect 35318 -13038 35330 -13004
rect 35514 -13038 35526 -13004
rect 35318 -13044 35526 -13038
rect 35394 -13390 35454 -13044
rect 35622 -13238 35682 -12954
rect 36086 -12954 36092 -12778
rect 36126 -12954 36132 -12778
rect 36086 -12966 36132 -12954
rect 36544 -12778 36590 -12766
rect 36544 -12954 36550 -12778
rect 36584 -12954 36590 -12778
rect 36544 -12966 36590 -12954
rect 37002 -12778 37048 -12766
rect 37002 -12954 37008 -12778
rect 37042 -12954 37048 -12778
rect 37002 -12966 37048 -12954
rect 37460 -12778 37506 -12766
rect 37460 -12954 37466 -12778
rect 37500 -12954 37506 -12778
rect 37460 -12966 37506 -12954
rect 37918 -12778 37964 -12766
rect 37918 -12954 37924 -12778
rect 37958 -12954 37964 -12778
rect 37918 -12966 37964 -12954
rect 38376 -12778 38422 -12766
rect 38376 -12954 38382 -12778
rect 38416 -12954 38422 -12778
rect 38376 -12966 38422 -12954
rect 38834 -12778 38880 -12766
rect 38834 -12954 38840 -12778
rect 38874 -12954 38880 -12778
rect 39286 -12778 39346 -12286
rect 39742 -12286 39756 -12266
rect 39790 -12140 39810 -12110
rect 39790 -12266 39796 -12140
rect 39790 -12286 39802 -12266
rect 39440 -12336 39648 -12330
rect 39440 -12370 39452 -12336
rect 39636 -12370 39648 -12336
rect 39440 -12376 39648 -12370
rect 39514 -12502 39574 -12376
rect 39742 -12502 39802 -12286
rect 39514 -12562 39802 -12502
rect 39514 -12688 39574 -12562
rect 39440 -12694 39648 -12688
rect 39440 -12728 39452 -12694
rect 39636 -12728 39648 -12694
rect 39440 -12734 39648 -12728
rect 39286 -12820 39298 -12778
rect 38834 -12966 38880 -12954
rect 39292 -12954 39298 -12820
rect 39332 -12820 39346 -12778
rect 39742 -12778 39802 -12562
rect 39742 -12818 39756 -12778
rect 39332 -12954 39338 -12820
rect 39750 -12914 39756 -12818
rect 39292 -12966 39338 -12954
rect 39742 -12954 39756 -12914
rect 39790 -12818 39802 -12778
rect 39790 -12914 39796 -12818
rect 39790 -12954 39802 -12914
rect 35776 -13004 35984 -12998
rect 35776 -13038 35788 -13004
rect 35972 -13038 35984 -13004
rect 35776 -13044 35984 -13038
rect 36234 -13004 36442 -12998
rect 36234 -13038 36246 -13004
rect 36430 -13038 36442 -13004
rect 36234 -13044 36442 -13038
rect 36692 -13004 36900 -12998
rect 36692 -13038 36704 -13004
rect 36888 -13038 36900 -13004
rect 36692 -13044 36900 -13038
rect 37150 -13004 37358 -12998
rect 37150 -13038 37162 -13004
rect 37346 -13038 37358 -13004
rect 37150 -13044 37358 -13038
rect 37608 -13004 37816 -12998
rect 37608 -13038 37620 -13004
rect 37804 -13038 37816 -13004
rect 37608 -13044 37816 -13038
rect 38066 -13004 38274 -12998
rect 38066 -13038 38078 -13004
rect 38262 -13038 38274 -13004
rect 38066 -13044 38274 -13038
rect 38524 -13004 38732 -12998
rect 38524 -13038 38536 -13004
rect 38720 -13038 38732 -13004
rect 38524 -13044 38732 -13038
rect 38982 -13004 39190 -12998
rect 38982 -13038 38994 -13004
rect 39178 -13038 39190 -13004
rect 38982 -13044 39190 -13038
rect 39440 -13004 39648 -12998
rect 39440 -13038 39452 -13004
rect 39636 -13038 39648 -13004
rect 39440 -13044 39648 -13038
rect 35850 -13110 35916 -13044
rect 36306 -13104 36372 -13044
rect 36306 -13110 36312 -13104
rect 35850 -13170 35856 -13110
rect 35916 -13164 36312 -13110
rect 36372 -13110 36378 -13104
rect 36772 -13110 36838 -13044
rect 37222 -13110 37288 -13044
rect 37676 -13110 37742 -13044
rect 38138 -13104 38204 -13044
rect 38138 -13110 38144 -13104
rect 36372 -13164 36778 -13110
rect 35916 -13170 36778 -13164
rect 36838 -13170 37228 -13110
rect 37288 -13170 37682 -13110
rect 37742 -13164 38144 -13110
rect 38204 -13110 38210 -13104
rect 38592 -13110 38658 -13044
rect 39054 -13104 39120 -13044
rect 39054 -13110 39060 -13104
rect 38204 -13164 38598 -13110
rect 37742 -13170 38598 -13164
rect 38658 -13164 39060 -13110
rect 39120 -13164 39126 -13104
rect 38658 -13170 39114 -13164
rect 35622 -13304 35682 -13298
rect 39512 -13390 39572 -13044
rect 39742 -13390 39802 -12954
rect 40110 -13266 40116 -11262
rect 40216 -13266 40222 -11262
rect 40110 -13390 40222 -13266
rect 29766 -13396 40222 -13390
rect 29766 -13496 29872 -13396
rect 40116 -13496 40222 -13396
rect 29766 -13502 40222 -13496
rect 29766 -13732 40222 -13726
rect 29766 -13832 29872 -13732
rect 40116 -13832 40222 -13732
rect 29766 -13838 40222 -13832
rect 29766 -14014 29878 -13838
rect 29766 -19186 29772 -14014
rect 29872 -15808 29878 -14014
rect 30164 -14271 30224 -13838
rect 30392 -14172 30452 -13838
rect 30622 -13912 30682 -13906
rect 30317 -14178 30525 -14172
rect 30317 -14212 30329 -14178
rect 30513 -14212 30525 -14178
rect 30317 -14218 30525 -14212
rect 30164 -14304 30175 -14271
rect 30169 -15394 30175 -14304
rect 30166 -15447 30175 -15394
rect 30209 -14304 30224 -14271
rect 30622 -14271 30682 -13972
rect 30854 -14042 30914 -14036
rect 31310 -14042 31370 -14036
rect 32226 -14042 32286 -14036
rect 30914 -14102 31310 -14044
rect 31776 -14044 31836 -14042
rect 31370 -14048 32226 -14044
rect 31370 -14102 31776 -14048
rect 30854 -14104 31776 -14102
rect 30854 -14172 30914 -14104
rect 31310 -14172 31370 -14104
rect 31836 -14102 32226 -14048
rect 32680 -14042 32740 -14036
rect 32286 -14102 32680 -14044
rect 33142 -14042 33202 -14036
rect 34058 -14040 34118 -14034
rect 32740 -14102 33142 -14044
rect 33596 -14044 33656 -14042
rect 33202 -14048 34058 -14044
rect 33202 -14102 33596 -14048
rect 31836 -14104 33596 -14102
rect 31776 -14172 31836 -14108
rect 32226 -14172 32286 -14104
rect 32680 -14172 32740 -14104
rect 33142 -14172 33202 -14104
rect 33656 -14100 34058 -14048
rect 33656 -14104 34118 -14100
rect 33596 -14172 33656 -14108
rect 34058 -14172 34118 -14104
rect 30775 -14178 30983 -14172
rect 30775 -14212 30787 -14178
rect 30971 -14212 30983 -14178
rect 30775 -14218 30983 -14212
rect 31233 -14178 31441 -14172
rect 31233 -14212 31245 -14178
rect 31429 -14212 31441 -14178
rect 31233 -14218 31441 -14212
rect 31691 -14178 31899 -14172
rect 31691 -14212 31703 -14178
rect 31887 -14212 31899 -14178
rect 31691 -14218 31899 -14212
rect 32149 -14178 32357 -14172
rect 32149 -14212 32161 -14178
rect 32345 -14212 32357 -14178
rect 32149 -14218 32357 -14212
rect 32607 -14178 32815 -14172
rect 32607 -14212 32619 -14178
rect 32803 -14212 32815 -14178
rect 32607 -14218 32815 -14212
rect 33065 -14178 33273 -14172
rect 33065 -14212 33077 -14178
rect 33261 -14212 33273 -14178
rect 33065 -14218 33273 -14212
rect 33523 -14178 33731 -14172
rect 33523 -14212 33535 -14178
rect 33719 -14212 33731 -14178
rect 33523 -14218 33731 -14212
rect 33981 -14178 34189 -14172
rect 33981 -14212 33993 -14178
rect 34177 -14212 34189 -14178
rect 33981 -14218 34189 -14212
rect 30622 -14278 30633 -14271
rect 30209 -15394 30215 -14304
rect 30209 -15447 30226 -15394
rect 30166 -15808 30226 -15447
rect 30627 -15447 30633 -14278
rect 30667 -14278 30682 -14271
rect 31085 -14271 31131 -14259
rect 30667 -15447 30673 -14278
rect 30627 -15459 30673 -15447
rect 31085 -15447 31091 -14271
rect 31125 -15447 31131 -14271
rect 31085 -15459 31131 -15447
rect 31543 -14271 31589 -14259
rect 31543 -15447 31549 -14271
rect 31583 -15447 31589 -14271
rect 31543 -15459 31589 -15447
rect 32001 -14271 32047 -14259
rect 32001 -15447 32007 -14271
rect 32041 -15447 32047 -14271
rect 32001 -15459 32047 -15447
rect 32459 -14271 32505 -14259
rect 32459 -15447 32465 -14271
rect 32499 -15447 32505 -14271
rect 32459 -15459 32505 -15447
rect 32917 -14271 32963 -14259
rect 32917 -15447 32923 -14271
rect 32957 -15447 32963 -14271
rect 32917 -15459 32963 -15447
rect 33375 -14271 33421 -14259
rect 33375 -15447 33381 -14271
rect 33415 -15447 33421 -14271
rect 33375 -15459 33421 -15447
rect 33833 -14271 33879 -14259
rect 33833 -15447 33839 -14271
rect 33873 -15447 33879 -14271
rect 34286 -14271 34346 -13838
rect 34516 -14172 34576 -13838
rect 34439 -14178 34647 -14172
rect 34439 -14212 34451 -14178
rect 34635 -14212 34647 -14178
rect 34439 -14218 34647 -14212
rect 34286 -14312 34297 -14271
rect 34291 -15404 34297 -14312
rect 33833 -15459 33879 -15447
rect 34284 -15447 34297 -15404
rect 34331 -14312 34346 -14271
rect 34744 -14271 34804 -13838
rect 34744 -14306 34755 -14271
rect 34331 -15404 34337 -14312
rect 34331 -15447 34344 -15404
rect 34749 -15426 34755 -14306
rect 30317 -15506 30525 -15500
rect 30317 -15540 30329 -15506
rect 30513 -15540 30525 -15506
rect 30317 -15546 30525 -15540
rect 30775 -15506 30983 -15500
rect 30775 -15540 30787 -15506
rect 30971 -15540 30983 -15506
rect 30775 -15546 30983 -15540
rect 31233 -15506 31441 -15500
rect 31233 -15540 31245 -15506
rect 31429 -15540 31441 -15506
rect 31233 -15546 31441 -15540
rect 31691 -15506 31899 -15500
rect 31691 -15540 31703 -15506
rect 31887 -15540 31899 -15506
rect 31691 -15546 31899 -15540
rect 32149 -15506 32357 -15500
rect 32149 -15540 32161 -15506
rect 32345 -15540 32357 -15506
rect 32149 -15546 32357 -15540
rect 32607 -15506 32815 -15500
rect 32607 -15540 32619 -15506
rect 32803 -15540 32815 -15506
rect 32607 -15546 32815 -15540
rect 33065 -15506 33273 -15500
rect 33065 -15540 33077 -15506
rect 33261 -15540 33273 -15506
rect 33065 -15546 33273 -15540
rect 33523 -15506 33731 -15500
rect 33523 -15540 33535 -15506
rect 33719 -15540 33731 -15506
rect 33523 -15546 33731 -15540
rect 33981 -15506 34189 -15500
rect 33981 -15540 33993 -15506
rect 34177 -15540 34189 -15506
rect 33981 -15546 34189 -15540
rect 30392 -15808 30452 -15546
rect 30854 -15616 30914 -15546
rect 31310 -15616 31370 -15546
rect 31776 -15616 31836 -15546
rect 32226 -15616 32286 -15546
rect 32680 -15616 32740 -15546
rect 33142 -15616 33202 -15546
rect 33596 -15616 33656 -15546
rect 34058 -15616 34118 -15546
rect 30854 -15676 34118 -15616
rect 34284 -15598 34344 -15447
rect 34742 -15447 34755 -15426
rect 34789 -14306 34804 -14271
rect 35164 -14271 35224 -13838
rect 35392 -14172 35452 -13838
rect 35616 -13978 35622 -13918
rect 35682 -13978 35688 -13918
rect 35317 -14178 35525 -14172
rect 35317 -14212 35329 -14178
rect 35513 -14212 35525 -14178
rect 35317 -14218 35525 -14212
rect 35164 -14306 35175 -14271
rect 34789 -15426 34795 -14306
rect 34789 -15447 34802 -15426
rect 35169 -15432 35175 -14306
rect 34439 -15506 34647 -15500
rect 34439 -15540 34451 -15506
rect 34635 -15540 34647 -15506
rect 34439 -15546 34647 -15540
rect 34510 -15598 34570 -15546
rect 34742 -15598 34802 -15447
rect 35162 -15447 35175 -15432
rect 35209 -14306 35224 -14271
rect 35622 -14271 35682 -13978
rect 35856 -14040 35916 -14034
rect 37228 -14038 37288 -14032
rect 36312 -14044 36372 -14038
rect 36778 -14044 36838 -14038
rect 35916 -14100 36312 -14044
rect 35856 -14104 36312 -14100
rect 36372 -14104 36778 -14044
rect 36838 -14098 37228 -14044
rect 37682 -14044 37742 -14038
rect 38144 -14044 38204 -14038
rect 38598 -14040 38658 -14034
rect 37288 -14098 37682 -14044
rect 36838 -14104 37682 -14098
rect 37742 -14104 38144 -14044
rect 38204 -14100 38598 -14044
rect 39060 -14040 39120 -14034
rect 38658 -14100 39060 -14044
rect 38204 -14104 39120 -14100
rect 35856 -14172 35916 -14104
rect 36312 -14172 36372 -14104
rect 36778 -14172 36838 -14104
rect 37228 -14172 37288 -14104
rect 37682 -14172 37742 -14104
rect 38144 -14172 38204 -14104
rect 38598 -14172 38658 -14104
rect 39060 -14172 39120 -14104
rect 39514 -14172 39574 -13838
rect 35775 -14178 35983 -14172
rect 35775 -14212 35787 -14178
rect 35971 -14212 35983 -14178
rect 35775 -14218 35983 -14212
rect 36233 -14178 36441 -14172
rect 36233 -14212 36245 -14178
rect 36429 -14212 36441 -14178
rect 36233 -14218 36441 -14212
rect 36691 -14178 36899 -14172
rect 36691 -14212 36703 -14178
rect 36887 -14212 36899 -14178
rect 36691 -14218 36899 -14212
rect 37149 -14178 37357 -14172
rect 37149 -14212 37161 -14178
rect 37345 -14212 37357 -14178
rect 37149 -14218 37357 -14212
rect 37607 -14178 37815 -14172
rect 37607 -14212 37619 -14178
rect 37803 -14212 37815 -14178
rect 37607 -14218 37815 -14212
rect 38065 -14178 38273 -14172
rect 38065 -14212 38077 -14178
rect 38261 -14212 38273 -14178
rect 38065 -14218 38273 -14212
rect 38523 -14178 38731 -14172
rect 38523 -14212 38535 -14178
rect 38719 -14212 38731 -14178
rect 38523 -14218 38731 -14212
rect 38981 -14178 39189 -14172
rect 38981 -14212 38993 -14178
rect 39177 -14212 39189 -14178
rect 38981 -14218 39189 -14212
rect 39439 -14178 39647 -14172
rect 39439 -14212 39451 -14178
rect 39635 -14212 39647 -14178
rect 39439 -14218 39647 -14212
rect 35209 -15432 35215 -14306
rect 35622 -14338 35633 -14271
rect 35209 -15447 35222 -15432
rect 35162 -15598 35222 -15447
rect 35627 -15447 35633 -14338
rect 35667 -14338 35682 -14271
rect 36085 -14271 36131 -14259
rect 35667 -15447 35673 -14338
rect 35627 -15459 35673 -15447
rect 36085 -15447 36091 -14271
rect 36125 -15447 36131 -14271
rect 36085 -15459 36131 -15447
rect 36543 -14271 36589 -14259
rect 36543 -15447 36549 -14271
rect 36583 -15447 36589 -14271
rect 36543 -15459 36589 -15447
rect 37001 -14271 37047 -14259
rect 37001 -15447 37007 -14271
rect 37041 -15447 37047 -14271
rect 37001 -15459 37047 -15447
rect 37459 -14271 37505 -14259
rect 37459 -15447 37465 -14271
rect 37499 -15447 37505 -14271
rect 37459 -15459 37505 -15447
rect 37917 -14271 37963 -14259
rect 37917 -15447 37923 -14271
rect 37957 -15447 37963 -14271
rect 37917 -15459 37963 -15447
rect 38375 -14271 38421 -14259
rect 38375 -15447 38381 -14271
rect 38415 -15447 38421 -14271
rect 38375 -15459 38421 -15447
rect 38833 -14271 38879 -14259
rect 38833 -15447 38839 -14271
rect 38873 -15447 38879 -14271
rect 39291 -14271 39337 -14259
rect 39291 -15380 39297 -14271
rect 38833 -15459 38879 -15447
rect 39284 -15447 39297 -15380
rect 39331 -15380 39337 -14271
rect 39742 -14271 39802 -13838
rect 39742 -14292 39755 -14271
rect 39331 -15447 39344 -15380
rect 39749 -15400 39755 -14292
rect 35317 -15506 35525 -15500
rect 35317 -15540 35329 -15506
rect 35513 -15540 35525 -15506
rect 35317 -15546 35525 -15540
rect 35775 -15506 35983 -15500
rect 35775 -15540 35787 -15506
rect 35971 -15540 35983 -15506
rect 35775 -15546 35983 -15540
rect 36233 -15506 36441 -15500
rect 36233 -15540 36245 -15506
rect 36429 -15540 36441 -15506
rect 36233 -15546 36441 -15540
rect 36691 -15506 36899 -15500
rect 36691 -15540 36703 -15506
rect 36887 -15540 36899 -15506
rect 36691 -15546 36899 -15540
rect 37149 -15506 37357 -15500
rect 37149 -15540 37161 -15506
rect 37345 -15540 37357 -15506
rect 37149 -15546 37357 -15540
rect 37607 -15506 37815 -15500
rect 37607 -15540 37619 -15506
rect 37803 -15540 37815 -15506
rect 37607 -15546 37815 -15540
rect 38065 -15506 38273 -15500
rect 38065 -15540 38077 -15506
rect 38261 -15540 38273 -15506
rect 38065 -15546 38273 -15540
rect 38523 -15506 38731 -15500
rect 38523 -15540 38535 -15506
rect 38719 -15540 38731 -15506
rect 38523 -15546 38731 -15540
rect 38981 -15506 39189 -15500
rect 38981 -15540 38993 -15506
rect 39177 -15540 39189 -15506
rect 38981 -15546 39189 -15540
rect 35392 -15598 35452 -15546
rect 34284 -15658 35452 -15598
rect 35848 -15616 35908 -15546
rect 36304 -15616 36364 -15546
rect 36770 -15616 36830 -15546
rect 37220 -15616 37280 -15546
rect 37674 -15616 37734 -15546
rect 38136 -15616 38196 -15546
rect 38590 -15616 38650 -15546
rect 39052 -15616 39112 -15546
rect 35848 -15676 39112 -15616
rect 39284 -15718 39344 -15447
rect 39742 -15447 39755 -15400
rect 39789 -14292 39802 -14271
rect 40110 -14014 40222 -13838
rect 39789 -15400 39795 -14292
rect 39789 -15447 39802 -15400
rect 39439 -15506 39647 -15500
rect 39439 -15540 39451 -15506
rect 39635 -15540 39647 -15506
rect 39439 -15546 39647 -15540
rect 39278 -15778 39284 -15718
rect 39344 -15778 39350 -15718
rect 29872 -15868 31002 -15808
rect 29872 -16302 29878 -15868
rect 30942 -16302 31002 -15868
rect 31854 -15884 38330 -15824
rect 39514 -15872 39574 -15546
rect 39742 -15872 39802 -15447
rect 40110 -15872 40116 -14014
rect 29872 -16362 31460 -16302
rect 29872 -19186 29878 -16362
rect 30942 -16536 31002 -16362
rect 31168 -16437 31228 -16362
rect 31094 -16443 31302 -16437
rect 31094 -16477 31106 -16443
rect 31290 -16477 31302 -16443
rect 31094 -16483 31302 -16477
rect 30942 -16580 30952 -16536
rect 30946 -18042 30952 -16580
rect 30938 -18112 30952 -18042
rect 30986 -16580 31002 -16536
rect 31400 -16536 31460 -16362
rect 31624 -16364 31630 -16304
rect 31690 -16364 31696 -16304
rect 31630 -16437 31690 -16364
rect 31552 -16443 31760 -16437
rect 31552 -16477 31564 -16443
rect 31748 -16477 31760 -16443
rect 31552 -16483 31760 -16477
rect 30986 -18042 30992 -16580
rect 31400 -16598 31410 -16536
rect 31404 -18036 31410 -16598
rect 30986 -18112 30998 -18042
rect 30938 -18900 30998 -18112
rect 31396 -18112 31410 -18036
rect 31444 -16598 31460 -16536
rect 31854 -16536 31914 -15884
rect 32768 -16014 37412 -15954
rect 32084 -16364 32090 -16304
rect 32150 -16364 32156 -16304
rect 32542 -16364 32548 -16304
rect 32608 -16364 32614 -16304
rect 32090 -16437 32150 -16364
rect 32548 -16437 32608 -16364
rect 32010 -16443 32218 -16437
rect 32010 -16477 32022 -16443
rect 32206 -16477 32218 -16443
rect 32010 -16483 32218 -16477
rect 32468 -16443 32676 -16437
rect 32468 -16477 32480 -16443
rect 32664 -16477 32676 -16443
rect 32468 -16483 32676 -16477
rect 31854 -16596 31868 -16536
rect 31444 -18036 31450 -16598
rect 31444 -18112 31456 -18036
rect 31094 -18171 31302 -18165
rect 31094 -18205 31106 -18171
rect 31290 -18205 31302 -18171
rect 31094 -18211 31302 -18205
rect 31166 -18900 31226 -18211
rect 31396 -18900 31456 -18112
rect 31862 -18112 31868 -16596
rect 31902 -16596 31914 -16536
rect 32320 -16536 32366 -16524
rect 31902 -18112 31908 -16596
rect 32320 -18056 32326 -16536
rect 31862 -18124 31908 -18112
rect 32312 -18112 32326 -18056
rect 32360 -18056 32366 -16536
rect 32768 -16536 32828 -16014
rect 33688 -16140 36504 -16080
rect 32998 -16364 33004 -16304
rect 33064 -16364 33070 -16304
rect 33454 -16364 33460 -16304
rect 33520 -16364 33526 -16304
rect 33004 -16437 33064 -16364
rect 33460 -16437 33520 -16364
rect 32926 -16443 33134 -16437
rect 32926 -16477 32938 -16443
rect 33122 -16477 33134 -16443
rect 32926 -16483 33134 -16477
rect 33384 -16443 33592 -16437
rect 33384 -16477 33396 -16443
rect 33580 -16477 33592 -16443
rect 33384 -16483 33592 -16477
rect 32768 -16604 32784 -16536
rect 32360 -18112 32372 -18056
rect 31552 -18171 31760 -18165
rect 31552 -18205 31564 -18171
rect 31748 -18205 31760 -18171
rect 31552 -18211 31760 -18205
rect 32010 -18171 32218 -18165
rect 32010 -18205 32022 -18171
rect 32206 -18205 32218 -18171
rect 32010 -18211 32218 -18205
rect 31626 -18278 31686 -18211
rect 32086 -18278 32146 -18211
rect 31620 -18338 31626 -18278
rect 31686 -18338 31692 -18278
rect 32080 -18338 32086 -18278
rect 32146 -18338 32152 -18278
rect 32312 -18646 32372 -18112
rect 32778 -18112 32784 -16604
rect 32818 -16604 32828 -16536
rect 33236 -16536 33282 -16524
rect 32818 -18112 32824 -16604
rect 33236 -18054 33242 -16536
rect 32778 -18124 32824 -18112
rect 33232 -18112 33242 -18054
rect 33276 -18054 33282 -16536
rect 33688 -16536 33748 -16140
rect 34602 -16256 35580 -16196
rect 33910 -16364 33916 -16304
rect 33976 -16364 33982 -16304
rect 34370 -16364 34376 -16304
rect 34436 -16364 34442 -16304
rect 33916 -16437 33976 -16364
rect 34376 -16437 34436 -16364
rect 33842 -16443 34050 -16437
rect 33842 -16477 33854 -16443
rect 34038 -16477 34050 -16443
rect 33842 -16483 34050 -16477
rect 34300 -16443 34508 -16437
rect 34300 -16477 34312 -16443
rect 34496 -16477 34508 -16443
rect 34300 -16483 34508 -16477
rect 33688 -16568 33700 -16536
rect 33276 -18112 33292 -18054
rect 32468 -18171 32676 -18165
rect 32468 -18205 32480 -18171
rect 32664 -18205 32676 -18171
rect 32468 -18211 32676 -18205
rect 32926 -18171 33134 -18165
rect 32926 -18205 32938 -18171
rect 33122 -18205 33134 -18171
rect 32926 -18211 33134 -18205
rect 32544 -18278 32604 -18211
rect 33000 -18278 33060 -18211
rect 32538 -18338 32544 -18278
rect 32604 -18338 32610 -18278
rect 32994 -18338 33000 -18278
rect 33060 -18338 33066 -18278
rect 33232 -18512 33292 -18112
rect 33694 -18112 33700 -16568
rect 33734 -16568 33748 -16536
rect 34152 -16536 34198 -16524
rect 33734 -18112 33740 -16568
rect 34152 -18068 34158 -16536
rect 33694 -18124 33740 -18112
rect 34148 -18112 34158 -18068
rect 34192 -18068 34198 -16536
rect 34602 -16536 34662 -16256
rect 34820 -16304 34904 -16300
rect 34820 -16366 34832 -16304
rect 34892 -16366 34904 -16304
rect 34820 -16372 34904 -16366
rect 35058 -16316 35118 -16310
rect 34832 -16437 34892 -16372
rect 35286 -16364 35292 -16304
rect 35352 -16364 35358 -16304
rect 35286 -16366 35358 -16364
rect 34758 -16443 34966 -16437
rect 34758 -16477 34770 -16443
rect 34954 -16477 34966 -16443
rect 34758 -16483 34966 -16477
rect 34602 -16564 34616 -16536
rect 34192 -18112 34208 -18068
rect 33384 -18171 33592 -18165
rect 33384 -18205 33396 -18171
rect 33580 -18205 33592 -18171
rect 33384 -18211 33592 -18205
rect 33842 -18171 34050 -18165
rect 33842 -18205 33854 -18171
rect 34038 -18205 34050 -18171
rect 33842 -18211 34050 -18205
rect 33456 -18278 33516 -18211
rect 33912 -18278 33972 -18211
rect 33450 -18338 33456 -18278
rect 33516 -18338 33522 -18278
rect 33906 -18338 33912 -18278
rect 33972 -18338 33978 -18278
rect 34148 -18388 34208 -18112
rect 34610 -18112 34616 -16564
rect 34650 -16564 34662 -16536
rect 35058 -16536 35118 -16376
rect 35292 -16437 35352 -16366
rect 35216 -16443 35424 -16437
rect 35216 -16477 35228 -16443
rect 35412 -16477 35424 -16443
rect 35216 -16483 35424 -16477
rect 35058 -16558 35074 -16536
rect 34650 -18112 34656 -16564
rect 34610 -18124 34656 -18112
rect 35068 -18112 35074 -16558
rect 35108 -16558 35118 -16536
rect 35520 -16536 35580 -16256
rect 35744 -16364 35750 -16304
rect 35810 -16364 35816 -16304
rect 36198 -16364 36204 -16304
rect 36264 -16364 36270 -16304
rect 35750 -16437 35810 -16364
rect 36204 -16437 36264 -16364
rect 35674 -16443 35882 -16437
rect 35674 -16477 35686 -16443
rect 35870 -16477 35882 -16443
rect 35674 -16483 35882 -16477
rect 36132 -16443 36340 -16437
rect 36132 -16477 36144 -16443
rect 36328 -16477 36340 -16443
rect 36132 -16483 36340 -16477
rect 36444 -16524 36504 -16140
rect 36662 -16364 36668 -16304
rect 36728 -16364 36734 -16304
rect 37120 -16364 37126 -16304
rect 37186 -16364 37192 -16304
rect 36668 -16437 36728 -16364
rect 37126 -16437 37186 -16364
rect 36590 -16443 36798 -16437
rect 36590 -16477 36602 -16443
rect 36786 -16477 36798 -16443
rect 36590 -16483 36798 -16477
rect 37048 -16443 37256 -16437
rect 37048 -16477 37060 -16443
rect 37244 -16477 37256 -16443
rect 37048 -16483 37256 -16477
rect 35108 -18112 35114 -16558
rect 35520 -16616 35532 -16536
rect 35068 -18124 35114 -18112
rect 35526 -18112 35532 -16616
rect 35566 -16616 35580 -16536
rect 35984 -16536 36030 -16524
rect 35566 -18112 35572 -16616
rect 35984 -18034 35990 -16536
rect 35526 -18124 35572 -18112
rect 35978 -18112 35990 -18034
rect 36024 -18034 36030 -16536
rect 36442 -16536 36504 -16524
rect 36024 -18112 36038 -18034
rect 34300 -18171 34508 -18165
rect 34300 -18205 34312 -18171
rect 34496 -18205 34508 -18171
rect 34300 -18211 34508 -18205
rect 34758 -18171 34966 -18165
rect 34758 -18205 34770 -18171
rect 34954 -18205 34966 -18171
rect 34758 -18211 34966 -18205
rect 35216 -18171 35424 -18165
rect 35216 -18205 35228 -18171
rect 35412 -18205 35424 -18171
rect 35216 -18211 35424 -18205
rect 35674 -18171 35882 -18165
rect 35674 -18205 35686 -18171
rect 35870 -18205 35882 -18171
rect 35674 -18211 35882 -18205
rect 34368 -18278 34428 -18211
rect 34826 -18278 34886 -18211
rect 35294 -18278 35354 -18211
rect 35750 -18278 35810 -18211
rect 34362 -18338 34368 -18278
rect 34428 -18338 34434 -18278
rect 34820 -18338 34826 -18278
rect 34886 -18338 34892 -18278
rect 35288 -18338 35294 -18278
rect 35354 -18338 35360 -18278
rect 35744 -18338 35750 -18278
rect 35810 -18338 35816 -18278
rect 35978 -18388 36038 -18112
rect 36442 -18112 36448 -16536
rect 36482 -16608 36504 -16536
rect 36900 -16536 36946 -16524
rect 36482 -18112 36488 -16608
rect 36900 -18052 36906 -16536
rect 36442 -18124 36488 -18112
rect 36894 -18112 36906 -18052
rect 36940 -18052 36946 -16536
rect 37352 -16536 37412 -16014
rect 37576 -16364 37582 -16304
rect 37642 -16364 37648 -16304
rect 38036 -16364 38042 -16304
rect 38102 -16364 38108 -16304
rect 37582 -16437 37642 -16364
rect 38042 -16437 38102 -16364
rect 37506 -16443 37714 -16437
rect 37506 -16477 37518 -16443
rect 37702 -16477 37714 -16443
rect 37506 -16483 37714 -16477
rect 37964 -16443 38172 -16437
rect 37964 -16477 37976 -16443
rect 38160 -16477 38172 -16443
rect 37964 -16483 38172 -16477
rect 37352 -16614 37364 -16536
rect 36940 -18112 36954 -18052
rect 36132 -18171 36340 -18165
rect 36132 -18205 36144 -18171
rect 36328 -18205 36340 -18171
rect 36132 -18211 36340 -18205
rect 36590 -18171 36798 -18165
rect 36590 -18205 36602 -18171
rect 36786 -18205 36798 -18171
rect 36590 -18211 36798 -18205
rect 36200 -18278 36260 -18211
rect 36664 -18278 36724 -18211
rect 36194 -18338 36200 -18278
rect 36260 -18338 36266 -18278
rect 36658 -18338 36664 -18278
rect 36724 -18338 36730 -18278
rect 34148 -18448 36038 -18388
rect 36894 -18512 36954 -18112
rect 37358 -18112 37364 -16614
rect 37398 -16614 37412 -16536
rect 37816 -16536 37862 -16524
rect 37398 -18112 37404 -16614
rect 37816 -18054 37822 -16536
rect 37358 -18124 37404 -18112
rect 37810 -18112 37822 -18054
rect 37856 -18054 37862 -16536
rect 38270 -16536 38330 -15884
rect 39182 -15932 40116 -15872
rect 39182 -16304 39242 -15932
rect 40110 -16304 40116 -15932
rect 38492 -16364 38498 -16304
rect 38558 -16364 38564 -16304
rect 38728 -16364 40116 -16304
rect 38498 -16437 38558 -16364
rect 38422 -16443 38630 -16437
rect 38422 -16477 38434 -16443
rect 38618 -16477 38630 -16443
rect 38422 -16483 38630 -16477
rect 38270 -16620 38280 -16536
rect 37856 -18112 37870 -18054
rect 37048 -18171 37256 -18165
rect 37048 -18205 37060 -18171
rect 37244 -18205 37256 -18171
rect 37048 -18211 37256 -18205
rect 37506 -18171 37714 -18165
rect 37506 -18205 37518 -18171
rect 37702 -18205 37714 -18171
rect 37506 -18211 37714 -18205
rect 37122 -18278 37182 -18211
rect 37578 -18278 37638 -18211
rect 37116 -18338 37122 -18278
rect 37182 -18338 37188 -18278
rect 37572 -18338 37578 -18278
rect 37638 -18338 37644 -18278
rect 33232 -18572 36954 -18512
rect 37810 -18646 37870 -18112
rect 38274 -18112 38280 -16620
rect 38314 -16620 38330 -16536
rect 38728 -16536 38788 -16364
rect 38954 -16437 39014 -16364
rect 38880 -16443 39088 -16437
rect 38880 -16477 38892 -16443
rect 39076 -16477 39088 -16443
rect 38880 -16483 39088 -16477
rect 38728 -16580 38738 -16536
rect 38314 -18112 38320 -16620
rect 38732 -18048 38738 -16580
rect 38274 -18124 38320 -18112
rect 38726 -18112 38738 -18048
rect 38772 -16580 38788 -16536
rect 39182 -16536 39242 -16364
rect 38772 -18048 38778 -16580
rect 39182 -16596 39196 -16536
rect 38772 -18112 38786 -18048
rect 39190 -18080 39196 -16596
rect 37964 -18171 38172 -18165
rect 37964 -18205 37976 -18171
rect 38160 -18205 38172 -18171
rect 37964 -18211 38172 -18205
rect 38422 -18171 38630 -18165
rect 38422 -18205 38434 -18171
rect 38618 -18205 38630 -18171
rect 38422 -18211 38630 -18205
rect 38038 -18278 38098 -18211
rect 38494 -18278 38554 -18211
rect 38032 -18338 38038 -18278
rect 38098 -18338 38104 -18278
rect 38488 -18338 38494 -18278
rect 38554 -18338 38560 -18278
rect 32312 -18706 37870 -18646
rect 38726 -18900 38786 -18112
rect 39184 -18112 39196 -18080
rect 39230 -16596 39242 -16536
rect 39230 -18080 39236 -16596
rect 39230 -18112 39244 -18080
rect 38880 -18171 39088 -18165
rect 38880 -18205 38892 -18171
rect 39076 -18205 39088 -18171
rect 38880 -18211 39088 -18205
rect 38952 -18900 39012 -18211
rect 39184 -18900 39244 -18112
rect 30916 -18910 39272 -18900
rect 30916 -18996 30942 -18910
rect 31038 -18996 31362 -18910
rect 31458 -18996 31962 -18910
rect 32058 -18996 32562 -18910
rect 32658 -18996 33162 -18910
rect 33258 -18996 33762 -18910
rect 33858 -18996 34362 -18910
rect 34458 -18996 34962 -18910
rect 35058 -18996 35562 -18910
rect 35658 -18996 36162 -18910
rect 36258 -18996 36762 -18910
rect 36858 -18996 37362 -18910
rect 37458 -18996 37962 -18910
rect 38058 -18996 38562 -18910
rect 38658 -18996 39162 -18910
rect 39258 -18996 39272 -18910
rect 30916 -19010 39272 -18996
rect 29766 -19470 29878 -19186
rect 30478 -19470 30488 -19170
rect 39500 -19470 39510 -19170
rect 40110 -19186 40116 -16364
rect 40216 -19186 40222 -14014
rect 40110 -19470 40222 -19186
rect 29766 -19476 40222 -19470
rect 29766 -19576 29872 -19476
rect 40116 -19576 40222 -19476
rect 29766 -19582 40222 -19576
rect 25812 -20028 36268 -20022
rect 25812 -20128 25918 -20028
rect 36162 -20128 36268 -20028
rect 25812 -20134 36268 -20128
rect 25812 -20418 25924 -20134
rect 25812 -25590 25818 -20418
rect 25918 -23240 25924 -20418
rect 26524 -20434 26534 -20134
rect 35546 -20434 35556 -20134
rect 36156 -20418 36268 -20134
rect 26762 -20608 35118 -20594
rect 26762 -20694 26776 -20608
rect 26872 -20694 27376 -20608
rect 27472 -20694 27976 -20608
rect 28072 -20694 28576 -20608
rect 28672 -20694 29176 -20608
rect 29272 -20694 29776 -20608
rect 29872 -20694 30376 -20608
rect 30472 -20694 30976 -20608
rect 31072 -20694 31576 -20608
rect 31672 -20694 32176 -20608
rect 32272 -20694 32776 -20608
rect 32872 -20694 33376 -20608
rect 33472 -20694 33976 -20608
rect 34072 -20694 34576 -20608
rect 34672 -20694 34996 -20608
rect 35092 -20694 35118 -20608
rect 26762 -20704 35118 -20694
rect 26790 -21492 26850 -20704
rect 27022 -21393 27082 -20704
rect 26946 -21399 27154 -21393
rect 26946 -21433 26958 -21399
rect 27142 -21433 27154 -21399
rect 26946 -21439 27154 -21433
rect 26790 -21524 26804 -21492
rect 26798 -23008 26804 -21524
rect 26792 -23068 26804 -23008
rect 26838 -21524 26850 -21492
rect 27248 -21492 27308 -20704
rect 28164 -20958 33722 -20898
rect 27474 -21326 27480 -21266
rect 27540 -21326 27546 -21266
rect 27930 -21326 27936 -21266
rect 27996 -21326 28002 -21266
rect 27480 -21393 27540 -21326
rect 27936 -21393 27996 -21326
rect 27404 -21399 27612 -21393
rect 27404 -21433 27416 -21399
rect 27600 -21433 27612 -21399
rect 27404 -21439 27612 -21433
rect 27862 -21399 28070 -21393
rect 27862 -21433 27874 -21399
rect 28058 -21433 28070 -21399
rect 27862 -21439 28070 -21433
rect 26838 -23008 26844 -21524
rect 27248 -21556 27262 -21492
rect 26838 -23068 26852 -23008
rect 27256 -23024 27262 -21556
rect 26792 -23240 26852 -23068
rect 27246 -23068 27262 -23024
rect 27296 -21556 27308 -21492
rect 27714 -21492 27760 -21480
rect 27296 -23024 27302 -21556
rect 27714 -22984 27720 -21492
rect 27296 -23068 27306 -23024
rect 26946 -23127 27154 -23121
rect 26946 -23161 26958 -23127
rect 27142 -23161 27154 -23127
rect 26946 -23167 27154 -23161
rect 27020 -23240 27080 -23167
rect 27246 -23240 27306 -23068
rect 27704 -23068 27720 -22984
rect 27754 -22984 27760 -21492
rect 28164 -21492 28224 -20958
rect 29080 -21092 32802 -21032
rect 28390 -21326 28396 -21266
rect 28456 -21326 28462 -21266
rect 28846 -21326 28852 -21266
rect 28912 -21326 28918 -21266
rect 28396 -21393 28456 -21326
rect 28852 -21393 28912 -21326
rect 28320 -21399 28528 -21393
rect 28320 -21433 28332 -21399
rect 28516 -21433 28528 -21399
rect 28320 -21439 28528 -21433
rect 28778 -21399 28986 -21393
rect 28778 -21433 28790 -21399
rect 28974 -21433 28986 -21399
rect 28778 -21439 28986 -21433
rect 28164 -21550 28178 -21492
rect 27754 -23068 27764 -22984
rect 27404 -23127 27612 -23121
rect 27404 -23161 27416 -23127
rect 27600 -23161 27612 -23127
rect 27404 -23167 27612 -23161
rect 27476 -23240 27536 -23167
rect 25918 -23300 27306 -23240
rect 27470 -23300 27476 -23240
rect 27536 -23300 27542 -23240
rect 25918 -23672 25924 -23300
rect 26792 -23672 26852 -23300
rect 25918 -23732 26852 -23672
rect 27704 -23720 27764 -23068
rect 28172 -23068 28178 -21550
rect 28212 -21550 28224 -21492
rect 28630 -21492 28676 -21480
rect 28212 -23068 28218 -21550
rect 28630 -22990 28636 -21492
rect 28172 -23080 28218 -23068
rect 28622 -23068 28636 -22990
rect 28670 -22990 28676 -21492
rect 29080 -21492 29140 -21092
rect 29996 -21216 31886 -21156
rect 29304 -21326 29310 -21266
rect 29370 -21326 29376 -21266
rect 29768 -21326 29774 -21266
rect 29834 -21326 29840 -21266
rect 29310 -21393 29370 -21326
rect 29774 -21393 29834 -21326
rect 29236 -21399 29444 -21393
rect 29236 -21433 29248 -21399
rect 29432 -21433 29444 -21399
rect 29236 -21439 29444 -21433
rect 29694 -21399 29902 -21393
rect 29694 -21433 29706 -21399
rect 29890 -21433 29902 -21399
rect 29694 -21439 29902 -21433
rect 29080 -21552 29094 -21492
rect 28670 -23068 28682 -22990
rect 27862 -23127 28070 -23121
rect 27862 -23161 27874 -23127
rect 28058 -23161 28070 -23127
rect 27862 -23167 28070 -23161
rect 28320 -23127 28528 -23121
rect 28320 -23161 28332 -23127
rect 28516 -23161 28528 -23127
rect 28320 -23167 28528 -23161
rect 27932 -23240 27992 -23167
rect 28392 -23240 28452 -23167
rect 27926 -23300 27932 -23240
rect 27992 -23300 27998 -23240
rect 28386 -23300 28392 -23240
rect 28452 -23300 28458 -23240
rect 28622 -23590 28682 -23068
rect 29088 -23068 29094 -21552
rect 29128 -21552 29140 -21492
rect 29546 -21492 29592 -21480
rect 29128 -23068 29134 -21552
rect 29546 -22996 29552 -21492
rect 29088 -23080 29134 -23068
rect 29530 -23068 29552 -22996
rect 29586 -23068 29592 -21492
rect 29996 -21492 30056 -21216
rect 30218 -21326 30224 -21266
rect 30284 -21326 30290 -21266
rect 30674 -21326 30680 -21266
rect 30740 -21326 30746 -21266
rect 31142 -21326 31148 -21266
rect 31208 -21326 31214 -21266
rect 31600 -21326 31606 -21266
rect 31666 -21326 31672 -21266
rect 30224 -21393 30284 -21326
rect 30680 -21393 30740 -21326
rect 31148 -21393 31208 -21326
rect 31606 -21393 31666 -21326
rect 30152 -21399 30360 -21393
rect 30152 -21433 30164 -21399
rect 30348 -21433 30360 -21399
rect 30152 -21439 30360 -21433
rect 30610 -21399 30818 -21393
rect 30610 -21433 30622 -21399
rect 30806 -21433 30818 -21399
rect 30610 -21439 30818 -21433
rect 31068 -21399 31276 -21393
rect 31068 -21433 31080 -21399
rect 31264 -21433 31276 -21399
rect 31068 -21439 31276 -21433
rect 31526 -21399 31734 -21393
rect 31526 -21433 31538 -21399
rect 31722 -21433 31734 -21399
rect 31526 -21439 31734 -21433
rect 29996 -21570 30010 -21492
rect 29530 -23080 29592 -23068
rect 30004 -23068 30010 -21570
rect 30044 -21570 30056 -21492
rect 30462 -21492 30508 -21480
rect 30044 -23068 30050 -21570
rect 30462 -22988 30468 -21492
rect 30004 -23080 30050 -23068
rect 30454 -23068 30468 -22988
rect 30502 -22988 30508 -21492
rect 30920 -21492 30966 -21480
rect 30502 -23068 30514 -22988
rect 30920 -23046 30926 -21492
rect 28778 -23127 28986 -23121
rect 28778 -23161 28790 -23127
rect 28974 -23161 28986 -23127
rect 28778 -23167 28986 -23161
rect 29236 -23127 29444 -23121
rect 29236 -23161 29248 -23127
rect 29432 -23161 29444 -23127
rect 29236 -23167 29444 -23161
rect 28848 -23240 28908 -23167
rect 29306 -23240 29366 -23167
rect 28842 -23300 28848 -23240
rect 28908 -23300 28914 -23240
rect 29300 -23300 29306 -23240
rect 29366 -23300 29372 -23240
rect 29530 -23464 29590 -23080
rect 29694 -23127 29902 -23121
rect 29694 -23161 29706 -23127
rect 29890 -23161 29902 -23127
rect 29694 -23167 29902 -23161
rect 30152 -23127 30360 -23121
rect 30152 -23161 30164 -23127
rect 30348 -23161 30360 -23127
rect 30152 -23167 30360 -23161
rect 29770 -23240 29830 -23167
rect 30224 -23240 30284 -23167
rect 29764 -23300 29770 -23240
rect 29830 -23300 29836 -23240
rect 30218 -23300 30224 -23240
rect 30284 -23300 30290 -23240
rect 30454 -23348 30514 -23068
rect 30916 -23068 30926 -23046
rect 30960 -23046 30966 -21492
rect 31378 -21492 31424 -21480
rect 31378 -23040 31384 -21492
rect 30960 -23068 30976 -23046
rect 30610 -23127 30818 -23121
rect 30610 -23161 30622 -23127
rect 30806 -23161 30818 -23127
rect 30610 -23167 30818 -23161
rect 30682 -23238 30742 -23167
rect 30916 -23228 30976 -23068
rect 31372 -23068 31384 -23040
rect 31418 -23040 31424 -21492
rect 31826 -21492 31886 -21216
rect 32056 -21326 32062 -21266
rect 32122 -21326 32128 -21266
rect 32512 -21326 32518 -21266
rect 32578 -21326 32584 -21266
rect 32062 -21393 32122 -21326
rect 32518 -21393 32578 -21326
rect 31984 -21399 32192 -21393
rect 31984 -21433 31996 -21399
rect 32180 -21433 32192 -21399
rect 31984 -21439 32192 -21433
rect 32442 -21399 32650 -21393
rect 32442 -21433 32454 -21399
rect 32638 -21433 32650 -21399
rect 32442 -21439 32650 -21433
rect 31826 -21536 31842 -21492
rect 31418 -23068 31432 -23040
rect 31068 -23127 31276 -23121
rect 31068 -23161 31080 -23127
rect 31264 -23161 31276 -23127
rect 31068 -23167 31276 -23161
rect 30676 -23240 30748 -23238
rect 30676 -23300 30682 -23240
rect 30742 -23300 30748 -23240
rect 31142 -23232 31202 -23167
rect 30916 -23294 30976 -23288
rect 31130 -23238 31214 -23232
rect 31130 -23300 31142 -23238
rect 31202 -23300 31214 -23238
rect 31130 -23304 31214 -23300
rect 31372 -23348 31432 -23068
rect 31836 -23068 31842 -21536
rect 31876 -21536 31886 -21492
rect 32294 -21492 32340 -21480
rect 31876 -23068 31882 -21536
rect 32294 -23036 32300 -21492
rect 31836 -23080 31882 -23068
rect 32286 -23068 32300 -23036
rect 32334 -23036 32340 -21492
rect 32742 -21492 32802 -21092
rect 32968 -21326 32974 -21266
rect 33034 -21326 33040 -21266
rect 33424 -21326 33430 -21266
rect 33490 -21326 33496 -21266
rect 32974 -21393 33034 -21326
rect 33430 -21393 33490 -21326
rect 32900 -21399 33108 -21393
rect 32900 -21433 32912 -21399
rect 33096 -21433 33108 -21399
rect 32900 -21439 33108 -21433
rect 33358 -21399 33566 -21393
rect 33358 -21433 33370 -21399
rect 33554 -21433 33566 -21399
rect 33358 -21439 33566 -21433
rect 32742 -21550 32758 -21492
rect 32334 -23068 32346 -23036
rect 31526 -23127 31734 -23121
rect 31526 -23161 31538 -23127
rect 31722 -23161 31734 -23127
rect 31526 -23167 31734 -23161
rect 31984 -23127 32192 -23121
rect 31984 -23161 31996 -23127
rect 32180 -23161 32192 -23127
rect 31984 -23167 32192 -23161
rect 31598 -23240 31658 -23167
rect 32058 -23240 32118 -23167
rect 31592 -23300 31598 -23240
rect 31658 -23300 31664 -23240
rect 32052 -23300 32058 -23240
rect 32118 -23300 32124 -23240
rect 30454 -23408 31432 -23348
rect 32286 -23464 32346 -23068
rect 32752 -23068 32758 -21550
rect 32792 -21550 32802 -21492
rect 33210 -21492 33256 -21480
rect 32792 -23068 32798 -21550
rect 33210 -23000 33216 -21492
rect 32752 -23080 32798 -23068
rect 33206 -23068 33216 -23000
rect 33250 -23000 33256 -21492
rect 33662 -21492 33722 -20958
rect 33882 -21326 33888 -21266
rect 33948 -21326 33954 -21266
rect 34342 -21326 34348 -21266
rect 34408 -21326 34414 -21266
rect 33888 -21393 33948 -21326
rect 34348 -21393 34408 -21326
rect 33816 -21399 34024 -21393
rect 33816 -21433 33828 -21399
rect 34012 -21433 34024 -21399
rect 33816 -21439 34024 -21433
rect 34274 -21399 34482 -21393
rect 34274 -21433 34286 -21399
rect 34470 -21433 34482 -21399
rect 34274 -21439 34482 -21433
rect 33662 -21548 33674 -21492
rect 33250 -23068 33266 -23000
rect 32442 -23127 32650 -23121
rect 32442 -23161 32454 -23127
rect 32638 -23161 32650 -23127
rect 32442 -23167 32650 -23161
rect 32900 -23127 33108 -23121
rect 32900 -23161 32912 -23127
rect 33096 -23161 33108 -23127
rect 32900 -23167 33108 -23161
rect 32514 -23240 32574 -23167
rect 32970 -23240 33030 -23167
rect 32508 -23300 32514 -23240
rect 32574 -23300 32580 -23240
rect 32964 -23300 32970 -23240
rect 33030 -23300 33036 -23240
rect 29530 -23524 32346 -23464
rect 33206 -23590 33266 -23068
rect 33668 -23068 33674 -21548
rect 33708 -21548 33722 -21492
rect 34126 -21492 34172 -21480
rect 33708 -23068 33714 -21548
rect 34126 -23008 34132 -21492
rect 33668 -23080 33714 -23068
rect 34120 -23068 34132 -23008
rect 34166 -23008 34172 -21492
rect 34578 -21492 34638 -20704
rect 34808 -21393 34868 -20704
rect 34732 -21399 34940 -21393
rect 34732 -21433 34744 -21399
rect 34928 -21433 34940 -21399
rect 34732 -21439 34940 -21433
rect 34578 -21568 34590 -21492
rect 34584 -23006 34590 -21568
rect 34166 -23068 34180 -23008
rect 33358 -23127 33566 -23121
rect 33358 -23161 33370 -23127
rect 33554 -23161 33566 -23127
rect 33358 -23167 33566 -23161
rect 33816 -23127 34024 -23121
rect 33816 -23161 33828 -23127
rect 34012 -23161 34024 -23127
rect 33816 -23167 34024 -23161
rect 33426 -23240 33486 -23167
rect 33884 -23240 33944 -23167
rect 33420 -23300 33426 -23240
rect 33486 -23300 33492 -23240
rect 33878 -23300 33884 -23240
rect 33944 -23300 33950 -23240
rect 28622 -23650 33266 -23590
rect 34120 -23720 34180 -23068
rect 34574 -23068 34590 -23006
rect 34624 -21568 34638 -21492
rect 35036 -21492 35096 -20704
rect 35036 -21562 35048 -21492
rect 34624 -23006 34630 -21568
rect 34624 -23068 34634 -23006
rect 35042 -23024 35048 -21562
rect 34274 -23127 34482 -23121
rect 34274 -23161 34286 -23127
rect 34470 -23161 34482 -23127
rect 34274 -23167 34482 -23161
rect 34344 -23240 34404 -23167
rect 34338 -23300 34344 -23240
rect 34404 -23300 34410 -23240
rect 34574 -23242 34634 -23068
rect 35032 -23068 35048 -23024
rect 35082 -21562 35096 -21492
rect 35082 -23024 35088 -21562
rect 35082 -23068 35092 -23024
rect 34732 -23127 34940 -23121
rect 34732 -23161 34744 -23127
rect 34928 -23161 34940 -23127
rect 34732 -23167 34940 -23161
rect 34806 -23242 34866 -23167
rect 35032 -23242 35092 -23068
rect 36156 -23242 36162 -20418
rect 34574 -23302 36162 -23242
rect 25918 -25590 25924 -23732
rect 26232 -24157 26292 -23732
rect 26460 -24058 26520 -23732
rect 27704 -23780 34180 -23720
rect 35032 -23736 35092 -23302
rect 36156 -23736 36162 -23302
rect 35032 -23796 36162 -23736
rect 26684 -23886 26690 -23826
rect 26750 -23886 26756 -23826
rect 26387 -24064 26595 -24058
rect 26387 -24098 26399 -24064
rect 26583 -24098 26595 -24064
rect 26387 -24104 26595 -24098
rect 26232 -24204 26245 -24157
rect 26239 -25312 26245 -24204
rect 25812 -25766 25924 -25590
rect 26232 -25333 26245 -25312
rect 26279 -24204 26292 -24157
rect 26690 -24157 26750 -23886
rect 26922 -23988 30186 -23928
rect 26922 -24058 26982 -23988
rect 27384 -24058 27444 -23988
rect 27838 -24058 27898 -23988
rect 28300 -24058 28360 -23988
rect 28754 -24058 28814 -23988
rect 29204 -24058 29264 -23988
rect 29670 -24058 29730 -23988
rect 30126 -24058 30186 -23988
rect 30582 -24006 31750 -23946
rect 30582 -24058 30642 -24006
rect 26845 -24064 27053 -24058
rect 26845 -24098 26857 -24064
rect 27041 -24098 27053 -24064
rect 26845 -24104 27053 -24098
rect 27303 -24064 27511 -24058
rect 27303 -24098 27315 -24064
rect 27499 -24098 27511 -24064
rect 27303 -24104 27511 -24098
rect 27761 -24064 27969 -24058
rect 27761 -24098 27773 -24064
rect 27957 -24098 27969 -24064
rect 27761 -24104 27969 -24098
rect 28219 -24064 28427 -24058
rect 28219 -24098 28231 -24064
rect 28415 -24098 28427 -24064
rect 28219 -24104 28427 -24098
rect 28677 -24064 28885 -24058
rect 28677 -24098 28689 -24064
rect 28873 -24098 28885 -24064
rect 28677 -24104 28885 -24098
rect 29135 -24064 29343 -24058
rect 29135 -24098 29147 -24064
rect 29331 -24098 29343 -24064
rect 29135 -24104 29343 -24098
rect 29593 -24064 29801 -24058
rect 29593 -24098 29605 -24064
rect 29789 -24098 29801 -24064
rect 29593 -24104 29801 -24098
rect 30051 -24064 30259 -24058
rect 30051 -24098 30063 -24064
rect 30247 -24098 30259 -24064
rect 30051 -24104 30259 -24098
rect 30509 -24064 30717 -24058
rect 30509 -24098 30521 -24064
rect 30705 -24098 30717 -24064
rect 30509 -24104 30717 -24098
rect 26279 -25312 26285 -24204
rect 26690 -24224 26703 -24157
rect 26279 -25333 26292 -25312
rect 26232 -25766 26292 -25333
rect 26697 -25333 26703 -24224
rect 26737 -24224 26750 -24157
rect 27155 -24157 27201 -24145
rect 26737 -25333 26743 -24224
rect 26697 -25345 26743 -25333
rect 27155 -25333 27161 -24157
rect 27195 -25333 27201 -24157
rect 27155 -25345 27201 -25333
rect 27613 -24157 27659 -24145
rect 27613 -25333 27619 -24157
rect 27653 -25333 27659 -24157
rect 27613 -25345 27659 -25333
rect 28071 -24157 28117 -24145
rect 28071 -25333 28077 -24157
rect 28111 -25333 28117 -24157
rect 28071 -25345 28117 -25333
rect 28529 -24157 28575 -24145
rect 28529 -25333 28535 -24157
rect 28569 -25333 28575 -24157
rect 28529 -25345 28575 -25333
rect 28987 -24157 29033 -24145
rect 28987 -25333 28993 -24157
rect 29027 -25333 29033 -24157
rect 28987 -25345 29033 -25333
rect 29445 -24157 29491 -24145
rect 29445 -25333 29451 -24157
rect 29485 -25333 29491 -24157
rect 29445 -25345 29491 -25333
rect 29903 -24157 29949 -24145
rect 29903 -25333 29909 -24157
rect 29943 -25333 29949 -24157
rect 30361 -24157 30407 -24145
rect 30361 -25266 30367 -24157
rect 29903 -25345 29949 -25333
rect 30352 -25333 30367 -25266
rect 30401 -25266 30407 -24157
rect 30812 -24157 30872 -24006
rect 30812 -24172 30825 -24157
rect 30401 -25333 30412 -25266
rect 30819 -25298 30825 -24172
rect 26387 -25392 26595 -25386
rect 26387 -25426 26399 -25392
rect 26583 -25426 26595 -25392
rect 26387 -25432 26595 -25426
rect 26845 -25392 27053 -25386
rect 26845 -25426 26857 -25392
rect 27041 -25426 27053 -25392
rect 26845 -25432 27053 -25426
rect 27303 -25392 27511 -25386
rect 27303 -25426 27315 -25392
rect 27499 -25426 27511 -25392
rect 27303 -25432 27511 -25426
rect 27761 -25392 27969 -25386
rect 27761 -25426 27773 -25392
rect 27957 -25426 27969 -25392
rect 27761 -25432 27969 -25426
rect 28219 -25392 28427 -25386
rect 28219 -25426 28231 -25392
rect 28415 -25426 28427 -25392
rect 28219 -25432 28427 -25426
rect 28677 -25392 28885 -25386
rect 28677 -25426 28689 -25392
rect 28873 -25426 28885 -25392
rect 28677 -25432 28885 -25426
rect 29135 -25392 29343 -25386
rect 29135 -25426 29147 -25392
rect 29331 -25426 29343 -25392
rect 29135 -25432 29343 -25426
rect 29593 -25392 29801 -25386
rect 29593 -25426 29605 -25392
rect 29789 -25426 29801 -25392
rect 29593 -25432 29801 -25426
rect 30051 -25392 30259 -25386
rect 30051 -25426 30063 -25392
rect 30247 -25426 30259 -25392
rect 30051 -25432 30259 -25426
rect 26460 -25766 26520 -25432
rect 26914 -25500 26974 -25432
rect 27376 -25500 27436 -25432
rect 27830 -25500 27890 -25432
rect 28292 -25500 28352 -25432
rect 28746 -25500 28806 -25432
rect 29196 -25500 29256 -25432
rect 29662 -25500 29722 -25432
rect 30118 -25500 30178 -25432
rect 26914 -25504 27830 -25500
rect 26974 -25560 27376 -25504
rect 26914 -25570 26974 -25564
rect 27436 -25560 27830 -25504
rect 27890 -25560 28292 -25500
rect 28352 -25506 29196 -25500
rect 28352 -25560 28746 -25506
rect 27376 -25570 27436 -25564
rect 27830 -25566 27890 -25560
rect 28292 -25566 28352 -25560
rect 28806 -25560 29196 -25506
rect 29256 -25560 29662 -25500
rect 29722 -25504 30178 -25500
rect 29722 -25560 30118 -25504
rect 29196 -25566 29256 -25560
rect 29662 -25566 29722 -25560
rect 28746 -25572 28806 -25566
rect 30118 -25570 30178 -25564
rect 30352 -25626 30412 -25333
rect 30810 -25333 30825 -25298
rect 30859 -24172 30872 -24157
rect 31232 -24157 31292 -24006
rect 31464 -24058 31524 -24006
rect 31387 -24064 31595 -24058
rect 31387 -24098 31399 -24064
rect 31583 -24098 31595 -24064
rect 31387 -24104 31595 -24098
rect 30859 -25298 30865 -24172
rect 31232 -24178 31245 -24157
rect 31239 -25298 31245 -24178
rect 30859 -25333 30870 -25298
rect 30509 -25392 30717 -25386
rect 30509 -25426 30521 -25392
rect 30705 -25426 30717 -25392
rect 30509 -25432 30717 -25426
rect 30346 -25686 30352 -25626
rect 30412 -25686 30418 -25626
rect 30582 -25766 30642 -25432
rect 30810 -25766 30870 -25333
rect 31230 -25333 31245 -25298
rect 31279 -24178 31292 -24157
rect 31690 -24157 31750 -24006
rect 31916 -23988 35180 -23928
rect 31916 -24058 31976 -23988
rect 32378 -24058 32438 -23988
rect 32832 -24058 32892 -23988
rect 33294 -24058 33354 -23988
rect 33748 -24058 33808 -23988
rect 34198 -24058 34258 -23988
rect 34664 -24058 34724 -23988
rect 35120 -24058 35180 -23988
rect 35582 -24058 35642 -23796
rect 31845 -24064 32053 -24058
rect 31845 -24098 31857 -24064
rect 32041 -24098 32053 -24064
rect 31845 -24104 32053 -24098
rect 32303 -24064 32511 -24058
rect 32303 -24098 32315 -24064
rect 32499 -24098 32511 -24064
rect 32303 -24104 32511 -24098
rect 32761 -24064 32969 -24058
rect 32761 -24098 32773 -24064
rect 32957 -24098 32969 -24064
rect 32761 -24104 32969 -24098
rect 33219 -24064 33427 -24058
rect 33219 -24098 33231 -24064
rect 33415 -24098 33427 -24064
rect 33219 -24104 33427 -24098
rect 33677 -24064 33885 -24058
rect 33677 -24098 33689 -24064
rect 33873 -24098 33885 -24064
rect 33677 -24104 33885 -24098
rect 34135 -24064 34343 -24058
rect 34135 -24098 34147 -24064
rect 34331 -24098 34343 -24064
rect 34135 -24104 34343 -24098
rect 34593 -24064 34801 -24058
rect 34593 -24098 34605 -24064
rect 34789 -24098 34801 -24064
rect 34593 -24104 34801 -24098
rect 35051 -24064 35259 -24058
rect 35051 -24098 35063 -24064
rect 35247 -24098 35259 -24064
rect 35051 -24104 35259 -24098
rect 35509 -24064 35717 -24058
rect 35509 -24098 35521 -24064
rect 35705 -24098 35717 -24064
rect 35509 -24104 35717 -24098
rect 31279 -25298 31285 -24178
rect 31690 -24200 31703 -24157
rect 31697 -25292 31703 -24200
rect 31279 -25333 31290 -25298
rect 31230 -25766 31290 -25333
rect 31688 -25333 31703 -25292
rect 31737 -24200 31750 -24157
rect 32155 -24157 32201 -24145
rect 31737 -25292 31743 -24200
rect 31737 -25333 31748 -25292
rect 31387 -25392 31595 -25386
rect 31387 -25426 31399 -25392
rect 31583 -25426 31595 -25392
rect 31387 -25432 31595 -25426
rect 31458 -25766 31518 -25432
rect 31688 -25766 31748 -25333
rect 32155 -25333 32161 -24157
rect 32195 -25333 32201 -24157
rect 32155 -25345 32201 -25333
rect 32613 -24157 32659 -24145
rect 32613 -25333 32619 -24157
rect 32653 -25333 32659 -24157
rect 32613 -25345 32659 -25333
rect 33071 -24157 33117 -24145
rect 33071 -25333 33077 -24157
rect 33111 -25333 33117 -24157
rect 33071 -25345 33117 -25333
rect 33529 -24157 33575 -24145
rect 33529 -25333 33535 -24157
rect 33569 -25333 33575 -24157
rect 33529 -25345 33575 -25333
rect 33987 -24157 34033 -24145
rect 33987 -25333 33993 -24157
rect 34027 -25333 34033 -24157
rect 33987 -25345 34033 -25333
rect 34445 -24157 34491 -24145
rect 34445 -25333 34451 -24157
rect 34485 -25333 34491 -24157
rect 34445 -25345 34491 -25333
rect 34903 -24157 34949 -24145
rect 34903 -25333 34909 -24157
rect 34943 -25333 34949 -24157
rect 35361 -24157 35407 -24145
rect 35361 -25326 35367 -24157
rect 34903 -25345 34949 -25333
rect 35352 -25333 35367 -25326
rect 35401 -25326 35407 -24157
rect 35808 -24157 35868 -23796
rect 35808 -24210 35825 -24157
rect 35819 -25300 35825 -24210
rect 35401 -25333 35412 -25326
rect 31845 -25392 32053 -25386
rect 31845 -25426 31857 -25392
rect 32041 -25426 32053 -25392
rect 31845 -25432 32053 -25426
rect 32303 -25392 32511 -25386
rect 32303 -25426 32315 -25392
rect 32499 -25426 32511 -25392
rect 32303 -25432 32511 -25426
rect 32761 -25392 32969 -25386
rect 32761 -25426 32773 -25392
rect 32957 -25426 32969 -25392
rect 32761 -25432 32969 -25426
rect 33219 -25392 33427 -25386
rect 33219 -25426 33231 -25392
rect 33415 -25426 33427 -25392
rect 33219 -25432 33427 -25426
rect 33677 -25392 33885 -25386
rect 33677 -25426 33689 -25392
rect 33873 -25426 33885 -25392
rect 33677 -25432 33885 -25426
rect 34135 -25392 34343 -25386
rect 34135 -25426 34147 -25392
rect 34331 -25426 34343 -25392
rect 34135 -25432 34343 -25426
rect 34593 -25392 34801 -25386
rect 34593 -25426 34605 -25392
rect 34789 -25426 34801 -25392
rect 34593 -25432 34801 -25426
rect 35051 -25392 35259 -25386
rect 35051 -25426 35063 -25392
rect 35247 -25426 35259 -25392
rect 35051 -25432 35259 -25426
rect 31916 -25500 31976 -25432
rect 32378 -25496 32438 -25432
rect 31916 -25504 32378 -25500
rect 31976 -25556 32378 -25504
rect 32832 -25500 32892 -25432
rect 33294 -25500 33354 -25432
rect 33748 -25500 33808 -25432
rect 34198 -25496 34258 -25432
rect 32438 -25502 34198 -25500
rect 32438 -25556 32832 -25502
rect 31976 -25560 32832 -25556
rect 32378 -25562 32438 -25560
rect 32892 -25560 33294 -25502
rect 31916 -25570 31976 -25564
rect 32832 -25568 32892 -25562
rect 33354 -25560 33748 -25502
rect 33294 -25568 33354 -25562
rect 33808 -25556 34198 -25502
rect 34664 -25500 34724 -25432
rect 35120 -25500 35180 -25432
rect 34258 -25502 35180 -25500
rect 34258 -25556 34664 -25502
rect 33808 -25560 34664 -25556
rect 34198 -25562 34258 -25560
rect 34724 -25560 35120 -25502
rect 33748 -25568 33808 -25562
rect 34664 -25568 34724 -25562
rect 35120 -25568 35180 -25562
rect 35352 -25632 35412 -25333
rect 35810 -25333 35825 -25300
rect 35859 -24210 35868 -24157
rect 35859 -25300 35865 -24210
rect 35859 -25333 35870 -25300
rect 35509 -25392 35717 -25386
rect 35509 -25426 35521 -25392
rect 35705 -25426 35717 -25392
rect 35509 -25432 35717 -25426
rect 35352 -25698 35412 -25692
rect 35582 -25766 35642 -25432
rect 35810 -25766 35870 -25333
rect 36156 -25590 36162 -23796
rect 36262 -25590 36268 -20418
rect 36156 -25766 36268 -25590
rect 25812 -25772 36268 -25766
rect 25812 -25872 25918 -25772
rect 36162 -25872 36268 -25772
rect 25812 -25878 36268 -25872
rect 25812 -26108 36268 -26102
rect 25812 -26208 25918 -26108
rect 36162 -26208 36268 -26108
rect 25812 -26214 36268 -26208
rect 25812 -26338 25924 -26214
rect 25540 -27710 25546 -27650
rect 25606 -27710 25612 -27650
rect 21156 -28466 21268 -28342
rect 10812 -28472 21268 -28466
rect 10812 -28572 10918 -28472
rect 21162 -28572 21268 -28472
rect 10812 -28578 21268 -28572
rect 25812 -28342 25818 -26338
rect 25918 -28342 25924 -26338
rect 26232 -26650 26292 -26214
rect 26462 -26560 26522 -26214
rect 30352 -26306 30412 -26300
rect 26920 -26440 27376 -26434
rect 26908 -26500 26914 -26440
rect 26974 -26494 27376 -26440
rect 27436 -26440 28292 -26434
rect 27436 -26494 27830 -26440
rect 26974 -26500 26980 -26494
rect 26914 -26560 26980 -26500
rect 27376 -26560 27442 -26494
rect 27824 -26500 27830 -26494
rect 27890 -26494 28292 -26440
rect 28352 -26494 28746 -26434
rect 28806 -26494 29196 -26434
rect 29256 -26440 30118 -26434
rect 29256 -26494 29662 -26440
rect 27890 -26500 27896 -26494
rect 27830 -26560 27896 -26500
rect 28292 -26560 28358 -26494
rect 28746 -26560 28812 -26494
rect 29196 -26560 29262 -26494
rect 29656 -26500 29662 -26494
rect 29722 -26494 30118 -26440
rect 30178 -26494 30184 -26434
rect 29722 -26500 29728 -26494
rect 29662 -26560 29728 -26500
rect 30118 -26560 30184 -26494
rect 26386 -26566 26594 -26560
rect 26386 -26600 26398 -26566
rect 26582 -26600 26594 -26566
rect 26386 -26606 26594 -26600
rect 26844 -26566 27052 -26560
rect 26844 -26600 26856 -26566
rect 27040 -26600 27052 -26566
rect 26844 -26606 27052 -26600
rect 27302 -26566 27510 -26560
rect 27302 -26600 27314 -26566
rect 27498 -26600 27510 -26566
rect 27302 -26606 27510 -26600
rect 27760 -26566 27968 -26560
rect 27760 -26600 27772 -26566
rect 27956 -26600 27968 -26566
rect 27760 -26606 27968 -26600
rect 28218 -26566 28426 -26560
rect 28218 -26600 28230 -26566
rect 28414 -26600 28426 -26566
rect 28218 -26606 28426 -26600
rect 28676 -26566 28884 -26560
rect 28676 -26600 28688 -26566
rect 28872 -26600 28884 -26566
rect 28676 -26606 28884 -26600
rect 29134 -26566 29342 -26560
rect 29134 -26600 29146 -26566
rect 29330 -26600 29342 -26566
rect 29134 -26606 29342 -26600
rect 29592 -26566 29800 -26560
rect 29592 -26600 29604 -26566
rect 29788 -26600 29800 -26566
rect 29592 -26606 29800 -26600
rect 30050 -26566 30258 -26560
rect 30050 -26600 30062 -26566
rect 30246 -26600 30258 -26566
rect 30050 -26606 30258 -26600
rect 26232 -26690 26244 -26650
rect 26238 -26786 26244 -26690
rect 26232 -26826 26244 -26786
rect 26278 -26690 26292 -26650
rect 26696 -26650 26742 -26638
rect 26278 -26786 26284 -26690
rect 26696 -26784 26702 -26650
rect 26278 -26826 26292 -26786
rect 26232 -27042 26292 -26826
rect 26688 -26826 26702 -26784
rect 26736 -26784 26742 -26650
rect 27154 -26650 27200 -26638
rect 26736 -26826 26748 -26784
rect 26386 -26876 26594 -26870
rect 26386 -26910 26398 -26876
rect 26582 -26910 26594 -26876
rect 26386 -26916 26594 -26910
rect 26460 -27042 26520 -26916
rect 26232 -27102 26520 -27042
rect 26232 -27318 26292 -27102
rect 26460 -27228 26520 -27102
rect 26386 -27234 26594 -27228
rect 26386 -27268 26398 -27234
rect 26582 -27268 26594 -27234
rect 26386 -27274 26594 -27268
rect 26232 -27338 26244 -27318
rect 26238 -27464 26244 -27338
rect 26224 -27494 26244 -27464
rect 26278 -27338 26292 -27318
rect 26688 -27318 26748 -26826
rect 27154 -26826 27160 -26650
rect 27194 -26826 27200 -26650
rect 27154 -26838 27200 -26826
rect 27612 -26650 27658 -26638
rect 27612 -26826 27618 -26650
rect 27652 -26826 27658 -26650
rect 27612 -26838 27658 -26826
rect 28070 -26650 28116 -26638
rect 28070 -26826 28076 -26650
rect 28110 -26826 28116 -26650
rect 28070 -26838 28116 -26826
rect 28528 -26650 28574 -26638
rect 28528 -26826 28534 -26650
rect 28568 -26826 28574 -26650
rect 28528 -26838 28574 -26826
rect 28986 -26650 29032 -26638
rect 28986 -26826 28992 -26650
rect 29026 -26826 29032 -26650
rect 28986 -26838 29032 -26826
rect 29444 -26650 29490 -26638
rect 29444 -26826 29450 -26650
rect 29484 -26826 29490 -26650
rect 29444 -26838 29490 -26826
rect 29902 -26650 29948 -26638
rect 29902 -26826 29908 -26650
rect 29942 -26826 29948 -26650
rect 30352 -26650 30412 -26366
rect 30580 -26560 30640 -26214
rect 30508 -26566 30716 -26560
rect 30508 -26600 30520 -26566
rect 30704 -26600 30716 -26566
rect 30508 -26606 30716 -26600
rect 30352 -26680 30366 -26650
rect 29902 -26838 29948 -26826
rect 30360 -26826 30366 -26680
rect 30400 -26680 30412 -26650
rect 30812 -26650 30872 -26214
rect 30812 -26678 30824 -26650
rect 30400 -26826 30406 -26680
rect 30818 -26770 30824 -26678
rect 30360 -26838 30406 -26826
rect 30812 -26826 30824 -26770
rect 30858 -26678 30872 -26650
rect 31232 -26650 31292 -26214
rect 31466 -26560 31526 -26214
rect 31386 -26566 31594 -26560
rect 31386 -26600 31398 -26566
rect 31582 -26600 31594 -26566
rect 31386 -26606 31594 -26600
rect 30858 -26770 30864 -26678
rect 31232 -26686 31244 -26650
rect 30858 -26826 30872 -26770
rect 31238 -26790 31244 -26686
rect 26844 -26876 27052 -26870
rect 26844 -26910 26856 -26876
rect 27040 -26910 27052 -26876
rect 26844 -26916 27052 -26910
rect 27302 -26876 27510 -26870
rect 27302 -26910 27314 -26876
rect 27498 -26910 27510 -26876
rect 27302 -26916 27510 -26910
rect 27760 -26876 27968 -26870
rect 27760 -26910 27772 -26876
rect 27956 -26910 27968 -26876
rect 27760 -26916 27968 -26910
rect 28218 -26876 28426 -26870
rect 28218 -26910 28230 -26876
rect 28414 -26910 28426 -26876
rect 28218 -26916 28426 -26910
rect 28676 -26876 28884 -26870
rect 28676 -26910 28688 -26876
rect 28872 -26910 28884 -26876
rect 28676 -26916 28884 -26910
rect 29134 -26876 29342 -26870
rect 29134 -26910 29146 -26876
rect 29330 -26910 29342 -26876
rect 29134 -26916 29342 -26910
rect 29592 -26876 29800 -26870
rect 29592 -26910 29604 -26876
rect 29788 -26910 29800 -26876
rect 29592 -26916 29800 -26910
rect 30050 -26876 30258 -26870
rect 30050 -26910 30062 -26876
rect 30246 -26910 30258 -26876
rect 30050 -26916 30258 -26910
rect 30508 -26876 30716 -26870
rect 30508 -26910 30520 -26876
rect 30704 -26910 30716 -26876
rect 30508 -26916 30716 -26910
rect 26914 -26982 26974 -26916
rect 27376 -26982 27436 -26916
rect 27830 -26982 27890 -26916
rect 28292 -26982 28352 -26916
rect 28746 -26982 28806 -26916
rect 29196 -26982 29256 -26916
rect 29662 -26982 29722 -26916
rect 30118 -26982 30178 -26916
rect 26914 -27042 30178 -26982
rect 26920 -27162 30184 -27102
rect 26920 -27228 26980 -27162
rect 27382 -27228 27442 -27162
rect 27836 -27228 27896 -27162
rect 28298 -27228 28358 -27162
rect 28752 -27228 28812 -27162
rect 29202 -27228 29262 -27162
rect 29668 -27228 29728 -27162
rect 30124 -27228 30184 -27162
rect 30580 -27228 30640 -26916
rect 26844 -27234 27052 -27228
rect 26844 -27268 26856 -27234
rect 27040 -27268 27052 -27234
rect 26844 -27274 27052 -27268
rect 27302 -27234 27510 -27228
rect 27302 -27268 27314 -27234
rect 27498 -27268 27510 -27234
rect 27302 -27274 27510 -27268
rect 27760 -27234 27968 -27228
rect 27760 -27268 27772 -27234
rect 27956 -27268 27968 -27234
rect 27760 -27274 27968 -27268
rect 28218 -27234 28426 -27228
rect 28218 -27268 28230 -27234
rect 28414 -27268 28426 -27234
rect 28218 -27274 28426 -27268
rect 28676 -27234 28884 -27228
rect 28676 -27268 28688 -27234
rect 28872 -27268 28884 -27234
rect 28676 -27274 28884 -27268
rect 29134 -27234 29342 -27228
rect 29134 -27268 29146 -27234
rect 29330 -27268 29342 -27234
rect 29134 -27274 29342 -27268
rect 29592 -27234 29800 -27228
rect 29592 -27268 29604 -27234
rect 29788 -27268 29800 -27234
rect 29592 -27274 29800 -27268
rect 30050 -27234 30258 -27228
rect 30050 -27268 30062 -27234
rect 30246 -27268 30258 -27234
rect 30050 -27274 30258 -27268
rect 30508 -27234 30716 -27228
rect 30508 -27268 30520 -27234
rect 30704 -27268 30716 -27234
rect 30508 -27274 30716 -27268
rect 26278 -27494 26284 -27338
rect 26688 -27346 26702 -27318
rect 26224 -27874 26284 -27494
rect 26696 -27494 26702 -27346
rect 26736 -27346 26748 -27318
rect 27154 -27318 27200 -27306
rect 26736 -27494 26742 -27346
rect 26696 -27506 26742 -27494
rect 27154 -27494 27160 -27318
rect 27194 -27494 27200 -27318
rect 27154 -27506 27200 -27494
rect 27612 -27318 27658 -27306
rect 27612 -27494 27618 -27318
rect 27652 -27494 27658 -27318
rect 27612 -27506 27658 -27494
rect 28070 -27318 28116 -27306
rect 28070 -27494 28076 -27318
rect 28110 -27494 28116 -27318
rect 28070 -27506 28116 -27494
rect 28528 -27318 28574 -27306
rect 28528 -27494 28534 -27318
rect 28568 -27494 28574 -27318
rect 28528 -27506 28574 -27494
rect 28986 -27318 29032 -27306
rect 28986 -27494 28992 -27318
rect 29026 -27494 29032 -27318
rect 28986 -27506 29032 -27494
rect 29444 -27318 29490 -27306
rect 29444 -27494 29450 -27318
rect 29484 -27494 29490 -27318
rect 29444 -27506 29490 -27494
rect 29902 -27318 29948 -27306
rect 29902 -27494 29908 -27318
rect 29942 -27494 29948 -27318
rect 30360 -27318 30406 -27306
rect 30360 -27466 30366 -27318
rect 29902 -27506 29948 -27494
rect 30352 -27494 30366 -27466
rect 30400 -27466 30406 -27318
rect 30812 -27318 30872 -26826
rect 30400 -27494 30412 -27466
rect 26386 -27544 26594 -27538
rect 26386 -27578 26398 -27544
rect 26582 -27578 26594 -27544
rect 26386 -27584 26594 -27578
rect 26844 -27544 27052 -27538
rect 26844 -27578 26856 -27544
rect 27040 -27578 27052 -27544
rect 26844 -27584 27052 -27578
rect 27302 -27544 27510 -27538
rect 27302 -27578 27314 -27544
rect 27498 -27578 27510 -27544
rect 27302 -27584 27510 -27578
rect 27760 -27544 27968 -27538
rect 27760 -27578 27772 -27544
rect 27956 -27578 27968 -27544
rect 27760 -27584 27968 -27578
rect 28218 -27544 28426 -27538
rect 28218 -27578 28230 -27544
rect 28414 -27578 28426 -27544
rect 28218 -27584 28426 -27578
rect 28676 -27544 28884 -27538
rect 28676 -27578 28688 -27544
rect 28872 -27578 28884 -27544
rect 28676 -27584 28884 -27578
rect 29134 -27544 29342 -27538
rect 29134 -27578 29146 -27544
rect 29330 -27578 29342 -27544
rect 29134 -27584 29342 -27578
rect 29592 -27544 29800 -27538
rect 29592 -27578 29604 -27544
rect 29788 -27578 29800 -27544
rect 29592 -27584 29800 -27578
rect 30050 -27544 30258 -27538
rect 30050 -27578 30062 -27544
rect 30246 -27578 30258 -27544
rect 30050 -27584 30258 -27578
rect 26464 -27874 26524 -27584
rect 26914 -27650 26974 -27584
rect 27376 -27650 27436 -27584
rect 27830 -27650 27890 -27584
rect 28292 -27650 28352 -27584
rect 28746 -27650 28806 -27584
rect 29196 -27650 29256 -27584
rect 29662 -27650 29722 -27584
rect 30118 -27650 30178 -27584
rect 26908 -27710 26914 -27650
rect 26974 -27710 30178 -27650
rect 30352 -27874 30412 -27494
rect 30812 -27494 30824 -27318
rect 30858 -27494 30872 -27318
rect 30508 -27544 30716 -27538
rect 30508 -27578 30520 -27544
rect 30704 -27578 30716 -27544
rect 30508 -27584 30716 -27578
rect 30578 -27874 30638 -27584
rect 30812 -27874 30872 -27494
rect 31228 -26826 31244 -26790
rect 31278 -26686 31292 -26650
rect 31688 -26650 31748 -26214
rect 35346 -26354 35352 -26294
rect 35412 -26354 35418 -26294
rect 34192 -26434 34198 -26430
rect 31910 -26494 31916 -26434
rect 31976 -26436 34198 -26434
rect 31976 -26494 32378 -26436
rect 31916 -26560 31980 -26494
rect 32372 -26496 32378 -26494
rect 32438 -26494 32832 -26436
rect 32438 -26496 32444 -26494
rect 32826 -26496 32832 -26494
rect 32892 -26494 33294 -26436
rect 32892 -26496 32898 -26494
rect 33288 -26496 33294 -26494
rect 33354 -26494 33748 -26436
rect 33354 -26496 33360 -26494
rect 33742 -26496 33748 -26494
rect 33808 -26490 34198 -26436
rect 34258 -26434 34264 -26430
rect 34258 -26490 34664 -26434
rect 33808 -26494 34664 -26490
rect 34724 -26494 35120 -26434
rect 35180 -26494 35186 -26434
rect 33808 -26496 33814 -26494
rect 32378 -26560 32442 -26496
rect 32832 -26560 32896 -26496
rect 33294 -26560 33358 -26496
rect 33748 -26560 33812 -26496
rect 34198 -26560 34262 -26494
rect 34664 -26560 34728 -26494
rect 35120 -26560 35184 -26494
rect 31844 -26566 32052 -26560
rect 31844 -26600 31856 -26566
rect 32040 -26600 32052 -26566
rect 31844 -26606 32052 -26600
rect 32302 -26566 32510 -26560
rect 32302 -26600 32314 -26566
rect 32498 -26600 32510 -26566
rect 32302 -26606 32510 -26600
rect 32760 -26566 32968 -26560
rect 32760 -26600 32772 -26566
rect 32956 -26600 32968 -26566
rect 32760 -26606 32968 -26600
rect 33218 -26566 33426 -26560
rect 33218 -26600 33230 -26566
rect 33414 -26600 33426 -26566
rect 33218 -26606 33426 -26600
rect 33676 -26566 33884 -26560
rect 33676 -26600 33688 -26566
rect 33872 -26600 33884 -26566
rect 33676 -26606 33884 -26600
rect 34134 -26566 34342 -26560
rect 34134 -26600 34146 -26566
rect 34330 -26600 34342 -26566
rect 34134 -26606 34342 -26600
rect 34592 -26566 34800 -26560
rect 34592 -26600 34604 -26566
rect 34788 -26600 34800 -26566
rect 34592 -26606 34800 -26600
rect 35050 -26566 35258 -26560
rect 35050 -26600 35062 -26566
rect 35246 -26600 35258 -26566
rect 35050 -26606 35258 -26600
rect 31278 -26790 31284 -26686
rect 31688 -26714 31702 -26650
rect 31696 -26782 31702 -26714
rect 31278 -26826 31288 -26790
rect 31228 -26980 31288 -26826
rect 31688 -26826 31702 -26782
rect 31736 -26714 31748 -26650
rect 32154 -26650 32200 -26638
rect 31736 -26782 31742 -26714
rect 31736 -26826 31748 -26782
rect 31386 -26876 31594 -26870
rect 31386 -26910 31398 -26876
rect 31582 -26910 31594 -26876
rect 31386 -26916 31594 -26910
rect 31456 -26980 31516 -26916
rect 31688 -26980 31748 -26826
rect 32154 -26826 32160 -26650
rect 32194 -26826 32200 -26650
rect 32154 -26838 32200 -26826
rect 32612 -26650 32658 -26638
rect 32612 -26826 32618 -26650
rect 32652 -26826 32658 -26650
rect 32612 -26838 32658 -26826
rect 33070 -26650 33116 -26638
rect 33070 -26826 33076 -26650
rect 33110 -26826 33116 -26650
rect 33070 -26838 33116 -26826
rect 33528 -26650 33574 -26638
rect 33528 -26826 33534 -26650
rect 33568 -26826 33574 -26650
rect 33528 -26838 33574 -26826
rect 33986 -26650 34032 -26638
rect 33986 -26826 33992 -26650
rect 34026 -26826 34032 -26650
rect 33986 -26838 34032 -26826
rect 34444 -26650 34490 -26638
rect 34444 -26826 34450 -26650
rect 34484 -26826 34490 -26650
rect 34444 -26838 34490 -26826
rect 34902 -26650 34948 -26638
rect 34902 -26826 34908 -26650
rect 34942 -26826 34948 -26650
rect 35352 -26650 35412 -26354
rect 35592 -26560 35652 -26214
rect 35508 -26566 35716 -26560
rect 35508 -26600 35520 -26566
rect 35704 -26600 35716 -26566
rect 35508 -26606 35716 -26600
rect 35352 -26692 35366 -26650
rect 34902 -26838 34948 -26826
rect 35360 -26826 35366 -26692
rect 35400 -26692 35412 -26650
rect 35810 -26650 35870 -26214
rect 35810 -26690 35824 -26650
rect 35400 -26826 35406 -26692
rect 35818 -26780 35824 -26690
rect 35360 -26838 35406 -26826
rect 35808 -26826 35824 -26780
rect 35858 -26690 35870 -26650
rect 36156 -26338 36268 -26214
rect 35858 -26780 35864 -26690
rect 35858 -26826 35868 -26780
rect 31844 -26876 32052 -26870
rect 31844 -26910 31856 -26876
rect 32040 -26910 32052 -26876
rect 31844 -26916 32052 -26910
rect 32302 -26876 32510 -26870
rect 32302 -26910 32314 -26876
rect 32498 -26910 32510 -26876
rect 32302 -26916 32510 -26910
rect 32760 -26876 32968 -26870
rect 32760 -26910 32772 -26876
rect 32956 -26910 32968 -26876
rect 32760 -26916 32968 -26910
rect 33218 -26876 33426 -26870
rect 33218 -26910 33230 -26876
rect 33414 -26910 33426 -26876
rect 33218 -26916 33426 -26910
rect 33676 -26876 33884 -26870
rect 33676 -26910 33688 -26876
rect 33872 -26910 33884 -26876
rect 33676 -26916 33884 -26910
rect 34134 -26876 34342 -26870
rect 34134 -26910 34146 -26876
rect 34330 -26910 34342 -26876
rect 34134 -26916 34342 -26910
rect 34592 -26876 34800 -26870
rect 34592 -26910 34604 -26876
rect 34788 -26910 34800 -26876
rect 34592 -26916 34800 -26910
rect 35050 -26876 35258 -26870
rect 35050 -26910 35062 -26876
rect 35246 -26910 35258 -26876
rect 35050 -26916 35258 -26910
rect 35508 -26876 35716 -26870
rect 35508 -26910 35520 -26876
rect 35704 -26910 35716 -26876
rect 35508 -26916 35716 -26910
rect 31228 -27040 31748 -26980
rect 31228 -27874 31288 -27040
rect 31456 -27874 31516 -27040
rect 31688 -27874 31748 -27040
rect 31914 -26982 31974 -26916
rect 32376 -26982 32436 -26916
rect 32830 -26982 32890 -26916
rect 33292 -26982 33352 -26916
rect 33746 -26982 33806 -26916
rect 34196 -26982 34256 -26916
rect 34662 -26982 34722 -26916
rect 35118 -26982 35178 -26916
rect 31914 -27042 35178 -26982
rect 35582 -27874 35642 -26916
rect 35808 -27874 35868 -26826
rect 26160 -27902 35930 -27874
rect 26160 -27988 26210 -27902
rect 26306 -27988 26790 -27902
rect 26886 -27988 27390 -27902
rect 27486 -27988 27990 -27902
rect 28086 -27988 28590 -27902
rect 28686 -27988 29190 -27902
rect 29286 -27988 29790 -27902
rect 29886 -27988 30390 -27902
rect 30486 -27988 30990 -27902
rect 31086 -27988 31590 -27902
rect 31686 -27988 32190 -27902
rect 32286 -27988 32790 -27902
rect 32886 -27988 33390 -27902
rect 33486 -27988 33990 -27902
rect 34086 -27988 34590 -27902
rect 34686 -27988 35190 -27902
rect 35286 -27988 35790 -27902
rect 35886 -27988 35930 -27902
rect 26160 -28018 35930 -27988
rect 25812 -28466 25924 -28342
rect 26524 -28466 26534 -28166
rect 35546 -28466 35556 -28166
rect 36156 -28342 36162 -26338
rect 36262 -28342 36268 -26338
rect 36156 -28466 36268 -28342
rect 25812 -28472 36268 -28466
rect 25812 -28572 25918 -28472
rect 36162 -28572 36268 -28472
rect 25812 -28578 36268 -28572
<< via1 >>
rect 15532 3904 15914 4204
rect 23666 3904 24344 4204
rect 17600 3640 17696 3726
rect 18180 3640 18276 3726
rect 18780 3640 18876 3726
rect 19380 3640 19476 3726
rect 19980 3640 20076 3726
rect 20580 3640 20676 3726
rect 21180 3640 21276 3726
rect 21780 3640 21876 3726
rect 22380 3640 22476 3726
rect 21514 3388 21574 3448
rect 18078 2708 18138 2768
rect 26114 3904 26714 4204
rect 30746 3904 31346 4204
rect 26362 3640 26458 3726
rect 26942 3640 27038 3726
rect 27542 3640 27638 3726
rect 28142 3640 28238 3726
rect 28742 3640 28838 3726
rect 29342 3640 29438 3726
rect 29942 3640 30038 3726
rect 30542 3640 30638 3726
rect 31142 3640 31238 3726
rect 27066 2834 27126 2894
rect 27528 2834 27588 2894
rect 27982 2836 28042 2896
rect 28444 2834 28504 2894
rect 28898 2834 28958 2894
rect 29348 2834 29408 2894
rect 29814 2834 29874 2894
rect 30270 2834 30330 2894
rect 30504 2626 30564 2686
rect 30504 2284 30564 2344
rect 16474 1554 16534 1614
rect 16930 1554 16990 1614
rect 17390 1554 17450 1614
rect 17846 1554 17906 1614
rect 18304 1554 18364 1614
rect 18768 1554 18828 1614
rect 19222 1554 19282 1614
rect 16478 -420 16538 -360
rect 16934 -420 16994 -360
rect 17394 -420 17454 -360
rect 17850 -420 17910 -360
rect 19682 1554 19742 1614
rect 19912 1554 19972 1614
rect 20140 1554 20200 1614
rect 18308 -420 18368 -360
rect 18772 -420 18832 -360
rect 20596 1554 20656 1614
rect 21056 1554 21116 1614
rect 21512 1554 21572 1614
rect 21968 1554 22028 1614
rect 19222 -420 19282 -360
rect 19678 -420 19738 -360
rect 20146 -420 20206 -360
rect 20604 -420 20664 -360
rect 22424 1554 22484 1614
rect 22882 1554 22942 1614
rect 21060 -420 21120 -360
rect 21516 -420 21576 -360
rect 23342 1554 23402 1614
rect 21972 -420 22032 -360
rect 22428 -420 22488 -360
rect 22886 -420 22946 -360
rect 23346 -420 23406 -360
rect 15774 -1078 15870 -992
rect 16374 -1078 16470 -992
rect 16974 -1078 17070 -992
rect 17574 -1078 17670 -992
rect 18174 -1078 18270 -992
rect 18774 -1078 18870 -992
rect 19374 -1078 19470 -992
rect 19974 -1078 20070 -992
rect 20574 -1078 20670 -992
rect 21174 -1078 21270 -992
rect 21774 -1078 21870 -992
rect 22374 -1078 22470 -992
rect 22974 -1078 23070 -992
rect 23574 -1078 23670 -992
rect 23994 -1078 24090 -992
rect 15532 -1552 15914 -1252
rect 23666 -1552 24344 -1252
rect 10924 -2434 11524 -2134
rect 20556 -2434 21156 -2134
rect 11776 -2694 11872 -2608
rect 12376 -2694 12472 -2608
rect 12976 -2694 13072 -2608
rect 13576 -2694 13672 -2608
rect 14176 -2694 14272 -2608
rect 14776 -2694 14872 -2608
rect 15376 -2694 15472 -2608
rect 15976 -2694 16072 -2608
rect 16576 -2694 16672 -2608
rect 17176 -2694 17272 -2608
rect 17776 -2694 17872 -2608
rect 18376 -2694 18472 -2608
rect 18976 -2694 19072 -2608
rect 19576 -2694 19672 -2608
rect 19996 -2694 20092 -2608
rect 12480 -3326 12540 -3266
rect 12936 -3326 12996 -3266
rect 13396 -3326 13456 -3266
rect 13852 -3326 13912 -3266
rect 12476 -5300 12536 -5240
rect 14310 -3326 14370 -3266
rect 14774 -3326 14834 -3266
rect 12932 -5300 12992 -5240
rect 13392 -5300 13452 -5240
rect 15224 -3326 15284 -3266
rect 15680 -3326 15740 -3266
rect 16148 -3326 16208 -3266
rect 16606 -3326 16666 -3266
rect 13848 -5300 13908 -5240
rect 14306 -5300 14366 -5240
rect 14770 -5300 14830 -5240
rect 15224 -5300 15284 -5240
rect 17062 -3326 17122 -3266
rect 17518 -3326 17578 -3266
rect 15682 -5244 15742 -5240
rect 15682 -5292 15688 -5244
rect 15688 -5292 15736 -5244
rect 15736 -5292 15742 -5244
rect 15682 -5300 15742 -5292
rect 15916 -5288 15976 -5228
rect 16142 -5298 16202 -5240
rect 16142 -5300 16202 -5298
rect 17974 -3326 18034 -3266
rect 18430 -3326 18490 -3266
rect 16598 -5300 16658 -5240
rect 17058 -5300 17118 -5240
rect 18888 -3326 18948 -3266
rect 19348 -3326 19408 -3266
rect 17514 -5300 17574 -5240
rect 17970 -5300 18030 -5240
rect 18426 -5300 18486 -5240
rect 18884 -5300 18944 -5240
rect 19344 -5300 19404 -5240
rect 11690 -5886 11750 -5826
rect 15124 -5988 15184 -5928
rect 11914 -7564 11974 -7504
rect 12376 -7564 12436 -7504
rect 12830 -7560 12890 -7500
rect 13292 -7560 13352 -7500
rect 13746 -7566 13806 -7506
rect 14196 -7560 14256 -7500
rect 14662 -7560 14722 -7500
rect 15118 -7564 15178 -7504
rect 15352 -7686 15412 -7626
rect 16916 -7564 16976 -7504
rect 17378 -7556 17438 -7496
rect 17832 -7562 17892 -7502
rect 18294 -7562 18354 -7502
rect 18748 -7562 18808 -7502
rect 19198 -7556 19258 -7496
rect 19664 -7562 19724 -7502
rect 20120 -7562 20180 -7502
rect 20352 -7692 20412 -7632
rect 25546 2140 25606 2200
rect 25406 -420 25466 -360
rect 25408 -3326 25468 -3266
rect 25234 -5724 25294 -5664
rect 15352 -8366 15412 -8306
rect 11914 -8500 11974 -8440
rect 12376 -8494 12436 -8434
rect 12830 -8500 12890 -8440
rect 13292 -8494 13352 -8434
rect 13746 -8494 13806 -8434
rect 14196 -8494 14256 -8434
rect 14662 -8500 14722 -8440
rect 15118 -8494 15178 -8434
rect 15116 -9710 15176 -9650
rect 20352 -8354 20412 -8294
rect 16916 -8494 16976 -8434
rect 17378 -8496 17438 -8436
rect 17832 -8496 17892 -8436
rect 18294 -8496 18354 -8436
rect 18748 -8496 18808 -8436
rect 19198 -8490 19258 -8430
rect 19664 -8494 19724 -8434
rect 20120 -8494 20180 -8434
rect 11210 -9988 11306 -9902
rect 11790 -9988 11886 -9902
rect 12390 -9988 12486 -9902
rect 12990 -9988 13086 -9902
rect 13590 -9988 13686 -9902
rect 14190 -9988 14286 -9902
rect 14790 -9988 14886 -9902
rect 15390 -9988 15486 -9902
rect 15990 -9988 16086 -9902
rect 16590 -9988 16686 -9902
rect 17190 -9988 17286 -9902
rect 17790 -9988 17886 -9902
rect 18390 -9988 18486 -9902
rect 18990 -9988 19086 -9902
rect 19590 -9988 19686 -9902
rect 20190 -9988 20286 -9902
rect 20790 -9988 20886 -9902
rect 10924 -10466 11524 -10166
rect 20556 -10466 21156 -10166
rect 14878 -11438 15478 -11138
rect 24510 -11438 25110 -11138
rect 15148 -11702 15244 -11616
rect 15748 -11702 15844 -11616
rect 16348 -11702 16444 -11616
rect 16948 -11702 17044 -11616
rect 17548 -11702 17644 -11616
rect 18148 -11702 18244 -11616
rect 18748 -11702 18844 -11616
rect 19348 -11702 19444 -11616
rect 19948 -11702 20044 -11616
rect 20548 -11702 20644 -11616
rect 21148 -11702 21244 -11616
rect 21748 -11702 21844 -11616
rect 22348 -11702 22444 -11616
rect 22948 -11702 23044 -11616
rect 23548 -11702 23644 -11616
rect 24148 -11702 24244 -11616
rect 24728 -11702 24824 -11616
rect 15854 -13170 15914 -13110
rect 16310 -13170 16370 -13110
rect 16776 -13174 16836 -13114
rect 17226 -13168 17286 -13108
rect 17680 -13168 17740 -13108
rect 18142 -13168 18202 -13108
rect 18596 -13168 18656 -13108
rect 19058 -13170 19118 -13110
rect 15622 -13310 15682 -13250
rect 24062 -11954 24122 -11894
rect 20856 -13170 20916 -13110
rect 21312 -13164 21372 -13104
rect 21778 -13170 21838 -13110
rect 22228 -13170 22288 -13110
rect 22682 -13170 22742 -13110
rect 23144 -13164 23204 -13104
rect 23598 -13170 23658 -13110
rect 24060 -13164 24120 -13104
rect 20622 -13298 20682 -13238
rect 15622 -13972 15682 -13912
rect 15854 -14102 15914 -14042
rect 16310 -14102 16370 -14042
rect 16776 -14108 16836 -14048
rect 17226 -14102 17286 -14042
rect 17680 -14102 17740 -14042
rect 18142 -14102 18202 -14042
rect 18596 -14108 18656 -14048
rect 19058 -14100 19118 -14040
rect 20622 -13978 20682 -13918
rect 20856 -14100 20916 -14040
rect 21312 -14104 21372 -14044
rect 21778 -14104 21838 -14044
rect 22228 -14098 22288 -14038
rect 22682 -14104 22742 -14044
rect 23144 -14104 23204 -14044
rect 23598 -14100 23658 -14040
rect 24060 -14100 24120 -14040
rect 24284 -15778 24344 -15718
rect 16630 -16364 16690 -16304
rect 17090 -16364 17150 -16304
rect 17548 -16364 17608 -16304
rect 18004 -16364 18064 -16304
rect 18460 -16364 18520 -16304
rect 16626 -18338 16686 -18278
rect 17086 -18338 17146 -18278
rect 18916 -16364 18976 -16304
rect 19376 -16364 19436 -16304
rect 17544 -18338 17604 -18278
rect 18000 -18338 18060 -18278
rect 19832 -16306 19892 -16304
rect 19832 -16364 19892 -16306
rect 20058 -16376 20118 -16316
rect 20292 -16312 20352 -16304
rect 20292 -16360 20298 -16312
rect 20298 -16360 20346 -16312
rect 20346 -16360 20352 -16312
rect 20292 -16364 20352 -16360
rect 18456 -18338 18516 -18278
rect 18912 -18338 18972 -18278
rect 20750 -16364 20810 -16304
rect 21204 -16364 21264 -16304
rect 21668 -16364 21728 -16304
rect 22126 -16364 22186 -16304
rect 19368 -18338 19428 -18278
rect 19826 -18338 19886 -18278
rect 20294 -18338 20354 -18278
rect 20750 -18338 20810 -18278
rect 22582 -16364 22642 -16304
rect 23042 -16364 23102 -16304
rect 21200 -18338 21260 -18278
rect 21664 -18338 21724 -18278
rect 23498 -16364 23558 -16304
rect 22122 -18338 22182 -18278
rect 22578 -18338 22638 -18278
rect 23038 -18338 23098 -18278
rect 23494 -18338 23554 -18278
rect 15942 -18996 16038 -18910
rect 16362 -18996 16458 -18910
rect 16962 -18996 17058 -18910
rect 17562 -18996 17658 -18910
rect 18162 -18996 18258 -18910
rect 18762 -18996 18858 -18910
rect 19362 -18996 19458 -18910
rect 19962 -18996 20058 -18910
rect 20562 -18996 20658 -18910
rect 21162 -18996 21258 -18910
rect 21762 -18996 21858 -18910
rect 22362 -18996 22458 -18910
rect 22962 -18996 23058 -18910
rect 23562 -18996 23658 -18910
rect 24162 -18996 24258 -18910
rect 14878 -19470 15478 -19170
rect 24510 -19470 25110 -19170
rect 27066 1966 27126 2026
rect 27528 1966 27588 2026
rect 27982 1966 28042 2026
rect 28444 1966 28504 2026
rect 28898 1966 28958 2026
rect 29348 1966 29408 2026
rect 29814 1966 29874 2026
rect 30270 1966 30330 2026
rect 30504 1972 30564 2032
rect 30278 394 30338 454
rect 26290 -1078 26386 -992
rect 26890 -1078 26986 -992
rect 27490 -1078 27586 -992
rect 28090 -1078 28186 -992
rect 28690 -1078 28786 -992
rect 29290 -1078 29386 -992
rect 29890 -1078 29986 -992
rect 30490 -1078 30586 -992
rect 31090 -1078 31186 -992
rect 26114 -1552 26714 -1252
rect 30746 -1552 31346 -1252
rect 25924 -2434 26524 -2134
rect 35556 -2434 36156 -2134
rect 26776 -2694 26872 -2608
rect 27376 -2694 27472 -2608
rect 27976 -2694 28072 -2608
rect 28576 -2694 28672 -2608
rect 29176 -2694 29272 -2608
rect 29776 -2694 29872 -2608
rect 30376 -2694 30472 -2608
rect 30976 -2694 31072 -2608
rect 31576 -2694 31672 -2608
rect 32176 -2694 32272 -2608
rect 32776 -2694 32872 -2608
rect 33376 -2694 33472 -2608
rect 33976 -2694 34072 -2608
rect 34576 -2694 34672 -2608
rect 34996 -2694 35092 -2608
rect 27480 -3326 27540 -3266
rect 27936 -3326 27996 -3266
rect 28396 -3326 28456 -3266
rect 28852 -3326 28912 -3266
rect 27476 -5300 27536 -5240
rect 29310 -3326 29370 -3266
rect 29774 -3326 29834 -3266
rect 27932 -5300 27992 -5240
rect 28392 -5300 28452 -5240
rect 30224 -3326 30284 -3266
rect 30680 -3326 30740 -3266
rect 31148 -3326 31208 -3266
rect 31606 -3326 31666 -3266
rect 28848 -5300 28908 -5240
rect 29306 -5300 29366 -5240
rect 29770 -5300 29830 -5240
rect 30224 -5300 30284 -5240
rect 32062 -3326 32122 -3266
rect 32518 -3326 32578 -3266
rect 30682 -5244 30742 -5240
rect 30682 -5292 30688 -5244
rect 30688 -5292 30736 -5244
rect 30736 -5292 30742 -5244
rect 30682 -5300 30742 -5292
rect 30916 -5288 30976 -5228
rect 31142 -5298 31202 -5240
rect 31142 -5300 31202 -5298
rect 32974 -3326 33034 -3266
rect 33430 -3326 33490 -3266
rect 31598 -5300 31658 -5240
rect 32058 -5300 32118 -5240
rect 33888 -3326 33948 -3266
rect 34348 -3326 34408 -3266
rect 32514 -5300 32574 -5240
rect 32970 -5300 33030 -5240
rect 33426 -5300 33486 -5240
rect 33884 -5300 33944 -5240
rect 34344 -5300 34404 -5240
rect 26690 -5886 26750 -5826
rect 26914 -7564 26974 -7504
rect 27376 -7564 27436 -7504
rect 27830 -7560 27890 -7500
rect 28292 -7560 28352 -7500
rect 28746 -7566 28806 -7506
rect 29196 -7560 29256 -7500
rect 29662 -7560 29722 -7500
rect 30118 -7564 30178 -7504
rect 30352 -7686 30412 -7626
rect 31916 -7564 31976 -7504
rect 32378 -7556 32438 -7496
rect 32832 -7562 32892 -7502
rect 33294 -7562 33354 -7502
rect 33748 -7562 33808 -7502
rect 34198 -7556 34258 -7496
rect 34664 -7562 34724 -7502
rect 35120 -7562 35180 -7502
rect 35352 -7692 35412 -7632
rect 25546 -9710 25606 -9650
rect 25406 -16364 25466 -16304
rect 10924 -20434 11524 -20134
rect 20556 -20434 21156 -20134
rect 11776 -20694 11872 -20608
rect 12376 -20694 12472 -20608
rect 12976 -20694 13072 -20608
rect 13576 -20694 13672 -20608
rect 14176 -20694 14272 -20608
rect 14776 -20694 14872 -20608
rect 15376 -20694 15472 -20608
rect 15976 -20694 16072 -20608
rect 16576 -20694 16672 -20608
rect 17176 -20694 17272 -20608
rect 17776 -20694 17872 -20608
rect 18376 -20694 18472 -20608
rect 18976 -20694 19072 -20608
rect 19576 -20694 19672 -20608
rect 19996 -20694 20092 -20608
rect 12480 -21326 12540 -21266
rect 12936 -21326 12996 -21266
rect 13396 -21326 13456 -21266
rect 13852 -21326 13912 -21266
rect 12476 -23300 12536 -23240
rect 14310 -21326 14370 -21266
rect 14774 -21326 14834 -21266
rect 12932 -23300 12992 -23240
rect 13392 -23300 13452 -23240
rect 15224 -21326 15284 -21266
rect 15680 -21326 15740 -21266
rect 16148 -21326 16208 -21266
rect 16606 -21326 16666 -21266
rect 13848 -23300 13908 -23240
rect 14306 -23300 14366 -23240
rect 14770 -23300 14830 -23240
rect 15224 -23300 15284 -23240
rect 17062 -21326 17122 -21266
rect 17518 -21326 17578 -21266
rect 15682 -23244 15742 -23240
rect 15682 -23292 15688 -23244
rect 15688 -23292 15736 -23244
rect 15736 -23292 15742 -23244
rect 15682 -23300 15742 -23292
rect 15916 -23288 15976 -23228
rect 16142 -23298 16202 -23240
rect 16142 -23300 16202 -23298
rect 17974 -21326 18034 -21266
rect 18430 -21326 18490 -21266
rect 16598 -23300 16658 -23240
rect 17058 -23300 17118 -23240
rect 18888 -21326 18948 -21266
rect 19348 -21326 19408 -21266
rect 17514 -23300 17574 -23240
rect 17970 -23300 18030 -23240
rect 18426 -23300 18486 -23240
rect 18884 -23300 18944 -23240
rect 19344 -23300 19404 -23240
rect 11690 -23886 11750 -23826
rect 11914 -25564 11974 -25504
rect 12376 -25564 12436 -25504
rect 12830 -25560 12890 -25500
rect 13292 -25560 13352 -25500
rect 13746 -25566 13806 -25506
rect 14196 -25560 14256 -25500
rect 14662 -25560 14722 -25500
rect 15118 -25564 15178 -25504
rect 15352 -25686 15412 -25626
rect 16916 -25564 16976 -25504
rect 17378 -25556 17438 -25496
rect 17832 -25562 17892 -25502
rect 18294 -25562 18354 -25502
rect 18748 -25562 18808 -25502
rect 19198 -25556 19258 -25496
rect 19664 -25562 19724 -25502
rect 20120 -25562 20180 -25502
rect 20352 -25692 20412 -25632
rect 30352 -8366 30412 -8306
rect 26914 -8500 26974 -8440
rect 27376 -8494 27436 -8434
rect 27830 -8500 27890 -8440
rect 28292 -8494 28352 -8434
rect 28746 -8494 28806 -8434
rect 29196 -8494 29256 -8434
rect 29662 -8500 29722 -8440
rect 30118 -8494 30178 -8434
rect 26914 -9710 26974 -9650
rect 35352 -8354 35412 -8294
rect 31916 -8494 31976 -8434
rect 32378 -8496 32438 -8436
rect 32832 -8496 32892 -8436
rect 33294 -8496 33354 -8436
rect 33748 -8496 33808 -8436
rect 34198 -8490 34258 -8430
rect 34664 -8494 34724 -8434
rect 35120 -8494 35180 -8434
rect 26210 -9988 26306 -9902
rect 26790 -9988 26886 -9902
rect 27390 -9988 27486 -9902
rect 27990 -9988 28086 -9902
rect 28590 -9988 28686 -9902
rect 29190 -9988 29286 -9902
rect 29790 -9988 29886 -9902
rect 30390 -9988 30486 -9902
rect 30990 -9988 31086 -9902
rect 31590 -9988 31686 -9902
rect 32190 -9988 32286 -9902
rect 32790 -9988 32886 -9902
rect 33390 -9988 33486 -9902
rect 33990 -9988 34086 -9902
rect 34590 -9988 34686 -9902
rect 35190 -9988 35286 -9902
rect 35790 -9988 35886 -9902
rect 25924 -10466 26524 -10166
rect 35556 -10466 36156 -10166
rect 25546 -11954 25606 -11894
rect 25406 -23300 25466 -23240
rect 15352 -26366 15412 -26306
rect 11914 -26500 11974 -26440
rect 12376 -26494 12436 -26434
rect 12830 -26500 12890 -26440
rect 13292 -26494 13352 -26434
rect 13746 -26494 13806 -26434
rect 14196 -26494 14256 -26434
rect 14662 -26500 14722 -26440
rect 15118 -26494 15178 -26434
rect 15118 -27710 15178 -27650
rect 20352 -26354 20412 -26294
rect 16916 -26494 16976 -26434
rect 17378 -26496 17438 -26436
rect 17832 -26496 17892 -26436
rect 18294 -26496 18354 -26436
rect 18748 -26496 18808 -26436
rect 19198 -26490 19258 -26430
rect 19664 -26494 19724 -26434
rect 20120 -26494 20180 -26434
rect 11210 -27988 11306 -27902
rect 11790 -27988 11886 -27902
rect 12390 -27988 12486 -27902
rect 12990 -27988 13086 -27902
rect 13590 -27988 13686 -27902
rect 14190 -27988 14286 -27902
rect 14790 -27988 14886 -27902
rect 15390 -27988 15486 -27902
rect 15990 -27988 16086 -27902
rect 16590 -27988 16686 -27902
rect 17190 -27988 17286 -27902
rect 17790 -27988 17886 -27902
rect 18390 -27988 18486 -27902
rect 18990 -27988 19086 -27902
rect 19590 -27988 19686 -27902
rect 20190 -27988 20286 -27902
rect 20790 -27988 20886 -27902
rect 10924 -28466 11524 -28166
rect 20556 -28466 21156 -28166
rect 29878 -11438 30478 -11138
rect 39510 -11438 40110 -11138
rect 30148 -11702 30244 -11616
rect 30748 -11702 30844 -11616
rect 31348 -11702 31444 -11616
rect 31948 -11702 32044 -11616
rect 32548 -11702 32644 -11616
rect 33148 -11702 33244 -11616
rect 33748 -11702 33844 -11616
rect 34348 -11702 34444 -11616
rect 34948 -11702 35044 -11616
rect 35548 -11702 35644 -11616
rect 36148 -11702 36244 -11616
rect 36748 -11702 36844 -11616
rect 37348 -11702 37444 -11616
rect 37948 -11702 38044 -11616
rect 38548 -11702 38644 -11616
rect 39148 -11702 39244 -11616
rect 39728 -11702 39824 -11616
rect 30854 -13170 30914 -13110
rect 31310 -13170 31370 -13110
rect 31776 -13174 31836 -13114
rect 32226 -13168 32286 -13108
rect 32680 -13168 32740 -13108
rect 33142 -13168 33202 -13108
rect 33596 -13168 33656 -13108
rect 34058 -13170 34118 -13110
rect 30622 -13310 30682 -13250
rect 35856 -11954 35916 -11894
rect 35856 -13170 35916 -13110
rect 36312 -13164 36372 -13104
rect 36778 -13170 36838 -13110
rect 37228 -13170 37288 -13110
rect 37682 -13170 37742 -13110
rect 38144 -13164 38204 -13104
rect 38598 -13170 38658 -13110
rect 39060 -13164 39120 -13104
rect 35622 -13298 35682 -13238
rect 30622 -13972 30682 -13912
rect 30854 -14102 30914 -14042
rect 31310 -14102 31370 -14042
rect 31776 -14108 31836 -14048
rect 32226 -14102 32286 -14042
rect 32680 -14102 32740 -14042
rect 33142 -14102 33202 -14042
rect 33596 -14108 33656 -14048
rect 34058 -14100 34118 -14040
rect 35622 -13978 35682 -13918
rect 35856 -14100 35916 -14040
rect 36312 -14104 36372 -14044
rect 36778 -14104 36838 -14044
rect 37228 -14098 37288 -14038
rect 37682 -14104 37742 -14044
rect 38144 -14104 38204 -14044
rect 38598 -14100 38658 -14040
rect 39060 -14100 39120 -14040
rect 39284 -15778 39344 -15718
rect 31630 -16364 31690 -16304
rect 32090 -16364 32150 -16304
rect 32548 -16364 32608 -16304
rect 33004 -16364 33064 -16304
rect 33460 -16364 33520 -16304
rect 31626 -18338 31686 -18278
rect 32086 -18338 32146 -18278
rect 33916 -16364 33976 -16304
rect 34376 -16364 34436 -16304
rect 32544 -18338 32604 -18278
rect 33000 -18338 33060 -18278
rect 34832 -16306 34892 -16304
rect 34832 -16364 34892 -16306
rect 35058 -16376 35118 -16316
rect 35292 -16312 35352 -16304
rect 35292 -16360 35298 -16312
rect 35298 -16360 35346 -16312
rect 35346 -16360 35352 -16312
rect 35292 -16364 35352 -16360
rect 33456 -18338 33516 -18278
rect 33912 -18338 33972 -18278
rect 35750 -16364 35810 -16304
rect 36204 -16364 36264 -16304
rect 36668 -16364 36728 -16304
rect 37126 -16364 37186 -16304
rect 34368 -18338 34428 -18278
rect 34826 -18338 34886 -18278
rect 35294 -18338 35354 -18278
rect 35750 -18338 35810 -18278
rect 37582 -16364 37642 -16304
rect 38042 -16364 38102 -16304
rect 36200 -18338 36260 -18278
rect 36664 -18338 36724 -18278
rect 38498 -16364 38558 -16304
rect 37122 -18338 37182 -18278
rect 37578 -18338 37638 -18278
rect 38038 -18338 38098 -18278
rect 38494 -18338 38554 -18278
rect 30942 -18996 31038 -18910
rect 31362 -18996 31458 -18910
rect 31962 -18996 32058 -18910
rect 32562 -18996 32658 -18910
rect 33162 -18996 33258 -18910
rect 33762 -18996 33858 -18910
rect 34362 -18996 34458 -18910
rect 34962 -18996 35058 -18910
rect 35562 -18996 35658 -18910
rect 36162 -18996 36258 -18910
rect 36762 -18996 36858 -18910
rect 37362 -18996 37458 -18910
rect 37962 -18996 38058 -18910
rect 38562 -18996 38658 -18910
rect 39162 -18996 39258 -18910
rect 29878 -19470 30478 -19170
rect 39510 -19470 40110 -19170
rect 25924 -20434 26524 -20134
rect 35556 -20434 36156 -20134
rect 26776 -20694 26872 -20608
rect 27376 -20694 27472 -20608
rect 27976 -20694 28072 -20608
rect 28576 -20694 28672 -20608
rect 29176 -20694 29272 -20608
rect 29776 -20694 29872 -20608
rect 30376 -20694 30472 -20608
rect 30976 -20694 31072 -20608
rect 31576 -20694 31672 -20608
rect 32176 -20694 32272 -20608
rect 32776 -20694 32872 -20608
rect 33376 -20694 33472 -20608
rect 33976 -20694 34072 -20608
rect 34576 -20694 34672 -20608
rect 34996 -20694 35092 -20608
rect 27480 -21326 27540 -21266
rect 27936 -21326 27996 -21266
rect 28396 -21326 28456 -21266
rect 28852 -21326 28912 -21266
rect 27476 -23300 27536 -23240
rect 29310 -21326 29370 -21266
rect 29774 -21326 29834 -21266
rect 27932 -23300 27992 -23240
rect 28392 -23300 28452 -23240
rect 30224 -21326 30284 -21266
rect 30680 -21326 30740 -21266
rect 31148 -21326 31208 -21266
rect 31606 -21326 31666 -21266
rect 28848 -23300 28908 -23240
rect 29306 -23300 29366 -23240
rect 29770 -23300 29830 -23240
rect 30224 -23300 30284 -23240
rect 32062 -21326 32122 -21266
rect 32518 -21326 32578 -21266
rect 30682 -23244 30742 -23240
rect 30682 -23292 30688 -23244
rect 30688 -23292 30736 -23244
rect 30736 -23292 30742 -23244
rect 30682 -23300 30742 -23292
rect 30916 -23288 30976 -23228
rect 31142 -23298 31202 -23240
rect 31142 -23300 31202 -23298
rect 32974 -21326 33034 -21266
rect 33430 -21326 33490 -21266
rect 31598 -23300 31658 -23240
rect 32058 -23300 32118 -23240
rect 33888 -21326 33948 -21266
rect 34348 -21326 34408 -21266
rect 32514 -23300 32574 -23240
rect 32970 -23300 33030 -23240
rect 33426 -23300 33486 -23240
rect 33884 -23300 33944 -23240
rect 34344 -23300 34404 -23240
rect 26690 -23886 26750 -23826
rect 26914 -25564 26974 -25504
rect 27376 -25564 27436 -25504
rect 27830 -25560 27890 -25500
rect 28292 -25560 28352 -25500
rect 28746 -25566 28806 -25506
rect 29196 -25560 29256 -25500
rect 29662 -25560 29722 -25500
rect 30118 -25564 30178 -25504
rect 30352 -25686 30412 -25626
rect 31916 -25564 31976 -25504
rect 32378 -25556 32438 -25496
rect 32832 -25562 32892 -25502
rect 33294 -25562 33354 -25502
rect 33748 -25562 33808 -25502
rect 34198 -25556 34258 -25496
rect 34664 -25562 34724 -25502
rect 35120 -25562 35180 -25502
rect 35352 -25692 35412 -25632
rect 25546 -27710 25606 -27650
rect 30352 -26366 30412 -26306
rect 26914 -26500 26974 -26440
rect 27376 -26494 27436 -26434
rect 27830 -26500 27890 -26440
rect 28292 -26494 28352 -26434
rect 28746 -26494 28806 -26434
rect 29196 -26494 29256 -26434
rect 29662 -26500 29722 -26440
rect 30118 -26494 30178 -26434
rect 26914 -27710 26974 -27650
rect 35352 -26354 35412 -26294
rect 31916 -26494 31976 -26434
rect 32378 -26496 32438 -26436
rect 32832 -26496 32892 -26436
rect 33294 -26496 33354 -26436
rect 33748 -26496 33808 -26436
rect 34198 -26490 34258 -26430
rect 34664 -26494 34724 -26434
rect 35120 -26494 35180 -26434
rect 26210 -27988 26306 -27902
rect 26790 -27988 26886 -27902
rect 27390 -27988 27486 -27902
rect 27990 -27988 28086 -27902
rect 28590 -27988 28686 -27902
rect 29190 -27988 29286 -27902
rect 29790 -27988 29886 -27902
rect 30390 -27988 30486 -27902
rect 30990 -27988 31086 -27902
rect 31590 -27988 31686 -27902
rect 32190 -27988 32286 -27902
rect 32790 -27988 32886 -27902
rect 33390 -27988 33486 -27902
rect 33990 -27988 34086 -27902
rect 34590 -27988 34686 -27902
rect 35190 -27988 35286 -27902
rect 35790 -27988 35886 -27902
rect 25924 -28466 26524 -28166
rect 35556 -28466 36156 -28166
<< metal2 >>
rect 15532 4204 15914 4214
rect 15532 3894 15914 3904
rect 23666 4204 24344 4214
rect 23666 3894 24344 3904
rect 26114 4204 26714 4214
rect 26114 3894 26714 3904
rect 30746 4204 31346 4214
rect 30746 3894 31346 3904
rect 17550 3726 22522 3756
rect 17550 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 22522 3726
rect 17550 3612 22522 3640
rect 26312 3726 31284 3756
rect 26312 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 31284 3726
rect 26312 3612 31284 3640
rect 21514 3448 21574 3454
rect 21574 3388 25606 3448
rect 21514 3382 21574 3388
rect 18072 2708 18078 2768
rect 18138 2708 18144 2768
rect 16474 1614 16534 1620
rect 16930 1614 16990 1620
rect 17390 1614 17450 1620
rect 17846 1614 17906 1620
rect 18078 1614 18138 2708
rect 25546 2200 25606 3388
rect 27066 2894 27126 2900
rect 25540 2140 25546 2200
rect 25606 2140 25612 2200
rect 27066 2026 27126 2834
rect 27066 1960 27126 1966
rect 27528 2894 27588 2900
rect 27528 2026 27588 2834
rect 27982 2896 28042 2902
rect 27982 2026 28042 2836
rect 28444 2894 28504 2900
rect 28444 2026 28504 2834
rect 28898 2894 28958 2900
rect 28898 2026 28958 2834
rect 29348 2894 29408 2900
rect 29348 2026 29408 2834
rect 29814 2894 29874 2900
rect 29814 2026 29874 2834
rect 30270 2894 30330 2900
rect 30270 2026 30330 2834
rect 30504 2686 30564 2692
rect 30504 2344 30564 2626
rect 30498 2284 30504 2344
rect 30564 2284 30570 2344
rect 30504 2032 30564 2284
rect 27976 1966 27982 2026
rect 28042 1966 28048 2026
rect 28438 1966 28444 2026
rect 28504 1966 28510 2026
rect 29342 1966 29348 2026
rect 29408 1966 29414 2026
rect 29808 1966 29814 2026
rect 29874 1966 29880 2026
rect 30498 1972 30504 2032
rect 30564 1972 30570 2032
rect 27528 1960 27588 1966
rect 28898 1960 28958 1966
rect 30270 1960 30330 1966
rect 18304 1614 18364 1620
rect 18768 1614 18828 1620
rect 19222 1614 19282 1620
rect 19682 1614 19742 1620
rect 19912 1614 19972 1620
rect 20140 1614 20200 1620
rect 20596 1614 20656 1620
rect 21056 1614 21116 1620
rect 21512 1614 21572 1620
rect 21968 1614 22028 1620
rect 22424 1614 22484 1620
rect 22882 1614 22942 1620
rect 23342 1614 23402 1620
rect 16534 1554 16930 1614
rect 16990 1554 17390 1614
rect 17450 1554 17846 1614
rect 17906 1554 18304 1614
rect 18364 1554 18768 1614
rect 18828 1554 19222 1614
rect 19282 1554 19682 1614
rect 19742 1554 19912 1614
rect 19972 1554 20140 1614
rect 20200 1554 20596 1614
rect 20656 1554 21056 1614
rect 21116 1554 21512 1614
rect 21572 1554 21968 1614
rect 22028 1554 22424 1614
rect 22484 1554 22882 1614
rect 22942 1554 23342 1614
rect 16474 1548 16534 1554
rect 16930 1548 16990 1554
rect 17390 1548 17450 1554
rect 17846 1548 17906 1554
rect 18304 1548 18364 1554
rect 18768 1548 18828 1554
rect 19222 1548 19282 1554
rect 19682 1548 19742 1554
rect 19912 1548 19972 1554
rect 20140 1548 20200 1554
rect 20596 1548 20656 1554
rect 21056 1548 21116 1554
rect 21512 1548 21572 1554
rect 21968 1548 22028 1554
rect 22424 1548 22484 1554
rect 22882 1548 22942 1554
rect 23342 1548 23402 1554
rect 30278 454 30338 460
rect 30338 394 31902 454
rect 30278 388 30338 394
rect 16478 -360 16538 -354
rect 16934 -360 16994 -354
rect 17394 -360 17454 -354
rect 17850 -360 17910 -354
rect 18308 -360 18368 -354
rect 18772 -360 18832 -354
rect 19222 -360 19282 -354
rect 19678 -360 19738 -354
rect 20146 -360 20206 -354
rect 20604 -360 20664 -354
rect 21060 -360 21120 -354
rect 21516 -360 21576 -354
rect 21972 -360 22032 -354
rect 22428 -360 22488 -354
rect 22886 -360 22946 -354
rect 23346 -360 23406 -354
rect 25406 -360 25466 -354
rect 16538 -420 16934 -360
rect 16994 -420 17394 -360
rect 17454 -420 17850 -360
rect 17910 -420 18308 -360
rect 18368 -420 18772 -360
rect 18832 -420 19222 -360
rect 19282 -420 19678 -360
rect 19738 -420 20146 -360
rect 20206 -420 20604 -360
rect 20664 -420 21060 -360
rect 21120 -420 21516 -360
rect 21576 -420 21972 -360
rect 22032 -420 22428 -360
rect 22488 -420 22886 -360
rect 22946 -420 23346 -360
rect 23406 -420 25406 -360
rect 16478 -426 16538 -420
rect 16934 -426 16994 -420
rect 17394 -426 17454 -420
rect 17850 -426 17910 -420
rect 18308 -426 18368 -420
rect 18772 -426 18832 -420
rect 19222 -426 19282 -420
rect 19678 -426 19738 -420
rect 20146 -426 20206 -420
rect 20604 -426 20664 -420
rect 21060 -426 21120 -420
rect 21516 -426 21576 -420
rect 21972 -426 22032 -420
rect 22428 -426 22488 -420
rect 22886 -426 22946 -420
rect 23346 -426 23406 -420
rect 25406 -426 25466 -420
rect 31802 -678 31902 394
rect 31802 -778 36438 -678
rect 15760 -992 24116 -982
rect 15760 -1078 15774 -992
rect 15870 -1078 16374 -992
rect 16470 -1078 16974 -992
rect 17070 -1078 17574 -992
rect 17670 -1078 18174 -992
rect 18270 -1078 18774 -992
rect 18870 -1078 19374 -992
rect 19470 -1078 19974 -992
rect 20070 -1078 20574 -992
rect 20670 -1078 21174 -992
rect 21270 -1078 21774 -992
rect 21870 -1078 22374 -992
rect 22470 -1078 22974 -992
rect 23070 -1078 23574 -992
rect 23670 -1078 23994 -992
rect 24090 -1078 24116 -992
rect 15760 -1092 24116 -1078
rect 26276 -992 31274 -982
rect 26276 -1078 26290 -992
rect 26386 -1078 26890 -992
rect 26986 -1078 27490 -992
rect 27586 -1078 28090 -992
rect 28186 -1078 28690 -992
rect 28786 -1078 29290 -992
rect 29386 -1078 29890 -992
rect 29986 -1078 30490 -992
rect 30586 -1078 31090 -992
rect 31186 -1078 31274 -992
rect 26276 -1092 31274 -1078
rect 15532 -1252 15914 -1242
rect 15532 -1562 15914 -1552
rect 23666 -1252 24344 -1242
rect 23666 -1562 24344 -1552
rect 26114 -1252 26714 -1242
rect 26114 -1562 26714 -1552
rect 30746 -1252 31346 -1242
rect 30746 -1562 31346 -1552
rect 10924 -2134 11524 -2124
rect 10924 -2444 11524 -2434
rect 20556 -2134 21156 -2124
rect 20556 -2444 21156 -2434
rect 25924 -2134 26524 -2124
rect 25924 -2444 26524 -2434
rect 35556 -2134 36156 -2124
rect 35556 -2444 36156 -2434
rect 11762 -2608 20118 -2594
rect 11762 -2694 11776 -2608
rect 11872 -2694 12376 -2608
rect 12472 -2694 12976 -2608
rect 13072 -2694 13576 -2608
rect 13672 -2694 14176 -2608
rect 14272 -2694 14776 -2608
rect 14872 -2694 15376 -2608
rect 15472 -2694 15976 -2608
rect 16072 -2694 16576 -2608
rect 16672 -2694 17176 -2608
rect 17272 -2694 17776 -2608
rect 17872 -2694 18376 -2608
rect 18472 -2694 18976 -2608
rect 19072 -2694 19576 -2608
rect 19672 -2694 19996 -2608
rect 20092 -2694 20118 -2608
rect 11762 -2704 20118 -2694
rect 26762 -2608 35118 -2594
rect 26762 -2694 26776 -2608
rect 26872 -2694 27376 -2608
rect 27472 -2694 27976 -2608
rect 28072 -2694 28576 -2608
rect 28672 -2694 29176 -2608
rect 29272 -2694 29776 -2608
rect 29872 -2694 30376 -2608
rect 30472 -2694 30976 -2608
rect 31072 -2694 31576 -2608
rect 31672 -2694 32176 -2608
rect 32272 -2694 32776 -2608
rect 32872 -2694 33376 -2608
rect 33472 -2694 33976 -2608
rect 34072 -2694 34576 -2608
rect 34672 -2694 34996 -2608
rect 35092 -2694 35118 -2608
rect 26762 -2704 35118 -2694
rect 12480 -3266 12540 -3260
rect 12936 -3266 12996 -3260
rect 13396 -3266 13456 -3260
rect 13852 -3266 13912 -3260
rect 14310 -3266 14370 -3260
rect 14774 -3266 14834 -3260
rect 15224 -3266 15284 -3260
rect 15680 -3266 15740 -3260
rect 16148 -3266 16208 -3260
rect 16606 -3266 16666 -3260
rect 17062 -3266 17122 -3260
rect 17518 -3266 17578 -3260
rect 17974 -3266 18034 -3260
rect 18430 -3266 18490 -3260
rect 18888 -3266 18948 -3260
rect 19348 -3266 19408 -3260
rect 27480 -3266 27540 -3260
rect 27936 -3266 27996 -3260
rect 28396 -3266 28456 -3260
rect 28852 -3266 28912 -3260
rect 29310 -3266 29370 -3260
rect 29774 -3266 29834 -3260
rect 30224 -3266 30284 -3260
rect 30680 -3266 30740 -3260
rect 31148 -3266 31208 -3260
rect 31606 -3266 31666 -3260
rect 32062 -3266 32122 -3260
rect 32518 -3266 32578 -3260
rect 32974 -3266 33034 -3260
rect 33430 -3266 33490 -3260
rect 33888 -3266 33948 -3260
rect 34348 -3266 34408 -3260
rect 12540 -3326 12936 -3266
rect 12996 -3326 13396 -3266
rect 13456 -3326 13852 -3266
rect 13912 -3326 14310 -3266
rect 14370 -3326 14774 -3266
rect 14834 -3326 15224 -3266
rect 15284 -3326 15680 -3266
rect 15740 -3326 16148 -3266
rect 16208 -3326 16606 -3266
rect 16666 -3326 17062 -3266
rect 17122 -3326 17518 -3266
rect 17578 -3326 17974 -3266
rect 18034 -3326 18430 -3266
rect 18490 -3326 18888 -3266
rect 18948 -3326 19348 -3266
rect 19408 -3326 25408 -3266
rect 25468 -3326 27480 -3266
rect 27540 -3326 27936 -3266
rect 27996 -3326 28396 -3266
rect 28456 -3326 28852 -3266
rect 28912 -3326 29310 -3266
rect 29370 -3326 29774 -3266
rect 29834 -3326 30224 -3266
rect 30284 -3326 30680 -3266
rect 30740 -3326 31148 -3266
rect 31208 -3326 31606 -3266
rect 31666 -3326 32062 -3266
rect 32122 -3326 32518 -3266
rect 32578 -3326 32974 -3266
rect 33034 -3326 33430 -3266
rect 33490 -3326 33888 -3266
rect 33948 -3326 34348 -3266
rect 12480 -3332 12540 -3326
rect 12936 -3332 12996 -3326
rect 13396 -3332 13456 -3326
rect 13852 -3332 13912 -3326
rect 14310 -3332 14370 -3326
rect 14774 -3332 14834 -3326
rect 15224 -3332 15284 -3326
rect 15680 -3332 15740 -3326
rect 16148 -3332 16208 -3326
rect 16606 -3332 16666 -3326
rect 17062 -3332 17122 -3326
rect 17518 -3332 17578 -3326
rect 17974 -3332 18034 -3326
rect 18430 -3332 18490 -3326
rect 18888 -3332 18948 -3326
rect 19348 -3332 19408 -3326
rect 27480 -3332 27540 -3326
rect 27936 -3332 27996 -3326
rect 28396 -3332 28456 -3326
rect 28852 -3332 28912 -3326
rect 29310 -3332 29370 -3326
rect 29774 -3332 29834 -3326
rect 30224 -3332 30284 -3326
rect 30680 -3332 30740 -3326
rect 31148 -3332 31208 -3326
rect 31606 -3332 31666 -3326
rect 32062 -3332 32122 -3326
rect 32518 -3332 32578 -3326
rect 32974 -3332 33034 -3326
rect 33430 -3332 33490 -3326
rect 33888 -3332 33948 -3326
rect 34348 -3332 34408 -3326
rect 12476 -5240 12536 -5234
rect 12932 -5240 12992 -5234
rect 13392 -5240 13452 -5234
rect 13848 -5240 13908 -5234
rect 14306 -5240 14366 -5234
rect 14770 -5240 14830 -5234
rect 15224 -5240 15284 -5234
rect 15682 -5240 15742 -5234
rect 12536 -5300 12932 -5240
rect 12992 -5300 13392 -5240
rect 13452 -5300 13848 -5240
rect 13908 -5300 14306 -5240
rect 14366 -5300 14770 -5240
rect 14830 -5300 15224 -5240
rect 15284 -5300 15682 -5240
rect 15910 -5288 15916 -5228
rect 15976 -5288 15982 -5228
rect 16142 -5240 16202 -5234
rect 16598 -5240 16658 -5234
rect 17058 -5240 17118 -5234
rect 17514 -5240 17574 -5234
rect 17970 -5240 18030 -5234
rect 18426 -5240 18486 -5234
rect 18884 -5240 18944 -5234
rect 19344 -5240 19404 -5234
rect 12476 -5306 12536 -5300
rect 12932 -5306 12992 -5300
rect 13392 -5306 13452 -5300
rect 13848 -5306 13908 -5300
rect 14306 -5306 14366 -5300
rect 14770 -5306 14830 -5300
rect 15224 -5306 15284 -5300
rect 15682 -5306 15742 -5300
rect 11690 -5826 11750 -5820
rect 15916 -5826 15976 -5288
rect 16202 -5300 16598 -5240
rect 16658 -5300 17058 -5240
rect 17118 -5300 17514 -5240
rect 17574 -5300 17970 -5240
rect 18030 -5300 18426 -5240
rect 18486 -5300 18884 -5240
rect 18944 -5300 19344 -5240
rect 16142 -5306 16202 -5300
rect 16598 -5306 16658 -5300
rect 17058 -5306 17118 -5300
rect 17514 -5306 17574 -5300
rect 17970 -5306 18030 -5300
rect 18426 -5306 18486 -5300
rect 18884 -5306 18944 -5300
rect 19344 -5306 19404 -5300
rect 27476 -5240 27536 -5234
rect 27932 -5240 27992 -5234
rect 28392 -5240 28452 -5234
rect 28848 -5240 28908 -5234
rect 29306 -5240 29366 -5234
rect 29770 -5240 29830 -5234
rect 30224 -5240 30284 -5234
rect 30682 -5240 30742 -5234
rect 27536 -5300 27932 -5240
rect 27992 -5300 28392 -5240
rect 28452 -5300 28848 -5240
rect 28908 -5300 29306 -5240
rect 29366 -5300 29770 -5240
rect 29830 -5300 30224 -5240
rect 30284 -5300 30682 -5240
rect 30910 -5288 30916 -5228
rect 30976 -5288 30982 -5228
rect 31142 -5240 31202 -5234
rect 31598 -5240 31658 -5234
rect 32058 -5240 32118 -5234
rect 32514 -5240 32574 -5234
rect 32970 -5240 33030 -5234
rect 33426 -5240 33486 -5234
rect 33884 -5240 33944 -5234
rect 34344 -5240 34404 -5234
rect 27476 -5306 27536 -5300
rect 27932 -5306 27992 -5300
rect 28392 -5306 28452 -5300
rect 28848 -5306 28908 -5300
rect 29306 -5306 29366 -5300
rect 29770 -5306 29830 -5300
rect 30224 -5306 30284 -5300
rect 30682 -5306 30742 -5300
rect 25234 -5664 25294 -5658
rect 11750 -5886 15976 -5826
rect 16180 -5724 25234 -5664
rect 11690 -5892 11750 -5886
rect 15124 -5928 15184 -5922
rect 16180 -5928 16240 -5724
rect 25234 -5730 25294 -5724
rect 26690 -5826 26750 -5820
rect 30916 -5826 30976 -5288
rect 31202 -5300 31598 -5240
rect 31658 -5300 32058 -5240
rect 32118 -5300 32514 -5240
rect 32574 -5300 32970 -5240
rect 33030 -5300 33426 -5240
rect 33486 -5300 33884 -5240
rect 33944 -5300 34344 -5240
rect 31142 -5306 31202 -5300
rect 31598 -5306 31658 -5300
rect 32058 -5306 32118 -5300
rect 32514 -5306 32574 -5300
rect 32970 -5306 33030 -5300
rect 33426 -5306 33486 -5300
rect 33884 -5306 33944 -5300
rect 34344 -5306 34404 -5300
rect 26750 -5886 30976 -5826
rect 26690 -5892 26750 -5886
rect 15184 -5988 16240 -5928
rect 15124 -5994 15184 -5988
rect 11908 -7564 11914 -7504
rect 11974 -7564 11980 -7504
rect 12370 -7564 12376 -7504
rect 12436 -7564 12442 -7504
rect 12824 -7560 12830 -7500
rect 12890 -7560 12896 -7500
rect 13286 -7560 13292 -7500
rect 13352 -7560 13358 -7500
rect 11914 -7958 11974 -7564
rect 12376 -7958 12436 -7564
rect 12830 -7958 12890 -7560
rect 13292 -7958 13352 -7560
rect 13740 -7566 13746 -7506
rect 13806 -7566 13812 -7506
rect 14190 -7560 14196 -7500
rect 14256 -7560 14262 -7500
rect 14656 -7560 14662 -7500
rect 14722 -7560 14728 -7500
rect 13746 -7958 13806 -7566
rect 14196 -7958 14256 -7560
rect 14662 -7958 14722 -7560
rect 15112 -7564 15118 -7504
rect 15178 -7564 15184 -7504
rect 16910 -7564 16916 -7504
rect 16976 -7564 16982 -7504
rect 17372 -7556 17378 -7496
rect 17438 -7556 17444 -7496
rect 15118 -7958 15178 -7564
rect 11912 -8018 15178 -7958
rect 11914 -8440 11974 -8018
rect 12376 -8434 12436 -8018
rect 12376 -8500 12436 -8494
rect 12830 -8440 12890 -8018
rect 13292 -8434 13352 -8018
rect 13292 -8500 13352 -8494
rect 13746 -8434 13806 -8018
rect 13746 -8500 13806 -8494
rect 14196 -8434 14256 -8018
rect 14196 -8500 14256 -8494
rect 14662 -8440 14722 -8018
rect 15118 -8434 15178 -8018
rect 15352 -7626 15412 -7620
rect 15352 -7964 15412 -7686
rect 16916 -7964 16976 -7564
rect 17378 -7964 17438 -7556
rect 17826 -7562 17832 -7502
rect 17892 -7562 17898 -7502
rect 18288 -7562 18294 -7502
rect 18354 -7562 18360 -7502
rect 18742 -7562 18748 -7502
rect 18808 -7562 18814 -7502
rect 19192 -7556 19198 -7496
rect 19258 -7556 19264 -7496
rect 17832 -7964 17892 -7562
rect 18294 -7964 18354 -7562
rect 18748 -7964 18808 -7562
rect 19198 -7964 19258 -7556
rect 19658 -7562 19664 -7502
rect 19724 -7562 19730 -7502
rect 20114 -7562 20120 -7502
rect 20180 -7562 20186 -7502
rect 19664 -7964 19724 -7562
rect 20120 -7964 20180 -7562
rect 26908 -7564 26914 -7504
rect 26974 -7564 26980 -7504
rect 27370 -7564 27376 -7504
rect 27436 -7564 27442 -7504
rect 27824 -7560 27830 -7500
rect 27890 -7560 27896 -7500
rect 28286 -7560 28292 -7500
rect 28352 -7560 28358 -7500
rect 20346 -7692 20352 -7632
rect 20412 -7692 20418 -7632
rect 15352 -8024 20180 -7964
rect 15352 -8306 15412 -8024
rect 15346 -8366 15352 -8306
rect 15412 -8366 15418 -8306
rect 15118 -8500 15178 -8494
rect 16916 -8434 16976 -8024
rect 16916 -8500 16976 -8494
rect 17378 -8436 17438 -8024
rect 11914 -8506 11974 -8500
rect 12830 -8506 12890 -8500
rect 14662 -8506 14722 -8500
rect 17378 -8502 17438 -8496
rect 17832 -8436 17892 -8024
rect 17832 -8502 17892 -8496
rect 18294 -8436 18354 -8024
rect 18294 -8502 18354 -8496
rect 18748 -8436 18808 -8024
rect 19198 -8430 19258 -8024
rect 19198 -8496 19258 -8490
rect 19664 -8434 19724 -8024
rect 18748 -8502 18808 -8496
rect 19664 -8500 19724 -8494
rect 20120 -8434 20180 -8024
rect 20352 -7968 20412 -7692
rect 25616 -7958 25676 -7949
rect 26914 -7958 26974 -7564
rect 27376 -7958 27436 -7564
rect 27830 -7958 27890 -7560
rect 28292 -7958 28352 -7560
rect 28740 -7566 28746 -7506
rect 28806 -7566 28812 -7506
rect 29190 -7560 29196 -7500
rect 29256 -7560 29262 -7500
rect 29656 -7560 29662 -7500
rect 29722 -7560 29728 -7500
rect 28746 -7958 28806 -7566
rect 29196 -7958 29256 -7560
rect 29662 -7958 29722 -7560
rect 30112 -7564 30118 -7504
rect 30178 -7564 30184 -7504
rect 31910 -7564 31916 -7504
rect 31976 -7564 31982 -7504
rect 32372 -7556 32378 -7496
rect 32438 -7556 32444 -7496
rect 30118 -7958 30178 -7564
rect 20352 -8028 21438 -7968
rect 25676 -8018 30178 -7958
rect 25616 -8027 25676 -8018
rect 20352 -8294 20412 -8028
rect 21338 -8157 21438 -8028
rect 21334 -8247 21343 -8157
rect 21433 -8247 21442 -8157
rect 21338 -8252 21438 -8247
rect 20352 -8360 20412 -8354
rect 20120 -8500 20180 -8494
rect 26914 -8440 26974 -8018
rect 27376 -8434 27436 -8018
rect 27376 -8500 27436 -8494
rect 27830 -8440 27890 -8018
rect 28292 -8434 28352 -8018
rect 28292 -8500 28352 -8494
rect 28746 -8434 28806 -8018
rect 28746 -8500 28806 -8494
rect 29196 -8434 29256 -8018
rect 29196 -8500 29256 -8494
rect 29662 -8440 29722 -8018
rect 30118 -8434 30178 -8018
rect 30352 -7626 30412 -7620
rect 30352 -7964 30412 -7686
rect 31916 -7964 31976 -7564
rect 32378 -7964 32438 -7556
rect 32826 -7562 32832 -7502
rect 32892 -7562 32898 -7502
rect 33288 -7562 33294 -7502
rect 33354 -7562 33360 -7502
rect 33742 -7562 33748 -7502
rect 33808 -7562 33814 -7502
rect 34192 -7556 34198 -7496
rect 34258 -7556 34264 -7496
rect 32832 -7964 32892 -7562
rect 33294 -7964 33354 -7562
rect 33748 -7964 33808 -7562
rect 34198 -7964 34258 -7556
rect 34658 -7562 34664 -7502
rect 34724 -7562 34730 -7502
rect 35114 -7562 35120 -7502
rect 35180 -7562 35186 -7502
rect 34664 -7964 34724 -7562
rect 35120 -7964 35180 -7562
rect 35346 -7692 35352 -7632
rect 35412 -7692 35418 -7632
rect 30352 -8024 35180 -7964
rect 30352 -8306 30412 -8024
rect 30346 -8366 30352 -8306
rect 30412 -8366 30418 -8306
rect 30118 -8500 30178 -8494
rect 31916 -8434 31976 -8024
rect 31916 -8500 31976 -8494
rect 32378 -8436 32438 -8024
rect 26914 -8506 26974 -8500
rect 27830 -8506 27890 -8500
rect 29662 -8506 29722 -8500
rect 32378 -8502 32438 -8496
rect 32832 -8436 32892 -8024
rect 32832 -8502 32892 -8496
rect 33294 -8436 33354 -8024
rect 33294 -8502 33354 -8496
rect 33748 -8436 33808 -8024
rect 34198 -8430 34258 -8024
rect 34198 -8496 34258 -8490
rect 34664 -8434 34724 -8024
rect 33748 -8502 33808 -8496
rect 34664 -8500 34724 -8494
rect 35120 -8434 35180 -8024
rect 35352 -7968 35412 -7692
rect 36338 -7968 36438 -778
rect 35352 -8028 36438 -7968
rect 35352 -8294 35412 -8028
rect 36338 -8157 36438 -8028
rect 36334 -8247 36343 -8157
rect 36433 -8247 36442 -8157
rect 36338 -8252 36438 -8247
rect 35352 -8360 35412 -8354
rect 35120 -8500 35180 -8494
rect 15116 -9650 15176 -9644
rect 25546 -9650 25606 -9644
rect 15176 -9710 25546 -9650
rect 25606 -9710 26914 -9650
rect 26974 -9710 26980 -9650
rect 15116 -9716 15176 -9710
rect 25546 -9716 25606 -9710
rect 11160 -9902 20930 -9874
rect 11160 -9988 11210 -9902
rect 11306 -9988 11790 -9902
rect 11886 -9988 12390 -9902
rect 12486 -9988 12990 -9902
rect 13086 -9988 13590 -9902
rect 13686 -9988 14190 -9902
rect 14286 -9988 14790 -9902
rect 14886 -9988 15390 -9902
rect 15486 -9988 15990 -9902
rect 16086 -9988 16590 -9902
rect 16686 -9988 17190 -9902
rect 17286 -9988 17790 -9902
rect 17886 -9988 18390 -9902
rect 18486 -9988 18990 -9902
rect 19086 -9988 19590 -9902
rect 19686 -9988 20190 -9902
rect 20286 -9988 20790 -9902
rect 20886 -9988 20930 -9902
rect 11160 -10018 20930 -9988
rect 26160 -9902 35930 -9874
rect 26160 -9988 26210 -9902
rect 26306 -9988 26790 -9902
rect 26886 -9988 27390 -9902
rect 27486 -9988 27990 -9902
rect 28086 -9988 28590 -9902
rect 28686 -9988 29190 -9902
rect 29286 -9988 29790 -9902
rect 29886 -9988 30390 -9902
rect 30486 -9988 30990 -9902
rect 31086 -9988 31590 -9902
rect 31686 -9988 32190 -9902
rect 32286 -9988 32790 -9902
rect 32886 -9988 33390 -9902
rect 33486 -9988 33990 -9902
rect 34086 -9988 34590 -9902
rect 34686 -9988 35190 -9902
rect 35286 -9988 35790 -9902
rect 35886 -9988 35930 -9902
rect 26160 -10018 35930 -9988
rect 10924 -10166 11524 -10156
rect 10924 -10476 11524 -10466
rect 20556 -10166 21156 -10156
rect 20556 -10476 21156 -10466
rect 25924 -10166 26524 -10156
rect 25924 -10476 26524 -10466
rect 35556 -10166 36156 -10156
rect 35556 -10476 36156 -10466
rect 14878 -11138 15478 -11128
rect 14878 -11448 15478 -11438
rect 24510 -11138 25110 -11128
rect 24510 -11448 25110 -11438
rect 29878 -11138 30478 -11128
rect 29878 -11448 30478 -11438
rect 39510 -11138 40110 -11128
rect 39510 -11448 40110 -11438
rect 15104 -11616 24874 -11586
rect 15104 -11702 15148 -11616
rect 15244 -11702 15748 -11616
rect 15844 -11702 16348 -11616
rect 16444 -11702 16948 -11616
rect 17044 -11702 17548 -11616
rect 17644 -11702 18148 -11616
rect 18244 -11702 18748 -11616
rect 18844 -11702 19348 -11616
rect 19444 -11702 19948 -11616
rect 20044 -11702 20548 -11616
rect 20644 -11702 21148 -11616
rect 21244 -11702 21748 -11616
rect 21844 -11702 22348 -11616
rect 22444 -11702 22948 -11616
rect 23044 -11702 23548 -11616
rect 23644 -11702 24148 -11616
rect 24244 -11702 24728 -11616
rect 24824 -11702 24874 -11616
rect 15104 -11730 24874 -11702
rect 30104 -11616 39874 -11586
rect 30104 -11702 30148 -11616
rect 30244 -11702 30748 -11616
rect 30844 -11702 31348 -11616
rect 31444 -11702 31948 -11616
rect 32044 -11702 32548 -11616
rect 32644 -11702 33148 -11616
rect 33244 -11702 33748 -11616
rect 33844 -11702 34348 -11616
rect 34444 -11702 34948 -11616
rect 35044 -11702 35548 -11616
rect 35644 -11702 36148 -11616
rect 36244 -11702 36748 -11616
rect 36844 -11702 37348 -11616
rect 37444 -11702 37948 -11616
rect 38044 -11702 38548 -11616
rect 38644 -11702 39148 -11616
rect 39244 -11702 39728 -11616
rect 39824 -11702 39874 -11616
rect 30104 -11730 39874 -11702
rect 24062 -11894 24122 -11888
rect 24122 -11954 25546 -11894
rect 25606 -11954 35856 -11894
rect 35916 -11954 35922 -11894
rect 24062 -11960 24122 -11954
rect 15854 -13110 15914 -13104
rect 15622 -13250 15682 -13244
rect 10630 -13357 10690 -13352
rect 14596 -13357 14696 -13352
rect 10600 -13447 10609 -13357
rect 10699 -13447 10708 -13357
rect 14592 -13447 14601 -13357
rect 14691 -13447 14700 -13357
rect 10630 -25958 10690 -13447
rect 14596 -13576 14696 -13447
rect 15622 -13576 15682 -13310
rect 14596 -13636 15682 -13576
rect 15622 -13912 15682 -13636
rect 15854 -13580 15914 -13170
rect 16310 -13110 16370 -13104
rect 17226 -13108 17286 -13102
rect 16310 -13580 16370 -13170
rect 16776 -13114 16836 -13108
rect 16776 -13580 16836 -13174
rect 17226 -13580 17286 -13168
rect 17680 -13108 17740 -13102
rect 17680 -13580 17740 -13168
rect 18142 -13108 18202 -13102
rect 18142 -13580 18202 -13168
rect 18596 -13108 18656 -13102
rect 21312 -13104 21372 -13098
rect 23144 -13104 23204 -13098
rect 24060 -13104 24120 -13098
rect 18596 -13580 18656 -13168
rect 19058 -13110 19118 -13104
rect 19058 -13580 19118 -13170
rect 20856 -13110 20916 -13104
rect 20616 -13298 20622 -13238
rect 20682 -13298 20688 -13238
rect 20622 -13580 20682 -13298
rect 15854 -13640 20682 -13580
rect 15616 -13972 15622 -13912
rect 15682 -13972 15688 -13912
rect 15854 -14042 15914 -13640
rect 16310 -14042 16370 -13640
rect 15848 -14102 15854 -14042
rect 15914 -14102 15920 -14042
rect 16304 -14102 16310 -14042
rect 16370 -14102 16376 -14042
rect 16776 -14048 16836 -13640
rect 17226 -14042 17286 -13640
rect 17680 -14042 17740 -13640
rect 18142 -14042 18202 -13640
rect 16770 -14108 16776 -14048
rect 16836 -14108 16842 -14048
rect 17220 -14102 17226 -14042
rect 17286 -14102 17292 -14042
rect 17674 -14102 17680 -14042
rect 17740 -14102 17746 -14042
rect 18136 -14102 18142 -14042
rect 18202 -14102 18208 -14042
rect 18596 -14048 18656 -13640
rect 19058 -14040 19118 -13640
rect 20622 -13918 20682 -13640
rect 20622 -13984 20682 -13978
rect 20856 -13586 20916 -13170
rect 21312 -13586 21372 -13164
rect 21778 -13110 21838 -13104
rect 21778 -13586 21838 -13170
rect 22228 -13110 22288 -13104
rect 22228 -13586 22288 -13170
rect 22682 -13110 22742 -13104
rect 22682 -13586 22742 -13170
rect 23144 -13586 23204 -13164
rect 23598 -13110 23658 -13104
rect 23598 -13586 23658 -13170
rect 24060 -13586 24120 -13164
rect 30854 -13110 30914 -13104
rect 30622 -13250 30682 -13244
rect 29596 -13357 29696 -13352
rect 29592 -13447 29601 -13357
rect 29691 -13447 29700 -13357
rect 29596 -13576 29696 -13447
rect 30622 -13576 30682 -13310
rect 25300 -13586 25360 -13577
rect 20856 -13646 25300 -13586
rect 29596 -13636 30682 -13576
rect 20856 -14040 20916 -13646
rect 18590 -14108 18596 -14048
rect 18656 -14108 18662 -14048
rect 19052 -14100 19058 -14040
rect 19118 -14100 19124 -14040
rect 20850 -14100 20856 -14040
rect 20916 -14100 20922 -14040
rect 21312 -14044 21372 -13646
rect 21778 -14044 21838 -13646
rect 22228 -14038 22288 -13646
rect 21306 -14104 21312 -14044
rect 21372 -14104 21378 -14044
rect 21772 -14104 21778 -14044
rect 21838 -14104 21844 -14044
rect 22222 -14098 22228 -14038
rect 22288 -14098 22294 -14038
rect 22682 -14044 22742 -13646
rect 23144 -14044 23204 -13646
rect 23598 -14040 23658 -13646
rect 24060 -14040 24120 -13646
rect 25300 -13655 25360 -13646
rect 30622 -13912 30682 -13636
rect 30854 -13580 30914 -13170
rect 31310 -13110 31370 -13104
rect 32226 -13108 32286 -13102
rect 31310 -13580 31370 -13170
rect 31776 -13114 31836 -13108
rect 31776 -13580 31836 -13174
rect 32226 -13580 32286 -13168
rect 32680 -13108 32740 -13102
rect 32680 -13580 32740 -13168
rect 33142 -13108 33202 -13102
rect 33142 -13580 33202 -13168
rect 33596 -13108 33656 -13102
rect 36312 -13104 36372 -13098
rect 38144 -13104 38204 -13098
rect 39060 -13104 39120 -13098
rect 33596 -13580 33656 -13168
rect 34058 -13110 34118 -13104
rect 34058 -13580 34118 -13170
rect 35856 -13110 35916 -13104
rect 35616 -13298 35622 -13238
rect 35682 -13298 35688 -13238
rect 35622 -13580 35682 -13298
rect 30854 -13640 35682 -13580
rect 30616 -13972 30622 -13912
rect 30682 -13972 30688 -13912
rect 22676 -14104 22682 -14044
rect 22742 -14104 22748 -14044
rect 23138 -14104 23144 -14044
rect 23204 -14104 23210 -14044
rect 23592 -14100 23598 -14040
rect 23658 -14100 23664 -14040
rect 24054 -14100 24060 -14040
rect 24120 -14100 24126 -14040
rect 30854 -14042 30914 -13640
rect 31310 -14042 31370 -13640
rect 30848 -14102 30854 -14042
rect 30914 -14102 30920 -14042
rect 31304 -14102 31310 -14042
rect 31370 -14102 31376 -14042
rect 31776 -14048 31836 -13640
rect 32226 -14042 32286 -13640
rect 32680 -14042 32740 -13640
rect 33142 -14042 33202 -13640
rect 31770 -14108 31776 -14048
rect 31836 -14108 31842 -14048
rect 32220 -14102 32226 -14042
rect 32286 -14102 32292 -14042
rect 32674 -14102 32680 -14042
rect 32740 -14102 32746 -14042
rect 33136 -14102 33142 -14042
rect 33202 -14102 33208 -14042
rect 33596 -14048 33656 -13640
rect 34058 -14040 34118 -13640
rect 35622 -13918 35682 -13640
rect 35622 -13984 35682 -13978
rect 35856 -13586 35916 -13170
rect 36312 -13586 36372 -13164
rect 36778 -13110 36838 -13104
rect 36778 -13586 36838 -13170
rect 37228 -13110 37288 -13104
rect 37228 -13586 37288 -13170
rect 37682 -13110 37742 -13104
rect 37682 -13586 37742 -13170
rect 38144 -13586 38204 -13164
rect 38598 -13110 38658 -13104
rect 38598 -13586 38658 -13170
rect 39060 -13586 39120 -13164
rect 35856 -13646 40380 -13586
rect 35856 -14040 35916 -13646
rect 33590 -14108 33596 -14048
rect 33656 -14108 33662 -14048
rect 34052 -14100 34058 -14040
rect 34118 -14100 34124 -14040
rect 35850 -14100 35856 -14040
rect 35916 -14100 35922 -14040
rect 36312 -14044 36372 -13646
rect 36778 -14044 36838 -13646
rect 37228 -14038 37288 -13646
rect 36306 -14104 36312 -14044
rect 36372 -14104 36378 -14044
rect 36772 -14104 36778 -14044
rect 36838 -14104 36844 -14044
rect 37222 -14098 37228 -14038
rect 37288 -14098 37294 -14038
rect 37682 -14044 37742 -13646
rect 38144 -14044 38204 -13646
rect 38598 -14040 38658 -13646
rect 39060 -14040 39120 -13646
rect 37676 -14104 37682 -14044
rect 37742 -14104 37748 -14044
rect 38138 -14104 38144 -14044
rect 38204 -14104 38210 -14044
rect 38592 -14100 38598 -14040
rect 38658 -14100 38664 -14040
rect 39054 -14100 39060 -14040
rect 39120 -14100 39126 -14040
rect 24284 -15718 24344 -15712
rect 39284 -15718 39344 -15712
rect 20058 -15778 24284 -15718
rect 16630 -16304 16690 -16298
rect 17090 -16304 17150 -16298
rect 17548 -16304 17608 -16298
rect 18004 -16304 18064 -16298
rect 18460 -16304 18520 -16298
rect 18916 -16304 18976 -16298
rect 19376 -16304 19436 -16298
rect 19832 -16304 19892 -16298
rect 16690 -16364 17090 -16304
rect 17150 -16364 17548 -16304
rect 17608 -16364 18004 -16304
rect 18064 -16364 18460 -16304
rect 18520 -16364 18916 -16304
rect 18976 -16364 19376 -16304
rect 19436 -16364 19832 -16304
rect 20058 -16316 20118 -15778
rect 24284 -15784 24344 -15778
rect 35058 -15778 39284 -15718
rect 20292 -16304 20352 -16298
rect 20750 -16304 20810 -16298
rect 21204 -16304 21264 -16298
rect 21668 -16304 21728 -16298
rect 22126 -16304 22186 -16298
rect 22582 -16304 22642 -16298
rect 23042 -16304 23102 -16298
rect 23498 -16304 23558 -16298
rect 31630 -16304 31690 -16298
rect 32090 -16304 32150 -16298
rect 32548 -16304 32608 -16298
rect 33004 -16304 33064 -16298
rect 33460 -16304 33520 -16298
rect 33916 -16304 33976 -16298
rect 34376 -16304 34436 -16298
rect 34832 -16304 34892 -16298
rect 16630 -16370 16690 -16364
rect 17090 -16370 17150 -16364
rect 17548 -16370 17608 -16364
rect 18004 -16370 18064 -16364
rect 18460 -16370 18520 -16364
rect 18916 -16370 18976 -16364
rect 19376 -16370 19436 -16364
rect 19832 -16370 19892 -16364
rect 20052 -16376 20058 -16316
rect 20118 -16376 20124 -16316
rect 20352 -16364 20750 -16304
rect 20810 -16364 21204 -16304
rect 21264 -16364 21668 -16304
rect 21728 -16364 22126 -16304
rect 22186 -16364 22582 -16304
rect 22642 -16364 23042 -16304
rect 23102 -16364 23498 -16304
rect 23558 -16364 25406 -16304
rect 25466 -16364 31630 -16304
rect 31690 -16364 32090 -16304
rect 32150 -16364 32548 -16304
rect 32608 -16364 33004 -16304
rect 33064 -16364 33460 -16304
rect 33520 -16364 33916 -16304
rect 33976 -16364 34376 -16304
rect 34436 -16364 34832 -16304
rect 35058 -16316 35118 -15778
rect 39284 -15784 39344 -15778
rect 35292 -16304 35352 -16298
rect 35750 -16304 35810 -16298
rect 36204 -16304 36264 -16298
rect 36668 -16304 36728 -16298
rect 37126 -16304 37186 -16298
rect 37582 -16304 37642 -16298
rect 38042 -16304 38102 -16298
rect 38498 -16304 38558 -16298
rect 20292 -16370 20352 -16364
rect 20750 -16370 20810 -16364
rect 21204 -16370 21264 -16364
rect 21668 -16370 21728 -16364
rect 22126 -16370 22186 -16364
rect 22582 -16370 22642 -16364
rect 23042 -16370 23102 -16364
rect 23498 -16370 23558 -16364
rect 31630 -16370 31690 -16364
rect 32090 -16370 32150 -16364
rect 32548 -16370 32608 -16364
rect 33004 -16370 33064 -16364
rect 33460 -16370 33520 -16364
rect 33916 -16370 33976 -16364
rect 34376 -16370 34436 -16364
rect 34832 -16370 34892 -16364
rect 35052 -16376 35058 -16316
rect 35118 -16376 35124 -16316
rect 35352 -16364 35750 -16304
rect 35810 -16364 36204 -16304
rect 36264 -16364 36668 -16304
rect 36728 -16364 37126 -16304
rect 37186 -16364 37582 -16304
rect 37642 -16364 38042 -16304
rect 38102 -16364 38498 -16304
rect 35292 -16370 35352 -16364
rect 35750 -16370 35810 -16364
rect 36204 -16370 36264 -16364
rect 36668 -16370 36728 -16364
rect 37126 -16370 37186 -16364
rect 37582 -16370 37642 -16364
rect 38042 -16370 38102 -16364
rect 38498 -16370 38558 -16364
rect 16626 -18278 16686 -18272
rect 17086 -18278 17146 -18272
rect 17544 -18278 17604 -18272
rect 18000 -18278 18060 -18272
rect 18456 -18278 18516 -18272
rect 18912 -18278 18972 -18272
rect 19368 -18278 19428 -18272
rect 19826 -18278 19886 -18272
rect 20294 -18278 20354 -18272
rect 20750 -18278 20810 -18272
rect 21200 -18278 21260 -18272
rect 21664 -18278 21724 -18272
rect 22122 -18278 22182 -18272
rect 22578 -18278 22638 -18272
rect 23038 -18278 23098 -18272
rect 23494 -18278 23554 -18272
rect 16686 -18338 17086 -18278
rect 17146 -18338 17544 -18278
rect 17604 -18338 18000 -18278
rect 18060 -18338 18456 -18278
rect 18516 -18338 18912 -18278
rect 18972 -18338 19368 -18278
rect 19428 -18338 19826 -18278
rect 19886 -18338 20294 -18278
rect 20354 -18338 20750 -18278
rect 20810 -18338 21200 -18278
rect 21260 -18338 21664 -18278
rect 21724 -18338 22122 -18278
rect 22182 -18338 22578 -18278
rect 22638 -18338 23038 -18278
rect 23098 -18338 23494 -18278
rect 16626 -18344 16686 -18338
rect 17086 -18344 17146 -18338
rect 17544 -18344 17604 -18338
rect 18000 -18344 18060 -18338
rect 18456 -18344 18516 -18338
rect 18912 -18344 18972 -18338
rect 19368 -18344 19428 -18338
rect 19826 -18344 19886 -18338
rect 20294 -18344 20354 -18338
rect 20750 -18344 20810 -18338
rect 21200 -18344 21260 -18338
rect 21664 -18344 21724 -18338
rect 22122 -18344 22182 -18338
rect 22578 -18344 22638 -18338
rect 23038 -18344 23098 -18338
rect 23494 -18344 23554 -18338
rect 31626 -18278 31686 -18272
rect 32086 -18278 32146 -18272
rect 32544 -18278 32604 -18272
rect 33000 -18278 33060 -18272
rect 33456 -18278 33516 -18272
rect 33912 -18278 33972 -18272
rect 34368 -18278 34428 -18272
rect 34826 -18278 34886 -18272
rect 35294 -18278 35354 -18272
rect 35750 -18278 35810 -18272
rect 36200 -18278 36260 -18272
rect 36664 -18278 36724 -18272
rect 37122 -18278 37182 -18272
rect 37578 -18278 37638 -18272
rect 38038 -18278 38098 -18272
rect 38494 -18278 38554 -18272
rect 31686 -18338 32086 -18278
rect 32146 -18338 32544 -18278
rect 32604 -18338 33000 -18278
rect 33060 -18338 33456 -18278
rect 33516 -18338 33912 -18278
rect 33972 -18338 34368 -18278
rect 34428 -18338 34826 -18278
rect 34886 -18338 35294 -18278
rect 35354 -18338 35750 -18278
rect 35810 -18338 36200 -18278
rect 36260 -18338 36664 -18278
rect 36724 -18338 37122 -18278
rect 37182 -18338 37578 -18278
rect 37638 -18338 38038 -18278
rect 38098 -18338 38494 -18278
rect 31626 -18344 31686 -18338
rect 32086 -18344 32146 -18338
rect 32544 -18344 32604 -18338
rect 33000 -18344 33060 -18338
rect 33456 -18344 33516 -18338
rect 33912 -18344 33972 -18338
rect 34368 -18344 34428 -18338
rect 34826 -18344 34886 -18338
rect 35294 -18344 35354 -18338
rect 35750 -18344 35810 -18338
rect 36200 -18344 36260 -18338
rect 36664 -18344 36724 -18338
rect 37122 -18344 37182 -18338
rect 37578 -18344 37638 -18338
rect 38038 -18344 38098 -18338
rect 38494 -18344 38554 -18338
rect 15916 -18910 24272 -18900
rect 15916 -18996 15942 -18910
rect 16038 -18996 16362 -18910
rect 16458 -18996 16962 -18910
rect 17058 -18996 17562 -18910
rect 17658 -18996 18162 -18910
rect 18258 -18996 18762 -18910
rect 18858 -18996 19362 -18910
rect 19458 -18996 19962 -18910
rect 20058 -18996 20562 -18910
rect 20658 -18996 21162 -18910
rect 21258 -18996 21762 -18910
rect 21858 -18996 22362 -18910
rect 22458 -18996 22962 -18910
rect 23058 -18996 23562 -18910
rect 23658 -18996 24162 -18910
rect 24258 -18996 24272 -18910
rect 15916 -19010 24272 -18996
rect 30916 -18910 39272 -18900
rect 30916 -18996 30942 -18910
rect 31038 -18996 31362 -18910
rect 31458 -18996 31962 -18910
rect 32058 -18996 32562 -18910
rect 32658 -18996 33162 -18910
rect 33258 -18996 33762 -18910
rect 33858 -18996 34362 -18910
rect 34458 -18996 34962 -18910
rect 35058 -18996 35562 -18910
rect 35658 -18996 36162 -18910
rect 36258 -18996 36762 -18910
rect 36858 -18996 37362 -18910
rect 37458 -18996 37962 -18910
rect 38058 -18996 38562 -18910
rect 38658 -18996 39162 -18910
rect 39258 -18996 39272 -18910
rect 30916 -19010 39272 -18996
rect 14878 -19170 15478 -19160
rect 14878 -19480 15478 -19470
rect 24510 -19170 25110 -19160
rect 24510 -19480 25110 -19470
rect 29878 -19170 30478 -19160
rect 29878 -19480 30478 -19470
rect 39510 -19170 40110 -19160
rect 39510 -19480 40110 -19470
rect 10924 -20134 11524 -20124
rect 10924 -20444 11524 -20434
rect 20556 -20134 21156 -20124
rect 20556 -20444 21156 -20434
rect 25924 -20134 26524 -20124
rect 25924 -20444 26524 -20434
rect 35556 -20134 36156 -20124
rect 35556 -20444 36156 -20434
rect 11762 -20608 20118 -20594
rect 11762 -20694 11776 -20608
rect 11872 -20694 12376 -20608
rect 12472 -20694 12976 -20608
rect 13072 -20694 13576 -20608
rect 13672 -20694 14176 -20608
rect 14272 -20694 14776 -20608
rect 14872 -20694 15376 -20608
rect 15472 -20694 15976 -20608
rect 16072 -20694 16576 -20608
rect 16672 -20694 17176 -20608
rect 17272 -20694 17776 -20608
rect 17872 -20694 18376 -20608
rect 18472 -20694 18976 -20608
rect 19072 -20694 19576 -20608
rect 19672 -20694 19996 -20608
rect 20092 -20694 20118 -20608
rect 11762 -20704 20118 -20694
rect 26762 -20608 35118 -20594
rect 26762 -20694 26776 -20608
rect 26872 -20694 27376 -20608
rect 27472 -20694 27976 -20608
rect 28072 -20694 28576 -20608
rect 28672 -20694 29176 -20608
rect 29272 -20694 29776 -20608
rect 29872 -20694 30376 -20608
rect 30472 -20694 30976 -20608
rect 31072 -20694 31576 -20608
rect 31672 -20694 32176 -20608
rect 32272 -20694 32776 -20608
rect 32872 -20694 33376 -20608
rect 33472 -20694 33976 -20608
rect 34072 -20694 34576 -20608
rect 34672 -20694 34996 -20608
rect 35092 -20694 35118 -20608
rect 26762 -20704 35118 -20694
rect 12480 -21266 12540 -21260
rect 12936 -21266 12996 -21260
rect 13396 -21266 13456 -21260
rect 13852 -21266 13912 -21260
rect 14310 -21266 14370 -21260
rect 14774 -21266 14834 -21260
rect 15224 -21266 15284 -21260
rect 15680 -21266 15740 -21260
rect 16148 -21266 16208 -21260
rect 16606 -21266 16666 -21260
rect 17062 -21266 17122 -21260
rect 17518 -21266 17578 -21260
rect 17974 -21266 18034 -21260
rect 18430 -21266 18490 -21260
rect 18888 -21266 18948 -21260
rect 19348 -21266 19408 -21260
rect 12540 -21326 12936 -21266
rect 12996 -21326 13396 -21266
rect 13456 -21326 13852 -21266
rect 13912 -21326 14310 -21266
rect 14370 -21326 14774 -21266
rect 14834 -21326 15224 -21266
rect 15284 -21326 15680 -21266
rect 15740 -21326 16148 -21266
rect 16208 -21326 16606 -21266
rect 16666 -21326 17062 -21266
rect 17122 -21326 17518 -21266
rect 17578 -21326 17974 -21266
rect 18034 -21326 18430 -21266
rect 18490 -21326 18888 -21266
rect 18948 -21326 19348 -21266
rect 12480 -21332 12540 -21326
rect 12936 -21332 12996 -21326
rect 13396 -21332 13456 -21326
rect 13852 -21332 13912 -21326
rect 14310 -21332 14370 -21326
rect 14774 -21332 14834 -21326
rect 15224 -21332 15284 -21326
rect 15680 -21332 15740 -21326
rect 16148 -21332 16208 -21326
rect 16606 -21332 16666 -21326
rect 17062 -21332 17122 -21326
rect 17518 -21332 17578 -21326
rect 17974 -21332 18034 -21326
rect 18430 -21332 18490 -21326
rect 18888 -21332 18948 -21326
rect 19348 -21332 19408 -21326
rect 27480 -21266 27540 -21260
rect 27936 -21266 27996 -21260
rect 28396 -21266 28456 -21260
rect 28852 -21266 28912 -21260
rect 29310 -21266 29370 -21260
rect 29774 -21266 29834 -21260
rect 30224 -21266 30284 -21260
rect 30680 -21266 30740 -21260
rect 31148 -21266 31208 -21260
rect 31606 -21266 31666 -21260
rect 32062 -21266 32122 -21260
rect 32518 -21266 32578 -21260
rect 32974 -21266 33034 -21260
rect 33430 -21266 33490 -21260
rect 33888 -21266 33948 -21260
rect 34348 -21266 34408 -21260
rect 27540 -21326 27936 -21266
rect 27996 -21326 28396 -21266
rect 28456 -21326 28852 -21266
rect 28912 -21326 29310 -21266
rect 29370 -21326 29774 -21266
rect 29834 -21326 30224 -21266
rect 30284 -21326 30680 -21266
rect 30740 -21326 31148 -21266
rect 31208 -21326 31606 -21266
rect 31666 -21326 32062 -21266
rect 32122 -21326 32518 -21266
rect 32578 -21326 32974 -21266
rect 33034 -21326 33430 -21266
rect 33490 -21326 33888 -21266
rect 33948 -21326 34348 -21266
rect 27480 -21332 27540 -21326
rect 27936 -21332 27996 -21326
rect 28396 -21332 28456 -21326
rect 28852 -21332 28912 -21326
rect 29310 -21332 29370 -21326
rect 29774 -21332 29834 -21326
rect 30224 -21332 30284 -21326
rect 30680 -21332 30740 -21326
rect 31148 -21332 31208 -21326
rect 31606 -21332 31666 -21326
rect 32062 -21332 32122 -21326
rect 32518 -21332 32578 -21326
rect 32974 -21332 33034 -21326
rect 33430 -21332 33490 -21326
rect 33888 -21332 33948 -21326
rect 34348 -21332 34408 -21326
rect 12476 -23240 12536 -23234
rect 12932 -23240 12992 -23234
rect 13392 -23240 13452 -23234
rect 13848 -23240 13908 -23234
rect 14306 -23240 14366 -23234
rect 14770 -23240 14830 -23234
rect 15224 -23240 15284 -23234
rect 15682 -23240 15742 -23234
rect 12536 -23300 12932 -23240
rect 12992 -23300 13392 -23240
rect 13452 -23300 13848 -23240
rect 13908 -23300 14306 -23240
rect 14366 -23300 14770 -23240
rect 14830 -23300 15224 -23240
rect 15284 -23300 15682 -23240
rect 15910 -23288 15916 -23228
rect 15976 -23288 15982 -23228
rect 16142 -23240 16202 -23234
rect 16598 -23240 16658 -23234
rect 17058 -23240 17118 -23234
rect 17514 -23240 17574 -23234
rect 17970 -23240 18030 -23234
rect 18426 -23240 18486 -23234
rect 18884 -23240 18944 -23234
rect 19344 -23240 19404 -23234
rect 25406 -23240 25466 -23234
rect 27476 -23240 27536 -23234
rect 27932 -23240 27992 -23234
rect 28392 -23240 28452 -23234
rect 28848 -23240 28908 -23234
rect 29306 -23240 29366 -23234
rect 29770 -23240 29830 -23234
rect 30224 -23240 30284 -23234
rect 30682 -23240 30742 -23234
rect 12476 -23306 12536 -23300
rect 12932 -23306 12992 -23300
rect 13392 -23306 13452 -23300
rect 13848 -23306 13908 -23300
rect 14306 -23306 14366 -23300
rect 14770 -23306 14830 -23300
rect 15224 -23306 15284 -23300
rect 15682 -23306 15742 -23300
rect 11690 -23826 11750 -23820
rect 15916 -23826 15976 -23288
rect 16202 -23300 16598 -23240
rect 16658 -23300 17058 -23240
rect 17118 -23300 17514 -23240
rect 17574 -23300 17970 -23240
rect 18030 -23300 18426 -23240
rect 18486 -23300 18884 -23240
rect 18944 -23300 19344 -23240
rect 19404 -23300 25406 -23240
rect 25466 -23300 27476 -23240
rect 27536 -23300 27932 -23240
rect 27992 -23300 28392 -23240
rect 28452 -23300 28848 -23240
rect 28908 -23300 29306 -23240
rect 29366 -23300 29770 -23240
rect 29830 -23300 30224 -23240
rect 30284 -23300 30682 -23240
rect 30910 -23288 30916 -23228
rect 30976 -23288 30982 -23228
rect 31142 -23240 31202 -23234
rect 31598 -23240 31658 -23234
rect 32058 -23240 32118 -23234
rect 32514 -23240 32574 -23234
rect 32970 -23240 33030 -23234
rect 33426 -23240 33486 -23234
rect 33884 -23240 33944 -23234
rect 34344 -23240 34404 -23234
rect 16142 -23306 16202 -23300
rect 16598 -23306 16658 -23300
rect 17058 -23306 17118 -23300
rect 17514 -23306 17574 -23300
rect 17970 -23306 18030 -23300
rect 18426 -23306 18486 -23300
rect 18884 -23306 18944 -23300
rect 19344 -23306 19404 -23300
rect 25406 -23306 25466 -23300
rect 27476 -23306 27536 -23300
rect 27932 -23306 27992 -23300
rect 28392 -23306 28452 -23300
rect 28848 -23306 28908 -23300
rect 29306 -23306 29366 -23300
rect 29770 -23306 29830 -23300
rect 30224 -23306 30284 -23300
rect 30682 -23306 30742 -23300
rect 11750 -23886 15976 -23826
rect 26690 -23826 26750 -23820
rect 30916 -23826 30976 -23288
rect 31202 -23300 31598 -23240
rect 31658 -23300 32058 -23240
rect 32118 -23300 32514 -23240
rect 32574 -23300 32970 -23240
rect 33030 -23300 33426 -23240
rect 33486 -23300 33884 -23240
rect 33944 -23300 34344 -23240
rect 31142 -23306 31202 -23300
rect 31598 -23306 31658 -23300
rect 32058 -23306 32118 -23300
rect 32514 -23306 32574 -23300
rect 32970 -23306 33030 -23300
rect 33426 -23306 33486 -23300
rect 33884 -23306 33944 -23300
rect 34344 -23306 34404 -23300
rect 26750 -23886 30976 -23826
rect 11690 -23892 11750 -23886
rect 26690 -23892 26750 -23886
rect 11908 -25564 11914 -25504
rect 11974 -25564 11980 -25504
rect 12370 -25564 12376 -25504
rect 12436 -25564 12442 -25504
rect 12824 -25560 12830 -25500
rect 12890 -25560 12896 -25500
rect 13286 -25560 13292 -25500
rect 13352 -25560 13358 -25500
rect 11914 -25958 11974 -25564
rect 12376 -25958 12436 -25564
rect 12830 -25958 12890 -25560
rect 13292 -25958 13352 -25560
rect 13740 -25566 13746 -25506
rect 13806 -25566 13812 -25506
rect 14190 -25560 14196 -25500
rect 14256 -25560 14262 -25500
rect 14656 -25560 14662 -25500
rect 14722 -25560 14728 -25500
rect 13746 -25958 13806 -25566
rect 14196 -25958 14256 -25560
rect 14662 -25958 14722 -25560
rect 15112 -25564 15118 -25504
rect 15178 -25564 15184 -25504
rect 16910 -25564 16916 -25504
rect 16976 -25564 16982 -25504
rect 17372 -25556 17378 -25496
rect 17438 -25556 17444 -25496
rect 15118 -25958 15178 -25564
rect 10630 -26018 15178 -25958
rect 11914 -26440 11974 -26018
rect 12376 -26434 12436 -26018
rect 12376 -26500 12436 -26494
rect 12830 -26440 12890 -26018
rect 13292 -26434 13352 -26018
rect 13292 -26500 13352 -26494
rect 13746 -26434 13806 -26018
rect 13746 -26500 13806 -26494
rect 14196 -26434 14256 -26018
rect 14196 -26500 14256 -26494
rect 14662 -26440 14722 -26018
rect 15118 -26434 15178 -26018
rect 15352 -25626 15412 -25620
rect 15352 -25964 15412 -25686
rect 16916 -25964 16976 -25564
rect 17378 -25964 17438 -25556
rect 17826 -25562 17832 -25502
rect 17892 -25562 17898 -25502
rect 18288 -25562 18294 -25502
rect 18354 -25562 18360 -25502
rect 18742 -25562 18748 -25502
rect 18808 -25562 18814 -25502
rect 19192 -25556 19198 -25496
rect 19258 -25556 19264 -25496
rect 17832 -25964 17892 -25562
rect 18294 -25964 18354 -25562
rect 18748 -25964 18808 -25562
rect 19198 -25964 19258 -25556
rect 19658 -25562 19664 -25502
rect 19724 -25562 19730 -25502
rect 20114 -25562 20120 -25502
rect 20180 -25562 20186 -25502
rect 19664 -25964 19724 -25562
rect 20120 -25964 20180 -25562
rect 26908 -25564 26914 -25504
rect 26974 -25564 26980 -25504
rect 27370 -25564 27376 -25504
rect 27436 -25564 27442 -25504
rect 27824 -25560 27830 -25500
rect 27890 -25560 27896 -25500
rect 28286 -25560 28292 -25500
rect 28352 -25560 28358 -25500
rect 20346 -25692 20352 -25632
rect 20412 -25692 20418 -25632
rect 15352 -26024 20180 -25964
rect 15352 -26306 15412 -26024
rect 15346 -26366 15352 -26306
rect 15412 -26366 15418 -26306
rect 15118 -26500 15178 -26494
rect 16916 -26434 16976 -26024
rect 16916 -26500 16976 -26494
rect 17378 -26436 17438 -26024
rect 11914 -26506 11974 -26500
rect 12830 -26506 12890 -26500
rect 14662 -26506 14722 -26500
rect 17378 -26502 17438 -26496
rect 17832 -26436 17892 -26024
rect 17832 -26502 17892 -26496
rect 18294 -26436 18354 -26024
rect 18294 -26502 18354 -26496
rect 18748 -26436 18808 -26024
rect 19198 -26430 19258 -26024
rect 19198 -26496 19258 -26490
rect 19664 -26434 19724 -26024
rect 18748 -26502 18808 -26496
rect 19664 -26500 19724 -26494
rect 20120 -26434 20180 -26024
rect 20352 -25968 20412 -25692
rect 26914 -25958 26974 -25564
rect 27376 -25958 27436 -25564
rect 27830 -25958 27890 -25560
rect 28292 -25958 28352 -25560
rect 28740 -25566 28746 -25506
rect 28806 -25566 28812 -25506
rect 29190 -25560 29196 -25500
rect 29256 -25560 29262 -25500
rect 29656 -25560 29662 -25500
rect 29722 -25560 29728 -25500
rect 28746 -25958 28806 -25566
rect 29196 -25958 29256 -25560
rect 29662 -25958 29722 -25560
rect 30112 -25564 30118 -25504
rect 30178 -25564 30184 -25504
rect 31910 -25564 31916 -25504
rect 31976 -25564 31982 -25504
rect 32372 -25556 32378 -25496
rect 32438 -25556 32444 -25496
rect 30118 -25958 30178 -25564
rect 20352 -26028 21438 -25968
rect 20352 -26294 20412 -26028
rect 21338 -26157 21438 -26028
rect 25420 -26018 30178 -25958
rect 25420 -26157 25480 -26018
rect 21334 -26247 21343 -26157
rect 21433 -26247 21442 -26157
rect 25398 -26247 25407 -26157
rect 25497 -26247 25506 -26157
rect 21338 -26252 21438 -26247
rect 25420 -26252 25480 -26247
rect 20352 -26360 20412 -26354
rect 20120 -26500 20180 -26494
rect 26914 -26440 26974 -26018
rect 27376 -26434 27436 -26018
rect 27376 -26500 27436 -26494
rect 27830 -26440 27890 -26018
rect 28292 -26434 28352 -26018
rect 28292 -26500 28352 -26494
rect 28746 -26434 28806 -26018
rect 28746 -26500 28806 -26494
rect 29196 -26434 29256 -26018
rect 29196 -26500 29256 -26494
rect 29662 -26440 29722 -26018
rect 30118 -26434 30178 -26018
rect 30352 -25626 30412 -25620
rect 30352 -25964 30412 -25686
rect 31916 -25964 31976 -25564
rect 32378 -25964 32438 -25556
rect 32826 -25562 32832 -25502
rect 32892 -25562 32898 -25502
rect 33288 -25562 33294 -25502
rect 33354 -25562 33360 -25502
rect 33742 -25562 33748 -25502
rect 33808 -25562 33814 -25502
rect 34192 -25556 34198 -25496
rect 34258 -25556 34264 -25496
rect 32832 -25964 32892 -25562
rect 33294 -25964 33354 -25562
rect 33748 -25964 33808 -25562
rect 34198 -25964 34258 -25556
rect 34658 -25562 34664 -25502
rect 34724 -25562 34730 -25502
rect 35114 -25562 35120 -25502
rect 35180 -25562 35186 -25502
rect 34664 -25964 34724 -25562
rect 35120 -25964 35180 -25562
rect 35346 -25692 35352 -25632
rect 35412 -25692 35418 -25632
rect 30352 -26024 35180 -25964
rect 30352 -26306 30412 -26024
rect 30346 -26366 30352 -26306
rect 30412 -26366 30418 -26306
rect 30118 -26500 30178 -26494
rect 31916 -26434 31976 -26024
rect 31916 -26500 31976 -26494
rect 32378 -26436 32438 -26024
rect 26914 -26506 26974 -26500
rect 27830 -26506 27890 -26500
rect 29662 -26506 29722 -26500
rect 32378 -26502 32438 -26496
rect 32832 -26436 32892 -26024
rect 32832 -26502 32892 -26496
rect 33294 -26436 33354 -26024
rect 33294 -26502 33354 -26496
rect 33748 -26436 33808 -26024
rect 34198 -26430 34258 -26024
rect 34198 -26496 34258 -26490
rect 34664 -26434 34724 -26024
rect 33748 -26502 33808 -26496
rect 34664 -26500 34724 -26494
rect 35120 -26434 35180 -26024
rect 35352 -25968 35412 -25692
rect 35352 -26028 36438 -25968
rect 35352 -26294 35412 -26028
rect 36338 -26157 36438 -26028
rect 40320 -26157 40380 -13646
rect 36334 -26247 36343 -26157
rect 36433 -26247 36442 -26157
rect 40296 -26247 40305 -26157
rect 40395 -26247 40404 -26157
rect 36338 -26252 36438 -26247
rect 40320 -26252 40380 -26247
rect 35352 -26360 35412 -26354
rect 35120 -26500 35180 -26494
rect 25546 -27650 25606 -27644
rect 26914 -27650 26974 -27644
rect 15112 -27710 15118 -27650
rect 15178 -27710 25546 -27650
rect 25606 -27710 26914 -27650
rect 25546 -27716 25606 -27710
rect 26914 -27716 26974 -27710
rect 11160 -27902 20930 -27874
rect 11160 -27988 11210 -27902
rect 11306 -27988 11790 -27902
rect 11886 -27988 12390 -27902
rect 12486 -27988 12990 -27902
rect 13086 -27988 13590 -27902
rect 13686 -27988 14190 -27902
rect 14286 -27988 14790 -27902
rect 14886 -27988 15390 -27902
rect 15486 -27988 15990 -27902
rect 16086 -27988 16590 -27902
rect 16686 -27988 17190 -27902
rect 17286 -27988 17790 -27902
rect 17886 -27988 18390 -27902
rect 18486 -27988 18990 -27902
rect 19086 -27988 19590 -27902
rect 19686 -27988 20190 -27902
rect 20286 -27988 20790 -27902
rect 20886 -27988 20930 -27902
rect 11160 -28018 20930 -27988
rect 26160 -27902 35930 -27874
rect 26160 -27988 26210 -27902
rect 26306 -27988 26790 -27902
rect 26886 -27988 27390 -27902
rect 27486 -27988 27990 -27902
rect 28086 -27988 28590 -27902
rect 28686 -27988 29190 -27902
rect 29286 -27988 29790 -27902
rect 29886 -27988 30390 -27902
rect 30486 -27988 30990 -27902
rect 31086 -27988 31590 -27902
rect 31686 -27988 32190 -27902
rect 32286 -27988 32790 -27902
rect 32886 -27988 33390 -27902
rect 33486 -27988 33990 -27902
rect 34086 -27988 34590 -27902
rect 34686 -27988 35190 -27902
rect 35286 -27988 35790 -27902
rect 35886 -27988 35930 -27902
rect 26160 -28018 35930 -27988
rect 10924 -28166 11524 -28156
rect 10924 -28476 11524 -28466
rect 20556 -28166 21156 -28156
rect 20556 -28476 21156 -28466
rect 25924 -28166 26524 -28156
rect 25924 -28476 26524 -28466
rect 35556 -28166 36156 -28156
rect 35556 -28476 36156 -28466
<< via2 >>
rect 15532 3904 15914 4204
rect 23666 3904 24344 4204
rect 26114 3904 26714 4204
rect 30746 3904 31346 4204
rect 17600 3640 17696 3726
rect 18180 3640 18276 3726
rect 18780 3640 18876 3726
rect 19380 3640 19476 3726
rect 19980 3640 20076 3726
rect 20580 3640 20676 3726
rect 21180 3640 21276 3726
rect 21780 3640 21876 3726
rect 22380 3640 22476 3726
rect 26362 3640 26458 3726
rect 26942 3640 27038 3726
rect 27542 3640 27638 3726
rect 28142 3640 28238 3726
rect 28742 3640 28838 3726
rect 29342 3640 29438 3726
rect 29942 3640 30038 3726
rect 30542 3640 30638 3726
rect 31142 3640 31238 3726
rect 15774 -1078 15870 -992
rect 16374 -1078 16470 -992
rect 16974 -1078 17070 -992
rect 17574 -1078 17670 -992
rect 18174 -1078 18270 -992
rect 18774 -1078 18870 -992
rect 19374 -1078 19470 -992
rect 19974 -1078 20070 -992
rect 20574 -1078 20670 -992
rect 21174 -1078 21270 -992
rect 21774 -1078 21870 -992
rect 22374 -1078 22470 -992
rect 22974 -1078 23070 -992
rect 23574 -1078 23670 -992
rect 23994 -1078 24090 -992
rect 26290 -1078 26386 -992
rect 26890 -1078 26986 -992
rect 27490 -1078 27586 -992
rect 28090 -1078 28186 -992
rect 28690 -1078 28786 -992
rect 29290 -1078 29386 -992
rect 29890 -1078 29986 -992
rect 30490 -1078 30586 -992
rect 31090 -1078 31186 -992
rect 15532 -1552 15914 -1252
rect 23666 -1552 24344 -1252
rect 26114 -1552 26714 -1252
rect 30746 -1552 31346 -1252
rect 10924 -2434 11524 -2134
rect 20556 -2434 21156 -2134
rect 25924 -2434 26524 -2134
rect 35556 -2434 36156 -2134
rect 11776 -2694 11872 -2608
rect 12376 -2694 12472 -2608
rect 12976 -2694 13072 -2608
rect 13576 -2694 13672 -2608
rect 14176 -2694 14272 -2608
rect 14776 -2694 14872 -2608
rect 15376 -2694 15472 -2608
rect 15976 -2694 16072 -2608
rect 16576 -2694 16672 -2608
rect 17176 -2694 17272 -2608
rect 17776 -2694 17872 -2608
rect 18376 -2694 18472 -2608
rect 18976 -2694 19072 -2608
rect 19576 -2694 19672 -2608
rect 19996 -2694 20092 -2608
rect 26776 -2694 26872 -2608
rect 27376 -2694 27472 -2608
rect 27976 -2694 28072 -2608
rect 28576 -2694 28672 -2608
rect 29176 -2694 29272 -2608
rect 29776 -2694 29872 -2608
rect 30376 -2694 30472 -2608
rect 30976 -2694 31072 -2608
rect 31576 -2694 31672 -2608
rect 32176 -2694 32272 -2608
rect 32776 -2694 32872 -2608
rect 33376 -2694 33472 -2608
rect 33976 -2694 34072 -2608
rect 34576 -2694 34672 -2608
rect 34996 -2694 35092 -2608
rect 25616 -8018 25676 -7958
rect 21343 -8247 21433 -8157
rect 36343 -8247 36433 -8157
rect 11210 -9988 11306 -9902
rect 11790 -9988 11886 -9902
rect 12390 -9988 12486 -9902
rect 12990 -9988 13086 -9902
rect 13590 -9988 13686 -9902
rect 14190 -9988 14286 -9902
rect 14790 -9988 14886 -9902
rect 15390 -9988 15486 -9902
rect 15990 -9988 16086 -9902
rect 16590 -9988 16686 -9902
rect 17190 -9988 17286 -9902
rect 17790 -9988 17886 -9902
rect 18390 -9988 18486 -9902
rect 18990 -9988 19086 -9902
rect 19590 -9988 19686 -9902
rect 20190 -9988 20286 -9902
rect 20790 -9988 20886 -9902
rect 26210 -9988 26306 -9902
rect 26790 -9988 26886 -9902
rect 27390 -9988 27486 -9902
rect 27990 -9988 28086 -9902
rect 28590 -9988 28686 -9902
rect 29190 -9988 29286 -9902
rect 29790 -9988 29886 -9902
rect 30390 -9988 30486 -9902
rect 30990 -9988 31086 -9902
rect 31590 -9988 31686 -9902
rect 32190 -9988 32286 -9902
rect 32790 -9988 32886 -9902
rect 33390 -9988 33486 -9902
rect 33990 -9988 34086 -9902
rect 34590 -9988 34686 -9902
rect 35190 -9988 35286 -9902
rect 35790 -9988 35886 -9902
rect 10924 -10466 11524 -10166
rect 20556 -10466 21156 -10166
rect 25924 -10466 26524 -10166
rect 35556 -10466 36156 -10166
rect 14878 -11438 15478 -11138
rect 24510 -11438 25110 -11138
rect 29878 -11438 30478 -11138
rect 39510 -11438 40110 -11138
rect 15148 -11702 15244 -11616
rect 15748 -11702 15844 -11616
rect 16348 -11702 16444 -11616
rect 16948 -11702 17044 -11616
rect 17548 -11702 17644 -11616
rect 18148 -11702 18244 -11616
rect 18748 -11702 18844 -11616
rect 19348 -11702 19444 -11616
rect 19948 -11702 20044 -11616
rect 20548 -11702 20644 -11616
rect 21148 -11702 21244 -11616
rect 21748 -11702 21844 -11616
rect 22348 -11702 22444 -11616
rect 22948 -11702 23044 -11616
rect 23548 -11702 23644 -11616
rect 24148 -11702 24244 -11616
rect 24728 -11702 24824 -11616
rect 30148 -11702 30244 -11616
rect 30748 -11702 30844 -11616
rect 31348 -11702 31444 -11616
rect 31948 -11702 32044 -11616
rect 32548 -11702 32644 -11616
rect 33148 -11702 33244 -11616
rect 33748 -11702 33844 -11616
rect 34348 -11702 34444 -11616
rect 34948 -11702 35044 -11616
rect 35548 -11702 35644 -11616
rect 36148 -11702 36244 -11616
rect 36748 -11702 36844 -11616
rect 37348 -11702 37444 -11616
rect 37948 -11702 38044 -11616
rect 38548 -11702 38644 -11616
rect 39148 -11702 39244 -11616
rect 39728 -11702 39824 -11616
rect 10609 -13447 10699 -13357
rect 14601 -13447 14691 -13357
rect 29601 -13447 29691 -13357
rect 25300 -13646 25360 -13586
rect 15942 -18996 16038 -18910
rect 16362 -18996 16458 -18910
rect 16962 -18996 17058 -18910
rect 17562 -18996 17658 -18910
rect 18162 -18996 18258 -18910
rect 18762 -18996 18858 -18910
rect 19362 -18996 19458 -18910
rect 19962 -18996 20058 -18910
rect 20562 -18996 20658 -18910
rect 21162 -18996 21258 -18910
rect 21762 -18996 21858 -18910
rect 22362 -18996 22458 -18910
rect 22962 -18996 23058 -18910
rect 23562 -18996 23658 -18910
rect 24162 -18996 24258 -18910
rect 30942 -18996 31038 -18910
rect 31362 -18996 31458 -18910
rect 31962 -18996 32058 -18910
rect 32562 -18996 32658 -18910
rect 33162 -18996 33258 -18910
rect 33762 -18996 33858 -18910
rect 34362 -18996 34458 -18910
rect 34962 -18996 35058 -18910
rect 35562 -18996 35658 -18910
rect 36162 -18996 36258 -18910
rect 36762 -18996 36858 -18910
rect 37362 -18996 37458 -18910
rect 37962 -18996 38058 -18910
rect 38562 -18996 38658 -18910
rect 39162 -18996 39258 -18910
rect 14878 -19470 15478 -19170
rect 24510 -19470 25110 -19170
rect 29878 -19470 30478 -19170
rect 39510 -19470 40110 -19170
rect 10924 -20434 11524 -20134
rect 20556 -20434 21156 -20134
rect 25924 -20434 26524 -20134
rect 35556 -20434 36156 -20134
rect 11776 -20694 11872 -20608
rect 12376 -20694 12472 -20608
rect 12976 -20694 13072 -20608
rect 13576 -20694 13672 -20608
rect 14176 -20694 14272 -20608
rect 14776 -20694 14872 -20608
rect 15376 -20694 15472 -20608
rect 15976 -20694 16072 -20608
rect 16576 -20694 16672 -20608
rect 17176 -20694 17272 -20608
rect 17776 -20694 17872 -20608
rect 18376 -20694 18472 -20608
rect 18976 -20694 19072 -20608
rect 19576 -20694 19672 -20608
rect 19996 -20694 20092 -20608
rect 26776 -20694 26872 -20608
rect 27376 -20694 27472 -20608
rect 27976 -20694 28072 -20608
rect 28576 -20694 28672 -20608
rect 29176 -20694 29272 -20608
rect 29776 -20694 29872 -20608
rect 30376 -20694 30472 -20608
rect 30976 -20694 31072 -20608
rect 31576 -20694 31672 -20608
rect 32176 -20694 32272 -20608
rect 32776 -20694 32872 -20608
rect 33376 -20694 33472 -20608
rect 33976 -20694 34072 -20608
rect 34576 -20694 34672 -20608
rect 34996 -20694 35092 -20608
rect 21343 -26247 21433 -26157
rect 25407 -26247 25497 -26157
rect 36343 -26247 36433 -26157
rect 40305 -26247 40395 -26157
rect 11210 -27988 11306 -27902
rect 11790 -27988 11886 -27902
rect 12390 -27988 12486 -27902
rect 12990 -27988 13086 -27902
rect 13590 -27988 13686 -27902
rect 14190 -27988 14286 -27902
rect 14790 -27988 14886 -27902
rect 15390 -27988 15486 -27902
rect 15990 -27988 16086 -27902
rect 16590 -27988 16686 -27902
rect 17190 -27988 17286 -27902
rect 17790 -27988 17886 -27902
rect 18390 -27988 18486 -27902
rect 18990 -27988 19086 -27902
rect 19590 -27988 19686 -27902
rect 20190 -27988 20286 -27902
rect 20790 -27988 20886 -27902
rect 26210 -27988 26306 -27902
rect 26790 -27988 26886 -27902
rect 27390 -27988 27486 -27902
rect 27990 -27988 28086 -27902
rect 28590 -27988 28686 -27902
rect 29190 -27988 29286 -27902
rect 29790 -27988 29886 -27902
rect 30390 -27988 30486 -27902
rect 30990 -27988 31086 -27902
rect 31590 -27988 31686 -27902
rect 32190 -27988 32286 -27902
rect 32790 -27988 32886 -27902
rect 33390 -27988 33486 -27902
rect 33990 -27988 34086 -27902
rect 34590 -27988 34686 -27902
rect 35190 -27988 35286 -27902
rect 35790 -27988 35886 -27902
rect 10924 -28466 11524 -28166
rect 20556 -28466 21156 -28166
rect 25924 -28466 26524 -28166
rect 35556 -28466 36156 -28166
<< metal3 >>
rect 15522 4204 15924 4209
rect 15522 3904 15532 4204
rect 15914 3904 15924 4204
rect 15522 3899 15924 3904
rect 23656 4204 24354 4209
rect 23656 3904 23666 4204
rect 24344 3904 24354 4204
rect 23656 3899 24354 3904
rect 26104 4204 26724 4209
rect 26104 3904 26114 4204
rect 26714 3904 26724 4204
rect 26104 3899 26724 3904
rect 30736 4204 31356 4209
rect 30736 3904 30746 4204
rect 31346 3904 31356 4204
rect 30736 3899 31356 3904
rect 17550 3726 22522 3756
rect 17550 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 22522 3726
rect 17550 3612 22522 3640
rect 26312 3726 31284 3756
rect 26312 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 31284 3726
rect 26312 3612 31284 3640
rect 15760 -992 24116 -982
rect 15760 -1078 15774 -992
rect 15870 -1078 16374 -992
rect 16470 -1078 16974 -992
rect 17070 -1078 17574 -992
rect 17670 -1078 18174 -992
rect 18270 -1078 18774 -992
rect 18870 -1078 19374 -992
rect 19470 -1078 19974 -992
rect 20070 -1078 20574 -992
rect 20670 -1078 21174 -992
rect 21270 -1078 21774 -992
rect 21870 -1078 22374 -992
rect 22470 -1078 22974 -992
rect 23070 -1078 23574 -992
rect 23670 -1078 23994 -992
rect 24090 -1078 24116 -992
rect 15760 -1092 24116 -1078
rect 26276 -992 31274 -982
rect 26276 -1078 26290 -992
rect 26386 -1078 26890 -992
rect 26986 -1078 27490 -992
rect 27586 -1078 28090 -992
rect 28186 -1078 28690 -992
rect 28786 -1078 29290 -992
rect 29386 -1078 29890 -992
rect 29986 -1078 30490 -992
rect 30586 -1078 31090 -992
rect 31186 -1078 31274 -992
rect 26276 -1092 31274 -1078
rect 15522 -1252 15924 -1247
rect 15522 -1552 15532 -1252
rect 15914 -1552 15924 -1252
rect 15522 -1557 15924 -1552
rect 23656 -1252 24354 -1247
rect 23656 -1552 23666 -1252
rect 24344 -1552 24354 -1252
rect 23656 -1557 24354 -1552
rect 26104 -1252 26724 -1247
rect 26104 -1552 26114 -1252
rect 26714 -1552 26724 -1252
rect 26104 -1557 26724 -1552
rect 30736 -1252 31356 -1247
rect 30736 -1552 30746 -1252
rect 31346 -1552 31356 -1252
rect 30736 -1557 31356 -1552
rect 10914 -2134 11534 -2129
rect 10914 -2434 10924 -2134
rect 11524 -2434 11534 -2134
rect 10914 -2439 11534 -2434
rect 20546 -2134 21166 -2129
rect 20546 -2434 20556 -2134
rect 21156 -2434 21166 -2134
rect 20546 -2439 21166 -2434
rect 25914 -2134 26534 -2129
rect 25914 -2434 25924 -2134
rect 26524 -2434 26534 -2134
rect 25914 -2439 26534 -2434
rect 35546 -2134 36166 -2129
rect 35546 -2434 35556 -2134
rect 36156 -2434 36166 -2134
rect 35546 -2439 36166 -2434
rect 11762 -2608 20118 -2594
rect 11762 -2694 11776 -2608
rect 11872 -2694 12376 -2608
rect 12472 -2694 12976 -2608
rect 13072 -2694 13576 -2608
rect 13672 -2694 14176 -2608
rect 14272 -2694 14776 -2608
rect 14872 -2694 15376 -2608
rect 15472 -2694 15976 -2608
rect 16072 -2694 16576 -2608
rect 16672 -2694 17176 -2608
rect 17272 -2694 17776 -2608
rect 17872 -2694 18376 -2608
rect 18472 -2694 18976 -2608
rect 19072 -2694 19576 -2608
rect 19672 -2694 19996 -2608
rect 20092 -2694 20118 -2608
rect 11762 -2704 20118 -2694
rect 26762 -2608 35118 -2594
rect 26762 -2694 26776 -2608
rect 26872 -2694 27376 -2608
rect 27472 -2694 27976 -2608
rect 28072 -2694 28576 -2608
rect 28672 -2694 29176 -2608
rect 29272 -2694 29776 -2608
rect 29872 -2694 30376 -2608
rect 30472 -2694 30976 -2608
rect 31072 -2694 31576 -2608
rect 31672 -2694 32176 -2608
rect 32272 -2694 32776 -2608
rect 32872 -2694 33376 -2608
rect 33472 -2694 33976 -2608
rect 34072 -2694 34576 -2608
rect 34672 -2694 34996 -2608
rect 35092 -2694 35118 -2608
rect 26762 -2704 35118 -2694
rect 21538 -6966 25166 -6832
rect 21538 -7338 22175 -6966
rect 22239 -6968 25166 -6966
rect 22239 -7338 22894 -6968
rect 22958 -7338 23613 -6968
rect 23677 -7338 24332 -6968
rect 24396 -7338 25051 -6968
rect 25115 -7338 25166 -6968
rect 21538 -7668 25166 -7338
rect 21538 -8036 22175 -7668
rect 22239 -8036 22894 -7668
rect 22958 -8036 23613 -7668
rect 23677 -8036 24332 -7668
rect 24396 -8036 25051 -7668
rect 25115 -8036 25166 -7668
rect 36538 -6966 40166 -6832
rect 36538 -7338 37175 -6966
rect 37239 -6968 40166 -6966
rect 37239 -7338 37894 -6968
rect 37958 -7338 38613 -6968
rect 38677 -7338 39332 -6968
rect 39396 -7338 40051 -6968
rect 40115 -7338 40166 -6968
rect 36538 -7668 40166 -7338
rect 25611 -7958 25681 -7953
rect 21338 -8153 21438 -8152
rect 21333 -8251 21339 -8153
rect 21437 -8251 21443 -8153
rect 21338 -8252 21438 -8251
rect 21538 -8368 25166 -8036
rect 25596 -8018 25616 -7958
rect 25676 -8018 25696 -7958
rect 25272 -8153 25372 -8152
rect 25267 -8251 25273 -8153
rect 25371 -8251 25377 -8153
rect 21538 -8736 22175 -8368
rect 22239 -8736 22894 -8368
rect 22958 -8736 23613 -8368
rect 23677 -8736 24332 -8368
rect 24396 -8736 25051 -8368
rect 25115 -8736 25166 -8368
rect 21538 -9068 25166 -8736
rect 21538 -9436 22175 -9068
rect 22239 -9436 22894 -9068
rect 22958 -9436 23613 -9068
rect 23677 -9436 24332 -9068
rect 24396 -9436 25051 -9068
rect 25115 -9436 25166 -9068
rect 21538 -9768 25166 -9436
rect 11160 -9902 20930 -9874
rect 11160 -9988 11210 -9902
rect 11306 -9988 11790 -9902
rect 11886 -9988 12390 -9902
rect 12486 -9988 12990 -9902
rect 13086 -9988 13590 -9902
rect 13686 -9988 14190 -9902
rect 14286 -9988 14790 -9902
rect 14886 -9988 15390 -9902
rect 15486 -9988 15990 -9902
rect 16086 -9988 16590 -9902
rect 16686 -9988 17190 -9902
rect 17286 -9988 17790 -9902
rect 17886 -9988 18390 -9902
rect 18486 -9988 18990 -9902
rect 19086 -9988 19590 -9902
rect 19686 -9988 20190 -9902
rect 20286 -9988 20790 -9902
rect 20886 -9988 20930 -9902
rect 11160 -10018 20930 -9988
rect 21538 -10136 22175 -9768
rect 22239 -10136 22894 -9768
rect 22958 -10136 23613 -9768
rect 23677 -10136 24332 -9768
rect 24396 -10136 25051 -9768
rect 25115 -10136 25166 -9768
rect 10914 -10166 11534 -10161
rect 10914 -10466 10924 -10166
rect 11524 -10466 11534 -10166
rect 10914 -10471 11534 -10466
rect 20546 -10166 21166 -10161
rect 20546 -10466 20556 -10166
rect 21156 -10466 21166 -10166
rect 21538 -10286 25166 -10136
rect 20546 -10471 21166 -10466
rect 14868 -11138 15488 -11133
rect 10868 -11468 14496 -11318
rect 14868 -11438 14878 -11138
rect 15478 -11438 15488 -11138
rect 14868 -11443 15488 -11438
rect 24500 -11138 25120 -11133
rect 24500 -11438 24510 -11138
rect 25110 -11438 25120 -11138
rect 24500 -11443 25120 -11438
rect 10868 -11836 10919 -11468
rect 10983 -11836 11638 -11468
rect 11702 -11836 12357 -11468
rect 12421 -11836 13076 -11468
rect 13140 -11836 13795 -11468
rect 13859 -11836 14496 -11468
rect 15104 -11616 24874 -11586
rect 15104 -11702 15148 -11616
rect 15244 -11702 15748 -11616
rect 15844 -11702 16348 -11616
rect 16444 -11702 16948 -11616
rect 17044 -11702 17548 -11616
rect 17644 -11702 18148 -11616
rect 18244 -11702 18748 -11616
rect 18844 -11702 19348 -11616
rect 19444 -11702 19948 -11616
rect 20044 -11702 20548 -11616
rect 20644 -11702 21148 -11616
rect 21244 -11702 21748 -11616
rect 21844 -11702 22348 -11616
rect 22444 -11702 22948 -11616
rect 23044 -11702 23548 -11616
rect 23644 -11702 24148 -11616
rect 24244 -11702 24728 -11616
rect 24824 -11702 24874 -11616
rect 15104 -11730 24874 -11702
rect 10868 -12168 14496 -11836
rect 10868 -12536 10919 -12168
rect 10983 -12536 11638 -12168
rect 11702 -12536 12357 -12168
rect 12421 -12536 13076 -12168
rect 13140 -12536 13795 -12168
rect 13859 -12536 14496 -12168
rect 10868 -12868 14496 -12536
rect 10868 -13236 10919 -12868
rect 10983 -13236 11638 -12868
rect 11702 -13236 12357 -12868
rect 12421 -13236 13076 -12868
rect 13140 -13236 13795 -12868
rect 13859 -13236 14496 -12868
rect 10604 -13353 10704 -13352
rect 10599 -13451 10605 -13353
rect 10703 -13451 10709 -13353
rect 10604 -13452 10704 -13451
rect 10868 -13568 14496 -13236
rect 14596 -13353 14696 -13352
rect 14591 -13451 14597 -13353
rect 14695 -13451 14701 -13353
rect 14596 -13452 14696 -13451
rect 10868 -13936 10919 -13568
rect 10983 -13936 11638 -13568
rect 11702 -13936 12357 -13568
rect 12421 -13936 13076 -13568
rect 13140 -13936 13795 -13568
rect 13859 -13936 14496 -13568
rect 25272 -13586 25372 -8251
rect 25596 -13353 25696 -8018
rect 36538 -8036 37175 -7668
rect 37239 -8036 37894 -7668
rect 37958 -8036 38613 -7668
rect 38677 -8036 39332 -7668
rect 39396 -8036 40051 -7668
rect 40115 -8036 40166 -7668
rect 36338 -8153 36438 -8152
rect 36333 -8251 36339 -8153
rect 36437 -8251 36443 -8153
rect 36338 -8252 36438 -8251
rect 36538 -8368 40166 -8036
rect 36538 -8736 37175 -8368
rect 37239 -8736 37894 -8368
rect 37958 -8736 38613 -8368
rect 38677 -8736 39332 -8368
rect 39396 -8736 40051 -8368
rect 40115 -8736 40166 -8368
rect 36538 -9068 40166 -8736
rect 36538 -9436 37175 -9068
rect 37239 -9436 37894 -9068
rect 37958 -9436 38613 -9068
rect 38677 -9436 39332 -9068
rect 39396 -9436 40051 -9068
rect 40115 -9436 40166 -9068
rect 36538 -9768 40166 -9436
rect 26160 -9902 35930 -9874
rect 26160 -9988 26210 -9902
rect 26306 -9988 26790 -9902
rect 26886 -9988 27390 -9902
rect 27486 -9988 27990 -9902
rect 28086 -9988 28590 -9902
rect 28686 -9988 29190 -9902
rect 29286 -9988 29790 -9902
rect 29886 -9988 30390 -9902
rect 30486 -9988 30990 -9902
rect 31086 -9988 31590 -9902
rect 31686 -9988 32190 -9902
rect 32286 -9988 32790 -9902
rect 32886 -9988 33390 -9902
rect 33486 -9988 33990 -9902
rect 34086 -9988 34590 -9902
rect 34686 -9988 35190 -9902
rect 35286 -9988 35790 -9902
rect 35886 -9988 35930 -9902
rect 26160 -10018 35930 -9988
rect 36538 -10136 37175 -9768
rect 37239 -10136 37894 -9768
rect 37958 -10136 38613 -9768
rect 38677 -10136 39332 -9768
rect 39396 -10136 40051 -9768
rect 40115 -10136 40166 -9768
rect 25914 -10166 26534 -10161
rect 25914 -10466 25924 -10166
rect 26524 -10466 26534 -10166
rect 25914 -10471 26534 -10466
rect 35546 -10166 36166 -10161
rect 35546 -10466 35556 -10166
rect 36156 -10466 36166 -10166
rect 36538 -10286 40166 -10136
rect 35546 -10471 36166 -10466
rect 29868 -11138 30488 -11133
rect 25868 -11468 29496 -11318
rect 29868 -11438 29878 -11138
rect 30478 -11438 30488 -11138
rect 29868 -11443 30488 -11438
rect 39500 -11138 40120 -11133
rect 39500 -11438 39510 -11138
rect 40110 -11438 40120 -11138
rect 39500 -11443 40120 -11438
rect 25868 -11836 25919 -11468
rect 25983 -11836 26638 -11468
rect 26702 -11836 27357 -11468
rect 27421 -11836 28076 -11468
rect 28140 -11836 28795 -11468
rect 28859 -11836 29496 -11468
rect 30104 -11616 39874 -11586
rect 30104 -11702 30148 -11616
rect 30244 -11702 30748 -11616
rect 30844 -11702 31348 -11616
rect 31444 -11702 31948 -11616
rect 32044 -11702 32548 -11616
rect 32644 -11702 33148 -11616
rect 33244 -11702 33748 -11616
rect 33844 -11702 34348 -11616
rect 34444 -11702 34948 -11616
rect 35044 -11702 35548 -11616
rect 35644 -11702 36148 -11616
rect 36244 -11702 36748 -11616
rect 36844 -11702 37348 -11616
rect 37444 -11702 37948 -11616
rect 38044 -11702 38548 -11616
rect 38644 -11702 39148 -11616
rect 39244 -11702 39728 -11616
rect 39824 -11702 39874 -11616
rect 30104 -11730 39874 -11702
rect 25868 -12168 29496 -11836
rect 25868 -12536 25919 -12168
rect 25983 -12536 26638 -12168
rect 26702 -12536 27357 -12168
rect 27421 -12536 28076 -12168
rect 28140 -12536 28795 -12168
rect 28859 -12536 29496 -12168
rect 25868 -12868 29496 -12536
rect 25868 -13236 25919 -12868
rect 25983 -13236 26638 -12868
rect 26702 -13236 27357 -12868
rect 27421 -13236 28076 -12868
rect 28140 -13236 28795 -12868
rect 28859 -13236 29496 -12868
rect 25591 -13451 25597 -13353
rect 25695 -13451 25701 -13353
rect 25596 -13452 25696 -13451
rect 25272 -13646 25300 -13586
rect 25360 -13646 25372 -13586
rect 25272 -13662 25372 -13646
rect 25868 -13568 29496 -13236
rect 29596 -13353 29696 -13352
rect 29591 -13451 29597 -13353
rect 29695 -13451 29701 -13353
rect 29596 -13452 29696 -13451
rect 10868 -14266 14496 -13936
rect 10868 -14636 10919 -14266
rect 10983 -14636 11638 -14266
rect 11702 -14636 12357 -14266
rect 12421 -14636 13076 -14266
rect 13140 -14636 13795 -14266
rect 10868 -14638 13795 -14636
rect 13859 -14638 14496 -14266
rect 10868 -14772 14496 -14638
rect 25868 -13936 25919 -13568
rect 25983 -13936 26638 -13568
rect 26702 -13936 27357 -13568
rect 27421 -13936 28076 -13568
rect 28140 -13936 28795 -13568
rect 28859 -13936 29496 -13568
rect 25868 -14266 29496 -13936
rect 25868 -14636 25919 -14266
rect 25983 -14636 26638 -14266
rect 26702 -14636 27357 -14266
rect 27421 -14636 28076 -14266
rect 28140 -14636 28795 -14266
rect 25868 -14638 28795 -14636
rect 28859 -14638 29496 -14266
rect 25868 -14772 29496 -14638
rect 15916 -18910 24272 -18900
rect 15916 -18996 15942 -18910
rect 16038 -18996 16362 -18910
rect 16458 -18996 16962 -18910
rect 17058 -18996 17562 -18910
rect 17658 -18996 18162 -18910
rect 18258 -18996 18762 -18910
rect 18858 -18996 19362 -18910
rect 19458 -18996 19962 -18910
rect 20058 -18996 20562 -18910
rect 20658 -18996 21162 -18910
rect 21258 -18996 21762 -18910
rect 21858 -18996 22362 -18910
rect 22458 -18996 22962 -18910
rect 23058 -18996 23562 -18910
rect 23658 -18996 24162 -18910
rect 24258 -18996 24272 -18910
rect 15916 -19010 24272 -18996
rect 30916 -18910 39272 -18900
rect 30916 -18996 30942 -18910
rect 31038 -18996 31362 -18910
rect 31458 -18996 31962 -18910
rect 32058 -18996 32562 -18910
rect 32658 -18996 33162 -18910
rect 33258 -18996 33762 -18910
rect 33858 -18996 34362 -18910
rect 34458 -18996 34962 -18910
rect 35058 -18996 35562 -18910
rect 35658 -18996 36162 -18910
rect 36258 -18996 36762 -18910
rect 36858 -18996 37362 -18910
rect 37458 -18996 37962 -18910
rect 38058 -18996 38562 -18910
rect 38658 -18996 39162 -18910
rect 39258 -18996 39272 -18910
rect 30916 -19010 39272 -18996
rect 14868 -19170 15488 -19165
rect 14868 -19470 14878 -19170
rect 15478 -19470 15488 -19170
rect 14868 -19475 15488 -19470
rect 24500 -19170 25120 -19165
rect 24500 -19470 24510 -19170
rect 25110 -19470 25120 -19170
rect 24500 -19475 25120 -19470
rect 29868 -19170 30488 -19165
rect 29868 -19470 29878 -19170
rect 30478 -19470 30488 -19170
rect 29868 -19475 30488 -19470
rect 39500 -19170 40120 -19165
rect 39500 -19470 39510 -19170
rect 40110 -19470 40120 -19170
rect 39500 -19475 40120 -19470
rect 10914 -20134 11534 -20129
rect 10914 -20434 10924 -20134
rect 11524 -20434 11534 -20134
rect 10914 -20439 11534 -20434
rect 20546 -20134 21166 -20129
rect 20546 -20434 20556 -20134
rect 21156 -20434 21166 -20134
rect 20546 -20439 21166 -20434
rect 25914 -20134 26534 -20129
rect 25914 -20434 25924 -20134
rect 26524 -20434 26534 -20134
rect 25914 -20439 26534 -20434
rect 35546 -20134 36166 -20129
rect 35546 -20434 35556 -20134
rect 36156 -20434 36166 -20134
rect 35546 -20439 36166 -20434
rect 11762 -20608 20118 -20594
rect 11762 -20694 11776 -20608
rect 11872 -20694 12376 -20608
rect 12472 -20694 12976 -20608
rect 13072 -20694 13576 -20608
rect 13672 -20694 14176 -20608
rect 14272 -20694 14776 -20608
rect 14872 -20694 15376 -20608
rect 15472 -20694 15976 -20608
rect 16072 -20694 16576 -20608
rect 16672 -20694 17176 -20608
rect 17272 -20694 17776 -20608
rect 17872 -20694 18376 -20608
rect 18472 -20694 18976 -20608
rect 19072 -20694 19576 -20608
rect 19672 -20694 19996 -20608
rect 20092 -20694 20118 -20608
rect 11762 -20704 20118 -20694
rect 26762 -20608 35118 -20594
rect 26762 -20694 26776 -20608
rect 26872 -20694 27376 -20608
rect 27472 -20694 27976 -20608
rect 28072 -20694 28576 -20608
rect 28672 -20694 29176 -20608
rect 29272 -20694 29776 -20608
rect 29872 -20694 30376 -20608
rect 30472 -20694 30976 -20608
rect 31072 -20694 31576 -20608
rect 31672 -20694 32176 -20608
rect 32272 -20694 32776 -20608
rect 32872 -20694 33376 -20608
rect 33472 -20694 33976 -20608
rect 34072 -20694 34576 -20608
rect 34672 -20694 34996 -20608
rect 35092 -20694 35118 -20608
rect 26762 -20704 35118 -20694
rect 21538 -24966 25166 -24832
rect 21538 -25338 22175 -24966
rect 22239 -24968 25166 -24966
rect 22239 -25338 22894 -24968
rect 22958 -25338 23613 -24968
rect 23677 -25338 24332 -24968
rect 24396 -25338 25051 -24968
rect 25115 -25338 25166 -24968
rect 21538 -25668 25166 -25338
rect 21538 -26036 22175 -25668
rect 22239 -26036 22894 -25668
rect 22958 -26036 23613 -25668
rect 23677 -26036 24332 -25668
rect 24396 -26036 25051 -25668
rect 25115 -26036 25166 -25668
rect 21338 -26153 21438 -26152
rect 21333 -26251 21339 -26153
rect 21437 -26251 21443 -26153
rect 21338 -26252 21438 -26251
rect 21538 -26368 25166 -26036
rect 36538 -24966 40166 -24832
rect 36538 -25338 37175 -24966
rect 37239 -24968 40166 -24966
rect 37239 -25338 37894 -24968
rect 37958 -25338 38613 -24968
rect 38677 -25338 39332 -24968
rect 39396 -25338 40051 -24968
rect 40115 -25338 40166 -24968
rect 36538 -25668 40166 -25338
rect 36538 -26036 37175 -25668
rect 37239 -26036 37894 -25668
rect 37958 -26036 38613 -25668
rect 38677 -26036 39332 -25668
rect 39396 -26036 40051 -25668
rect 40115 -26036 40166 -25668
rect 25402 -26153 25502 -26152
rect 36338 -26153 36438 -26152
rect 25397 -26251 25403 -26153
rect 25501 -26251 25507 -26153
rect 36333 -26251 36339 -26153
rect 36437 -26251 36443 -26153
rect 25402 -26252 25502 -26251
rect 36338 -26252 36438 -26251
rect 21538 -26736 22175 -26368
rect 22239 -26736 22894 -26368
rect 22958 -26736 23613 -26368
rect 23677 -26736 24332 -26368
rect 24396 -26736 25051 -26368
rect 25115 -26736 25166 -26368
rect 21538 -27068 25166 -26736
rect 21538 -27436 22175 -27068
rect 22239 -27436 22894 -27068
rect 22958 -27436 23613 -27068
rect 23677 -27436 24332 -27068
rect 24396 -27436 25051 -27068
rect 25115 -27436 25166 -27068
rect 21538 -27768 25166 -27436
rect 11160 -27902 20930 -27874
rect 11160 -27988 11210 -27902
rect 11306 -27988 11790 -27902
rect 11886 -27988 12390 -27902
rect 12486 -27988 12990 -27902
rect 13086 -27988 13590 -27902
rect 13686 -27988 14190 -27902
rect 14286 -27988 14790 -27902
rect 14886 -27988 15390 -27902
rect 15486 -27988 15990 -27902
rect 16086 -27988 16590 -27902
rect 16686 -27988 17190 -27902
rect 17286 -27988 17790 -27902
rect 17886 -27988 18390 -27902
rect 18486 -27988 18990 -27902
rect 19086 -27988 19590 -27902
rect 19686 -27988 20190 -27902
rect 20286 -27988 20790 -27902
rect 20886 -27988 20930 -27902
rect 11160 -28018 20930 -27988
rect 21538 -28136 22175 -27768
rect 22239 -28136 22894 -27768
rect 22958 -28136 23613 -27768
rect 23677 -28136 24332 -27768
rect 24396 -28136 25051 -27768
rect 25115 -28136 25166 -27768
rect 36538 -26368 40166 -26036
rect 40300 -26153 40400 -26152
rect 40295 -26251 40301 -26153
rect 40399 -26251 40405 -26153
rect 40300 -26252 40400 -26251
rect 36538 -26736 37175 -26368
rect 37239 -26736 37894 -26368
rect 37958 -26736 38613 -26368
rect 38677 -26736 39332 -26368
rect 39396 -26736 40051 -26368
rect 40115 -26736 40166 -26368
rect 36538 -27068 40166 -26736
rect 36538 -27436 37175 -27068
rect 37239 -27436 37894 -27068
rect 37958 -27436 38613 -27068
rect 38677 -27436 39332 -27068
rect 39396 -27436 40051 -27068
rect 40115 -27436 40166 -27068
rect 36538 -27768 40166 -27436
rect 26160 -27902 35930 -27874
rect 26160 -27988 26210 -27902
rect 26306 -27988 26790 -27902
rect 26886 -27988 27390 -27902
rect 27486 -27988 27990 -27902
rect 28086 -27988 28590 -27902
rect 28686 -27988 29190 -27902
rect 29286 -27988 29790 -27902
rect 29886 -27988 30390 -27902
rect 30486 -27988 30990 -27902
rect 31086 -27988 31590 -27902
rect 31686 -27988 32190 -27902
rect 32286 -27988 32790 -27902
rect 32886 -27988 33390 -27902
rect 33486 -27988 33990 -27902
rect 34086 -27988 34590 -27902
rect 34686 -27988 35190 -27902
rect 35286 -27988 35790 -27902
rect 35886 -27988 35930 -27902
rect 26160 -28018 35930 -27988
rect 10914 -28166 11534 -28161
rect 10914 -28466 10924 -28166
rect 11524 -28466 11534 -28166
rect 10914 -28471 11534 -28466
rect 20546 -28166 21166 -28161
rect 20546 -28466 20556 -28166
rect 21156 -28466 21166 -28166
rect 21538 -28286 25166 -28136
rect 36538 -28136 37175 -27768
rect 37239 -28136 37894 -27768
rect 37958 -28136 38613 -27768
rect 38677 -28136 39332 -27768
rect 39396 -28136 40051 -27768
rect 40115 -28136 40166 -27768
rect 25914 -28166 26534 -28161
rect 20546 -28471 21166 -28466
rect 25914 -28466 25924 -28166
rect 26524 -28466 26534 -28166
rect 25914 -28471 26534 -28466
rect 35546 -28166 36166 -28161
rect 35546 -28466 35556 -28166
rect 36156 -28466 36166 -28166
rect 36538 -28286 40166 -28136
rect 35546 -28471 36166 -28466
<< via3 >>
rect 15532 3904 15914 4204
rect 23666 3904 24344 4204
rect 26114 3904 26714 4204
rect 30746 3904 31346 4204
rect 17600 3640 17696 3726
rect 18180 3640 18276 3726
rect 18780 3640 18876 3726
rect 19380 3640 19476 3726
rect 19980 3640 20076 3726
rect 20580 3640 20676 3726
rect 21180 3640 21276 3726
rect 21780 3640 21876 3726
rect 22380 3640 22476 3726
rect 26362 3640 26458 3726
rect 26942 3640 27038 3726
rect 27542 3640 27638 3726
rect 28142 3640 28238 3726
rect 28742 3640 28838 3726
rect 29342 3640 29438 3726
rect 29942 3640 30038 3726
rect 30542 3640 30638 3726
rect 31142 3640 31238 3726
rect 15532 -1552 15914 -1252
rect 23666 -1552 24344 -1252
rect 26114 -1552 26714 -1252
rect 30746 -1552 31346 -1252
rect 10924 -2434 11524 -2134
rect 20556 -2434 21156 -2134
rect 25924 -2434 26524 -2134
rect 35556 -2434 36156 -2134
rect 11776 -2694 11872 -2608
rect 12376 -2694 12472 -2608
rect 12976 -2694 13072 -2608
rect 13576 -2694 13672 -2608
rect 14176 -2694 14272 -2608
rect 14776 -2694 14872 -2608
rect 15376 -2694 15472 -2608
rect 15976 -2694 16072 -2608
rect 16576 -2694 16672 -2608
rect 17176 -2694 17272 -2608
rect 17776 -2694 17872 -2608
rect 18376 -2694 18472 -2608
rect 18976 -2694 19072 -2608
rect 19576 -2694 19672 -2608
rect 19996 -2694 20092 -2608
rect 26776 -2694 26872 -2608
rect 27376 -2694 27472 -2608
rect 27976 -2694 28072 -2608
rect 28576 -2694 28672 -2608
rect 29176 -2694 29272 -2608
rect 29776 -2694 29872 -2608
rect 30376 -2694 30472 -2608
rect 30976 -2694 31072 -2608
rect 31576 -2694 31672 -2608
rect 32176 -2694 32272 -2608
rect 32776 -2694 32872 -2608
rect 33376 -2694 33472 -2608
rect 33976 -2694 34072 -2608
rect 34576 -2694 34672 -2608
rect 34996 -2694 35092 -2608
rect 22175 -7338 22239 -6966
rect 22894 -7338 22958 -6968
rect 23613 -7338 23677 -6968
rect 24332 -7338 24396 -6968
rect 25051 -7338 25115 -6968
rect 22175 -8036 22239 -7668
rect 22894 -8036 22958 -7668
rect 23613 -8036 23677 -7668
rect 24332 -8036 24396 -7668
rect 25051 -8036 25115 -7668
rect 37175 -7338 37239 -6966
rect 37894 -7338 37958 -6968
rect 38613 -7338 38677 -6968
rect 39332 -7338 39396 -6968
rect 40051 -7338 40115 -6968
rect 21339 -8157 21437 -8153
rect 21339 -8247 21343 -8157
rect 21343 -8247 21433 -8157
rect 21433 -8247 21437 -8157
rect 21339 -8251 21437 -8247
rect 25273 -8251 25371 -8153
rect 22175 -8736 22239 -8368
rect 22894 -8736 22958 -8368
rect 23613 -8736 23677 -8368
rect 24332 -8736 24396 -8368
rect 25051 -8736 25115 -8368
rect 22175 -9436 22239 -9068
rect 22894 -9436 22958 -9068
rect 23613 -9436 23677 -9068
rect 24332 -9436 24396 -9068
rect 25051 -9436 25115 -9068
rect 11210 -9988 11306 -9902
rect 11790 -9988 11886 -9902
rect 12390 -9988 12486 -9902
rect 12990 -9988 13086 -9902
rect 13590 -9988 13686 -9902
rect 14190 -9988 14286 -9902
rect 14790 -9988 14886 -9902
rect 15390 -9988 15486 -9902
rect 15990 -9988 16086 -9902
rect 16590 -9988 16686 -9902
rect 17190 -9988 17286 -9902
rect 17790 -9988 17886 -9902
rect 18390 -9988 18486 -9902
rect 18990 -9988 19086 -9902
rect 19590 -9988 19686 -9902
rect 20190 -9988 20286 -9902
rect 20790 -9988 20886 -9902
rect 22175 -10136 22239 -9768
rect 22894 -10136 22958 -9768
rect 23613 -10136 23677 -9768
rect 24332 -10136 24396 -9768
rect 25051 -10136 25115 -9768
rect 10924 -10466 11524 -10166
rect 20556 -10466 21156 -10166
rect 14878 -11438 15478 -11138
rect 24510 -11438 25110 -11138
rect 10919 -11836 10983 -11468
rect 11638 -11836 11702 -11468
rect 12357 -11836 12421 -11468
rect 13076 -11836 13140 -11468
rect 13795 -11836 13859 -11468
rect 15148 -11702 15244 -11616
rect 15748 -11702 15844 -11616
rect 16348 -11702 16444 -11616
rect 16948 -11702 17044 -11616
rect 17548 -11702 17644 -11616
rect 18148 -11702 18244 -11616
rect 18748 -11702 18844 -11616
rect 19348 -11702 19444 -11616
rect 19948 -11702 20044 -11616
rect 20548 -11702 20644 -11616
rect 21148 -11702 21244 -11616
rect 21748 -11702 21844 -11616
rect 22348 -11702 22444 -11616
rect 22948 -11702 23044 -11616
rect 23548 -11702 23644 -11616
rect 24148 -11702 24244 -11616
rect 24728 -11702 24824 -11616
rect 10919 -12536 10983 -12168
rect 11638 -12536 11702 -12168
rect 12357 -12536 12421 -12168
rect 13076 -12536 13140 -12168
rect 13795 -12536 13859 -12168
rect 10919 -13236 10983 -12868
rect 11638 -13236 11702 -12868
rect 12357 -13236 12421 -12868
rect 13076 -13236 13140 -12868
rect 13795 -13236 13859 -12868
rect 10605 -13357 10703 -13353
rect 10605 -13447 10609 -13357
rect 10609 -13447 10699 -13357
rect 10699 -13447 10703 -13357
rect 10605 -13451 10703 -13447
rect 14597 -13357 14695 -13353
rect 14597 -13447 14601 -13357
rect 14601 -13447 14691 -13357
rect 14691 -13447 14695 -13357
rect 14597 -13451 14695 -13447
rect 10919 -13936 10983 -13568
rect 11638 -13936 11702 -13568
rect 12357 -13936 12421 -13568
rect 13076 -13936 13140 -13568
rect 13795 -13936 13859 -13568
rect 37175 -8036 37239 -7668
rect 37894 -8036 37958 -7668
rect 38613 -8036 38677 -7668
rect 39332 -8036 39396 -7668
rect 40051 -8036 40115 -7668
rect 36339 -8157 36437 -8153
rect 36339 -8247 36343 -8157
rect 36343 -8247 36433 -8157
rect 36433 -8247 36437 -8157
rect 36339 -8251 36437 -8247
rect 37175 -8736 37239 -8368
rect 37894 -8736 37958 -8368
rect 38613 -8736 38677 -8368
rect 39332 -8736 39396 -8368
rect 40051 -8736 40115 -8368
rect 37175 -9436 37239 -9068
rect 37894 -9436 37958 -9068
rect 38613 -9436 38677 -9068
rect 39332 -9436 39396 -9068
rect 40051 -9436 40115 -9068
rect 26210 -9988 26306 -9902
rect 26790 -9988 26886 -9902
rect 27390 -9988 27486 -9902
rect 27990 -9988 28086 -9902
rect 28590 -9988 28686 -9902
rect 29190 -9988 29286 -9902
rect 29790 -9988 29886 -9902
rect 30390 -9988 30486 -9902
rect 30990 -9988 31086 -9902
rect 31590 -9988 31686 -9902
rect 32190 -9988 32286 -9902
rect 32790 -9988 32886 -9902
rect 33390 -9988 33486 -9902
rect 33990 -9988 34086 -9902
rect 34590 -9988 34686 -9902
rect 35190 -9988 35286 -9902
rect 35790 -9988 35886 -9902
rect 37175 -10136 37239 -9768
rect 37894 -10136 37958 -9768
rect 38613 -10136 38677 -9768
rect 39332 -10136 39396 -9768
rect 40051 -10136 40115 -9768
rect 25924 -10466 26524 -10166
rect 35556 -10466 36156 -10166
rect 29878 -11438 30478 -11138
rect 39510 -11438 40110 -11138
rect 25919 -11836 25983 -11468
rect 26638 -11836 26702 -11468
rect 27357 -11836 27421 -11468
rect 28076 -11836 28140 -11468
rect 28795 -11836 28859 -11468
rect 30148 -11702 30244 -11616
rect 30748 -11702 30844 -11616
rect 31348 -11702 31444 -11616
rect 31948 -11702 32044 -11616
rect 32548 -11702 32644 -11616
rect 33148 -11702 33244 -11616
rect 33748 -11702 33844 -11616
rect 34348 -11702 34444 -11616
rect 34948 -11702 35044 -11616
rect 35548 -11702 35644 -11616
rect 36148 -11702 36244 -11616
rect 36748 -11702 36844 -11616
rect 37348 -11702 37444 -11616
rect 37948 -11702 38044 -11616
rect 38548 -11702 38644 -11616
rect 39148 -11702 39244 -11616
rect 39728 -11702 39824 -11616
rect 25919 -12536 25983 -12168
rect 26638 -12536 26702 -12168
rect 27357 -12536 27421 -12168
rect 28076 -12536 28140 -12168
rect 28795 -12536 28859 -12168
rect 25919 -13236 25983 -12868
rect 26638 -13236 26702 -12868
rect 27357 -13236 27421 -12868
rect 28076 -13236 28140 -12868
rect 28795 -13236 28859 -12868
rect 25597 -13451 25695 -13353
rect 29597 -13357 29695 -13353
rect 29597 -13447 29601 -13357
rect 29601 -13447 29691 -13357
rect 29691 -13447 29695 -13357
rect 29597 -13451 29695 -13447
rect 10919 -14636 10983 -14266
rect 11638 -14636 11702 -14266
rect 12357 -14636 12421 -14266
rect 13076 -14636 13140 -14266
rect 13795 -14638 13859 -14266
rect 25919 -13936 25983 -13568
rect 26638 -13936 26702 -13568
rect 27357 -13936 27421 -13568
rect 28076 -13936 28140 -13568
rect 28795 -13936 28859 -13568
rect 25919 -14636 25983 -14266
rect 26638 -14636 26702 -14266
rect 27357 -14636 27421 -14266
rect 28076 -14636 28140 -14266
rect 28795 -14638 28859 -14266
rect 15942 -18996 16038 -18910
rect 16362 -18996 16458 -18910
rect 16962 -18996 17058 -18910
rect 17562 -18996 17658 -18910
rect 18162 -18996 18258 -18910
rect 18762 -18996 18858 -18910
rect 19362 -18996 19458 -18910
rect 19962 -18996 20058 -18910
rect 20562 -18996 20658 -18910
rect 21162 -18996 21258 -18910
rect 21762 -18996 21858 -18910
rect 22362 -18996 22458 -18910
rect 22962 -18996 23058 -18910
rect 23562 -18996 23658 -18910
rect 24162 -18996 24258 -18910
rect 30942 -18996 31038 -18910
rect 31362 -18996 31458 -18910
rect 31962 -18996 32058 -18910
rect 32562 -18996 32658 -18910
rect 33162 -18996 33258 -18910
rect 33762 -18996 33858 -18910
rect 34362 -18996 34458 -18910
rect 34962 -18996 35058 -18910
rect 35562 -18996 35658 -18910
rect 36162 -18996 36258 -18910
rect 36762 -18996 36858 -18910
rect 37362 -18996 37458 -18910
rect 37962 -18996 38058 -18910
rect 38562 -18996 38658 -18910
rect 39162 -18996 39258 -18910
rect 14878 -19470 15478 -19170
rect 24510 -19470 25110 -19170
rect 29878 -19470 30478 -19170
rect 39510 -19470 40110 -19170
rect 10924 -20434 11524 -20134
rect 20556 -20434 21156 -20134
rect 25924 -20434 26524 -20134
rect 35556 -20434 36156 -20134
rect 11776 -20694 11872 -20608
rect 12376 -20694 12472 -20608
rect 12976 -20694 13072 -20608
rect 13576 -20694 13672 -20608
rect 14176 -20694 14272 -20608
rect 14776 -20694 14872 -20608
rect 15376 -20694 15472 -20608
rect 15976 -20694 16072 -20608
rect 16576 -20694 16672 -20608
rect 17176 -20694 17272 -20608
rect 17776 -20694 17872 -20608
rect 18376 -20694 18472 -20608
rect 18976 -20694 19072 -20608
rect 19576 -20694 19672 -20608
rect 19996 -20694 20092 -20608
rect 26776 -20694 26872 -20608
rect 27376 -20694 27472 -20608
rect 27976 -20694 28072 -20608
rect 28576 -20694 28672 -20608
rect 29176 -20694 29272 -20608
rect 29776 -20694 29872 -20608
rect 30376 -20694 30472 -20608
rect 30976 -20694 31072 -20608
rect 31576 -20694 31672 -20608
rect 32176 -20694 32272 -20608
rect 32776 -20694 32872 -20608
rect 33376 -20694 33472 -20608
rect 33976 -20694 34072 -20608
rect 34576 -20694 34672 -20608
rect 34996 -20694 35092 -20608
rect 22175 -25338 22239 -24966
rect 22894 -25338 22958 -24968
rect 23613 -25338 23677 -24968
rect 24332 -25338 24396 -24968
rect 25051 -25338 25115 -24968
rect 22175 -26036 22239 -25668
rect 22894 -26036 22958 -25668
rect 23613 -26036 23677 -25668
rect 24332 -26036 24396 -25668
rect 25051 -26036 25115 -25668
rect 21339 -26157 21437 -26153
rect 21339 -26247 21343 -26157
rect 21343 -26247 21433 -26157
rect 21433 -26247 21437 -26157
rect 21339 -26251 21437 -26247
rect 37175 -25338 37239 -24966
rect 37894 -25338 37958 -24968
rect 38613 -25338 38677 -24968
rect 39332 -25338 39396 -24968
rect 40051 -25338 40115 -24968
rect 37175 -26036 37239 -25668
rect 37894 -26036 37958 -25668
rect 38613 -26036 38677 -25668
rect 39332 -26036 39396 -25668
rect 40051 -26036 40115 -25668
rect 25403 -26157 25501 -26153
rect 25403 -26247 25407 -26157
rect 25407 -26247 25497 -26157
rect 25497 -26247 25501 -26157
rect 25403 -26251 25501 -26247
rect 36339 -26157 36437 -26153
rect 36339 -26247 36343 -26157
rect 36343 -26247 36433 -26157
rect 36433 -26247 36437 -26157
rect 36339 -26251 36437 -26247
rect 22175 -26736 22239 -26368
rect 22894 -26736 22958 -26368
rect 23613 -26736 23677 -26368
rect 24332 -26736 24396 -26368
rect 25051 -26736 25115 -26368
rect 22175 -27436 22239 -27068
rect 22894 -27436 22958 -27068
rect 23613 -27436 23677 -27068
rect 24332 -27436 24396 -27068
rect 25051 -27436 25115 -27068
rect 11210 -27988 11306 -27902
rect 11790 -27988 11886 -27902
rect 12390 -27988 12486 -27902
rect 12990 -27988 13086 -27902
rect 13590 -27988 13686 -27902
rect 14190 -27988 14286 -27902
rect 14790 -27988 14886 -27902
rect 15390 -27988 15486 -27902
rect 15990 -27988 16086 -27902
rect 16590 -27988 16686 -27902
rect 17190 -27988 17286 -27902
rect 17790 -27988 17886 -27902
rect 18390 -27988 18486 -27902
rect 18990 -27988 19086 -27902
rect 19590 -27988 19686 -27902
rect 20190 -27988 20286 -27902
rect 20790 -27988 20886 -27902
rect 22175 -28136 22239 -27768
rect 22894 -28136 22958 -27768
rect 23613 -28136 23677 -27768
rect 24332 -28136 24396 -27768
rect 25051 -28136 25115 -27768
rect 40301 -26157 40399 -26153
rect 40301 -26247 40305 -26157
rect 40305 -26247 40395 -26157
rect 40395 -26247 40399 -26157
rect 40301 -26251 40399 -26247
rect 37175 -26736 37239 -26368
rect 37894 -26736 37958 -26368
rect 38613 -26736 38677 -26368
rect 39332 -26736 39396 -26368
rect 40051 -26736 40115 -26368
rect 37175 -27436 37239 -27068
rect 37894 -27436 37958 -27068
rect 38613 -27436 38677 -27068
rect 39332 -27436 39396 -27068
rect 40051 -27436 40115 -27068
rect 26210 -27988 26306 -27902
rect 26790 -27988 26886 -27902
rect 27390 -27988 27486 -27902
rect 27990 -27988 28086 -27902
rect 28590 -27988 28686 -27902
rect 29190 -27988 29286 -27902
rect 29790 -27988 29886 -27902
rect 30390 -27988 30486 -27902
rect 30990 -27988 31086 -27902
rect 31590 -27988 31686 -27902
rect 32190 -27988 32286 -27902
rect 32790 -27988 32886 -27902
rect 33390 -27988 33486 -27902
rect 33990 -27988 34086 -27902
rect 34590 -27988 34686 -27902
rect 35190 -27988 35286 -27902
rect 35790 -27988 35886 -27902
rect 10924 -28466 11524 -28166
rect 20556 -28466 21156 -28166
rect 37175 -28136 37239 -27768
rect 37894 -28136 37958 -27768
rect 38613 -28136 38677 -27768
rect 39332 -28136 39396 -27768
rect 40051 -28136 40115 -27768
rect 25924 -28466 26524 -28166
rect 35556 -28466 36156 -28166
<< mimcap >>
rect 21660 -6990 22060 -6950
rect 21660 -7310 21700 -6990
rect 22020 -7310 22060 -6990
rect 21660 -7350 22060 -7310
rect 22379 -6990 22779 -6950
rect 22379 -7310 22419 -6990
rect 22739 -7310 22779 -6990
rect 22379 -7350 22779 -7310
rect 23098 -6990 23498 -6950
rect 23098 -7310 23138 -6990
rect 23458 -7310 23498 -6990
rect 23098 -7350 23498 -7310
rect 23817 -6990 24217 -6950
rect 23817 -7310 23857 -6990
rect 24177 -7310 24217 -6990
rect 23817 -7350 24217 -7310
rect 24536 -6990 24936 -6950
rect 24536 -7310 24576 -6990
rect 24896 -7310 24936 -6990
rect 24536 -7350 24936 -7310
rect 36660 -6990 37060 -6950
rect 36660 -7310 36700 -6990
rect 37020 -7310 37060 -6990
rect 36660 -7350 37060 -7310
rect 37379 -6990 37779 -6950
rect 37379 -7310 37419 -6990
rect 37739 -7310 37779 -6990
rect 37379 -7350 37779 -7310
rect 38098 -6990 38498 -6950
rect 38098 -7310 38138 -6990
rect 38458 -7310 38498 -6990
rect 38098 -7350 38498 -7310
rect 38817 -6990 39217 -6950
rect 38817 -7310 38857 -6990
rect 39177 -7310 39217 -6990
rect 38817 -7350 39217 -7310
rect 39536 -6990 39936 -6950
rect 39536 -7310 39576 -6990
rect 39896 -7310 39936 -6990
rect 39536 -7350 39936 -7310
rect 21660 -7690 22060 -7650
rect 21660 -8010 21700 -7690
rect 22020 -8010 22060 -7690
rect 21660 -8050 22060 -8010
rect 22379 -7690 22779 -7650
rect 22379 -8010 22419 -7690
rect 22739 -8010 22779 -7690
rect 22379 -8050 22779 -8010
rect 23098 -7690 23498 -7650
rect 23098 -8010 23138 -7690
rect 23458 -8010 23498 -7690
rect 23098 -8050 23498 -8010
rect 23817 -7690 24217 -7650
rect 23817 -8010 23857 -7690
rect 24177 -8010 24217 -7690
rect 23817 -8050 24217 -8010
rect 24536 -7690 24936 -7650
rect 24536 -8010 24576 -7690
rect 24896 -8010 24936 -7690
rect 24536 -8050 24936 -8010
rect 36660 -7690 37060 -7650
rect 36660 -8010 36700 -7690
rect 37020 -8010 37060 -7690
rect 36660 -8050 37060 -8010
rect 37379 -7690 37779 -7650
rect 37379 -8010 37419 -7690
rect 37739 -8010 37779 -7690
rect 37379 -8050 37779 -8010
rect 38098 -7690 38498 -7650
rect 38098 -8010 38138 -7690
rect 38458 -8010 38498 -7690
rect 38098 -8050 38498 -8010
rect 38817 -7690 39217 -7650
rect 38817 -8010 38857 -7690
rect 39177 -8010 39217 -7690
rect 38817 -8050 39217 -8010
rect 39536 -7690 39936 -7650
rect 39536 -8010 39576 -7690
rect 39896 -8010 39936 -7690
rect 39536 -8050 39936 -8010
rect 21660 -8390 22060 -8350
rect 21660 -8710 21700 -8390
rect 22020 -8710 22060 -8390
rect 21660 -8750 22060 -8710
rect 22379 -8390 22779 -8350
rect 22379 -8710 22419 -8390
rect 22739 -8710 22779 -8390
rect 22379 -8750 22779 -8710
rect 23098 -8390 23498 -8350
rect 23098 -8710 23138 -8390
rect 23458 -8710 23498 -8390
rect 23098 -8750 23498 -8710
rect 23817 -8390 24217 -8350
rect 23817 -8710 23857 -8390
rect 24177 -8710 24217 -8390
rect 23817 -8750 24217 -8710
rect 24536 -8390 24936 -8350
rect 24536 -8710 24576 -8390
rect 24896 -8710 24936 -8390
rect 24536 -8750 24936 -8710
rect 36660 -8390 37060 -8350
rect 36660 -8710 36700 -8390
rect 37020 -8710 37060 -8390
rect 36660 -8750 37060 -8710
rect 37379 -8390 37779 -8350
rect 37379 -8710 37419 -8390
rect 37739 -8710 37779 -8390
rect 37379 -8750 37779 -8710
rect 38098 -8390 38498 -8350
rect 38098 -8710 38138 -8390
rect 38458 -8710 38498 -8390
rect 38098 -8750 38498 -8710
rect 38817 -8390 39217 -8350
rect 38817 -8710 38857 -8390
rect 39177 -8710 39217 -8390
rect 38817 -8750 39217 -8710
rect 39536 -8390 39936 -8350
rect 39536 -8710 39576 -8390
rect 39896 -8710 39936 -8390
rect 39536 -8750 39936 -8710
rect 21660 -9090 22060 -9050
rect 21660 -9410 21700 -9090
rect 22020 -9410 22060 -9090
rect 21660 -9450 22060 -9410
rect 22379 -9090 22779 -9050
rect 22379 -9410 22419 -9090
rect 22739 -9410 22779 -9090
rect 22379 -9450 22779 -9410
rect 23098 -9090 23498 -9050
rect 23098 -9410 23138 -9090
rect 23458 -9410 23498 -9090
rect 23098 -9450 23498 -9410
rect 23817 -9090 24217 -9050
rect 23817 -9410 23857 -9090
rect 24177 -9410 24217 -9090
rect 23817 -9450 24217 -9410
rect 24536 -9090 24936 -9050
rect 24536 -9410 24576 -9090
rect 24896 -9410 24936 -9090
rect 24536 -9450 24936 -9410
rect 36660 -9090 37060 -9050
rect 36660 -9410 36700 -9090
rect 37020 -9410 37060 -9090
rect 36660 -9450 37060 -9410
rect 37379 -9090 37779 -9050
rect 37379 -9410 37419 -9090
rect 37739 -9410 37779 -9090
rect 37379 -9450 37779 -9410
rect 38098 -9090 38498 -9050
rect 38098 -9410 38138 -9090
rect 38458 -9410 38498 -9090
rect 38098 -9450 38498 -9410
rect 38817 -9090 39217 -9050
rect 38817 -9410 38857 -9090
rect 39177 -9410 39217 -9090
rect 38817 -9450 39217 -9410
rect 39536 -9090 39936 -9050
rect 39536 -9410 39576 -9090
rect 39896 -9410 39936 -9090
rect 39536 -9450 39936 -9410
rect 21660 -9790 22060 -9750
rect 21660 -10110 21700 -9790
rect 22020 -10110 22060 -9790
rect 21660 -10150 22060 -10110
rect 22379 -9790 22779 -9750
rect 22379 -10110 22419 -9790
rect 22739 -10110 22779 -9790
rect 22379 -10150 22779 -10110
rect 23098 -9790 23498 -9750
rect 23098 -10110 23138 -9790
rect 23458 -10110 23498 -9790
rect 23098 -10150 23498 -10110
rect 23817 -9790 24217 -9750
rect 23817 -10110 23857 -9790
rect 24177 -10110 24217 -9790
rect 23817 -10150 24217 -10110
rect 24536 -9790 24936 -9750
rect 24536 -10110 24576 -9790
rect 24896 -10110 24936 -9790
rect 24536 -10150 24936 -10110
rect 36660 -9790 37060 -9750
rect 36660 -10110 36700 -9790
rect 37020 -10110 37060 -9790
rect 36660 -10150 37060 -10110
rect 37379 -9790 37779 -9750
rect 37379 -10110 37419 -9790
rect 37739 -10110 37779 -9790
rect 37379 -10150 37779 -10110
rect 38098 -9790 38498 -9750
rect 38098 -10110 38138 -9790
rect 38458 -10110 38498 -9790
rect 38098 -10150 38498 -10110
rect 38817 -9790 39217 -9750
rect 38817 -10110 38857 -9790
rect 39177 -10110 39217 -9790
rect 38817 -10150 39217 -10110
rect 39536 -9790 39936 -9750
rect 39536 -10110 39576 -9790
rect 39896 -10110 39936 -9790
rect 39536 -10150 39936 -10110
rect 11098 -11494 11498 -11454
rect 11098 -11814 11138 -11494
rect 11458 -11814 11498 -11494
rect 11098 -11854 11498 -11814
rect 11817 -11494 12217 -11454
rect 11817 -11814 11857 -11494
rect 12177 -11814 12217 -11494
rect 11817 -11854 12217 -11814
rect 12536 -11494 12936 -11454
rect 12536 -11814 12576 -11494
rect 12896 -11814 12936 -11494
rect 12536 -11854 12936 -11814
rect 13255 -11494 13655 -11454
rect 13255 -11814 13295 -11494
rect 13615 -11814 13655 -11494
rect 13255 -11854 13655 -11814
rect 13974 -11494 14374 -11454
rect 13974 -11814 14014 -11494
rect 14334 -11814 14374 -11494
rect 13974 -11854 14374 -11814
rect 26098 -11494 26498 -11454
rect 26098 -11814 26138 -11494
rect 26458 -11814 26498 -11494
rect 26098 -11854 26498 -11814
rect 26817 -11494 27217 -11454
rect 26817 -11814 26857 -11494
rect 27177 -11814 27217 -11494
rect 26817 -11854 27217 -11814
rect 27536 -11494 27936 -11454
rect 27536 -11814 27576 -11494
rect 27896 -11814 27936 -11494
rect 27536 -11854 27936 -11814
rect 28255 -11494 28655 -11454
rect 28255 -11814 28295 -11494
rect 28615 -11814 28655 -11494
rect 28255 -11854 28655 -11814
rect 28974 -11494 29374 -11454
rect 28974 -11814 29014 -11494
rect 29334 -11814 29374 -11494
rect 28974 -11854 29374 -11814
rect 11098 -12194 11498 -12154
rect 11098 -12514 11138 -12194
rect 11458 -12514 11498 -12194
rect 11098 -12554 11498 -12514
rect 11817 -12194 12217 -12154
rect 11817 -12514 11857 -12194
rect 12177 -12514 12217 -12194
rect 11817 -12554 12217 -12514
rect 12536 -12194 12936 -12154
rect 12536 -12514 12576 -12194
rect 12896 -12514 12936 -12194
rect 12536 -12554 12936 -12514
rect 13255 -12194 13655 -12154
rect 13255 -12514 13295 -12194
rect 13615 -12514 13655 -12194
rect 13255 -12554 13655 -12514
rect 13974 -12194 14374 -12154
rect 13974 -12514 14014 -12194
rect 14334 -12514 14374 -12194
rect 13974 -12554 14374 -12514
rect 26098 -12194 26498 -12154
rect 26098 -12514 26138 -12194
rect 26458 -12514 26498 -12194
rect 26098 -12554 26498 -12514
rect 26817 -12194 27217 -12154
rect 26817 -12514 26857 -12194
rect 27177 -12514 27217 -12194
rect 26817 -12554 27217 -12514
rect 27536 -12194 27936 -12154
rect 27536 -12514 27576 -12194
rect 27896 -12514 27936 -12194
rect 27536 -12554 27936 -12514
rect 28255 -12194 28655 -12154
rect 28255 -12514 28295 -12194
rect 28615 -12514 28655 -12194
rect 28255 -12554 28655 -12514
rect 28974 -12194 29374 -12154
rect 28974 -12514 29014 -12194
rect 29334 -12514 29374 -12194
rect 28974 -12554 29374 -12514
rect 11098 -12894 11498 -12854
rect 11098 -13214 11138 -12894
rect 11458 -13214 11498 -12894
rect 11098 -13254 11498 -13214
rect 11817 -12894 12217 -12854
rect 11817 -13214 11857 -12894
rect 12177 -13214 12217 -12894
rect 11817 -13254 12217 -13214
rect 12536 -12894 12936 -12854
rect 12536 -13214 12576 -12894
rect 12896 -13214 12936 -12894
rect 12536 -13254 12936 -13214
rect 13255 -12894 13655 -12854
rect 13255 -13214 13295 -12894
rect 13615 -13214 13655 -12894
rect 13255 -13254 13655 -13214
rect 13974 -12894 14374 -12854
rect 13974 -13214 14014 -12894
rect 14334 -13214 14374 -12894
rect 13974 -13254 14374 -13214
rect 26098 -12894 26498 -12854
rect 26098 -13214 26138 -12894
rect 26458 -13214 26498 -12894
rect 26098 -13254 26498 -13214
rect 26817 -12894 27217 -12854
rect 26817 -13214 26857 -12894
rect 27177 -13214 27217 -12894
rect 26817 -13254 27217 -13214
rect 27536 -12894 27936 -12854
rect 27536 -13214 27576 -12894
rect 27896 -13214 27936 -12894
rect 27536 -13254 27936 -13214
rect 28255 -12894 28655 -12854
rect 28255 -13214 28295 -12894
rect 28615 -13214 28655 -12894
rect 28255 -13254 28655 -13214
rect 28974 -12894 29374 -12854
rect 28974 -13214 29014 -12894
rect 29334 -13214 29374 -12894
rect 28974 -13254 29374 -13214
rect 11098 -13594 11498 -13554
rect 11098 -13914 11138 -13594
rect 11458 -13914 11498 -13594
rect 11098 -13954 11498 -13914
rect 11817 -13594 12217 -13554
rect 11817 -13914 11857 -13594
rect 12177 -13914 12217 -13594
rect 11817 -13954 12217 -13914
rect 12536 -13594 12936 -13554
rect 12536 -13914 12576 -13594
rect 12896 -13914 12936 -13594
rect 12536 -13954 12936 -13914
rect 13255 -13594 13655 -13554
rect 13255 -13914 13295 -13594
rect 13615 -13914 13655 -13594
rect 13255 -13954 13655 -13914
rect 13974 -13594 14374 -13554
rect 13974 -13914 14014 -13594
rect 14334 -13914 14374 -13594
rect 13974 -13954 14374 -13914
rect 26098 -13594 26498 -13554
rect 26098 -13914 26138 -13594
rect 26458 -13914 26498 -13594
rect 26098 -13954 26498 -13914
rect 26817 -13594 27217 -13554
rect 26817 -13914 26857 -13594
rect 27177 -13914 27217 -13594
rect 26817 -13954 27217 -13914
rect 27536 -13594 27936 -13554
rect 27536 -13914 27576 -13594
rect 27896 -13914 27936 -13594
rect 27536 -13954 27936 -13914
rect 28255 -13594 28655 -13554
rect 28255 -13914 28295 -13594
rect 28615 -13914 28655 -13594
rect 28255 -13954 28655 -13914
rect 28974 -13594 29374 -13554
rect 28974 -13914 29014 -13594
rect 29334 -13914 29374 -13594
rect 28974 -13954 29374 -13914
rect 11098 -14294 11498 -14254
rect 11098 -14614 11138 -14294
rect 11458 -14614 11498 -14294
rect 11098 -14654 11498 -14614
rect 11817 -14294 12217 -14254
rect 11817 -14614 11857 -14294
rect 12177 -14614 12217 -14294
rect 11817 -14654 12217 -14614
rect 12536 -14294 12936 -14254
rect 12536 -14614 12576 -14294
rect 12896 -14614 12936 -14294
rect 12536 -14654 12936 -14614
rect 13255 -14294 13655 -14254
rect 13255 -14614 13295 -14294
rect 13615 -14614 13655 -14294
rect 13255 -14654 13655 -14614
rect 13974 -14294 14374 -14254
rect 13974 -14614 14014 -14294
rect 14334 -14614 14374 -14294
rect 13974 -14654 14374 -14614
rect 26098 -14294 26498 -14254
rect 26098 -14614 26138 -14294
rect 26458 -14614 26498 -14294
rect 26098 -14654 26498 -14614
rect 26817 -14294 27217 -14254
rect 26817 -14614 26857 -14294
rect 27177 -14614 27217 -14294
rect 26817 -14654 27217 -14614
rect 27536 -14294 27936 -14254
rect 27536 -14614 27576 -14294
rect 27896 -14614 27936 -14294
rect 27536 -14654 27936 -14614
rect 28255 -14294 28655 -14254
rect 28255 -14614 28295 -14294
rect 28615 -14614 28655 -14294
rect 28255 -14654 28655 -14614
rect 28974 -14294 29374 -14254
rect 28974 -14614 29014 -14294
rect 29334 -14614 29374 -14294
rect 28974 -14654 29374 -14614
rect 21660 -24990 22060 -24950
rect 21660 -25310 21700 -24990
rect 22020 -25310 22060 -24990
rect 21660 -25350 22060 -25310
rect 22379 -24990 22779 -24950
rect 22379 -25310 22419 -24990
rect 22739 -25310 22779 -24990
rect 22379 -25350 22779 -25310
rect 23098 -24990 23498 -24950
rect 23098 -25310 23138 -24990
rect 23458 -25310 23498 -24990
rect 23098 -25350 23498 -25310
rect 23817 -24990 24217 -24950
rect 23817 -25310 23857 -24990
rect 24177 -25310 24217 -24990
rect 23817 -25350 24217 -25310
rect 24536 -24990 24936 -24950
rect 24536 -25310 24576 -24990
rect 24896 -25310 24936 -24990
rect 24536 -25350 24936 -25310
rect 36660 -24990 37060 -24950
rect 36660 -25310 36700 -24990
rect 37020 -25310 37060 -24990
rect 36660 -25350 37060 -25310
rect 37379 -24990 37779 -24950
rect 37379 -25310 37419 -24990
rect 37739 -25310 37779 -24990
rect 37379 -25350 37779 -25310
rect 38098 -24990 38498 -24950
rect 38098 -25310 38138 -24990
rect 38458 -25310 38498 -24990
rect 38098 -25350 38498 -25310
rect 38817 -24990 39217 -24950
rect 38817 -25310 38857 -24990
rect 39177 -25310 39217 -24990
rect 38817 -25350 39217 -25310
rect 39536 -24990 39936 -24950
rect 39536 -25310 39576 -24990
rect 39896 -25310 39936 -24990
rect 39536 -25350 39936 -25310
rect 21660 -25690 22060 -25650
rect 21660 -26010 21700 -25690
rect 22020 -26010 22060 -25690
rect 21660 -26050 22060 -26010
rect 22379 -25690 22779 -25650
rect 22379 -26010 22419 -25690
rect 22739 -26010 22779 -25690
rect 22379 -26050 22779 -26010
rect 23098 -25690 23498 -25650
rect 23098 -26010 23138 -25690
rect 23458 -26010 23498 -25690
rect 23098 -26050 23498 -26010
rect 23817 -25690 24217 -25650
rect 23817 -26010 23857 -25690
rect 24177 -26010 24217 -25690
rect 23817 -26050 24217 -26010
rect 24536 -25690 24936 -25650
rect 24536 -26010 24576 -25690
rect 24896 -26010 24936 -25690
rect 24536 -26050 24936 -26010
rect 36660 -25690 37060 -25650
rect 36660 -26010 36700 -25690
rect 37020 -26010 37060 -25690
rect 36660 -26050 37060 -26010
rect 37379 -25690 37779 -25650
rect 37379 -26010 37419 -25690
rect 37739 -26010 37779 -25690
rect 37379 -26050 37779 -26010
rect 38098 -25690 38498 -25650
rect 38098 -26010 38138 -25690
rect 38458 -26010 38498 -25690
rect 38098 -26050 38498 -26010
rect 38817 -25690 39217 -25650
rect 38817 -26010 38857 -25690
rect 39177 -26010 39217 -25690
rect 38817 -26050 39217 -26010
rect 39536 -25690 39936 -25650
rect 39536 -26010 39576 -25690
rect 39896 -26010 39936 -25690
rect 39536 -26050 39936 -26010
rect 21660 -26390 22060 -26350
rect 21660 -26710 21700 -26390
rect 22020 -26710 22060 -26390
rect 21660 -26750 22060 -26710
rect 22379 -26390 22779 -26350
rect 22379 -26710 22419 -26390
rect 22739 -26710 22779 -26390
rect 22379 -26750 22779 -26710
rect 23098 -26390 23498 -26350
rect 23098 -26710 23138 -26390
rect 23458 -26710 23498 -26390
rect 23098 -26750 23498 -26710
rect 23817 -26390 24217 -26350
rect 23817 -26710 23857 -26390
rect 24177 -26710 24217 -26390
rect 23817 -26750 24217 -26710
rect 24536 -26390 24936 -26350
rect 24536 -26710 24576 -26390
rect 24896 -26710 24936 -26390
rect 24536 -26750 24936 -26710
rect 36660 -26390 37060 -26350
rect 36660 -26710 36700 -26390
rect 37020 -26710 37060 -26390
rect 36660 -26750 37060 -26710
rect 37379 -26390 37779 -26350
rect 37379 -26710 37419 -26390
rect 37739 -26710 37779 -26390
rect 37379 -26750 37779 -26710
rect 38098 -26390 38498 -26350
rect 38098 -26710 38138 -26390
rect 38458 -26710 38498 -26390
rect 38098 -26750 38498 -26710
rect 38817 -26390 39217 -26350
rect 38817 -26710 38857 -26390
rect 39177 -26710 39217 -26390
rect 38817 -26750 39217 -26710
rect 39536 -26390 39936 -26350
rect 39536 -26710 39576 -26390
rect 39896 -26710 39936 -26390
rect 39536 -26750 39936 -26710
rect 21660 -27090 22060 -27050
rect 21660 -27410 21700 -27090
rect 22020 -27410 22060 -27090
rect 21660 -27450 22060 -27410
rect 22379 -27090 22779 -27050
rect 22379 -27410 22419 -27090
rect 22739 -27410 22779 -27090
rect 22379 -27450 22779 -27410
rect 23098 -27090 23498 -27050
rect 23098 -27410 23138 -27090
rect 23458 -27410 23498 -27090
rect 23098 -27450 23498 -27410
rect 23817 -27090 24217 -27050
rect 23817 -27410 23857 -27090
rect 24177 -27410 24217 -27090
rect 23817 -27450 24217 -27410
rect 24536 -27090 24936 -27050
rect 24536 -27410 24576 -27090
rect 24896 -27410 24936 -27090
rect 24536 -27450 24936 -27410
rect 36660 -27090 37060 -27050
rect 36660 -27410 36700 -27090
rect 37020 -27410 37060 -27090
rect 36660 -27450 37060 -27410
rect 37379 -27090 37779 -27050
rect 37379 -27410 37419 -27090
rect 37739 -27410 37779 -27090
rect 37379 -27450 37779 -27410
rect 38098 -27090 38498 -27050
rect 38098 -27410 38138 -27090
rect 38458 -27410 38498 -27090
rect 38098 -27450 38498 -27410
rect 38817 -27090 39217 -27050
rect 38817 -27410 38857 -27090
rect 39177 -27410 39217 -27090
rect 38817 -27450 39217 -27410
rect 39536 -27090 39936 -27050
rect 39536 -27410 39576 -27090
rect 39896 -27410 39936 -27090
rect 39536 -27450 39936 -27410
rect 21660 -27790 22060 -27750
rect 21660 -28110 21700 -27790
rect 22020 -28110 22060 -27790
rect 21660 -28150 22060 -28110
rect 22379 -27790 22779 -27750
rect 22379 -28110 22419 -27790
rect 22739 -28110 22779 -27790
rect 22379 -28150 22779 -28110
rect 23098 -27790 23498 -27750
rect 23098 -28110 23138 -27790
rect 23458 -28110 23498 -27790
rect 23098 -28150 23498 -28110
rect 23817 -27790 24217 -27750
rect 23817 -28110 23857 -27790
rect 24177 -28110 24217 -27790
rect 23817 -28150 24217 -28110
rect 24536 -27790 24936 -27750
rect 24536 -28110 24576 -27790
rect 24896 -28110 24936 -27790
rect 24536 -28150 24936 -28110
rect 36660 -27790 37060 -27750
rect 36660 -28110 36700 -27790
rect 37020 -28110 37060 -27790
rect 36660 -28150 37060 -28110
rect 37379 -27790 37779 -27750
rect 37379 -28110 37419 -27790
rect 37739 -28110 37779 -27790
rect 37379 -28150 37779 -28110
rect 38098 -27790 38498 -27750
rect 38098 -28110 38138 -27790
rect 38458 -28110 38498 -27790
rect 38098 -28150 38498 -28110
rect 38817 -27790 39217 -27750
rect 38817 -28110 38857 -27790
rect 39177 -28110 39217 -27790
rect 38817 -28150 39217 -28110
rect 39536 -27790 39936 -27750
rect 39536 -28110 39576 -27790
rect 39896 -28110 39936 -27790
rect 39536 -28150 39936 -28110
<< mimcapcontact >>
rect 21700 -7310 22020 -6990
rect 22419 -7310 22739 -6990
rect 23138 -7310 23458 -6990
rect 23857 -7310 24177 -6990
rect 24576 -7310 24896 -6990
rect 36700 -7310 37020 -6990
rect 37419 -7310 37739 -6990
rect 38138 -7310 38458 -6990
rect 38857 -7310 39177 -6990
rect 39576 -7310 39896 -6990
rect 21700 -8010 22020 -7690
rect 22419 -8010 22739 -7690
rect 23138 -8010 23458 -7690
rect 23857 -8010 24177 -7690
rect 24576 -8010 24896 -7690
rect 36700 -8010 37020 -7690
rect 37419 -8010 37739 -7690
rect 38138 -8010 38458 -7690
rect 38857 -8010 39177 -7690
rect 39576 -8010 39896 -7690
rect 21700 -8710 22020 -8390
rect 22419 -8710 22739 -8390
rect 23138 -8710 23458 -8390
rect 23857 -8710 24177 -8390
rect 24576 -8710 24896 -8390
rect 36700 -8710 37020 -8390
rect 37419 -8710 37739 -8390
rect 38138 -8710 38458 -8390
rect 38857 -8710 39177 -8390
rect 39576 -8710 39896 -8390
rect 21700 -9410 22020 -9090
rect 22419 -9410 22739 -9090
rect 23138 -9410 23458 -9090
rect 23857 -9410 24177 -9090
rect 24576 -9410 24896 -9090
rect 36700 -9410 37020 -9090
rect 37419 -9410 37739 -9090
rect 38138 -9410 38458 -9090
rect 38857 -9410 39177 -9090
rect 39576 -9410 39896 -9090
rect 21700 -10110 22020 -9790
rect 22419 -10110 22739 -9790
rect 23138 -10110 23458 -9790
rect 23857 -10110 24177 -9790
rect 24576 -10110 24896 -9790
rect 36700 -10110 37020 -9790
rect 37419 -10110 37739 -9790
rect 38138 -10110 38458 -9790
rect 38857 -10110 39177 -9790
rect 39576 -10110 39896 -9790
rect 11138 -11814 11458 -11494
rect 11857 -11814 12177 -11494
rect 12576 -11814 12896 -11494
rect 13295 -11814 13615 -11494
rect 14014 -11814 14334 -11494
rect 26138 -11814 26458 -11494
rect 26857 -11814 27177 -11494
rect 27576 -11814 27896 -11494
rect 28295 -11814 28615 -11494
rect 29014 -11814 29334 -11494
rect 11138 -12514 11458 -12194
rect 11857 -12514 12177 -12194
rect 12576 -12514 12896 -12194
rect 13295 -12514 13615 -12194
rect 14014 -12514 14334 -12194
rect 26138 -12514 26458 -12194
rect 26857 -12514 27177 -12194
rect 27576 -12514 27896 -12194
rect 28295 -12514 28615 -12194
rect 29014 -12514 29334 -12194
rect 11138 -13214 11458 -12894
rect 11857 -13214 12177 -12894
rect 12576 -13214 12896 -12894
rect 13295 -13214 13615 -12894
rect 14014 -13214 14334 -12894
rect 26138 -13214 26458 -12894
rect 26857 -13214 27177 -12894
rect 27576 -13214 27896 -12894
rect 28295 -13214 28615 -12894
rect 29014 -13214 29334 -12894
rect 11138 -13914 11458 -13594
rect 11857 -13914 12177 -13594
rect 12576 -13914 12896 -13594
rect 13295 -13914 13615 -13594
rect 14014 -13914 14334 -13594
rect 26138 -13914 26458 -13594
rect 26857 -13914 27177 -13594
rect 27576 -13914 27896 -13594
rect 28295 -13914 28615 -13594
rect 29014 -13914 29334 -13594
rect 11138 -14614 11458 -14294
rect 11857 -14614 12177 -14294
rect 12576 -14614 12896 -14294
rect 13295 -14614 13615 -14294
rect 14014 -14614 14334 -14294
rect 26138 -14614 26458 -14294
rect 26857 -14614 27177 -14294
rect 27576 -14614 27896 -14294
rect 28295 -14614 28615 -14294
rect 29014 -14614 29334 -14294
rect 21700 -25310 22020 -24990
rect 22419 -25310 22739 -24990
rect 23138 -25310 23458 -24990
rect 23857 -25310 24177 -24990
rect 24576 -25310 24896 -24990
rect 36700 -25310 37020 -24990
rect 37419 -25310 37739 -24990
rect 38138 -25310 38458 -24990
rect 38857 -25310 39177 -24990
rect 39576 -25310 39896 -24990
rect 21700 -26010 22020 -25690
rect 22419 -26010 22739 -25690
rect 23138 -26010 23458 -25690
rect 23857 -26010 24177 -25690
rect 24576 -26010 24896 -25690
rect 36700 -26010 37020 -25690
rect 37419 -26010 37739 -25690
rect 38138 -26010 38458 -25690
rect 38857 -26010 39177 -25690
rect 39576 -26010 39896 -25690
rect 21700 -26710 22020 -26390
rect 22419 -26710 22739 -26390
rect 23138 -26710 23458 -26390
rect 23857 -26710 24177 -26390
rect 24576 -26710 24896 -26390
rect 36700 -26710 37020 -26390
rect 37419 -26710 37739 -26390
rect 38138 -26710 38458 -26390
rect 38857 -26710 39177 -26390
rect 39576 -26710 39896 -26390
rect 21700 -27410 22020 -27090
rect 22419 -27410 22739 -27090
rect 23138 -27410 23458 -27090
rect 23857 -27410 24177 -27090
rect 24576 -27410 24896 -27090
rect 36700 -27410 37020 -27090
rect 37419 -27410 37739 -27090
rect 38138 -27410 38458 -27090
rect 38857 -27410 39177 -27090
rect 39576 -27410 39896 -27090
rect 21700 -28110 22020 -27790
rect 22419 -28110 22739 -27790
rect 23138 -28110 23458 -27790
rect 23857 -28110 24177 -27790
rect 24576 -28110 24896 -27790
rect 36700 -28110 37020 -27790
rect 37419 -28110 37739 -27790
rect 38138 -28110 38458 -27790
rect 38857 -28110 39177 -27790
rect 39576 -28110 39896 -27790
<< metal4 >>
rect 10584 4204 40288 4388
rect 10584 3904 15532 4204
rect 15914 3904 23666 4204
rect 24344 3904 26114 4204
rect 26714 3904 30746 4204
rect 31346 3904 40288 4204
rect 10584 3726 40288 3904
rect 10584 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 40288 3726
rect 10584 3588 40288 3640
rect 15348 -940 31530 -936
rect 10744 -974 41209 -940
rect 10744 -1252 40432 -974
rect 10744 -1552 15532 -1252
rect 15914 -1552 23666 -1252
rect 24344 -1552 26114 -1252
rect 26714 -1552 30746 -1252
rect 31346 -1552 40432 -1252
rect 10744 -1950 40432 -1552
rect 10740 -2134 40432 -1950
rect 10740 -2434 10924 -2134
rect 11524 -2434 20556 -2134
rect 21156 -2434 25924 -2134
rect 26524 -2434 35556 -2134
rect 36156 -2434 40432 -2134
rect 10740 -2608 40432 -2434
rect 10740 -2694 11776 -2608
rect 11872 -2694 12376 -2608
rect 12472 -2694 12976 -2608
rect 13072 -2694 13576 -2608
rect 13672 -2694 14176 -2608
rect 14272 -2694 14776 -2608
rect 14872 -2694 15376 -2608
rect 15472 -2694 15976 -2608
rect 16072 -2694 16576 -2608
rect 16672 -2694 17176 -2608
rect 17272 -2694 17776 -2608
rect 17872 -2694 18376 -2608
rect 18472 -2694 18976 -2608
rect 19072 -2694 19576 -2608
rect 19672 -2694 19996 -2608
rect 20092 -2694 26776 -2608
rect 26872 -2694 27376 -2608
rect 27472 -2694 27976 -2608
rect 28072 -2694 28576 -2608
rect 28672 -2694 29176 -2608
rect 29272 -2694 29776 -2608
rect 29872 -2694 30376 -2608
rect 30472 -2694 30976 -2608
rect 31072 -2694 31576 -2608
rect 31672 -2694 32176 -2608
rect 32272 -2694 32776 -2608
rect 32872 -2694 33376 -2608
rect 33472 -2694 33976 -2608
rect 34072 -2694 34576 -2608
rect 34672 -2694 34996 -2608
rect 35092 -2694 40432 -2608
rect 10740 -2722 40432 -2694
rect 41178 -2722 41209 -974
rect 10740 -2750 41209 -2722
rect 22159 -6966 22255 -6950
rect 21699 -6990 22021 -6989
rect 21699 -7310 21700 -6990
rect 22020 -7106 22021 -6990
rect 22159 -7106 22175 -6966
rect 22020 -7206 22175 -7106
rect 22020 -7310 22021 -7206
rect 21699 -7311 22021 -7310
rect 21814 -7689 21914 -7311
rect 22150 -7338 22175 -7206
rect 22239 -7106 22255 -6966
rect 22878 -6968 22974 -6952
rect 22418 -6990 22740 -6989
rect 22418 -7106 22419 -6990
rect 22239 -7206 22419 -7106
rect 22239 -7338 22255 -7206
rect 22418 -7310 22419 -7206
rect 22739 -7106 22740 -6990
rect 22878 -7106 22894 -6968
rect 22739 -7206 22894 -7106
rect 22739 -7310 22740 -7206
rect 22418 -7311 22740 -7310
rect 22150 -7354 22255 -7338
rect 22878 -7338 22894 -7206
rect 22958 -7106 22974 -6968
rect 23597 -6968 23693 -6952
rect 23137 -6990 23459 -6989
rect 23137 -7106 23138 -6990
rect 22958 -7206 23138 -7106
rect 22958 -7338 22974 -7206
rect 23137 -7310 23138 -7206
rect 23458 -7106 23459 -6990
rect 23597 -7106 23613 -6968
rect 23458 -7206 23613 -7106
rect 23458 -7310 23459 -7206
rect 23137 -7311 23459 -7310
rect 22878 -7354 22974 -7338
rect 23597 -7338 23613 -7206
rect 23677 -7106 23693 -6968
rect 24316 -6968 24412 -6952
rect 23856 -6990 24178 -6989
rect 23856 -7106 23857 -6990
rect 23677 -7206 23857 -7106
rect 23677 -7338 23693 -7206
rect 23856 -7310 23857 -7206
rect 24177 -7106 24178 -6990
rect 24316 -7106 24332 -6968
rect 24177 -7206 24332 -7106
rect 24177 -7310 24178 -7206
rect 23856 -7311 24178 -7310
rect 23597 -7354 23693 -7338
rect 24316 -7338 24332 -7206
rect 24396 -7106 24412 -6968
rect 25035 -6968 25131 -6952
rect 24575 -6990 24897 -6989
rect 24575 -7106 24576 -6990
rect 24396 -7206 24576 -7106
rect 24396 -7338 24418 -7206
rect 24575 -7310 24576 -7206
rect 24896 -7106 24897 -6990
rect 25035 -7106 25051 -6968
rect 24896 -7206 25051 -7106
rect 24896 -7310 24897 -7206
rect 24575 -7311 24897 -7310
rect 22150 -7652 22250 -7354
rect 22528 -7560 24072 -7460
rect 22150 -7668 22255 -7652
rect 21699 -7690 22021 -7689
rect 21699 -8010 21700 -7690
rect 22020 -7796 22021 -7690
rect 22150 -7796 22175 -7668
rect 22020 -7896 22175 -7796
rect 22020 -8010 22021 -7896
rect 22150 -8010 22175 -7896
rect 21699 -8011 22021 -8010
rect 22159 -8036 22175 -8010
rect 22239 -8036 22255 -7668
rect 22528 -7689 22628 -7560
rect 22878 -7668 22974 -7652
rect 22418 -7690 22740 -7689
rect 22418 -8010 22419 -7690
rect 22739 -8010 22740 -7690
rect 22418 -8011 22740 -8010
rect 22159 -8056 22255 -8036
rect 22528 -8152 22628 -8011
rect 22878 -8036 22894 -7668
rect 22958 -8036 22974 -7668
rect 23248 -7689 23348 -7560
rect 23597 -7668 23693 -7652
rect 23137 -7690 23459 -7689
rect 23137 -8010 23138 -7690
rect 23458 -8010 23459 -7690
rect 23137 -8011 23459 -8010
rect 22878 -8056 22974 -8036
rect 23248 -8152 23348 -8011
rect 23597 -8036 23613 -7668
rect 23677 -8036 23693 -7668
rect 23970 -7689 24071 -7560
rect 24316 -7668 24418 -7338
rect 23856 -7690 24178 -7689
rect 23856 -8010 23857 -7690
rect 24177 -8010 24178 -7690
rect 23856 -8011 24178 -8010
rect 23597 -8056 23693 -8036
rect 23970 -8152 24071 -8011
rect 24316 -8036 24332 -7668
rect 24396 -7800 24418 -7668
rect 24690 -7689 24790 -7311
rect 25028 -7338 25051 -7206
rect 25115 -7338 25131 -6968
rect 37159 -6966 37255 -6950
rect 36699 -6990 37021 -6989
rect 36699 -7310 36700 -6990
rect 37020 -7106 37021 -6990
rect 37159 -7106 37175 -6966
rect 37020 -7206 37175 -7106
rect 37020 -7310 37021 -7206
rect 36699 -7311 37021 -7310
rect 25028 -7668 25131 -7338
rect 24575 -7690 24897 -7689
rect 24575 -7800 24576 -7690
rect 24396 -7900 24576 -7800
rect 24396 -8036 24418 -7900
rect 24575 -8010 24576 -7900
rect 24896 -7800 24897 -7690
rect 25028 -7800 25051 -7668
rect 24896 -7900 25051 -7800
rect 24896 -8010 24897 -7900
rect 24575 -8011 24897 -8010
rect 24690 -8012 24790 -8011
rect 24316 -8050 24418 -8036
rect 25028 -8036 25051 -7900
rect 25115 -8036 25131 -7668
rect 36814 -7689 36914 -7311
rect 37150 -7338 37175 -7206
rect 37239 -7106 37255 -6966
rect 37878 -6968 37974 -6952
rect 37418 -6990 37740 -6989
rect 37418 -7106 37419 -6990
rect 37239 -7206 37419 -7106
rect 37239 -7338 37255 -7206
rect 37418 -7310 37419 -7206
rect 37739 -7106 37740 -6990
rect 37878 -7106 37894 -6968
rect 37739 -7206 37894 -7106
rect 37739 -7310 37740 -7206
rect 37418 -7311 37740 -7310
rect 37150 -7354 37255 -7338
rect 37878 -7338 37894 -7206
rect 37958 -7106 37974 -6968
rect 38597 -6968 38693 -6952
rect 38137 -6990 38459 -6989
rect 38137 -7106 38138 -6990
rect 37958 -7206 38138 -7106
rect 37958 -7338 37974 -7206
rect 38137 -7310 38138 -7206
rect 38458 -7106 38459 -6990
rect 38597 -7106 38613 -6968
rect 38458 -7206 38613 -7106
rect 38458 -7310 38459 -7206
rect 38137 -7311 38459 -7310
rect 37878 -7354 37974 -7338
rect 38597 -7338 38613 -7206
rect 38677 -7106 38693 -6968
rect 39316 -6968 39412 -6952
rect 38856 -6990 39178 -6989
rect 38856 -7106 38857 -6990
rect 38677 -7206 38857 -7106
rect 38677 -7338 38693 -7206
rect 38856 -7310 38857 -7206
rect 39177 -7106 39178 -6990
rect 39316 -7106 39332 -6968
rect 39177 -7206 39332 -7106
rect 39177 -7310 39178 -7206
rect 38856 -7311 39178 -7310
rect 38597 -7354 38693 -7338
rect 39316 -7338 39332 -7206
rect 39396 -7106 39412 -6968
rect 40035 -6968 40131 -6952
rect 39575 -6990 39897 -6989
rect 39575 -7106 39576 -6990
rect 39396 -7206 39576 -7106
rect 39396 -7338 39418 -7206
rect 39575 -7310 39576 -7206
rect 39896 -7106 39897 -6990
rect 40035 -7106 40051 -6968
rect 39896 -7206 40051 -7106
rect 39896 -7310 39897 -7206
rect 39575 -7311 39897 -7310
rect 37150 -7652 37250 -7354
rect 37528 -7560 39072 -7460
rect 37150 -7668 37255 -7652
rect 36699 -7690 37021 -7689
rect 36699 -8010 36700 -7690
rect 37020 -7796 37021 -7690
rect 37150 -7796 37175 -7668
rect 37020 -7896 37175 -7796
rect 37020 -8010 37021 -7896
rect 37150 -8010 37175 -7896
rect 36699 -8011 37021 -8010
rect 25028 -8050 25131 -8036
rect 24316 -8056 24412 -8050
rect 25035 -8056 25131 -8050
rect 37159 -8036 37175 -8010
rect 37239 -8036 37255 -7668
rect 37528 -7689 37628 -7560
rect 37878 -7668 37974 -7652
rect 37418 -7690 37740 -7689
rect 37418 -8010 37419 -7690
rect 37739 -8010 37740 -7690
rect 37418 -8011 37740 -8010
rect 37159 -8056 37255 -8036
rect 37528 -8152 37628 -8011
rect 37878 -8036 37894 -7668
rect 37958 -8036 37974 -7668
rect 38248 -7689 38348 -7560
rect 38597 -7668 38693 -7652
rect 38137 -7690 38459 -7689
rect 38137 -8010 38138 -7690
rect 38458 -8010 38459 -7690
rect 38137 -8011 38459 -8010
rect 37878 -8056 37974 -8036
rect 38248 -8152 38348 -8011
rect 38597 -8036 38613 -7668
rect 38677 -8036 38693 -7668
rect 38970 -7689 39071 -7560
rect 39316 -7668 39418 -7338
rect 38856 -7690 39178 -7689
rect 38856 -8010 38857 -7690
rect 39177 -8010 39178 -7690
rect 38856 -8011 39178 -8010
rect 38597 -8056 38693 -8036
rect 38970 -8152 39071 -8011
rect 39316 -8036 39332 -7668
rect 39396 -7800 39418 -7668
rect 39690 -7689 39790 -7311
rect 40028 -7338 40051 -7206
rect 40115 -7338 40131 -6968
rect 40028 -7668 40131 -7338
rect 39575 -7690 39897 -7689
rect 39575 -7800 39576 -7690
rect 39396 -7900 39576 -7800
rect 39396 -8036 39418 -7900
rect 39575 -8010 39576 -7900
rect 39896 -7800 39897 -7690
rect 40028 -7800 40051 -7668
rect 39896 -7900 40051 -7800
rect 39896 -8010 39897 -7900
rect 39575 -8011 39897 -8010
rect 39690 -8012 39790 -8011
rect 39316 -8050 39418 -8036
rect 40028 -8036 40051 -7900
rect 40115 -8036 40131 -7668
rect 40028 -8050 40131 -8036
rect 39316 -8056 39412 -8050
rect 40035 -8056 40131 -8050
rect 21338 -8153 25372 -8152
rect 21338 -8251 21339 -8153
rect 21437 -8251 25273 -8153
rect 25371 -8251 25372 -8153
rect 21338 -8252 25372 -8251
rect 36338 -8153 40290 -8152
rect 36338 -8251 36339 -8153
rect 36437 -8251 40290 -8153
rect 36338 -8252 40290 -8251
rect 22159 -8368 22255 -8352
rect 22159 -8388 22175 -8368
rect 21814 -8389 21914 -8388
rect 21699 -8390 22021 -8389
rect 21699 -8710 21700 -8390
rect 22020 -8498 22021 -8390
rect 22150 -8498 22175 -8388
rect 22020 -8598 22175 -8498
rect 22020 -8710 22021 -8598
rect 21699 -8711 22021 -8710
rect 21814 -9089 21914 -8711
rect 22150 -8736 22175 -8598
rect 22239 -8736 22255 -8368
rect 22528 -8389 22628 -8252
rect 22878 -8368 22974 -8352
rect 22418 -8390 22740 -8389
rect 22418 -8710 22419 -8390
rect 22739 -8710 22740 -8390
rect 22418 -8711 22740 -8710
rect 22150 -8754 22255 -8736
rect 22150 -9052 22250 -8754
rect 22528 -8854 22628 -8711
rect 22878 -8736 22894 -8368
rect 22958 -8736 22974 -8368
rect 23248 -8389 23348 -8252
rect 23597 -8368 23693 -8352
rect 23137 -8390 23459 -8389
rect 23137 -8710 23138 -8390
rect 23458 -8710 23459 -8390
rect 23137 -8711 23459 -8710
rect 22878 -8754 22974 -8736
rect 23248 -8854 23348 -8711
rect 23597 -8736 23613 -8368
rect 23677 -8736 23693 -8368
rect 23970 -8389 24071 -8252
rect 24318 -8352 24418 -8350
rect 24316 -8368 24418 -8352
rect 23856 -8390 24178 -8389
rect 23856 -8710 23857 -8390
rect 24177 -8710 24178 -8390
rect 23856 -8711 24178 -8710
rect 23597 -8754 23693 -8736
rect 23970 -8854 24071 -8711
rect 24316 -8736 24332 -8368
rect 24396 -8504 24418 -8368
rect 25028 -8352 25128 -8350
rect 25028 -8368 25131 -8352
rect 24690 -8389 24790 -8388
rect 24575 -8390 24897 -8389
rect 24575 -8504 24576 -8390
rect 24396 -8604 24576 -8504
rect 24396 -8736 24418 -8604
rect 24575 -8710 24576 -8604
rect 24896 -8504 24897 -8390
rect 25028 -8504 25051 -8368
rect 24896 -8604 25051 -8504
rect 24896 -8710 24897 -8604
rect 24575 -8711 24897 -8710
rect 24316 -8754 24418 -8736
rect 22528 -8954 24071 -8854
rect 22150 -9068 22255 -9052
rect 21699 -9090 22021 -9089
rect 21699 -9410 21700 -9090
rect 22020 -9204 22021 -9090
rect 22150 -9204 22175 -9068
rect 22020 -9304 22175 -9204
rect 22020 -9410 22021 -9304
rect 21699 -9411 22021 -9410
rect 21814 -9789 21914 -9411
rect 22150 -9436 22175 -9304
rect 22239 -9436 22255 -9068
rect 22528 -9089 22628 -8954
rect 22878 -9068 22974 -9052
rect 22418 -9090 22740 -9089
rect 22418 -9410 22419 -9090
rect 22739 -9410 22740 -9090
rect 22418 -9411 22740 -9410
rect 22150 -9454 22255 -9436
rect 22150 -9752 22250 -9454
rect 22528 -9554 22628 -9411
rect 22878 -9436 22894 -9068
rect 22958 -9436 22974 -9068
rect 23248 -9089 23348 -8954
rect 23597 -9068 23693 -9052
rect 23137 -9090 23459 -9089
rect 23137 -9410 23138 -9090
rect 23458 -9410 23459 -9090
rect 23137 -9411 23459 -9410
rect 22878 -9454 22974 -9436
rect 23248 -9554 23348 -9411
rect 23597 -9436 23613 -9068
rect 23677 -9436 23693 -9068
rect 23970 -9089 24071 -8954
rect 24318 -9052 24418 -8754
rect 24316 -9068 24418 -9052
rect 23856 -9090 24178 -9089
rect 23856 -9410 23857 -9090
rect 24177 -9410 24178 -9090
rect 23856 -9411 24178 -9410
rect 23597 -9454 23693 -9436
rect 23970 -9554 24071 -9411
rect 24316 -9436 24332 -9068
rect 24396 -9196 24418 -9068
rect 24690 -9089 24790 -8711
rect 25028 -8736 25051 -8604
rect 25115 -8736 25131 -8368
rect 37159 -8368 37255 -8352
rect 37159 -8388 37175 -8368
rect 36814 -8389 36914 -8388
rect 36699 -8390 37021 -8389
rect 36699 -8710 36700 -8390
rect 37020 -8498 37021 -8390
rect 37150 -8498 37175 -8388
rect 37020 -8598 37175 -8498
rect 37020 -8710 37021 -8598
rect 36699 -8711 37021 -8710
rect 25028 -8754 25131 -8736
rect 25028 -9052 25128 -8754
rect 25028 -9068 25131 -9052
rect 24575 -9090 24897 -9089
rect 24575 -9196 24576 -9090
rect 24396 -9296 24576 -9196
rect 24396 -9436 24418 -9296
rect 24575 -9410 24576 -9296
rect 24896 -9196 24897 -9090
rect 25028 -9196 25051 -9068
rect 24896 -9296 25051 -9196
rect 24896 -9410 24897 -9296
rect 24575 -9411 24897 -9410
rect 22528 -9654 24072 -9554
rect 22150 -9768 22255 -9752
rect 21699 -9790 22021 -9789
rect 21699 -9850 21700 -9790
rect 9780 -9878 21700 -9850
rect 9780 -11722 9814 -9878
rect 10548 -9902 21700 -9878
rect 10548 -9988 11210 -9902
rect 11306 -9988 11790 -9902
rect 11886 -9988 12390 -9902
rect 12486 -9988 12990 -9902
rect 13086 -9988 13590 -9902
rect 13686 -9988 14190 -9902
rect 14286 -9988 14790 -9902
rect 14886 -9988 15390 -9902
rect 15486 -9988 15990 -9902
rect 16086 -9988 16590 -9902
rect 16686 -9988 17190 -9902
rect 17286 -9988 17790 -9902
rect 17886 -9988 18390 -9902
rect 18486 -9988 18990 -9902
rect 19086 -9988 19590 -9902
rect 19686 -9988 20190 -9902
rect 20286 -9988 20790 -9902
rect 20886 -9988 21700 -9902
rect 10548 -10110 21700 -9988
rect 22020 -9850 22021 -9790
rect 22150 -9850 22175 -9768
rect 22020 -10110 22175 -9850
rect 10548 -10136 22175 -10110
rect 22239 -9850 22255 -9768
rect 22878 -9768 22974 -9752
rect 22418 -9790 22740 -9789
rect 22418 -9850 22419 -9790
rect 22239 -10110 22419 -9850
rect 22739 -9850 22740 -9790
rect 22878 -9850 22894 -9768
rect 22739 -10110 22894 -9850
rect 22239 -10136 22894 -10110
rect 22958 -9850 22974 -9768
rect 23597 -9768 23693 -9752
rect 23137 -9790 23459 -9789
rect 23137 -9850 23138 -9790
rect 22958 -10110 23138 -9850
rect 23458 -9850 23459 -9790
rect 23597 -9850 23613 -9768
rect 23458 -10110 23613 -9850
rect 22958 -10136 23613 -10110
rect 23677 -9850 23693 -9768
rect 24316 -9768 24418 -9436
rect 23856 -9790 24178 -9789
rect 23856 -9850 23857 -9790
rect 23677 -10110 23857 -9850
rect 24177 -9850 24178 -9790
rect 24316 -9850 24332 -9768
rect 24177 -10110 24332 -9850
rect 23677 -10136 24332 -10110
rect 24396 -9850 24418 -9768
rect 24690 -9789 24790 -9411
rect 25028 -9436 25051 -9296
rect 25115 -9436 25131 -9068
rect 36814 -9089 36914 -8711
rect 37150 -8736 37175 -8598
rect 37239 -8736 37255 -8368
rect 37528 -8389 37628 -8252
rect 37878 -8368 37974 -8352
rect 37418 -8390 37740 -8389
rect 37418 -8710 37419 -8390
rect 37739 -8710 37740 -8390
rect 37418 -8711 37740 -8710
rect 37150 -8754 37255 -8736
rect 37150 -9052 37250 -8754
rect 37528 -8854 37628 -8711
rect 37878 -8736 37894 -8368
rect 37958 -8736 37974 -8368
rect 38248 -8389 38348 -8252
rect 38597 -8368 38693 -8352
rect 38137 -8390 38459 -8389
rect 38137 -8710 38138 -8390
rect 38458 -8710 38459 -8390
rect 38137 -8711 38459 -8710
rect 37878 -8754 37974 -8736
rect 38248 -8854 38348 -8711
rect 38597 -8736 38613 -8368
rect 38677 -8736 38693 -8368
rect 38970 -8389 39071 -8252
rect 39318 -8352 39418 -8350
rect 39316 -8368 39418 -8352
rect 38856 -8390 39178 -8389
rect 38856 -8710 38857 -8390
rect 39177 -8710 39178 -8390
rect 38856 -8711 39178 -8710
rect 38597 -8754 38693 -8736
rect 38970 -8854 39071 -8711
rect 39316 -8736 39332 -8368
rect 39396 -8504 39418 -8368
rect 40028 -8352 40128 -8350
rect 40028 -8368 40131 -8352
rect 39690 -8389 39790 -8388
rect 39575 -8390 39897 -8389
rect 39575 -8504 39576 -8390
rect 39396 -8604 39576 -8504
rect 39396 -8736 39418 -8604
rect 39575 -8710 39576 -8604
rect 39896 -8504 39897 -8390
rect 40028 -8504 40051 -8368
rect 39896 -8604 40051 -8504
rect 39896 -8710 39897 -8604
rect 39575 -8711 39897 -8710
rect 39316 -8754 39418 -8736
rect 37528 -8954 39071 -8854
rect 37150 -9068 37255 -9052
rect 36699 -9090 37021 -9089
rect 36699 -9410 36700 -9090
rect 37020 -9204 37021 -9090
rect 37150 -9204 37175 -9068
rect 37020 -9304 37175 -9204
rect 37020 -9410 37021 -9304
rect 36699 -9411 37021 -9410
rect 25028 -9768 25131 -9436
rect 24575 -9790 24897 -9789
rect 24575 -9850 24576 -9790
rect 24396 -10110 24576 -9850
rect 24896 -9850 24897 -9790
rect 25028 -9850 25051 -9768
rect 24896 -10110 25051 -9850
rect 24396 -10136 25051 -10110
rect 25115 -9850 25131 -9768
rect 36814 -9789 36914 -9411
rect 37150 -9436 37175 -9304
rect 37239 -9436 37255 -9068
rect 37528 -9089 37628 -8954
rect 37878 -9068 37974 -9052
rect 37418 -9090 37740 -9089
rect 37418 -9410 37419 -9090
rect 37739 -9410 37740 -9090
rect 37418 -9411 37740 -9410
rect 37150 -9454 37255 -9436
rect 37150 -9752 37250 -9454
rect 37528 -9554 37628 -9411
rect 37878 -9436 37894 -9068
rect 37958 -9436 37974 -9068
rect 38248 -9089 38348 -8954
rect 38597 -9068 38693 -9052
rect 38137 -9090 38459 -9089
rect 38137 -9410 38138 -9090
rect 38458 -9410 38459 -9090
rect 38137 -9411 38459 -9410
rect 37878 -9454 37974 -9436
rect 38248 -9554 38348 -9411
rect 38597 -9436 38613 -9068
rect 38677 -9436 38693 -9068
rect 38970 -9089 39071 -8954
rect 39318 -9052 39418 -8754
rect 39316 -9068 39418 -9052
rect 38856 -9090 39178 -9089
rect 38856 -9410 38857 -9090
rect 39177 -9410 39178 -9090
rect 38856 -9411 39178 -9410
rect 38597 -9454 38693 -9436
rect 38970 -9554 39071 -9411
rect 39316 -9436 39332 -9068
rect 39396 -9196 39418 -9068
rect 39690 -9089 39790 -8711
rect 40028 -8736 40051 -8604
rect 40115 -8736 40131 -8368
rect 40028 -8754 40131 -8736
rect 40028 -9052 40128 -8754
rect 40028 -9068 40131 -9052
rect 39575 -9090 39897 -9089
rect 39575 -9196 39576 -9090
rect 39396 -9296 39576 -9196
rect 39396 -9436 39418 -9296
rect 39575 -9410 39576 -9296
rect 39896 -9196 39897 -9090
rect 40028 -9196 40051 -9068
rect 39896 -9296 40051 -9196
rect 39896 -9410 39897 -9296
rect 39575 -9411 39897 -9410
rect 37528 -9654 39072 -9554
rect 37150 -9768 37255 -9752
rect 36699 -9790 37021 -9789
rect 36699 -9850 36700 -9790
rect 25115 -9902 36700 -9850
rect 25115 -9988 26210 -9902
rect 26306 -9988 26790 -9902
rect 26886 -9988 27390 -9902
rect 27486 -9988 27990 -9902
rect 28086 -9988 28590 -9902
rect 28686 -9988 29190 -9902
rect 29286 -9988 29790 -9902
rect 29886 -9988 30390 -9902
rect 30486 -9988 30990 -9902
rect 31086 -9988 31590 -9902
rect 31686 -9988 32190 -9902
rect 32286 -9988 32790 -9902
rect 32886 -9988 33390 -9902
rect 33486 -9988 33990 -9902
rect 34086 -9988 34590 -9902
rect 34686 -9988 35190 -9902
rect 35286 -9988 35790 -9902
rect 35886 -9988 36700 -9902
rect 25115 -10110 36700 -9988
rect 37020 -9850 37021 -9790
rect 37150 -9850 37175 -9768
rect 37020 -10110 37175 -9850
rect 25115 -10136 37175 -10110
rect 37239 -9850 37255 -9768
rect 37878 -9768 37974 -9752
rect 37418 -9790 37740 -9789
rect 37418 -9850 37419 -9790
rect 37239 -10110 37419 -9850
rect 37739 -9850 37740 -9790
rect 37878 -9850 37894 -9768
rect 37739 -10110 37894 -9850
rect 37239 -10136 37894 -10110
rect 37958 -9850 37974 -9768
rect 38597 -9768 38693 -9752
rect 38137 -9790 38459 -9789
rect 38137 -9850 38138 -9790
rect 37958 -10110 38138 -9850
rect 38458 -9850 38459 -9790
rect 38597 -9850 38613 -9768
rect 38458 -10110 38613 -9850
rect 37958 -10136 38613 -10110
rect 38677 -9850 38693 -9768
rect 39316 -9768 39418 -9436
rect 38856 -9790 39178 -9789
rect 38856 -9850 38857 -9790
rect 38677 -10110 38857 -9850
rect 39177 -9850 39178 -9790
rect 39316 -9850 39332 -9768
rect 39177 -10110 39332 -9850
rect 38677 -10136 39332 -10110
rect 39396 -9850 39418 -9768
rect 39690 -9789 39790 -9411
rect 40028 -9436 40051 -9296
rect 40115 -9436 40131 -9068
rect 40028 -9768 40131 -9436
rect 39575 -9790 39897 -9789
rect 39575 -9850 39576 -9790
rect 39396 -10110 39576 -9850
rect 39896 -9850 39897 -9790
rect 40028 -9850 40051 -9768
rect 39896 -10110 40051 -9850
rect 39396 -10136 40051 -10110
rect 40115 -9850 40131 -9768
rect 40115 -9856 40288 -9850
rect 40115 -10136 40292 -9856
rect 10548 -10166 40292 -10136
rect 10548 -10466 10924 -10166
rect 11524 -10466 20556 -10166
rect 21156 -10466 25924 -10166
rect 26524 -10466 35556 -10166
rect 36156 -10466 40292 -10166
rect 10548 -10954 40292 -10466
rect 10548 -11138 40294 -10954
rect 10548 -11438 14878 -11138
rect 15478 -11438 24510 -11138
rect 25110 -11438 29878 -11138
rect 30478 -11438 39510 -11138
rect 40110 -11438 40294 -11138
rect 10548 -11468 40294 -11438
rect 10548 -11722 10919 -11468
rect 9780 -11754 10919 -11722
rect 10903 -11836 10919 -11754
rect 10983 -11494 11638 -11468
rect 10983 -11754 11138 -11494
rect 10983 -11836 11006 -11754
rect 11137 -11814 11138 -11754
rect 11458 -11754 11638 -11494
rect 11458 -11814 11459 -11754
rect 11137 -11815 11459 -11814
rect 10903 -12168 11006 -11836
rect 10903 -12536 10919 -12168
rect 10983 -12308 11006 -12168
rect 11244 -12193 11344 -11815
rect 11616 -11836 11638 -11754
rect 11702 -11494 12357 -11468
rect 11702 -11754 11857 -11494
rect 11702 -11836 11718 -11754
rect 11856 -11814 11857 -11754
rect 12177 -11754 12357 -11494
rect 12177 -11814 12178 -11754
rect 11856 -11815 12178 -11814
rect 11616 -12168 11718 -11836
rect 12341 -11836 12357 -11754
rect 12421 -11494 13076 -11468
rect 12421 -11754 12576 -11494
rect 12421 -11836 12437 -11754
rect 12575 -11814 12576 -11754
rect 12896 -11754 13076 -11494
rect 12896 -11814 12897 -11754
rect 12575 -11815 12897 -11814
rect 12341 -11852 12437 -11836
rect 13060 -11836 13076 -11754
rect 13140 -11494 13795 -11468
rect 13140 -11754 13295 -11494
rect 13140 -11836 13156 -11754
rect 13294 -11814 13295 -11754
rect 13615 -11754 13795 -11494
rect 13615 -11814 13616 -11754
rect 13294 -11815 13616 -11814
rect 13060 -11852 13156 -11836
rect 13779 -11836 13795 -11754
rect 13859 -11494 25919 -11468
rect 13859 -11754 14014 -11494
rect 13859 -11836 13884 -11754
rect 14013 -11814 14014 -11754
rect 14334 -11616 25919 -11494
rect 14334 -11702 15148 -11616
rect 15244 -11702 15748 -11616
rect 15844 -11702 16348 -11616
rect 16444 -11702 16948 -11616
rect 17044 -11702 17548 -11616
rect 17644 -11702 18148 -11616
rect 18244 -11702 18748 -11616
rect 18844 -11702 19348 -11616
rect 19444 -11702 19948 -11616
rect 20044 -11702 20548 -11616
rect 20644 -11702 21148 -11616
rect 21244 -11702 21748 -11616
rect 21844 -11702 22348 -11616
rect 22444 -11702 22948 -11616
rect 23044 -11702 23548 -11616
rect 23644 -11702 24148 -11616
rect 24244 -11702 24728 -11616
rect 24824 -11702 25919 -11616
rect 14334 -11754 25919 -11702
rect 14334 -11814 14335 -11754
rect 14013 -11815 14335 -11814
rect 13779 -11852 13884 -11836
rect 11962 -12050 13506 -11950
rect 11137 -12194 11459 -12193
rect 11137 -12308 11138 -12194
rect 10983 -12408 11138 -12308
rect 10983 -12536 11006 -12408
rect 11137 -12514 11138 -12408
rect 11458 -12308 11459 -12194
rect 11616 -12308 11638 -12168
rect 11458 -12408 11638 -12308
rect 11458 -12514 11459 -12408
rect 11137 -12515 11459 -12514
rect 10903 -12552 11006 -12536
rect 10906 -12850 11006 -12552
rect 10903 -12868 11006 -12850
rect 10903 -13236 10919 -12868
rect 10983 -13000 11006 -12868
rect 11244 -12893 11344 -12515
rect 11616 -12536 11638 -12408
rect 11702 -12536 11718 -12168
rect 11963 -12193 12064 -12050
rect 12341 -12168 12437 -12150
rect 11856 -12194 12178 -12193
rect 11856 -12514 11857 -12194
rect 12177 -12514 12178 -12194
rect 11856 -12515 12178 -12514
rect 11616 -12552 11718 -12536
rect 11616 -12850 11716 -12552
rect 11963 -12650 12064 -12515
rect 12341 -12536 12357 -12168
rect 12421 -12536 12437 -12168
rect 12686 -12193 12786 -12050
rect 13060 -12168 13156 -12150
rect 12575 -12194 12897 -12193
rect 12575 -12514 12576 -12194
rect 12896 -12514 12897 -12194
rect 12575 -12515 12897 -12514
rect 12341 -12552 12437 -12536
rect 12686 -12650 12786 -12515
rect 13060 -12536 13076 -12168
rect 13140 -12536 13156 -12168
rect 13406 -12193 13506 -12050
rect 13784 -12150 13884 -11852
rect 13779 -12168 13884 -12150
rect 13294 -12194 13616 -12193
rect 13294 -12514 13295 -12194
rect 13615 -12514 13616 -12194
rect 13294 -12515 13616 -12514
rect 13060 -12552 13156 -12536
rect 13406 -12650 13506 -12515
rect 13779 -12536 13795 -12168
rect 13859 -12300 13884 -12168
rect 14120 -12193 14220 -11815
rect 25903 -11836 25919 -11754
rect 25983 -11494 26638 -11468
rect 25983 -11754 26138 -11494
rect 25983 -11836 26006 -11754
rect 26137 -11814 26138 -11754
rect 26458 -11754 26638 -11494
rect 26458 -11814 26459 -11754
rect 26137 -11815 26459 -11814
rect 25903 -12168 26006 -11836
rect 14013 -12194 14335 -12193
rect 14013 -12300 14014 -12194
rect 13859 -12400 14014 -12300
rect 13859 -12536 13884 -12400
rect 14013 -12514 14014 -12400
rect 14334 -12514 14335 -12194
rect 14013 -12515 14335 -12514
rect 13779 -12552 13884 -12536
rect 11963 -12750 13506 -12650
rect 11616 -12868 11718 -12850
rect 11137 -12894 11459 -12893
rect 11137 -13000 11138 -12894
rect 10983 -13100 11138 -13000
rect 10983 -13236 11006 -13100
rect 11137 -13214 11138 -13100
rect 11458 -13000 11459 -12894
rect 11616 -13000 11638 -12868
rect 11458 -13100 11638 -13000
rect 11458 -13214 11459 -13100
rect 11137 -13215 11459 -13214
rect 11244 -13216 11344 -13215
rect 10903 -13252 11006 -13236
rect 10906 -13254 11006 -13252
rect 11616 -13236 11638 -13100
rect 11702 -13236 11718 -12868
rect 11963 -12893 12064 -12750
rect 12341 -12868 12437 -12850
rect 11856 -12894 12178 -12893
rect 11856 -13214 11857 -12894
rect 12177 -13214 12178 -12894
rect 11856 -13215 12178 -13214
rect 11616 -13252 11718 -13236
rect 11616 -13254 11716 -13252
rect 11963 -13352 12064 -13215
rect 12341 -13236 12357 -12868
rect 12421 -13236 12437 -12868
rect 12686 -12893 12786 -12750
rect 13060 -12868 13156 -12850
rect 12575 -12894 12897 -12893
rect 12575 -13214 12576 -12894
rect 12896 -13214 12897 -12894
rect 12575 -13215 12897 -13214
rect 12341 -13252 12437 -13236
rect 12686 -13352 12786 -13215
rect 13060 -13236 13076 -12868
rect 13140 -13236 13156 -12868
rect 13406 -12893 13506 -12750
rect 13784 -12850 13884 -12552
rect 13779 -12868 13884 -12850
rect 13294 -12894 13616 -12893
rect 13294 -13214 13295 -12894
rect 13615 -13214 13616 -12894
rect 13294 -13215 13616 -13214
rect 13060 -13252 13156 -13236
rect 13406 -13352 13506 -13215
rect 13779 -13236 13795 -12868
rect 13859 -13006 13884 -12868
rect 14120 -12893 14220 -12515
rect 25903 -12536 25919 -12168
rect 25983 -12308 26006 -12168
rect 26244 -12193 26344 -11815
rect 26616 -11836 26638 -11754
rect 26702 -11494 27357 -11468
rect 26702 -11754 26857 -11494
rect 26702 -11836 26718 -11754
rect 26856 -11814 26857 -11754
rect 27177 -11754 27357 -11494
rect 27177 -11814 27178 -11754
rect 26856 -11815 27178 -11814
rect 26616 -12168 26718 -11836
rect 27341 -11836 27357 -11754
rect 27421 -11494 28076 -11468
rect 27421 -11754 27576 -11494
rect 27421 -11836 27437 -11754
rect 27575 -11814 27576 -11754
rect 27896 -11754 28076 -11494
rect 27896 -11814 27897 -11754
rect 27575 -11815 27897 -11814
rect 27341 -11852 27437 -11836
rect 28060 -11836 28076 -11754
rect 28140 -11494 28795 -11468
rect 28140 -11754 28295 -11494
rect 28140 -11836 28156 -11754
rect 28294 -11814 28295 -11754
rect 28615 -11754 28795 -11494
rect 28615 -11814 28616 -11754
rect 28294 -11815 28616 -11814
rect 28060 -11852 28156 -11836
rect 28779 -11836 28795 -11754
rect 28859 -11494 40294 -11468
rect 28859 -11754 29014 -11494
rect 28859 -11836 28884 -11754
rect 29013 -11814 29014 -11754
rect 29334 -11616 40294 -11494
rect 29334 -11702 30148 -11616
rect 30244 -11702 30748 -11616
rect 30844 -11702 31348 -11616
rect 31444 -11702 31948 -11616
rect 32044 -11702 32548 -11616
rect 32644 -11702 33148 -11616
rect 33244 -11702 33748 -11616
rect 33844 -11702 34348 -11616
rect 34444 -11702 34948 -11616
rect 35044 -11702 35548 -11616
rect 35644 -11702 36148 -11616
rect 36244 -11702 36748 -11616
rect 36844 -11702 37348 -11616
rect 37444 -11702 37948 -11616
rect 38044 -11702 38548 -11616
rect 38644 -11702 39148 -11616
rect 39244 -11702 39728 -11616
rect 39824 -11702 40294 -11616
rect 29334 -11754 40294 -11702
rect 29334 -11814 29335 -11754
rect 29013 -11815 29335 -11814
rect 28779 -11852 28884 -11836
rect 26962 -12050 28506 -11950
rect 26137 -12194 26459 -12193
rect 26137 -12308 26138 -12194
rect 25983 -12408 26138 -12308
rect 25983 -12536 26006 -12408
rect 26137 -12514 26138 -12408
rect 26458 -12308 26459 -12194
rect 26616 -12308 26638 -12168
rect 26458 -12408 26638 -12308
rect 26458 -12514 26459 -12408
rect 26137 -12515 26459 -12514
rect 25903 -12552 26006 -12536
rect 25906 -12850 26006 -12552
rect 25903 -12868 26006 -12850
rect 14013 -12894 14335 -12893
rect 14013 -13006 14014 -12894
rect 13859 -13106 14014 -13006
rect 13859 -13216 13884 -13106
rect 14013 -13214 14014 -13106
rect 14334 -13214 14335 -12894
rect 14013 -13215 14335 -13214
rect 14120 -13216 14220 -13215
rect 13859 -13236 13875 -13216
rect 13779 -13252 13875 -13236
rect 25903 -13236 25919 -12868
rect 25983 -13000 26006 -12868
rect 26244 -12893 26344 -12515
rect 26616 -12536 26638 -12408
rect 26702 -12536 26718 -12168
rect 26963 -12193 27064 -12050
rect 27341 -12168 27437 -12150
rect 26856 -12194 27178 -12193
rect 26856 -12514 26857 -12194
rect 27177 -12514 27178 -12194
rect 26856 -12515 27178 -12514
rect 26616 -12552 26718 -12536
rect 26616 -12850 26716 -12552
rect 26963 -12650 27064 -12515
rect 27341 -12536 27357 -12168
rect 27421 -12536 27437 -12168
rect 27686 -12193 27786 -12050
rect 28060 -12168 28156 -12150
rect 27575 -12194 27897 -12193
rect 27575 -12514 27576 -12194
rect 27896 -12514 27897 -12194
rect 27575 -12515 27897 -12514
rect 27341 -12552 27437 -12536
rect 27686 -12650 27786 -12515
rect 28060 -12536 28076 -12168
rect 28140 -12536 28156 -12168
rect 28406 -12193 28506 -12050
rect 28784 -12150 28884 -11852
rect 28779 -12168 28884 -12150
rect 28294 -12194 28616 -12193
rect 28294 -12514 28295 -12194
rect 28615 -12514 28616 -12194
rect 28294 -12515 28616 -12514
rect 28060 -12552 28156 -12536
rect 28406 -12650 28506 -12515
rect 28779 -12536 28795 -12168
rect 28859 -12300 28884 -12168
rect 29120 -12193 29220 -11815
rect 29013 -12194 29335 -12193
rect 29013 -12300 29014 -12194
rect 28859 -12400 29014 -12300
rect 28859 -12536 28884 -12400
rect 29013 -12514 29014 -12400
rect 29334 -12514 29335 -12194
rect 29013 -12515 29335 -12514
rect 28779 -12552 28884 -12536
rect 26963 -12750 28506 -12650
rect 26616 -12868 26718 -12850
rect 26137 -12894 26459 -12893
rect 26137 -13000 26138 -12894
rect 25983 -13100 26138 -13000
rect 25983 -13236 26006 -13100
rect 26137 -13214 26138 -13100
rect 26458 -13000 26459 -12894
rect 26616 -13000 26638 -12868
rect 26458 -13100 26638 -13000
rect 26458 -13214 26459 -13100
rect 26137 -13215 26459 -13214
rect 26244 -13216 26344 -13215
rect 25903 -13252 26006 -13236
rect 25906 -13254 26006 -13252
rect 26616 -13236 26638 -13100
rect 26702 -13236 26718 -12868
rect 26963 -12893 27064 -12750
rect 27341 -12868 27437 -12850
rect 26856 -12894 27178 -12893
rect 26856 -13214 26857 -12894
rect 27177 -13214 27178 -12894
rect 26856 -13215 27178 -13214
rect 26616 -13252 26718 -13236
rect 26616 -13254 26716 -13252
rect 26963 -13352 27064 -13215
rect 27341 -13236 27357 -12868
rect 27421 -13236 27437 -12868
rect 27686 -12893 27786 -12750
rect 28060 -12868 28156 -12850
rect 27575 -12894 27897 -12893
rect 27575 -13214 27576 -12894
rect 27896 -13214 27897 -12894
rect 27575 -13215 27897 -13214
rect 27341 -13252 27437 -13236
rect 27686 -13352 27786 -13215
rect 28060 -13236 28076 -12868
rect 28140 -13236 28156 -12868
rect 28406 -12893 28506 -12750
rect 28784 -12850 28884 -12552
rect 28779 -12868 28884 -12850
rect 28294 -12894 28616 -12893
rect 28294 -13214 28295 -12894
rect 28615 -13214 28616 -12894
rect 28294 -13215 28616 -13214
rect 28060 -13252 28156 -13236
rect 28406 -13352 28506 -13215
rect 28779 -13236 28795 -12868
rect 28859 -13006 28884 -12868
rect 29120 -12893 29220 -12515
rect 29013 -12894 29335 -12893
rect 29013 -13006 29014 -12894
rect 28859 -13106 29014 -13006
rect 28859 -13216 28884 -13106
rect 29013 -13214 29014 -13106
rect 29334 -13214 29335 -12894
rect 29013 -13215 29335 -13214
rect 29120 -13216 29220 -13215
rect 28859 -13236 28875 -13216
rect 28779 -13252 28875 -13236
rect 10604 -13353 14696 -13352
rect 10604 -13451 10605 -13353
rect 10703 -13451 14597 -13353
rect 14695 -13451 14696 -13353
rect 10604 -13452 14696 -13451
rect 25596 -13353 29696 -13352
rect 25596 -13451 25597 -13353
rect 25695 -13451 29597 -13353
rect 29695 -13451 29696 -13353
rect 25596 -13452 29696 -13451
rect 10903 -13554 10999 -13548
rect 11622 -13554 11718 -13548
rect 10903 -13568 11006 -13554
rect 10903 -13936 10919 -13568
rect 10983 -13704 11006 -13568
rect 11616 -13568 11718 -13554
rect 11244 -13593 11344 -13592
rect 11137 -13594 11459 -13593
rect 11137 -13704 11138 -13594
rect 10983 -13804 11138 -13704
rect 10983 -13936 11006 -13804
rect 11137 -13914 11138 -13804
rect 11458 -13704 11459 -13594
rect 11616 -13704 11638 -13568
rect 11458 -13804 11638 -13704
rect 11458 -13914 11459 -13804
rect 11137 -13915 11459 -13914
rect 10903 -14266 11006 -13936
rect 10903 -14636 10919 -14266
rect 10983 -14398 11006 -14266
rect 11244 -14293 11344 -13915
rect 11616 -13936 11638 -13804
rect 11702 -13936 11718 -13568
rect 11963 -13593 12064 -13452
rect 12341 -13568 12437 -13548
rect 11856 -13594 12178 -13593
rect 11856 -13914 11857 -13594
rect 12177 -13914 12178 -13594
rect 11856 -13915 12178 -13914
rect 11616 -14266 11718 -13936
rect 11963 -14044 12064 -13915
rect 12341 -13936 12357 -13568
rect 12421 -13936 12437 -13568
rect 12686 -13593 12786 -13452
rect 13060 -13568 13156 -13548
rect 12575 -13594 12897 -13593
rect 12575 -13914 12576 -13594
rect 12896 -13914 12897 -13594
rect 12575 -13915 12897 -13914
rect 12341 -13952 12437 -13936
rect 12686 -14044 12786 -13915
rect 13060 -13936 13076 -13568
rect 13140 -13936 13156 -13568
rect 13406 -13593 13506 -13452
rect 13779 -13568 13875 -13548
rect 13294 -13594 13616 -13593
rect 13294 -13914 13295 -13594
rect 13615 -13914 13616 -13594
rect 13294 -13915 13616 -13914
rect 13060 -13952 13156 -13936
rect 13406 -14044 13506 -13915
rect 13779 -13936 13795 -13568
rect 13859 -13594 13875 -13568
rect 25903 -13554 25999 -13548
rect 26622 -13554 26718 -13548
rect 25903 -13568 26006 -13554
rect 14013 -13594 14335 -13593
rect 13859 -13708 13884 -13594
rect 14013 -13708 14014 -13594
rect 13859 -13808 14014 -13708
rect 13859 -13936 13884 -13808
rect 14013 -13914 14014 -13808
rect 14334 -13914 14335 -13594
rect 14013 -13915 14335 -13914
rect 13779 -13952 13884 -13936
rect 11962 -14144 13506 -14044
rect 13784 -14250 13884 -13952
rect 11137 -14294 11459 -14293
rect 11137 -14398 11138 -14294
rect 10983 -14498 11138 -14398
rect 10983 -14636 10999 -14498
rect 11137 -14614 11138 -14498
rect 11458 -14398 11459 -14294
rect 11616 -14398 11638 -14266
rect 11458 -14498 11638 -14398
rect 11458 -14614 11459 -14498
rect 11137 -14615 11459 -14614
rect 10903 -14652 10999 -14636
rect 11622 -14636 11638 -14498
rect 11702 -14398 11718 -14266
rect 12341 -14266 12437 -14250
rect 11856 -14294 12178 -14293
rect 11856 -14398 11857 -14294
rect 11702 -14498 11857 -14398
rect 11702 -14636 11718 -14498
rect 11856 -14614 11857 -14498
rect 12177 -14398 12178 -14294
rect 12341 -14398 12357 -14266
rect 12177 -14498 12357 -14398
rect 12177 -14614 12178 -14498
rect 11856 -14615 12178 -14614
rect 11622 -14652 11718 -14636
rect 12341 -14636 12357 -14498
rect 12421 -14398 12437 -14266
rect 13060 -14266 13156 -14250
rect 12575 -14294 12897 -14293
rect 12575 -14398 12576 -14294
rect 12421 -14498 12576 -14398
rect 12421 -14636 12437 -14498
rect 12575 -14614 12576 -14498
rect 12896 -14398 12897 -14294
rect 13060 -14398 13076 -14266
rect 12896 -14498 13076 -14398
rect 12896 -14614 12897 -14498
rect 12575 -14615 12897 -14614
rect 12341 -14652 12437 -14636
rect 13060 -14636 13076 -14498
rect 13140 -14398 13156 -14266
rect 13779 -14266 13884 -14250
rect 13294 -14294 13616 -14293
rect 13294 -14398 13295 -14294
rect 13140 -14498 13295 -14398
rect 13140 -14636 13156 -14498
rect 13294 -14614 13295 -14498
rect 13615 -14398 13616 -14294
rect 13779 -14398 13795 -14266
rect 13615 -14498 13795 -14398
rect 13615 -14614 13616 -14498
rect 13294 -14615 13616 -14614
rect 13060 -14652 13156 -14636
rect 13779 -14638 13795 -14498
rect 13859 -14398 13884 -14266
rect 14120 -14293 14220 -13915
rect 25903 -13936 25919 -13568
rect 25983 -13704 26006 -13568
rect 26616 -13568 26718 -13554
rect 26244 -13593 26344 -13592
rect 26137 -13594 26459 -13593
rect 26137 -13704 26138 -13594
rect 25983 -13804 26138 -13704
rect 25983 -13936 26006 -13804
rect 26137 -13914 26138 -13804
rect 26458 -13704 26459 -13594
rect 26616 -13704 26638 -13568
rect 26458 -13804 26638 -13704
rect 26458 -13914 26459 -13804
rect 26137 -13915 26459 -13914
rect 25903 -14266 26006 -13936
rect 14013 -14294 14335 -14293
rect 14013 -14398 14014 -14294
rect 13859 -14498 14014 -14398
rect 13859 -14638 13875 -14498
rect 14013 -14614 14014 -14498
rect 14334 -14614 14335 -14294
rect 14013 -14615 14335 -14614
rect 13779 -14654 13875 -14638
rect 25903 -14636 25919 -14266
rect 25983 -14398 26006 -14266
rect 26244 -14293 26344 -13915
rect 26616 -13936 26638 -13804
rect 26702 -13936 26718 -13568
rect 26963 -13593 27064 -13452
rect 27341 -13568 27437 -13548
rect 26856 -13594 27178 -13593
rect 26856 -13914 26857 -13594
rect 27177 -13914 27178 -13594
rect 26856 -13915 27178 -13914
rect 26616 -14266 26718 -13936
rect 26963 -14044 27064 -13915
rect 27341 -13936 27357 -13568
rect 27421 -13936 27437 -13568
rect 27686 -13593 27786 -13452
rect 28060 -13568 28156 -13548
rect 27575 -13594 27897 -13593
rect 27575 -13914 27576 -13594
rect 27896 -13914 27897 -13594
rect 27575 -13915 27897 -13914
rect 27341 -13952 27437 -13936
rect 27686 -14044 27786 -13915
rect 28060 -13936 28076 -13568
rect 28140 -13936 28156 -13568
rect 28406 -13593 28506 -13452
rect 28779 -13568 28875 -13548
rect 28294 -13594 28616 -13593
rect 28294 -13914 28295 -13594
rect 28615 -13914 28616 -13594
rect 28294 -13915 28616 -13914
rect 28060 -13952 28156 -13936
rect 28406 -14044 28506 -13915
rect 28779 -13936 28795 -13568
rect 28859 -13594 28875 -13568
rect 29013 -13594 29335 -13593
rect 28859 -13708 28884 -13594
rect 29013 -13708 29014 -13594
rect 28859 -13808 29014 -13708
rect 28859 -13936 28884 -13808
rect 29013 -13914 29014 -13808
rect 29334 -13914 29335 -13594
rect 29013 -13915 29335 -13914
rect 28779 -13952 28884 -13936
rect 26962 -14144 28506 -14044
rect 28784 -14250 28884 -13952
rect 26137 -14294 26459 -14293
rect 26137 -14398 26138 -14294
rect 25983 -14498 26138 -14398
rect 25983 -14636 25999 -14498
rect 26137 -14614 26138 -14498
rect 26458 -14398 26459 -14294
rect 26616 -14398 26638 -14266
rect 26458 -14498 26638 -14398
rect 26458 -14614 26459 -14498
rect 26137 -14615 26459 -14614
rect 25903 -14652 25999 -14636
rect 26622 -14636 26638 -14498
rect 26702 -14398 26718 -14266
rect 27341 -14266 27437 -14250
rect 26856 -14294 27178 -14293
rect 26856 -14398 26857 -14294
rect 26702 -14498 26857 -14398
rect 26702 -14636 26718 -14498
rect 26856 -14614 26857 -14498
rect 27177 -14398 27178 -14294
rect 27341 -14398 27357 -14266
rect 27177 -14498 27357 -14398
rect 27177 -14614 27178 -14498
rect 26856 -14615 27178 -14614
rect 26622 -14652 26718 -14636
rect 27341 -14636 27357 -14498
rect 27421 -14398 27437 -14266
rect 28060 -14266 28156 -14250
rect 27575 -14294 27897 -14293
rect 27575 -14398 27576 -14294
rect 27421 -14498 27576 -14398
rect 27421 -14636 27437 -14498
rect 27575 -14614 27576 -14498
rect 27896 -14398 27897 -14294
rect 28060 -14398 28076 -14266
rect 27896 -14498 28076 -14398
rect 27896 -14614 27897 -14498
rect 27575 -14615 27897 -14614
rect 27341 -14652 27437 -14636
rect 28060 -14636 28076 -14498
rect 28140 -14398 28156 -14266
rect 28779 -14266 28884 -14250
rect 28294 -14294 28616 -14293
rect 28294 -14398 28295 -14294
rect 28140 -14498 28295 -14398
rect 28140 -14636 28156 -14498
rect 28294 -14614 28295 -14498
rect 28615 -14398 28616 -14294
rect 28779 -14398 28795 -14266
rect 28615 -14498 28795 -14398
rect 28615 -14614 28616 -14498
rect 28294 -14615 28616 -14614
rect 28060 -14652 28156 -14636
rect 28779 -14638 28795 -14498
rect 28859 -14398 28884 -14266
rect 29120 -14293 29220 -13915
rect 29013 -14294 29335 -14293
rect 29013 -14398 29014 -14294
rect 28859 -14498 29014 -14398
rect 28859 -14638 28875 -14498
rect 29013 -14614 29014 -14498
rect 29334 -14614 29335 -14294
rect 29013 -14615 29335 -14614
rect 28779 -14654 28875 -14638
rect 10740 -18880 41204 -18850
rect 10740 -18910 40432 -18880
rect 10740 -18996 15942 -18910
rect 16038 -18996 16362 -18910
rect 16458 -18996 16962 -18910
rect 17058 -18996 17562 -18910
rect 17658 -18996 18162 -18910
rect 18258 -18996 18762 -18910
rect 18858 -18996 19362 -18910
rect 19458 -18996 19962 -18910
rect 20058 -18996 20562 -18910
rect 20658 -18996 21162 -18910
rect 21258 -18996 21762 -18910
rect 21858 -18996 22362 -18910
rect 22458 -18996 22962 -18910
rect 23058 -18996 23562 -18910
rect 23658 -18996 24162 -18910
rect 24258 -18996 30942 -18910
rect 31038 -18996 31362 -18910
rect 31458 -18996 31962 -18910
rect 32058 -18996 32562 -18910
rect 32658 -18996 33162 -18910
rect 33258 -18996 33762 -18910
rect 33858 -18996 34362 -18910
rect 34458 -18996 34962 -18910
rect 35058 -18996 35562 -18910
rect 35658 -18996 36162 -18910
rect 36258 -18996 36762 -18910
rect 36858 -18996 37362 -18910
rect 37458 -18996 37962 -18910
rect 38058 -18996 38562 -18910
rect 38658 -18996 39162 -18910
rect 39258 -18996 40432 -18910
rect 10740 -19170 40432 -18996
rect 10740 -19470 14878 -19170
rect 15478 -19470 24510 -19170
rect 25110 -19470 29878 -19170
rect 30478 -19470 39510 -19170
rect 40110 -19470 40432 -19170
rect 10740 -20134 40432 -19470
rect 10740 -20434 10924 -20134
rect 11524 -20434 20556 -20134
rect 21156 -20434 25924 -20134
rect 26524 -20434 35556 -20134
rect 36156 -20434 40432 -20134
rect 10740 -20608 40432 -20434
rect 10740 -20694 11776 -20608
rect 11872 -20694 12376 -20608
rect 12472 -20694 12976 -20608
rect 13072 -20694 13576 -20608
rect 13672 -20694 14176 -20608
rect 14272 -20694 14776 -20608
rect 14872 -20694 15376 -20608
rect 15472 -20694 15976 -20608
rect 16072 -20694 16576 -20608
rect 16672 -20694 17176 -20608
rect 17272 -20694 17776 -20608
rect 17872 -20694 18376 -20608
rect 18472 -20694 18976 -20608
rect 19072 -20694 19576 -20608
rect 19672 -20694 19996 -20608
rect 20092 -20694 26776 -20608
rect 26872 -20694 27376 -20608
rect 27472 -20694 27976 -20608
rect 28072 -20694 28576 -20608
rect 28672 -20694 29176 -20608
rect 29272 -20694 29776 -20608
rect 29872 -20694 30376 -20608
rect 30472 -20694 30976 -20608
rect 31072 -20694 31576 -20608
rect 31672 -20694 32176 -20608
rect 32272 -20694 32776 -20608
rect 32872 -20694 33376 -20608
rect 33472 -20694 33976 -20608
rect 34072 -20694 34576 -20608
rect 34672 -20694 34996 -20608
rect 35092 -20694 40432 -20608
rect 10740 -20726 40432 -20694
rect 41166 -20726 41204 -18880
rect 10740 -20752 41204 -20726
rect 22159 -24966 22255 -24950
rect 21699 -24990 22021 -24989
rect 21699 -25310 21700 -24990
rect 22020 -25106 22021 -24990
rect 22159 -25106 22175 -24966
rect 22020 -25206 22175 -25106
rect 22020 -25310 22021 -25206
rect 21699 -25311 22021 -25310
rect 21814 -25689 21914 -25311
rect 22150 -25338 22175 -25206
rect 22239 -25106 22255 -24966
rect 22878 -24968 22974 -24952
rect 22418 -24990 22740 -24989
rect 22418 -25106 22419 -24990
rect 22239 -25206 22419 -25106
rect 22239 -25338 22255 -25206
rect 22418 -25310 22419 -25206
rect 22739 -25106 22740 -24990
rect 22878 -25106 22894 -24968
rect 22739 -25206 22894 -25106
rect 22739 -25310 22740 -25206
rect 22418 -25311 22740 -25310
rect 22150 -25354 22255 -25338
rect 22878 -25338 22894 -25206
rect 22958 -25106 22974 -24968
rect 23597 -24968 23693 -24952
rect 23137 -24990 23459 -24989
rect 23137 -25106 23138 -24990
rect 22958 -25206 23138 -25106
rect 22958 -25338 22974 -25206
rect 23137 -25310 23138 -25206
rect 23458 -25106 23459 -24990
rect 23597 -25106 23613 -24968
rect 23458 -25206 23613 -25106
rect 23458 -25310 23459 -25206
rect 23137 -25311 23459 -25310
rect 22878 -25354 22974 -25338
rect 23597 -25338 23613 -25206
rect 23677 -25106 23693 -24968
rect 24316 -24968 24412 -24952
rect 23856 -24990 24178 -24989
rect 23856 -25106 23857 -24990
rect 23677 -25206 23857 -25106
rect 23677 -25338 23693 -25206
rect 23856 -25310 23857 -25206
rect 24177 -25106 24178 -24990
rect 24316 -25106 24332 -24968
rect 24177 -25206 24332 -25106
rect 24177 -25310 24178 -25206
rect 23856 -25311 24178 -25310
rect 23597 -25354 23693 -25338
rect 24316 -25338 24332 -25206
rect 24396 -25106 24412 -24968
rect 25035 -24968 25131 -24952
rect 24575 -24990 24897 -24989
rect 24575 -25106 24576 -24990
rect 24396 -25206 24576 -25106
rect 24396 -25338 24418 -25206
rect 24575 -25310 24576 -25206
rect 24896 -25106 24897 -24990
rect 25035 -25106 25051 -24968
rect 24896 -25206 25051 -25106
rect 24896 -25310 24897 -25206
rect 24575 -25311 24897 -25310
rect 22150 -25652 22250 -25354
rect 22528 -25560 24072 -25460
rect 22150 -25668 22255 -25652
rect 21699 -25690 22021 -25689
rect 21699 -26010 21700 -25690
rect 22020 -25796 22021 -25690
rect 22150 -25796 22175 -25668
rect 22020 -25896 22175 -25796
rect 22020 -26010 22021 -25896
rect 22150 -26010 22175 -25896
rect 21699 -26011 22021 -26010
rect 22159 -26036 22175 -26010
rect 22239 -26036 22255 -25668
rect 22528 -25689 22628 -25560
rect 22878 -25668 22974 -25652
rect 22418 -25690 22740 -25689
rect 22418 -26010 22419 -25690
rect 22739 -26010 22740 -25690
rect 22418 -26011 22740 -26010
rect 22159 -26056 22255 -26036
rect 22528 -26152 22628 -26011
rect 22878 -26036 22894 -25668
rect 22958 -26036 22974 -25668
rect 23248 -25689 23348 -25560
rect 23597 -25668 23693 -25652
rect 23137 -25690 23459 -25689
rect 23137 -26010 23138 -25690
rect 23458 -26010 23459 -25690
rect 23137 -26011 23459 -26010
rect 22878 -26056 22974 -26036
rect 23248 -26152 23348 -26011
rect 23597 -26036 23613 -25668
rect 23677 -26036 23693 -25668
rect 23970 -25689 24071 -25560
rect 24316 -25668 24418 -25338
rect 23856 -25690 24178 -25689
rect 23856 -26010 23857 -25690
rect 24177 -26010 24178 -25690
rect 23856 -26011 24178 -26010
rect 23597 -26056 23693 -26036
rect 23970 -26152 24071 -26011
rect 24316 -26036 24332 -25668
rect 24396 -25800 24418 -25668
rect 24690 -25689 24790 -25311
rect 25028 -25338 25051 -25206
rect 25115 -25338 25131 -24968
rect 37159 -24966 37255 -24950
rect 36699 -24990 37021 -24989
rect 36699 -25310 36700 -24990
rect 37020 -25106 37021 -24990
rect 37159 -25106 37175 -24966
rect 37020 -25206 37175 -25106
rect 37020 -25310 37021 -25206
rect 36699 -25311 37021 -25310
rect 25028 -25668 25131 -25338
rect 24575 -25690 24897 -25689
rect 24575 -25800 24576 -25690
rect 24396 -25900 24576 -25800
rect 24396 -26036 24418 -25900
rect 24575 -26010 24576 -25900
rect 24896 -25800 24897 -25690
rect 25028 -25800 25051 -25668
rect 24896 -25900 25051 -25800
rect 24896 -26010 24897 -25900
rect 24575 -26011 24897 -26010
rect 24690 -26012 24790 -26011
rect 24316 -26050 24418 -26036
rect 25028 -26036 25051 -25900
rect 25115 -26036 25131 -25668
rect 36814 -25689 36914 -25311
rect 37150 -25338 37175 -25206
rect 37239 -25106 37255 -24966
rect 37878 -24968 37974 -24952
rect 37418 -24990 37740 -24989
rect 37418 -25106 37419 -24990
rect 37239 -25206 37419 -25106
rect 37239 -25338 37255 -25206
rect 37418 -25310 37419 -25206
rect 37739 -25106 37740 -24990
rect 37878 -25106 37894 -24968
rect 37739 -25206 37894 -25106
rect 37739 -25310 37740 -25206
rect 37418 -25311 37740 -25310
rect 37150 -25354 37255 -25338
rect 37878 -25338 37894 -25206
rect 37958 -25106 37974 -24968
rect 38597 -24968 38693 -24952
rect 38137 -24990 38459 -24989
rect 38137 -25106 38138 -24990
rect 37958 -25206 38138 -25106
rect 37958 -25338 37974 -25206
rect 38137 -25310 38138 -25206
rect 38458 -25106 38459 -24990
rect 38597 -25106 38613 -24968
rect 38458 -25206 38613 -25106
rect 38458 -25310 38459 -25206
rect 38137 -25311 38459 -25310
rect 37878 -25354 37974 -25338
rect 38597 -25338 38613 -25206
rect 38677 -25106 38693 -24968
rect 39316 -24968 39412 -24952
rect 38856 -24990 39178 -24989
rect 38856 -25106 38857 -24990
rect 38677 -25206 38857 -25106
rect 38677 -25338 38693 -25206
rect 38856 -25310 38857 -25206
rect 39177 -25106 39178 -24990
rect 39316 -25106 39332 -24968
rect 39177 -25206 39332 -25106
rect 39177 -25310 39178 -25206
rect 38856 -25311 39178 -25310
rect 38597 -25354 38693 -25338
rect 39316 -25338 39332 -25206
rect 39396 -25106 39412 -24968
rect 40035 -24968 40131 -24952
rect 39575 -24990 39897 -24989
rect 39575 -25106 39576 -24990
rect 39396 -25206 39576 -25106
rect 39396 -25338 39418 -25206
rect 39575 -25310 39576 -25206
rect 39896 -25106 39897 -24990
rect 40035 -25106 40051 -24968
rect 39896 -25206 40051 -25106
rect 39896 -25310 39897 -25206
rect 39575 -25311 39897 -25310
rect 37150 -25652 37250 -25354
rect 37528 -25560 39072 -25460
rect 37150 -25668 37255 -25652
rect 36699 -25690 37021 -25689
rect 36699 -26010 36700 -25690
rect 37020 -25796 37021 -25690
rect 37150 -25796 37175 -25668
rect 37020 -25896 37175 -25796
rect 37020 -26010 37021 -25896
rect 37150 -26010 37175 -25896
rect 36699 -26011 37021 -26010
rect 25028 -26050 25131 -26036
rect 24316 -26056 24412 -26050
rect 25035 -26056 25131 -26050
rect 37159 -26036 37175 -26010
rect 37239 -26036 37255 -25668
rect 37528 -25689 37628 -25560
rect 37878 -25668 37974 -25652
rect 37418 -25690 37740 -25689
rect 37418 -26010 37419 -25690
rect 37739 -26010 37740 -25690
rect 37418 -26011 37740 -26010
rect 37159 -26056 37255 -26036
rect 37528 -26152 37628 -26011
rect 37878 -26036 37894 -25668
rect 37958 -26036 37974 -25668
rect 38248 -25689 38348 -25560
rect 38597 -25668 38693 -25652
rect 38137 -25690 38459 -25689
rect 38137 -26010 38138 -25690
rect 38458 -26010 38459 -25690
rect 38137 -26011 38459 -26010
rect 37878 -26056 37974 -26036
rect 38248 -26152 38348 -26011
rect 38597 -26036 38613 -25668
rect 38677 -26036 38693 -25668
rect 38970 -25689 39071 -25560
rect 39316 -25668 39418 -25338
rect 38856 -25690 39178 -25689
rect 38856 -26010 38857 -25690
rect 39177 -26010 39178 -25690
rect 38856 -26011 39178 -26010
rect 38597 -26056 38693 -26036
rect 38970 -26152 39071 -26011
rect 39316 -26036 39332 -25668
rect 39396 -25800 39418 -25668
rect 39690 -25689 39790 -25311
rect 40028 -25338 40051 -25206
rect 40115 -25338 40131 -24968
rect 40028 -25668 40131 -25338
rect 39575 -25690 39897 -25689
rect 39575 -25800 39576 -25690
rect 39396 -25900 39576 -25800
rect 39396 -26036 39418 -25900
rect 39575 -26010 39576 -25900
rect 39896 -25800 39897 -25690
rect 40028 -25800 40051 -25668
rect 39896 -25900 40051 -25800
rect 39896 -26010 39897 -25900
rect 39575 -26011 39897 -26010
rect 39690 -26012 39790 -26011
rect 39316 -26050 39418 -26036
rect 40028 -26036 40051 -25900
rect 40115 -26036 40131 -25668
rect 40028 -26050 40131 -26036
rect 39316 -26056 39412 -26050
rect 40035 -26056 40131 -26050
rect 21338 -26153 25502 -26152
rect 21338 -26251 21339 -26153
rect 21437 -26251 25403 -26153
rect 25501 -26251 25502 -26153
rect 21338 -26252 25502 -26251
rect 36338 -26153 40400 -26152
rect 36338 -26251 36339 -26153
rect 36437 -26251 40301 -26153
rect 40399 -26251 40400 -26153
rect 36338 -26252 40400 -26251
rect 22159 -26368 22255 -26352
rect 22159 -26388 22175 -26368
rect 21814 -26389 21914 -26388
rect 21699 -26390 22021 -26389
rect 21699 -26710 21700 -26390
rect 22020 -26498 22021 -26390
rect 22150 -26498 22175 -26388
rect 22020 -26598 22175 -26498
rect 22020 -26710 22021 -26598
rect 21699 -26711 22021 -26710
rect 21814 -27089 21914 -26711
rect 22150 -26736 22175 -26598
rect 22239 -26736 22255 -26368
rect 22528 -26389 22628 -26252
rect 22878 -26368 22974 -26352
rect 22418 -26390 22740 -26389
rect 22418 -26710 22419 -26390
rect 22739 -26710 22740 -26390
rect 22418 -26711 22740 -26710
rect 22150 -26754 22255 -26736
rect 22150 -27052 22250 -26754
rect 22528 -26854 22628 -26711
rect 22878 -26736 22894 -26368
rect 22958 -26736 22974 -26368
rect 23248 -26389 23348 -26252
rect 23597 -26368 23693 -26352
rect 23137 -26390 23459 -26389
rect 23137 -26710 23138 -26390
rect 23458 -26710 23459 -26390
rect 23137 -26711 23459 -26710
rect 22878 -26754 22974 -26736
rect 23248 -26854 23348 -26711
rect 23597 -26736 23613 -26368
rect 23677 -26736 23693 -26368
rect 23970 -26389 24071 -26252
rect 24318 -26352 24418 -26350
rect 24316 -26368 24418 -26352
rect 23856 -26390 24178 -26389
rect 23856 -26710 23857 -26390
rect 24177 -26710 24178 -26390
rect 23856 -26711 24178 -26710
rect 23597 -26754 23693 -26736
rect 23970 -26854 24071 -26711
rect 24316 -26736 24332 -26368
rect 24396 -26504 24418 -26368
rect 25028 -26352 25128 -26350
rect 25028 -26368 25131 -26352
rect 24690 -26389 24790 -26388
rect 24575 -26390 24897 -26389
rect 24575 -26504 24576 -26390
rect 24396 -26604 24576 -26504
rect 24396 -26736 24418 -26604
rect 24575 -26710 24576 -26604
rect 24896 -26504 24897 -26390
rect 25028 -26504 25051 -26368
rect 24896 -26604 25051 -26504
rect 24896 -26710 24897 -26604
rect 24575 -26711 24897 -26710
rect 24316 -26754 24418 -26736
rect 22528 -26954 24071 -26854
rect 22150 -27068 22255 -27052
rect 21699 -27090 22021 -27089
rect 21699 -27410 21700 -27090
rect 22020 -27204 22021 -27090
rect 22150 -27204 22175 -27068
rect 22020 -27304 22175 -27204
rect 22020 -27410 22021 -27304
rect 21699 -27411 22021 -27410
rect 21814 -27789 21914 -27411
rect 22150 -27436 22175 -27304
rect 22239 -27436 22255 -27068
rect 22528 -27089 22628 -26954
rect 22878 -27068 22974 -27052
rect 22418 -27090 22740 -27089
rect 22418 -27410 22419 -27090
rect 22739 -27410 22740 -27090
rect 22418 -27411 22740 -27410
rect 22150 -27454 22255 -27436
rect 22150 -27752 22250 -27454
rect 22528 -27554 22628 -27411
rect 22878 -27436 22894 -27068
rect 22958 -27436 22974 -27068
rect 23248 -27089 23348 -26954
rect 23597 -27068 23693 -27052
rect 23137 -27090 23459 -27089
rect 23137 -27410 23138 -27090
rect 23458 -27410 23459 -27090
rect 23137 -27411 23459 -27410
rect 22878 -27454 22974 -27436
rect 23248 -27554 23348 -27411
rect 23597 -27436 23613 -27068
rect 23677 -27436 23693 -27068
rect 23970 -27089 24071 -26954
rect 24318 -27052 24418 -26754
rect 24316 -27068 24418 -27052
rect 23856 -27090 24178 -27089
rect 23856 -27410 23857 -27090
rect 24177 -27410 24178 -27090
rect 23856 -27411 24178 -27410
rect 23597 -27454 23693 -27436
rect 23970 -27554 24071 -27411
rect 24316 -27436 24332 -27068
rect 24396 -27196 24418 -27068
rect 24690 -27089 24790 -26711
rect 25028 -26736 25051 -26604
rect 25115 -26736 25131 -26368
rect 37159 -26368 37255 -26352
rect 37159 -26388 37175 -26368
rect 36814 -26389 36914 -26388
rect 36699 -26390 37021 -26389
rect 36699 -26710 36700 -26390
rect 37020 -26498 37021 -26390
rect 37150 -26498 37175 -26388
rect 37020 -26598 37175 -26498
rect 37020 -26710 37021 -26598
rect 36699 -26711 37021 -26710
rect 25028 -26754 25131 -26736
rect 25028 -27052 25128 -26754
rect 25028 -27068 25131 -27052
rect 24575 -27090 24897 -27089
rect 24575 -27196 24576 -27090
rect 24396 -27296 24576 -27196
rect 24396 -27436 24418 -27296
rect 24575 -27410 24576 -27296
rect 24896 -27196 24897 -27090
rect 25028 -27196 25051 -27068
rect 24896 -27296 25051 -27196
rect 24896 -27410 24897 -27296
rect 24575 -27411 24897 -27410
rect 22528 -27654 24072 -27554
rect 22150 -27768 22255 -27752
rect 21699 -27790 22021 -27789
rect 21699 -27850 21700 -27790
rect 10586 -27902 21700 -27850
rect 10586 -27988 11210 -27902
rect 11306 -27988 11790 -27902
rect 11886 -27988 12390 -27902
rect 12486 -27988 12990 -27902
rect 13086 -27988 13590 -27902
rect 13686 -27988 14190 -27902
rect 14286 -27988 14790 -27902
rect 14886 -27988 15390 -27902
rect 15486 -27988 15990 -27902
rect 16086 -27988 16590 -27902
rect 16686 -27988 17190 -27902
rect 17286 -27988 17790 -27902
rect 17886 -27988 18390 -27902
rect 18486 -27988 18990 -27902
rect 19086 -27988 19590 -27902
rect 19686 -27988 20190 -27902
rect 20286 -27988 20790 -27902
rect 20886 -27988 21700 -27902
rect 10586 -28110 21700 -27988
rect 22020 -27850 22021 -27790
rect 22150 -27850 22175 -27768
rect 22020 -28110 22175 -27850
rect 10586 -28136 22175 -28110
rect 22239 -27850 22255 -27768
rect 22878 -27768 22974 -27752
rect 22418 -27790 22740 -27789
rect 22418 -27850 22419 -27790
rect 22239 -28110 22419 -27850
rect 22739 -27850 22740 -27790
rect 22878 -27850 22894 -27768
rect 22739 -28110 22894 -27850
rect 22239 -28136 22894 -28110
rect 22958 -27850 22974 -27768
rect 23597 -27768 23693 -27752
rect 23137 -27790 23459 -27789
rect 23137 -27850 23138 -27790
rect 22958 -28110 23138 -27850
rect 23458 -27850 23459 -27790
rect 23597 -27850 23613 -27768
rect 23458 -28110 23613 -27850
rect 22958 -28136 23613 -28110
rect 23677 -27850 23693 -27768
rect 24316 -27768 24418 -27436
rect 23856 -27790 24178 -27789
rect 23856 -27850 23857 -27790
rect 23677 -28110 23857 -27850
rect 24177 -27850 24178 -27790
rect 24316 -27850 24332 -27768
rect 24177 -28110 24332 -27850
rect 23677 -28136 24332 -28110
rect 24396 -27850 24418 -27768
rect 24690 -27789 24790 -27411
rect 25028 -27436 25051 -27296
rect 25115 -27436 25131 -27068
rect 36814 -27089 36914 -26711
rect 37150 -26736 37175 -26598
rect 37239 -26736 37255 -26368
rect 37528 -26389 37628 -26252
rect 37878 -26368 37974 -26352
rect 37418 -26390 37740 -26389
rect 37418 -26710 37419 -26390
rect 37739 -26710 37740 -26390
rect 37418 -26711 37740 -26710
rect 37150 -26754 37255 -26736
rect 37150 -27052 37250 -26754
rect 37528 -26854 37628 -26711
rect 37878 -26736 37894 -26368
rect 37958 -26736 37974 -26368
rect 38248 -26389 38348 -26252
rect 38597 -26368 38693 -26352
rect 38137 -26390 38459 -26389
rect 38137 -26710 38138 -26390
rect 38458 -26710 38459 -26390
rect 38137 -26711 38459 -26710
rect 37878 -26754 37974 -26736
rect 38248 -26854 38348 -26711
rect 38597 -26736 38613 -26368
rect 38677 -26736 38693 -26368
rect 38970 -26389 39071 -26252
rect 39318 -26352 39418 -26350
rect 39316 -26368 39418 -26352
rect 38856 -26390 39178 -26389
rect 38856 -26710 38857 -26390
rect 39177 -26710 39178 -26390
rect 38856 -26711 39178 -26710
rect 38597 -26754 38693 -26736
rect 38970 -26854 39071 -26711
rect 39316 -26736 39332 -26368
rect 39396 -26504 39418 -26368
rect 40028 -26352 40128 -26350
rect 40028 -26368 40131 -26352
rect 39690 -26389 39790 -26388
rect 39575 -26390 39897 -26389
rect 39575 -26504 39576 -26390
rect 39396 -26604 39576 -26504
rect 39396 -26736 39418 -26604
rect 39575 -26710 39576 -26604
rect 39896 -26504 39897 -26390
rect 40028 -26504 40051 -26368
rect 39896 -26604 40051 -26504
rect 39896 -26710 39897 -26604
rect 39575 -26711 39897 -26710
rect 39316 -26754 39418 -26736
rect 37528 -26954 39071 -26854
rect 37150 -27068 37255 -27052
rect 36699 -27090 37021 -27089
rect 36699 -27410 36700 -27090
rect 37020 -27204 37021 -27090
rect 37150 -27204 37175 -27068
rect 37020 -27304 37175 -27204
rect 37020 -27410 37021 -27304
rect 36699 -27411 37021 -27410
rect 25028 -27768 25131 -27436
rect 24575 -27790 24897 -27789
rect 24575 -27850 24576 -27790
rect 24396 -28110 24576 -27850
rect 24896 -27850 24897 -27790
rect 25028 -27850 25051 -27768
rect 24896 -28110 25051 -27850
rect 24396 -28136 25051 -28110
rect 25115 -27850 25131 -27768
rect 36814 -27789 36914 -27411
rect 37150 -27436 37175 -27304
rect 37239 -27436 37255 -27068
rect 37528 -27089 37628 -26954
rect 37878 -27068 37974 -27052
rect 37418 -27090 37740 -27089
rect 37418 -27410 37419 -27090
rect 37739 -27410 37740 -27090
rect 37418 -27411 37740 -27410
rect 37150 -27454 37255 -27436
rect 37150 -27752 37250 -27454
rect 37528 -27554 37628 -27411
rect 37878 -27436 37894 -27068
rect 37958 -27436 37974 -27068
rect 38248 -27089 38348 -26954
rect 38597 -27068 38693 -27052
rect 38137 -27090 38459 -27089
rect 38137 -27410 38138 -27090
rect 38458 -27410 38459 -27090
rect 38137 -27411 38459 -27410
rect 37878 -27454 37974 -27436
rect 38248 -27554 38348 -27411
rect 38597 -27436 38613 -27068
rect 38677 -27436 38693 -27068
rect 38970 -27089 39071 -26954
rect 39318 -27052 39418 -26754
rect 39316 -27068 39418 -27052
rect 38856 -27090 39178 -27089
rect 38856 -27410 38857 -27090
rect 39177 -27410 39178 -27090
rect 38856 -27411 39178 -27410
rect 38597 -27454 38693 -27436
rect 38970 -27554 39071 -27411
rect 39316 -27436 39332 -27068
rect 39396 -27196 39418 -27068
rect 39690 -27089 39790 -26711
rect 40028 -26736 40051 -26604
rect 40115 -26736 40131 -26368
rect 40028 -26754 40131 -26736
rect 40028 -27052 40128 -26754
rect 40028 -27068 40131 -27052
rect 39575 -27090 39897 -27089
rect 39575 -27196 39576 -27090
rect 39396 -27296 39576 -27196
rect 39396 -27436 39418 -27296
rect 39575 -27410 39576 -27296
rect 39896 -27196 39897 -27090
rect 40028 -27196 40051 -27068
rect 39896 -27296 40051 -27196
rect 39896 -27410 39897 -27296
rect 39575 -27411 39897 -27410
rect 37528 -27654 39072 -27554
rect 37150 -27768 37255 -27752
rect 36699 -27790 37021 -27789
rect 36699 -27850 36700 -27790
rect 25115 -27902 36700 -27850
rect 25115 -27988 26210 -27902
rect 26306 -27988 26790 -27902
rect 26886 -27988 27390 -27902
rect 27486 -27988 27990 -27902
rect 28086 -27988 28590 -27902
rect 28686 -27988 29190 -27902
rect 29286 -27988 29790 -27902
rect 29886 -27988 30390 -27902
rect 30486 -27988 30990 -27902
rect 31086 -27988 31590 -27902
rect 31686 -27988 32190 -27902
rect 32286 -27988 32790 -27902
rect 32886 -27988 33390 -27902
rect 33486 -27988 33990 -27902
rect 34086 -27988 34590 -27902
rect 34686 -27988 35190 -27902
rect 35286 -27988 35790 -27902
rect 35886 -27988 36700 -27902
rect 25115 -28110 36700 -27988
rect 37020 -27850 37021 -27790
rect 37150 -27850 37175 -27768
rect 37020 -28110 37175 -27850
rect 25115 -28136 37175 -28110
rect 37239 -27850 37255 -27768
rect 37878 -27768 37974 -27752
rect 37418 -27790 37740 -27789
rect 37418 -27850 37419 -27790
rect 37239 -28110 37419 -27850
rect 37739 -27850 37740 -27790
rect 37878 -27850 37894 -27768
rect 37739 -28110 37894 -27850
rect 37239 -28136 37894 -28110
rect 37958 -27850 37974 -27768
rect 38597 -27768 38693 -27752
rect 38137 -27790 38459 -27789
rect 38137 -27850 38138 -27790
rect 37958 -28110 38138 -27850
rect 38458 -27850 38459 -27790
rect 38597 -27850 38613 -27768
rect 38458 -28110 38613 -27850
rect 37958 -28136 38613 -28110
rect 38677 -27850 38693 -27768
rect 39316 -27768 39418 -27436
rect 38856 -27790 39178 -27789
rect 38856 -27850 38857 -27790
rect 38677 -28110 38857 -27850
rect 39177 -27850 39178 -27790
rect 39316 -27850 39332 -27768
rect 39177 -28110 39332 -27850
rect 38677 -28136 39332 -28110
rect 39396 -27850 39418 -27768
rect 39690 -27789 39790 -27411
rect 40028 -27436 40051 -27296
rect 40115 -27436 40131 -27068
rect 40028 -27768 40131 -27436
rect 39575 -27790 39897 -27789
rect 39575 -27850 39576 -27790
rect 39396 -28110 39576 -27850
rect 39896 -27850 39897 -27790
rect 40028 -27850 40051 -27768
rect 39896 -28110 40051 -27850
rect 39396 -28136 40051 -28110
rect 40115 -27850 40131 -27768
rect 40115 -28136 40288 -27850
rect 10586 -28166 40288 -28136
rect 10586 -28466 10924 -28166
rect 11524 -28466 20556 -28166
rect 21156 -28466 25924 -28166
rect 26524 -28466 35556 -28166
rect 36156 -28466 40288 -28166
rect 10586 -28650 40288 -28466
rect 24318 -28654 24418 -28650
rect 39318 -28654 39418 -28650
<< via4 >>
rect 9784 3588 10584 4388
rect 40432 -2722 41178 -974
rect 9814 -11722 10548 -9878
rect 40432 -20726 41166 -18880
rect 9786 -28650 10586 -27850
<< metal5 >>
rect 9786 4412 10586 4472
rect 9760 4388 10608 4412
rect 9760 3588 9784 4388
rect 10584 3588 10608 4388
rect 9760 3564 10608 3588
rect 9786 -9878 10586 3564
rect 9786 -11722 9814 -9878
rect 10548 -11722 10586 -9878
rect 9786 -27826 10586 -11722
rect 40402 -974 41202 4472
rect 40402 -2722 40432 -974
rect 41178 -2722 41202 -974
rect 40402 -18880 41202 -2722
rect 40402 -20726 40432 -18880
rect 41166 -20726 41202 -18880
rect 9762 -27850 10610 -27826
rect 9762 -28650 9786 -27850
rect 10586 -28650 10610 -27850
rect 9762 -28674 10610 -28650
rect 9786 -28686 10586 -28674
rect 40402 -28686 41202 -20726
<< labels >>
flabel metal2 16596 1582 16604 1588 5 FreeSans 480 0 0 0 vpbias
flabel metal1 18498 3414 18504 3422 5 FreeSans 480 0 0 0 vctrl
port 3 s
flabel metal1 32398 2246 32414 2260 1 FreeSans 480 0 0 0 voscbuf
port 4 n
flabel metal1 31098 2304 31114 2316 1 FreeSans 480 0 0 0 vosc
port 5 n
flabel metal1 31796 2256 31804 2260 1 FreeSans 480 0 0 0 vosc2
flabel metal4 13612 3930 13632 3948 1 FreeSans 480 0 0 0 VSS
port 2 n ground bidirectional
flabel metal4 13272 -1542 13284 -1524 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel locali 31706 2167 31740 2201 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 31706 2235 31740 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 31614 2235 31648 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 31571 1929 31605 1963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 31571 2473 31605 2507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 31571 2473 31605 2507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 31571 1929 31605 1963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 31542 2490 31542 2490 2 sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali 32215 2303 32249 2337 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 32215 2235 32249 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 32215 2167 32249 2201 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 31847 2235 31881 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 31939 2235 31973 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 32031 2235 32065 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 32123 2235 32157 2269 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel nwell 31847 1929 31881 1963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VPB
flabel pwell 31847 2473 31881 2507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VNB
flabel metal1 31847 1929 31881 1963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VPWR
flabel metal1 31847 2473 31881 2507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VGND
rlabel comment 31818 2490 31818 2490 2 sky130_fd_sc_hd__inv_4_0/inv_4
flabel metal4 28540 -10248 28560 -10228 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/VSS
flabel metal4 28306 -2344 28340 -2320 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/VDD
flabel metal2 27140 -7994 27154 -7980 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/vin
flabel metal1 27142 -9688 27150 -9678 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/vbiasn
flabel metal2 27612 -5272 27622 -5266 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/vbiasp
flabel metal2 34966 -8000 34978 -7986 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/voutcs
flabel metal2 35372 -7970 35384 -7960 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/vout
flabel metal1 26706 -9098 26718 -9080 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/csinvn
flabel metal2 27256 -5870 27266 -5856 1 FreeSans 480 0 0 0 cs_ring_osc_stage_5/csinvp
flabel metal4 13540 -10248 13560 -10228 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/VSS
flabel metal4 13306 -2344 13340 -2320 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/VDD
flabel metal2 12140 -7994 12154 -7980 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/vin
flabel metal1 12142 -9688 12150 -9678 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/vbiasn
flabel metal2 12612 -5272 12622 -5266 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/vbiasp
flabel metal2 19966 -8000 19978 -7986 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/voutcs
flabel metal2 20372 -7970 20384 -7960 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/vout
flabel metal1 11706 -9098 11718 -9080 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/csinvn
flabel metal2 12256 -5870 12266 -5856 1 FreeSans 480 0 0 0 cs_ring_osc_stage_0/csinvp
flabel metal4 37474 -11376 37494 -11356 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/VSS
flabel metal4 37694 -19284 37728 -19260 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/VDD
flabel metal2 38880 -13624 38894 -13610 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/vin
flabel metal1 38884 -11926 38892 -11916 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/vbiasn
flabel metal2 38412 -16338 38422 -16332 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/vbiasp
flabel metal2 31056 -13618 31068 -13604 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/voutcs
flabel metal2 30650 -13644 30662 -13634 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/vout
flabel metal1 39316 -12524 39328 -12506 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/csinvn
flabel metal2 38768 -15748 38778 -15734 5 FreeSans 480 0 0 0 cs_ring_osc_stage_4/csinvp
flabel metal4 22474 -11376 22494 -11356 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/VSS
flabel metal4 22694 -19284 22728 -19260 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/VDD
flabel metal2 23880 -13624 23894 -13610 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/vin
flabel metal1 23884 -11926 23892 -11916 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/vbiasn
flabel metal2 23412 -16338 23422 -16332 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/vbiasp
flabel metal2 16056 -13618 16068 -13604 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/voutcs
flabel metal2 15650 -13644 15662 -13634 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/vout
flabel metal1 24316 -12524 24328 -12506 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/csinvn
flabel metal2 23768 -15748 23778 -15734 5 FreeSans 480 0 0 0 cs_ring_osc_stage_1/csinvp
flabel metal4 28540 -28248 28560 -28228 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/VSS
flabel metal4 28306 -20344 28340 -20320 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/VDD
flabel metal2 27140 -25994 27154 -25980 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/vin
flabel metal1 27142 -27688 27150 -27678 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/vbiasn
flabel metal2 27612 -23272 27622 -23266 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/vbiasp
flabel metal2 34966 -26000 34978 -25986 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/voutcs
flabel metal2 35372 -25970 35384 -25960 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/vout
flabel metal1 26706 -27098 26718 -27080 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/csinvn
flabel metal2 27256 -23870 27266 -23856 1 FreeSans 480 0 0 0 cs_ring_osc_stage_3/csinvp
flabel metal4 13540 -28248 13560 -28228 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/VSS
flabel metal4 13306 -20344 13340 -20320 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/VDD
flabel metal2 12140 -25994 12154 -25980 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/vin
flabel metal1 12142 -27688 12150 -27678 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/vbiasn
flabel metal2 12612 -23272 12622 -23266 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/vbiasp
flabel metal2 19966 -26000 19978 -25986 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/voutcs
flabel metal2 20372 -25970 20384 -25960 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/vout
flabel metal1 11706 -27098 11718 -27080 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/csinvn
flabel metal2 12256 -23870 12266 -23856 1 FreeSans 480 0 0 0 cs_ring_osc_stage_2/csinvp
<< end >>
