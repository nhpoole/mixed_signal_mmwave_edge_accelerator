magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1298 -1308 1758 1852
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 439 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 247 177
rect 193 127 203 161
rect 237 127 247 161
rect 193 93 247 127
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 47 331 131
rect 361 93 413 177
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 417 413 451
rect 361 383 371 417
rect 405 383 413 417
rect 361 297 413 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 203 127 237 161
rect 203 59 237 93
rect 287 131 321 165
rect 371 59 405 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 79 265 109 297
rect 163 265 193 297
rect 79 249 193 265
rect 79 215 119 249
rect 153 215 193 249
rect 79 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 265 277 297
rect 331 265 361 297
rect 247 249 361 265
rect 247 215 287 249
rect 321 215 361 249
rect 247 199 361 215
rect 247 177 277 199
rect 331 177 361 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
<< polycont >>
rect 119 215 153 249
rect 287 215 321 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 422 527
rect 405 451 422 485
rect 371 417 422 451
rect 405 383 422 417
rect 371 367 422 383
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 321 315 443 333
rect 103 299 443 315
rect 17 249 169 265
rect 17 215 119 249
rect 153 215 169 249
rect 203 249 353 265
rect 203 215 287 249
rect 321 215 353 249
rect 387 181 443 299
rect 17 161 237 177
rect 17 127 35 161
rect 69 143 203 161
rect 69 127 85 143
rect 17 93 85 127
rect 187 127 203 143
rect 271 165 443 181
rect 271 131 287 165
rect 321 131 443 165
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 119 93 153 109
rect 119 17 153 59
rect 187 93 237 127
rect 355 93 421 97
rect 187 59 203 93
rect 237 59 371 93
rect 405 59 421 93
rect 187 51 421 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 398 153 432 187 0 FreeSans 250 0 0 0 Y
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 Y
flabel locali s 398 289 432 323 0 FreeSans 250 0 0 0 Y
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 A
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
rlabel comment s 0 0 0 0 4 nand2_2
<< properties >>
string FIXED_BBOX 0 0 460 544
string path 0.000 0.000 11.500 0.000 
<< end >>
