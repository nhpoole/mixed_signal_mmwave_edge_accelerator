magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -36 679 1160 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 1124 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 918 1130 952 1397
rect 1022 1322 1056 1397
rect 64 674 98 740
rect 490 724 524 1096
rect 490 690 541 724
rect 490 318 524 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 918 17 952 218
rect 1022 17 1056 92
rect 0 -17 1124 17
use nmos_m8_w2_000_sli_dli_da_p  nmos_m8_w2_000_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 51
box -26 -26 932 456
use pmos_m8_w2_000_sli_dli_da_p  pmos_m8_w2_000_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 963
box -59 -56 965 454
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 48 0 1 674
box 0 0 66 66
use contact_28  contact_28_0
timestamp 1624494425
transform 1 0 1014 0 1 51
box -26 -26 76 108
use contact_27  contact_27_0
timestamp 1624494425
transform 1 0 1014 0 1 1281
box -59 -43 109 125
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 524 707 524 707 4 Z
rlabel locali s 562 0 562 0 4 gnd
rlabel locali s 562 1414 562 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1124 1414
<< end >>
