magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1296 -1277 1880 2731
<< nwell >>
rect -36 679 620 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 584 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 482 1322 516 1397
rect 64 674 98 740
rect 272 724 306 1096
rect 272 690 323 724
rect 272 318 306 690
rect 62 17 96 218
rect 274 17 308 218
rect 482 17 516 92
rect 0 -17 584 17
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m3_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m3_w2_000_sli_dli_da_p_0
timestamp 1626065694
transform 1 0 54 0 1 963
box -59 -56 425 454
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m3_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m3_w2_000_sli_dli_da_p_0
timestamp 1626065694
transform 1 0 54 0 1 51
box -26 -26 392 456
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1626065694
transform 1 0 48 0 1 674
box 0 0 66 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1626065694
transform 1 0 474 0 1 51
box -26 -26 76 108
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1626065694
transform 1 0 474 0 1 1281
box -59 -43 109 125
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 306 707 306 707 4 Z
rlabel locali s 292 0 292 0 4 gnd
rlabel locali s 292 1414 292 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 584 1414
<< end >>
