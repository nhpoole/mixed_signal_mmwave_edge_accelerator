magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 1935 517 1969 551
rect 21903 517 21937 551
rect 41871 517 41905 551
rect 61839 517 61873 551
rect 1374 253 1503 287
rect 21342 253 21471 287
rect 41310 253 41439 287
rect 61278 253 61407 287
<< metal1 >>
rect -32 1134 32 1146
rect 81214 1134 81278 1146
rect -32 1106 81278 1134
rect -32 1094 32 1106
rect 81214 1094 81278 1106
rect 1571 492 1635 544
rect 21539 492 21603 544
rect 41507 492 41571 544
rect 61475 492 61539 544
rect 1342 244 1406 296
rect 21310 244 21374 296
rect 41278 244 41342 296
rect 61246 244 61310 296
rect -32 14 32 26
rect 81214 14 81278 26
rect -32 -14 81278 14
rect -32 -26 32 -14
rect 81214 -26 81278 -14
<< metal2 >>
rect -28 1096 28 1144
rect 81218 1096 81274 1144
rect 1575 494 1631 542
rect 21543 494 21599 542
rect 41511 494 41567 542
rect 61479 494 61535 542
rect 1360 256 1388 284
rect 21328 256 21356 284
rect 41296 256 41324 284
rect 61264 256 61292 284
rect -28 -24 28 24
rect 81218 -24 81274 24
<< metal3 >>
rect -49 1071 49 1169
rect 81197 1071 81295 1169
rect 0 488 81246 548
rect -49 -49 49 49
rect 81197 -49 81295 49
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 -33 0 1 -37
box 0 0 66 74
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 -32 0 1 -32
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 -29 0 1 -33
box 0 0 58 66
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 -29 0 1 -33
box 0 0 58 66
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 1570 0 1 481
box 0 0 66 74
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 1571 0 1 486
box 0 0 64 64
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 1574 0 1 485
box 0 0 58 66
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 1342 0 1 238
box 0 0 64 64
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 1345 0 1 237
box 0 0 58 66
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 -33 0 1 1083
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 -32 0 1 1088
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 -29 0 1 1087
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 -29 0 1 1087
box 0 0 58 66
use pand2  pand2_3
timestamp 1624494425
transform 1 0 1374 0 1 0
box -36 -17 890 1177
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 1772 0 1 -33
box 0 0 58 66
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 1772 0 1 1087
box 0 0 58 66
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 21313 0 1 237
box 0 0 58 66
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 21310 0 1 238
box 0 0 64 64
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 21542 0 1 485
box 0 0 58 66
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 21539 0 1 486
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 21538 0 1 481
box 0 0 66 74
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 21740 0 1 -33
box 0 0 58 66
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 21740 0 1 1087
box 0 0 58 66
use pand2  pand2_2
timestamp 1624494425
transform 1 0 21342 0 1 0
box -36 -17 890 1177
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 41281 0 1 237
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 41278 0 1 238
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 41510 0 1 485
box 0 0 58 66
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 41507 0 1 486
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 41506 0 1 481
box 0 0 66 74
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 41708 0 1 -33
box 0 0 58 66
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 41708 0 1 1087
box 0 0 58 66
use pand2  pand2_1
timestamp 1624494425
transform 1 0 41310 0 1 0
box -36 -17 890 1177
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 61249 0 1 237
box 0 0 58 66
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 61246 0 1 238
box 0 0 64 64
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 61478 0 1 485
box 0 0 58 66
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 61475 0 1 486
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 61474 0 1 481
box 0 0 66 74
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 61676 0 1 -33
box 0 0 58 66
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 61676 0 1 1087
box 0 0 58 66
use pand2  pand2_0
timestamp 1624494425
transform 1 0 61278 0 1 0
box -36 -17 890 1177
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 81217 0 1 -33
box 0 0 58 66
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 81217 0 1 -33
box 0 0 58 66
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 81214 0 1 -32
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 81213 0 1 -37
box 0 0 66 74
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 81217 0 1 1087
box 0 0 58 66
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 81217 0 1 1087
box 0 0 58 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 81214 0 1 1088
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 81213 0 1 1083
box 0 0 66 74
<< labels >>
rlabel metal3 s 0 488 81246 548 4 en
rlabel metal2 s 1360 256 1388 284 4 wmask_in_0
rlabel locali s 1952 534 1952 534 4 wmask_out_0
rlabel metal2 s 21328 256 21356 284 4 wmask_in_1
rlabel locali s 21920 534 21920 534 4 wmask_out_1
rlabel metal2 s 41296 256 41324 284 4 wmask_in_2
rlabel locali s 41888 534 41888 534 4 wmask_out_2
rlabel metal2 s 61264 256 61292 284 4 wmask_in_3
rlabel locali s 61856 534 61856 534 4 wmask_out_3
rlabel metal3 s 81197 -49 81295 49 4 gnd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal3 s -49 1071 49 1169 4 vdd
rlabel metal3 s 81197 1071 81295 1169 4 vdd
<< properties >>
string FIXED_BBOX 0 0 81246 1120
<< end >>
