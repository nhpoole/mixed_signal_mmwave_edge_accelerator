magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -54 -54 312 454
<< scpmos >>
rect 60 0 90 400
rect 168 0 198 400
<< pdiff >>
rect 0 0 60 400
rect 90 0 168 400
rect 198 0 258 400
<< poly >>
rect 60 400 90 426
rect 168 400 198 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 60 -56 198 -26
<< locali >>
rect 8 167 42 233
rect 112 167 146 233
rect 216 167 250 233
use contact_12  contact_12_2
timestamp 1624494425
transform 1 0 0 0 1 167
box -59 -51 109 117
use contact_12  contact_12_1
timestamp 1624494425
transform 1 0 104 0 1 167
box -59 -51 109 117
use contact_12  contact_12_0
timestamp 1624494425
transform 1 0 208 0 1 167
box -59 -51 109 117
<< labels >>
rlabel poly s 129 -41 129 -41 4 G
rlabel locali s 25 200 25 200 4 S
rlabel locali s 233 200 233 200 4 S
rlabel locali s 129 200 129 200 4 D
<< properties >>
string FIXED_BBOX -54 -56 312 454
<< end >>
