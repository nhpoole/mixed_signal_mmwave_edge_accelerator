magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1403 -200 -1345 200
rect -945 -200 -887 200
rect -487 -200 -429 200
rect -29 -200 29 200
rect 429 -200 487 200
rect 887 -200 945 200
rect 1345 -200 1403 200
<< nmos >>
rect -1345 -200 -945 200
rect -887 -200 -487 200
rect -429 -200 -29 200
rect 29 -200 429 200
rect 487 -200 887 200
rect 945 -200 1345 200
<< ndiff >>
rect -1403 188 -1345 200
rect -1403 -188 -1391 188
rect -1357 -188 -1345 188
rect -1403 -200 -1345 -188
rect -945 188 -887 200
rect -945 -188 -933 188
rect -899 -188 -887 188
rect -945 -200 -887 -188
rect -487 188 -429 200
rect -487 -188 -475 188
rect -441 -188 -429 188
rect -487 -200 -429 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 429 188 487 200
rect 429 -188 441 188
rect 475 -188 487 188
rect 429 -200 487 -188
rect 887 188 945 200
rect 887 -188 899 188
rect 933 -188 945 188
rect 887 -200 945 -188
rect 1345 188 1403 200
rect 1345 -188 1357 188
rect 1391 -188 1403 188
rect 1345 -200 1403 -188
<< ndiffc >>
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
<< poly >>
rect -1271 272 -1019 288
rect -1271 255 -1255 272
rect -1345 238 -1255 255
rect -1035 255 -1019 272
rect -813 272 -561 288
rect -813 255 -797 272
rect -1035 238 -945 255
rect -1345 200 -945 238
rect -887 238 -797 255
rect -577 255 -561 272
rect -355 272 -103 288
rect -355 255 -339 272
rect -577 238 -487 255
rect -887 200 -487 238
rect -429 238 -339 255
rect -119 255 -103 272
rect 103 272 355 288
rect 103 255 119 272
rect -119 238 -29 255
rect -429 200 -29 238
rect 29 238 119 255
rect 339 255 355 272
rect 561 272 813 288
rect 561 255 577 272
rect 339 238 429 255
rect 29 200 429 238
rect 487 238 577 255
rect 797 255 813 272
rect 1019 272 1271 288
rect 1019 255 1035 272
rect 797 238 887 255
rect 487 200 887 238
rect 945 238 1035 255
rect 1255 255 1271 272
rect 1255 238 1345 255
rect 945 200 1345 238
rect -1345 -238 -945 -200
rect -1345 -255 -1255 -238
rect -1271 -272 -1255 -255
rect -1035 -255 -945 -238
rect -887 -238 -487 -200
rect -887 -255 -797 -238
rect -1035 -272 -1019 -255
rect -1271 -288 -1019 -272
rect -813 -272 -797 -255
rect -577 -255 -487 -238
rect -429 -238 -29 -200
rect -429 -255 -339 -238
rect -577 -272 -561 -255
rect -813 -288 -561 -272
rect -355 -272 -339 -255
rect -119 -255 -29 -238
rect 29 -238 429 -200
rect 29 -255 119 -238
rect -119 -272 -103 -255
rect -355 -288 -103 -272
rect 103 -272 119 -255
rect 339 -255 429 -238
rect 487 -238 887 -200
rect 487 -255 577 -238
rect 339 -272 355 -255
rect 103 -288 355 -272
rect 561 -272 577 -255
rect 797 -255 887 -238
rect 945 -238 1345 -200
rect 945 -255 1035 -238
rect 797 -272 813 -255
rect 561 -288 813 -272
rect 1019 -272 1035 -255
rect 1255 -255 1345 -238
rect 1255 -272 1271 -255
rect 1019 -288 1271 -272
<< polycont >>
rect -1255 238 -1035 272
rect -797 238 -577 272
rect -339 238 -119 272
rect 119 238 339 272
rect 577 238 797 272
rect 1035 238 1255 272
rect -1255 -272 -1035 -238
rect -797 -272 -577 -238
rect -339 -272 -119 -238
rect 119 -272 339 -238
rect 577 -272 797 -238
rect 1035 -272 1255 -238
<< locali >>
rect -1271 238 -1255 272
rect -1035 238 -1019 272
rect -813 238 -797 272
rect -577 238 -561 272
rect -355 238 -339 272
rect -119 238 -103 272
rect 103 238 119 272
rect 339 238 355 272
rect 561 238 577 272
rect 797 238 813 272
rect 1019 238 1035 272
rect 1255 238 1271 272
rect -1391 188 -1357 204
rect -1391 -204 -1357 -188
rect -933 188 -899 204
rect -933 -204 -899 -188
rect -475 188 -441 204
rect -475 -204 -441 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 441 188 475 204
rect 441 -204 475 -188
rect 899 188 933 204
rect 899 -204 933 -188
rect 1357 188 1391 204
rect 1357 -204 1391 -188
rect -1271 -272 -1255 -238
rect -1035 -272 -1019 -238
rect -813 -272 -797 -238
rect -577 -272 -561 -238
rect -355 -272 -339 -238
rect -119 -272 -103 -238
rect 103 -272 119 -238
rect 339 -272 355 -238
rect 561 -272 577 -238
rect 797 -272 813 -238
rect 1019 -272 1035 -238
rect 1255 -272 1271 -238
<< viali >>
rect -1237 238 -1053 272
rect -779 238 -595 272
rect -321 238 -137 272
rect 137 238 321 272
rect 595 238 779 272
rect 1053 238 1237 272
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect -1237 -272 -1053 -238
rect -779 -272 -595 -238
rect -321 -272 -137 -238
rect 137 -272 321 -238
rect 595 -272 779 -238
rect 1053 -272 1237 -238
<< metal1 >>
rect -1249 272 -1041 278
rect -1249 238 -1237 272
rect -1053 238 -1041 272
rect -1249 232 -1041 238
rect -791 272 -583 278
rect -791 238 -779 272
rect -595 238 -583 272
rect -791 232 -583 238
rect -333 272 -125 278
rect -333 238 -321 272
rect -137 238 -125 272
rect -333 232 -125 238
rect 125 272 333 278
rect 125 238 137 272
rect 321 238 333 272
rect 125 232 333 238
rect 583 272 791 278
rect 583 238 595 272
rect 779 238 791 272
rect 583 232 791 238
rect 1041 272 1249 278
rect 1041 238 1053 272
rect 1237 238 1249 272
rect 1041 232 1249 238
rect -1397 188 -1351 200
rect -1397 -188 -1391 188
rect -1357 -188 -1351 188
rect -1397 -200 -1351 -188
rect -939 188 -893 200
rect -939 -188 -933 188
rect -899 -188 -893 188
rect -939 -200 -893 -188
rect -481 188 -435 200
rect -481 -188 -475 188
rect -441 -188 -435 188
rect -481 -200 -435 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 435 188 481 200
rect 435 -188 441 188
rect 475 -188 481 188
rect 435 -200 481 -188
rect 893 188 939 200
rect 893 -188 899 188
rect 933 -188 939 188
rect 893 -200 939 -188
rect 1351 188 1397 200
rect 1351 -188 1357 188
rect 1391 -188 1397 188
rect 1351 -200 1397 -188
rect -1249 -238 -1041 -232
rect -1249 -272 -1237 -238
rect -1053 -272 -1041 -238
rect -1249 -278 -1041 -272
rect -791 -238 -583 -232
rect -791 -272 -779 -238
rect -595 -272 -583 -238
rect -791 -278 -583 -272
rect -333 -238 -125 -232
rect -333 -272 -321 -238
rect -137 -272 -125 -238
rect -333 -278 -125 -272
rect 125 -238 333 -232
rect 125 -272 137 -238
rect 321 -272 333 -238
rect 125 -278 333 -272
rect 583 -238 791 -232
rect 583 -272 595 -238
rect 779 -272 791 -238
rect 583 -278 791 -272
rect 1041 -238 1249 -232
rect 1041 -272 1053 -238
rect 1237 -272 1249 -238
rect 1041 -278 1249 -272
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 2 l 2 m 1 nf 6 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
