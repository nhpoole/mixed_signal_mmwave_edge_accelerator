magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -599 -572 728 755
<< pwell >>
rect 31 58 98 125
<< psubdiff >>
rect 44 100 85 112
rect 44 83 56 100
rect 73 83 85 100
rect 44 71 85 83
<< psubdiffcont >>
rect 56 83 73 100
<< locali >>
rect 44 100 85 112
rect 44 83 56 100
rect 73 83 85 100
rect 44 71 85 83
<< end >>
