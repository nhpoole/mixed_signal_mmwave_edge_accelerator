magic
tech sky130A
magscale 1 2
timestamp 1621056506
<< metal3 >>
rect -350 1072 349 1100
rect -350 -1072 265 1072
rect 329 -1072 349 1072
rect -350 -1100 349 -1072
<< via3 >>
rect 265 -1072 329 1072
<< mimcap >>
rect -250 960 150 1000
rect -250 -960 -210 960
rect 110 -960 150 960
rect -250 -1000 150 -960
<< mimcapcontact >>
rect -210 -960 110 960
<< metal4 >>
rect 249 1072 345 1088
rect -211 960 111 961
rect -211 -960 -210 960
rect 110 -960 111 960
rect -211 -961 111 -960
rect 249 -1072 265 1072
rect 329 -1072 345 1072
rect 249 -1088 345 -1072
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -350 -1100 250 1100
string parameters w 2.00 l 10.00 val 44.56 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
