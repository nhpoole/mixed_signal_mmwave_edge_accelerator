magic
tech sky130A
magscale 1 2
timestamp 1621053618
<< error_p >>
rect -2389 2350 -2329 4550
rect -2309 2350 -2249 4550
rect -70 2350 -10 4550
rect 10 2350 70 4550
rect 2249 2350 2309 4550
rect 2329 2350 2389 4550
rect -2389 50 -2329 2250
rect -2309 50 -2249 2250
rect -70 50 -10 2250
rect 10 50 70 2250
rect 2249 50 2309 2250
rect 2329 50 2389 2250
rect -2389 -2250 -2329 -50
rect -2309 -2250 -2249 -50
rect -70 -2250 -10 -50
rect 10 -2250 70 -50
rect 2249 -2250 2309 -50
rect 2329 -2250 2389 -50
rect -2389 -4550 -2329 -2350
rect -2309 -4550 -2249 -2350
rect -70 -4550 -10 -2350
rect 10 -4550 70 -2350
rect 2249 -4550 2309 -2350
rect 2329 -4550 2389 -2350
<< metal3 >>
rect -4628 4522 -2329 4550
rect -4628 2378 -2413 4522
rect -2349 2378 -2329 4522
rect -4628 2350 -2329 2378
rect -2309 4522 -10 4550
rect -2309 2378 -94 4522
rect -30 2378 -10 4522
rect -2309 2350 -10 2378
rect 10 4522 2309 4550
rect 10 2378 2225 4522
rect 2289 2378 2309 4522
rect 10 2350 2309 2378
rect 2329 4522 4628 4550
rect 2329 2378 4544 4522
rect 4608 2378 4628 4522
rect 2329 2350 4628 2378
rect -4628 2222 -2329 2250
rect -4628 78 -2413 2222
rect -2349 78 -2329 2222
rect -4628 50 -2329 78
rect -2309 2222 -10 2250
rect -2309 78 -94 2222
rect -30 78 -10 2222
rect -2309 50 -10 78
rect 10 2222 2309 2250
rect 10 78 2225 2222
rect 2289 78 2309 2222
rect 10 50 2309 78
rect 2329 2222 4628 2250
rect 2329 78 4544 2222
rect 4608 78 4628 2222
rect 2329 50 4628 78
rect -4628 -78 -2329 -50
rect -4628 -2222 -2413 -78
rect -2349 -2222 -2329 -78
rect -4628 -2250 -2329 -2222
rect -2309 -78 -10 -50
rect -2309 -2222 -94 -78
rect -30 -2222 -10 -78
rect -2309 -2250 -10 -2222
rect 10 -78 2309 -50
rect 10 -2222 2225 -78
rect 2289 -2222 2309 -78
rect 10 -2250 2309 -2222
rect 2329 -78 4628 -50
rect 2329 -2222 4544 -78
rect 4608 -2222 4628 -78
rect 2329 -2250 4628 -2222
rect -4628 -2378 -2329 -2350
rect -4628 -4522 -2413 -2378
rect -2349 -4522 -2329 -2378
rect -4628 -4550 -2329 -4522
rect -2309 -2378 -10 -2350
rect -2309 -4522 -94 -2378
rect -30 -4522 -10 -2378
rect -2309 -4550 -10 -4522
rect 10 -2378 2309 -2350
rect 10 -4522 2225 -2378
rect 2289 -4522 2309 -2378
rect 10 -4550 2309 -4522
rect 2329 -2378 4628 -2350
rect 2329 -4522 4544 -2378
rect 4608 -4522 4628 -2378
rect 2329 -4550 4628 -4522
<< via3 >>
rect -2413 2378 -2349 4522
rect -94 2378 -30 4522
rect 2225 2378 2289 4522
rect 4544 2378 4608 4522
rect -2413 78 -2349 2222
rect -94 78 -30 2222
rect 2225 78 2289 2222
rect 4544 78 4608 2222
rect -2413 -2222 -2349 -78
rect -94 -2222 -30 -78
rect 2225 -2222 2289 -78
rect 4544 -2222 4608 -78
rect -2413 -4522 -2349 -2378
rect -94 -4522 -30 -2378
rect 2225 -4522 2289 -2378
rect 4544 -4522 4608 -2378
<< mimcap >>
rect -4528 4410 -2528 4450
rect -4528 2490 -4488 4410
rect -2568 2490 -2528 4410
rect -4528 2450 -2528 2490
rect -2209 4410 -209 4450
rect -2209 2490 -2169 4410
rect -249 2490 -209 4410
rect -2209 2450 -209 2490
rect 110 4410 2110 4450
rect 110 2490 150 4410
rect 2070 2490 2110 4410
rect 110 2450 2110 2490
rect 2429 4410 4429 4450
rect 2429 2490 2469 4410
rect 4389 2490 4429 4410
rect 2429 2450 4429 2490
rect -4528 2110 -2528 2150
rect -4528 190 -4488 2110
rect -2568 190 -2528 2110
rect -4528 150 -2528 190
rect -2209 2110 -209 2150
rect -2209 190 -2169 2110
rect -249 190 -209 2110
rect -2209 150 -209 190
rect 110 2110 2110 2150
rect 110 190 150 2110
rect 2070 190 2110 2110
rect 110 150 2110 190
rect 2429 2110 4429 2150
rect 2429 190 2469 2110
rect 4389 190 4429 2110
rect 2429 150 4429 190
rect -4528 -190 -2528 -150
rect -4528 -2110 -4488 -190
rect -2568 -2110 -2528 -190
rect -4528 -2150 -2528 -2110
rect -2209 -190 -209 -150
rect -2209 -2110 -2169 -190
rect -249 -2110 -209 -190
rect -2209 -2150 -209 -2110
rect 110 -190 2110 -150
rect 110 -2110 150 -190
rect 2070 -2110 2110 -190
rect 110 -2150 2110 -2110
rect 2429 -190 4429 -150
rect 2429 -2110 2469 -190
rect 4389 -2110 4429 -190
rect 2429 -2150 4429 -2110
rect -4528 -2490 -2528 -2450
rect -4528 -4410 -4488 -2490
rect -2568 -4410 -2528 -2490
rect -4528 -4450 -2528 -4410
rect -2209 -2490 -209 -2450
rect -2209 -4410 -2169 -2490
rect -249 -4410 -209 -2490
rect -2209 -4450 -209 -4410
rect 110 -2490 2110 -2450
rect 110 -4410 150 -2490
rect 2070 -4410 2110 -2490
rect 110 -4450 2110 -4410
rect 2429 -2490 4429 -2450
rect 2429 -4410 2469 -2490
rect 4389 -4410 4429 -2490
rect 2429 -4450 4429 -4410
<< mimcapcontact >>
rect -4488 2490 -2568 4410
rect -2169 2490 -249 4410
rect 150 2490 2070 4410
rect 2469 2490 4389 4410
rect -4488 190 -2568 2110
rect -2169 190 -249 2110
rect 150 190 2070 2110
rect 2469 190 4389 2110
rect -4488 -2110 -2568 -190
rect -2169 -2110 -249 -190
rect 150 -2110 2070 -190
rect 2469 -2110 4389 -190
rect -4488 -4410 -2568 -2490
rect -2169 -4410 -249 -2490
rect 150 -4410 2070 -2490
rect 2469 -4410 4389 -2490
<< metal4 >>
rect -3580 4411 -3476 4600
rect -2460 4538 -2356 4600
rect -2460 4522 -2333 4538
rect -4489 4410 -2567 4411
rect -4489 2490 -4488 4410
rect -2568 2490 -2567 4410
rect -4489 2489 -2567 2490
rect -3580 2111 -3476 2489
rect -2460 2378 -2413 4522
rect -2349 2378 -2333 4522
rect -1261 4411 -1157 4600
rect -141 4538 -37 4600
rect -141 4522 -14 4538
rect -2170 4410 -248 4411
rect -2170 2490 -2169 4410
rect -249 2490 -248 4410
rect -2170 2489 -248 2490
rect -2460 2362 -2333 2378
rect -2460 2238 -2356 2362
rect -2460 2222 -2333 2238
rect -4489 2110 -2567 2111
rect -4489 190 -4488 2110
rect -2568 190 -2567 2110
rect -4489 189 -2567 190
rect -3580 -189 -3476 189
rect -2460 78 -2413 2222
rect -2349 78 -2333 2222
rect -1261 2111 -1157 2489
rect -141 2378 -94 4522
rect -30 2378 -14 4522
rect 1058 4411 1162 4600
rect 2178 4538 2282 4600
rect 2178 4522 2305 4538
rect 149 4410 2071 4411
rect 149 2490 150 4410
rect 2070 2490 2071 4410
rect 149 2489 2071 2490
rect -141 2362 -14 2378
rect -141 2238 -37 2362
rect -141 2222 -14 2238
rect -2170 2110 -248 2111
rect -2170 190 -2169 2110
rect -249 190 -248 2110
rect -2170 189 -248 190
rect -2460 62 -2333 78
rect -2460 -62 -2356 62
rect -2460 -78 -2333 -62
rect -4489 -190 -2567 -189
rect -4489 -2110 -4488 -190
rect -2568 -2110 -2567 -190
rect -4489 -2111 -2567 -2110
rect -3580 -2489 -3476 -2111
rect -2460 -2222 -2413 -78
rect -2349 -2222 -2333 -78
rect -1261 -189 -1157 189
rect -141 78 -94 2222
rect -30 78 -14 2222
rect 1058 2111 1162 2489
rect 2178 2378 2225 4522
rect 2289 2378 2305 4522
rect 3377 4411 3481 4600
rect 4497 4538 4601 4600
rect 4497 4522 4624 4538
rect 2468 4410 4390 4411
rect 2468 2490 2469 4410
rect 4389 2490 4390 4410
rect 2468 2489 4390 2490
rect 2178 2362 2305 2378
rect 2178 2238 2282 2362
rect 2178 2222 2305 2238
rect 149 2110 2071 2111
rect 149 190 150 2110
rect 2070 190 2071 2110
rect 149 189 2071 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -2170 -190 -248 -189
rect -2170 -2110 -2169 -190
rect -249 -2110 -248 -190
rect -2170 -2111 -248 -2110
rect -2460 -2238 -2333 -2222
rect -2460 -2362 -2356 -2238
rect -2460 -2378 -2333 -2362
rect -4489 -2490 -2567 -2489
rect -4489 -4410 -4488 -2490
rect -2568 -4410 -2567 -2490
rect -4489 -4411 -2567 -4410
rect -3580 -4600 -3476 -4411
rect -2460 -4522 -2413 -2378
rect -2349 -4522 -2333 -2378
rect -1261 -2489 -1157 -2111
rect -141 -2222 -94 -78
rect -30 -2222 -14 -78
rect 1058 -189 1162 189
rect 2178 78 2225 2222
rect 2289 78 2305 2222
rect 3377 2111 3481 2489
rect 4497 2378 4544 4522
rect 4608 2378 4624 4522
rect 4497 2362 4624 2378
rect 4497 2238 4601 2362
rect 4497 2222 4624 2238
rect 2468 2110 4390 2111
rect 2468 190 2469 2110
rect 4389 190 4390 2110
rect 2468 189 4390 190
rect 2178 62 2305 78
rect 2178 -62 2282 62
rect 2178 -78 2305 -62
rect 149 -190 2071 -189
rect 149 -2110 150 -190
rect 2070 -2110 2071 -190
rect 149 -2111 2071 -2110
rect -141 -2238 -14 -2222
rect -141 -2362 -37 -2238
rect -141 -2378 -14 -2362
rect -2170 -2490 -248 -2489
rect -2170 -4410 -2169 -2490
rect -249 -4410 -248 -2490
rect -2170 -4411 -248 -4410
rect -2460 -4538 -2333 -4522
rect -2460 -4600 -2356 -4538
rect -1261 -4600 -1157 -4411
rect -141 -4522 -94 -2378
rect -30 -4522 -14 -2378
rect 1058 -2489 1162 -2111
rect 2178 -2222 2225 -78
rect 2289 -2222 2305 -78
rect 3377 -189 3481 189
rect 4497 78 4544 2222
rect 4608 78 4624 2222
rect 4497 62 4624 78
rect 4497 -62 4601 62
rect 4497 -78 4624 -62
rect 2468 -190 4390 -189
rect 2468 -2110 2469 -190
rect 4389 -2110 4390 -190
rect 2468 -2111 4390 -2110
rect 2178 -2238 2305 -2222
rect 2178 -2362 2282 -2238
rect 2178 -2378 2305 -2362
rect 149 -2490 2071 -2489
rect 149 -4410 150 -2490
rect 2070 -4410 2071 -2490
rect 149 -4411 2071 -4410
rect -141 -4538 -14 -4522
rect -141 -4600 -37 -4538
rect 1058 -4600 1162 -4411
rect 2178 -4522 2225 -2378
rect 2289 -4522 2305 -2378
rect 3377 -2489 3481 -2111
rect 4497 -2222 4544 -78
rect 4608 -2222 4624 -78
rect 4497 -2238 4624 -2222
rect 4497 -2362 4601 -2238
rect 4497 -2378 4624 -2362
rect 2468 -2490 4390 -2489
rect 2468 -4410 2469 -2490
rect 4389 -4410 4390 -2490
rect 2468 -4411 4390 -4410
rect 2178 -4538 2305 -4522
rect 2178 -4600 2282 -4538
rect 3377 -4600 3481 -4411
rect 4497 -4522 4544 -2378
rect 4608 -4522 4624 -2378
rect 4497 -4538 4624 -4522
rect 4497 -4600 4601 -4538
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2329 2350 4529 4550
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
