magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1296 -1303 3850 2731
<< locali >>
rect 0 1396 2554 1432
rect 1855 724 1889 885
rect 1855 698 2051 724
rect 1694 690 2051 698
rect 2276 690 2395 724
rect 1694 664 1889 690
rect 2361 503 2395 690
rect 0 -18 2554 18
<< metal1 >>
rect 1841 859 1905 911
rect 1543 655 1607 707
rect 2346 477 2410 529
<< metal2 >>
rect 1858 871 1886 899
rect 369 692 423 756
rect 1549 661 1601 681
rect 1115 609 1601 661
rect 137 538 203 590
rect 2364 489 2392 517
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_3  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_3_0
timestamp 1626065694
transform 1 0 1970 0 1 0
box -36 -17 620 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_2  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_2_0
timestamp 1626065694
transform 1 0 1494 0 1 0
box -36 -17 512 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626065694
transform 1 0 1840 0 1 853
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626065694
transform 1 0 1844 0 1 852
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626065694
transform 1 0 2346 0 1 471
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626065694
transform 1 0 2349 0 1 470
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626065694
transform 1 0 1543 0 1 649
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626065694
transform 1 0 1546 0 1 648
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1626065694
transform 1 0 0 0 1 0
box -36 -43 1204 1467
<< labels >>
rlabel metal2 s 369 692 423 756 4 clk
rlabel metal2 s 137 538 203 590 4 D
rlabel metal2 s 2364 489 2392 517 4 Q
rlabel metal2 s 1858 871 1886 899 4 Qb
rlabel locali s 1277 1414 1277 1414 4 vdd
rlabel locali s 1277 0 1277 0 4 gnd
<< properties >>
string FIXED_BBOX 0 0 2554 1414
<< end >>
