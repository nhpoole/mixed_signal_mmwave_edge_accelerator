

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO sar_adc_controller 
  PIN clk 
    ANTENNAPARTIALMETALAREA 5.3802 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.74 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 11.4156 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.824 LAYER met3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9825 LAYER met3 ; 
    ANTENNAMAXAREACAR 14.4443 LAYER met3 ;
    ANTENNAMAXSIDEAREACAR 74.5771 LAYER met3 ;
    ANTENNAMAXCUTCAR 0.228125 LAYER via3 ;
  END clk
  PIN rst_n 
    ANTENNAPARTIALMETALAREA 9.8095 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 48.0025 LAYER met2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.503 LAYER met2 ; 
    ANTENNAMAXAREACAR 25.6 LAYER met2 ;
    ANTENNAMAXSIDEAREACAR 120.2 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAMAXCUTCAR 0.613121 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3 ;
    ANTENNAGATEAREA 2.889 LAYER met3 ; 
    ANTENNAMAXAREACAR 26.1666 LAYER met3 ;
    ANTENNAMAXSIDEAREACAR 123.384 LAYER met3 ;
    ANTENNAMAXCUTCAR 0.615368 LAYER via3 ;
  END rst_n
  PIN adc_start 
    ANTENNAPARTIALMETALAREA 5.1169 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.4765 LAYER met2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2 ; 
    ANTENNAMAXAREACAR 37.6333 LAYER met2 ;
    ANTENNAMAXSIDEAREACAR 185.956 LAYER met2 ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2 ;
  END adc_start
  PIN comparator_val 
    ANTENNAPARTIALMETALAREA 1.5784 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.784 LAYER met2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2 ; 
    ANTENNAMAXAREACAR 26.1226 LAYER met2 ;
    ANTENNAMAXSIDEAREACAR 128.495 LAYER met2 ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2 ;
  END comparator_val
  PIN run_adc_n 
    ANTENNADIFFAREA 0.429 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2 ;
  END run_adc_n
  PIN adc_val[7] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 2.9007 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3955 LAYER met2 ;
  END adc_val[7]
  PIN adc_val[6] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2 ;
  END adc_val[6]
  PIN adc_val[5] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2 ;
  END adc_val[5]
  PIN adc_val[4] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2 ;
  END adc_val[4]
  PIN adc_val[3] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 1.5308 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.546 LAYER met2 ;
  END adc_val[3]
  PIN adc_val[2] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 0.2414 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.099 LAYER met2 ;
  END adc_val[2]
  PIN adc_val[1] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 1.3362 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.573 LAYER met2 ;
  END adc_val[1]
  PIN adc_val[0] 
    ANTENNADIFFAREA 0.336 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 0.6222 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.003 LAYER met2 ;
  END adc_val[0]
  PIN out_valid 
    ANTENNADIFFAREA 0.429 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 4.5443 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6135 LAYER met2 ;
  END out_valid
END sar_adc_controller

END LIBRARY
