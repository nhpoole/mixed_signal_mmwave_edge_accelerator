magic
tech sky130A
magscale 1 2
timestamp 1622599880
<< metal3 >>
rect -950 -300 818 300
<< mimcap >>
rect -850 160 750 200
rect -850 -160 -810 160
rect 710 -160 750 160
rect -850 -200 750 -160
<< mimcapcontact >>
rect -810 -160 710 160
<< metal4 >>
rect -811 160 711 161
rect -811 -160 -810 160
rect 710 -160 711 160
rect -811 -161 711 -160
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -950 -300 850 300
string parameters w 8.00 l 2.00 val 35.8 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
