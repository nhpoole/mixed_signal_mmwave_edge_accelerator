magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -5896 -2875 5896 2875
<< pwell >>
rect -4636 -1553 4636 1553
<< nmoslvt >>
rect -4552 927 -3592 1527
rect -3534 927 -2574 1527
rect -2516 927 -1556 1527
rect -1498 927 -538 1527
rect -480 927 480 1527
rect 538 927 1498 1527
rect 1556 927 2516 1527
rect 2574 927 3534 1527
rect 3592 927 4552 1527
rect -4552 109 -3592 709
rect -3534 109 -2574 709
rect -2516 109 -1556 709
rect -1498 109 -538 709
rect -480 109 480 709
rect 538 109 1498 709
rect 1556 109 2516 709
rect 2574 109 3534 709
rect 3592 109 4552 709
rect -4552 -709 -3592 -109
rect -3534 -709 -2574 -109
rect -2516 -709 -1556 -109
rect -1498 -709 -538 -109
rect -480 -709 480 -109
rect 538 -709 1498 -109
rect 1556 -709 2516 -109
rect 2574 -709 3534 -109
rect 3592 -709 4552 -109
rect -4552 -1527 -3592 -927
rect -3534 -1527 -2574 -927
rect -2516 -1527 -1556 -927
rect -1498 -1527 -538 -927
rect -480 -1527 480 -927
rect 538 -1527 1498 -927
rect 1556 -1527 2516 -927
rect 2574 -1527 3534 -927
rect 3592 -1527 4552 -927
<< ndiff >>
rect -4610 1482 -4552 1527
rect -4610 1448 -4598 1482
rect -4564 1448 -4552 1482
rect -4610 1414 -4552 1448
rect -4610 1380 -4598 1414
rect -4564 1380 -4552 1414
rect -4610 1346 -4552 1380
rect -4610 1312 -4598 1346
rect -4564 1312 -4552 1346
rect -4610 1278 -4552 1312
rect -4610 1244 -4598 1278
rect -4564 1244 -4552 1278
rect -4610 1210 -4552 1244
rect -4610 1176 -4598 1210
rect -4564 1176 -4552 1210
rect -4610 1142 -4552 1176
rect -4610 1108 -4598 1142
rect -4564 1108 -4552 1142
rect -4610 1074 -4552 1108
rect -4610 1040 -4598 1074
rect -4564 1040 -4552 1074
rect -4610 1006 -4552 1040
rect -4610 972 -4598 1006
rect -4564 972 -4552 1006
rect -4610 927 -4552 972
rect -3592 1482 -3534 1527
rect -3592 1448 -3580 1482
rect -3546 1448 -3534 1482
rect -3592 1414 -3534 1448
rect -3592 1380 -3580 1414
rect -3546 1380 -3534 1414
rect -3592 1346 -3534 1380
rect -3592 1312 -3580 1346
rect -3546 1312 -3534 1346
rect -3592 1278 -3534 1312
rect -3592 1244 -3580 1278
rect -3546 1244 -3534 1278
rect -3592 1210 -3534 1244
rect -3592 1176 -3580 1210
rect -3546 1176 -3534 1210
rect -3592 1142 -3534 1176
rect -3592 1108 -3580 1142
rect -3546 1108 -3534 1142
rect -3592 1074 -3534 1108
rect -3592 1040 -3580 1074
rect -3546 1040 -3534 1074
rect -3592 1006 -3534 1040
rect -3592 972 -3580 1006
rect -3546 972 -3534 1006
rect -3592 927 -3534 972
rect -2574 1482 -2516 1527
rect -2574 1448 -2562 1482
rect -2528 1448 -2516 1482
rect -2574 1414 -2516 1448
rect -2574 1380 -2562 1414
rect -2528 1380 -2516 1414
rect -2574 1346 -2516 1380
rect -2574 1312 -2562 1346
rect -2528 1312 -2516 1346
rect -2574 1278 -2516 1312
rect -2574 1244 -2562 1278
rect -2528 1244 -2516 1278
rect -2574 1210 -2516 1244
rect -2574 1176 -2562 1210
rect -2528 1176 -2516 1210
rect -2574 1142 -2516 1176
rect -2574 1108 -2562 1142
rect -2528 1108 -2516 1142
rect -2574 1074 -2516 1108
rect -2574 1040 -2562 1074
rect -2528 1040 -2516 1074
rect -2574 1006 -2516 1040
rect -2574 972 -2562 1006
rect -2528 972 -2516 1006
rect -2574 927 -2516 972
rect -1556 1482 -1498 1527
rect -1556 1448 -1544 1482
rect -1510 1448 -1498 1482
rect -1556 1414 -1498 1448
rect -1556 1380 -1544 1414
rect -1510 1380 -1498 1414
rect -1556 1346 -1498 1380
rect -1556 1312 -1544 1346
rect -1510 1312 -1498 1346
rect -1556 1278 -1498 1312
rect -1556 1244 -1544 1278
rect -1510 1244 -1498 1278
rect -1556 1210 -1498 1244
rect -1556 1176 -1544 1210
rect -1510 1176 -1498 1210
rect -1556 1142 -1498 1176
rect -1556 1108 -1544 1142
rect -1510 1108 -1498 1142
rect -1556 1074 -1498 1108
rect -1556 1040 -1544 1074
rect -1510 1040 -1498 1074
rect -1556 1006 -1498 1040
rect -1556 972 -1544 1006
rect -1510 972 -1498 1006
rect -1556 927 -1498 972
rect -538 1482 -480 1527
rect -538 1448 -526 1482
rect -492 1448 -480 1482
rect -538 1414 -480 1448
rect -538 1380 -526 1414
rect -492 1380 -480 1414
rect -538 1346 -480 1380
rect -538 1312 -526 1346
rect -492 1312 -480 1346
rect -538 1278 -480 1312
rect -538 1244 -526 1278
rect -492 1244 -480 1278
rect -538 1210 -480 1244
rect -538 1176 -526 1210
rect -492 1176 -480 1210
rect -538 1142 -480 1176
rect -538 1108 -526 1142
rect -492 1108 -480 1142
rect -538 1074 -480 1108
rect -538 1040 -526 1074
rect -492 1040 -480 1074
rect -538 1006 -480 1040
rect -538 972 -526 1006
rect -492 972 -480 1006
rect -538 927 -480 972
rect 480 1482 538 1527
rect 480 1448 492 1482
rect 526 1448 538 1482
rect 480 1414 538 1448
rect 480 1380 492 1414
rect 526 1380 538 1414
rect 480 1346 538 1380
rect 480 1312 492 1346
rect 526 1312 538 1346
rect 480 1278 538 1312
rect 480 1244 492 1278
rect 526 1244 538 1278
rect 480 1210 538 1244
rect 480 1176 492 1210
rect 526 1176 538 1210
rect 480 1142 538 1176
rect 480 1108 492 1142
rect 526 1108 538 1142
rect 480 1074 538 1108
rect 480 1040 492 1074
rect 526 1040 538 1074
rect 480 1006 538 1040
rect 480 972 492 1006
rect 526 972 538 1006
rect 480 927 538 972
rect 1498 1482 1556 1527
rect 1498 1448 1510 1482
rect 1544 1448 1556 1482
rect 1498 1414 1556 1448
rect 1498 1380 1510 1414
rect 1544 1380 1556 1414
rect 1498 1346 1556 1380
rect 1498 1312 1510 1346
rect 1544 1312 1556 1346
rect 1498 1278 1556 1312
rect 1498 1244 1510 1278
rect 1544 1244 1556 1278
rect 1498 1210 1556 1244
rect 1498 1176 1510 1210
rect 1544 1176 1556 1210
rect 1498 1142 1556 1176
rect 1498 1108 1510 1142
rect 1544 1108 1556 1142
rect 1498 1074 1556 1108
rect 1498 1040 1510 1074
rect 1544 1040 1556 1074
rect 1498 1006 1556 1040
rect 1498 972 1510 1006
rect 1544 972 1556 1006
rect 1498 927 1556 972
rect 2516 1482 2574 1527
rect 2516 1448 2528 1482
rect 2562 1448 2574 1482
rect 2516 1414 2574 1448
rect 2516 1380 2528 1414
rect 2562 1380 2574 1414
rect 2516 1346 2574 1380
rect 2516 1312 2528 1346
rect 2562 1312 2574 1346
rect 2516 1278 2574 1312
rect 2516 1244 2528 1278
rect 2562 1244 2574 1278
rect 2516 1210 2574 1244
rect 2516 1176 2528 1210
rect 2562 1176 2574 1210
rect 2516 1142 2574 1176
rect 2516 1108 2528 1142
rect 2562 1108 2574 1142
rect 2516 1074 2574 1108
rect 2516 1040 2528 1074
rect 2562 1040 2574 1074
rect 2516 1006 2574 1040
rect 2516 972 2528 1006
rect 2562 972 2574 1006
rect 2516 927 2574 972
rect 3534 1482 3592 1527
rect 3534 1448 3546 1482
rect 3580 1448 3592 1482
rect 3534 1414 3592 1448
rect 3534 1380 3546 1414
rect 3580 1380 3592 1414
rect 3534 1346 3592 1380
rect 3534 1312 3546 1346
rect 3580 1312 3592 1346
rect 3534 1278 3592 1312
rect 3534 1244 3546 1278
rect 3580 1244 3592 1278
rect 3534 1210 3592 1244
rect 3534 1176 3546 1210
rect 3580 1176 3592 1210
rect 3534 1142 3592 1176
rect 3534 1108 3546 1142
rect 3580 1108 3592 1142
rect 3534 1074 3592 1108
rect 3534 1040 3546 1074
rect 3580 1040 3592 1074
rect 3534 1006 3592 1040
rect 3534 972 3546 1006
rect 3580 972 3592 1006
rect 3534 927 3592 972
rect 4552 1482 4610 1527
rect 4552 1448 4564 1482
rect 4598 1448 4610 1482
rect 4552 1414 4610 1448
rect 4552 1380 4564 1414
rect 4598 1380 4610 1414
rect 4552 1346 4610 1380
rect 4552 1312 4564 1346
rect 4598 1312 4610 1346
rect 4552 1278 4610 1312
rect 4552 1244 4564 1278
rect 4598 1244 4610 1278
rect 4552 1210 4610 1244
rect 4552 1176 4564 1210
rect 4598 1176 4610 1210
rect 4552 1142 4610 1176
rect 4552 1108 4564 1142
rect 4598 1108 4610 1142
rect 4552 1074 4610 1108
rect 4552 1040 4564 1074
rect 4598 1040 4610 1074
rect 4552 1006 4610 1040
rect 4552 972 4564 1006
rect 4598 972 4610 1006
rect 4552 927 4610 972
rect -4610 664 -4552 709
rect -4610 630 -4598 664
rect -4564 630 -4552 664
rect -4610 596 -4552 630
rect -4610 562 -4598 596
rect -4564 562 -4552 596
rect -4610 528 -4552 562
rect -4610 494 -4598 528
rect -4564 494 -4552 528
rect -4610 460 -4552 494
rect -4610 426 -4598 460
rect -4564 426 -4552 460
rect -4610 392 -4552 426
rect -4610 358 -4598 392
rect -4564 358 -4552 392
rect -4610 324 -4552 358
rect -4610 290 -4598 324
rect -4564 290 -4552 324
rect -4610 256 -4552 290
rect -4610 222 -4598 256
rect -4564 222 -4552 256
rect -4610 188 -4552 222
rect -4610 154 -4598 188
rect -4564 154 -4552 188
rect -4610 109 -4552 154
rect -3592 664 -3534 709
rect -3592 630 -3580 664
rect -3546 630 -3534 664
rect -3592 596 -3534 630
rect -3592 562 -3580 596
rect -3546 562 -3534 596
rect -3592 528 -3534 562
rect -3592 494 -3580 528
rect -3546 494 -3534 528
rect -3592 460 -3534 494
rect -3592 426 -3580 460
rect -3546 426 -3534 460
rect -3592 392 -3534 426
rect -3592 358 -3580 392
rect -3546 358 -3534 392
rect -3592 324 -3534 358
rect -3592 290 -3580 324
rect -3546 290 -3534 324
rect -3592 256 -3534 290
rect -3592 222 -3580 256
rect -3546 222 -3534 256
rect -3592 188 -3534 222
rect -3592 154 -3580 188
rect -3546 154 -3534 188
rect -3592 109 -3534 154
rect -2574 664 -2516 709
rect -2574 630 -2562 664
rect -2528 630 -2516 664
rect -2574 596 -2516 630
rect -2574 562 -2562 596
rect -2528 562 -2516 596
rect -2574 528 -2516 562
rect -2574 494 -2562 528
rect -2528 494 -2516 528
rect -2574 460 -2516 494
rect -2574 426 -2562 460
rect -2528 426 -2516 460
rect -2574 392 -2516 426
rect -2574 358 -2562 392
rect -2528 358 -2516 392
rect -2574 324 -2516 358
rect -2574 290 -2562 324
rect -2528 290 -2516 324
rect -2574 256 -2516 290
rect -2574 222 -2562 256
rect -2528 222 -2516 256
rect -2574 188 -2516 222
rect -2574 154 -2562 188
rect -2528 154 -2516 188
rect -2574 109 -2516 154
rect -1556 664 -1498 709
rect -1556 630 -1544 664
rect -1510 630 -1498 664
rect -1556 596 -1498 630
rect -1556 562 -1544 596
rect -1510 562 -1498 596
rect -1556 528 -1498 562
rect -1556 494 -1544 528
rect -1510 494 -1498 528
rect -1556 460 -1498 494
rect -1556 426 -1544 460
rect -1510 426 -1498 460
rect -1556 392 -1498 426
rect -1556 358 -1544 392
rect -1510 358 -1498 392
rect -1556 324 -1498 358
rect -1556 290 -1544 324
rect -1510 290 -1498 324
rect -1556 256 -1498 290
rect -1556 222 -1544 256
rect -1510 222 -1498 256
rect -1556 188 -1498 222
rect -1556 154 -1544 188
rect -1510 154 -1498 188
rect -1556 109 -1498 154
rect -538 664 -480 709
rect -538 630 -526 664
rect -492 630 -480 664
rect -538 596 -480 630
rect -538 562 -526 596
rect -492 562 -480 596
rect -538 528 -480 562
rect -538 494 -526 528
rect -492 494 -480 528
rect -538 460 -480 494
rect -538 426 -526 460
rect -492 426 -480 460
rect -538 392 -480 426
rect -538 358 -526 392
rect -492 358 -480 392
rect -538 324 -480 358
rect -538 290 -526 324
rect -492 290 -480 324
rect -538 256 -480 290
rect -538 222 -526 256
rect -492 222 -480 256
rect -538 188 -480 222
rect -538 154 -526 188
rect -492 154 -480 188
rect -538 109 -480 154
rect 480 664 538 709
rect 480 630 492 664
rect 526 630 538 664
rect 480 596 538 630
rect 480 562 492 596
rect 526 562 538 596
rect 480 528 538 562
rect 480 494 492 528
rect 526 494 538 528
rect 480 460 538 494
rect 480 426 492 460
rect 526 426 538 460
rect 480 392 538 426
rect 480 358 492 392
rect 526 358 538 392
rect 480 324 538 358
rect 480 290 492 324
rect 526 290 538 324
rect 480 256 538 290
rect 480 222 492 256
rect 526 222 538 256
rect 480 188 538 222
rect 480 154 492 188
rect 526 154 538 188
rect 480 109 538 154
rect 1498 664 1556 709
rect 1498 630 1510 664
rect 1544 630 1556 664
rect 1498 596 1556 630
rect 1498 562 1510 596
rect 1544 562 1556 596
rect 1498 528 1556 562
rect 1498 494 1510 528
rect 1544 494 1556 528
rect 1498 460 1556 494
rect 1498 426 1510 460
rect 1544 426 1556 460
rect 1498 392 1556 426
rect 1498 358 1510 392
rect 1544 358 1556 392
rect 1498 324 1556 358
rect 1498 290 1510 324
rect 1544 290 1556 324
rect 1498 256 1556 290
rect 1498 222 1510 256
rect 1544 222 1556 256
rect 1498 188 1556 222
rect 1498 154 1510 188
rect 1544 154 1556 188
rect 1498 109 1556 154
rect 2516 664 2574 709
rect 2516 630 2528 664
rect 2562 630 2574 664
rect 2516 596 2574 630
rect 2516 562 2528 596
rect 2562 562 2574 596
rect 2516 528 2574 562
rect 2516 494 2528 528
rect 2562 494 2574 528
rect 2516 460 2574 494
rect 2516 426 2528 460
rect 2562 426 2574 460
rect 2516 392 2574 426
rect 2516 358 2528 392
rect 2562 358 2574 392
rect 2516 324 2574 358
rect 2516 290 2528 324
rect 2562 290 2574 324
rect 2516 256 2574 290
rect 2516 222 2528 256
rect 2562 222 2574 256
rect 2516 188 2574 222
rect 2516 154 2528 188
rect 2562 154 2574 188
rect 2516 109 2574 154
rect 3534 664 3592 709
rect 3534 630 3546 664
rect 3580 630 3592 664
rect 3534 596 3592 630
rect 3534 562 3546 596
rect 3580 562 3592 596
rect 3534 528 3592 562
rect 3534 494 3546 528
rect 3580 494 3592 528
rect 3534 460 3592 494
rect 3534 426 3546 460
rect 3580 426 3592 460
rect 3534 392 3592 426
rect 3534 358 3546 392
rect 3580 358 3592 392
rect 3534 324 3592 358
rect 3534 290 3546 324
rect 3580 290 3592 324
rect 3534 256 3592 290
rect 3534 222 3546 256
rect 3580 222 3592 256
rect 3534 188 3592 222
rect 3534 154 3546 188
rect 3580 154 3592 188
rect 3534 109 3592 154
rect 4552 664 4610 709
rect 4552 630 4564 664
rect 4598 630 4610 664
rect 4552 596 4610 630
rect 4552 562 4564 596
rect 4598 562 4610 596
rect 4552 528 4610 562
rect 4552 494 4564 528
rect 4598 494 4610 528
rect 4552 460 4610 494
rect 4552 426 4564 460
rect 4598 426 4610 460
rect 4552 392 4610 426
rect 4552 358 4564 392
rect 4598 358 4610 392
rect 4552 324 4610 358
rect 4552 290 4564 324
rect 4598 290 4610 324
rect 4552 256 4610 290
rect 4552 222 4564 256
rect 4598 222 4610 256
rect 4552 188 4610 222
rect 4552 154 4564 188
rect 4598 154 4610 188
rect 4552 109 4610 154
rect -4610 -154 -4552 -109
rect -4610 -188 -4598 -154
rect -4564 -188 -4552 -154
rect -4610 -222 -4552 -188
rect -4610 -256 -4598 -222
rect -4564 -256 -4552 -222
rect -4610 -290 -4552 -256
rect -4610 -324 -4598 -290
rect -4564 -324 -4552 -290
rect -4610 -358 -4552 -324
rect -4610 -392 -4598 -358
rect -4564 -392 -4552 -358
rect -4610 -426 -4552 -392
rect -4610 -460 -4598 -426
rect -4564 -460 -4552 -426
rect -4610 -494 -4552 -460
rect -4610 -528 -4598 -494
rect -4564 -528 -4552 -494
rect -4610 -562 -4552 -528
rect -4610 -596 -4598 -562
rect -4564 -596 -4552 -562
rect -4610 -630 -4552 -596
rect -4610 -664 -4598 -630
rect -4564 -664 -4552 -630
rect -4610 -709 -4552 -664
rect -3592 -154 -3534 -109
rect -3592 -188 -3580 -154
rect -3546 -188 -3534 -154
rect -3592 -222 -3534 -188
rect -3592 -256 -3580 -222
rect -3546 -256 -3534 -222
rect -3592 -290 -3534 -256
rect -3592 -324 -3580 -290
rect -3546 -324 -3534 -290
rect -3592 -358 -3534 -324
rect -3592 -392 -3580 -358
rect -3546 -392 -3534 -358
rect -3592 -426 -3534 -392
rect -3592 -460 -3580 -426
rect -3546 -460 -3534 -426
rect -3592 -494 -3534 -460
rect -3592 -528 -3580 -494
rect -3546 -528 -3534 -494
rect -3592 -562 -3534 -528
rect -3592 -596 -3580 -562
rect -3546 -596 -3534 -562
rect -3592 -630 -3534 -596
rect -3592 -664 -3580 -630
rect -3546 -664 -3534 -630
rect -3592 -709 -3534 -664
rect -2574 -154 -2516 -109
rect -2574 -188 -2562 -154
rect -2528 -188 -2516 -154
rect -2574 -222 -2516 -188
rect -2574 -256 -2562 -222
rect -2528 -256 -2516 -222
rect -2574 -290 -2516 -256
rect -2574 -324 -2562 -290
rect -2528 -324 -2516 -290
rect -2574 -358 -2516 -324
rect -2574 -392 -2562 -358
rect -2528 -392 -2516 -358
rect -2574 -426 -2516 -392
rect -2574 -460 -2562 -426
rect -2528 -460 -2516 -426
rect -2574 -494 -2516 -460
rect -2574 -528 -2562 -494
rect -2528 -528 -2516 -494
rect -2574 -562 -2516 -528
rect -2574 -596 -2562 -562
rect -2528 -596 -2516 -562
rect -2574 -630 -2516 -596
rect -2574 -664 -2562 -630
rect -2528 -664 -2516 -630
rect -2574 -709 -2516 -664
rect -1556 -154 -1498 -109
rect -1556 -188 -1544 -154
rect -1510 -188 -1498 -154
rect -1556 -222 -1498 -188
rect -1556 -256 -1544 -222
rect -1510 -256 -1498 -222
rect -1556 -290 -1498 -256
rect -1556 -324 -1544 -290
rect -1510 -324 -1498 -290
rect -1556 -358 -1498 -324
rect -1556 -392 -1544 -358
rect -1510 -392 -1498 -358
rect -1556 -426 -1498 -392
rect -1556 -460 -1544 -426
rect -1510 -460 -1498 -426
rect -1556 -494 -1498 -460
rect -1556 -528 -1544 -494
rect -1510 -528 -1498 -494
rect -1556 -562 -1498 -528
rect -1556 -596 -1544 -562
rect -1510 -596 -1498 -562
rect -1556 -630 -1498 -596
rect -1556 -664 -1544 -630
rect -1510 -664 -1498 -630
rect -1556 -709 -1498 -664
rect -538 -154 -480 -109
rect -538 -188 -526 -154
rect -492 -188 -480 -154
rect -538 -222 -480 -188
rect -538 -256 -526 -222
rect -492 -256 -480 -222
rect -538 -290 -480 -256
rect -538 -324 -526 -290
rect -492 -324 -480 -290
rect -538 -358 -480 -324
rect -538 -392 -526 -358
rect -492 -392 -480 -358
rect -538 -426 -480 -392
rect -538 -460 -526 -426
rect -492 -460 -480 -426
rect -538 -494 -480 -460
rect -538 -528 -526 -494
rect -492 -528 -480 -494
rect -538 -562 -480 -528
rect -538 -596 -526 -562
rect -492 -596 -480 -562
rect -538 -630 -480 -596
rect -538 -664 -526 -630
rect -492 -664 -480 -630
rect -538 -709 -480 -664
rect 480 -154 538 -109
rect 480 -188 492 -154
rect 526 -188 538 -154
rect 480 -222 538 -188
rect 480 -256 492 -222
rect 526 -256 538 -222
rect 480 -290 538 -256
rect 480 -324 492 -290
rect 526 -324 538 -290
rect 480 -358 538 -324
rect 480 -392 492 -358
rect 526 -392 538 -358
rect 480 -426 538 -392
rect 480 -460 492 -426
rect 526 -460 538 -426
rect 480 -494 538 -460
rect 480 -528 492 -494
rect 526 -528 538 -494
rect 480 -562 538 -528
rect 480 -596 492 -562
rect 526 -596 538 -562
rect 480 -630 538 -596
rect 480 -664 492 -630
rect 526 -664 538 -630
rect 480 -709 538 -664
rect 1498 -154 1556 -109
rect 1498 -188 1510 -154
rect 1544 -188 1556 -154
rect 1498 -222 1556 -188
rect 1498 -256 1510 -222
rect 1544 -256 1556 -222
rect 1498 -290 1556 -256
rect 1498 -324 1510 -290
rect 1544 -324 1556 -290
rect 1498 -358 1556 -324
rect 1498 -392 1510 -358
rect 1544 -392 1556 -358
rect 1498 -426 1556 -392
rect 1498 -460 1510 -426
rect 1544 -460 1556 -426
rect 1498 -494 1556 -460
rect 1498 -528 1510 -494
rect 1544 -528 1556 -494
rect 1498 -562 1556 -528
rect 1498 -596 1510 -562
rect 1544 -596 1556 -562
rect 1498 -630 1556 -596
rect 1498 -664 1510 -630
rect 1544 -664 1556 -630
rect 1498 -709 1556 -664
rect 2516 -154 2574 -109
rect 2516 -188 2528 -154
rect 2562 -188 2574 -154
rect 2516 -222 2574 -188
rect 2516 -256 2528 -222
rect 2562 -256 2574 -222
rect 2516 -290 2574 -256
rect 2516 -324 2528 -290
rect 2562 -324 2574 -290
rect 2516 -358 2574 -324
rect 2516 -392 2528 -358
rect 2562 -392 2574 -358
rect 2516 -426 2574 -392
rect 2516 -460 2528 -426
rect 2562 -460 2574 -426
rect 2516 -494 2574 -460
rect 2516 -528 2528 -494
rect 2562 -528 2574 -494
rect 2516 -562 2574 -528
rect 2516 -596 2528 -562
rect 2562 -596 2574 -562
rect 2516 -630 2574 -596
rect 2516 -664 2528 -630
rect 2562 -664 2574 -630
rect 2516 -709 2574 -664
rect 3534 -154 3592 -109
rect 3534 -188 3546 -154
rect 3580 -188 3592 -154
rect 3534 -222 3592 -188
rect 3534 -256 3546 -222
rect 3580 -256 3592 -222
rect 3534 -290 3592 -256
rect 3534 -324 3546 -290
rect 3580 -324 3592 -290
rect 3534 -358 3592 -324
rect 3534 -392 3546 -358
rect 3580 -392 3592 -358
rect 3534 -426 3592 -392
rect 3534 -460 3546 -426
rect 3580 -460 3592 -426
rect 3534 -494 3592 -460
rect 3534 -528 3546 -494
rect 3580 -528 3592 -494
rect 3534 -562 3592 -528
rect 3534 -596 3546 -562
rect 3580 -596 3592 -562
rect 3534 -630 3592 -596
rect 3534 -664 3546 -630
rect 3580 -664 3592 -630
rect 3534 -709 3592 -664
rect 4552 -154 4610 -109
rect 4552 -188 4564 -154
rect 4598 -188 4610 -154
rect 4552 -222 4610 -188
rect 4552 -256 4564 -222
rect 4598 -256 4610 -222
rect 4552 -290 4610 -256
rect 4552 -324 4564 -290
rect 4598 -324 4610 -290
rect 4552 -358 4610 -324
rect 4552 -392 4564 -358
rect 4598 -392 4610 -358
rect 4552 -426 4610 -392
rect 4552 -460 4564 -426
rect 4598 -460 4610 -426
rect 4552 -494 4610 -460
rect 4552 -528 4564 -494
rect 4598 -528 4610 -494
rect 4552 -562 4610 -528
rect 4552 -596 4564 -562
rect 4598 -596 4610 -562
rect 4552 -630 4610 -596
rect 4552 -664 4564 -630
rect 4598 -664 4610 -630
rect 4552 -709 4610 -664
rect -4610 -972 -4552 -927
rect -4610 -1006 -4598 -972
rect -4564 -1006 -4552 -972
rect -4610 -1040 -4552 -1006
rect -4610 -1074 -4598 -1040
rect -4564 -1074 -4552 -1040
rect -4610 -1108 -4552 -1074
rect -4610 -1142 -4598 -1108
rect -4564 -1142 -4552 -1108
rect -4610 -1176 -4552 -1142
rect -4610 -1210 -4598 -1176
rect -4564 -1210 -4552 -1176
rect -4610 -1244 -4552 -1210
rect -4610 -1278 -4598 -1244
rect -4564 -1278 -4552 -1244
rect -4610 -1312 -4552 -1278
rect -4610 -1346 -4598 -1312
rect -4564 -1346 -4552 -1312
rect -4610 -1380 -4552 -1346
rect -4610 -1414 -4598 -1380
rect -4564 -1414 -4552 -1380
rect -4610 -1448 -4552 -1414
rect -4610 -1482 -4598 -1448
rect -4564 -1482 -4552 -1448
rect -4610 -1527 -4552 -1482
rect -3592 -972 -3534 -927
rect -3592 -1006 -3580 -972
rect -3546 -1006 -3534 -972
rect -3592 -1040 -3534 -1006
rect -3592 -1074 -3580 -1040
rect -3546 -1074 -3534 -1040
rect -3592 -1108 -3534 -1074
rect -3592 -1142 -3580 -1108
rect -3546 -1142 -3534 -1108
rect -3592 -1176 -3534 -1142
rect -3592 -1210 -3580 -1176
rect -3546 -1210 -3534 -1176
rect -3592 -1244 -3534 -1210
rect -3592 -1278 -3580 -1244
rect -3546 -1278 -3534 -1244
rect -3592 -1312 -3534 -1278
rect -3592 -1346 -3580 -1312
rect -3546 -1346 -3534 -1312
rect -3592 -1380 -3534 -1346
rect -3592 -1414 -3580 -1380
rect -3546 -1414 -3534 -1380
rect -3592 -1448 -3534 -1414
rect -3592 -1482 -3580 -1448
rect -3546 -1482 -3534 -1448
rect -3592 -1527 -3534 -1482
rect -2574 -972 -2516 -927
rect -2574 -1006 -2562 -972
rect -2528 -1006 -2516 -972
rect -2574 -1040 -2516 -1006
rect -2574 -1074 -2562 -1040
rect -2528 -1074 -2516 -1040
rect -2574 -1108 -2516 -1074
rect -2574 -1142 -2562 -1108
rect -2528 -1142 -2516 -1108
rect -2574 -1176 -2516 -1142
rect -2574 -1210 -2562 -1176
rect -2528 -1210 -2516 -1176
rect -2574 -1244 -2516 -1210
rect -2574 -1278 -2562 -1244
rect -2528 -1278 -2516 -1244
rect -2574 -1312 -2516 -1278
rect -2574 -1346 -2562 -1312
rect -2528 -1346 -2516 -1312
rect -2574 -1380 -2516 -1346
rect -2574 -1414 -2562 -1380
rect -2528 -1414 -2516 -1380
rect -2574 -1448 -2516 -1414
rect -2574 -1482 -2562 -1448
rect -2528 -1482 -2516 -1448
rect -2574 -1527 -2516 -1482
rect -1556 -972 -1498 -927
rect -1556 -1006 -1544 -972
rect -1510 -1006 -1498 -972
rect -1556 -1040 -1498 -1006
rect -1556 -1074 -1544 -1040
rect -1510 -1074 -1498 -1040
rect -1556 -1108 -1498 -1074
rect -1556 -1142 -1544 -1108
rect -1510 -1142 -1498 -1108
rect -1556 -1176 -1498 -1142
rect -1556 -1210 -1544 -1176
rect -1510 -1210 -1498 -1176
rect -1556 -1244 -1498 -1210
rect -1556 -1278 -1544 -1244
rect -1510 -1278 -1498 -1244
rect -1556 -1312 -1498 -1278
rect -1556 -1346 -1544 -1312
rect -1510 -1346 -1498 -1312
rect -1556 -1380 -1498 -1346
rect -1556 -1414 -1544 -1380
rect -1510 -1414 -1498 -1380
rect -1556 -1448 -1498 -1414
rect -1556 -1482 -1544 -1448
rect -1510 -1482 -1498 -1448
rect -1556 -1527 -1498 -1482
rect -538 -972 -480 -927
rect -538 -1006 -526 -972
rect -492 -1006 -480 -972
rect -538 -1040 -480 -1006
rect -538 -1074 -526 -1040
rect -492 -1074 -480 -1040
rect -538 -1108 -480 -1074
rect -538 -1142 -526 -1108
rect -492 -1142 -480 -1108
rect -538 -1176 -480 -1142
rect -538 -1210 -526 -1176
rect -492 -1210 -480 -1176
rect -538 -1244 -480 -1210
rect -538 -1278 -526 -1244
rect -492 -1278 -480 -1244
rect -538 -1312 -480 -1278
rect -538 -1346 -526 -1312
rect -492 -1346 -480 -1312
rect -538 -1380 -480 -1346
rect -538 -1414 -526 -1380
rect -492 -1414 -480 -1380
rect -538 -1448 -480 -1414
rect -538 -1482 -526 -1448
rect -492 -1482 -480 -1448
rect -538 -1527 -480 -1482
rect 480 -972 538 -927
rect 480 -1006 492 -972
rect 526 -1006 538 -972
rect 480 -1040 538 -1006
rect 480 -1074 492 -1040
rect 526 -1074 538 -1040
rect 480 -1108 538 -1074
rect 480 -1142 492 -1108
rect 526 -1142 538 -1108
rect 480 -1176 538 -1142
rect 480 -1210 492 -1176
rect 526 -1210 538 -1176
rect 480 -1244 538 -1210
rect 480 -1278 492 -1244
rect 526 -1278 538 -1244
rect 480 -1312 538 -1278
rect 480 -1346 492 -1312
rect 526 -1346 538 -1312
rect 480 -1380 538 -1346
rect 480 -1414 492 -1380
rect 526 -1414 538 -1380
rect 480 -1448 538 -1414
rect 480 -1482 492 -1448
rect 526 -1482 538 -1448
rect 480 -1527 538 -1482
rect 1498 -972 1556 -927
rect 1498 -1006 1510 -972
rect 1544 -1006 1556 -972
rect 1498 -1040 1556 -1006
rect 1498 -1074 1510 -1040
rect 1544 -1074 1556 -1040
rect 1498 -1108 1556 -1074
rect 1498 -1142 1510 -1108
rect 1544 -1142 1556 -1108
rect 1498 -1176 1556 -1142
rect 1498 -1210 1510 -1176
rect 1544 -1210 1556 -1176
rect 1498 -1244 1556 -1210
rect 1498 -1278 1510 -1244
rect 1544 -1278 1556 -1244
rect 1498 -1312 1556 -1278
rect 1498 -1346 1510 -1312
rect 1544 -1346 1556 -1312
rect 1498 -1380 1556 -1346
rect 1498 -1414 1510 -1380
rect 1544 -1414 1556 -1380
rect 1498 -1448 1556 -1414
rect 1498 -1482 1510 -1448
rect 1544 -1482 1556 -1448
rect 1498 -1527 1556 -1482
rect 2516 -972 2574 -927
rect 2516 -1006 2528 -972
rect 2562 -1006 2574 -972
rect 2516 -1040 2574 -1006
rect 2516 -1074 2528 -1040
rect 2562 -1074 2574 -1040
rect 2516 -1108 2574 -1074
rect 2516 -1142 2528 -1108
rect 2562 -1142 2574 -1108
rect 2516 -1176 2574 -1142
rect 2516 -1210 2528 -1176
rect 2562 -1210 2574 -1176
rect 2516 -1244 2574 -1210
rect 2516 -1278 2528 -1244
rect 2562 -1278 2574 -1244
rect 2516 -1312 2574 -1278
rect 2516 -1346 2528 -1312
rect 2562 -1346 2574 -1312
rect 2516 -1380 2574 -1346
rect 2516 -1414 2528 -1380
rect 2562 -1414 2574 -1380
rect 2516 -1448 2574 -1414
rect 2516 -1482 2528 -1448
rect 2562 -1482 2574 -1448
rect 2516 -1527 2574 -1482
rect 3534 -972 3592 -927
rect 3534 -1006 3546 -972
rect 3580 -1006 3592 -972
rect 3534 -1040 3592 -1006
rect 3534 -1074 3546 -1040
rect 3580 -1074 3592 -1040
rect 3534 -1108 3592 -1074
rect 3534 -1142 3546 -1108
rect 3580 -1142 3592 -1108
rect 3534 -1176 3592 -1142
rect 3534 -1210 3546 -1176
rect 3580 -1210 3592 -1176
rect 3534 -1244 3592 -1210
rect 3534 -1278 3546 -1244
rect 3580 -1278 3592 -1244
rect 3534 -1312 3592 -1278
rect 3534 -1346 3546 -1312
rect 3580 -1346 3592 -1312
rect 3534 -1380 3592 -1346
rect 3534 -1414 3546 -1380
rect 3580 -1414 3592 -1380
rect 3534 -1448 3592 -1414
rect 3534 -1482 3546 -1448
rect 3580 -1482 3592 -1448
rect 3534 -1527 3592 -1482
rect 4552 -972 4610 -927
rect 4552 -1006 4564 -972
rect 4598 -1006 4610 -972
rect 4552 -1040 4610 -1006
rect 4552 -1074 4564 -1040
rect 4598 -1074 4610 -1040
rect 4552 -1108 4610 -1074
rect 4552 -1142 4564 -1108
rect 4598 -1142 4610 -1108
rect 4552 -1176 4610 -1142
rect 4552 -1210 4564 -1176
rect 4598 -1210 4610 -1176
rect 4552 -1244 4610 -1210
rect 4552 -1278 4564 -1244
rect 4598 -1278 4610 -1244
rect 4552 -1312 4610 -1278
rect 4552 -1346 4564 -1312
rect 4598 -1346 4610 -1312
rect 4552 -1380 4610 -1346
rect 4552 -1414 4564 -1380
rect 4598 -1414 4610 -1380
rect 4552 -1448 4610 -1414
rect 4552 -1482 4564 -1448
rect 4598 -1482 4610 -1448
rect 4552 -1527 4610 -1482
<< ndiffc >>
rect -4598 1448 -4564 1482
rect -4598 1380 -4564 1414
rect -4598 1312 -4564 1346
rect -4598 1244 -4564 1278
rect -4598 1176 -4564 1210
rect -4598 1108 -4564 1142
rect -4598 1040 -4564 1074
rect -4598 972 -4564 1006
rect -3580 1448 -3546 1482
rect -3580 1380 -3546 1414
rect -3580 1312 -3546 1346
rect -3580 1244 -3546 1278
rect -3580 1176 -3546 1210
rect -3580 1108 -3546 1142
rect -3580 1040 -3546 1074
rect -3580 972 -3546 1006
rect -2562 1448 -2528 1482
rect -2562 1380 -2528 1414
rect -2562 1312 -2528 1346
rect -2562 1244 -2528 1278
rect -2562 1176 -2528 1210
rect -2562 1108 -2528 1142
rect -2562 1040 -2528 1074
rect -2562 972 -2528 1006
rect -1544 1448 -1510 1482
rect -1544 1380 -1510 1414
rect -1544 1312 -1510 1346
rect -1544 1244 -1510 1278
rect -1544 1176 -1510 1210
rect -1544 1108 -1510 1142
rect -1544 1040 -1510 1074
rect -1544 972 -1510 1006
rect -526 1448 -492 1482
rect -526 1380 -492 1414
rect -526 1312 -492 1346
rect -526 1244 -492 1278
rect -526 1176 -492 1210
rect -526 1108 -492 1142
rect -526 1040 -492 1074
rect -526 972 -492 1006
rect 492 1448 526 1482
rect 492 1380 526 1414
rect 492 1312 526 1346
rect 492 1244 526 1278
rect 492 1176 526 1210
rect 492 1108 526 1142
rect 492 1040 526 1074
rect 492 972 526 1006
rect 1510 1448 1544 1482
rect 1510 1380 1544 1414
rect 1510 1312 1544 1346
rect 1510 1244 1544 1278
rect 1510 1176 1544 1210
rect 1510 1108 1544 1142
rect 1510 1040 1544 1074
rect 1510 972 1544 1006
rect 2528 1448 2562 1482
rect 2528 1380 2562 1414
rect 2528 1312 2562 1346
rect 2528 1244 2562 1278
rect 2528 1176 2562 1210
rect 2528 1108 2562 1142
rect 2528 1040 2562 1074
rect 2528 972 2562 1006
rect 3546 1448 3580 1482
rect 3546 1380 3580 1414
rect 3546 1312 3580 1346
rect 3546 1244 3580 1278
rect 3546 1176 3580 1210
rect 3546 1108 3580 1142
rect 3546 1040 3580 1074
rect 3546 972 3580 1006
rect 4564 1448 4598 1482
rect 4564 1380 4598 1414
rect 4564 1312 4598 1346
rect 4564 1244 4598 1278
rect 4564 1176 4598 1210
rect 4564 1108 4598 1142
rect 4564 1040 4598 1074
rect 4564 972 4598 1006
rect -4598 630 -4564 664
rect -4598 562 -4564 596
rect -4598 494 -4564 528
rect -4598 426 -4564 460
rect -4598 358 -4564 392
rect -4598 290 -4564 324
rect -4598 222 -4564 256
rect -4598 154 -4564 188
rect -3580 630 -3546 664
rect -3580 562 -3546 596
rect -3580 494 -3546 528
rect -3580 426 -3546 460
rect -3580 358 -3546 392
rect -3580 290 -3546 324
rect -3580 222 -3546 256
rect -3580 154 -3546 188
rect -2562 630 -2528 664
rect -2562 562 -2528 596
rect -2562 494 -2528 528
rect -2562 426 -2528 460
rect -2562 358 -2528 392
rect -2562 290 -2528 324
rect -2562 222 -2528 256
rect -2562 154 -2528 188
rect -1544 630 -1510 664
rect -1544 562 -1510 596
rect -1544 494 -1510 528
rect -1544 426 -1510 460
rect -1544 358 -1510 392
rect -1544 290 -1510 324
rect -1544 222 -1510 256
rect -1544 154 -1510 188
rect -526 630 -492 664
rect -526 562 -492 596
rect -526 494 -492 528
rect -526 426 -492 460
rect -526 358 -492 392
rect -526 290 -492 324
rect -526 222 -492 256
rect -526 154 -492 188
rect 492 630 526 664
rect 492 562 526 596
rect 492 494 526 528
rect 492 426 526 460
rect 492 358 526 392
rect 492 290 526 324
rect 492 222 526 256
rect 492 154 526 188
rect 1510 630 1544 664
rect 1510 562 1544 596
rect 1510 494 1544 528
rect 1510 426 1544 460
rect 1510 358 1544 392
rect 1510 290 1544 324
rect 1510 222 1544 256
rect 1510 154 1544 188
rect 2528 630 2562 664
rect 2528 562 2562 596
rect 2528 494 2562 528
rect 2528 426 2562 460
rect 2528 358 2562 392
rect 2528 290 2562 324
rect 2528 222 2562 256
rect 2528 154 2562 188
rect 3546 630 3580 664
rect 3546 562 3580 596
rect 3546 494 3580 528
rect 3546 426 3580 460
rect 3546 358 3580 392
rect 3546 290 3580 324
rect 3546 222 3580 256
rect 3546 154 3580 188
rect 4564 630 4598 664
rect 4564 562 4598 596
rect 4564 494 4598 528
rect 4564 426 4598 460
rect 4564 358 4598 392
rect 4564 290 4598 324
rect 4564 222 4598 256
rect 4564 154 4598 188
rect -4598 -188 -4564 -154
rect -4598 -256 -4564 -222
rect -4598 -324 -4564 -290
rect -4598 -392 -4564 -358
rect -4598 -460 -4564 -426
rect -4598 -528 -4564 -494
rect -4598 -596 -4564 -562
rect -4598 -664 -4564 -630
rect -3580 -188 -3546 -154
rect -3580 -256 -3546 -222
rect -3580 -324 -3546 -290
rect -3580 -392 -3546 -358
rect -3580 -460 -3546 -426
rect -3580 -528 -3546 -494
rect -3580 -596 -3546 -562
rect -3580 -664 -3546 -630
rect -2562 -188 -2528 -154
rect -2562 -256 -2528 -222
rect -2562 -324 -2528 -290
rect -2562 -392 -2528 -358
rect -2562 -460 -2528 -426
rect -2562 -528 -2528 -494
rect -2562 -596 -2528 -562
rect -2562 -664 -2528 -630
rect -1544 -188 -1510 -154
rect -1544 -256 -1510 -222
rect -1544 -324 -1510 -290
rect -1544 -392 -1510 -358
rect -1544 -460 -1510 -426
rect -1544 -528 -1510 -494
rect -1544 -596 -1510 -562
rect -1544 -664 -1510 -630
rect -526 -188 -492 -154
rect -526 -256 -492 -222
rect -526 -324 -492 -290
rect -526 -392 -492 -358
rect -526 -460 -492 -426
rect -526 -528 -492 -494
rect -526 -596 -492 -562
rect -526 -664 -492 -630
rect 492 -188 526 -154
rect 492 -256 526 -222
rect 492 -324 526 -290
rect 492 -392 526 -358
rect 492 -460 526 -426
rect 492 -528 526 -494
rect 492 -596 526 -562
rect 492 -664 526 -630
rect 1510 -188 1544 -154
rect 1510 -256 1544 -222
rect 1510 -324 1544 -290
rect 1510 -392 1544 -358
rect 1510 -460 1544 -426
rect 1510 -528 1544 -494
rect 1510 -596 1544 -562
rect 1510 -664 1544 -630
rect 2528 -188 2562 -154
rect 2528 -256 2562 -222
rect 2528 -324 2562 -290
rect 2528 -392 2562 -358
rect 2528 -460 2562 -426
rect 2528 -528 2562 -494
rect 2528 -596 2562 -562
rect 2528 -664 2562 -630
rect 3546 -188 3580 -154
rect 3546 -256 3580 -222
rect 3546 -324 3580 -290
rect 3546 -392 3580 -358
rect 3546 -460 3580 -426
rect 3546 -528 3580 -494
rect 3546 -596 3580 -562
rect 3546 -664 3580 -630
rect 4564 -188 4598 -154
rect 4564 -256 4598 -222
rect 4564 -324 4598 -290
rect 4564 -392 4598 -358
rect 4564 -460 4598 -426
rect 4564 -528 4598 -494
rect 4564 -596 4598 -562
rect 4564 -664 4598 -630
rect -4598 -1006 -4564 -972
rect -4598 -1074 -4564 -1040
rect -4598 -1142 -4564 -1108
rect -4598 -1210 -4564 -1176
rect -4598 -1278 -4564 -1244
rect -4598 -1346 -4564 -1312
rect -4598 -1414 -4564 -1380
rect -4598 -1482 -4564 -1448
rect -3580 -1006 -3546 -972
rect -3580 -1074 -3546 -1040
rect -3580 -1142 -3546 -1108
rect -3580 -1210 -3546 -1176
rect -3580 -1278 -3546 -1244
rect -3580 -1346 -3546 -1312
rect -3580 -1414 -3546 -1380
rect -3580 -1482 -3546 -1448
rect -2562 -1006 -2528 -972
rect -2562 -1074 -2528 -1040
rect -2562 -1142 -2528 -1108
rect -2562 -1210 -2528 -1176
rect -2562 -1278 -2528 -1244
rect -2562 -1346 -2528 -1312
rect -2562 -1414 -2528 -1380
rect -2562 -1482 -2528 -1448
rect -1544 -1006 -1510 -972
rect -1544 -1074 -1510 -1040
rect -1544 -1142 -1510 -1108
rect -1544 -1210 -1510 -1176
rect -1544 -1278 -1510 -1244
rect -1544 -1346 -1510 -1312
rect -1544 -1414 -1510 -1380
rect -1544 -1482 -1510 -1448
rect -526 -1006 -492 -972
rect -526 -1074 -492 -1040
rect -526 -1142 -492 -1108
rect -526 -1210 -492 -1176
rect -526 -1278 -492 -1244
rect -526 -1346 -492 -1312
rect -526 -1414 -492 -1380
rect -526 -1482 -492 -1448
rect 492 -1006 526 -972
rect 492 -1074 526 -1040
rect 492 -1142 526 -1108
rect 492 -1210 526 -1176
rect 492 -1278 526 -1244
rect 492 -1346 526 -1312
rect 492 -1414 526 -1380
rect 492 -1482 526 -1448
rect 1510 -1006 1544 -972
rect 1510 -1074 1544 -1040
rect 1510 -1142 1544 -1108
rect 1510 -1210 1544 -1176
rect 1510 -1278 1544 -1244
rect 1510 -1346 1544 -1312
rect 1510 -1414 1544 -1380
rect 1510 -1482 1544 -1448
rect 2528 -1006 2562 -972
rect 2528 -1074 2562 -1040
rect 2528 -1142 2562 -1108
rect 2528 -1210 2562 -1176
rect 2528 -1278 2562 -1244
rect 2528 -1346 2562 -1312
rect 2528 -1414 2562 -1380
rect 2528 -1482 2562 -1448
rect 3546 -1006 3580 -972
rect 3546 -1074 3580 -1040
rect 3546 -1142 3580 -1108
rect 3546 -1210 3580 -1176
rect 3546 -1278 3580 -1244
rect 3546 -1346 3580 -1312
rect 3546 -1414 3580 -1380
rect 3546 -1482 3580 -1448
rect 4564 -1006 4598 -972
rect 4564 -1074 4598 -1040
rect 4564 -1142 4598 -1108
rect 4564 -1210 4598 -1176
rect 4564 -1278 4598 -1244
rect 4564 -1346 4598 -1312
rect 4564 -1414 4598 -1380
rect 4564 -1482 4598 -1448
<< poly >>
rect -4366 1599 -3778 1615
rect -4366 1582 -4327 1599
rect -4552 1565 -4327 1582
rect -4293 1565 -4259 1599
rect -4225 1565 -4191 1599
rect -4157 1565 -4123 1599
rect -4089 1565 -4055 1599
rect -4021 1565 -3987 1599
rect -3953 1565 -3919 1599
rect -3885 1565 -3851 1599
rect -3817 1582 -3778 1599
rect -3348 1599 -2760 1615
rect -3348 1582 -3309 1599
rect -3817 1565 -3592 1582
rect -4552 1527 -3592 1565
rect -3534 1565 -3309 1582
rect -3275 1565 -3241 1599
rect -3207 1565 -3173 1599
rect -3139 1565 -3105 1599
rect -3071 1565 -3037 1599
rect -3003 1565 -2969 1599
rect -2935 1565 -2901 1599
rect -2867 1565 -2833 1599
rect -2799 1582 -2760 1599
rect -2330 1599 -1742 1615
rect -2330 1582 -2291 1599
rect -2799 1565 -2574 1582
rect -3534 1527 -2574 1565
rect -2516 1565 -2291 1582
rect -2257 1565 -2223 1599
rect -2189 1565 -2155 1599
rect -2121 1565 -2087 1599
rect -2053 1565 -2019 1599
rect -1985 1565 -1951 1599
rect -1917 1565 -1883 1599
rect -1849 1565 -1815 1599
rect -1781 1582 -1742 1599
rect -1312 1599 -724 1615
rect -1312 1582 -1273 1599
rect -1781 1565 -1556 1582
rect -2516 1527 -1556 1565
rect -1498 1565 -1273 1582
rect -1239 1565 -1205 1599
rect -1171 1565 -1137 1599
rect -1103 1565 -1069 1599
rect -1035 1565 -1001 1599
rect -967 1565 -933 1599
rect -899 1565 -865 1599
rect -831 1565 -797 1599
rect -763 1582 -724 1599
rect -294 1599 294 1615
rect -294 1582 -255 1599
rect -763 1565 -538 1582
rect -1498 1527 -538 1565
rect -480 1565 -255 1582
rect -221 1565 -187 1599
rect -153 1565 -119 1599
rect -85 1565 -51 1599
rect -17 1565 17 1599
rect 51 1565 85 1599
rect 119 1565 153 1599
rect 187 1565 221 1599
rect 255 1582 294 1599
rect 724 1599 1312 1615
rect 724 1582 763 1599
rect 255 1565 480 1582
rect -480 1527 480 1565
rect 538 1565 763 1582
rect 797 1565 831 1599
rect 865 1565 899 1599
rect 933 1565 967 1599
rect 1001 1565 1035 1599
rect 1069 1565 1103 1599
rect 1137 1565 1171 1599
rect 1205 1565 1239 1599
rect 1273 1582 1312 1599
rect 1742 1599 2330 1615
rect 1742 1582 1781 1599
rect 1273 1565 1498 1582
rect 538 1527 1498 1565
rect 1556 1565 1781 1582
rect 1815 1565 1849 1599
rect 1883 1565 1917 1599
rect 1951 1565 1985 1599
rect 2019 1565 2053 1599
rect 2087 1565 2121 1599
rect 2155 1565 2189 1599
rect 2223 1565 2257 1599
rect 2291 1582 2330 1599
rect 2760 1599 3348 1615
rect 2760 1582 2799 1599
rect 2291 1565 2516 1582
rect 1556 1527 2516 1565
rect 2574 1565 2799 1582
rect 2833 1565 2867 1599
rect 2901 1565 2935 1599
rect 2969 1565 3003 1599
rect 3037 1565 3071 1599
rect 3105 1565 3139 1599
rect 3173 1565 3207 1599
rect 3241 1565 3275 1599
rect 3309 1582 3348 1599
rect 3778 1599 4366 1615
rect 3778 1582 3817 1599
rect 3309 1565 3534 1582
rect 2574 1527 3534 1565
rect 3592 1565 3817 1582
rect 3851 1565 3885 1599
rect 3919 1565 3953 1599
rect 3987 1565 4021 1599
rect 4055 1565 4089 1599
rect 4123 1565 4157 1599
rect 4191 1565 4225 1599
rect 4259 1565 4293 1599
rect 4327 1582 4366 1599
rect 4327 1565 4552 1582
rect 3592 1527 4552 1565
rect -4552 889 -3592 927
rect -4552 872 -4327 889
rect -4366 855 -4327 872
rect -4293 855 -4259 889
rect -4225 855 -4191 889
rect -4157 855 -4123 889
rect -4089 855 -4055 889
rect -4021 855 -3987 889
rect -3953 855 -3919 889
rect -3885 855 -3851 889
rect -3817 872 -3592 889
rect -3534 889 -2574 927
rect -3534 872 -3309 889
rect -3817 855 -3778 872
rect -4366 839 -3778 855
rect -3348 855 -3309 872
rect -3275 855 -3241 889
rect -3207 855 -3173 889
rect -3139 855 -3105 889
rect -3071 855 -3037 889
rect -3003 855 -2969 889
rect -2935 855 -2901 889
rect -2867 855 -2833 889
rect -2799 872 -2574 889
rect -2516 889 -1556 927
rect -2516 872 -2291 889
rect -2799 855 -2760 872
rect -3348 839 -2760 855
rect -2330 855 -2291 872
rect -2257 855 -2223 889
rect -2189 855 -2155 889
rect -2121 855 -2087 889
rect -2053 855 -2019 889
rect -1985 855 -1951 889
rect -1917 855 -1883 889
rect -1849 855 -1815 889
rect -1781 872 -1556 889
rect -1498 889 -538 927
rect -1498 872 -1273 889
rect -1781 855 -1742 872
rect -2330 839 -1742 855
rect -1312 855 -1273 872
rect -1239 855 -1205 889
rect -1171 855 -1137 889
rect -1103 855 -1069 889
rect -1035 855 -1001 889
rect -967 855 -933 889
rect -899 855 -865 889
rect -831 855 -797 889
rect -763 872 -538 889
rect -480 889 480 927
rect -480 872 -255 889
rect -763 855 -724 872
rect -1312 839 -724 855
rect -294 855 -255 872
rect -221 855 -187 889
rect -153 855 -119 889
rect -85 855 -51 889
rect -17 855 17 889
rect 51 855 85 889
rect 119 855 153 889
rect 187 855 221 889
rect 255 872 480 889
rect 538 889 1498 927
rect 538 872 763 889
rect 255 855 294 872
rect -294 839 294 855
rect 724 855 763 872
rect 797 855 831 889
rect 865 855 899 889
rect 933 855 967 889
rect 1001 855 1035 889
rect 1069 855 1103 889
rect 1137 855 1171 889
rect 1205 855 1239 889
rect 1273 872 1498 889
rect 1556 889 2516 927
rect 1556 872 1781 889
rect 1273 855 1312 872
rect 724 839 1312 855
rect 1742 855 1781 872
rect 1815 855 1849 889
rect 1883 855 1917 889
rect 1951 855 1985 889
rect 2019 855 2053 889
rect 2087 855 2121 889
rect 2155 855 2189 889
rect 2223 855 2257 889
rect 2291 872 2516 889
rect 2574 889 3534 927
rect 2574 872 2799 889
rect 2291 855 2330 872
rect 1742 839 2330 855
rect 2760 855 2799 872
rect 2833 855 2867 889
rect 2901 855 2935 889
rect 2969 855 3003 889
rect 3037 855 3071 889
rect 3105 855 3139 889
rect 3173 855 3207 889
rect 3241 855 3275 889
rect 3309 872 3534 889
rect 3592 889 4552 927
rect 3592 872 3817 889
rect 3309 855 3348 872
rect 2760 839 3348 855
rect 3778 855 3817 872
rect 3851 855 3885 889
rect 3919 855 3953 889
rect 3987 855 4021 889
rect 4055 855 4089 889
rect 4123 855 4157 889
rect 4191 855 4225 889
rect 4259 855 4293 889
rect 4327 872 4552 889
rect 4327 855 4366 872
rect 3778 839 4366 855
rect -4366 781 -3778 797
rect -4366 764 -4327 781
rect -4552 747 -4327 764
rect -4293 747 -4259 781
rect -4225 747 -4191 781
rect -4157 747 -4123 781
rect -4089 747 -4055 781
rect -4021 747 -3987 781
rect -3953 747 -3919 781
rect -3885 747 -3851 781
rect -3817 764 -3778 781
rect -3348 781 -2760 797
rect -3348 764 -3309 781
rect -3817 747 -3592 764
rect -4552 709 -3592 747
rect -3534 747 -3309 764
rect -3275 747 -3241 781
rect -3207 747 -3173 781
rect -3139 747 -3105 781
rect -3071 747 -3037 781
rect -3003 747 -2969 781
rect -2935 747 -2901 781
rect -2867 747 -2833 781
rect -2799 764 -2760 781
rect -2330 781 -1742 797
rect -2330 764 -2291 781
rect -2799 747 -2574 764
rect -3534 709 -2574 747
rect -2516 747 -2291 764
rect -2257 747 -2223 781
rect -2189 747 -2155 781
rect -2121 747 -2087 781
rect -2053 747 -2019 781
rect -1985 747 -1951 781
rect -1917 747 -1883 781
rect -1849 747 -1815 781
rect -1781 764 -1742 781
rect -1312 781 -724 797
rect -1312 764 -1273 781
rect -1781 747 -1556 764
rect -2516 709 -1556 747
rect -1498 747 -1273 764
rect -1239 747 -1205 781
rect -1171 747 -1137 781
rect -1103 747 -1069 781
rect -1035 747 -1001 781
rect -967 747 -933 781
rect -899 747 -865 781
rect -831 747 -797 781
rect -763 764 -724 781
rect -294 781 294 797
rect -294 764 -255 781
rect -763 747 -538 764
rect -1498 709 -538 747
rect -480 747 -255 764
rect -221 747 -187 781
rect -153 747 -119 781
rect -85 747 -51 781
rect -17 747 17 781
rect 51 747 85 781
rect 119 747 153 781
rect 187 747 221 781
rect 255 764 294 781
rect 724 781 1312 797
rect 724 764 763 781
rect 255 747 480 764
rect -480 709 480 747
rect 538 747 763 764
rect 797 747 831 781
rect 865 747 899 781
rect 933 747 967 781
rect 1001 747 1035 781
rect 1069 747 1103 781
rect 1137 747 1171 781
rect 1205 747 1239 781
rect 1273 764 1312 781
rect 1742 781 2330 797
rect 1742 764 1781 781
rect 1273 747 1498 764
rect 538 709 1498 747
rect 1556 747 1781 764
rect 1815 747 1849 781
rect 1883 747 1917 781
rect 1951 747 1985 781
rect 2019 747 2053 781
rect 2087 747 2121 781
rect 2155 747 2189 781
rect 2223 747 2257 781
rect 2291 764 2330 781
rect 2760 781 3348 797
rect 2760 764 2799 781
rect 2291 747 2516 764
rect 1556 709 2516 747
rect 2574 747 2799 764
rect 2833 747 2867 781
rect 2901 747 2935 781
rect 2969 747 3003 781
rect 3037 747 3071 781
rect 3105 747 3139 781
rect 3173 747 3207 781
rect 3241 747 3275 781
rect 3309 764 3348 781
rect 3778 781 4366 797
rect 3778 764 3817 781
rect 3309 747 3534 764
rect 2574 709 3534 747
rect 3592 747 3817 764
rect 3851 747 3885 781
rect 3919 747 3953 781
rect 3987 747 4021 781
rect 4055 747 4089 781
rect 4123 747 4157 781
rect 4191 747 4225 781
rect 4259 747 4293 781
rect 4327 764 4366 781
rect 4327 747 4552 764
rect 3592 709 4552 747
rect -4552 71 -3592 109
rect -4552 54 -4327 71
rect -4366 37 -4327 54
rect -4293 37 -4259 71
rect -4225 37 -4191 71
rect -4157 37 -4123 71
rect -4089 37 -4055 71
rect -4021 37 -3987 71
rect -3953 37 -3919 71
rect -3885 37 -3851 71
rect -3817 54 -3592 71
rect -3534 71 -2574 109
rect -3534 54 -3309 71
rect -3817 37 -3778 54
rect -4366 21 -3778 37
rect -3348 37 -3309 54
rect -3275 37 -3241 71
rect -3207 37 -3173 71
rect -3139 37 -3105 71
rect -3071 37 -3037 71
rect -3003 37 -2969 71
rect -2935 37 -2901 71
rect -2867 37 -2833 71
rect -2799 54 -2574 71
rect -2516 71 -1556 109
rect -2516 54 -2291 71
rect -2799 37 -2760 54
rect -3348 21 -2760 37
rect -2330 37 -2291 54
rect -2257 37 -2223 71
rect -2189 37 -2155 71
rect -2121 37 -2087 71
rect -2053 37 -2019 71
rect -1985 37 -1951 71
rect -1917 37 -1883 71
rect -1849 37 -1815 71
rect -1781 54 -1556 71
rect -1498 71 -538 109
rect -1498 54 -1273 71
rect -1781 37 -1742 54
rect -2330 21 -1742 37
rect -1312 37 -1273 54
rect -1239 37 -1205 71
rect -1171 37 -1137 71
rect -1103 37 -1069 71
rect -1035 37 -1001 71
rect -967 37 -933 71
rect -899 37 -865 71
rect -831 37 -797 71
rect -763 54 -538 71
rect -480 71 480 109
rect -480 54 -255 71
rect -763 37 -724 54
rect -1312 21 -724 37
rect -294 37 -255 54
rect -221 37 -187 71
rect -153 37 -119 71
rect -85 37 -51 71
rect -17 37 17 71
rect 51 37 85 71
rect 119 37 153 71
rect 187 37 221 71
rect 255 54 480 71
rect 538 71 1498 109
rect 538 54 763 71
rect 255 37 294 54
rect -294 21 294 37
rect 724 37 763 54
rect 797 37 831 71
rect 865 37 899 71
rect 933 37 967 71
rect 1001 37 1035 71
rect 1069 37 1103 71
rect 1137 37 1171 71
rect 1205 37 1239 71
rect 1273 54 1498 71
rect 1556 71 2516 109
rect 1556 54 1781 71
rect 1273 37 1312 54
rect 724 21 1312 37
rect 1742 37 1781 54
rect 1815 37 1849 71
rect 1883 37 1917 71
rect 1951 37 1985 71
rect 2019 37 2053 71
rect 2087 37 2121 71
rect 2155 37 2189 71
rect 2223 37 2257 71
rect 2291 54 2516 71
rect 2574 71 3534 109
rect 2574 54 2799 71
rect 2291 37 2330 54
rect 1742 21 2330 37
rect 2760 37 2799 54
rect 2833 37 2867 71
rect 2901 37 2935 71
rect 2969 37 3003 71
rect 3037 37 3071 71
rect 3105 37 3139 71
rect 3173 37 3207 71
rect 3241 37 3275 71
rect 3309 54 3534 71
rect 3592 71 4552 109
rect 3592 54 3817 71
rect 3309 37 3348 54
rect 2760 21 3348 37
rect 3778 37 3817 54
rect 3851 37 3885 71
rect 3919 37 3953 71
rect 3987 37 4021 71
rect 4055 37 4089 71
rect 4123 37 4157 71
rect 4191 37 4225 71
rect 4259 37 4293 71
rect 4327 54 4552 71
rect 4327 37 4366 54
rect 3778 21 4366 37
rect -4366 -37 -3778 -21
rect -4366 -54 -4327 -37
rect -4552 -71 -4327 -54
rect -4293 -71 -4259 -37
rect -4225 -71 -4191 -37
rect -4157 -71 -4123 -37
rect -4089 -71 -4055 -37
rect -4021 -71 -3987 -37
rect -3953 -71 -3919 -37
rect -3885 -71 -3851 -37
rect -3817 -54 -3778 -37
rect -3348 -37 -2760 -21
rect -3348 -54 -3309 -37
rect -3817 -71 -3592 -54
rect -4552 -109 -3592 -71
rect -3534 -71 -3309 -54
rect -3275 -71 -3241 -37
rect -3207 -71 -3173 -37
rect -3139 -71 -3105 -37
rect -3071 -71 -3037 -37
rect -3003 -71 -2969 -37
rect -2935 -71 -2901 -37
rect -2867 -71 -2833 -37
rect -2799 -54 -2760 -37
rect -2330 -37 -1742 -21
rect -2330 -54 -2291 -37
rect -2799 -71 -2574 -54
rect -3534 -109 -2574 -71
rect -2516 -71 -2291 -54
rect -2257 -71 -2223 -37
rect -2189 -71 -2155 -37
rect -2121 -71 -2087 -37
rect -2053 -71 -2019 -37
rect -1985 -71 -1951 -37
rect -1917 -71 -1883 -37
rect -1849 -71 -1815 -37
rect -1781 -54 -1742 -37
rect -1312 -37 -724 -21
rect -1312 -54 -1273 -37
rect -1781 -71 -1556 -54
rect -2516 -109 -1556 -71
rect -1498 -71 -1273 -54
rect -1239 -71 -1205 -37
rect -1171 -71 -1137 -37
rect -1103 -71 -1069 -37
rect -1035 -71 -1001 -37
rect -967 -71 -933 -37
rect -899 -71 -865 -37
rect -831 -71 -797 -37
rect -763 -54 -724 -37
rect -294 -37 294 -21
rect -294 -54 -255 -37
rect -763 -71 -538 -54
rect -1498 -109 -538 -71
rect -480 -71 -255 -54
rect -221 -71 -187 -37
rect -153 -71 -119 -37
rect -85 -71 -51 -37
rect -17 -71 17 -37
rect 51 -71 85 -37
rect 119 -71 153 -37
rect 187 -71 221 -37
rect 255 -54 294 -37
rect 724 -37 1312 -21
rect 724 -54 763 -37
rect 255 -71 480 -54
rect -480 -109 480 -71
rect 538 -71 763 -54
rect 797 -71 831 -37
rect 865 -71 899 -37
rect 933 -71 967 -37
rect 1001 -71 1035 -37
rect 1069 -71 1103 -37
rect 1137 -71 1171 -37
rect 1205 -71 1239 -37
rect 1273 -54 1312 -37
rect 1742 -37 2330 -21
rect 1742 -54 1781 -37
rect 1273 -71 1498 -54
rect 538 -109 1498 -71
rect 1556 -71 1781 -54
rect 1815 -71 1849 -37
rect 1883 -71 1917 -37
rect 1951 -71 1985 -37
rect 2019 -71 2053 -37
rect 2087 -71 2121 -37
rect 2155 -71 2189 -37
rect 2223 -71 2257 -37
rect 2291 -54 2330 -37
rect 2760 -37 3348 -21
rect 2760 -54 2799 -37
rect 2291 -71 2516 -54
rect 1556 -109 2516 -71
rect 2574 -71 2799 -54
rect 2833 -71 2867 -37
rect 2901 -71 2935 -37
rect 2969 -71 3003 -37
rect 3037 -71 3071 -37
rect 3105 -71 3139 -37
rect 3173 -71 3207 -37
rect 3241 -71 3275 -37
rect 3309 -54 3348 -37
rect 3778 -37 4366 -21
rect 3778 -54 3817 -37
rect 3309 -71 3534 -54
rect 2574 -109 3534 -71
rect 3592 -71 3817 -54
rect 3851 -71 3885 -37
rect 3919 -71 3953 -37
rect 3987 -71 4021 -37
rect 4055 -71 4089 -37
rect 4123 -71 4157 -37
rect 4191 -71 4225 -37
rect 4259 -71 4293 -37
rect 4327 -54 4366 -37
rect 4327 -71 4552 -54
rect 3592 -109 4552 -71
rect -4552 -747 -3592 -709
rect -4552 -764 -4327 -747
rect -4366 -781 -4327 -764
rect -4293 -781 -4259 -747
rect -4225 -781 -4191 -747
rect -4157 -781 -4123 -747
rect -4089 -781 -4055 -747
rect -4021 -781 -3987 -747
rect -3953 -781 -3919 -747
rect -3885 -781 -3851 -747
rect -3817 -764 -3592 -747
rect -3534 -747 -2574 -709
rect -3534 -764 -3309 -747
rect -3817 -781 -3778 -764
rect -4366 -797 -3778 -781
rect -3348 -781 -3309 -764
rect -3275 -781 -3241 -747
rect -3207 -781 -3173 -747
rect -3139 -781 -3105 -747
rect -3071 -781 -3037 -747
rect -3003 -781 -2969 -747
rect -2935 -781 -2901 -747
rect -2867 -781 -2833 -747
rect -2799 -764 -2574 -747
rect -2516 -747 -1556 -709
rect -2516 -764 -2291 -747
rect -2799 -781 -2760 -764
rect -3348 -797 -2760 -781
rect -2330 -781 -2291 -764
rect -2257 -781 -2223 -747
rect -2189 -781 -2155 -747
rect -2121 -781 -2087 -747
rect -2053 -781 -2019 -747
rect -1985 -781 -1951 -747
rect -1917 -781 -1883 -747
rect -1849 -781 -1815 -747
rect -1781 -764 -1556 -747
rect -1498 -747 -538 -709
rect -1498 -764 -1273 -747
rect -1781 -781 -1742 -764
rect -2330 -797 -1742 -781
rect -1312 -781 -1273 -764
rect -1239 -781 -1205 -747
rect -1171 -781 -1137 -747
rect -1103 -781 -1069 -747
rect -1035 -781 -1001 -747
rect -967 -781 -933 -747
rect -899 -781 -865 -747
rect -831 -781 -797 -747
rect -763 -764 -538 -747
rect -480 -747 480 -709
rect -480 -764 -255 -747
rect -763 -781 -724 -764
rect -1312 -797 -724 -781
rect -294 -781 -255 -764
rect -221 -781 -187 -747
rect -153 -781 -119 -747
rect -85 -781 -51 -747
rect -17 -781 17 -747
rect 51 -781 85 -747
rect 119 -781 153 -747
rect 187 -781 221 -747
rect 255 -764 480 -747
rect 538 -747 1498 -709
rect 538 -764 763 -747
rect 255 -781 294 -764
rect -294 -797 294 -781
rect 724 -781 763 -764
rect 797 -781 831 -747
rect 865 -781 899 -747
rect 933 -781 967 -747
rect 1001 -781 1035 -747
rect 1069 -781 1103 -747
rect 1137 -781 1171 -747
rect 1205 -781 1239 -747
rect 1273 -764 1498 -747
rect 1556 -747 2516 -709
rect 1556 -764 1781 -747
rect 1273 -781 1312 -764
rect 724 -797 1312 -781
rect 1742 -781 1781 -764
rect 1815 -781 1849 -747
rect 1883 -781 1917 -747
rect 1951 -781 1985 -747
rect 2019 -781 2053 -747
rect 2087 -781 2121 -747
rect 2155 -781 2189 -747
rect 2223 -781 2257 -747
rect 2291 -764 2516 -747
rect 2574 -747 3534 -709
rect 2574 -764 2799 -747
rect 2291 -781 2330 -764
rect 1742 -797 2330 -781
rect 2760 -781 2799 -764
rect 2833 -781 2867 -747
rect 2901 -781 2935 -747
rect 2969 -781 3003 -747
rect 3037 -781 3071 -747
rect 3105 -781 3139 -747
rect 3173 -781 3207 -747
rect 3241 -781 3275 -747
rect 3309 -764 3534 -747
rect 3592 -747 4552 -709
rect 3592 -764 3817 -747
rect 3309 -781 3348 -764
rect 2760 -797 3348 -781
rect 3778 -781 3817 -764
rect 3851 -781 3885 -747
rect 3919 -781 3953 -747
rect 3987 -781 4021 -747
rect 4055 -781 4089 -747
rect 4123 -781 4157 -747
rect 4191 -781 4225 -747
rect 4259 -781 4293 -747
rect 4327 -764 4552 -747
rect 4327 -781 4366 -764
rect 3778 -797 4366 -781
rect -4366 -855 -3778 -839
rect -4366 -872 -4327 -855
rect -4552 -889 -4327 -872
rect -4293 -889 -4259 -855
rect -4225 -889 -4191 -855
rect -4157 -889 -4123 -855
rect -4089 -889 -4055 -855
rect -4021 -889 -3987 -855
rect -3953 -889 -3919 -855
rect -3885 -889 -3851 -855
rect -3817 -872 -3778 -855
rect -3348 -855 -2760 -839
rect -3348 -872 -3309 -855
rect -3817 -889 -3592 -872
rect -4552 -927 -3592 -889
rect -3534 -889 -3309 -872
rect -3275 -889 -3241 -855
rect -3207 -889 -3173 -855
rect -3139 -889 -3105 -855
rect -3071 -889 -3037 -855
rect -3003 -889 -2969 -855
rect -2935 -889 -2901 -855
rect -2867 -889 -2833 -855
rect -2799 -872 -2760 -855
rect -2330 -855 -1742 -839
rect -2330 -872 -2291 -855
rect -2799 -889 -2574 -872
rect -3534 -927 -2574 -889
rect -2516 -889 -2291 -872
rect -2257 -889 -2223 -855
rect -2189 -889 -2155 -855
rect -2121 -889 -2087 -855
rect -2053 -889 -2019 -855
rect -1985 -889 -1951 -855
rect -1917 -889 -1883 -855
rect -1849 -889 -1815 -855
rect -1781 -872 -1742 -855
rect -1312 -855 -724 -839
rect -1312 -872 -1273 -855
rect -1781 -889 -1556 -872
rect -2516 -927 -1556 -889
rect -1498 -889 -1273 -872
rect -1239 -889 -1205 -855
rect -1171 -889 -1137 -855
rect -1103 -889 -1069 -855
rect -1035 -889 -1001 -855
rect -967 -889 -933 -855
rect -899 -889 -865 -855
rect -831 -889 -797 -855
rect -763 -872 -724 -855
rect -294 -855 294 -839
rect -294 -872 -255 -855
rect -763 -889 -538 -872
rect -1498 -927 -538 -889
rect -480 -889 -255 -872
rect -221 -889 -187 -855
rect -153 -889 -119 -855
rect -85 -889 -51 -855
rect -17 -889 17 -855
rect 51 -889 85 -855
rect 119 -889 153 -855
rect 187 -889 221 -855
rect 255 -872 294 -855
rect 724 -855 1312 -839
rect 724 -872 763 -855
rect 255 -889 480 -872
rect -480 -927 480 -889
rect 538 -889 763 -872
rect 797 -889 831 -855
rect 865 -889 899 -855
rect 933 -889 967 -855
rect 1001 -889 1035 -855
rect 1069 -889 1103 -855
rect 1137 -889 1171 -855
rect 1205 -889 1239 -855
rect 1273 -872 1312 -855
rect 1742 -855 2330 -839
rect 1742 -872 1781 -855
rect 1273 -889 1498 -872
rect 538 -927 1498 -889
rect 1556 -889 1781 -872
rect 1815 -889 1849 -855
rect 1883 -889 1917 -855
rect 1951 -889 1985 -855
rect 2019 -889 2053 -855
rect 2087 -889 2121 -855
rect 2155 -889 2189 -855
rect 2223 -889 2257 -855
rect 2291 -872 2330 -855
rect 2760 -855 3348 -839
rect 2760 -872 2799 -855
rect 2291 -889 2516 -872
rect 1556 -927 2516 -889
rect 2574 -889 2799 -872
rect 2833 -889 2867 -855
rect 2901 -889 2935 -855
rect 2969 -889 3003 -855
rect 3037 -889 3071 -855
rect 3105 -889 3139 -855
rect 3173 -889 3207 -855
rect 3241 -889 3275 -855
rect 3309 -872 3348 -855
rect 3778 -855 4366 -839
rect 3778 -872 3817 -855
rect 3309 -889 3534 -872
rect 2574 -927 3534 -889
rect 3592 -889 3817 -872
rect 3851 -889 3885 -855
rect 3919 -889 3953 -855
rect 3987 -889 4021 -855
rect 4055 -889 4089 -855
rect 4123 -889 4157 -855
rect 4191 -889 4225 -855
rect 4259 -889 4293 -855
rect 4327 -872 4366 -855
rect 4327 -889 4552 -872
rect 3592 -927 4552 -889
rect -4552 -1565 -3592 -1527
rect -4552 -1582 -4327 -1565
rect -4366 -1599 -4327 -1582
rect -4293 -1599 -4259 -1565
rect -4225 -1599 -4191 -1565
rect -4157 -1599 -4123 -1565
rect -4089 -1599 -4055 -1565
rect -4021 -1599 -3987 -1565
rect -3953 -1599 -3919 -1565
rect -3885 -1599 -3851 -1565
rect -3817 -1582 -3592 -1565
rect -3534 -1565 -2574 -1527
rect -3534 -1582 -3309 -1565
rect -3817 -1599 -3778 -1582
rect -4366 -1615 -3778 -1599
rect -3348 -1599 -3309 -1582
rect -3275 -1599 -3241 -1565
rect -3207 -1599 -3173 -1565
rect -3139 -1599 -3105 -1565
rect -3071 -1599 -3037 -1565
rect -3003 -1599 -2969 -1565
rect -2935 -1599 -2901 -1565
rect -2867 -1599 -2833 -1565
rect -2799 -1582 -2574 -1565
rect -2516 -1565 -1556 -1527
rect -2516 -1582 -2291 -1565
rect -2799 -1599 -2760 -1582
rect -3348 -1615 -2760 -1599
rect -2330 -1599 -2291 -1582
rect -2257 -1599 -2223 -1565
rect -2189 -1599 -2155 -1565
rect -2121 -1599 -2087 -1565
rect -2053 -1599 -2019 -1565
rect -1985 -1599 -1951 -1565
rect -1917 -1599 -1883 -1565
rect -1849 -1599 -1815 -1565
rect -1781 -1582 -1556 -1565
rect -1498 -1565 -538 -1527
rect -1498 -1582 -1273 -1565
rect -1781 -1599 -1742 -1582
rect -2330 -1615 -1742 -1599
rect -1312 -1599 -1273 -1582
rect -1239 -1599 -1205 -1565
rect -1171 -1599 -1137 -1565
rect -1103 -1599 -1069 -1565
rect -1035 -1599 -1001 -1565
rect -967 -1599 -933 -1565
rect -899 -1599 -865 -1565
rect -831 -1599 -797 -1565
rect -763 -1582 -538 -1565
rect -480 -1565 480 -1527
rect -480 -1582 -255 -1565
rect -763 -1599 -724 -1582
rect -1312 -1615 -724 -1599
rect -294 -1599 -255 -1582
rect -221 -1599 -187 -1565
rect -153 -1599 -119 -1565
rect -85 -1599 -51 -1565
rect -17 -1599 17 -1565
rect 51 -1599 85 -1565
rect 119 -1599 153 -1565
rect 187 -1599 221 -1565
rect 255 -1582 480 -1565
rect 538 -1565 1498 -1527
rect 538 -1582 763 -1565
rect 255 -1599 294 -1582
rect -294 -1615 294 -1599
rect 724 -1599 763 -1582
rect 797 -1599 831 -1565
rect 865 -1599 899 -1565
rect 933 -1599 967 -1565
rect 1001 -1599 1035 -1565
rect 1069 -1599 1103 -1565
rect 1137 -1599 1171 -1565
rect 1205 -1599 1239 -1565
rect 1273 -1582 1498 -1565
rect 1556 -1565 2516 -1527
rect 1556 -1582 1781 -1565
rect 1273 -1599 1312 -1582
rect 724 -1615 1312 -1599
rect 1742 -1599 1781 -1582
rect 1815 -1599 1849 -1565
rect 1883 -1599 1917 -1565
rect 1951 -1599 1985 -1565
rect 2019 -1599 2053 -1565
rect 2087 -1599 2121 -1565
rect 2155 -1599 2189 -1565
rect 2223 -1599 2257 -1565
rect 2291 -1582 2516 -1565
rect 2574 -1565 3534 -1527
rect 2574 -1582 2799 -1565
rect 2291 -1599 2330 -1582
rect 1742 -1615 2330 -1599
rect 2760 -1599 2799 -1582
rect 2833 -1599 2867 -1565
rect 2901 -1599 2935 -1565
rect 2969 -1599 3003 -1565
rect 3037 -1599 3071 -1565
rect 3105 -1599 3139 -1565
rect 3173 -1599 3207 -1565
rect 3241 -1599 3275 -1565
rect 3309 -1582 3534 -1565
rect 3592 -1565 4552 -1527
rect 3592 -1582 3817 -1565
rect 3309 -1599 3348 -1582
rect 2760 -1615 3348 -1599
rect 3778 -1599 3817 -1582
rect 3851 -1599 3885 -1565
rect 3919 -1599 3953 -1565
rect 3987 -1599 4021 -1565
rect 4055 -1599 4089 -1565
rect 4123 -1599 4157 -1565
rect 4191 -1599 4225 -1565
rect 4259 -1599 4293 -1565
rect 4327 -1582 4552 -1565
rect 4327 -1599 4366 -1582
rect 3778 -1615 4366 -1599
<< polycont >>
rect -4327 1565 -4293 1599
rect -4259 1565 -4225 1599
rect -4191 1565 -4157 1599
rect -4123 1565 -4089 1599
rect -4055 1565 -4021 1599
rect -3987 1565 -3953 1599
rect -3919 1565 -3885 1599
rect -3851 1565 -3817 1599
rect -3309 1565 -3275 1599
rect -3241 1565 -3207 1599
rect -3173 1565 -3139 1599
rect -3105 1565 -3071 1599
rect -3037 1565 -3003 1599
rect -2969 1565 -2935 1599
rect -2901 1565 -2867 1599
rect -2833 1565 -2799 1599
rect -2291 1565 -2257 1599
rect -2223 1565 -2189 1599
rect -2155 1565 -2121 1599
rect -2087 1565 -2053 1599
rect -2019 1565 -1985 1599
rect -1951 1565 -1917 1599
rect -1883 1565 -1849 1599
rect -1815 1565 -1781 1599
rect -1273 1565 -1239 1599
rect -1205 1565 -1171 1599
rect -1137 1565 -1103 1599
rect -1069 1565 -1035 1599
rect -1001 1565 -967 1599
rect -933 1565 -899 1599
rect -865 1565 -831 1599
rect -797 1565 -763 1599
rect -255 1565 -221 1599
rect -187 1565 -153 1599
rect -119 1565 -85 1599
rect -51 1565 -17 1599
rect 17 1565 51 1599
rect 85 1565 119 1599
rect 153 1565 187 1599
rect 221 1565 255 1599
rect 763 1565 797 1599
rect 831 1565 865 1599
rect 899 1565 933 1599
rect 967 1565 1001 1599
rect 1035 1565 1069 1599
rect 1103 1565 1137 1599
rect 1171 1565 1205 1599
rect 1239 1565 1273 1599
rect 1781 1565 1815 1599
rect 1849 1565 1883 1599
rect 1917 1565 1951 1599
rect 1985 1565 2019 1599
rect 2053 1565 2087 1599
rect 2121 1565 2155 1599
rect 2189 1565 2223 1599
rect 2257 1565 2291 1599
rect 2799 1565 2833 1599
rect 2867 1565 2901 1599
rect 2935 1565 2969 1599
rect 3003 1565 3037 1599
rect 3071 1565 3105 1599
rect 3139 1565 3173 1599
rect 3207 1565 3241 1599
rect 3275 1565 3309 1599
rect 3817 1565 3851 1599
rect 3885 1565 3919 1599
rect 3953 1565 3987 1599
rect 4021 1565 4055 1599
rect 4089 1565 4123 1599
rect 4157 1565 4191 1599
rect 4225 1565 4259 1599
rect 4293 1565 4327 1599
rect -4327 855 -4293 889
rect -4259 855 -4225 889
rect -4191 855 -4157 889
rect -4123 855 -4089 889
rect -4055 855 -4021 889
rect -3987 855 -3953 889
rect -3919 855 -3885 889
rect -3851 855 -3817 889
rect -3309 855 -3275 889
rect -3241 855 -3207 889
rect -3173 855 -3139 889
rect -3105 855 -3071 889
rect -3037 855 -3003 889
rect -2969 855 -2935 889
rect -2901 855 -2867 889
rect -2833 855 -2799 889
rect -2291 855 -2257 889
rect -2223 855 -2189 889
rect -2155 855 -2121 889
rect -2087 855 -2053 889
rect -2019 855 -1985 889
rect -1951 855 -1917 889
rect -1883 855 -1849 889
rect -1815 855 -1781 889
rect -1273 855 -1239 889
rect -1205 855 -1171 889
rect -1137 855 -1103 889
rect -1069 855 -1035 889
rect -1001 855 -967 889
rect -933 855 -899 889
rect -865 855 -831 889
rect -797 855 -763 889
rect -255 855 -221 889
rect -187 855 -153 889
rect -119 855 -85 889
rect -51 855 -17 889
rect 17 855 51 889
rect 85 855 119 889
rect 153 855 187 889
rect 221 855 255 889
rect 763 855 797 889
rect 831 855 865 889
rect 899 855 933 889
rect 967 855 1001 889
rect 1035 855 1069 889
rect 1103 855 1137 889
rect 1171 855 1205 889
rect 1239 855 1273 889
rect 1781 855 1815 889
rect 1849 855 1883 889
rect 1917 855 1951 889
rect 1985 855 2019 889
rect 2053 855 2087 889
rect 2121 855 2155 889
rect 2189 855 2223 889
rect 2257 855 2291 889
rect 2799 855 2833 889
rect 2867 855 2901 889
rect 2935 855 2969 889
rect 3003 855 3037 889
rect 3071 855 3105 889
rect 3139 855 3173 889
rect 3207 855 3241 889
rect 3275 855 3309 889
rect 3817 855 3851 889
rect 3885 855 3919 889
rect 3953 855 3987 889
rect 4021 855 4055 889
rect 4089 855 4123 889
rect 4157 855 4191 889
rect 4225 855 4259 889
rect 4293 855 4327 889
rect -4327 747 -4293 781
rect -4259 747 -4225 781
rect -4191 747 -4157 781
rect -4123 747 -4089 781
rect -4055 747 -4021 781
rect -3987 747 -3953 781
rect -3919 747 -3885 781
rect -3851 747 -3817 781
rect -3309 747 -3275 781
rect -3241 747 -3207 781
rect -3173 747 -3139 781
rect -3105 747 -3071 781
rect -3037 747 -3003 781
rect -2969 747 -2935 781
rect -2901 747 -2867 781
rect -2833 747 -2799 781
rect -2291 747 -2257 781
rect -2223 747 -2189 781
rect -2155 747 -2121 781
rect -2087 747 -2053 781
rect -2019 747 -1985 781
rect -1951 747 -1917 781
rect -1883 747 -1849 781
rect -1815 747 -1781 781
rect -1273 747 -1239 781
rect -1205 747 -1171 781
rect -1137 747 -1103 781
rect -1069 747 -1035 781
rect -1001 747 -967 781
rect -933 747 -899 781
rect -865 747 -831 781
rect -797 747 -763 781
rect -255 747 -221 781
rect -187 747 -153 781
rect -119 747 -85 781
rect -51 747 -17 781
rect 17 747 51 781
rect 85 747 119 781
rect 153 747 187 781
rect 221 747 255 781
rect 763 747 797 781
rect 831 747 865 781
rect 899 747 933 781
rect 967 747 1001 781
rect 1035 747 1069 781
rect 1103 747 1137 781
rect 1171 747 1205 781
rect 1239 747 1273 781
rect 1781 747 1815 781
rect 1849 747 1883 781
rect 1917 747 1951 781
rect 1985 747 2019 781
rect 2053 747 2087 781
rect 2121 747 2155 781
rect 2189 747 2223 781
rect 2257 747 2291 781
rect 2799 747 2833 781
rect 2867 747 2901 781
rect 2935 747 2969 781
rect 3003 747 3037 781
rect 3071 747 3105 781
rect 3139 747 3173 781
rect 3207 747 3241 781
rect 3275 747 3309 781
rect 3817 747 3851 781
rect 3885 747 3919 781
rect 3953 747 3987 781
rect 4021 747 4055 781
rect 4089 747 4123 781
rect 4157 747 4191 781
rect 4225 747 4259 781
rect 4293 747 4327 781
rect -4327 37 -4293 71
rect -4259 37 -4225 71
rect -4191 37 -4157 71
rect -4123 37 -4089 71
rect -4055 37 -4021 71
rect -3987 37 -3953 71
rect -3919 37 -3885 71
rect -3851 37 -3817 71
rect -3309 37 -3275 71
rect -3241 37 -3207 71
rect -3173 37 -3139 71
rect -3105 37 -3071 71
rect -3037 37 -3003 71
rect -2969 37 -2935 71
rect -2901 37 -2867 71
rect -2833 37 -2799 71
rect -2291 37 -2257 71
rect -2223 37 -2189 71
rect -2155 37 -2121 71
rect -2087 37 -2053 71
rect -2019 37 -1985 71
rect -1951 37 -1917 71
rect -1883 37 -1849 71
rect -1815 37 -1781 71
rect -1273 37 -1239 71
rect -1205 37 -1171 71
rect -1137 37 -1103 71
rect -1069 37 -1035 71
rect -1001 37 -967 71
rect -933 37 -899 71
rect -865 37 -831 71
rect -797 37 -763 71
rect -255 37 -221 71
rect -187 37 -153 71
rect -119 37 -85 71
rect -51 37 -17 71
rect 17 37 51 71
rect 85 37 119 71
rect 153 37 187 71
rect 221 37 255 71
rect 763 37 797 71
rect 831 37 865 71
rect 899 37 933 71
rect 967 37 1001 71
rect 1035 37 1069 71
rect 1103 37 1137 71
rect 1171 37 1205 71
rect 1239 37 1273 71
rect 1781 37 1815 71
rect 1849 37 1883 71
rect 1917 37 1951 71
rect 1985 37 2019 71
rect 2053 37 2087 71
rect 2121 37 2155 71
rect 2189 37 2223 71
rect 2257 37 2291 71
rect 2799 37 2833 71
rect 2867 37 2901 71
rect 2935 37 2969 71
rect 3003 37 3037 71
rect 3071 37 3105 71
rect 3139 37 3173 71
rect 3207 37 3241 71
rect 3275 37 3309 71
rect 3817 37 3851 71
rect 3885 37 3919 71
rect 3953 37 3987 71
rect 4021 37 4055 71
rect 4089 37 4123 71
rect 4157 37 4191 71
rect 4225 37 4259 71
rect 4293 37 4327 71
rect -4327 -71 -4293 -37
rect -4259 -71 -4225 -37
rect -4191 -71 -4157 -37
rect -4123 -71 -4089 -37
rect -4055 -71 -4021 -37
rect -3987 -71 -3953 -37
rect -3919 -71 -3885 -37
rect -3851 -71 -3817 -37
rect -3309 -71 -3275 -37
rect -3241 -71 -3207 -37
rect -3173 -71 -3139 -37
rect -3105 -71 -3071 -37
rect -3037 -71 -3003 -37
rect -2969 -71 -2935 -37
rect -2901 -71 -2867 -37
rect -2833 -71 -2799 -37
rect -2291 -71 -2257 -37
rect -2223 -71 -2189 -37
rect -2155 -71 -2121 -37
rect -2087 -71 -2053 -37
rect -2019 -71 -1985 -37
rect -1951 -71 -1917 -37
rect -1883 -71 -1849 -37
rect -1815 -71 -1781 -37
rect -1273 -71 -1239 -37
rect -1205 -71 -1171 -37
rect -1137 -71 -1103 -37
rect -1069 -71 -1035 -37
rect -1001 -71 -967 -37
rect -933 -71 -899 -37
rect -865 -71 -831 -37
rect -797 -71 -763 -37
rect -255 -71 -221 -37
rect -187 -71 -153 -37
rect -119 -71 -85 -37
rect -51 -71 -17 -37
rect 17 -71 51 -37
rect 85 -71 119 -37
rect 153 -71 187 -37
rect 221 -71 255 -37
rect 763 -71 797 -37
rect 831 -71 865 -37
rect 899 -71 933 -37
rect 967 -71 1001 -37
rect 1035 -71 1069 -37
rect 1103 -71 1137 -37
rect 1171 -71 1205 -37
rect 1239 -71 1273 -37
rect 1781 -71 1815 -37
rect 1849 -71 1883 -37
rect 1917 -71 1951 -37
rect 1985 -71 2019 -37
rect 2053 -71 2087 -37
rect 2121 -71 2155 -37
rect 2189 -71 2223 -37
rect 2257 -71 2291 -37
rect 2799 -71 2833 -37
rect 2867 -71 2901 -37
rect 2935 -71 2969 -37
rect 3003 -71 3037 -37
rect 3071 -71 3105 -37
rect 3139 -71 3173 -37
rect 3207 -71 3241 -37
rect 3275 -71 3309 -37
rect 3817 -71 3851 -37
rect 3885 -71 3919 -37
rect 3953 -71 3987 -37
rect 4021 -71 4055 -37
rect 4089 -71 4123 -37
rect 4157 -71 4191 -37
rect 4225 -71 4259 -37
rect 4293 -71 4327 -37
rect -4327 -781 -4293 -747
rect -4259 -781 -4225 -747
rect -4191 -781 -4157 -747
rect -4123 -781 -4089 -747
rect -4055 -781 -4021 -747
rect -3987 -781 -3953 -747
rect -3919 -781 -3885 -747
rect -3851 -781 -3817 -747
rect -3309 -781 -3275 -747
rect -3241 -781 -3207 -747
rect -3173 -781 -3139 -747
rect -3105 -781 -3071 -747
rect -3037 -781 -3003 -747
rect -2969 -781 -2935 -747
rect -2901 -781 -2867 -747
rect -2833 -781 -2799 -747
rect -2291 -781 -2257 -747
rect -2223 -781 -2189 -747
rect -2155 -781 -2121 -747
rect -2087 -781 -2053 -747
rect -2019 -781 -1985 -747
rect -1951 -781 -1917 -747
rect -1883 -781 -1849 -747
rect -1815 -781 -1781 -747
rect -1273 -781 -1239 -747
rect -1205 -781 -1171 -747
rect -1137 -781 -1103 -747
rect -1069 -781 -1035 -747
rect -1001 -781 -967 -747
rect -933 -781 -899 -747
rect -865 -781 -831 -747
rect -797 -781 -763 -747
rect -255 -781 -221 -747
rect -187 -781 -153 -747
rect -119 -781 -85 -747
rect -51 -781 -17 -747
rect 17 -781 51 -747
rect 85 -781 119 -747
rect 153 -781 187 -747
rect 221 -781 255 -747
rect 763 -781 797 -747
rect 831 -781 865 -747
rect 899 -781 933 -747
rect 967 -781 1001 -747
rect 1035 -781 1069 -747
rect 1103 -781 1137 -747
rect 1171 -781 1205 -747
rect 1239 -781 1273 -747
rect 1781 -781 1815 -747
rect 1849 -781 1883 -747
rect 1917 -781 1951 -747
rect 1985 -781 2019 -747
rect 2053 -781 2087 -747
rect 2121 -781 2155 -747
rect 2189 -781 2223 -747
rect 2257 -781 2291 -747
rect 2799 -781 2833 -747
rect 2867 -781 2901 -747
rect 2935 -781 2969 -747
rect 3003 -781 3037 -747
rect 3071 -781 3105 -747
rect 3139 -781 3173 -747
rect 3207 -781 3241 -747
rect 3275 -781 3309 -747
rect 3817 -781 3851 -747
rect 3885 -781 3919 -747
rect 3953 -781 3987 -747
rect 4021 -781 4055 -747
rect 4089 -781 4123 -747
rect 4157 -781 4191 -747
rect 4225 -781 4259 -747
rect 4293 -781 4327 -747
rect -4327 -889 -4293 -855
rect -4259 -889 -4225 -855
rect -4191 -889 -4157 -855
rect -4123 -889 -4089 -855
rect -4055 -889 -4021 -855
rect -3987 -889 -3953 -855
rect -3919 -889 -3885 -855
rect -3851 -889 -3817 -855
rect -3309 -889 -3275 -855
rect -3241 -889 -3207 -855
rect -3173 -889 -3139 -855
rect -3105 -889 -3071 -855
rect -3037 -889 -3003 -855
rect -2969 -889 -2935 -855
rect -2901 -889 -2867 -855
rect -2833 -889 -2799 -855
rect -2291 -889 -2257 -855
rect -2223 -889 -2189 -855
rect -2155 -889 -2121 -855
rect -2087 -889 -2053 -855
rect -2019 -889 -1985 -855
rect -1951 -889 -1917 -855
rect -1883 -889 -1849 -855
rect -1815 -889 -1781 -855
rect -1273 -889 -1239 -855
rect -1205 -889 -1171 -855
rect -1137 -889 -1103 -855
rect -1069 -889 -1035 -855
rect -1001 -889 -967 -855
rect -933 -889 -899 -855
rect -865 -889 -831 -855
rect -797 -889 -763 -855
rect -255 -889 -221 -855
rect -187 -889 -153 -855
rect -119 -889 -85 -855
rect -51 -889 -17 -855
rect 17 -889 51 -855
rect 85 -889 119 -855
rect 153 -889 187 -855
rect 221 -889 255 -855
rect 763 -889 797 -855
rect 831 -889 865 -855
rect 899 -889 933 -855
rect 967 -889 1001 -855
rect 1035 -889 1069 -855
rect 1103 -889 1137 -855
rect 1171 -889 1205 -855
rect 1239 -889 1273 -855
rect 1781 -889 1815 -855
rect 1849 -889 1883 -855
rect 1917 -889 1951 -855
rect 1985 -889 2019 -855
rect 2053 -889 2087 -855
rect 2121 -889 2155 -855
rect 2189 -889 2223 -855
rect 2257 -889 2291 -855
rect 2799 -889 2833 -855
rect 2867 -889 2901 -855
rect 2935 -889 2969 -855
rect 3003 -889 3037 -855
rect 3071 -889 3105 -855
rect 3139 -889 3173 -855
rect 3207 -889 3241 -855
rect 3275 -889 3309 -855
rect 3817 -889 3851 -855
rect 3885 -889 3919 -855
rect 3953 -889 3987 -855
rect 4021 -889 4055 -855
rect 4089 -889 4123 -855
rect 4157 -889 4191 -855
rect 4225 -889 4259 -855
rect 4293 -889 4327 -855
rect -4327 -1599 -4293 -1565
rect -4259 -1599 -4225 -1565
rect -4191 -1599 -4157 -1565
rect -4123 -1599 -4089 -1565
rect -4055 -1599 -4021 -1565
rect -3987 -1599 -3953 -1565
rect -3919 -1599 -3885 -1565
rect -3851 -1599 -3817 -1565
rect -3309 -1599 -3275 -1565
rect -3241 -1599 -3207 -1565
rect -3173 -1599 -3139 -1565
rect -3105 -1599 -3071 -1565
rect -3037 -1599 -3003 -1565
rect -2969 -1599 -2935 -1565
rect -2901 -1599 -2867 -1565
rect -2833 -1599 -2799 -1565
rect -2291 -1599 -2257 -1565
rect -2223 -1599 -2189 -1565
rect -2155 -1599 -2121 -1565
rect -2087 -1599 -2053 -1565
rect -2019 -1599 -1985 -1565
rect -1951 -1599 -1917 -1565
rect -1883 -1599 -1849 -1565
rect -1815 -1599 -1781 -1565
rect -1273 -1599 -1239 -1565
rect -1205 -1599 -1171 -1565
rect -1137 -1599 -1103 -1565
rect -1069 -1599 -1035 -1565
rect -1001 -1599 -967 -1565
rect -933 -1599 -899 -1565
rect -865 -1599 -831 -1565
rect -797 -1599 -763 -1565
rect -255 -1599 -221 -1565
rect -187 -1599 -153 -1565
rect -119 -1599 -85 -1565
rect -51 -1599 -17 -1565
rect 17 -1599 51 -1565
rect 85 -1599 119 -1565
rect 153 -1599 187 -1565
rect 221 -1599 255 -1565
rect 763 -1599 797 -1565
rect 831 -1599 865 -1565
rect 899 -1599 933 -1565
rect 967 -1599 1001 -1565
rect 1035 -1599 1069 -1565
rect 1103 -1599 1137 -1565
rect 1171 -1599 1205 -1565
rect 1239 -1599 1273 -1565
rect 1781 -1599 1815 -1565
rect 1849 -1599 1883 -1565
rect 1917 -1599 1951 -1565
rect 1985 -1599 2019 -1565
rect 2053 -1599 2087 -1565
rect 2121 -1599 2155 -1565
rect 2189 -1599 2223 -1565
rect 2257 -1599 2291 -1565
rect 2799 -1599 2833 -1565
rect 2867 -1599 2901 -1565
rect 2935 -1599 2969 -1565
rect 3003 -1599 3037 -1565
rect 3071 -1599 3105 -1565
rect 3139 -1599 3173 -1565
rect 3207 -1599 3241 -1565
rect 3275 -1599 3309 -1565
rect 3817 -1599 3851 -1565
rect 3885 -1599 3919 -1565
rect 3953 -1599 3987 -1565
rect 4021 -1599 4055 -1565
rect 4089 -1599 4123 -1565
rect 4157 -1599 4191 -1565
rect 4225 -1599 4259 -1565
rect 4293 -1599 4327 -1565
<< locali >>
rect -4366 1565 -4327 1599
rect -4293 1565 -4269 1599
rect -4225 1565 -4197 1599
rect -4157 1565 -4125 1599
rect -4089 1565 -4055 1599
rect -4019 1565 -3987 1599
rect -3947 1565 -3919 1599
rect -3875 1565 -3851 1599
rect -3817 1565 -3778 1599
rect -3348 1565 -3309 1599
rect -3275 1565 -3251 1599
rect -3207 1565 -3179 1599
rect -3139 1565 -3107 1599
rect -3071 1565 -3037 1599
rect -3001 1565 -2969 1599
rect -2929 1565 -2901 1599
rect -2857 1565 -2833 1599
rect -2799 1565 -2760 1599
rect -2330 1565 -2291 1599
rect -2257 1565 -2233 1599
rect -2189 1565 -2161 1599
rect -2121 1565 -2089 1599
rect -2053 1565 -2019 1599
rect -1983 1565 -1951 1599
rect -1911 1565 -1883 1599
rect -1839 1565 -1815 1599
rect -1781 1565 -1742 1599
rect -1312 1565 -1273 1599
rect -1239 1565 -1215 1599
rect -1171 1565 -1143 1599
rect -1103 1565 -1071 1599
rect -1035 1565 -1001 1599
rect -965 1565 -933 1599
rect -893 1565 -865 1599
rect -821 1565 -797 1599
rect -763 1565 -724 1599
rect -294 1565 -255 1599
rect -221 1565 -197 1599
rect -153 1565 -125 1599
rect -85 1565 -53 1599
rect -17 1565 17 1599
rect 53 1565 85 1599
rect 125 1565 153 1599
rect 197 1565 221 1599
rect 255 1565 294 1599
rect 724 1565 763 1599
rect 797 1565 821 1599
rect 865 1565 893 1599
rect 933 1565 965 1599
rect 1001 1565 1035 1599
rect 1071 1565 1103 1599
rect 1143 1565 1171 1599
rect 1215 1565 1239 1599
rect 1273 1565 1312 1599
rect 1742 1565 1781 1599
rect 1815 1565 1839 1599
rect 1883 1565 1911 1599
rect 1951 1565 1983 1599
rect 2019 1565 2053 1599
rect 2089 1565 2121 1599
rect 2161 1565 2189 1599
rect 2233 1565 2257 1599
rect 2291 1565 2330 1599
rect 2760 1565 2799 1599
rect 2833 1565 2857 1599
rect 2901 1565 2929 1599
rect 2969 1565 3001 1599
rect 3037 1565 3071 1599
rect 3107 1565 3139 1599
rect 3179 1565 3207 1599
rect 3251 1565 3275 1599
rect 3309 1565 3348 1599
rect 3778 1565 3817 1599
rect 3851 1565 3875 1599
rect 3919 1565 3947 1599
rect 3987 1565 4019 1599
rect 4055 1565 4089 1599
rect 4125 1565 4157 1599
rect 4197 1565 4225 1599
rect 4269 1565 4293 1599
rect 4327 1565 4366 1599
rect -4598 1496 -4564 1531
rect -4598 1424 -4564 1448
rect -4598 1352 -4564 1380
rect -4598 1280 -4564 1312
rect -4598 1210 -4564 1244
rect -4598 1142 -4564 1174
rect -4598 1074 -4564 1102
rect -4598 1006 -4564 1030
rect -4598 923 -4564 958
rect -3580 1496 -3546 1531
rect -3580 1424 -3546 1448
rect -3580 1352 -3546 1380
rect -3580 1280 -3546 1312
rect -3580 1210 -3546 1244
rect -3580 1142 -3546 1174
rect -3580 1074 -3546 1102
rect -3580 1006 -3546 1030
rect -3580 923 -3546 958
rect -2562 1496 -2528 1531
rect -2562 1424 -2528 1448
rect -2562 1352 -2528 1380
rect -2562 1280 -2528 1312
rect -2562 1210 -2528 1244
rect -2562 1142 -2528 1174
rect -2562 1074 -2528 1102
rect -2562 1006 -2528 1030
rect -2562 923 -2528 958
rect -1544 1496 -1510 1531
rect -1544 1424 -1510 1448
rect -1544 1352 -1510 1380
rect -1544 1280 -1510 1312
rect -1544 1210 -1510 1244
rect -1544 1142 -1510 1174
rect -1544 1074 -1510 1102
rect -1544 1006 -1510 1030
rect -1544 923 -1510 958
rect -526 1496 -492 1531
rect -526 1424 -492 1448
rect -526 1352 -492 1380
rect -526 1280 -492 1312
rect -526 1210 -492 1244
rect -526 1142 -492 1174
rect -526 1074 -492 1102
rect -526 1006 -492 1030
rect -526 923 -492 958
rect 492 1496 526 1531
rect 492 1424 526 1448
rect 492 1352 526 1380
rect 492 1280 526 1312
rect 492 1210 526 1244
rect 492 1142 526 1174
rect 492 1074 526 1102
rect 492 1006 526 1030
rect 492 923 526 958
rect 1510 1496 1544 1531
rect 1510 1424 1544 1448
rect 1510 1352 1544 1380
rect 1510 1280 1544 1312
rect 1510 1210 1544 1244
rect 1510 1142 1544 1174
rect 1510 1074 1544 1102
rect 1510 1006 1544 1030
rect 1510 923 1544 958
rect 2528 1496 2562 1531
rect 2528 1424 2562 1448
rect 2528 1352 2562 1380
rect 2528 1280 2562 1312
rect 2528 1210 2562 1244
rect 2528 1142 2562 1174
rect 2528 1074 2562 1102
rect 2528 1006 2562 1030
rect 2528 923 2562 958
rect 3546 1496 3580 1531
rect 3546 1424 3580 1448
rect 3546 1352 3580 1380
rect 3546 1280 3580 1312
rect 3546 1210 3580 1244
rect 3546 1142 3580 1174
rect 3546 1074 3580 1102
rect 3546 1006 3580 1030
rect 3546 923 3580 958
rect 4564 1496 4598 1531
rect 4564 1424 4598 1448
rect 4564 1352 4598 1380
rect 4564 1280 4598 1312
rect 4564 1210 4598 1244
rect 4564 1142 4598 1174
rect 4564 1074 4598 1102
rect 4564 1006 4598 1030
rect 4564 923 4598 958
rect -4366 855 -4327 889
rect -4293 855 -4269 889
rect -4225 855 -4197 889
rect -4157 855 -4125 889
rect -4089 855 -4055 889
rect -4019 855 -3987 889
rect -3947 855 -3919 889
rect -3875 855 -3851 889
rect -3817 855 -3778 889
rect -3348 855 -3309 889
rect -3275 855 -3251 889
rect -3207 855 -3179 889
rect -3139 855 -3107 889
rect -3071 855 -3037 889
rect -3001 855 -2969 889
rect -2929 855 -2901 889
rect -2857 855 -2833 889
rect -2799 855 -2760 889
rect -2330 855 -2291 889
rect -2257 855 -2233 889
rect -2189 855 -2161 889
rect -2121 855 -2089 889
rect -2053 855 -2019 889
rect -1983 855 -1951 889
rect -1911 855 -1883 889
rect -1839 855 -1815 889
rect -1781 855 -1742 889
rect -1312 855 -1273 889
rect -1239 855 -1215 889
rect -1171 855 -1143 889
rect -1103 855 -1071 889
rect -1035 855 -1001 889
rect -965 855 -933 889
rect -893 855 -865 889
rect -821 855 -797 889
rect -763 855 -724 889
rect -294 855 -255 889
rect -221 855 -197 889
rect -153 855 -125 889
rect -85 855 -53 889
rect -17 855 17 889
rect 53 855 85 889
rect 125 855 153 889
rect 197 855 221 889
rect 255 855 294 889
rect 724 855 763 889
rect 797 855 821 889
rect 865 855 893 889
rect 933 855 965 889
rect 1001 855 1035 889
rect 1071 855 1103 889
rect 1143 855 1171 889
rect 1215 855 1239 889
rect 1273 855 1312 889
rect 1742 855 1781 889
rect 1815 855 1839 889
rect 1883 855 1911 889
rect 1951 855 1983 889
rect 2019 855 2053 889
rect 2089 855 2121 889
rect 2161 855 2189 889
rect 2233 855 2257 889
rect 2291 855 2330 889
rect 2760 855 2799 889
rect 2833 855 2857 889
rect 2901 855 2929 889
rect 2969 855 3001 889
rect 3037 855 3071 889
rect 3107 855 3139 889
rect 3179 855 3207 889
rect 3251 855 3275 889
rect 3309 855 3348 889
rect 3778 855 3817 889
rect 3851 855 3875 889
rect 3919 855 3947 889
rect 3987 855 4019 889
rect 4055 855 4089 889
rect 4125 855 4157 889
rect 4197 855 4225 889
rect 4269 855 4293 889
rect 4327 855 4366 889
rect -4366 747 -4327 781
rect -4293 747 -4269 781
rect -4225 747 -4197 781
rect -4157 747 -4125 781
rect -4089 747 -4055 781
rect -4019 747 -3987 781
rect -3947 747 -3919 781
rect -3875 747 -3851 781
rect -3817 747 -3778 781
rect -3348 747 -3309 781
rect -3275 747 -3251 781
rect -3207 747 -3179 781
rect -3139 747 -3107 781
rect -3071 747 -3037 781
rect -3001 747 -2969 781
rect -2929 747 -2901 781
rect -2857 747 -2833 781
rect -2799 747 -2760 781
rect -2330 747 -2291 781
rect -2257 747 -2233 781
rect -2189 747 -2161 781
rect -2121 747 -2089 781
rect -2053 747 -2019 781
rect -1983 747 -1951 781
rect -1911 747 -1883 781
rect -1839 747 -1815 781
rect -1781 747 -1742 781
rect -1312 747 -1273 781
rect -1239 747 -1215 781
rect -1171 747 -1143 781
rect -1103 747 -1071 781
rect -1035 747 -1001 781
rect -965 747 -933 781
rect -893 747 -865 781
rect -821 747 -797 781
rect -763 747 -724 781
rect -294 747 -255 781
rect -221 747 -197 781
rect -153 747 -125 781
rect -85 747 -53 781
rect -17 747 17 781
rect 53 747 85 781
rect 125 747 153 781
rect 197 747 221 781
rect 255 747 294 781
rect 724 747 763 781
rect 797 747 821 781
rect 865 747 893 781
rect 933 747 965 781
rect 1001 747 1035 781
rect 1071 747 1103 781
rect 1143 747 1171 781
rect 1215 747 1239 781
rect 1273 747 1312 781
rect 1742 747 1781 781
rect 1815 747 1839 781
rect 1883 747 1911 781
rect 1951 747 1983 781
rect 2019 747 2053 781
rect 2089 747 2121 781
rect 2161 747 2189 781
rect 2233 747 2257 781
rect 2291 747 2330 781
rect 2760 747 2799 781
rect 2833 747 2857 781
rect 2901 747 2929 781
rect 2969 747 3001 781
rect 3037 747 3071 781
rect 3107 747 3139 781
rect 3179 747 3207 781
rect 3251 747 3275 781
rect 3309 747 3348 781
rect 3778 747 3817 781
rect 3851 747 3875 781
rect 3919 747 3947 781
rect 3987 747 4019 781
rect 4055 747 4089 781
rect 4125 747 4157 781
rect 4197 747 4225 781
rect 4269 747 4293 781
rect 4327 747 4366 781
rect -4598 678 -4564 713
rect -4598 606 -4564 630
rect -4598 534 -4564 562
rect -4598 462 -4564 494
rect -4598 392 -4564 426
rect -4598 324 -4564 356
rect -4598 256 -4564 284
rect -4598 188 -4564 212
rect -4598 105 -4564 140
rect -3580 678 -3546 713
rect -3580 606 -3546 630
rect -3580 534 -3546 562
rect -3580 462 -3546 494
rect -3580 392 -3546 426
rect -3580 324 -3546 356
rect -3580 256 -3546 284
rect -3580 188 -3546 212
rect -3580 105 -3546 140
rect -2562 678 -2528 713
rect -2562 606 -2528 630
rect -2562 534 -2528 562
rect -2562 462 -2528 494
rect -2562 392 -2528 426
rect -2562 324 -2528 356
rect -2562 256 -2528 284
rect -2562 188 -2528 212
rect -2562 105 -2528 140
rect -1544 678 -1510 713
rect -1544 606 -1510 630
rect -1544 534 -1510 562
rect -1544 462 -1510 494
rect -1544 392 -1510 426
rect -1544 324 -1510 356
rect -1544 256 -1510 284
rect -1544 188 -1510 212
rect -1544 105 -1510 140
rect -526 678 -492 713
rect -526 606 -492 630
rect -526 534 -492 562
rect -526 462 -492 494
rect -526 392 -492 426
rect -526 324 -492 356
rect -526 256 -492 284
rect -526 188 -492 212
rect -526 105 -492 140
rect 492 678 526 713
rect 492 606 526 630
rect 492 534 526 562
rect 492 462 526 494
rect 492 392 526 426
rect 492 324 526 356
rect 492 256 526 284
rect 492 188 526 212
rect 492 105 526 140
rect 1510 678 1544 713
rect 1510 606 1544 630
rect 1510 534 1544 562
rect 1510 462 1544 494
rect 1510 392 1544 426
rect 1510 324 1544 356
rect 1510 256 1544 284
rect 1510 188 1544 212
rect 1510 105 1544 140
rect 2528 678 2562 713
rect 2528 606 2562 630
rect 2528 534 2562 562
rect 2528 462 2562 494
rect 2528 392 2562 426
rect 2528 324 2562 356
rect 2528 256 2562 284
rect 2528 188 2562 212
rect 2528 105 2562 140
rect 3546 678 3580 713
rect 3546 606 3580 630
rect 3546 534 3580 562
rect 3546 462 3580 494
rect 3546 392 3580 426
rect 3546 324 3580 356
rect 3546 256 3580 284
rect 3546 188 3580 212
rect 3546 105 3580 140
rect 4564 678 4598 713
rect 4564 606 4598 630
rect 4564 534 4598 562
rect 4564 462 4598 494
rect 4564 392 4598 426
rect 4564 324 4598 356
rect 4564 256 4598 284
rect 4564 188 4598 212
rect 4564 105 4598 140
rect -4366 37 -4327 71
rect -4293 37 -4269 71
rect -4225 37 -4197 71
rect -4157 37 -4125 71
rect -4089 37 -4055 71
rect -4019 37 -3987 71
rect -3947 37 -3919 71
rect -3875 37 -3851 71
rect -3817 37 -3778 71
rect -3348 37 -3309 71
rect -3275 37 -3251 71
rect -3207 37 -3179 71
rect -3139 37 -3107 71
rect -3071 37 -3037 71
rect -3001 37 -2969 71
rect -2929 37 -2901 71
rect -2857 37 -2833 71
rect -2799 37 -2760 71
rect -2330 37 -2291 71
rect -2257 37 -2233 71
rect -2189 37 -2161 71
rect -2121 37 -2089 71
rect -2053 37 -2019 71
rect -1983 37 -1951 71
rect -1911 37 -1883 71
rect -1839 37 -1815 71
rect -1781 37 -1742 71
rect -1312 37 -1273 71
rect -1239 37 -1215 71
rect -1171 37 -1143 71
rect -1103 37 -1071 71
rect -1035 37 -1001 71
rect -965 37 -933 71
rect -893 37 -865 71
rect -821 37 -797 71
rect -763 37 -724 71
rect -294 37 -255 71
rect -221 37 -197 71
rect -153 37 -125 71
rect -85 37 -53 71
rect -17 37 17 71
rect 53 37 85 71
rect 125 37 153 71
rect 197 37 221 71
rect 255 37 294 71
rect 724 37 763 71
rect 797 37 821 71
rect 865 37 893 71
rect 933 37 965 71
rect 1001 37 1035 71
rect 1071 37 1103 71
rect 1143 37 1171 71
rect 1215 37 1239 71
rect 1273 37 1312 71
rect 1742 37 1781 71
rect 1815 37 1839 71
rect 1883 37 1911 71
rect 1951 37 1983 71
rect 2019 37 2053 71
rect 2089 37 2121 71
rect 2161 37 2189 71
rect 2233 37 2257 71
rect 2291 37 2330 71
rect 2760 37 2799 71
rect 2833 37 2857 71
rect 2901 37 2929 71
rect 2969 37 3001 71
rect 3037 37 3071 71
rect 3107 37 3139 71
rect 3179 37 3207 71
rect 3251 37 3275 71
rect 3309 37 3348 71
rect 3778 37 3817 71
rect 3851 37 3875 71
rect 3919 37 3947 71
rect 3987 37 4019 71
rect 4055 37 4089 71
rect 4125 37 4157 71
rect 4197 37 4225 71
rect 4269 37 4293 71
rect 4327 37 4366 71
rect -4366 -71 -4327 -37
rect -4293 -71 -4269 -37
rect -4225 -71 -4197 -37
rect -4157 -71 -4125 -37
rect -4089 -71 -4055 -37
rect -4019 -71 -3987 -37
rect -3947 -71 -3919 -37
rect -3875 -71 -3851 -37
rect -3817 -71 -3778 -37
rect -3348 -71 -3309 -37
rect -3275 -71 -3251 -37
rect -3207 -71 -3179 -37
rect -3139 -71 -3107 -37
rect -3071 -71 -3037 -37
rect -3001 -71 -2969 -37
rect -2929 -71 -2901 -37
rect -2857 -71 -2833 -37
rect -2799 -71 -2760 -37
rect -2330 -71 -2291 -37
rect -2257 -71 -2233 -37
rect -2189 -71 -2161 -37
rect -2121 -71 -2089 -37
rect -2053 -71 -2019 -37
rect -1983 -71 -1951 -37
rect -1911 -71 -1883 -37
rect -1839 -71 -1815 -37
rect -1781 -71 -1742 -37
rect -1312 -71 -1273 -37
rect -1239 -71 -1215 -37
rect -1171 -71 -1143 -37
rect -1103 -71 -1071 -37
rect -1035 -71 -1001 -37
rect -965 -71 -933 -37
rect -893 -71 -865 -37
rect -821 -71 -797 -37
rect -763 -71 -724 -37
rect -294 -71 -255 -37
rect -221 -71 -197 -37
rect -153 -71 -125 -37
rect -85 -71 -53 -37
rect -17 -71 17 -37
rect 53 -71 85 -37
rect 125 -71 153 -37
rect 197 -71 221 -37
rect 255 -71 294 -37
rect 724 -71 763 -37
rect 797 -71 821 -37
rect 865 -71 893 -37
rect 933 -71 965 -37
rect 1001 -71 1035 -37
rect 1071 -71 1103 -37
rect 1143 -71 1171 -37
rect 1215 -71 1239 -37
rect 1273 -71 1312 -37
rect 1742 -71 1781 -37
rect 1815 -71 1839 -37
rect 1883 -71 1911 -37
rect 1951 -71 1983 -37
rect 2019 -71 2053 -37
rect 2089 -71 2121 -37
rect 2161 -71 2189 -37
rect 2233 -71 2257 -37
rect 2291 -71 2330 -37
rect 2760 -71 2799 -37
rect 2833 -71 2857 -37
rect 2901 -71 2929 -37
rect 2969 -71 3001 -37
rect 3037 -71 3071 -37
rect 3107 -71 3139 -37
rect 3179 -71 3207 -37
rect 3251 -71 3275 -37
rect 3309 -71 3348 -37
rect 3778 -71 3817 -37
rect 3851 -71 3875 -37
rect 3919 -71 3947 -37
rect 3987 -71 4019 -37
rect 4055 -71 4089 -37
rect 4125 -71 4157 -37
rect 4197 -71 4225 -37
rect 4269 -71 4293 -37
rect 4327 -71 4366 -37
rect -4598 -140 -4564 -105
rect -4598 -212 -4564 -188
rect -4598 -284 -4564 -256
rect -4598 -356 -4564 -324
rect -4598 -426 -4564 -392
rect -4598 -494 -4564 -462
rect -4598 -562 -4564 -534
rect -4598 -630 -4564 -606
rect -4598 -713 -4564 -678
rect -3580 -140 -3546 -105
rect -3580 -212 -3546 -188
rect -3580 -284 -3546 -256
rect -3580 -356 -3546 -324
rect -3580 -426 -3546 -392
rect -3580 -494 -3546 -462
rect -3580 -562 -3546 -534
rect -3580 -630 -3546 -606
rect -3580 -713 -3546 -678
rect -2562 -140 -2528 -105
rect -2562 -212 -2528 -188
rect -2562 -284 -2528 -256
rect -2562 -356 -2528 -324
rect -2562 -426 -2528 -392
rect -2562 -494 -2528 -462
rect -2562 -562 -2528 -534
rect -2562 -630 -2528 -606
rect -2562 -713 -2528 -678
rect -1544 -140 -1510 -105
rect -1544 -212 -1510 -188
rect -1544 -284 -1510 -256
rect -1544 -356 -1510 -324
rect -1544 -426 -1510 -392
rect -1544 -494 -1510 -462
rect -1544 -562 -1510 -534
rect -1544 -630 -1510 -606
rect -1544 -713 -1510 -678
rect -526 -140 -492 -105
rect -526 -212 -492 -188
rect -526 -284 -492 -256
rect -526 -356 -492 -324
rect -526 -426 -492 -392
rect -526 -494 -492 -462
rect -526 -562 -492 -534
rect -526 -630 -492 -606
rect -526 -713 -492 -678
rect 492 -140 526 -105
rect 492 -212 526 -188
rect 492 -284 526 -256
rect 492 -356 526 -324
rect 492 -426 526 -392
rect 492 -494 526 -462
rect 492 -562 526 -534
rect 492 -630 526 -606
rect 492 -713 526 -678
rect 1510 -140 1544 -105
rect 1510 -212 1544 -188
rect 1510 -284 1544 -256
rect 1510 -356 1544 -324
rect 1510 -426 1544 -392
rect 1510 -494 1544 -462
rect 1510 -562 1544 -534
rect 1510 -630 1544 -606
rect 1510 -713 1544 -678
rect 2528 -140 2562 -105
rect 2528 -212 2562 -188
rect 2528 -284 2562 -256
rect 2528 -356 2562 -324
rect 2528 -426 2562 -392
rect 2528 -494 2562 -462
rect 2528 -562 2562 -534
rect 2528 -630 2562 -606
rect 2528 -713 2562 -678
rect 3546 -140 3580 -105
rect 3546 -212 3580 -188
rect 3546 -284 3580 -256
rect 3546 -356 3580 -324
rect 3546 -426 3580 -392
rect 3546 -494 3580 -462
rect 3546 -562 3580 -534
rect 3546 -630 3580 -606
rect 3546 -713 3580 -678
rect 4564 -140 4598 -105
rect 4564 -212 4598 -188
rect 4564 -284 4598 -256
rect 4564 -356 4598 -324
rect 4564 -426 4598 -392
rect 4564 -494 4598 -462
rect 4564 -562 4598 -534
rect 4564 -630 4598 -606
rect 4564 -713 4598 -678
rect -4366 -781 -4327 -747
rect -4293 -781 -4269 -747
rect -4225 -781 -4197 -747
rect -4157 -781 -4125 -747
rect -4089 -781 -4055 -747
rect -4019 -781 -3987 -747
rect -3947 -781 -3919 -747
rect -3875 -781 -3851 -747
rect -3817 -781 -3778 -747
rect -3348 -781 -3309 -747
rect -3275 -781 -3251 -747
rect -3207 -781 -3179 -747
rect -3139 -781 -3107 -747
rect -3071 -781 -3037 -747
rect -3001 -781 -2969 -747
rect -2929 -781 -2901 -747
rect -2857 -781 -2833 -747
rect -2799 -781 -2760 -747
rect -2330 -781 -2291 -747
rect -2257 -781 -2233 -747
rect -2189 -781 -2161 -747
rect -2121 -781 -2089 -747
rect -2053 -781 -2019 -747
rect -1983 -781 -1951 -747
rect -1911 -781 -1883 -747
rect -1839 -781 -1815 -747
rect -1781 -781 -1742 -747
rect -1312 -781 -1273 -747
rect -1239 -781 -1215 -747
rect -1171 -781 -1143 -747
rect -1103 -781 -1071 -747
rect -1035 -781 -1001 -747
rect -965 -781 -933 -747
rect -893 -781 -865 -747
rect -821 -781 -797 -747
rect -763 -781 -724 -747
rect -294 -781 -255 -747
rect -221 -781 -197 -747
rect -153 -781 -125 -747
rect -85 -781 -53 -747
rect -17 -781 17 -747
rect 53 -781 85 -747
rect 125 -781 153 -747
rect 197 -781 221 -747
rect 255 -781 294 -747
rect 724 -781 763 -747
rect 797 -781 821 -747
rect 865 -781 893 -747
rect 933 -781 965 -747
rect 1001 -781 1035 -747
rect 1071 -781 1103 -747
rect 1143 -781 1171 -747
rect 1215 -781 1239 -747
rect 1273 -781 1312 -747
rect 1742 -781 1781 -747
rect 1815 -781 1839 -747
rect 1883 -781 1911 -747
rect 1951 -781 1983 -747
rect 2019 -781 2053 -747
rect 2089 -781 2121 -747
rect 2161 -781 2189 -747
rect 2233 -781 2257 -747
rect 2291 -781 2330 -747
rect 2760 -781 2799 -747
rect 2833 -781 2857 -747
rect 2901 -781 2929 -747
rect 2969 -781 3001 -747
rect 3037 -781 3071 -747
rect 3107 -781 3139 -747
rect 3179 -781 3207 -747
rect 3251 -781 3275 -747
rect 3309 -781 3348 -747
rect 3778 -781 3817 -747
rect 3851 -781 3875 -747
rect 3919 -781 3947 -747
rect 3987 -781 4019 -747
rect 4055 -781 4089 -747
rect 4125 -781 4157 -747
rect 4197 -781 4225 -747
rect 4269 -781 4293 -747
rect 4327 -781 4366 -747
rect -4366 -889 -4327 -855
rect -4293 -889 -4269 -855
rect -4225 -889 -4197 -855
rect -4157 -889 -4125 -855
rect -4089 -889 -4055 -855
rect -4019 -889 -3987 -855
rect -3947 -889 -3919 -855
rect -3875 -889 -3851 -855
rect -3817 -889 -3778 -855
rect -3348 -889 -3309 -855
rect -3275 -889 -3251 -855
rect -3207 -889 -3179 -855
rect -3139 -889 -3107 -855
rect -3071 -889 -3037 -855
rect -3001 -889 -2969 -855
rect -2929 -889 -2901 -855
rect -2857 -889 -2833 -855
rect -2799 -889 -2760 -855
rect -2330 -889 -2291 -855
rect -2257 -889 -2233 -855
rect -2189 -889 -2161 -855
rect -2121 -889 -2089 -855
rect -2053 -889 -2019 -855
rect -1983 -889 -1951 -855
rect -1911 -889 -1883 -855
rect -1839 -889 -1815 -855
rect -1781 -889 -1742 -855
rect -1312 -889 -1273 -855
rect -1239 -889 -1215 -855
rect -1171 -889 -1143 -855
rect -1103 -889 -1071 -855
rect -1035 -889 -1001 -855
rect -965 -889 -933 -855
rect -893 -889 -865 -855
rect -821 -889 -797 -855
rect -763 -889 -724 -855
rect -294 -889 -255 -855
rect -221 -889 -197 -855
rect -153 -889 -125 -855
rect -85 -889 -53 -855
rect -17 -889 17 -855
rect 53 -889 85 -855
rect 125 -889 153 -855
rect 197 -889 221 -855
rect 255 -889 294 -855
rect 724 -889 763 -855
rect 797 -889 821 -855
rect 865 -889 893 -855
rect 933 -889 965 -855
rect 1001 -889 1035 -855
rect 1071 -889 1103 -855
rect 1143 -889 1171 -855
rect 1215 -889 1239 -855
rect 1273 -889 1312 -855
rect 1742 -889 1781 -855
rect 1815 -889 1839 -855
rect 1883 -889 1911 -855
rect 1951 -889 1983 -855
rect 2019 -889 2053 -855
rect 2089 -889 2121 -855
rect 2161 -889 2189 -855
rect 2233 -889 2257 -855
rect 2291 -889 2330 -855
rect 2760 -889 2799 -855
rect 2833 -889 2857 -855
rect 2901 -889 2929 -855
rect 2969 -889 3001 -855
rect 3037 -889 3071 -855
rect 3107 -889 3139 -855
rect 3179 -889 3207 -855
rect 3251 -889 3275 -855
rect 3309 -889 3348 -855
rect 3778 -889 3817 -855
rect 3851 -889 3875 -855
rect 3919 -889 3947 -855
rect 3987 -889 4019 -855
rect 4055 -889 4089 -855
rect 4125 -889 4157 -855
rect 4197 -889 4225 -855
rect 4269 -889 4293 -855
rect 4327 -889 4366 -855
rect -4598 -958 -4564 -923
rect -4598 -1030 -4564 -1006
rect -4598 -1102 -4564 -1074
rect -4598 -1174 -4564 -1142
rect -4598 -1244 -4564 -1210
rect -4598 -1312 -4564 -1280
rect -4598 -1380 -4564 -1352
rect -4598 -1448 -4564 -1424
rect -4598 -1531 -4564 -1496
rect -3580 -958 -3546 -923
rect -3580 -1030 -3546 -1006
rect -3580 -1102 -3546 -1074
rect -3580 -1174 -3546 -1142
rect -3580 -1244 -3546 -1210
rect -3580 -1312 -3546 -1280
rect -3580 -1380 -3546 -1352
rect -3580 -1448 -3546 -1424
rect -3580 -1531 -3546 -1496
rect -2562 -958 -2528 -923
rect -2562 -1030 -2528 -1006
rect -2562 -1102 -2528 -1074
rect -2562 -1174 -2528 -1142
rect -2562 -1244 -2528 -1210
rect -2562 -1312 -2528 -1280
rect -2562 -1380 -2528 -1352
rect -2562 -1448 -2528 -1424
rect -2562 -1531 -2528 -1496
rect -1544 -958 -1510 -923
rect -1544 -1030 -1510 -1006
rect -1544 -1102 -1510 -1074
rect -1544 -1174 -1510 -1142
rect -1544 -1244 -1510 -1210
rect -1544 -1312 -1510 -1280
rect -1544 -1380 -1510 -1352
rect -1544 -1448 -1510 -1424
rect -1544 -1531 -1510 -1496
rect -526 -958 -492 -923
rect -526 -1030 -492 -1006
rect -526 -1102 -492 -1074
rect -526 -1174 -492 -1142
rect -526 -1244 -492 -1210
rect -526 -1312 -492 -1280
rect -526 -1380 -492 -1352
rect -526 -1448 -492 -1424
rect -526 -1531 -492 -1496
rect 492 -958 526 -923
rect 492 -1030 526 -1006
rect 492 -1102 526 -1074
rect 492 -1174 526 -1142
rect 492 -1244 526 -1210
rect 492 -1312 526 -1280
rect 492 -1380 526 -1352
rect 492 -1448 526 -1424
rect 492 -1531 526 -1496
rect 1510 -958 1544 -923
rect 1510 -1030 1544 -1006
rect 1510 -1102 1544 -1074
rect 1510 -1174 1544 -1142
rect 1510 -1244 1544 -1210
rect 1510 -1312 1544 -1280
rect 1510 -1380 1544 -1352
rect 1510 -1448 1544 -1424
rect 1510 -1531 1544 -1496
rect 2528 -958 2562 -923
rect 2528 -1030 2562 -1006
rect 2528 -1102 2562 -1074
rect 2528 -1174 2562 -1142
rect 2528 -1244 2562 -1210
rect 2528 -1312 2562 -1280
rect 2528 -1380 2562 -1352
rect 2528 -1448 2562 -1424
rect 2528 -1531 2562 -1496
rect 3546 -958 3580 -923
rect 3546 -1030 3580 -1006
rect 3546 -1102 3580 -1074
rect 3546 -1174 3580 -1142
rect 3546 -1244 3580 -1210
rect 3546 -1312 3580 -1280
rect 3546 -1380 3580 -1352
rect 3546 -1448 3580 -1424
rect 3546 -1531 3580 -1496
rect 4564 -958 4598 -923
rect 4564 -1030 4598 -1006
rect 4564 -1102 4598 -1074
rect 4564 -1174 4598 -1142
rect 4564 -1244 4598 -1210
rect 4564 -1312 4598 -1280
rect 4564 -1380 4598 -1352
rect 4564 -1448 4598 -1424
rect 4564 -1531 4598 -1496
rect -4366 -1599 -4327 -1565
rect -4293 -1599 -4269 -1565
rect -4225 -1599 -4197 -1565
rect -4157 -1599 -4125 -1565
rect -4089 -1599 -4055 -1565
rect -4019 -1599 -3987 -1565
rect -3947 -1599 -3919 -1565
rect -3875 -1599 -3851 -1565
rect -3817 -1599 -3778 -1565
rect -3348 -1599 -3309 -1565
rect -3275 -1599 -3251 -1565
rect -3207 -1599 -3179 -1565
rect -3139 -1599 -3107 -1565
rect -3071 -1599 -3037 -1565
rect -3001 -1599 -2969 -1565
rect -2929 -1599 -2901 -1565
rect -2857 -1599 -2833 -1565
rect -2799 -1599 -2760 -1565
rect -2330 -1599 -2291 -1565
rect -2257 -1599 -2233 -1565
rect -2189 -1599 -2161 -1565
rect -2121 -1599 -2089 -1565
rect -2053 -1599 -2019 -1565
rect -1983 -1599 -1951 -1565
rect -1911 -1599 -1883 -1565
rect -1839 -1599 -1815 -1565
rect -1781 -1599 -1742 -1565
rect -1312 -1599 -1273 -1565
rect -1239 -1599 -1215 -1565
rect -1171 -1599 -1143 -1565
rect -1103 -1599 -1071 -1565
rect -1035 -1599 -1001 -1565
rect -965 -1599 -933 -1565
rect -893 -1599 -865 -1565
rect -821 -1599 -797 -1565
rect -763 -1599 -724 -1565
rect -294 -1599 -255 -1565
rect -221 -1599 -197 -1565
rect -153 -1599 -125 -1565
rect -85 -1599 -53 -1565
rect -17 -1599 17 -1565
rect 53 -1599 85 -1565
rect 125 -1599 153 -1565
rect 197 -1599 221 -1565
rect 255 -1599 294 -1565
rect 724 -1599 763 -1565
rect 797 -1599 821 -1565
rect 865 -1599 893 -1565
rect 933 -1599 965 -1565
rect 1001 -1599 1035 -1565
rect 1071 -1599 1103 -1565
rect 1143 -1599 1171 -1565
rect 1215 -1599 1239 -1565
rect 1273 -1599 1312 -1565
rect 1742 -1599 1781 -1565
rect 1815 -1599 1839 -1565
rect 1883 -1599 1911 -1565
rect 1951 -1599 1983 -1565
rect 2019 -1599 2053 -1565
rect 2089 -1599 2121 -1565
rect 2161 -1599 2189 -1565
rect 2233 -1599 2257 -1565
rect 2291 -1599 2330 -1565
rect 2760 -1599 2799 -1565
rect 2833 -1599 2857 -1565
rect 2901 -1599 2929 -1565
rect 2969 -1599 3001 -1565
rect 3037 -1599 3071 -1565
rect 3107 -1599 3139 -1565
rect 3179 -1599 3207 -1565
rect 3251 -1599 3275 -1565
rect 3309 -1599 3348 -1565
rect 3778 -1599 3817 -1565
rect 3851 -1599 3875 -1565
rect 3919 -1599 3947 -1565
rect 3987 -1599 4019 -1565
rect 4055 -1599 4089 -1565
rect 4125 -1599 4157 -1565
rect 4197 -1599 4225 -1565
rect 4269 -1599 4293 -1565
rect 4327 -1599 4366 -1565
<< viali >>
rect -4269 1565 -4259 1599
rect -4259 1565 -4235 1599
rect -4197 1565 -4191 1599
rect -4191 1565 -4163 1599
rect -4125 1565 -4123 1599
rect -4123 1565 -4091 1599
rect -4053 1565 -4021 1599
rect -4021 1565 -4019 1599
rect -3981 1565 -3953 1599
rect -3953 1565 -3947 1599
rect -3909 1565 -3885 1599
rect -3885 1565 -3875 1599
rect -3251 1565 -3241 1599
rect -3241 1565 -3217 1599
rect -3179 1565 -3173 1599
rect -3173 1565 -3145 1599
rect -3107 1565 -3105 1599
rect -3105 1565 -3073 1599
rect -3035 1565 -3003 1599
rect -3003 1565 -3001 1599
rect -2963 1565 -2935 1599
rect -2935 1565 -2929 1599
rect -2891 1565 -2867 1599
rect -2867 1565 -2857 1599
rect -2233 1565 -2223 1599
rect -2223 1565 -2199 1599
rect -2161 1565 -2155 1599
rect -2155 1565 -2127 1599
rect -2089 1565 -2087 1599
rect -2087 1565 -2055 1599
rect -2017 1565 -1985 1599
rect -1985 1565 -1983 1599
rect -1945 1565 -1917 1599
rect -1917 1565 -1911 1599
rect -1873 1565 -1849 1599
rect -1849 1565 -1839 1599
rect -1215 1565 -1205 1599
rect -1205 1565 -1181 1599
rect -1143 1565 -1137 1599
rect -1137 1565 -1109 1599
rect -1071 1565 -1069 1599
rect -1069 1565 -1037 1599
rect -999 1565 -967 1599
rect -967 1565 -965 1599
rect -927 1565 -899 1599
rect -899 1565 -893 1599
rect -855 1565 -831 1599
rect -831 1565 -821 1599
rect -197 1565 -187 1599
rect -187 1565 -163 1599
rect -125 1565 -119 1599
rect -119 1565 -91 1599
rect -53 1565 -51 1599
rect -51 1565 -19 1599
rect 19 1565 51 1599
rect 51 1565 53 1599
rect 91 1565 119 1599
rect 119 1565 125 1599
rect 163 1565 187 1599
rect 187 1565 197 1599
rect 821 1565 831 1599
rect 831 1565 855 1599
rect 893 1565 899 1599
rect 899 1565 927 1599
rect 965 1565 967 1599
rect 967 1565 999 1599
rect 1037 1565 1069 1599
rect 1069 1565 1071 1599
rect 1109 1565 1137 1599
rect 1137 1565 1143 1599
rect 1181 1565 1205 1599
rect 1205 1565 1215 1599
rect 1839 1565 1849 1599
rect 1849 1565 1873 1599
rect 1911 1565 1917 1599
rect 1917 1565 1945 1599
rect 1983 1565 1985 1599
rect 1985 1565 2017 1599
rect 2055 1565 2087 1599
rect 2087 1565 2089 1599
rect 2127 1565 2155 1599
rect 2155 1565 2161 1599
rect 2199 1565 2223 1599
rect 2223 1565 2233 1599
rect 2857 1565 2867 1599
rect 2867 1565 2891 1599
rect 2929 1565 2935 1599
rect 2935 1565 2963 1599
rect 3001 1565 3003 1599
rect 3003 1565 3035 1599
rect 3073 1565 3105 1599
rect 3105 1565 3107 1599
rect 3145 1565 3173 1599
rect 3173 1565 3179 1599
rect 3217 1565 3241 1599
rect 3241 1565 3251 1599
rect 3875 1565 3885 1599
rect 3885 1565 3909 1599
rect 3947 1565 3953 1599
rect 3953 1565 3981 1599
rect 4019 1565 4021 1599
rect 4021 1565 4053 1599
rect 4091 1565 4123 1599
rect 4123 1565 4125 1599
rect 4163 1565 4191 1599
rect 4191 1565 4197 1599
rect 4235 1565 4259 1599
rect 4259 1565 4269 1599
rect -4598 1482 -4564 1496
rect -4598 1462 -4564 1482
rect -4598 1414 -4564 1424
rect -4598 1390 -4564 1414
rect -4598 1346 -4564 1352
rect -4598 1318 -4564 1346
rect -4598 1278 -4564 1280
rect -4598 1246 -4564 1278
rect -4598 1176 -4564 1208
rect -4598 1174 -4564 1176
rect -4598 1108 -4564 1136
rect -4598 1102 -4564 1108
rect -4598 1040 -4564 1064
rect -4598 1030 -4564 1040
rect -4598 972 -4564 992
rect -4598 958 -4564 972
rect -3580 1482 -3546 1496
rect -3580 1462 -3546 1482
rect -3580 1414 -3546 1424
rect -3580 1390 -3546 1414
rect -3580 1346 -3546 1352
rect -3580 1318 -3546 1346
rect -3580 1278 -3546 1280
rect -3580 1246 -3546 1278
rect -3580 1176 -3546 1208
rect -3580 1174 -3546 1176
rect -3580 1108 -3546 1136
rect -3580 1102 -3546 1108
rect -3580 1040 -3546 1064
rect -3580 1030 -3546 1040
rect -3580 972 -3546 992
rect -3580 958 -3546 972
rect -2562 1482 -2528 1496
rect -2562 1462 -2528 1482
rect -2562 1414 -2528 1424
rect -2562 1390 -2528 1414
rect -2562 1346 -2528 1352
rect -2562 1318 -2528 1346
rect -2562 1278 -2528 1280
rect -2562 1246 -2528 1278
rect -2562 1176 -2528 1208
rect -2562 1174 -2528 1176
rect -2562 1108 -2528 1136
rect -2562 1102 -2528 1108
rect -2562 1040 -2528 1064
rect -2562 1030 -2528 1040
rect -2562 972 -2528 992
rect -2562 958 -2528 972
rect -1544 1482 -1510 1496
rect -1544 1462 -1510 1482
rect -1544 1414 -1510 1424
rect -1544 1390 -1510 1414
rect -1544 1346 -1510 1352
rect -1544 1318 -1510 1346
rect -1544 1278 -1510 1280
rect -1544 1246 -1510 1278
rect -1544 1176 -1510 1208
rect -1544 1174 -1510 1176
rect -1544 1108 -1510 1136
rect -1544 1102 -1510 1108
rect -1544 1040 -1510 1064
rect -1544 1030 -1510 1040
rect -1544 972 -1510 992
rect -1544 958 -1510 972
rect -526 1482 -492 1496
rect -526 1462 -492 1482
rect -526 1414 -492 1424
rect -526 1390 -492 1414
rect -526 1346 -492 1352
rect -526 1318 -492 1346
rect -526 1278 -492 1280
rect -526 1246 -492 1278
rect -526 1176 -492 1208
rect -526 1174 -492 1176
rect -526 1108 -492 1136
rect -526 1102 -492 1108
rect -526 1040 -492 1064
rect -526 1030 -492 1040
rect -526 972 -492 992
rect -526 958 -492 972
rect 492 1482 526 1496
rect 492 1462 526 1482
rect 492 1414 526 1424
rect 492 1390 526 1414
rect 492 1346 526 1352
rect 492 1318 526 1346
rect 492 1278 526 1280
rect 492 1246 526 1278
rect 492 1176 526 1208
rect 492 1174 526 1176
rect 492 1108 526 1136
rect 492 1102 526 1108
rect 492 1040 526 1064
rect 492 1030 526 1040
rect 492 972 526 992
rect 492 958 526 972
rect 1510 1482 1544 1496
rect 1510 1462 1544 1482
rect 1510 1414 1544 1424
rect 1510 1390 1544 1414
rect 1510 1346 1544 1352
rect 1510 1318 1544 1346
rect 1510 1278 1544 1280
rect 1510 1246 1544 1278
rect 1510 1176 1544 1208
rect 1510 1174 1544 1176
rect 1510 1108 1544 1136
rect 1510 1102 1544 1108
rect 1510 1040 1544 1064
rect 1510 1030 1544 1040
rect 1510 972 1544 992
rect 1510 958 1544 972
rect 2528 1482 2562 1496
rect 2528 1462 2562 1482
rect 2528 1414 2562 1424
rect 2528 1390 2562 1414
rect 2528 1346 2562 1352
rect 2528 1318 2562 1346
rect 2528 1278 2562 1280
rect 2528 1246 2562 1278
rect 2528 1176 2562 1208
rect 2528 1174 2562 1176
rect 2528 1108 2562 1136
rect 2528 1102 2562 1108
rect 2528 1040 2562 1064
rect 2528 1030 2562 1040
rect 2528 972 2562 992
rect 2528 958 2562 972
rect 3546 1482 3580 1496
rect 3546 1462 3580 1482
rect 3546 1414 3580 1424
rect 3546 1390 3580 1414
rect 3546 1346 3580 1352
rect 3546 1318 3580 1346
rect 3546 1278 3580 1280
rect 3546 1246 3580 1278
rect 3546 1176 3580 1208
rect 3546 1174 3580 1176
rect 3546 1108 3580 1136
rect 3546 1102 3580 1108
rect 3546 1040 3580 1064
rect 3546 1030 3580 1040
rect 3546 972 3580 992
rect 3546 958 3580 972
rect 4564 1482 4598 1496
rect 4564 1462 4598 1482
rect 4564 1414 4598 1424
rect 4564 1390 4598 1414
rect 4564 1346 4598 1352
rect 4564 1318 4598 1346
rect 4564 1278 4598 1280
rect 4564 1246 4598 1278
rect 4564 1176 4598 1208
rect 4564 1174 4598 1176
rect 4564 1108 4598 1136
rect 4564 1102 4598 1108
rect 4564 1040 4598 1064
rect 4564 1030 4598 1040
rect 4564 972 4598 992
rect 4564 958 4598 972
rect -4269 855 -4259 889
rect -4259 855 -4235 889
rect -4197 855 -4191 889
rect -4191 855 -4163 889
rect -4125 855 -4123 889
rect -4123 855 -4091 889
rect -4053 855 -4021 889
rect -4021 855 -4019 889
rect -3981 855 -3953 889
rect -3953 855 -3947 889
rect -3909 855 -3885 889
rect -3885 855 -3875 889
rect -3251 855 -3241 889
rect -3241 855 -3217 889
rect -3179 855 -3173 889
rect -3173 855 -3145 889
rect -3107 855 -3105 889
rect -3105 855 -3073 889
rect -3035 855 -3003 889
rect -3003 855 -3001 889
rect -2963 855 -2935 889
rect -2935 855 -2929 889
rect -2891 855 -2867 889
rect -2867 855 -2857 889
rect -2233 855 -2223 889
rect -2223 855 -2199 889
rect -2161 855 -2155 889
rect -2155 855 -2127 889
rect -2089 855 -2087 889
rect -2087 855 -2055 889
rect -2017 855 -1985 889
rect -1985 855 -1983 889
rect -1945 855 -1917 889
rect -1917 855 -1911 889
rect -1873 855 -1849 889
rect -1849 855 -1839 889
rect -1215 855 -1205 889
rect -1205 855 -1181 889
rect -1143 855 -1137 889
rect -1137 855 -1109 889
rect -1071 855 -1069 889
rect -1069 855 -1037 889
rect -999 855 -967 889
rect -967 855 -965 889
rect -927 855 -899 889
rect -899 855 -893 889
rect -855 855 -831 889
rect -831 855 -821 889
rect -197 855 -187 889
rect -187 855 -163 889
rect -125 855 -119 889
rect -119 855 -91 889
rect -53 855 -51 889
rect -51 855 -19 889
rect 19 855 51 889
rect 51 855 53 889
rect 91 855 119 889
rect 119 855 125 889
rect 163 855 187 889
rect 187 855 197 889
rect 821 855 831 889
rect 831 855 855 889
rect 893 855 899 889
rect 899 855 927 889
rect 965 855 967 889
rect 967 855 999 889
rect 1037 855 1069 889
rect 1069 855 1071 889
rect 1109 855 1137 889
rect 1137 855 1143 889
rect 1181 855 1205 889
rect 1205 855 1215 889
rect 1839 855 1849 889
rect 1849 855 1873 889
rect 1911 855 1917 889
rect 1917 855 1945 889
rect 1983 855 1985 889
rect 1985 855 2017 889
rect 2055 855 2087 889
rect 2087 855 2089 889
rect 2127 855 2155 889
rect 2155 855 2161 889
rect 2199 855 2223 889
rect 2223 855 2233 889
rect 2857 855 2867 889
rect 2867 855 2891 889
rect 2929 855 2935 889
rect 2935 855 2963 889
rect 3001 855 3003 889
rect 3003 855 3035 889
rect 3073 855 3105 889
rect 3105 855 3107 889
rect 3145 855 3173 889
rect 3173 855 3179 889
rect 3217 855 3241 889
rect 3241 855 3251 889
rect 3875 855 3885 889
rect 3885 855 3909 889
rect 3947 855 3953 889
rect 3953 855 3981 889
rect 4019 855 4021 889
rect 4021 855 4053 889
rect 4091 855 4123 889
rect 4123 855 4125 889
rect 4163 855 4191 889
rect 4191 855 4197 889
rect 4235 855 4259 889
rect 4259 855 4269 889
rect -4269 747 -4259 781
rect -4259 747 -4235 781
rect -4197 747 -4191 781
rect -4191 747 -4163 781
rect -4125 747 -4123 781
rect -4123 747 -4091 781
rect -4053 747 -4021 781
rect -4021 747 -4019 781
rect -3981 747 -3953 781
rect -3953 747 -3947 781
rect -3909 747 -3885 781
rect -3885 747 -3875 781
rect -3251 747 -3241 781
rect -3241 747 -3217 781
rect -3179 747 -3173 781
rect -3173 747 -3145 781
rect -3107 747 -3105 781
rect -3105 747 -3073 781
rect -3035 747 -3003 781
rect -3003 747 -3001 781
rect -2963 747 -2935 781
rect -2935 747 -2929 781
rect -2891 747 -2867 781
rect -2867 747 -2857 781
rect -2233 747 -2223 781
rect -2223 747 -2199 781
rect -2161 747 -2155 781
rect -2155 747 -2127 781
rect -2089 747 -2087 781
rect -2087 747 -2055 781
rect -2017 747 -1985 781
rect -1985 747 -1983 781
rect -1945 747 -1917 781
rect -1917 747 -1911 781
rect -1873 747 -1849 781
rect -1849 747 -1839 781
rect -1215 747 -1205 781
rect -1205 747 -1181 781
rect -1143 747 -1137 781
rect -1137 747 -1109 781
rect -1071 747 -1069 781
rect -1069 747 -1037 781
rect -999 747 -967 781
rect -967 747 -965 781
rect -927 747 -899 781
rect -899 747 -893 781
rect -855 747 -831 781
rect -831 747 -821 781
rect -197 747 -187 781
rect -187 747 -163 781
rect -125 747 -119 781
rect -119 747 -91 781
rect -53 747 -51 781
rect -51 747 -19 781
rect 19 747 51 781
rect 51 747 53 781
rect 91 747 119 781
rect 119 747 125 781
rect 163 747 187 781
rect 187 747 197 781
rect 821 747 831 781
rect 831 747 855 781
rect 893 747 899 781
rect 899 747 927 781
rect 965 747 967 781
rect 967 747 999 781
rect 1037 747 1069 781
rect 1069 747 1071 781
rect 1109 747 1137 781
rect 1137 747 1143 781
rect 1181 747 1205 781
rect 1205 747 1215 781
rect 1839 747 1849 781
rect 1849 747 1873 781
rect 1911 747 1917 781
rect 1917 747 1945 781
rect 1983 747 1985 781
rect 1985 747 2017 781
rect 2055 747 2087 781
rect 2087 747 2089 781
rect 2127 747 2155 781
rect 2155 747 2161 781
rect 2199 747 2223 781
rect 2223 747 2233 781
rect 2857 747 2867 781
rect 2867 747 2891 781
rect 2929 747 2935 781
rect 2935 747 2963 781
rect 3001 747 3003 781
rect 3003 747 3035 781
rect 3073 747 3105 781
rect 3105 747 3107 781
rect 3145 747 3173 781
rect 3173 747 3179 781
rect 3217 747 3241 781
rect 3241 747 3251 781
rect 3875 747 3885 781
rect 3885 747 3909 781
rect 3947 747 3953 781
rect 3953 747 3981 781
rect 4019 747 4021 781
rect 4021 747 4053 781
rect 4091 747 4123 781
rect 4123 747 4125 781
rect 4163 747 4191 781
rect 4191 747 4197 781
rect 4235 747 4259 781
rect 4259 747 4269 781
rect -4598 664 -4564 678
rect -4598 644 -4564 664
rect -4598 596 -4564 606
rect -4598 572 -4564 596
rect -4598 528 -4564 534
rect -4598 500 -4564 528
rect -4598 460 -4564 462
rect -4598 428 -4564 460
rect -4598 358 -4564 390
rect -4598 356 -4564 358
rect -4598 290 -4564 318
rect -4598 284 -4564 290
rect -4598 222 -4564 246
rect -4598 212 -4564 222
rect -4598 154 -4564 174
rect -4598 140 -4564 154
rect -3580 664 -3546 678
rect -3580 644 -3546 664
rect -3580 596 -3546 606
rect -3580 572 -3546 596
rect -3580 528 -3546 534
rect -3580 500 -3546 528
rect -3580 460 -3546 462
rect -3580 428 -3546 460
rect -3580 358 -3546 390
rect -3580 356 -3546 358
rect -3580 290 -3546 318
rect -3580 284 -3546 290
rect -3580 222 -3546 246
rect -3580 212 -3546 222
rect -3580 154 -3546 174
rect -3580 140 -3546 154
rect -2562 664 -2528 678
rect -2562 644 -2528 664
rect -2562 596 -2528 606
rect -2562 572 -2528 596
rect -2562 528 -2528 534
rect -2562 500 -2528 528
rect -2562 460 -2528 462
rect -2562 428 -2528 460
rect -2562 358 -2528 390
rect -2562 356 -2528 358
rect -2562 290 -2528 318
rect -2562 284 -2528 290
rect -2562 222 -2528 246
rect -2562 212 -2528 222
rect -2562 154 -2528 174
rect -2562 140 -2528 154
rect -1544 664 -1510 678
rect -1544 644 -1510 664
rect -1544 596 -1510 606
rect -1544 572 -1510 596
rect -1544 528 -1510 534
rect -1544 500 -1510 528
rect -1544 460 -1510 462
rect -1544 428 -1510 460
rect -1544 358 -1510 390
rect -1544 356 -1510 358
rect -1544 290 -1510 318
rect -1544 284 -1510 290
rect -1544 222 -1510 246
rect -1544 212 -1510 222
rect -1544 154 -1510 174
rect -1544 140 -1510 154
rect -526 664 -492 678
rect -526 644 -492 664
rect -526 596 -492 606
rect -526 572 -492 596
rect -526 528 -492 534
rect -526 500 -492 528
rect -526 460 -492 462
rect -526 428 -492 460
rect -526 358 -492 390
rect -526 356 -492 358
rect -526 290 -492 318
rect -526 284 -492 290
rect -526 222 -492 246
rect -526 212 -492 222
rect -526 154 -492 174
rect -526 140 -492 154
rect 492 664 526 678
rect 492 644 526 664
rect 492 596 526 606
rect 492 572 526 596
rect 492 528 526 534
rect 492 500 526 528
rect 492 460 526 462
rect 492 428 526 460
rect 492 358 526 390
rect 492 356 526 358
rect 492 290 526 318
rect 492 284 526 290
rect 492 222 526 246
rect 492 212 526 222
rect 492 154 526 174
rect 492 140 526 154
rect 1510 664 1544 678
rect 1510 644 1544 664
rect 1510 596 1544 606
rect 1510 572 1544 596
rect 1510 528 1544 534
rect 1510 500 1544 528
rect 1510 460 1544 462
rect 1510 428 1544 460
rect 1510 358 1544 390
rect 1510 356 1544 358
rect 1510 290 1544 318
rect 1510 284 1544 290
rect 1510 222 1544 246
rect 1510 212 1544 222
rect 1510 154 1544 174
rect 1510 140 1544 154
rect 2528 664 2562 678
rect 2528 644 2562 664
rect 2528 596 2562 606
rect 2528 572 2562 596
rect 2528 528 2562 534
rect 2528 500 2562 528
rect 2528 460 2562 462
rect 2528 428 2562 460
rect 2528 358 2562 390
rect 2528 356 2562 358
rect 2528 290 2562 318
rect 2528 284 2562 290
rect 2528 222 2562 246
rect 2528 212 2562 222
rect 2528 154 2562 174
rect 2528 140 2562 154
rect 3546 664 3580 678
rect 3546 644 3580 664
rect 3546 596 3580 606
rect 3546 572 3580 596
rect 3546 528 3580 534
rect 3546 500 3580 528
rect 3546 460 3580 462
rect 3546 428 3580 460
rect 3546 358 3580 390
rect 3546 356 3580 358
rect 3546 290 3580 318
rect 3546 284 3580 290
rect 3546 222 3580 246
rect 3546 212 3580 222
rect 3546 154 3580 174
rect 3546 140 3580 154
rect 4564 664 4598 678
rect 4564 644 4598 664
rect 4564 596 4598 606
rect 4564 572 4598 596
rect 4564 528 4598 534
rect 4564 500 4598 528
rect 4564 460 4598 462
rect 4564 428 4598 460
rect 4564 358 4598 390
rect 4564 356 4598 358
rect 4564 290 4598 318
rect 4564 284 4598 290
rect 4564 222 4598 246
rect 4564 212 4598 222
rect 4564 154 4598 174
rect 4564 140 4598 154
rect -4269 37 -4259 71
rect -4259 37 -4235 71
rect -4197 37 -4191 71
rect -4191 37 -4163 71
rect -4125 37 -4123 71
rect -4123 37 -4091 71
rect -4053 37 -4021 71
rect -4021 37 -4019 71
rect -3981 37 -3953 71
rect -3953 37 -3947 71
rect -3909 37 -3885 71
rect -3885 37 -3875 71
rect -3251 37 -3241 71
rect -3241 37 -3217 71
rect -3179 37 -3173 71
rect -3173 37 -3145 71
rect -3107 37 -3105 71
rect -3105 37 -3073 71
rect -3035 37 -3003 71
rect -3003 37 -3001 71
rect -2963 37 -2935 71
rect -2935 37 -2929 71
rect -2891 37 -2867 71
rect -2867 37 -2857 71
rect -2233 37 -2223 71
rect -2223 37 -2199 71
rect -2161 37 -2155 71
rect -2155 37 -2127 71
rect -2089 37 -2087 71
rect -2087 37 -2055 71
rect -2017 37 -1985 71
rect -1985 37 -1983 71
rect -1945 37 -1917 71
rect -1917 37 -1911 71
rect -1873 37 -1849 71
rect -1849 37 -1839 71
rect -1215 37 -1205 71
rect -1205 37 -1181 71
rect -1143 37 -1137 71
rect -1137 37 -1109 71
rect -1071 37 -1069 71
rect -1069 37 -1037 71
rect -999 37 -967 71
rect -967 37 -965 71
rect -927 37 -899 71
rect -899 37 -893 71
rect -855 37 -831 71
rect -831 37 -821 71
rect -197 37 -187 71
rect -187 37 -163 71
rect -125 37 -119 71
rect -119 37 -91 71
rect -53 37 -51 71
rect -51 37 -19 71
rect 19 37 51 71
rect 51 37 53 71
rect 91 37 119 71
rect 119 37 125 71
rect 163 37 187 71
rect 187 37 197 71
rect 821 37 831 71
rect 831 37 855 71
rect 893 37 899 71
rect 899 37 927 71
rect 965 37 967 71
rect 967 37 999 71
rect 1037 37 1069 71
rect 1069 37 1071 71
rect 1109 37 1137 71
rect 1137 37 1143 71
rect 1181 37 1205 71
rect 1205 37 1215 71
rect 1839 37 1849 71
rect 1849 37 1873 71
rect 1911 37 1917 71
rect 1917 37 1945 71
rect 1983 37 1985 71
rect 1985 37 2017 71
rect 2055 37 2087 71
rect 2087 37 2089 71
rect 2127 37 2155 71
rect 2155 37 2161 71
rect 2199 37 2223 71
rect 2223 37 2233 71
rect 2857 37 2867 71
rect 2867 37 2891 71
rect 2929 37 2935 71
rect 2935 37 2963 71
rect 3001 37 3003 71
rect 3003 37 3035 71
rect 3073 37 3105 71
rect 3105 37 3107 71
rect 3145 37 3173 71
rect 3173 37 3179 71
rect 3217 37 3241 71
rect 3241 37 3251 71
rect 3875 37 3885 71
rect 3885 37 3909 71
rect 3947 37 3953 71
rect 3953 37 3981 71
rect 4019 37 4021 71
rect 4021 37 4053 71
rect 4091 37 4123 71
rect 4123 37 4125 71
rect 4163 37 4191 71
rect 4191 37 4197 71
rect 4235 37 4259 71
rect 4259 37 4269 71
rect -4269 -71 -4259 -37
rect -4259 -71 -4235 -37
rect -4197 -71 -4191 -37
rect -4191 -71 -4163 -37
rect -4125 -71 -4123 -37
rect -4123 -71 -4091 -37
rect -4053 -71 -4021 -37
rect -4021 -71 -4019 -37
rect -3981 -71 -3953 -37
rect -3953 -71 -3947 -37
rect -3909 -71 -3885 -37
rect -3885 -71 -3875 -37
rect -3251 -71 -3241 -37
rect -3241 -71 -3217 -37
rect -3179 -71 -3173 -37
rect -3173 -71 -3145 -37
rect -3107 -71 -3105 -37
rect -3105 -71 -3073 -37
rect -3035 -71 -3003 -37
rect -3003 -71 -3001 -37
rect -2963 -71 -2935 -37
rect -2935 -71 -2929 -37
rect -2891 -71 -2867 -37
rect -2867 -71 -2857 -37
rect -2233 -71 -2223 -37
rect -2223 -71 -2199 -37
rect -2161 -71 -2155 -37
rect -2155 -71 -2127 -37
rect -2089 -71 -2087 -37
rect -2087 -71 -2055 -37
rect -2017 -71 -1985 -37
rect -1985 -71 -1983 -37
rect -1945 -71 -1917 -37
rect -1917 -71 -1911 -37
rect -1873 -71 -1849 -37
rect -1849 -71 -1839 -37
rect -1215 -71 -1205 -37
rect -1205 -71 -1181 -37
rect -1143 -71 -1137 -37
rect -1137 -71 -1109 -37
rect -1071 -71 -1069 -37
rect -1069 -71 -1037 -37
rect -999 -71 -967 -37
rect -967 -71 -965 -37
rect -927 -71 -899 -37
rect -899 -71 -893 -37
rect -855 -71 -831 -37
rect -831 -71 -821 -37
rect -197 -71 -187 -37
rect -187 -71 -163 -37
rect -125 -71 -119 -37
rect -119 -71 -91 -37
rect -53 -71 -51 -37
rect -51 -71 -19 -37
rect 19 -71 51 -37
rect 51 -71 53 -37
rect 91 -71 119 -37
rect 119 -71 125 -37
rect 163 -71 187 -37
rect 187 -71 197 -37
rect 821 -71 831 -37
rect 831 -71 855 -37
rect 893 -71 899 -37
rect 899 -71 927 -37
rect 965 -71 967 -37
rect 967 -71 999 -37
rect 1037 -71 1069 -37
rect 1069 -71 1071 -37
rect 1109 -71 1137 -37
rect 1137 -71 1143 -37
rect 1181 -71 1205 -37
rect 1205 -71 1215 -37
rect 1839 -71 1849 -37
rect 1849 -71 1873 -37
rect 1911 -71 1917 -37
rect 1917 -71 1945 -37
rect 1983 -71 1985 -37
rect 1985 -71 2017 -37
rect 2055 -71 2087 -37
rect 2087 -71 2089 -37
rect 2127 -71 2155 -37
rect 2155 -71 2161 -37
rect 2199 -71 2223 -37
rect 2223 -71 2233 -37
rect 2857 -71 2867 -37
rect 2867 -71 2891 -37
rect 2929 -71 2935 -37
rect 2935 -71 2963 -37
rect 3001 -71 3003 -37
rect 3003 -71 3035 -37
rect 3073 -71 3105 -37
rect 3105 -71 3107 -37
rect 3145 -71 3173 -37
rect 3173 -71 3179 -37
rect 3217 -71 3241 -37
rect 3241 -71 3251 -37
rect 3875 -71 3885 -37
rect 3885 -71 3909 -37
rect 3947 -71 3953 -37
rect 3953 -71 3981 -37
rect 4019 -71 4021 -37
rect 4021 -71 4053 -37
rect 4091 -71 4123 -37
rect 4123 -71 4125 -37
rect 4163 -71 4191 -37
rect 4191 -71 4197 -37
rect 4235 -71 4259 -37
rect 4259 -71 4269 -37
rect -4598 -154 -4564 -140
rect -4598 -174 -4564 -154
rect -4598 -222 -4564 -212
rect -4598 -246 -4564 -222
rect -4598 -290 -4564 -284
rect -4598 -318 -4564 -290
rect -4598 -358 -4564 -356
rect -4598 -390 -4564 -358
rect -4598 -460 -4564 -428
rect -4598 -462 -4564 -460
rect -4598 -528 -4564 -500
rect -4598 -534 -4564 -528
rect -4598 -596 -4564 -572
rect -4598 -606 -4564 -596
rect -4598 -664 -4564 -644
rect -4598 -678 -4564 -664
rect -3580 -154 -3546 -140
rect -3580 -174 -3546 -154
rect -3580 -222 -3546 -212
rect -3580 -246 -3546 -222
rect -3580 -290 -3546 -284
rect -3580 -318 -3546 -290
rect -3580 -358 -3546 -356
rect -3580 -390 -3546 -358
rect -3580 -460 -3546 -428
rect -3580 -462 -3546 -460
rect -3580 -528 -3546 -500
rect -3580 -534 -3546 -528
rect -3580 -596 -3546 -572
rect -3580 -606 -3546 -596
rect -3580 -664 -3546 -644
rect -3580 -678 -3546 -664
rect -2562 -154 -2528 -140
rect -2562 -174 -2528 -154
rect -2562 -222 -2528 -212
rect -2562 -246 -2528 -222
rect -2562 -290 -2528 -284
rect -2562 -318 -2528 -290
rect -2562 -358 -2528 -356
rect -2562 -390 -2528 -358
rect -2562 -460 -2528 -428
rect -2562 -462 -2528 -460
rect -2562 -528 -2528 -500
rect -2562 -534 -2528 -528
rect -2562 -596 -2528 -572
rect -2562 -606 -2528 -596
rect -2562 -664 -2528 -644
rect -2562 -678 -2528 -664
rect -1544 -154 -1510 -140
rect -1544 -174 -1510 -154
rect -1544 -222 -1510 -212
rect -1544 -246 -1510 -222
rect -1544 -290 -1510 -284
rect -1544 -318 -1510 -290
rect -1544 -358 -1510 -356
rect -1544 -390 -1510 -358
rect -1544 -460 -1510 -428
rect -1544 -462 -1510 -460
rect -1544 -528 -1510 -500
rect -1544 -534 -1510 -528
rect -1544 -596 -1510 -572
rect -1544 -606 -1510 -596
rect -1544 -664 -1510 -644
rect -1544 -678 -1510 -664
rect -526 -154 -492 -140
rect -526 -174 -492 -154
rect -526 -222 -492 -212
rect -526 -246 -492 -222
rect -526 -290 -492 -284
rect -526 -318 -492 -290
rect -526 -358 -492 -356
rect -526 -390 -492 -358
rect -526 -460 -492 -428
rect -526 -462 -492 -460
rect -526 -528 -492 -500
rect -526 -534 -492 -528
rect -526 -596 -492 -572
rect -526 -606 -492 -596
rect -526 -664 -492 -644
rect -526 -678 -492 -664
rect 492 -154 526 -140
rect 492 -174 526 -154
rect 492 -222 526 -212
rect 492 -246 526 -222
rect 492 -290 526 -284
rect 492 -318 526 -290
rect 492 -358 526 -356
rect 492 -390 526 -358
rect 492 -460 526 -428
rect 492 -462 526 -460
rect 492 -528 526 -500
rect 492 -534 526 -528
rect 492 -596 526 -572
rect 492 -606 526 -596
rect 492 -664 526 -644
rect 492 -678 526 -664
rect 1510 -154 1544 -140
rect 1510 -174 1544 -154
rect 1510 -222 1544 -212
rect 1510 -246 1544 -222
rect 1510 -290 1544 -284
rect 1510 -318 1544 -290
rect 1510 -358 1544 -356
rect 1510 -390 1544 -358
rect 1510 -460 1544 -428
rect 1510 -462 1544 -460
rect 1510 -528 1544 -500
rect 1510 -534 1544 -528
rect 1510 -596 1544 -572
rect 1510 -606 1544 -596
rect 1510 -664 1544 -644
rect 1510 -678 1544 -664
rect 2528 -154 2562 -140
rect 2528 -174 2562 -154
rect 2528 -222 2562 -212
rect 2528 -246 2562 -222
rect 2528 -290 2562 -284
rect 2528 -318 2562 -290
rect 2528 -358 2562 -356
rect 2528 -390 2562 -358
rect 2528 -460 2562 -428
rect 2528 -462 2562 -460
rect 2528 -528 2562 -500
rect 2528 -534 2562 -528
rect 2528 -596 2562 -572
rect 2528 -606 2562 -596
rect 2528 -664 2562 -644
rect 2528 -678 2562 -664
rect 3546 -154 3580 -140
rect 3546 -174 3580 -154
rect 3546 -222 3580 -212
rect 3546 -246 3580 -222
rect 3546 -290 3580 -284
rect 3546 -318 3580 -290
rect 3546 -358 3580 -356
rect 3546 -390 3580 -358
rect 3546 -460 3580 -428
rect 3546 -462 3580 -460
rect 3546 -528 3580 -500
rect 3546 -534 3580 -528
rect 3546 -596 3580 -572
rect 3546 -606 3580 -596
rect 3546 -664 3580 -644
rect 3546 -678 3580 -664
rect 4564 -154 4598 -140
rect 4564 -174 4598 -154
rect 4564 -222 4598 -212
rect 4564 -246 4598 -222
rect 4564 -290 4598 -284
rect 4564 -318 4598 -290
rect 4564 -358 4598 -356
rect 4564 -390 4598 -358
rect 4564 -460 4598 -428
rect 4564 -462 4598 -460
rect 4564 -528 4598 -500
rect 4564 -534 4598 -528
rect 4564 -596 4598 -572
rect 4564 -606 4598 -596
rect 4564 -664 4598 -644
rect 4564 -678 4598 -664
rect -4269 -781 -4259 -747
rect -4259 -781 -4235 -747
rect -4197 -781 -4191 -747
rect -4191 -781 -4163 -747
rect -4125 -781 -4123 -747
rect -4123 -781 -4091 -747
rect -4053 -781 -4021 -747
rect -4021 -781 -4019 -747
rect -3981 -781 -3953 -747
rect -3953 -781 -3947 -747
rect -3909 -781 -3885 -747
rect -3885 -781 -3875 -747
rect -3251 -781 -3241 -747
rect -3241 -781 -3217 -747
rect -3179 -781 -3173 -747
rect -3173 -781 -3145 -747
rect -3107 -781 -3105 -747
rect -3105 -781 -3073 -747
rect -3035 -781 -3003 -747
rect -3003 -781 -3001 -747
rect -2963 -781 -2935 -747
rect -2935 -781 -2929 -747
rect -2891 -781 -2867 -747
rect -2867 -781 -2857 -747
rect -2233 -781 -2223 -747
rect -2223 -781 -2199 -747
rect -2161 -781 -2155 -747
rect -2155 -781 -2127 -747
rect -2089 -781 -2087 -747
rect -2087 -781 -2055 -747
rect -2017 -781 -1985 -747
rect -1985 -781 -1983 -747
rect -1945 -781 -1917 -747
rect -1917 -781 -1911 -747
rect -1873 -781 -1849 -747
rect -1849 -781 -1839 -747
rect -1215 -781 -1205 -747
rect -1205 -781 -1181 -747
rect -1143 -781 -1137 -747
rect -1137 -781 -1109 -747
rect -1071 -781 -1069 -747
rect -1069 -781 -1037 -747
rect -999 -781 -967 -747
rect -967 -781 -965 -747
rect -927 -781 -899 -747
rect -899 -781 -893 -747
rect -855 -781 -831 -747
rect -831 -781 -821 -747
rect -197 -781 -187 -747
rect -187 -781 -163 -747
rect -125 -781 -119 -747
rect -119 -781 -91 -747
rect -53 -781 -51 -747
rect -51 -781 -19 -747
rect 19 -781 51 -747
rect 51 -781 53 -747
rect 91 -781 119 -747
rect 119 -781 125 -747
rect 163 -781 187 -747
rect 187 -781 197 -747
rect 821 -781 831 -747
rect 831 -781 855 -747
rect 893 -781 899 -747
rect 899 -781 927 -747
rect 965 -781 967 -747
rect 967 -781 999 -747
rect 1037 -781 1069 -747
rect 1069 -781 1071 -747
rect 1109 -781 1137 -747
rect 1137 -781 1143 -747
rect 1181 -781 1205 -747
rect 1205 -781 1215 -747
rect 1839 -781 1849 -747
rect 1849 -781 1873 -747
rect 1911 -781 1917 -747
rect 1917 -781 1945 -747
rect 1983 -781 1985 -747
rect 1985 -781 2017 -747
rect 2055 -781 2087 -747
rect 2087 -781 2089 -747
rect 2127 -781 2155 -747
rect 2155 -781 2161 -747
rect 2199 -781 2223 -747
rect 2223 -781 2233 -747
rect 2857 -781 2867 -747
rect 2867 -781 2891 -747
rect 2929 -781 2935 -747
rect 2935 -781 2963 -747
rect 3001 -781 3003 -747
rect 3003 -781 3035 -747
rect 3073 -781 3105 -747
rect 3105 -781 3107 -747
rect 3145 -781 3173 -747
rect 3173 -781 3179 -747
rect 3217 -781 3241 -747
rect 3241 -781 3251 -747
rect 3875 -781 3885 -747
rect 3885 -781 3909 -747
rect 3947 -781 3953 -747
rect 3953 -781 3981 -747
rect 4019 -781 4021 -747
rect 4021 -781 4053 -747
rect 4091 -781 4123 -747
rect 4123 -781 4125 -747
rect 4163 -781 4191 -747
rect 4191 -781 4197 -747
rect 4235 -781 4259 -747
rect 4259 -781 4269 -747
rect -4269 -889 -4259 -855
rect -4259 -889 -4235 -855
rect -4197 -889 -4191 -855
rect -4191 -889 -4163 -855
rect -4125 -889 -4123 -855
rect -4123 -889 -4091 -855
rect -4053 -889 -4021 -855
rect -4021 -889 -4019 -855
rect -3981 -889 -3953 -855
rect -3953 -889 -3947 -855
rect -3909 -889 -3885 -855
rect -3885 -889 -3875 -855
rect -3251 -889 -3241 -855
rect -3241 -889 -3217 -855
rect -3179 -889 -3173 -855
rect -3173 -889 -3145 -855
rect -3107 -889 -3105 -855
rect -3105 -889 -3073 -855
rect -3035 -889 -3003 -855
rect -3003 -889 -3001 -855
rect -2963 -889 -2935 -855
rect -2935 -889 -2929 -855
rect -2891 -889 -2867 -855
rect -2867 -889 -2857 -855
rect -2233 -889 -2223 -855
rect -2223 -889 -2199 -855
rect -2161 -889 -2155 -855
rect -2155 -889 -2127 -855
rect -2089 -889 -2087 -855
rect -2087 -889 -2055 -855
rect -2017 -889 -1985 -855
rect -1985 -889 -1983 -855
rect -1945 -889 -1917 -855
rect -1917 -889 -1911 -855
rect -1873 -889 -1849 -855
rect -1849 -889 -1839 -855
rect -1215 -889 -1205 -855
rect -1205 -889 -1181 -855
rect -1143 -889 -1137 -855
rect -1137 -889 -1109 -855
rect -1071 -889 -1069 -855
rect -1069 -889 -1037 -855
rect -999 -889 -967 -855
rect -967 -889 -965 -855
rect -927 -889 -899 -855
rect -899 -889 -893 -855
rect -855 -889 -831 -855
rect -831 -889 -821 -855
rect -197 -889 -187 -855
rect -187 -889 -163 -855
rect -125 -889 -119 -855
rect -119 -889 -91 -855
rect -53 -889 -51 -855
rect -51 -889 -19 -855
rect 19 -889 51 -855
rect 51 -889 53 -855
rect 91 -889 119 -855
rect 119 -889 125 -855
rect 163 -889 187 -855
rect 187 -889 197 -855
rect 821 -889 831 -855
rect 831 -889 855 -855
rect 893 -889 899 -855
rect 899 -889 927 -855
rect 965 -889 967 -855
rect 967 -889 999 -855
rect 1037 -889 1069 -855
rect 1069 -889 1071 -855
rect 1109 -889 1137 -855
rect 1137 -889 1143 -855
rect 1181 -889 1205 -855
rect 1205 -889 1215 -855
rect 1839 -889 1849 -855
rect 1849 -889 1873 -855
rect 1911 -889 1917 -855
rect 1917 -889 1945 -855
rect 1983 -889 1985 -855
rect 1985 -889 2017 -855
rect 2055 -889 2087 -855
rect 2087 -889 2089 -855
rect 2127 -889 2155 -855
rect 2155 -889 2161 -855
rect 2199 -889 2223 -855
rect 2223 -889 2233 -855
rect 2857 -889 2867 -855
rect 2867 -889 2891 -855
rect 2929 -889 2935 -855
rect 2935 -889 2963 -855
rect 3001 -889 3003 -855
rect 3003 -889 3035 -855
rect 3073 -889 3105 -855
rect 3105 -889 3107 -855
rect 3145 -889 3173 -855
rect 3173 -889 3179 -855
rect 3217 -889 3241 -855
rect 3241 -889 3251 -855
rect 3875 -889 3885 -855
rect 3885 -889 3909 -855
rect 3947 -889 3953 -855
rect 3953 -889 3981 -855
rect 4019 -889 4021 -855
rect 4021 -889 4053 -855
rect 4091 -889 4123 -855
rect 4123 -889 4125 -855
rect 4163 -889 4191 -855
rect 4191 -889 4197 -855
rect 4235 -889 4259 -855
rect 4259 -889 4269 -855
rect -4598 -972 -4564 -958
rect -4598 -992 -4564 -972
rect -4598 -1040 -4564 -1030
rect -4598 -1064 -4564 -1040
rect -4598 -1108 -4564 -1102
rect -4598 -1136 -4564 -1108
rect -4598 -1176 -4564 -1174
rect -4598 -1208 -4564 -1176
rect -4598 -1278 -4564 -1246
rect -4598 -1280 -4564 -1278
rect -4598 -1346 -4564 -1318
rect -4598 -1352 -4564 -1346
rect -4598 -1414 -4564 -1390
rect -4598 -1424 -4564 -1414
rect -4598 -1482 -4564 -1462
rect -4598 -1496 -4564 -1482
rect -3580 -972 -3546 -958
rect -3580 -992 -3546 -972
rect -3580 -1040 -3546 -1030
rect -3580 -1064 -3546 -1040
rect -3580 -1108 -3546 -1102
rect -3580 -1136 -3546 -1108
rect -3580 -1176 -3546 -1174
rect -3580 -1208 -3546 -1176
rect -3580 -1278 -3546 -1246
rect -3580 -1280 -3546 -1278
rect -3580 -1346 -3546 -1318
rect -3580 -1352 -3546 -1346
rect -3580 -1414 -3546 -1390
rect -3580 -1424 -3546 -1414
rect -3580 -1482 -3546 -1462
rect -3580 -1496 -3546 -1482
rect -2562 -972 -2528 -958
rect -2562 -992 -2528 -972
rect -2562 -1040 -2528 -1030
rect -2562 -1064 -2528 -1040
rect -2562 -1108 -2528 -1102
rect -2562 -1136 -2528 -1108
rect -2562 -1176 -2528 -1174
rect -2562 -1208 -2528 -1176
rect -2562 -1278 -2528 -1246
rect -2562 -1280 -2528 -1278
rect -2562 -1346 -2528 -1318
rect -2562 -1352 -2528 -1346
rect -2562 -1414 -2528 -1390
rect -2562 -1424 -2528 -1414
rect -2562 -1482 -2528 -1462
rect -2562 -1496 -2528 -1482
rect -1544 -972 -1510 -958
rect -1544 -992 -1510 -972
rect -1544 -1040 -1510 -1030
rect -1544 -1064 -1510 -1040
rect -1544 -1108 -1510 -1102
rect -1544 -1136 -1510 -1108
rect -1544 -1176 -1510 -1174
rect -1544 -1208 -1510 -1176
rect -1544 -1278 -1510 -1246
rect -1544 -1280 -1510 -1278
rect -1544 -1346 -1510 -1318
rect -1544 -1352 -1510 -1346
rect -1544 -1414 -1510 -1390
rect -1544 -1424 -1510 -1414
rect -1544 -1482 -1510 -1462
rect -1544 -1496 -1510 -1482
rect -526 -972 -492 -958
rect -526 -992 -492 -972
rect -526 -1040 -492 -1030
rect -526 -1064 -492 -1040
rect -526 -1108 -492 -1102
rect -526 -1136 -492 -1108
rect -526 -1176 -492 -1174
rect -526 -1208 -492 -1176
rect -526 -1278 -492 -1246
rect -526 -1280 -492 -1278
rect -526 -1346 -492 -1318
rect -526 -1352 -492 -1346
rect -526 -1414 -492 -1390
rect -526 -1424 -492 -1414
rect -526 -1482 -492 -1462
rect -526 -1496 -492 -1482
rect 492 -972 526 -958
rect 492 -992 526 -972
rect 492 -1040 526 -1030
rect 492 -1064 526 -1040
rect 492 -1108 526 -1102
rect 492 -1136 526 -1108
rect 492 -1176 526 -1174
rect 492 -1208 526 -1176
rect 492 -1278 526 -1246
rect 492 -1280 526 -1278
rect 492 -1346 526 -1318
rect 492 -1352 526 -1346
rect 492 -1414 526 -1390
rect 492 -1424 526 -1414
rect 492 -1482 526 -1462
rect 492 -1496 526 -1482
rect 1510 -972 1544 -958
rect 1510 -992 1544 -972
rect 1510 -1040 1544 -1030
rect 1510 -1064 1544 -1040
rect 1510 -1108 1544 -1102
rect 1510 -1136 1544 -1108
rect 1510 -1176 1544 -1174
rect 1510 -1208 1544 -1176
rect 1510 -1278 1544 -1246
rect 1510 -1280 1544 -1278
rect 1510 -1346 1544 -1318
rect 1510 -1352 1544 -1346
rect 1510 -1414 1544 -1390
rect 1510 -1424 1544 -1414
rect 1510 -1482 1544 -1462
rect 1510 -1496 1544 -1482
rect 2528 -972 2562 -958
rect 2528 -992 2562 -972
rect 2528 -1040 2562 -1030
rect 2528 -1064 2562 -1040
rect 2528 -1108 2562 -1102
rect 2528 -1136 2562 -1108
rect 2528 -1176 2562 -1174
rect 2528 -1208 2562 -1176
rect 2528 -1278 2562 -1246
rect 2528 -1280 2562 -1278
rect 2528 -1346 2562 -1318
rect 2528 -1352 2562 -1346
rect 2528 -1414 2562 -1390
rect 2528 -1424 2562 -1414
rect 2528 -1482 2562 -1462
rect 2528 -1496 2562 -1482
rect 3546 -972 3580 -958
rect 3546 -992 3580 -972
rect 3546 -1040 3580 -1030
rect 3546 -1064 3580 -1040
rect 3546 -1108 3580 -1102
rect 3546 -1136 3580 -1108
rect 3546 -1176 3580 -1174
rect 3546 -1208 3580 -1176
rect 3546 -1278 3580 -1246
rect 3546 -1280 3580 -1278
rect 3546 -1346 3580 -1318
rect 3546 -1352 3580 -1346
rect 3546 -1414 3580 -1390
rect 3546 -1424 3580 -1414
rect 3546 -1482 3580 -1462
rect 3546 -1496 3580 -1482
rect 4564 -972 4598 -958
rect 4564 -992 4598 -972
rect 4564 -1040 4598 -1030
rect 4564 -1064 4598 -1040
rect 4564 -1108 4598 -1102
rect 4564 -1136 4598 -1108
rect 4564 -1176 4598 -1174
rect 4564 -1208 4598 -1176
rect 4564 -1278 4598 -1246
rect 4564 -1280 4598 -1278
rect 4564 -1346 4598 -1318
rect 4564 -1352 4598 -1346
rect 4564 -1414 4598 -1390
rect 4564 -1424 4598 -1414
rect 4564 -1482 4598 -1462
rect 4564 -1496 4598 -1482
rect -4269 -1599 -4259 -1565
rect -4259 -1599 -4235 -1565
rect -4197 -1599 -4191 -1565
rect -4191 -1599 -4163 -1565
rect -4125 -1599 -4123 -1565
rect -4123 -1599 -4091 -1565
rect -4053 -1599 -4021 -1565
rect -4021 -1599 -4019 -1565
rect -3981 -1599 -3953 -1565
rect -3953 -1599 -3947 -1565
rect -3909 -1599 -3885 -1565
rect -3885 -1599 -3875 -1565
rect -3251 -1599 -3241 -1565
rect -3241 -1599 -3217 -1565
rect -3179 -1599 -3173 -1565
rect -3173 -1599 -3145 -1565
rect -3107 -1599 -3105 -1565
rect -3105 -1599 -3073 -1565
rect -3035 -1599 -3003 -1565
rect -3003 -1599 -3001 -1565
rect -2963 -1599 -2935 -1565
rect -2935 -1599 -2929 -1565
rect -2891 -1599 -2867 -1565
rect -2867 -1599 -2857 -1565
rect -2233 -1599 -2223 -1565
rect -2223 -1599 -2199 -1565
rect -2161 -1599 -2155 -1565
rect -2155 -1599 -2127 -1565
rect -2089 -1599 -2087 -1565
rect -2087 -1599 -2055 -1565
rect -2017 -1599 -1985 -1565
rect -1985 -1599 -1983 -1565
rect -1945 -1599 -1917 -1565
rect -1917 -1599 -1911 -1565
rect -1873 -1599 -1849 -1565
rect -1849 -1599 -1839 -1565
rect -1215 -1599 -1205 -1565
rect -1205 -1599 -1181 -1565
rect -1143 -1599 -1137 -1565
rect -1137 -1599 -1109 -1565
rect -1071 -1599 -1069 -1565
rect -1069 -1599 -1037 -1565
rect -999 -1599 -967 -1565
rect -967 -1599 -965 -1565
rect -927 -1599 -899 -1565
rect -899 -1599 -893 -1565
rect -855 -1599 -831 -1565
rect -831 -1599 -821 -1565
rect -197 -1599 -187 -1565
rect -187 -1599 -163 -1565
rect -125 -1599 -119 -1565
rect -119 -1599 -91 -1565
rect -53 -1599 -51 -1565
rect -51 -1599 -19 -1565
rect 19 -1599 51 -1565
rect 51 -1599 53 -1565
rect 91 -1599 119 -1565
rect 119 -1599 125 -1565
rect 163 -1599 187 -1565
rect 187 -1599 197 -1565
rect 821 -1599 831 -1565
rect 831 -1599 855 -1565
rect 893 -1599 899 -1565
rect 899 -1599 927 -1565
rect 965 -1599 967 -1565
rect 967 -1599 999 -1565
rect 1037 -1599 1069 -1565
rect 1069 -1599 1071 -1565
rect 1109 -1599 1137 -1565
rect 1137 -1599 1143 -1565
rect 1181 -1599 1205 -1565
rect 1205 -1599 1215 -1565
rect 1839 -1599 1849 -1565
rect 1849 -1599 1873 -1565
rect 1911 -1599 1917 -1565
rect 1917 -1599 1945 -1565
rect 1983 -1599 1985 -1565
rect 1985 -1599 2017 -1565
rect 2055 -1599 2087 -1565
rect 2087 -1599 2089 -1565
rect 2127 -1599 2155 -1565
rect 2155 -1599 2161 -1565
rect 2199 -1599 2223 -1565
rect 2223 -1599 2233 -1565
rect 2857 -1599 2867 -1565
rect 2867 -1599 2891 -1565
rect 2929 -1599 2935 -1565
rect 2935 -1599 2963 -1565
rect 3001 -1599 3003 -1565
rect 3003 -1599 3035 -1565
rect 3073 -1599 3105 -1565
rect 3105 -1599 3107 -1565
rect 3145 -1599 3173 -1565
rect 3173 -1599 3179 -1565
rect 3217 -1599 3241 -1565
rect 3241 -1599 3251 -1565
rect 3875 -1599 3885 -1565
rect 3885 -1599 3909 -1565
rect 3947 -1599 3953 -1565
rect 3953 -1599 3981 -1565
rect 4019 -1599 4021 -1565
rect 4021 -1599 4053 -1565
rect 4091 -1599 4123 -1565
rect 4123 -1599 4125 -1565
rect 4163 -1599 4191 -1565
rect 4191 -1599 4197 -1565
rect 4235 -1599 4259 -1565
rect 4259 -1599 4269 -1565
<< metal1 >>
rect -4316 1599 -3828 1605
rect -4316 1565 -4269 1599
rect -4235 1565 -4197 1599
rect -4163 1565 -4125 1599
rect -4091 1565 -4053 1599
rect -4019 1565 -3981 1599
rect -3947 1565 -3909 1599
rect -3875 1565 -3828 1599
rect -4316 1559 -3828 1565
rect -3298 1599 -2810 1605
rect -3298 1565 -3251 1599
rect -3217 1565 -3179 1599
rect -3145 1565 -3107 1599
rect -3073 1565 -3035 1599
rect -3001 1565 -2963 1599
rect -2929 1565 -2891 1599
rect -2857 1565 -2810 1599
rect -3298 1559 -2810 1565
rect -2280 1599 -1792 1605
rect -2280 1565 -2233 1599
rect -2199 1565 -2161 1599
rect -2127 1565 -2089 1599
rect -2055 1565 -2017 1599
rect -1983 1565 -1945 1599
rect -1911 1565 -1873 1599
rect -1839 1565 -1792 1599
rect -2280 1559 -1792 1565
rect -1262 1599 -774 1605
rect -1262 1565 -1215 1599
rect -1181 1565 -1143 1599
rect -1109 1565 -1071 1599
rect -1037 1565 -999 1599
rect -965 1565 -927 1599
rect -893 1565 -855 1599
rect -821 1565 -774 1599
rect -1262 1559 -774 1565
rect -244 1599 244 1605
rect -244 1565 -197 1599
rect -163 1565 -125 1599
rect -91 1565 -53 1599
rect -19 1565 19 1599
rect 53 1565 91 1599
rect 125 1565 163 1599
rect 197 1565 244 1599
rect -244 1559 244 1565
rect 774 1599 1262 1605
rect 774 1565 821 1599
rect 855 1565 893 1599
rect 927 1565 965 1599
rect 999 1565 1037 1599
rect 1071 1565 1109 1599
rect 1143 1565 1181 1599
rect 1215 1565 1262 1599
rect 774 1559 1262 1565
rect 1792 1599 2280 1605
rect 1792 1565 1839 1599
rect 1873 1565 1911 1599
rect 1945 1565 1983 1599
rect 2017 1565 2055 1599
rect 2089 1565 2127 1599
rect 2161 1565 2199 1599
rect 2233 1565 2280 1599
rect 1792 1559 2280 1565
rect 2810 1599 3298 1605
rect 2810 1565 2857 1599
rect 2891 1565 2929 1599
rect 2963 1565 3001 1599
rect 3035 1565 3073 1599
rect 3107 1565 3145 1599
rect 3179 1565 3217 1599
rect 3251 1565 3298 1599
rect 2810 1559 3298 1565
rect 3828 1599 4316 1605
rect 3828 1565 3875 1599
rect 3909 1565 3947 1599
rect 3981 1565 4019 1599
rect 4053 1565 4091 1599
rect 4125 1565 4163 1599
rect 4197 1565 4235 1599
rect 4269 1565 4316 1599
rect 3828 1559 4316 1565
rect -4604 1496 -4558 1527
rect -4604 1462 -4598 1496
rect -4564 1462 -4558 1496
rect -4604 1424 -4558 1462
rect -4604 1390 -4598 1424
rect -4564 1390 -4558 1424
rect -4604 1352 -4558 1390
rect -4604 1318 -4598 1352
rect -4564 1318 -4558 1352
rect -4604 1280 -4558 1318
rect -4604 1246 -4598 1280
rect -4564 1246 -4558 1280
rect -4604 1208 -4558 1246
rect -4604 1174 -4598 1208
rect -4564 1174 -4558 1208
rect -4604 1136 -4558 1174
rect -4604 1102 -4598 1136
rect -4564 1102 -4558 1136
rect -4604 1064 -4558 1102
rect -4604 1030 -4598 1064
rect -4564 1030 -4558 1064
rect -4604 992 -4558 1030
rect -4604 958 -4598 992
rect -4564 958 -4558 992
rect -4604 927 -4558 958
rect -3586 1496 -3540 1527
rect -3586 1462 -3580 1496
rect -3546 1462 -3540 1496
rect -3586 1424 -3540 1462
rect -3586 1390 -3580 1424
rect -3546 1390 -3540 1424
rect -3586 1352 -3540 1390
rect -3586 1318 -3580 1352
rect -3546 1318 -3540 1352
rect -3586 1280 -3540 1318
rect -3586 1246 -3580 1280
rect -3546 1246 -3540 1280
rect -3586 1208 -3540 1246
rect -3586 1174 -3580 1208
rect -3546 1174 -3540 1208
rect -3586 1136 -3540 1174
rect -3586 1102 -3580 1136
rect -3546 1102 -3540 1136
rect -3586 1064 -3540 1102
rect -3586 1030 -3580 1064
rect -3546 1030 -3540 1064
rect -3586 992 -3540 1030
rect -3586 958 -3580 992
rect -3546 958 -3540 992
rect -3586 927 -3540 958
rect -2568 1496 -2522 1527
rect -2568 1462 -2562 1496
rect -2528 1462 -2522 1496
rect -2568 1424 -2522 1462
rect -2568 1390 -2562 1424
rect -2528 1390 -2522 1424
rect -2568 1352 -2522 1390
rect -2568 1318 -2562 1352
rect -2528 1318 -2522 1352
rect -2568 1280 -2522 1318
rect -2568 1246 -2562 1280
rect -2528 1246 -2522 1280
rect -2568 1208 -2522 1246
rect -2568 1174 -2562 1208
rect -2528 1174 -2522 1208
rect -2568 1136 -2522 1174
rect -2568 1102 -2562 1136
rect -2528 1102 -2522 1136
rect -2568 1064 -2522 1102
rect -2568 1030 -2562 1064
rect -2528 1030 -2522 1064
rect -2568 992 -2522 1030
rect -2568 958 -2562 992
rect -2528 958 -2522 992
rect -2568 927 -2522 958
rect -1550 1496 -1504 1527
rect -1550 1462 -1544 1496
rect -1510 1462 -1504 1496
rect -1550 1424 -1504 1462
rect -1550 1390 -1544 1424
rect -1510 1390 -1504 1424
rect -1550 1352 -1504 1390
rect -1550 1318 -1544 1352
rect -1510 1318 -1504 1352
rect -1550 1280 -1504 1318
rect -1550 1246 -1544 1280
rect -1510 1246 -1504 1280
rect -1550 1208 -1504 1246
rect -1550 1174 -1544 1208
rect -1510 1174 -1504 1208
rect -1550 1136 -1504 1174
rect -1550 1102 -1544 1136
rect -1510 1102 -1504 1136
rect -1550 1064 -1504 1102
rect -1550 1030 -1544 1064
rect -1510 1030 -1504 1064
rect -1550 992 -1504 1030
rect -1550 958 -1544 992
rect -1510 958 -1504 992
rect -1550 927 -1504 958
rect -532 1496 -486 1527
rect -532 1462 -526 1496
rect -492 1462 -486 1496
rect -532 1424 -486 1462
rect -532 1390 -526 1424
rect -492 1390 -486 1424
rect -532 1352 -486 1390
rect -532 1318 -526 1352
rect -492 1318 -486 1352
rect -532 1280 -486 1318
rect -532 1246 -526 1280
rect -492 1246 -486 1280
rect -532 1208 -486 1246
rect -532 1174 -526 1208
rect -492 1174 -486 1208
rect -532 1136 -486 1174
rect -532 1102 -526 1136
rect -492 1102 -486 1136
rect -532 1064 -486 1102
rect -532 1030 -526 1064
rect -492 1030 -486 1064
rect -532 992 -486 1030
rect -532 958 -526 992
rect -492 958 -486 992
rect -532 927 -486 958
rect 486 1496 532 1527
rect 486 1462 492 1496
rect 526 1462 532 1496
rect 486 1424 532 1462
rect 486 1390 492 1424
rect 526 1390 532 1424
rect 486 1352 532 1390
rect 486 1318 492 1352
rect 526 1318 532 1352
rect 486 1280 532 1318
rect 486 1246 492 1280
rect 526 1246 532 1280
rect 486 1208 532 1246
rect 486 1174 492 1208
rect 526 1174 532 1208
rect 486 1136 532 1174
rect 486 1102 492 1136
rect 526 1102 532 1136
rect 486 1064 532 1102
rect 486 1030 492 1064
rect 526 1030 532 1064
rect 486 992 532 1030
rect 486 958 492 992
rect 526 958 532 992
rect 486 927 532 958
rect 1504 1496 1550 1527
rect 1504 1462 1510 1496
rect 1544 1462 1550 1496
rect 1504 1424 1550 1462
rect 1504 1390 1510 1424
rect 1544 1390 1550 1424
rect 1504 1352 1550 1390
rect 1504 1318 1510 1352
rect 1544 1318 1550 1352
rect 1504 1280 1550 1318
rect 1504 1246 1510 1280
rect 1544 1246 1550 1280
rect 1504 1208 1550 1246
rect 1504 1174 1510 1208
rect 1544 1174 1550 1208
rect 1504 1136 1550 1174
rect 1504 1102 1510 1136
rect 1544 1102 1550 1136
rect 1504 1064 1550 1102
rect 1504 1030 1510 1064
rect 1544 1030 1550 1064
rect 1504 992 1550 1030
rect 1504 958 1510 992
rect 1544 958 1550 992
rect 1504 927 1550 958
rect 2522 1496 2568 1527
rect 2522 1462 2528 1496
rect 2562 1462 2568 1496
rect 2522 1424 2568 1462
rect 2522 1390 2528 1424
rect 2562 1390 2568 1424
rect 2522 1352 2568 1390
rect 2522 1318 2528 1352
rect 2562 1318 2568 1352
rect 2522 1280 2568 1318
rect 2522 1246 2528 1280
rect 2562 1246 2568 1280
rect 2522 1208 2568 1246
rect 2522 1174 2528 1208
rect 2562 1174 2568 1208
rect 2522 1136 2568 1174
rect 2522 1102 2528 1136
rect 2562 1102 2568 1136
rect 2522 1064 2568 1102
rect 2522 1030 2528 1064
rect 2562 1030 2568 1064
rect 2522 992 2568 1030
rect 2522 958 2528 992
rect 2562 958 2568 992
rect 2522 927 2568 958
rect 3540 1496 3586 1527
rect 3540 1462 3546 1496
rect 3580 1462 3586 1496
rect 3540 1424 3586 1462
rect 3540 1390 3546 1424
rect 3580 1390 3586 1424
rect 3540 1352 3586 1390
rect 3540 1318 3546 1352
rect 3580 1318 3586 1352
rect 3540 1280 3586 1318
rect 3540 1246 3546 1280
rect 3580 1246 3586 1280
rect 3540 1208 3586 1246
rect 3540 1174 3546 1208
rect 3580 1174 3586 1208
rect 3540 1136 3586 1174
rect 3540 1102 3546 1136
rect 3580 1102 3586 1136
rect 3540 1064 3586 1102
rect 3540 1030 3546 1064
rect 3580 1030 3586 1064
rect 3540 992 3586 1030
rect 3540 958 3546 992
rect 3580 958 3586 992
rect 3540 927 3586 958
rect 4558 1496 4604 1527
rect 4558 1462 4564 1496
rect 4598 1462 4604 1496
rect 4558 1424 4604 1462
rect 4558 1390 4564 1424
rect 4598 1390 4604 1424
rect 4558 1352 4604 1390
rect 4558 1318 4564 1352
rect 4598 1318 4604 1352
rect 4558 1280 4604 1318
rect 4558 1246 4564 1280
rect 4598 1246 4604 1280
rect 4558 1208 4604 1246
rect 4558 1174 4564 1208
rect 4598 1174 4604 1208
rect 4558 1136 4604 1174
rect 4558 1102 4564 1136
rect 4598 1102 4604 1136
rect 4558 1064 4604 1102
rect 4558 1030 4564 1064
rect 4598 1030 4604 1064
rect 4558 992 4604 1030
rect 4558 958 4564 992
rect 4598 958 4604 992
rect 4558 927 4604 958
rect -4316 889 -3828 895
rect -4316 855 -4269 889
rect -4235 855 -4197 889
rect -4163 855 -4125 889
rect -4091 855 -4053 889
rect -4019 855 -3981 889
rect -3947 855 -3909 889
rect -3875 855 -3828 889
rect -4316 849 -3828 855
rect -3298 889 -2810 895
rect -3298 855 -3251 889
rect -3217 855 -3179 889
rect -3145 855 -3107 889
rect -3073 855 -3035 889
rect -3001 855 -2963 889
rect -2929 855 -2891 889
rect -2857 855 -2810 889
rect -3298 849 -2810 855
rect -2280 889 -1792 895
rect -2280 855 -2233 889
rect -2199 855 -2161 889
rect -2127 855 -2089 889
rect -2055 855 -2017 889
rect -1983 855 -1945 889
rect -1911 855 -1873 889
rect -1839 855 -1792 889
rect -2280 849 -1792 855
rect -1262 889 -774 895
rect -1262 855 -1215 889
rect -1181 855 -1143 889
rect -1109 855 -1071 889
rect -1037 855 -999 889
rect -965 855 -927 889
rect -893 855 -855 889
rect -821 855 -774 889
rect -1262 849 -774 855
rect -244 889 244 895
rect -244 855 -197 889
rect -163 855 -125 889
rect -91 855 -53 889
rect -19 855 19 889
rect 53 855 91 889
rect 125 855 163 889
rect 197 855 244 889
rect -244 849 244 855
rect 774 889 1262 895
rect 774 855 821 889
rect 855 855 893 889
rect 927 855 965 889
rect 999 855 1037 889
rect 1071 855 1109 889
rect 1143 855 1181 889
rect 1215 855 1262 889
rect 774 849 1262 855
rect 1792 889 2280 895
rect 1792 855 1839 889
rect 1873 855 1911 889
rect 1945 855 1983 889
rect 2017 855 2055 889
rect 2089 855 2127 889
rect 2161 855 2199 889
rect 2233 855 2280 889
rect 1792 849 2280 855
rect 2810 889 3298 895
rect 2810 855 2857 889
rect 2891 855 2929 889
rect 2963 855 3001 889
rect 3035 855 3073 889
rect 3107 855 3145 889
rect 3179 855 3217 889
rect 3251 855 3298 889
rect 2810 849 3298 855
rect 3828 889 4316 895
rect 3828 855 3875 889
rect 3909 855 3947 889
rect 3981 855 4019 889
rect 4053 855 4091 889
rect 4125 855 4163 889
rect 4197 855 4235 889
rect 4269 855 4316 889
rect 3828 849 4316 855
rect -4316 781 -3828 787
rect -4316 747 -4269 781
rect -4235 747 -4197 781
rect -4163 747 -4125 781
rect -4091 747 -4053 781
rect -4019 747 -3981 781
rect -3947 747 -3909 781
rect -3875 747 -3828 781
rect -4316 741 -3828 747
rect -3298 781 -2810 787
rect -3298 747 -3251 781
rect -3217 747 -3179 781
rect -3145 747 -3107 781
rect -3073 747 -3035 781
rect -3001 747 -2963 781
rect -2929 747 -2891 781
rect -2857 747 -2810 781
rect -3298 741 -2810 747
rect -2280 781 -1792 787
rect -2280 747 -2233 781
rect -2199 747 -2161 781
rect -2127 747 -2089 781
rect -2055 747 -2017 781
rect -1983 747 -1945 781
rect -1911 747 -1873 781
rect -1839 747 -1792 781
rect -2280 741 -1792 747
rect -1262 781 -774 787
rect -1262 747 -1215 781
rect -1181 747 -1143 781
rect -1109 747 -1071 781
rect -1037 747 -999 781
rect -965 747 -927 781
rect -893 747 -855 781
rect -821 747 -774 781
rect -1262 741 -774 747
rect -244 781 244 787
rect -244 747 -197 781
rect -163 747 -125 781
rect -91 747 -53 781
rect -19 747 19 781
rect 53 747 91 781
rect 125 747 163 781
rect 197 747 244 781
rect -244 741 244 747
rect 774 781 1262 787
rect 774 747 821 781
rect 855 747 893 781
rect 927 747 965 781
rect 999 747 1037 781
rect 1071 747 1109 781
rect 1143 747 1181 781
rect 1215 747 1262 781
rect 774 741 1262 747
rect 1792 781 2280 787
rect 1792 747 1839 781
rect 1873 747 1911 781
rect 1945 747 1983 781
rect 2017 747 2055 781
rect 2089 747 2127 781
rect 2161 747 2199 781
rect 2233 747 2280 781
rect 1792 741 2280 747
rect 2810 781 3298 787
rect 2810 747 2857 781
rect 2891 747 2929 781
rect 2963 747 3001 781
rect 3035 747 3073 781
rect 3107 747 3145 781
rect 3179 747 3217 781
rect 3251 747 3298 781
rect 2810 741 3298 747
rect 3828 781 4316 787
rect 3828 747 3875 781
rect 3909 747 3947 781
rect 3981 747 4019 781
rect 4053 747 4091 781
rect 4125 747 4163 781
rect 4197 747 4235 781
rect 4269 747 4316 781
rect 3828 741 4316 747
rect -4604 678 -4558 709
rect -4604 644 -4598 678
rect -4564 644 -4558 678
rect -4604 606 -4558 644
rect -4604 572 -4598 606
rect -4564 572 -4558 606
rect -4604 534 -4558 572
rect -4604 500 -4598 534
rect -4564 500 -4558 534
rect -4604 462 -4558 500
rect -4604 428 -4598 462
rect -4564 428 -4558 462
rect -4604 390 -4558 428
rect -4604 356 -4598 390
rect -4564 356 -4558 390
rect -4604 318 -4558 356
rect -4604 284 -4598 318
rect -4564 284 -4558 318
rect -4604 246 -4558 284
rect -4604 212 -4598 246
rect -4564 212 -4558 246
rect -4604 174 -4558 212
rect -4604 140 -4598 174
rect -4564 140 -4558 174
rect -4604 109 -4558 140
rect -3586 678 -3540 709
rect -3586 644 -3580 678
rect -3546 644 -3540 678
rect -3586 606 -3540 644
rect -3586 572 -3580 606
rect -3546 572 -3540 606
rect -3586 534 -3540 572
rect -3586 500 -3580 534
rect -3546 500 -3540 534
rect -3586 462 -3540 500
rect -3586 428 -3580 462
rect -3546 428 -3540 462
rect -3586 390 -3540 428
rect -3586 356 -3580 390
rect -3546 356 -3540 390
rect -3586 318 -3540 356
rect -3586 284 -3580 318
rect -3546 284 -3540 318
rect -3586 246 -3540 284
rect -3586 212 -3580 246
rect -3546 212 -3540 246
rect -3586 174 -3540 212
rect -3586 140 -3580 174
rect -3546 140 -3540 174
rect -3586 109 -3540 140
rect -2568 678 -2522 709
rect -2568 644 -2562 678
rect -2528 644 -2522 678
rect -2568 606 -2522 644
rect -2568 572 -2562 606
rect -2528 572 -2522 606
rect -2568 534 -2522 572
rect -2568 500 -2562 534
rect -2528 500 -2522 534
rect -2568 462 -2522 500
rect -2568 428 -2562 462
rect -2528 428 -2522 462
rect -2568 390 -2522 428
rect -2568 356 -2562 390
rect -2528 356 -2522 390
rect -2568 318 -2522 356
rect -2568 284 -2562 318
rect -2528 284 -2522 318
rect -2568 246 -2522 284
rect -2568 212 -2562 246
rect -2528 212 -2522 246
rect -2568 174 -2522 212
rect -2568 140 -2562 174
rect -2528 140 -2522 174
rect -2568 109 -2522 140
rect -1550 678 -1504 709
rect -1550 644 -1544 678
rect -1510 644 -1504 678
rect -1550 606 -1504 644
rect -1550 572 -1544 606
rect -1510 572 -1504 606
rect -1550 534 -1504 572
rect -1550 500 -1544 534
rect -1510 500 -1504 534
rect -1550 462 -1504 500
rect -1550 428 -1544 462
rect -1510 428 -1504 462
rect -1550 390 -1504 428
rect -1550 356 -1544 390
rect -1510 356 -1504 390
rect -1550 318 -1504 356
rect -1550 284 -1544 318
rect -1510 284 -1504 318
rect -1550 246 -1504 284
rect -1550 212 -1544 246
rect -1510 212 -1504 246
rect -1550 174 -1504 212
rect -1550 140 -1544 174
rect -1510 140 -1504 174
rect -1550 109 -1504 140
rect -532 678 -486 709
rect -532 644 -526 678
rect -492 644 -486 678
rect -532 606 -486 644
rect -532 572 -526 606
rect -492 572 -486 606
rect -532 534 -486 572
rect -532 500 -526 534
rect -492 500 -486 534
rect -532 462 -486 500
rect -532 428 -526 462
rect -492 428 -486 462
rect -532 390 -486 428
rect -532 356 -526 390
rect -492 356 -486 390
rect -532 318 -486 356
rect -532 284 -526 318
rect -492 284 -486 318
rect -532 246 -486 284
rect -532 212 -526 246
rect -492 212 -486 246
rect -532 174 -486 212
rect -532 140 -526 174
rect -492 140 -486 174
rect -532 109 -486 140
rect 486 678 532 709
rect 486 644 492 678
rect 526 644 532 678
rect 486 606 532 644
rect 486 572 492 606
rect 526 572 532 606
rect 486 534 532 572
rect 486 500 492 534
rect 526 500 532 534
rect 486 462 532 500
rect 486 428 492 462
rect 526 428 532 462
rect 486 390 532 428
rect 486 356 492 390
rect 526 356 532 390
rect 486 318 532 356
rect 486 284 492 318
rect 526 284 532 318
rect 486 246 532 284
rect 486 212 492 246
rect 526 212 532 246
rect 486 174 532 212
rect 486 140 492 174
rect 526 140 532 174
rect 486 109 532 140
rect 1504 678 1550 709
rect 1504 644 1510 678
rect 1544 644 1550 678
rect 1504 606 1550 644
rect 1504 572 1510 606
rect 1544 572 1550 606
rect 1504 534 1550 572
rect 1504 500 1510 534
rect 1544 500 1550 534
rect 1504 462 1550 500
rect 1504 428 1510 462
rect 1544 428 1550 462
rect 1504 390 1550 428
rect 1504 356 1510 390
rect 1544 356 1550 390
rect 1504 318 1550 356
rect 1504 284 1510 318
rect 1544 284 1550 318
rect 1504 246 1550 284
rect 1504 212 1510 246
rect 1544 212 1550 246
rect 1504 174 1550 212
rect 1504 140 1510 174
rect 1544 140 1550 174
rect 1504 109 1550 140
rect 2522 678 2568 709
rect 2522 644 2528 678
rect 2562 644 2568 678
rect 2522 606 2568 644
rect 2522 572 2528 606
rect 2562 572 2568 606
rect 2522 534 2568 572
rect 2522 500 2528 534
rect 2562 500 2568 534
rect 2522 462 2568 500
rect 2522 428 2528 462
rect 2562 428 2568 462
rect 2522 390 2568 428
rect 2522 356 2528 390
rect 2562 356 2568 390
rect 2522 318 2568 356
rect 2522 284 2528 318
rect 2562 284 2568 318
rect 2522 246 2568 284
rect 2522 212 2528 246
rect 2562 212 2568 246
rect 2522 174 2568 212
rect 2522 140 2528 174
rect 2562 140 2568 174
rect 2522 109 2568 140
rect 3540 678 3586 709
rect 3540 644 3546 678
rect 3580 644 3586 678
rect 3540 606 3586 644
rect 3540 572 3546 606
rect 3580 572 3586 606
rect 3540 534 3586 572
rect 3540 500 3546 534
rect 3580 500 3586 534
rect 3540 462 3586 500
rect 3540 428 3546 462
rect 3580 428 3586 462
rect 3540 390 3586 428
rect 3540 356 3546 390
rect 3580 356 3586 390
rect 3540 318 3586 356
rect 3540 284 3546 318
rect 3580 284 3586 318
rect 3540 246 3586 284
rect 3540 212 3546 246
rect 3580 212 3586 246
rect 3540 174 3586 212
rect 3540 140 3546 174
rect 3580 140 3586 174
rect 3540 109 3586 140
rect 4558 678 4604 709
rect 4558 644 4564 678
rect 4598 644 4604 678
rect 4558 606 4604 644
rect 4558 572 4564 606
rect 4598 572 4604 606
rect 4558 534 4604 572
rect 4558 500 4564 534
rect 4598 500 4604 534
rect 4558 462 4604 500
rect 4558 428 4564 462
rect 4598 428 4604 462
rect 4558 390 4604 428
rect 4558 356 4564 390
rect 4598 356 4604 390
rect 4558 318 4604 356
rect 4558 284 4564 318
rect 4598 284 4604 318
rect 4558 246 4604 284
rect 4558 212 4564 246
rect 4598 212 4604 246
rect 4558 174 4604 212
rect 4558 140 4564 174
rect 4598 140 4604 174
rect 4558 109 4604 140
rect -4316 71 -3828 77
rect -4316 37 -4269 71
rect -4235 37 -4197 71
rect -4163 37 -4125 71
rect -4091 37 -4053 71
rect -4019 37 -3981 71
rect -3947 37 -3909 71
rect -3875 37 -3828 71
rect -4316 31 -3828 37
rect -3298 71 -2810 77
rect -3298 37 -3251 71
rect -3217 37 -3179 71
rect -3145 37 -3107 71
rect -3073 37 -3035 71
rect -3001 37 -2963 71
rect -2929 37 -2891 71
rect -2857 37 -2810 71
rect -3298 31 -2810 37
rect -2280 71 -1792 77
rect -2280 37 -2233 71
rect -2199 37 -2161 71
rect -2127 37 -2089 71
rect -2055 37 -2017 71
rect -1983 37 -1945 71
rect -1911 37 -1873 71
rect -1839 37 -1792 71
rect -2280 31 -1792 37
rect -1262 71 -774 77
rect -1262 37 -1215 71
rect -1181 37 -1143 71
rect -1109 37 -1071 71
rect -1037 37 -999 71
rect -965 37 -927 71
rect -893 37 -855 71
rect -821 37 -774 71
rect -1262 31 -774 37
rect -244 71 244 77
rect -244 37 -197 71
rect -163 37 -125 71
rect -91 37 -53 71
rect -19 37 19 71
rect 53 37 91 71
rect 125 37 163 71
rect 197 37 244 71
rect -244 31 244 37
rect 774 71 1262 77
rect 774 37 821 71
rect 855 37 893 71
rect 927 37 965 71
rect 999 37 1037 71
rect 1071 37 1109 71
rect 1143 37 1181 71
rect 1215 37 1262 71
rect 774 31 1262 37
rect 1792 71 2280 77
rect 1792 37 1839 71
rect 1873 37 1911 71
rect 1945 37 1983 71
rect 2017 37 2055 71
rect 2089 37 2127 71
rect 2161 37 2199 71
rect 2233 37 2280 71
rect 1792 31 2280 37
rect 2810 71 3298 77
rect 2810 37 2857 71
rect 2891 37 2929 71
rect 2963 37 3001 71
rect 3035 37 3073 71
rect 3107 37 3145 71
rect 3179 37 3217 71
rect 3251 37 3298 71
rect 2810 31 3298 37
rect 3828 71 4316 77
rect 3828 37 3875 71
rect 3909 37 3947 71
rect 3981 37 4019 71
rect 4053 37 4091 71
rect 4125 37 4163 71
rect 4197 37 4235 71
rect 4269 37 4316 71
rect 3828 31 4316 37
rect -4316 -37 -3828 -31
rect -4316 -71 -4269 -37
rect -4235 -71 -4197 -37
rect -4163 -71 -4125 -37
rect -4091 -71 -4053 -37
rect -4019 -71 -3981 -37
rect -3947 -71 -3909 -37
rect -3875 -71 -3828 -37
rect -4316 -77 -3828 -71
rect -3298 -37 -2810 -31
rect -3298 -71 -3251 -37
rect -3217 -71 -3179 -37
rect -3145 -71 -3107 -37
rect -3073 -71 -3035 -37
rect -3001 -71 -2963 -37
rect -2929 -71 -2891 -37
rect -2857 -71 -2810 -37
rect -3298 -77 -2810 -71
rect -2280 -37 -1792 -31
rect -2280 -71 -2233 -37
rect -2199 -71 -2161 -37
rect -2127 -71 -2089 -37
rect -2055 -71 -2017 -37
rect -1983 -71 -1945 -37
rect -1911 -71 -1873 -37
rect -1839 -71 -1792 -37
rect -2280 -77 -1792 -71
rect -1262 -37 -774 -31
rect -1262 -71 -1215 -37
rect -1181 -71 -1143 -37
rect -1109 -71 -1071 -37
rect -1037 -71 -999 -37
rect -965 -71 -927 -37
rect -893 -71 -855 -37
rect -821 -71 -774 -37
rect -1262 -77 -774 -71
rect -244 -37 244 -31
rect -244 -71 -197 -37
rect -163 -71 -125 -37
rect -91 -71 -53 -37
rect -19 -71 19 -37
rect 53 -71 91 -37
rect 125 -71 163 -37
rect 197 -71 244 -37
rect -244 -77 244 -71
rect 774 -37 1262 -31
rect 774 -71 821 -37
rect 855 -71 893 -37
rect 927 -71 965 -37
rect 999 -71 1037 -37
rect 1071 -71 1109 -37
rect 1143 -71 1181 -37
rect 1215 -71 1262 -37
rect 774 -77 1262 -71
rect 1792 -37 2280 -31
rect 1792 -71 1839 -37
rect 1873 -71 1911 -37
rect 1945 -71 1983 -37
rect 2017 -71 2055 -37
rect 2089 -71 2127 -37
rect 2161 -71 2199 -37
rect 2233 -71 2280 -37
rect 1792 -77 2280 -71
rect 2810 -37 3298 -31
rect 2810 -71 2857 -37
rect 2891 -71 2929 -37
rect 2963 -71 3001 -37
rect 3035 -71 3073 -37
rect 3107 -71 3145 -37
rect 3179 -71 3217 -37
rect 3251 -71 3298 -37
rect 2810 -77 3298 -71
rect 3828 -37 4316 -31
rect 3828 -71 3875 -37
rect 3909 -71 3947 -37
rect 3981 -71 4019 -37
rect 4053 -71 4091 -37
rect 4125 -71 4163 -37
rect 4197 -71 4235 -37
rect 4269 -71 4316 -37
rect 3828 -77 4316 -71
rect -4604 -140 -4558 -109
rect -4604 -174 -4598 -140
rect -4564 -174 -4558 -140
rect -4604 -212 -4558 -174
rect -4604 -246 -4598 -212
rect -4564 -246 -4558 -212
rect -4604 -284 -4558 -246
rect -4604 -318 -4598 -284
rect -4564 -318 -4558 -284
rect -4604 -356 -4558 -318
rect -4604 -390 -4598 -356
rect -4564 -390 -4558 -356
rect -4604 -428 -4558 -390
rect -4604 -462 -4598 -428
rect -4564 -462 -4558 -428
rect -4604 -500 -4558 -462
rect -4604 -534 -4598 -500
rect -4564 -534 -4558 -500
rect -4604 -572 -4558 -534
rect -4604 -606 -4598 -572
rect -4564 -606 -4558 -572
rect -4604 -644 -4558 -606
rect -4604 -678 -4598 -644
rect -4564 -678 -4558 -644
rect -4604 -709 -4558 -678
rect -3586 -140 -3540 -109
rect -3586 -174 -3580 -140
rect -3546 -174 -3540 -140
rect -3586 -212 -3540 -174
rect -3586 -246 -3580 -212
rect -3546 -246 -3540 -212
rect -3586 -284 -3540 -246
rect -3586 -318 -3580 -284
rect -3546 -318 -3540 -284
rect -3586 -356 -3540 -318
rect -3586 -390 -3580 -356
rect -3546 -390 -3540 -356
rect -3586 -428 -3540 -390
rect -3586 -462 -3580 -428
rect -3546 -462 -3540 -428
rect -3586 -500 -3540 -462
rect -3586 -534 -3580 -500
rect -3546 -534 -3540 -500
rect -3586 -572 -3540 -534
rect -3586 -606 -3580 -572
rect -3546 -606 -3540 -572
rect -3586 -644 -3540 -606
rect -3586 -678 -3580 -644
rect -3546 -678 -3540 -644
rect -3586 -709 -3540 -678
rect -2568 -140 -2522 -109
rect -2568 -174 -2562 -140
rect -2528 -174 -2522 -140
rect -2568 -212 -2522 -174
rect -2568 -246 -2562 -212
rect -2528 -246 -2522 -212
rect -2568 -284 -2522 -246
rect -2568 -318 -2562 -284
rect -2528 -318 -2522 -284
rect -2568 -356 -2522 -318
rect -2568 -390 -2562 -356
rect -2528 -390 -2522 -356
rect -2568 -428 -2522 -390
rect -2568 -462 -2562 -428
rect -2528 -462 -2522 -428
rect -2568 -500 -2522 -462
rect -2568 -534 -2562 -500
rect -2528 -534 -2522 -500
rect -2568 -572 -2522 -534
rect -2568 -606 -2562 -572
rect -2528 -606 -2522 -572
rect -2568 -644 -2522 -606
rect -2568 -678 -2562 -644
rect -2528 -678 -2522 -644
rect -2568 -709 -2522 -678
rect -1550 -140 -1504 -109
rect -1550 -174 -1544 -140
rect -1510 -174 -1504 -140
rect -1550 -212 -1504 -174
rect -1550 -246 -1544 -212
rect -1510 -246 -1504 -212
rect -1550 -284 -1504 -246
rect -1550 -318 -1544 -284
rect -1510 -318 -1504 -284
rect -1550 -356 -1504 -318
rect -1550 -390 -1544 -356
rect -1510 -390 -1504 -356
rect -1550 -428 -1504 -390
rect -1550 -462 -1544 -428
rect -1510 -462 -1504 -428
rect -1550 -500 -1504 -462
rect -1550 -534 -1544 -500
rect -1510 -534 -1504 -500
rect -1550 -572 -1504 -534
rect -1550 -606 -1544 -572
rect -1510 -606 -1504 -572
rect -1550 -644 -1504 -606
rect -1550 -678 -1544 -644
rect -1510 -678 -1504 -644
rect -1550 -709 -1504 -678
rect -532 -140 -486 -109
rect -532 -174 -526 -140
rect -492 -174 -486 -140
rect -532 -212 -486 -174
rect -532 -246 -526 -212
rect -492 -246 -486 -212
rect -532 -284 -486 -246
rect -532 -318 -526 -284
rect -492 -318 -486 -284
rect -532 -356 -486 -318
rect -532 -390 -526 -356
rect -492 -390 -486 -356
rect -532 -428 -486 -390
rect -532 -462 -526 -428
rect -492 -462 -486 -428
rect -532 -500 -486 -462
rect -532 -534 -526 -500
rect -492 -534 -486 -500
rect -532 -572 -486 -534
rect -532 -606 -526 -572
rect -492 -606 -486 -572
rect -532 -644 -486 -606
rect -532 -678 -526 -644
rect -492 -678 -486 -644
rect -532 -709 -486 -678
rect 486 -140 532 -109
rect 486 -174 492 -140
rect 526 -174 532 -140
rect 486 -212 532 -174
rect 486 -246 492 -212
rect 526 -246 532 -212
rect 486 -284 532 -246
rect 486 -318 492 -284
rect 526 -318 532 -284
rect 486 -356 532 -318
rect 486 -390 492 -356
rect 526 -390 532 -356
rect 486 -428 532 -390
rect 486 -462 492 -428
rect 526 -462 532 -428
rect 486 -500 532 -462
rect 486 -534 492 -500
rect 526 -534 532 -500
rect 486 -572 532 -534
rect 486 -606 492 -572
rect 526 -606 532 -572
rect 486 -644 532 -606
rect 486 -678 492 -644
rect 526 -678 532 -644
rect 486 -709 532 -678
rect 1504 -140 1550 -109
rect 1504 -174 1510 -140
rect 1544 -174 1550 -140
rect 1504 -212 1550 -174
rect 1504 -246 1510 -212
rect 1544 -246 1550 -212
rect 1504 -284 1550 -246
rect 1504 -318 1510 -284
rect 1544 -318 1550 -284
rect 1504 -356 1550 -318
rect 1504 -390 1510 -356
rect 1544 -390 1550 -356
rect 1504 -428 1550 -390
rect 1504 -462 1510 -428
rect 1544 -462 1550 -428
rect 1504 -500 1550 -462
rect 1504 -534 1510 -500
rect 1544 -534 1550 -500
rect 1504 -572 1550 -534
rect 1504 -606 1510 -572
rect 1544 -606 1550 -572
rect 1504 -644 1550 -606
rect 1504 -678 1510 -644
rect 1544 -678 1550 -644
rect 1504 -709 1550 -678
rect 2522 -140 2568 -109
rect 2522 -174 2528 -140
rect 2562 -174 2568 -140
rect 2522 -212 2568 -174
rect 2522 -246 2528 -212
rect 2562 -246 2568 -212
rect 2522 -284 2568 -246
rect 2522 -318 2528 -284
rect 2562 -318 2568 -284
rect 2522 -356 2568 -318
rect 2522 -390 2528 -356
rect 2562 -390 2568 -356
rect 2522 -428 2568 -390
rect 2522 -462 2528 -428
rect 2562 -462 2568 -428
rect 2522 -500 2568 -462
rect 2522 -534 2528 -500
rect 2562 -534 2568 -500
rect 2522 -572 2568 -534
rect 2522 -606 2528 -572
rect 2562 -606 2568 -572
rect 2522 -644 2568 -606
rect 2522 -678 2528 -644
rect 2562 -678 2568 -644
rect 2522 -709 2568 -678
rect 3540 -140 3586 -109
rect 3540 -174 3546 -140
rect 3580 -174 3586 -140
rect 3540 -212 3586 -174
rect 3540 -246 3546 -212
rect 3580 -246 3586 -212
rect 3540 -284 3586 -246
rect 3540 -318 3546 -284
rect 3580 -318 3586 -284
rect 3540 -356 3586 -318
rect 3540 -390 3546 -356
rect 3580 -390 3586 -356
rect 3540 -428 3586 -390
rect 3540 -462 3546 -428
rect 3580 -462 3586 -428
rect 3540 -500 3586 -462
rect 3540 -534 3546 -500
rect 3580 -534 3586 -500
rect 3540 -572 3586 -534
rect 3540 -606 3546 -572
rect 3580 -606 3586 -572
rect 3540 -644 3586 -606
rect 3540 -678 3546 -644
rect 3580 -678 3586 -644
rect 3540 -709 3586 -678
rect 4558 -140 4604 -109
rect 4558 -174 4564 -140
rect 4598 -174 4604 -140
rect 4558 -212 4604 -174
rect 4558 -246 4564 -212
rect 4598 -246 4604 -212
rect 4558 -284 4604 -246
rect 4558 -318 4564 -284
rect 4598 -318 4604 -284
rect 4558 -356 4604 -318
rect 4558 -390 4564 -356
rect 4598 -390 4604 -356
rect 4558 -428 4604 -390
rect 4558 -462 4564 -428
rect 4598 -462 4604 -428
rect 4558 -500 4604 -462
rect 4558 -534 4564 -500
rect 4598 -534 4604 -500
rect 4558 -572 4604 -534
rect 4558 -606 4564 -572
rect 4598 -606 4604 -572
rect 4558 -644 4604 -606
rect 4558 -678 4564 -644
rect 4598 -678 4604 -644
rect 4558 -709 4604 -678
rect -4316 -747 -3828 -741
rect -4316 -781 -4269 -747
rect -4235 -781 -4197 -747
rect -4163 -781 -4125 -747
rect -4091 -781 -4053 -747
rect -4019 -781 -3981 -747
rect -3947 -781 -3909 -747
rect -3875 -781 -3828 -747
rect -4316 -787 -3828 -781
rect -3298 -747 -2810 -741
rect -3298 -781 -3251 -747
rect -3217 -781 -3179 -747
rect -3145 -781 -3107 -747
rect -3073 -781 -3035 -747
rect -3001 -781 -2963 -747
rect -2929 -781 -2891 -747
rect -2857 -781 -2810 -747
rect -3298 -787 -2810 -781
rect -2280 -747 -1792 -741
rect -2280 -781 -2233 -747
rect -2199 -781 -2161 -747
rect -2127 -781 -2089 -747
rect -2055 -781 -2017 -747
rect -1983 -781 -1945 -747
rect -1911 -781 -1873 -747
rect -1839 -781 -1792 -747
rect -2280 -787 -1792 -781
rect -1262 -747 -774 -741
rect -1262 -781 -1215 -747
rect -1181 -781 -1143 -747
rect -1109 -781 -1071 -747
rect -1037 -781 -999 -747
rect -965 -781 -927 -747
rect -893 -781 -855 -747
rect -821 -781 -774 -747
rect -1262 -787 -774 -781
rect -244 -747 244 -741
rect -244 -781 -197 -747
rect -163 -781 -125 -747
rect -91 -781 -53 -747
rect -19 -781 19 -747
rect 53 -781 91 -747
rect 125 -781 163 -747
rect 197 -781 244 -747
rect -244 -787 244 -781
rect 774 -747 1262 -741
rect 774 -781 821 -747
rect 855 -781 893 -747
rect 927 -781 965 -747
rect 999 -781 1037 -747
rect 1071 -781 1109 -747
rect 1143 -781 1181 -747
rect 1215 -781 1262 -747
rect 774 -787 1262 -781
rect 1792 -747 2280 -741
rect 1792 -781 1839 -747
rect 1873 -781 1911 -747
rect 1945 -781 1983 -747
rect 2017 -781 2055 -747
rect 2089 -781 2127 -747
rect 2161 -781 2199 -747
rect 2233 -781 2280 -747
rect 1792 -787 2280 -781
rect 2810 -747 3298 -741
rect 2810 -781 2857 -747
rect 2891 -781 2929 -747
rect 2963 -781 3001 -747
rect 3035 -781 3073 -747
rect 3107 -781 3145 -747
rect 3179 -781 3217 -747
rect 3251 -781 3298 -747
rect 2810 -787 3298 -781
rect 3828 -747 4316 -741
rect 3828 -781 3875 -747
rect 3909 -781 3947 -747
rect 3981 -781 4019 -747
rect 4053 -781 4091 -747
rect 4125 -781 4163 -747
rect 4197 -781 4235 -747
rect 4269 -781 4316 -747
rect 3828 -787 4316 -781
rect -4316 -855 -3828 -849
rect -4316 -889 -4269 -855
rect -4235 -889 -4197 -855
rect -4163 -889 -4125 -855
rect -4091 -889 -4053 -855
rect -4019 -889 -3981 -855
rect -3947 -889 -3909 -855
rect -3875 -889 -3828 -855
rect -4316 -895 -3828 -889
rect -3298 -855 -2810 -849
rect -3298 -889 -3251 -855
rect -3217 -889 -3179 -855
rect -3145 -889 -3107 -855
rect -3073 -889 -3035 -855
rect -3001 -889 -2963 -855
rect -2929 -889 -2891 -855
rect -2857 -889 -2810 -855
rect -3298 -895 -2810 -889
rect -2280 -855 -1792 -849
rect -2280 -889 -2233 -855
rect -2199 -889 -2161 -855
rect -2127 -889 -2089 -855
rect -2055 -889 -2017 -855
rect -1983 -889 -1945 -855
rect -1911 -889 -1873 -855
rect -1839 -889 -1792 -855
rect -2280 -895 -1792 -889
rect -1262 -855 -774 -849
rect -1262 -889 -1215 -855
rect -1181 -889 -1143 -855
rect -1109 -889 -1071 -855
rect -1037 -889 -999 -855
rect -965 -889 -927 -855
rect -893 -889 -855 -855
rect -821 -889 -774 -855
rect -1262 -895 -774 -889
rect -244 -855 244 -849
rect -244 -889 -197 -855
rect -163 -889 -125 -855
rect -91 -889 -53 -855
rect -19 -889 19 -855
rect 53 -889 91 -855
rect 125 -889 163 -855
rect 197 -889 244 -855
rect -244 -895 244 -889
rect 774 -855 1262 -849
rect 774 -889 821 -855
rect 855 -889 893 -855
rect 927 -889 965 -855
rect 999 -889 1037 -855
rect 1071 -889 1109 -855
rect 1143 -889 1181 -855
rect 1215 -889 1262 -855
rect 774 -895 1262 -889
rect 1792 -855 2280 -849
rect 1792 -889 1839 -855
rect 1873 -889 1911 -855
rect 1945 -889 1983 -855
rect 2017 -889 2055 -855
rect 2089 -889 2127 -855
rect 2161 -889 2199 -855
rect 2233 -889 2280 -855
rect 1792 -895 2280 -889
rect 2810 -855 3298 -849
rect 2810 -889 2857 -855
rect 2891 -889 2929 -855
rect 2963 -889 3001 -855
rect 3035 -889 3073 -855
rect 3107 -889 3145 -855
rect 3179 -889 3217 -855
rect 3251 -889 3298 -855
rect 2810 -895 3298 -889
rect 3828 -855 4316 -849
rect 3828 -889 3875 -855
rect 3909 -889 3947 -855
rect 3981 -889 4019 -855
rect 4053 -889 4091 -855
rect 4125 -889 4163 -855
rect 4197 -889 4235 -855
rect 4269 -889 4316 -855
rect 3828 -895 4316 -889
rect -4604 -958 -4558 -927
rect -4604 -992 -4598 -958
rect -4564 -992 -4558 -958
rect -4604 -1030 -4558 -992
rect -4604 -1064 -4598 -1030
rect -4564 -1064 -4558 -1030
rect -4604 -1102 -4558 -1064
rect -4604 -1136 -4598 -1102
rect -4564 -1136 -4558 -1102
rect -4604 -1174 -4558 -1136
rect -4604 -1208 -4598 -1174
rect -4564 -1208 -4558 -1174
rect -4604 -1246 -4558 -1208
rect -4604 -1280 -4598 -1246
rect -4564 -1280 -4558 -1246
rect -4604 -1318 -4558 -1280
rect -4604 -1352 -4598 -1318
rect -4564 -1352 -4558 -1318
rect -4604 -1390 -4558 -1352
rect -4604 -1424 -4598 -1390
rect -4564 -1424 -4558 -1390
rect -4604 -1462 -4558 -1424
rect -4604 -1496 -4598 -1462
rect -4564 -1496 -4558 -1462
rect -4604 -1527 -4558 -1496
rect -3586 -958 -3540 -927
rect -3586 -992 -3580 -958
rect -3546 -992 -3540 -958
rect -3586 -1030 -3540 -992
rect -3586 -1064 -3580 -1030
rect -3546 -1064 -3540 -1030
rect -3586 -1102 -3540 -1064
rect -3586 -1136 -3580 -1102
rect -3546 -1136 -3540 -1102
rect -3586 -1174 -3540 -1136
rect -3586 -1208 -3580 -1174
rect -3546 -1208 -3540 -1174
rect -3586 -1246 -3540 -1208
rect -3586 -1280 -3580 -1246
rect -3546 -1280 -3540 -1246
rect -3586 -1318 -3540 -1280
rect -3586 -1352 -3580 -1318
rect -3546 -1352 -3540 -1318
rect -3586 -1390 -3540 -1352
rect -3586 -1424 -3580 -1390
rect -3546 -1424 -3540 -1390
rect -3586 -1462 -3540 -1424
rect -3586 -1496 -3580 -1462
rect -3546 -1496 -3540 -1462
rect -3586 -1527 -3540 -1496
rect -2568 -958 -2522 -927
rect -2568 -992 -2562 -958
rect -2528 -992 -2522 -958
rect -2568 -1030 -2522 -992
rect -2568 -1064 -2562 -1030
rect -2528 -1064 -2522 -1030
rect -2568 -1102 -2522 -1064
rect -2568 -1136 -2562 -1102
rect -2528 -1136 -2522 -1102
rect -2568 -1174 -2522 -1136
rect -2568 -1208 -2562 -1174
rect -2528 -1208 -2522 -1174
rect -2568 -1246 -2522 -1208
rect -2568 -1280 -2562 -1246
rect -2528 -1280 -2522 -1246
rect -2568 -1318 -2522 -1280
rect -2568 -1352 -2562 -1318
rect -2528 -1352 -2522 -1318
rect -2568 -1390 -2522 -1352
rect -2568 -1424 -2562 -1390
rect -2528 -1424 -2522 -1390
rect -2568 -1462 -2522 -1424
rect -2568 -1496 -2562 -1462
rect -2528 -1496 -2522 -1462
rect -2568 -1527 -2522 -1496
rect -1550 -958 -1504 -927
rect -1550 -992 -1544 -958
rect -1510 -992 -1504 -958
rect -1550 -1030 -1504 -992
rect -1550 -1064 -1544 -1030
rect -1510 -1064 -1504 -1030
rect -1550 -1102 -1504 -1064
rect -1550 -1136 -1544 -1102
rect -1510 -1136 -1504 -1102
rect -1550 -1174 -1504 -1136
rect -1550 -1208 -1544 -1174
rect -1510 -1208 -1504 -1174
rect -1550 -1246 -1504 -1208
rect -1550 -1280 -1544 -1246
rect -1510 -1280 -1504 -1246
rect -1550 -1318 -1504 -1280
rect -1550 -1352 -1544 -1318
rect -1510 -1352 -1504 -1318
rect -1550 -1390 -1504 -1352
rect -1550 -1424 -1544 -1390
rect -1510 -1424 -1504 -1390
rect -1550 -1462 -1504 -1424
rect -1550 -1496 -1544 -1462
rect -1510 -1496 -1504 -1462
rect -1550 -1527 -1504 -1496
rect -532 -958 -486 -927
rect -532 -992 -526 -958
rect -492 -992 -486 -958
rect -532 -1030 -486 -992
rect -532 -1064 -526 -1030
rect -492 -1064 -486 -1030
rect -532 -1102 -486 -1064
rect -532 -1136 -526 -1102
rect -492 -1136 -486 -1102
rect -532 -1174 -486 -1136
rect -532 -1208 -526 -1174
rect -492 -1208 -486 -1174
rect -532 -1246 -486 -1208
rect -532 -1280 -526 -1246
rect -492 -1280 -486 -1246
rect -532 -1318 -486 -1280
rect -532 -1352 -526 -1318
rect -492 -1352 -486 -1318
rect -532 -1390 -486 -1352
rect -532 -1424 -526 -1390
rect -492 -1424 -486 -1390
rect -532 -1462 -486 -1424
rect -532 -1496 -526 -1462
rect -492 -1496 -486 -1462
rect -532 -1527 -486 -1496
rect 486 -958 532 -927
rect 486 -992 492 -958
rect 526 -992 532 -958
rect 486 -1030 532 -992
rect 486 -1064 492 -1030
rect 526 -1064 532 -1030
rect 486 -1102 532 -1064
rect 486 -1136 492 -1102
rect 526 -1136 532 -1102
rect 486 -1174 532 -1136
rect 486 -1208 492 -1174
rect 526 -1208 532 -1174
rect 486 -1246 532 -1208
rect 486 -1280 492 -1246
rect 526 -1280 532 -1246
rect 486 -1318 532 -1280
rect 486 -1352 492 -1318
rect 526 -1352 532 -1318
rect 486 -1390 532 -1352
rect 486 -1424 492 -1390
rect 526 -1424 532 -1390
rect 486 -1462 532 -1424
rect 486 -1496 492 -1462
rect 526 -1496 532 -1462
rect 486 -1527 532 -1496
rect 1504 -958 1550 -927
rect 1504 -992 1510 -958
rect 1544 -992 1550 -958
rect 1504 -1030 1550 -992
rect 1504 -1064 1510 -1030
rect 1544 -1064 1550 -1030
rect 1504 -1102 1550 -1064
rect 1504 -1136 1510 -1102
rect 1544 -1136 1550 -1102
rect 1504 -1174 1550 -1136
rect 1504 -1208 1510 -1174
rect 1544 -1208 1550 -1174
rect 1504 -1246 1550 -1208
rect 1504 -1280 1510 -1246
rect 1544 -1280 1550 -1246
rect 1504 -1318 1550 -1280
rect 1504 -1352 1510 -1318
rect 1544 -1352 1550 -1318
rect 1504 -1390 1550 -1352
rect 1504 -1424 1510 -1390
rect 1544 -1424 1550 -1390
rect 1504 -1462 1550 -1424
rect 1504 -1496 1510 -1462
rect 1544 -1496 1550 -1462
rect 1504 -1527 1550 -1496
rect 2522 -958 2568 -927
rect 2522 -992 2528 -958
rect 2562 -992 2568 -958
rect 2522 -1030 2568 -992
rect 2522 -1064 2528 -1030
rect 2562 -1064 2568 -1030
rect 2522 -1102 2568 -1064
rect 2522 -1136 2528 -1102
rect 2562 -1136 2568 -1102
rect 2522 -1174 2568 -1136
rect 2522 -1208 2528 -1174
rect 2562 -1208 2568 -1174
rect 2522 -1246 2568 -1208
rect 2522 -1280 2528 -1246
rect 2562 -1280 2568 -1246
rect 2522 -1318 2568 -1280
rect 2522 -1352 2528 -1318
rect 2562 -1352 2568 -1318
rect 2522 -1390 2568 -1352
rect 2522 -1424 2528 -1390
rect 2562 -1424 2568 -1390
rect 2522 -1462 2568 -1424
rect 2522 -1496 2528 -1462
rect 2562 -1496 2568 -1462
rect 2522 -1527 2568 -1496
rect 3540 -958 3586 -927
rect 3540 -992 3546 -958
rect 3580 -992 3586 -958
rect 3540 -1030 3586 -992
rect 3540 -1064 3546 -1030
rect 3580 -1064 3586 -1030
rect 3540 -1102 3586 -1064
rect 3540 -1136 3546 -1102
rect 3580 -1136 3586 -1102
rect 3540 -1174 3586 -1136
rect 3540 -1208 3546 -1174
rect 3580 -1208 3586 -1174
rect 3540 -1246 3586 -1208
rect 3540 -1280 3546 -1246
rect 3580 -1280 3586 -1246
rect 3540 -1318 3586 -1280
rect 3540 -1352 3546 -1318
rect 3580 -1352 3586 -1318
rect 3540 -1390 3586 -1352
rect 3540 -1424 3546 -1390
rect 3580 -1424 3586 -1390
rect 3540 -1462 3586 -1424
rect 3540 -1496 3546 -1462
rect 3580 -1496 3586 -1462
rect 3540 -1527 3586 -1496
rect 4558 -958 4604 -927
rect 4558 -992 4564 -958
rect 4598 -992 4604 -958
rect 4558 -1030 4604 -992
rect 4558 -1064 4564 -1030
rect 4598 -1064 4604 -1030
rect 4558 -1102 4604 -1064
rect 4558 -1136 4564 -1102
rect 4598 -1136 4604 -1102
rect 4558 -1174 4604 -1136
rect 4558 -1208 4564 -1174
rect 4598 -1208 4604 -1174
rect 4558 -1246 4604 -1208
rect 4558 -1280 4564 -1246
rect 4598 -1280 4604 -1246
rect 4558 -1318 4604 -1280
rect 4558 -1352 4564 -1318
rect 4598 -1352 4604 -1318
rect 4558 -1390 4604 -1352
rect 4558 -1424 4564 -1390
rect 4598 -1424 4604 -1390
rect 4558 -1462 4604 -1424
rect 4558 -1496 4564 -1462
rect 4598 -1496 4604 -1462
rect 4558 -1527 4604 -1496
rect -4316 -1565 -3828 -1559
rect -4316 -1599 -4269 -1565
rect -4235 -1599 -4197 -1565
rect -4163 -1599 -4125 -1565
rect -4091 -1599 -4053 -1565
rect -4019 -1599 -3981 -1565
rect -3947 -1599 -3909 -1565
rect -3875 -1599 -3828 -1565
rect -4316 -1605 -3828 -1599
rect -3298 -1565 -2810 -1559
rect -3298 -1599 -3251 -1565
rect -3217 -1599 -3179 -1565
rect -3145 -1599 -3107 -1565
rect -3073 -1599 -3035 -1565
rect -3001 -1599 -2963 -1565
rect -2929 -1599 -2891 -1565
rect -2857 -1599 -2810 -1565
rect -3298 -1605 -2810 -1599
rect -2280 -1565 -1792 -1559
rect -2280 -1599 -2233 -1565
rect -2199 -1599 -2161 -1565
rect -2127 -1599 -2089 -1565
rect -2055 -1599 -2017 -1565
rect -1983 -1599 -1945 -1565
rect -1911 -1599 -1873 -1565
rect -1839 -1599 -1792 -1565
rect -2280 -1605 -1792 -1599
rect -1262 -1565 -774 -1559
rect -1262 -1599 -1215 -1565
rect -1181 -1599 -1143 -1565
rect -1109 -1599 -1071 -1565
rect -1037 -1599 -999 -1565
rect -965 -1599 -927 -1565
rect -893 -1599 -855 -1565
rect -821 -1599 -774 -1565
rect -1262 -1605 -774 -1599
rect -244 -1565 244 -1559
rect -244 -1599 -197 -1565
rect -163 -1599 -125 -1565
rect -91 -1599 -53 -1565
rect -19 -1599 19 -1565
rect 53 -1599 91 -1565
rect 125 -1599 163 -1565
rect 197 -1599 244 -1565
rect -244 -1605 244 -1599
rect 774 -1565 1262 -1559
rect 774 -1599 821 -1565
rect 855 -1599 893 -1565
rect 927 -1599 965 -1565
rect 999 -1599 1037 -1565
rect 1071 -1599 1109 -1565
rect 1143 -1599 1181 -1565
rect 1215 -1599 1262 -1565
rect 774 -1605 1262 -1599
rect 1792 -1565 2280 -1559
rect 1792 -1599 1839 -1565
rect 1873 -1599 1911 -1565
rect 1945 -1599 1983 -1565
rect 2017 -1599 2055 -1565
rect 2089 -1599 2127 -1565
rect 2161 -1599 2199 -1565
rect 2233 -1599 2280 -1565
rect 1792 -1605 2280 -1599
rect 2810 -1565 3298 -1559
rect 2810 -1599 2857 -1565
rect 2891 -1599 2929 -1565
rect 2963 -1599 3001 -1565
rect 3035 -1599 3073 -1565
rect 3107 -1599 3145 -1565
rect 3179 -1599 3217 -1565
rect 3251 -1599 3298 -1565
rect 2810 -1605 3298 -1599
rect 3828 -1565 4316 -1559
rect 3828 -1599 3875 -1565
rect 3909 -1599 3947 -1565
rect 3981 -1599 4019 -1565
rect 4053 -1599 4091 -1565
rect 4125 -1599 4163 -1565
rect 4197 -1599 4235 -1565
rect 4269 -1599 4316 -1565
rect 3828 -1605 4316 -1599
<< end >>
