magic
tech sky130A
magscale 1 2
timestamp 1622700284
<< nwell >>
rect 30 3318 23246 5174
rect 30 -5978 23246 -4122
<< pwell >>
rect 30 -322 11446 3154
rect 11830 -322 23246 3154
rect 30 -3958 11446 -482
rect 11830 -3958 23246 -482
<< nmos >>
rect 1170 2158 1370 2558
rect 1428 2158 1628 2558
rect 1686 2158 1886 2558
rect 1944 2158 2144 2558
rect 2202 2158 2402 2558
rect 2460 2158 2660 2558
rect 2718 2158 2918 2558
rect 2976 2158 3176 2558
rect 3234 2158 3434 2558
rect 3492 2158 3692 2558
rect 7762 2158 7962 2558
rect 8020 2158 8220 2558
rect 8278 2158 8478 2558
rect 8536 2158 8736 2558
rect 8794 2158 8994 2558
rect 9052 2158 9252 2558
rect 9310 2158 9510 2558
rect 9568 2158 9768 2558
rect 9826 2158 10026 2558
rect 10084 2158 10284 2558
rect 622 1250 1422 1450
rect 1480 1250 2280 1450
rect 2338 1250 3138 1450
rect 3196 1250 3996 1450
rect 4054 1250 4854 1450
rect 4912 1250 5712 1450
rect 5770 1250 6570 1450
rect 6628 1250 7428 1450
rect 7486 1250 8286 1450
rect 8344 1250 9144 1450
rect 9202 1250 10002 1450
rect 10060 1250 10860 1450
rect 622 710 1422 910
rect 1480 710 2280 910
rect 2338 710 3138 910
rect 3196 710 3996 910
rect 4054 710 4854 910
rect 4912 710 5712 910
rect 5770 710 6570 910
rect 6628 710 7428 910
rect 7486 710 8286 910
rect 8344 710 9144 910
rect 9202 710 10002 910
rect 10060 710 10860 910
rect 12970 2158 13170 2558
rect 13228 2158 13428 2558
rect 13486 2158 13686 2558
rect 13744 2158 13944 2558
rect 14002 2158 14202 2558
rect 14260 2158 14460 2558
rect 14518 2158 14718 2558
rect 14776 2158 14976 2558
rect 15034 2158 15234 2558
rect 15292 2158 15492 2558
rect 19562 2158 19762 2558
rect 19820 2158 20020 2558
rect 20078 2158 20278 2558
rect 20336 2158 20536 2558
rect 20594 2158 20794 2558
rect 20852 2158 21052 2558
rect 21110 2158 21310 2558
rect 21368 2158 21568 2558
rect 21626 2158 21826 2558
rect 21884 2158 22084 2558
rect 12422 1250 13222 1450
rect 13280 1250 14080 1450
rect 14138 1250 14938 1450
rect 14996 1250 15796 1450
rect 15854 1250 16654 1450
rect 16712 1250 17512 1450
rect 17570 1250 18370 1450
rect 18428 1250 19228 1450
rect 19286 1250 20086 1450
rect 20144 1250 20944 1450
rect 21002 1250 21802 1450
rect 21860 1250 22660 1450
rect 12422 710 13222 910
rect 13280 710 14080 910
rect 14138 710 14938 910
rect 14996 710 15796 910
rect 15854 710 16654 910
rect 16712 710 17512 910
rect 17570 710 18370 910
rect 18428 710 19228 910
rect 19286 710 20086 910
rect 20144 710 20944 910
rect 21002 710 21802 910
rect 21860 710 22660 910
rect 622 -1714 1422 -1514
rect 1480 -1714 2280 -1514
rect 2338 -1714 3138 -1514
rect 3196 -1714 3996 -1514
rect 4054 -1714 4854 -1514
rect 4912 -1714 5712 -1514
rect 5770 -1714 6570 -1514
rect 6628 -1714 7428 -1514
rect 7486 -1714 8286 -1514
rect 8344 -1714 9144 -1514
rect 9202 -1714 10002 -1514
rect 10060 -1714 10860 -1514
rect 622 -2254 1422 -2054
rect 1480 -2254 2280 -2054
rect 2338 -2254 3138 -2054
rect 3196 -2254 3996 -2054
rect 4054 -2254 4854 -2054
rect 4912 -2254 5712 -2054
rect 5770 -2254 6570 -2054
rect 6628 -2254 7428 -2054
rect 7486 -2254 8286 -2054
rect 8344 -2254 9144 -2054
rect 9202 -2254 10002 -2054
rect 10060 -2254 10860 -2054
rect 1170 -3362 1370 -2962
rect 1428 -3362 1628 -2962
rect 1686 -3362 1886 -2962
rect 1944 -3362 2144 -2962
rect 2202 -3362 2402 -2962
rect 2460 -3362 2660 -2962
rect 2718 -3362 2918 -2962
rect 2976 -3362 3176 -2962
rect 3234 -3362 3434 -2962
rect 3492 -3362 3692 -2962
rect 7762 -3362 7962 -2962
rect 8020 -3362 8220 -2962
rect 8278 -3362 8478 -2962
rect 8536 -3362 8736 -2962
rect 8794 -3362 8994 -2962
rect 9052 -3362 9252 -2962
rect 9310 -3362 9510 -2962
rect 9568 -3362 9768 -2962
rect 9826 -3362 10026 -2962
rect 10084 -3362 10284 -2962
rect 12422 -1714 13222 -1514
rect 13280 -1714 14080 -1514
rect 14138 -1714 14938 -1514
rect 14996 -1714 15796 -1514
rect 15854 -1714 16654 -1514
rect 16712 -1714 17512 -1514
rect 17570 -1714 18370 -1514
rect 18428 -1714 19228 -1514
rect 19286 -1714 20086 -1514
rect 20144 -1714 20944 -1514
rect 21002 -1714 21802 -1514
rect 21860 -1714 22660 -1514
rect 12422 -2254 13222 -2054
rect 13280 -2254 14080 -2054
rect 14138 -2254 14938 -2054
rect 14996 -2254 15796 -2054
rect 15854 -2254 16654 -2054
rect 16712 -2254 17512 -2054
rect 17570 -2254 18370 -2054
rect 18428 -2254 19228 -2054
rect 19286 -2254 20086 -2054
rect 20144 -2254 20944 -2054
rect 21002 -2254 21802 -2054
rect 21860 -2254 22660 -2054
rect 12970 -3362 13170 -2962
rect 13228 -3362 13428 -2962
rect 13486 -3362 13686 -2962
rect 13744 -3362 13944 -2962
rect 14002 -3362 14202 -2962
rect 14260 -3362 14460 -2962
rect 14518 -3362 14718 -2962
rect 14776 -3362 14976 -2962
rect 15034 -3362 15234 -2962
rect 15292 -3362 15492 -2962
rect 19562 -3362 19762 -2962
rect 19820 -3362 20020 -2962
rect 20078 -3362 20278 -2962
rect 20336 -3362 20536 -2962
rect 20594 -3362 20794 -2962
rect 20852 -3362 21052 -2962
rect 21110 -3362 21310 -2962
rect 21368 -3362 21568 -2962
rect 21626 -3362 21826 -2962
rect 21884 -3362 22084 -2962
<< pmos >>
rect 3954 3826 4154 4026
rect 4212 3826 4412 4026
rect 4470 3826 4670 4026
rect 4728 3826 4928 4026
rect 4986 3826 5186 4026
rect 5244 3826 5444 4026
rect 5502 3826 5702 4026
rect 5760 3826 5960 4026
rect 6018 3826 6218 4026
rect 6276 3826 6476 4026
rect 6534 3826 6734 4026
rect 6792 3826 6992 4026
rect 7050 3826 7250 4026
rect 7308 3826 7508 4026
rect 15754 3826 15954 4026
rect 16012 3826 16212 4026
rect 16270 3826 16470 4026
rect 16528 3826 16728 4026
rect 16786 3826 16986 4026
rect 17044 3826 17244 4026
rect 17302 3826 17502 4026
rect 17560 3826 17760 4026
rect 17818 3826 18018 4026
rect 18076 3826 18276 4026
rect 18334 3826 18534 4026
rect 18592 3826 18792 4026
rect 18850 3826 19050 4026
rect 19108 3826 19308 4026
rect 3954 -4830 4154 -4630
rect 4212 -4830 4412 -4630
rect 4470 -4830 4670 -4630
rect 4728 -4830 4928 -4630
rect 4986 -4830 5186 -4630
rect 5244 -4830 5444 -4630
rect 5502 -4830 5702 -4630
rect 5760 -4830 5960 -4630
rect 6018 -4830 6218 -4630
rect 6276 -4830 6476 -4630
rect 6534 -4830 6734 -4630
rect 6792 -4830 6992 -4630
rect 7050 -4830 7250 -4630
rect 7308 -4830 7508 -4630
rect 15754 -4830 15954 -4630
rect 16012 -4830 16212 -4630
rect 16270 -4830 16470 -4630
rect 16528 -4830 16728 -4630
rect 16786 -4830 16986 -4630
rect 17044 -4830 17244 -4630
rect 17302 -4830 17502 -4630
rect 17560 -4830 17760 -4630
rect 17818 -4830 18018 -4630
rect 18076 -4830 18276 -4630
rect 18334 -4830 18534 -4630
rect 18592 -4830 18792 -4630
rect 18850 -4830 19050 -4630
rect 19108 -4830 19308 -4630
<< nmoslvt >>
rect 4466 2158 4666 2558
rect 4724 2158 4924 2558
rect 4982 2158 5182 2558
rect 5240 2158 5440 2558
rect 5498 2158 5698 2558
rect 5756 2158 5956 2558
rect 6014 2158 6214 2558
rect 6272 2158 6472 2558
rect 6530 2158 6730 2558
rect 6788 2158 6988 2558
rect 16266 2158 16466 2558
rect 16524 2158 16724 2558
rect 16782 2158 16982 2558
rect 17040 2158 17240 2558
rect 17298 2158 17498 2558
rect 17556 2158 17756 2558
rect 17814 2158 18014 2558
rect 18072 2158 18272 2558
rect 18330 2158 18530 2558
rect 18588 2158 18788 2558
rect 4466 -3362 4666 -2962
rect 4724 -3362 4924 -2962
rect 4982 -3362 5182 -2962
rect 5240 -3362 5440 -2962
rect 5498 -3362 5698 -2962
rect 5756 -3362 5956 -2962
rect 6014 -3362 6214 -2962
rect 6272 -3362 6472 -2962
rect 6530 -3362 6730 -2962
rect 6788 -3362 6988 -2962
rect 16266 -3362 16466 -2962
rect 16524 -3362 16724 -2962
rect 16782 -3362 16982 -2962
rect 17040 -3362 17240 -2962
rect 17298 -3362 17498 -2962
rect 17556 -3362 17756 -2962
rect 17814 -3362 18014 -2962
rect 18072 -3362 18272 -2962
rect 18330 -3362 18530 -2962
rect 18588 -3362 18788 -2962
<< ndiff >>
rect 1112 2546 1170 2558
rect 1112 2170 1124 2546
rect 1158 2170 1170 2546
rect 1112 2158 1170 2170
rect 1370 2546 1428 2558
rect 1370 2170 1382 2546
rect 1416 2170 1428 2546
rect 1370 2158 1428 2170
rect 1628 2546 1686 2558
rect 1628 2170 1640 2546
rect 1674 2170 1686 2546
rect 1628 2158 1686 2170
rect 1886 2546 1944 2558
rect 1886 2170 1898 2546
rect 1932 2170 1944 2546
rect 1886 2158 1944 2170
rect 2144 2546 2202 2558
rect 2144 2170 2156 2546
rect 2190 2170 2202 2546
rect 2144 2158 2202 2170
rect 2402 2546 2460 2558
rect 2402 2170 2414 2546
rect 2448 2170 2460 2546
rect 2402 2158 2460 2170
rect 2660 2546 2718 2558
rect 2660 2170 2672 2546
rect 2706 2170 2718 2546
rect 2660 2158 2718 2170
rect 2918 2546 2976 2558
rect 2918 2170 2930 2546
rect 2964 2170 2976 2546
rect 2918 2158 2976 2170
rect 3176 2546 3234 2558
rect 3176 2170 3188 2546
rect 3222 2170 3234 2546
rect 3176 2158 3234 2170
rect 3434 2546 3492 2558
rect 3434 2170 3446 2546
rect 3480 2170 3492 2546
rect 3434 2158 3492 2170
rect 3692 2546 3750 2558
rect 3692 2170 3704 2546
rect 3738 2170 3750 2546
rect 3692 2158 3750 2170
rect 4408 2546 4466 2558
rect 4408 2170 4420 2546
rect 4454 2170 4466 2546
rect 4408 2158 4466 2170
rect 4666 2546 4724 2558
rect 4666 2170 4678 2546
rect 4712 2170 4724 2546
rect 4666 2158 4724 2170
rect 4924 2546 4982 2558
rect 4924 2170 4936 2546
rect 4970 2170 4982 2546
rect 4924 2158 4982 2170
rect 5182 2546 5240 2558
rect 5182 2170 5194 2546
rect 5228 2170 5240 2546
rect 5182 2158 5240 2170
rect 5440 2546 5498 2558
rect 5440 2170 5452 2546
rect 5486 2170 5498 2546
rect 5440 2158 5498 2170
rect 5698 2546 5756 2558
rect 5698 2170 5710 2546
rect 5744 2170 5756 2546
rect 5698 2158 5756 2170
rect 5956 2546 6014 2558
rect 5956 2170 5968 2546
rect 6002 2170 6014 2546
rect 5956 2158 6014 2170
rect 6214 2546 6272 2558
rect 6214 2170 6226 2546
rect 6260 2170 6272 2546
rect 6214 2158 6272 2170
rect 6472 2546 6530 2558
rect 6472 2170 6484 2546
rect 6518 2170 6530 2546
rect 6472 2158 6530 2170
rect 6730 2546 6788 2558
rect 6730 2170 6742 2546
rect 6776 2170 6788 2546
rect 6730 2158 6788 2170
rect 6988 2546 7046 2558
rect 6988 2170 7000 2546
rect 7034 2170 7046 2546
rect 6988 2158 7046 2170
rect 7704 2546 7762 2558
rect 7704 2170 7716 2546
rect 7750 2170 7762 2546
rect 7704 2158 7762 2170
rect 7962 2546 8020 2558
rect 7962 2170 7974 2546
rect 8008 2170 8020 2546
rect 7962 2158 8020 2170
rect 8220 2546 8278 2558
rect 8220 2170 8232 2546
rect 8266 2170 8278 2546
rect 8220 2158 8278 2170
rect 8478 2546 8536 2558
rect 8478 2170 8490 2546
rect 8524 2170 8536 2546
rect 8478 2158 8536 2170
rect 8736 2546 8794 2558
rect 8736 2170 8748 2546
rect 8782 2170 8794 2546
rect 8736 2158 8794 2170
rect 8994 2546 9052 2558
rect 8994 2170 9006 2546
rect 9040 2170 9052 2546
rect 8994 2158 9052 2170
rect 9252 2546 9310 2558
rect 9252 2170 9264 2546
rect 9298 2170 9310 2546
rect 9252 2158 9310 2170
rect 9510 2546 9568 2558
rect 9510 2170 9522 2546
rect 9556 2170 9568 2546
rect 9510 2158 9568 2170
rect 9768 2546 9826 2558
rect 9768 2170 9780 2546
rect 9814 2170 9826 2546
rect 9768 2158 9826 2170
rect 10026 2546 10084 2558
rect 10026 2170 10038 2546
rect 10072 2170 10084 2546
rect 10026 2158 10084 2170
rect 10284 2546 10342 2558
rect 10284 2170 10296 2546
rect 10330 2170 10342 2546
rect 10284 2158 10342 2170
rect 564 1438 622 1450
rect 564 1262 576 1438
rect 610 1262 622 1438
rect 564 1250 622 1262
rect 1422 1438 1480 1450
rect 1422 1262 1434 1438
rect 1468 1262 1480 1438
rect 1422 1250 1480 1262
rect 2280 1438 2338 1450
rect 2280 1262 2292 1438
rect 2326 1262 2338 1438
rect 2280 1250 2338 1262
rect 3138 1438 3196 1450
rect 3138 1262 3150 1438
rect 3184 1262 3196 1438
rect 3138 1250 3196 1262
rect 3996 1438 4054 1450
rect 3996 1262 4008 1438
rect 4042 1262 4054 1438
rect 3996 1250 4054 1262
rect 4854 1438 4912 1450
rect 4854 1262 4866 1438
rect 4900 1262 4912 1438
rect 4854 1250 4912 1262
rect 5712 1438 5770 1450
rect 5712 1262 5724 1438
rect 5758 1262 5770 1438
rect 5712 1250 5770 1262
rect 6570 1438 6628 1450
rect 6570 1262 6582 1438
rect 6616 1262 6628 1438
rect 6570 1250 6628 1262
rect 7428 1438 7486 1450
rect 7428 1262 7440 1438
rect 7474 1262 7486 1438
rect 7428 1250 7486 1262
rect 8286 1438 8344 1450
rect 8286 1262 8298 1438
rect 8332 1262 8344 1438
rect 8286 1250 8344 1262
rect 9144 1438 9202 1450
rect 9144 1262 9156 1438
rect 9190 1262 9202 1438
rect 9144 1250 9202 1262
rect 10002 1438 10060 1450
rect 10002 1262 10014 1438
rect 10048 1262 10060 1438
rect 10002 1250 10060 1262
rect 10860 1438 10918 1450
rect 10860 1262 10872 1438
rect 10906 1262 10918 1438
rect 10860 1250 10918 1262
rect 564 898 622 910
rect 564 722 576 898
rect 610 722 622 898
rect 564 710 622 722
rect 1422 898 1480 910
rect 1422 722 1434 898
rect 1468 722 1480 898
rect 1422 710 1480 722
rect 2280 898 2338 910
rect 2280 722 2292 898
rect 2326 722 2338 898
rect 2280 710 2338 722
rect 3138 898 3196 910
rect 3138 722 3150 898
rect 3184 722 3196 898
rect 3138 710 3196 722
rect 3996 898 4054 910
rect 3996 722 4008 898
rect 4042 722 4054 898
rect 3996 710 4054 722
rect 4854 898 4912 910
rect 4854 722 4866 898
rect 4900 722 4912 898
rect 4854 710 4912 722
rect 5712 898 5770 910
rect 5712 722 5724 898
rect 5758 722 5770 898
rect 5712 710 5770 722
rect 6570 898 6628 910
rect 6570 722 6582 898
rect 6616 722 6628 898
rect 6570 710 6628 722
rect 7428 898 7486 910
rect 7428 722 7440 898
rect 7474 722 7486 898
rect 7428 710 7486 722
rect 8286 898 8344 910
rect 8286 722 8298 898
rect 8332 722 8344 898
rect 8286 710 8344 722
rect 9144 898 9202 910
rect 9144 722 9156 898
rect 9190 722 9202 898
rect 9144 710 9202 722
rect 10002 898 10060 910
rect 10002 722 10014 898
rect 10048 722 10060 898
rect 10002 710 10060 722
rect 10860 898 10918 910
rect 10860 722 10872 898
rect 10906 722 10918 898
rect 10860 710 10918 722
rect 12912 2546 12970 2558
rect 12912 2170 12924 2546
rect 12958 2170 12970 2546
rect 12912 2158 12970 2170
rect 13170 2546 13228 2558
rect 13170 2170 13182 2546
rect 13216 2170 13228 2546
rect 13170 2158 13228 2170
rect 13428 2546 13486 2558
rect 13428 2170 13440 2546
rect 13474 2170 13486 2546
rect 13428 2158 13486 2170
rect 13686 2546 13744 2558
rect 13686 2170 13698 2546
rect 13732 2170 13744 2546
rect 13686 2158 13744 2170
rect 13944 2546 14002 2558
rect 13944 2170 13956 2546
rect 13990 2170 14002 2546
rect 13944 2158 14002 2170
rect 14202 2546 14260 2558
rect 14202 2170 14214 2546
rect 14248 2170 14260 2546
rect 14202 2158 14260 2170
rect 14460 2546 14518 2558
rect 14460 2170 14472 2546
rect 14506 2170 14518 2546
rect 14460 2158 14518 2170
rect 14718 2546 14776 2558
rect 14718 2170 14730 2546
rect 14764 2170 14776 2546
rect 14718 2158 14776 2170
rect 14976 2546 15034 2558
rect 14976 2170 14988 2546
rect 15022 2170 15034 2546
rect 14976 2158 15034 2170
rect 15234 2546 15292 2558
rect 15234 2170 15246 2546
rect 15280 2170 15292 2546
rect 15234 2158 15292 2170
rect 15492 2546 15550 2558
rect 15492 2170 15504 2546
rect 15538 2170 15550 2546
rect 15492 2158 15550 2170
rect 16208 2546 16266 2558
rect 16208 2170 16220 2546
rect 16254 2170 16266 2546
rect 16208 2158 16266 2170
rect 16466 2546 16524 2558
rect 16466 2170 16478 2546
rect 16512 2170 16524 2546
rect 16466 2158 16524 2170
rect 16724 2546 16782 2558
rect 16724 2170 16736 2546
rect 16770 2170 16782 2546
rect 16724 2158 16782 2170
rect 16982 2546 17040 2558
rect 16982 2170 16994 2546
rect 17028 2170 17040 2546
rect 16982 2158 17040 2170
rect 17240 2546 17298 2558
rect 17240 2170 17252 2546
rect 17286 2170 17298 2546
rect 17240 2158 17298 2170
rect 17498 2546 17556 2558
rect 17498 2170 17510 2546
rect 17544 2170 17556 2546
rect 17498 2158 17556 2170
rect 17756 2546 17814 2558
rect 17756 2170 17768 2546
rect 17802 2170 17814 2546
rect 17756 2158 17814 2170
rect 18014 2546 18072 2558
rect 18014 2170 18026 2546
rect 18060 2170 18072 2546
rect 18014 2158 18072 2170
rect 18272 2546 18330 2558
rect 18272 2170 18284 2546
rect 18318 2170 18330 2546
rect 18272 2158 18330 2170
rect 18530 2546 18588 2558
rect 18530 2170 18542 2546
rect 18576 2170 18588 2546
rect 18530 2158 18588 2170
rect 18788 2546 18846 2558
rect 18788 2170 18800 2546
rect 18834 2170 18846 2546
rect 18788 2158 18846 2170
rect 19504 2546 19562 2558
rect 19504 2170 19516 2546
rect 19550 2170 19562 2546
rect 19504 2158 19562 2170
rect 19762 2546 19820 2558
rect 19762 2170 19774 2546
rect 19808 2170 19820 2546
rect 19762 2158 19820 2170
rect 20020 2546 20078 2558
rect 20020 2170 20032 2546
rect 20066 2170 20078 2546
rect 20020 2158 20078 2170
rect 20278 2546 20336 2558
rect 20278 2170 20290 2546
rect 20324 2170 20336 2546
rect 20278 2158 20336 2170
rect 20536 2546 20594 2558
rect 20536 2170 20548 2546
rect 20582 2170 20594 2546
rect 20536 2158 20594 2170
rect 20794 2546 20852 2558
rect 20794 2170 20806 2546
rect 20840 2170 20852 2546
rect 20794 2158 20852 2170
rect 21052 2546 21110 2558
rect 21052 2170 21064 2546
rect 21098 2170 21110 2546
rect 21052 2158 21110 2170
rect 21310 2546 21368 2558
rect 21310 2170 21322 2546
rect 21356 2170 21368 2546
rect 21310 2158 21368 2170
rect 21568 2546 21626 2558
rect 21568 2170 21580 2546
rect 21614 2170 21626 2546
rect 21568 2158 21626 2170
rect 21826 2546 21884 2558
rect 21826 2170 21838 2546
rect 21872 2170 21884 2546
rect 21826 2158 21884 2170
rect 22084 2546 22142 2558
rect 22084 2170 22096 2546
rect 22130 2170 22142 2546
rect 22084 2158 22142 2170
rect 12364 1438 12422 1450
rect 12364 1262 12376 1438
rect 12410 1262 12422 1438
rect 12364 1250 12422 1262
rect 13222 1438 13280 1450
rect 13222 1262 13234 1438
rect 13268 1262 13280 1438
rect 13222 1250 13280 1262
rect 14080 1438 14138 1450
rect 14080 1262 14092 1438
rect 14126 1262 14138 1438
rect 14080 1250 14138 1262
rect 14938 1438 14996 1450
rect 14938 1262 14950 1438
rect 14984 1262 14996 1438
rect 14938 1250 14996 1262
rect 15796 1438 15854 1450
rect 15796 1262 15808 1438
rect 15842 1262 15854 1438
rect 15796 1250 15854 1262
rect 16654 1438 16712 1450
rect 16654 1262 16666 1438
rect 16700 1262 16712 1438
rect 16654 1250 16712 1262
rect 17512 1438 17570 1450
rect 17512 1262 17524 1438
rect 17558 1262 17570 1438
rect 17512 1250 17570 1262
rect 18370 1438 18428 1450
rect 18370 1262 18382 1438
rect 18416 1262 18428 1438
rect 18370 1250 18428 1262
rect 19228 1438 19286 1450
rect 19228 1262 19240 1438
rect 19274 1262 19286 1438
rect 19228 1250 19286 1262
rect 20086 1438 20144 1450
rect 20086 1262 20098 1438
rect 20132 1262 20144 1438
rect 20086 1250 20144 1262
rect 20944 1438 21002 1450
rect 20944 1262 20956 1438
rect 20990 1262 21002 1438
rect 20944 1250 21002 1262
rect 21802 1438 21860 1450
rect 21802 1262 21814 1438
rect 21848 1262 21860 1438
rect 21802 1250 21860 1262
rect 22660 1438 22718 1450
rect 22660 1262 22672 1438
rect 22706 1262 22718 1438
rect 22660 1250 22718 1262
rect 12364 898 12422 910
rect 12364 722 12376 898
rect 12410 722 12422 898
rect 12364 710 12422 722
rect 13222 898 13280 910
rect 13222 722 13234 898
rect 13268 722 13280 898
rect 13222 710 13280 722
rect 14080 898 14138 910
rect 14080 722 14092 898
rect 14126 722 14138 898
rect 14080 710 14138 722
rect 14938 898 14996 910
rect 14938 722 14950 898
rect 14984 722 14996 898
rect 14938 710 14996 722
rect 15796 898 15854 910
rect 15796 722 15808 898
rect 15842 722 15854 898
rect 15796 710 15854 722
rect 16654 898 16712 910
rect 16654 722 16666 898
rect 16700 722 16712 898
rect 16654 710 16712 722
rect 17512 898 17570 910
rect 17512 722 17524 898
rect 17558 722 17570 898
rect 17512 710 17570 722
rect 18370 898 18428 910
rect 18370 722 18382 898
rect 18416 722 18428 898
rect 18370 710 18428 722
rect 19228 898 19286 910
rect 19228 722 19240 898
rect 19274 722 19286 898
rect 19228 710 19286 722
rect 20086 898 20144 910
rect 20086 722 20098 898
rect 20132 722 20144 898
rect 20086 710 20144 722
rect 20944 898 21002 910
rect 20944 722 20956 898
rect 20990 722 21002 898
rect 20944 710 21002 722
rect 21802 898 21860 910
rect 21802 722 21814 898
rect 21848 722 21860 898
rect 21802 710 21860 722
rect 22660 898 22718 910
rect 22660 722 22672 898
rect 22706 722 22718 898
rect 22660 710 22718 722
rect 564 -1526 622 -1514
rect 564 -1702 576 -1526
rect 610 -1702 622 -1526
rect 564 -1714 622 -1702
rect 1422 -1526 1480 -1514
rect 1422 -1702 1434 -1526
rect 1468 -1702 1480 -1526
rect 1422 -1714 1480 -1702
rect 2280 -1526 2338 -1514
rect 2280 -1702 2292 -1526
rect 2326 -1702 2338 -1526
rect 2280 -1714 2338 -1702
rect 3138 -1526 3196 -1514
rect 3138 -1702 3150 -1526
rect 3184 -1702 3196 -1526
rect 3138 -1714 3196 -1702
rect 3996 -1526 4054 -1514
rect 3996 -1702 4008 -1526
rect 4042 -1702 4054 -1526
rect 3996 -1714 4054 -1702
rect 4854 -1526 4912 -1514
rect 4854 -1702 4866 -1526
rect 4900 -1702 4912 -1526
rect 4854 -1714 4912 -1702
rect 5712 -1526 5770 -1514
rect 5712 -1702 5724 -1526
rect 5758 -1702 5770 -1526
rect 5712 -1714 5770 -1702
rect 6570 -1526 6628 -1514
rect 6570 -1702 6582 -1526
rect 6616 -1702 6628 -1526
rect 6570 -1714 6628 -1702
rect 7428 -1526 7486 -1514
rect 7428 -1702 7440 -1526
rect 7474 -1702 7486 -1526
rect 7428 -1714 7486 -1702
rect 8286 -1526 8344 -1514
rect 8286 -1702 8298 -1526
rect 8332 -1702 8344 -1526
rect 8286 -1714 8344 -1702
rect 9144 -1526 9202 -1514
rect 9144 -1702 9156 -1526
rect 9190 -1702 9202 -1526
rect 9144 -1714 9202 -1702
rect 10002 -1526 10060 -1514
rect 10002 -1702 10014 -1526
rect 10048 -1702 10060 -1526
rect 10002 -1714 10060 -1702
rect 10860 -1526 10918 -1514
rect 10860 -1702 10872 -1526
rect 10906 -1702 10918 -1526
rect 10860 -1714 10918 -1702
rect 564 -2066 622 -2054
rect 564 -2242 576 -2066
rect 610 -2242 622 -2066
rect 564 -2254 622 -2242
rect 1422 -2066 1480 -2054
rect 1422 -2242 1434 -2066
rect 1468 -2242 1480 -2066
rect 1422 -2254 1480 -2242
rect 2280 -2066 2338 -2054
rect 2280 -2242 2292 -2066
rect 2326 -2242 2338 -2066
rect 2280 -2254 2338 -2242
rect 3138 -2066 3196 -2054
rect 3138 -2242 3150 -2066
rect 3184 -2242 3196 -2066
rect 3138 -2254 3196 -2242
rect 3996 -2066 4054 -2054
rect 3996 -2242 4008 -2066
rect 4042 -2242 4054 -2066
rect 3996 -2254 4054 -2242
rect 4854 -2066 4912 -2054
rect 4854 -2242 4866 -2066
rect 4900 -2242 4912 -2066
rect 4854 -2254 4912 -2242
rect 5712 -2066 5770 -2054
rect 5712 -2242 5724 -2066
rect 5758 -2242 5770 -2066
rect 5712 -2254 5770 -2242
rect 6570 -2066 6628 -2054
rect 6570 -2242 6582 -2066
rect 6616 -2242 6628 -2066
rect 6570 -2254 6628 -2242
rect 7428 -2066 7486 -2054
rect 7428 -2242 7440 -2066
rect 7474 -2242 7486 -2066
rect 7428 -2254 7486 -2242
rect 8286 -2066 8344 -2054
rect 8286 -2242 8298 -2066
rect 8332 -2242 8344 -2066
rect 8286 -2254 8344 -2242
rect 9144 -2066 9202 -2054
rect 9144 -2242 9156 -2066
rect 9190 -2242 9202 -2066
rect 9144 -2254 9202 -2242
rect 10002 -2066 10060 -2054
rect 10002 -2242 10014 -2066
rect 10048 -2242 10060 -2066
rect 10002 -2254 10060 -2242
rect 10860 -2066 10918 -2054
rect 10860 -2242 10872 -2066
rect 10906 -2242 10918 -2066
rect 10860 -2254 10918 -2242
rect 1112 -2974 1170 -2962
rect 1112 -3350 1124 -2974
rect 1158 -3350 1170 -2974
rect 1112 -3362 1170 -3350
rect 1370 -2974 1428 -2962
rect 1370 -3350 1382 -2974
rect 1416 -3350 1428 -2974
rect 1370 -3362 1428 -3350
rect 1628 -2974 1686 -2962
rect 1628 -3350 1640 -2974
rect 1674 -3350 1686 -2974
rect 1628 -3362 1686 -3350
rect 1886 -2974 1944 -2962
rect 1886 -3350 1898 -2974
rect 1932 -3350 1944 -2974
rect 1886 -3362 1944 -3350
rect 2144 -2974 2202 -2962
rect 2144 -3350 2156 -2974
rect 2190 -3350 2202 -2974
rect 2144 -3362 2202 -3350
rect 2402 -2974 2460 -2962
rect 2402 -3350 2414 -2974
rect 2448 -3350 2460 -2974
rect 2402 -3362 2460 -3350
rect 2660 -2974 2718 -2962
rect 2660 -3350 2672 -2974
rect 2706 -3350 2718 -2974
rect 2660 -3362 2718 -3350
rect 2918 -2974 2976 -2962
rect 2918 -3350 2930 -2974
rect 2964 -3350 2976 -2974
rect 2918 -3362 2976 -3350
rect 3176 -2974 3234 -2962
rect 3176 -3350 3188 -2974
rect 3222 -3350 3234 -2974
rect 3176 -3362 3234 -3350
rect 3434 -2974 3492 -2962
rect 3434 -3350 3446 -2974
rect 3480 -3350 3492 -2974
rect 3434 -3362 3492 -3350
rect 3692 -2974 3750 -2962
rect 3692 -3350 3704 -2974
rect 3738 -3350 3750 -2974
rect 3692 -3362 3750 -3350
rect 4408 -2974 4466 -2962
rect 4408 -3350 4420 -2974
rect 4454 -3350 4466 -2974
rect 4408 -3362 4466 -3350
rect 4666 -2974 4724 -2962
rect 4666 -3350 4678 -2974
rect 4712 -3350 4724 -2974
rect 4666 -3362 4724 -3350
rect 4924 -2974 4982 -2962
rect 4924 -3350 4936 -2974
rect 4970 -3350 4982 -2974
rect 4924 -3362 4982 -3350
rect 5182 -2974 5240 -2962
rect 5182 -3350 5194 -2974
rect 5228 -3350 5240 -2974
rect 5182 -3362 5240 -3350
rect 5440 -2974 5498 -2962
rect 5440 -3350 5452 -2974
rect 5486 -3350 5498 -2974
rect 5440 -3362 5498 -3350
rect 5698 -2974 5756 -2962
rect 5698 -3350 5710 -2974
rect 5744 -3350 5756 -2974
rect 5698 -3362 5756 -3350
rect 5956 -2974 6014 -2962
rect 5956 -3350 5968 -2974
rect 6002 -3350 6014 -2974
rect 5956 -3362 6014 -3350
rect 6214 -2974 6272 -2962
rect 6214 -3350 6226 -2974
rect 6260 -3350 6272 -2974
rect 6214 -3362 6272 -3350
rect 6472 -2974 6530 -2962
rect 6472 -3350 6484 -2974
rect 6518 -3350 6530 -2974
rect 6472 -3362 6530 -3350
rect 6730 -2974 6788 -2962
rect 6730 -3350 6742 -2974
rect 6776 -3350 6788 -2974
rect 6730 -3362 6788 -3350
rect 6988 -2974 7046 -2962
rect 6988 -3350 7000 -2974
rect 7034 -3350 7046 -2974
rect 6988 -3362 7046 -3350
rect 7704 -2974 7762 -2962
rect 7704 -3350 7716 -2974
rect 7750 -3350 7762 -2974
rect 7704 -3362 7762 -3350
rect 7962 -2974 8020 -2962
rect 7962 -3350 7974 -2974
rect 8008 -3350 8020 -2974
rect 7962 -3362 8020 -3350
rect 8220 -2974 8278 -2962
rect 8220 -3350 8232 -2974
rect 8266 -3350 8278 -2974
rect 8220 -3362 8278 -3350
rect 8478 -2974 8536 -2962
rect 8478 -3350 8490 -2974
rect 8524 -3350 8536 -2974
rect 8478 -3362 8536 -3350
rect 8736 -2974 8794 -2962
rect 8736 -3350 8748 -2974
rect 8782 -3350 8794 -2974
rect 8736 -3362 8794 -3350
rect 8994 -2974 9052 -2962
rect 8994 -3350 9006 -2974
rect 9040 -3350 9052 -2974
rect 8994 -3362 9052 -3350
rect 9252 -2974 9310 -2962
rect 9252 -3350 9264 -2974
rect 9298 -3350 9310 -2974
rect 9252 -3362 9310 -3350
rect 9510 -2974 9568 -2962
rect 9510 -3350 9522 -2974
rect 9556 -3350 9568 -2974
rect 9510 -3362 9568 -3350
rect 9768 -2974 9826 -2962
rect 9768 -3350 9780 -2974
rect 9814 -3350 9826 -2974
rect 9768 -3362 9826 -3350
rect 10026 -2974 10084 -2962
rect 10026 -3350 10038 -2974
rect 10072 -3350 10084 -2974
rect 10026 -3362 10084 -3350
rect 10284 -2974 10342 -2962
rect 10284 -3350 10296 -2974
rect 10330 -3350 10342 -2974
rect 10284 -3362 10342 -3350
rect 12364 -1526 12422 -1514
rect 12364 -1702 12376 -1526
rect 12410 -1702 12422 -1526
rect 12364 -1714 12422 -1702
rect 13222 -1526 13280 -1514
rect 13222 -1702 13234 -1526
rect 13268 -1702 13280 -1526
rect 13222 -1714 13280 -1702
rect 14080 -1526 14138 -1514
rect 14080 -1702 14092 -1526
rect 14126 -1702 14138 -1526
rect 14080 -1714 14138 -1702
rect 14938 -1526 14996 -1514
rect 14938 -1702 14950 -1526
rect 14984 -1702 14996 -1526
rect 14938 -1714 14996 -1702
rect 15796 -1526 15854 -1514
rect 15796 -1702 15808 -1526
rect 15842 -1702 15854 -1526
rect 15796 -1714 15854 -1702
rect 16654 -1526 16712 -1514
rect 16654 -1702 16666 -1526
rect 16700 -1702 16712 -1526
rect 16654 -1714 16712 -1702
rect 17512 -1526 17570 -1514
rect 17512 -1702 17524 -1526
rect 17558 -1702 17570 -1526
rect 17512 -1714 17570 -1702
rect 18370 -1526 18428 -1514
rect 18370 -1702 18382 -1526
rect 18416 -1702 18428 -1526
rect 18370 -1714 18428 -1702
rect 19228 -1526 19286 -1514
rect 19228 -1702 19240 -1526
rect 19274 -1702 19286 -1526
rect 19228 -1714 19286 -1702
rect 20086 -1526 20144 -1514
rect 20086 -1702 20098 -1526
rect 20132 -1702 20144 -1526
rect 20086 -1714 20144 -1702
rect 20944 -1526 21002 -1514
rect 20944 -1702 20956 -1526
rect 20990 -1702 21002 -1526
rect 20944 -1714 21002 -1702
rect 21802 -1526 21860 -1514
rect 21802 -1702 21814 -1526
rect 21848 -1702 21860 -1526
rect 21802 -1714 21860 -1702
rect 22660 -1526 22718 -1514
rect 22660 -1702 22672 -1526
rect 22706 -1702 22718 -1526
rect 22660 -1714 22718 -1702
rect 12364 -2066 12422 -2054
rect 12364 -2242 12376 -2066
rect 12410 -2242 12422 -2066
rect 12364 -2254 12422 -2242
rect 13222 -2066 13280 -2054
rect 13222 -2242 13234 -2066
rect 13268 -2242 13280 -2066
rect 13222 -2254 13280 -2242
rect 14080 -2066 14138 -2054
rect 14080 -2242 14092 -2066
rect 14126 -2242 14138 -2066
rect 14080 -2254 14138 -2242
rect 14938 -2066 14996 -2054
rect 14938 -2242 14950 -2066
rect 14984 -2242 14996 -2066
rect 14938 -2254 14996 -2242
rect 15796 -2066 15854 -2054
rect 15796 -2242 15808 -2066
rect 15842 -2242 15854 -2066
rect 15796 -2254 15854 -2242
rect 16654 -2066 16712 -2054
rect 16654 -2242 16666 -2066
rect 16700 -2242 16712 -2066
rect 16654 -2254 16712 -2242
rect 17512 -2066 17570 -2054
rect 17512 -2242 17524 -2066
rect 17558 -2242 17570 -2066
rect 17512 -2254 17570 -2242
rect 18370 -2066 18428 -2054
rect 18370 -2242 18382 -2066
rect 18416 -2242 18428 -2066
rect 18370 -2254 18428 -2242
rect 19228 -2066 19286 -2054
rect 19228 -2242 19240 -2066
rect 19274 -2242 19286 -2066
rect 19228 -2254 19286 -2242
rect 20086 -2066 20144 -2054
rect 20086 -2242 20098 -2066
rect 20132 -2242 20144 -2066
rect 20086 -2254 20144 -2242
rect 20944 -2066 21002 -2054
rect 20944 -2242 20956 -2066
rect 20990 -2242 21002 -2066
rect 20944 -2254 21002 -2242
rect 21802 -2066 21860 -2054
rect 21802 -2242 21814 -2066
rect 21848 -2242 21860 -2066
rect 21802 -2254 21860 -2242
rect 22660 -2066 22718 -2054
rect 22660 -2242 22672 -2066
rect 22706 -2242 22718 -2066
rect 22660 -2254 22718 -2242
rect 12912 -2974 12970 -2962
rect 12912 -3350 12924 -2974
rect 12958 -3350 12970 -2974
rect 12912 -3362 12970 -3350
rect 13170 -2974 13228 -2962
rect 13170 -3350 13182 -2974
rect 13216 -3350 13228 -2974
rect 13170 -3362 13228 -3350
rect 13428 -2974 13486 -2962
rect 13428 -3350 13440 -2974
rect 13474 -3350 13486 -2974
rect 13428 -3362 13486 -3350
rect 13686 -2974 13744 -2962
rect 13686 -3350 13698 -2974
rect 13732 -3350 13744 -2974
rect 13686 -3362 13744 -3350
rect 13944 -2974 14002 -2962
rect 13944 -3350 13956 -2974
rect 13990 -3350 14002 -2974
rect 13944 -3362 14002 -3350
rect 14202 -2974 14260 -2962
rect 14202 -3350 14214 -2974
rect 14248 -3350 14260 -2974
rect 14202 -3362 14260 -3350
rect 14460 -2974 14518 -2962
rect 14460 -3350 14472 -2974
rect 14506 -3350 14518 -2974
rect 14460 -3362 14518 -3350
rect 14718 -2974 14776 -2962
rect 14718 -3350 14730 -2974
rect 14764 -3350 14776 -2974
rect 14718 -3362 14776 -3350
rect 14976 -2974 15034 -2962
rect 14976 -3350 14988 -2974
rect 15022 -3350 15034 -2974
rect 14976 -3362 15034 -3350
rect 15234 -2974 15292 -2962
rect 15234 -3350 15246 -2974
rect 15280 -3350 15292 -2974
rect 15234 -3362 15292 -3350
rect 15492 -2974 15550 -2962
rect 15492 -3350 15504 -2974
rect 15538 -3350 15550 -2974
rect 15492 -3362 15550 -3350
rect 16208 -2974 16266 -2962
rect 16208 -3350 16220 -2974
rect 16254 -3350 16266 -2974
rect 16208 -3362 16266 -3350
rect 16466 -2974 16524 -2962
rect 16466 -3350 16478 -2974
rect 16512 -3350 16524 -2974
rect 16466 -3362 16524 -3350
rect 16724 -2974 16782 -2962
rect 16724 -3350 16736 -2974
rect 16770 -3350 16782 -2974
rect 16724 -3362 16782 -3350
rect 16982 -2974 17040 -2962
rect 16982 -3350 16994 -2974
rect 17028 -3350 17040 -2974
rect 16982 -3362 17040 -3350
rect 17240 -2974 17298 -2962
rect 17240 -3350 17252 -2974
rect 17286 -3350 17298 -2974
rect 17240 -3362 17298 -3350
rect 17498 -2974 17556 -2962
rect 17498 -3350 17510 -2974
rect 17544 -3350 17556 -2974
rect 17498 -3362 17556 -3350
rect 17756 -2974 17814 -2962
rect 17756 -3350 17768 -2974
rect 17802 -3350 17814 -2974
rect 17756 -3362 17814 -3350
rect 18014 -2974 18072 -2962
rect 18014 -3350 18026 -2974
rect 18060 -3350 18072 -2974
rect 18014 -3362 18072 -3350
rect 18272 -2974 18330 -2962
rect 18272 -3350 18284 -2974
rect 18318 -3350 18330 -2974
rect 18272 -3362 18330 -3350
rect 18530 -2974 18588 -2962
rect 18530 -3350 18542 -2974
rect 18576 -3350 18588 -2974
rect 18530 -3362 18588 -3350
rect 18788 -2974 18846 -2962
rect 18788 -3350 18800 -2974
rect 18834 -3350 18846 -2974
rect 18788 -3362 18846 -3350
rect 19504 -2974 19562 -2962
rect 19504 -3350 19516 -2974
rect 19550 -3350 19562 -2974
rect 19504 -3362 19562 -3350
rect 19762 -2974 19820 -2962
rect 19762 -3350 19774 -2974
rect 19808 -3350 19820 -2974
rect 19762 -3362 19820 -3350
rect 20020 -2974 20078 -2962
rect 20020 -3350 20032 -2974
rect 20066 -3350 20078 -2974
rect 20020 -3362 20078 -3350
rect 20278 -2974 20336 -2962
rect 20278 -3350 20290 -2974
rect 20324 -3350 20336 -2974
rect 20278 -3362 20336 -3350
rect 20536 -2974 20594 -2962
rect 20536 -3350 20548 -2974
rect 20582 -3350 20594 -2974
rect 20536 -3362 20594 -3350
rect 20794 -2974 20852 -2962
rect 20794 -3350 20806 -2974
rect 20840 -3350 20852 -2974
rect 20794 -3362 20852 -3350
rect 21052 -2974 21110 -2962
rect 21052 -3350 21064 -2974
rect 21098 -3350 21110 -2974
rect 21052 -3362 21110 -3350
rect 21310 -2974 21368 -2962
rect 21310 -3350 21322 -2974
rect 21356 -3350 21368 -2974
rect 21310 -3362 21368 -3350
rect 21568 -2974 21626 -2962
rect 21568 -3350 21580 -2974
rect 21614 -3350 21626 -2974
rect 21568 -3362 21626 -3350
rect 21826 -2974 21884 -2962
rect 21826 -3350 21838 -2974
rect 21872 -3350 21884 -2974
rect 21826 -3362 21884 -3350
rect 22084 -2974 22142 -2962
rect 22084 -3350 22096 -2974
rect 22130 -3350 22142 -2974
rect 22084 -3362 22142 -3350
<< pdiff >>
rect 3896 4014 3954 4026
rect 3896 3838 3908 4014
rect 3942 3838 3954 4014
rect 3896 3826 3954 3838
rect 4154 4014 4212 4026
rect 4154 3838 4166 4014
rect 4200 3838 4212 4014
rect 4154 3826 4212 3838
rect 4412 4014 4470 4026
rect 4412 3838 4424 4014
rect 4458 3838 4470 4014
rect 4412 3826 4470 3838
rect 4670 4014 4728 4026
rect 4670 3838 4682 4014
rect 4716 3838 4728 4014
rect 4670 3826 4728 3838
rect 4928 4014 4986 4026
rect 4928 3838 4940 4014
rect 4974 3838 4986 4014
rect 4928 3826 4986 3838
rect 5186 4014 5244 4026
rect 5186 3838 5198 4014
rect 5232 3838 5244 4014
rect 5186 3826 5244 3838
rect 5444 4014 5502 4026
rect 5444 3838 5456 4014
rect 5490 3838 5502 4014
rect 5444 3826 5502 3838
rect 5702 4014 5760 4026
rect 5702 3838 5714 4014
rect 5748 3838 5760 4014
rect 5702 3826 5760 3838
rect 5960 4014 6018 4026
rect 5960 3838 5972 4014
rect 6006 3838 6018 4014
rect 5960 3826 6018 3838
rect 6218 4014 6276 4026
rect 6218 3838 6230 4014
rect 6264 3838 6276 4014
rect 6218 3826 6276 3838
rect 6476 4014 6534 4026
rect 6476 3838 6488 4014
rect 6522 3838 6534 4014
rect 6476 3826 6534 3838
rect 6734 4014 6792 4026
rect 6734 3838 6746 4014
rect 6780 3838 6792 4014
rect 6734 3826 6792 3838
rect 6992 4014 7050 4026
rect 6992 3838 7004 4014
rect 7038 3838 7050 4014
rect 6992 3826 7050 3838
rect 7250 4014 7308 4026
rect 7250 3838 7262 4014
rect 7296 3838 7308 4014
rect 7250 3826 7308 3838
rect 7508 4014 7566 4026
rect 7508 3838 7520 4014
rect 7554 3838 7566 4014
rect 7508 3826 7566 3838
rect 15696 4014 15754 4026
rect 15696 3838 15708 4014
rect 15742 3838 15754 4014
rect 15696 3826 15754 3838
rect 15954 4014 16012 4026
rect 15954 3838 15966 4014
rect 16000 3838 16012 4014
rect 15954 3826 16012 3838
rect 16212 4014 16270 4026
rect 16212 3838 16224 4014
rect 16258 3838 16270 4014
rect 16212 3826 16270 3838
rect 16470 4014 16528 4026
rect 16470 3838 16482 4014
rect 16516 3838 16528 4014
rect 16470 3826 16528 3838
rect 16728 4014 16786 4026
rect 16728 3838 16740 4014
rect 16774 3838 16786 4014
rect 16728 3826 16786 3838
rect 16986 4014 17044 4026
rect 16986 3838 16998 4014
rect 17032 3838 17044 4014
rect 16986 3826 17044 3838
rect 17244 4014 17302 4026
rect 17244 3838 17256 4014
rect 17290 3838 17302 4014
rect 17244 3826 17302 3838
rect 17502 4014 17560 4026
rect 17502 3838 17514 4014
rect 17548 3838 17560 4014
rect 17502 3826 17560 3838
rect 17760 4014 17818 4026
rect 17760 3838 17772 4014
rect 17806 3838 17818 4014
rect 17760 3826 17818 3838
rect 18018 4014 18076 4026
rect 18018 3838 18030 4014
rect 18064 3838 18076 4014
rect 18018 3826 18076 3838
rect 18276 4014 18334 4026
rect 18276 3838 18288 4014
rect 18322 3838 18334 4014
rect 18276 3826 18334 3838
rect 18534 4014 18592 4026
rect 18534 3838 18546 4014
rect 18580 3838 18592 4014
rect 18534 3826 18592 3838
rect 18792 4014 18850 4026
rect 18792 3838 18804 4014
rect 18838 3838 18850 4014
rect 18792 3826 18850 3838
rect 19050 4014 19108 4026
rect 19050 3838 19062 4014
rect 19096 3838 19108 4014
rect 19050 3826 19108 3838
rect 19308 4014 19366 4026
rect 19308 3838 19320 4014
rect 19354 3838 19366 4014
rect 19308 3826 19366 3838
rect 3896 -4642 3954 -4630
rect 3896 -4818 3908 -4642
rect 3942 -4818 3954 -4642
rect 3896 -4830 3954 -4818
rect 4154 -4642 4212 -4630
rect 4154 -4818 4166 -4642
rect 4200 -4818 4212 -4642
rect 4154 -4830 4212 -4818
rect 4412 -4642 4470 -4630
rect 4412 -4818 4424 -4642
rect 4458 -4818 4470 -4642
rect 4412 -4830 4470 -4818
rect 4670 -4642 4728 -4630
rect 4670 -4818 4682 -4642
rect 4716 -4818 4728 -4642
rect 4670 -4830 4728 -4818
rect 4928 -4642 4986 -4630
rect 4928 -4818 4940 -4642
rect 4974 -4818 4986 -4642
rect 4928 -4830 4986 -4818
rect 5186 -4642 5244 -4630
rect 5186 -4818 5198 -4642
rect 5232 -4818 5244 -4642
rect 5186 -4830 5244 -4818
rect 5444 -4642 5502 -4630
rect 5444 -4818 5456 -4642
rect 5490 -4818 5502 -4642
rect 5444 -4830 5502 -4818
rect 5702 -4642 5760 -4630
rect 5702 -4818 5714 -4642
rect 5748 -4818 5760 -4642
rect 5702 -4830 5760 -4818
rect 5960 -4642 6018 -4630
rect 5960 -4818 5972 -4642
rect 6006 -4818 6018 -4642
rect 5960 -4830 6018 -4818
rect 6218 -4642 6276 -4630
rect 6218 -4818 6230 -4642
rect 6264 -4818 6276 -4642
rect 6218 -4830 6276 -4818
rect 6476 -4642 6534 -4630
rect 6476 -4818 6488 -4642
rect 6522 -4818 6534 -4642
rect 6476 -4830 6534 -4818
rect 6734 -4642 6792 -4630
rect 6734 -4818 6746 -4642
rect 6780 -4818 6792 -4642
rect 6734 -4830 6792 -4818
rect 6992 -4642 7050 -4630
rect 6992 -4818 7004 -4642
rect 7038 -4818 7050 -4642
rect 6992 -4830 7050 -4818
rect 7250 -4642 7308 -4630
rect 7250 -4818 7262 -4642
rect 7296 -4818 7308 -4642
rect 7250 -4830 7308 -4818
rect 7508 -4642 7566 -4630
rect 7508 -4818 7520 -4642
rect 7554 -4818 7566 -4642
rect 7508 -4830 7566 -4818
rect 15696 -4642 15754 -4630
rect 15696 -4818 15708 -4642
rect 15742 -4818 15754 -4642
rect 15696 -4830 15754 -4818
rect 15954 -4642 16012 -4630
rect 15954 -4818 15966 -4642
rect 16000 -4818 16012 -4642
rect 15954 -4830 16012 -4818
rect 16212 -4642 16270 -4630
rect 16212 -4818 16224 -4642
rect 16258 -4818 16270 -4642
rect 16212 -4830 16270 -4818
rect 16470 -4642 16528 -4630
rect 16470 -4818 16482 -4642
rect 16516 -4818 16528 -4642
rect 16470 -4830 16528 -4818
rect 16728 -4642 16786 -4630
rect 16728 -4818 16740 -4642
rect 16774 -4818 16786 -4642
rect 16728 -4830 16786 -4818
rect 16986 -4642 17044 -4630
rect 16986 -4818 16998 -4642
rect 17032 -4818 17044 -4642
rect 16986 -4830 17044 -4818
rect 17244 -4642 17302 -4630
rect 17244 -4818 17256 -4642
rect 17290 -4818 17302 -4642
rect 17244 -4830 17302 -4818
rect 17502 -4642 17560 -4630
rect 17502 -4818 17514 -4642
rect 17548 -4818 17560 -4642
rect 17502 -4830 17560 -4818
rect 17760 -4642 17818 -4630
rect 17760 -4818 17772 -4642
rect 17806 -4818 17818 -4642
rect 17760 -4830 17818 -4818
rect 18018 -4642 18076 -4630
rect 18018 -4818 18030 -4642
rect 18064 -4818 18076 -4642
rect 18018 -4830 18076 -4818
rect 18276 -4642 18334 -4630
rect 18276 -4818 18288 -4642
rect 18322 -4818 18334 -4642
rect 18276 -4830 18334 -4818
rect 18534 -4642 18592 -4630
rect 18534 -4818 18546 -4642
rect 18580 -4818 18592 -4642
rect 18534 -4830 18592 -4818
rect 18792 -4642 18850 -4630
rect 18792 -4818 18804 -4642
rect 18838 -4818 18850 -4642
rect 18792 -4830 18850 -4818
rect 19050 -4642 19108 -4630
rect 19050 -4818 19062 -4642
rect 19096 -4818 19108 -4642
rect 19050 -4830 19108 -4818
rect 19308 -4642 19366 -4630
rect 19308 -4818 19320 -4642
rect 19354 -4818 19366 -4642
rect 19308 -4830 19366 -4818
<< ndiffc >>
rect 1124 2170 1158 2546
rect 1382 2170 1416 2546
rect 1640 2170 1674 2546
rect 1898 2170 1932 2546
rect 2156 2170 2190 2546
rect 2414 2170 2448 2546
rect 2672 2170 2706 2546
rect 2930 2170 2964 2546
rect 3188 2170 3222 2546
rect 3446 2170 3480 2546
rect 3704 2170 3738 2546
rect 4420 2170 4454 2546
rect 4678 2170 4712 2546
rect 4936 2170 4970 2546
rect 5194 2170 5228 2546
rect 5452 2170 5486 2546
rect 5710 2170 5744 2546
rect 5968 2170 6002 2546
rect 6226 2170 6260 2546
rect 6484 2170 6518 2546
rect 6742 2170 6776 2546
rect 7000 2170 7034 2546
rect 7716 2170 7750 2546
rect 7974 2170 8008 2546
rect 8232 2170 8266 2546
rect 8490 2170 8524 2546
rect 8748 2170 8782 2546
rect 9006 2170 9040 2546
rect 9264 2170 9298 2546
rect 9522 2170 9556 2546
rect 9780 2170 9814 2546
rect 10038 2170 10072 2546
rect 10296 2170 10330 2546
rect 576 1262 610 1438
rect 1434 1262 1468 1438
rect 2292 1262 2326 1438
rect 3150 1262 3184 1438
rect 4008 1262 4042 1438
rect 4866 1262 4900 1438
rect 5724 1262 5758 1438
rect 6582 1262 6616 1438
rect 7440 1262 7474 1438
rect 8298 1262 8332 1438
rect 9156 1262 9190 1438
rect 10014 1262 10048 1438
rect 10872 1262 10906 1438
rect 576 722 610 898
rect 1434 722 1468 898
rect 2292 722 2326 898
rect 3150 722 3184 898
rect 4008 722 4042 898
rect 4866 722 4900 898
rect 5724 722 5758 898
rect 6582 722 6616 898
rect 7440 722 7474 898
rect 8298 722 8332 898
rect 9156 722 9190 898
rect 10014 722 10048 898
rect 10872 722 10906 898
rect 12924 2170 12958 2546
rect 13182 2170 13216 2546
rect 13440 2170 13474 2546
rect 13698 2170 13732 2546
rect 13956 2170 13990 2546
rect 14214 2170 14248 2546
rect 14472 2170 14506 2546
rect 14730 2170 14764 2546
rect 14988 2170 15022 2546
rect 15246 2170 15280 2546
rect 15504 2170 15538 2546
rect 16220 2170 16254 2546
rect 16478 2170 16512 2546
rect 16736 2170 16770 2546
rect 16994 2170 17028 2546
rect 17252 2170 17286 2546
rect 17510 2170 17544 2546
rect 17768 2170 17802 2546
rect 18026 2170 18060 2546
rect 18284 2170 18318 2546
rect 18542 2170 18576 2546
rect 18800 2170 18834 2546
rect 19516 2170 19550 2546
rect 19774 2170 19808 2546
rect 20032 2170 20066 2546
rect 20290 2170 20324 2546
rect 20548 2170 20582 2546
rect 20806 2170 20840 2546
rect 21064 2170 21098 2546
rect 21322 2170 21356 2546
rect 21580 2170 21614 2546
rect 21838 2170 21872 2546
rect 22096 2170 22130 2546
rect 12376 1262 12410 1438
rect 13234 1262 13268 1438
rect 14092 1262 14126 1438
rect 14950 1262 14984 1438
rect 15808 1262 15842 1438
rect 16666 1262 16700 1438
rect 17524 1262 17558 1438
rect 18382 1262 18416 1438
rect 19240 1262 19274 1438
rect 20098 1262 20132 1438
rect 20956 1262 20990 1438
rect 21814 1262 21848 1438
rect 22672 1262 22706 1438
rect 12376 722 12410 898
rect 13234 722 13268 898
rect 14092 722 14126 898
rect 14950 722 14984 898
rect 15808 722 15842 898
rect 16666 722 16700 898
rect 17524 722 17558 898
rect 18382 722 18416 898
rect 19240 722 19274 898
rect 20098 722 20132 898
rect 20956 722 20990 898
rect 21814 722 21848 898
rect 22672 722 22706 898
rect 576 -1702 610 -1526
rect 1434 -1702 1468 -1526
rect 2292 -1702 2326 -1526
rect 3150 -1702 3184 -1526
rect 4008 -1702 4042 -1526
rect 4866 -1702 4900 -1526
rect 5724 -1702 5758 -1526
rect 6582 -1702 6616 -1526
rect 7440 -1702 7474 -1526
rect 8298 -1702 8332 -1526
rect 9156 -1702 9190 -1526
rect 10014 -1702 10048 -1526
rect 10872 -1702 10906 -1526
rect 576 -2242 610 -2066
rect 1434 -2242 1468 -2066
rect 2292 -2242 2326 -2066
rect 3150 -2242 3184 -2066
rect 4008 -2242 4042 -2066
rect 4866 -2242 4900 -2066
rect 5724 -2242 5758 -2066
rect 6582 -2242 6616 -2066
rect 7440 -2242 7474 -2066
rect 8298 -2242 8332 -2066
rect 9156 -2242 9190 -2066
rect 10014 -2242 10048 -2066
rect 10872 -2242 10906 -2066
rect 1124 -3350 1158 -2974
rect 1382 -3350 1416 -2974
rect 1640 -3350 1674 -2974
rect 1898 -3350 1932 -2974
rect 2156 -3350 2190 -2974
rect 2414 -3350 2448 -2974
rect 2672 -3350 2706 -2974
rect 2930 -3350 2964 -2974
rect 3188 -3350 3222 -2974
rect 3446 -3350 3480 -2974
rect 3704 -3350 3738 -2974
rect 4420 -3350 4454 -2974
rect 4678 -3350 4712 -2974
rect 4936 -3350 4970 -2974
rect 5194 -3350 5228 -2974
rect 5452 -3350 5486 -2974
rect 5710 -3350 5744 -2974
rect 5968 -3350 6002 -2974
rect 6226 -3350 6260 -2974
rect 6484 -3350 6518 -2974
rect 6742 -3350 6776 -2974
rect 7000 -3350 7034 -2974
rect 7716 -3350 7750 -2974
rect 7974 -3350 8008 -2974
rect 8232 -3350 8266 -2974
rect 8490 -3350 8524 -2974
rect 8748 -3350 8782 -2974
rect 9006 -3350 9040 -2974
rect 9264 -3350 9298 -2974
rect 9522 -3350 9556 -2974
rect 9780 -3350 9814 -2974
rect 10038 -3350 10072 -2974
rect 10296 -3350 10330 -2974
rect 12376 -1702 12410 -1526
rect 13234 -1702 13268 -1526
rect 14092 -1702 14126 -1526
rect 14950 -1702 14984 -1526
rect 15808 -1702 15842 -1526
rect 16666 -1702 16700 -1526
rect 17524 -1702 17558 -1526
rect 18382 -1702 18416 -1526
rect 19240 -1702 19274 -1526
rect 20098 -1702 20132 -1526
rect 20956 -1702 20990 -1526
rect 21814 -1702 21848 -1526
rect 22672 -1702 22706 -1526
rect 12376 -2242 12410 -2066
rect 13234 -2242 13268 -2066
rect 14092 -2242 14126 -2066
rect 14950 -2242 14984 -2066
rect 15808 -2242 15842 -2066
rect 16666 -2242 16700 -2066
rect 17524 -2242 17558 -2066
rect 18382 -2242 18416 -2066
rect 19240 -2242 19274 -2066
rect 20098 -2242 20132 -2066
rect 20956 -2242 20990 -2066
rect 21814 -2242 21848 -2066
rect 22672 -2242 22706 -2066
rect 12924 -3350 12958 -2974
rect 13182 -3350 13216 -2974
rect 13440 -3350 13474 -2974
rect 13698 -3350 13732 -2974
rect 13956 -3350 13990 -2974
rect 14214 -3350 14248 -2974
rect 14472 -3350 14506 -2974
rect 14730 -3350 14764 -2974
rect 14988 -3350 15022 -2974
rect 15246 -3350 15280 -2974
rect 15504 -3350 15538 -2974
rect 16220 -3350 16254 -2974
rect 16478 -3350 16512 -2974
rect 16736 -3350 16770 -2974
rect 16994 -3350 17028 -2974
rect 17252 -3350 17286 -2974
rect 17510 -3350 17544 -2974
rect 17768 -3350 17802 -2974
rect 18026 -3350 18060 -2974
rect 18284 -3350 18318 -2974
rect 18542 -3350 18576 -2974
rect 18800 -3350 18834 -2974
rect 19516 -3350 19550 -2974
rect 19774 -3350 19808 -2974
rect 20032 -3350 20066 -2974
rect 20290 -3350 20324 -2974
rect 20548 -3350 20582 -2974
rect 20806 -3350 20840 -2974
rect 21064 -3350 21098 -2974
rect 21322 -3350 21356 -2974
rect 21580 -3350 21614 -2974
rect 21838 -3350 21872 -2974
rect 22096 -3350 22130 -2974
<< pdiffc >>
rect 3908 3838 3942 4014
rect 4166 3838 4200 4014
rect 4424 3838 4458 4014
rect 4682 3838 4716 4014
rect 4940 3838 4974 4014
rect 5198 3838 5232 4014
rect 5456 3838 5490 4014
rect 5714 3838 5748 4014
rect 5972 3838 6006 4014
rect 6230 3838 6264 4014
rect 6488 3838 6522 4014
rect 6746 3838 6780 4014
rect 7004 3838 7038 4014
rect 7262 3838 7296 4014
rect 7520 3838 7554 4014
rect 15708 3838 15742 4014
rect 15966 3838 16000 4014
rect 16224 3838 16258 4014
rect 16482 3838 16516 4014
rect 16740 3838 16774 4014
rect 16998 3838 17032 4014
rect 17256 3838 17290 4014
rect 17514 3838 17548 4014
rect 17772 3838 17806 4014
rect 18030 3838 18064 4014
rect 18288 3838 18322 4014
rect 18546 3838 18580 4014
rect 18804 3838 18838 4014
rect 19062 3838 19096 4014
rect 19320 3838 19354 4014
rect 3908 -4818 3942 -4642
rect 4166 -4818 4200 -4642
rect 4424 -4818 4458 -4642
rect 4682 -4818 4716 -4642
rect 4940 -4818 4974 -4642
rect 5198 -4818 5232 -4642
rect 5456 -4818 5490 -4642
rect 5714 -4818 5748 -4642
rect 5972 -4818 6006 -4642
rect 6230 -4818 6264 -4642
rect 6488 -4818 6522 -4642
rect 6746 -4818 6780 -4642
rect 7004 -4818 7038 -4642
rect 7262 -4818 7296 -4642
rect 7520 -4818 7554 -4642
rect 15708 -4818 15742 -4642
rect 15966 -4818 16000 -4642
rect 16224 -4818 16258 -4642
rect 16482 -4818 16516 -4642
rect 16740 -4818 16774 -4642
rect 16998 -4818 17032 -4642
rect 17256 -4818 17290 -4642
rect 17514 -4818 17548 -4642
rect 17772 -4818 17806 -4642
rect 18030 -4818 18064 -4642
rect 18288 -4818 18322 -4642
rect 18546 -4818 18580 -4642
rect 18804 -4818 18838 -4642
rect 19062 -4818 19096 -4642
rect 19320 -4818 19354 -4642
<< psubdiff >>
rect 66 3018 228 3118
rect 11248 3018 11410 3118
rect 66 2956 166 3018
rect 11310 2956 11410 3018
rect 66 -186 166 -124
rect 11310 -186 11410 -124
rect 66 -286 228 -186
rect 11248 -286 11410 -186
rect 11866 3018 12028 3118
rect 23048 3018 23210 3118
rect 11866 2956 11966 3018
rect 23110 2956 23210 3018
rect 11866 -186 11966 -124
rect 23110 -186 23210 -124
rect 11866 -286 12028 -186
rect 23048 -286 23210 -186
rect 66 -618 228 -518
rect 11248 -618 11410 -518
rect 66 -680 166 -618
rect 11310 -680 11410 -618
rect 66 -3822 166 -3760
rect 11310 -3822 11410 -3760
rect 66 -3922 228 -3822
rect 11248 -3922 11410 -3822
rect 11866 -618 12028 -518
rect 23048 -618 23210 -518
rect 11866 -680 11966 -618
rect 23110 -680 23210 -618
rect 11866 -3822 11966 -3760
rect 23110 -3822 23210 -3760
rect 11866 -3922 12028 -3822
rect 23048 -3922 23210 -3822
<< nsubdiff >>
rect 66 5038 228 5138
rect 11248 5038 11410 5138
rect 66 4976 166 5038
rect 11310 4976 11410 5038
rect 66 3454 166 3516
rect 11310 3454 11410 3516
rect 66 3354 228 3454
rect 11248 3354 11410 3454
rect 11866 5038 12028 5138
rect 23048 5038 23210 5138
rect 11866 4976 11966 5038
rect 23110 4976 23210 5038
rect 11866 3454 11966 3516
rect 23110 3454 23210 3516
rect 11866 3354 12028 3454
rect 23048 3354 23210 3454
rect 66 -4258 228 -4158
rect 11248 -4258 11410 -4158
rect 66 -4320 166 -4258
rect 11310 -4320 11410 -4258
rect 66 -5842 166 -5780
rect 11310 -5842 11410 -5780
rect 66 -5942 228 -5842
rect 11248 -5942 11410 -5842
rect 11866 -4258 12028 -4158
rect 23048 -4258 23210 -4158
rect 11866 -4320 11966 -4258
rect 23110 -4320 23210 -4258
rect 11866 -5842 11966 -5780
rect 23110 -5842 23210 -5780
rect 11866 -5942 12028 -5842
rect 23048 -5942 23210 -5842
<< psubdiffcont >>
rect 228 3018 11248 3118
rect 66 -124 166 2956
rect 11310 -124 11410 2956
rect 228 -286 11248 -186
rect 12028 3018 23048 3118
rect 11866 -124 11966 2956
rect 23110 -124 23210 2956
rect 12028 -286 23048 -186
rect 228 -618 11248 -518
rect 66 -3760 166 -680
rect 11310 -3760 11410 -680
rect 228 -3922 11248 -3822
rect 12028 -618 23048 -518
rect 11866 -3760 11966 -680
rect 23110 -3760 23210 -680
rect 12028 -3922 23048 -3822
<< nsubdiffcont >>
rect 228 5038 11248 5138
rect 66 3516 166 4976
rect 11310 3516 11410 4976
rect 228 3354 11248 3454
rect 12028 5038 23048 5138
rect 11866 3516 11966 4976
rect 23110 3516 23210 4976
rect 12028 3354 23048 3454
rect 228 -4258 11248 -4158
rect 66 -5780 166 -4320
rect 11310 -5780 11410 -4320
rect 228 -5942 11248 -5842
rect 12028 -4258 23048 -4158
rect 11866 -5780 11966 -4320
rect 23110 -5780 23210 -4320
rect 12028 -5942 23048 -5842
<< poly >>
rect 3988 4107 4120 4123
rect 3988 4090 4004 4107
rect 3954 4073 4004 4090
rect 4104 4090 4120 4107
rect 4246 4107 4378 4123
rect 4246 4090 4262 4107
rect 4104 4073 4154 4090
rect 3954 4026 4154 4073
rect 4212 4073 4262 4090
rect 4362 4090 4378 4107
rect 4504 4107 4636 4123
rect 4504 4090 4520 4107
rect 4362 4073 4412 4090
rect 4212 4026 4412 4073
rect 4470 4073 4520 4090
rect 4620 4090 4636 4107
rect 4762 4107 4894 4123
rect 4762 4090 4778 4107
rect 4620 4073 4670 4090
rect 4470 4026 4670 4073
rect 4728 4073 4778 4090
rect 4878 4090 4894 4107
rect 5020 4107 5152 4123
rect 5020 4090 5036 4107
rect 4878 4073 4928 4090
rect 4728 4026 4928 4073
rect 4986 4073 5036 4090
rect 5136 4090 5152 4107
rect 5278 4107 5410 4123
rect 5278 4090 5294 4107
rect 5136 4073 5186 4090
rect 4986 4026 5186 4073
rect 5244 4073 5294 4090
rect 5394 4090 5410 4107
rect 5536 4107 5668 4123
rect 5536 4090 5552 4107
rect 5394 4073 5444 4090
rect 5244 4026 5444 4073
rect 5502 4073 5552 4090
rect 5652 4090 5668 4107
rect 5794 4107 5926 4123
rect 5794 4090 5810 4107
rect 5652 4073 5702 4090
rect 5502 4026 5702 4073
rect 5760 4073 5810 4090
rect 5910 4090 5926 4107
rect 6052 4107 6184 4123
rect 6052 4090 6068 4107
rect 5910 4073 5960 4090
rect 5760 4026 5960 4073
rect 6018 4073 6068 4090
rect 6168 4090 6184 4107
rect 6310 4107 6442 4123
rect 6310 4090 6326 4107
rect 6168 4073 6218 4090
rect 6018 4026 6218 4073
rect 6276 4073 6326 4090
rect 6426 4090 6442 4107
rect 6568 4107 6700 4123
rect 6568 4090 6584 4107
rect 6426 4073 6476 4090
rect 6276 4026 6476 4073
rect 6534 4073 6584 4090
rect 6684 4090 6700 4107
rect 6826 4107 6958 4123
rect 6826 4090 6842 4107
rect 6684 4073 6734 4090
rect 6534 4026 6734 4073
rect 6792 4073 6842 4090
rect 6942 4090 6958 4107
rect 7084 4107 7216 4123
rect 7084 4090 7100 4107
rect 6942 4073 6992 4090
rect 6792 4026 6992 4073
rect 7050 4073 7100 4090
rect 7200 4090 7216 4107
rect 7342 4107 7474 4123
rect 7342 4090 7358 4107
rect 7200 4073 7250 4090
rect 7050 4026 7250 4073
rect 7308 4073 7358 4090
rect 7458 4090 7474 4107
rect 7458 4073 7508 4090
rect 7308 4026 7508 4073
rect 3954 3779 4154 3826
rect 3954 3762 4004 3779
rect 3988 3745 4004 3762
rect 4104 3762 4154 3779
rect 4212 3779 4412 3826
rect 4212 3762 4262 3779
rect 4104 3745 4120 3762
rect 3988 3729 4120 3745
rect 4246 3745 4262 3762
rect 4362 3762 4412 3779
rect 4470 3779 4670 3826
rect 4470 3762 4520 3779
rect 4362 3745 4378 3762
rect 4246 3729 4378 3745
rect 4504 3745 4520 3762
rect 4620 3762 4670 3779
rect 4728 3779 4928 3826
rect 4728 3762 4778 3779
rect 4620 3745 4636 3762
rect 4504 3729 4636 3745
rect 4762 3745 4778 3762
rect 4878 3762 4928 3779
rect 4986 3779 5186 3826
rect 4986 3762 5036 3779
rect 4878 3745 4894 3762
rect 4762 3729 4894 3745
rect 5020 3745 5036 3762
rect 5136 3762 5186 3779
rect 5244 3779 5444 3826
rect 5244 3762 5294 3779
rect 5136 3745 5152 3762
rect 5020 3729 5152 3745
rect 5278 3745 5294 3762
rect 5394 3762 5444 3779
rect 5502 3779 5702 3826
rect 5502 3762 5552 3779
rect 5394 3745 5410 3762
rect 5278 3729 5410 3745
rect 5536 3745 5552 3762
rect 5652 3762 5702 3779
rect 5760 3779 5960 3826
rect 5760 3762 5810 3779
rect 5652 3745 5668 3762
rect 5536 3729 5668 3745
rect 5794 3745 5810 3762
rect 5910 3762 5960 3779
rect 6018 3779 6218 3826
rect 6018 3762 6068 3779
rect 5910 3745 5926 3762
rect 5794 3729 5926 3745
rect 6052 3745 6068 3762
rect 6168 3762 6218 3779
rect 6276 3779 6476 3826
rect 6276 3762 6326 3779
rect 6168 3745 6184 3762
rect 6052 3729 6184 3745
rect 6310 3745 6326 3762
rect 6426 3762 6476 3779
rect 6534 3779 6734 3826
rect 6534 3762 6584 3779
rect 6426 3745 6442 3762
rect 6310 3729 6442 3745
rect 6568 3745 6584 3762
rect 6684 3762 6734 3779
rect 6792 3779 6992 3826
rect 6792 3762 6842 3779
rect 6684 3745 6700 3762
rect 6568 3729 6700 3745
rect 6826 3745 6842 3762
rect 6942 3762 6992 3779
rect 7050 3779 7250 3826
rect 7050 3762 7100 3779
rect 6942 3745 6958 3762
rect 6826 3729 6958 3745
rect 7084 3745 7100 3762
rect 7200 3762 7250 3779
rect 7308 3779 7508 3826
rect 7308 3762 7358 3779
rect 7200 3745 7216 3762
rect 7084 3729 7216 3745
rect 7342 3745 7358 3762
rect 7458 3762 7508 3779
rect 7458 3745 7474 3762
rect 7342 3729 7474 3745
rect 15788 4107 15920 4123
rect 15788 4090 15804 4107
rect 15754 4073 15804 4090
rect 15904 4090 15920 4107
rect 16046 4107 16178 4123
rect 16046 4090 16062 4107
rect 15904 4073 15954 4090
rect 15754 4026 15954 4073
rect 16012 4073 16062 4090
rect 16162 4090 16178 4107
rect 16304 4107 16436 4123
rect 16304 4090 16320 4107
rect 16162 4073 16212 4090
rect 16012 4026 16212 4073
rect 16270 4073 16320 4090
rect 16420 4090 16436 4107
rect 16562 4107 16694 4123
rect 16562 4090 16578 4107
rect 16420 4073 16470 4090
rect 16270 4026 16470 4073
rect 16528 4073 16578 4090
rect 16678 4090 16694 4107
rect 16820 4107 16952 4123
rect 16820 4090 16836 4107
rect 16678 4073 16728 4090
rect 16528 4026 16728 4073
rect 16786 4073 16836 4090
rect 16936 4090 16952 4107
rect 17078 4107 17210 4123
rect 17078 4090 17094 4107
rect 16936 4073 16986 4090
rect 16786 4026 16986 4073
rect 17044 4073 17094 4090
rect 17194 4090 17210 4107
rect 17336 4107 17468 4123
rect 17336 4090 17352 4107
rect 17194 4073 17244 4090
rect 17044 4026 17244 4073
rect 17302 4073 17352 4090
rect 17452 4090 17468 4107
rect 17594 4107 17726 4123
rect 17594 4090 17610 4107
rect 17452 4073 17502 4090
rect 17302 4026 17502 4073
rect 17560 4073 17610 4090
rect 17710 4090 17726 4107
rect 17852 4107 17984 4123
rect 17852 4090 17868 4107
rect 17710 4073 17760 4090
rect 17560 4026 17760 4073
rect 17818 4073 17868 4090
rect 17968 4090 17984 4107
rect 18110 4107 18242 4123
rect 18110 4090 18126 4107
rect 17968 4073 18018 4090
rect 17818 4026 18018 4073
rect 18076 4073 18126 4090
rect 18226 4090 18242 4107
rect 18368 4107 18500 4123
rect 18368 4090 18384 4107
rect 18226 4073 18276 4090
rect 18076 4026 18276 4073
rect 18334 4073 18384 4090
rect 18484 4090 18500 4107
rect 18626 4107 18758 4123
rect 18626 4090 18642 4107
rect 18484 4073 18534 4090
rect 18334 4026 18534 4073
rect 18592 4073 18642 4090
rect 18742 4090 18758 4107
rect 18884 4107 19016 4123
rect 18884 4090 18900 4107
rect 18742 4073 18792 4090
rect 18592 4026 18792 4073
rect 18850 4073 18900 4090
rect 19000 4090 19016 4107
rect 19142 4107 19274 4123
rect 19142 4090 19158 4107
rect 19000 4073 19050 4090
rect 18850 4026 19050 4073
rect 19108 4073 19158 4090
rect 19258 4090 19274 4107
rect 19258 4073 19308 4090
rect 19108 4026 19308 4073
rect 15754 3779 15954 3826
rect 15754 3762 15804 3779
rect 15788 3745 15804 3762
rect 15904 3762 15954 3779
rect 16012 3779 16212 3826
rect 16012 3762 16062 3779
rect 15904 3745 15920 3762
rect 15788 3729 15920 3745
rect 16046 3745 16062 3762
rect 16162 3762 16212 3779
rect 16270 3779 16470 3826
rect 16270 3762 16320 3779
rect 16162 3745 16178 3762
rect 16046 3729 16178 3745
rect 16304 3745 16320 3762
rect 16420 3762 16470 3779
rect 16528 3779 16728 3826
rect 16528 3762 16578 3779
rect 16420 3745 16436 3762
rect 16304 3729 16436 3745
rect 16562 3745 16578 3762
rect 16678 3762 16728 3779
rect 16786 3779 16986 3826
rect 16786 3762 16836 3779
rect 16678 3745 16694 3762
rect 16562 3729 16694 3745
rect 16820 3745 16836 3762
rect 16936 3762 16986 3779
rect 17044 3779 17244 3826
rect 17044 3762 17094 3779
rect 16936 3745 16952 3762
rect 16820 3729 16952 3745
rect 17078 3745 17094 3762
rect 17194 3762 17244 3779
rect 17302 3779 17502 3826
rect 17302 3762 17352 3779
rect 17194 3745 17210 3762
rect 17078 3729 17210 3745
rect 17336 3745 17352 3762
rect 17452 3762 17502 3779
rect 17560 3779 17760 3826
rect 17560 3762 17610 3779
rect 17452 3745 17468 3762
rect 17336 3729 17468 3745
rect 17594 3745 17610 3762
rect 17710 3762 17760 3779
rect 17818 3779 18018 3826
rect 17818 3762 17868 3779
rect 17710 3745 17726 3762
rect 17594 3729 17726 3745
rect 17852 3745 17868 3762
rect 17968 3762 18018 3779
rect 18076 3779 18276 3826
rect 18076 3762 18126 3779
rect 17968 3745 17984 3762
rect 17852 3729 17984 3745
rect 18110 3745 18126 3762
rect 18226 3762 18276 3779
rect 18334 3779 18534 3826
rect 18334 3762 18384 3779
rect 18226 3745 18242 3762
rect 18110 3729 18242 3745
rect 18368 3745 18384 3762
rect 18484 3762 18534 3779
rect 18592 3779 18792 3826
rect 18592 3762 18642 3779
rect 18484 3745 18500 3762
rect 18368 3729 18500 3745
rect 18626 3745 18642 3762
rect 18742 3762 18792 3779
rect 18850 3779 19050 3826
rect 18850 3762 18900 3779
rect 18742 3745 18758 3762
rect 18626 3729 18758 3745
rect 18884 3745 18900 3762
rect 19000 3762 19050 3779
rect 19108 3779 19308 3826
rect 19108 3762 19158 3779
rect 19000 3745 19016 3762
rect 18884 3729 19016 3745
rect 19142 3745 19158 3762
rect 19258 3762 19308 3779
rect 19258 3745 19274 3762
rect 19142 3729 19274 3745
rect 1204 2630 1336 2646
rect 1204 2613 1220 2630
rect 1170 2596 1220 2613
rect 1320 2613 1336 2630
rect 1462 2630 1594 2646
rect 1462 2613 1478 2630
rect 1320 2596 1370 2613
rect 1170 2558 1370 2596
rect 1428 2596 1478 2613
rect 1578 2613 1594 2630
rect 1720 2630 1852 2646
rect 1720 2613 1736 2630
rect 1578 2596 1628 2613
rect 1428 2558 1628 2596
rect 1686 2596 1736 2613
rect 1836 2613 1852 2630
rect 1978 2630 2110 2646
rect 1978 2613 1994 2630
rect 1836 2596 1886 2613
rect 1686 2558 1886 2596
rect 1944 2596 1994 2613
rect 2094 2613 2110 2630
rect 2236 2630 2368 2646
rect 2236 2613 2252 2630
rect 2094 2596 2144 2613
rect 1944 2558 2144 2596
rect 2202 2596 2252 2613
rect 2352 2613 2368 2630
rect 2494 2630 2626 2646
rect 2494 2613 2510 2630
rect 2352 2596 2402 2613
rect 2202 2558 2402 2596
rect 2460 2596 2510 2613
rect 2610 2613 2626 2630
rect 2752 2630 2884 2646
rect 2752 2613 2768 2630
rect 2610 2596 2660 2613
rect 2460 2558 2660 2596
rect 2718 2596 2768 2613
rect 2868 2613 2884 2630
rect 3010 2630 3142 2646
rect 3010 2613 3026 2630
rect 2868 2596 2918 2613
rect 2718 2558 2918 2596
rect 2976 2596 3026 2613
rect 3126 2613 3142 2630
rect 3268 2630 3400 2646
rect 3268 2613 3284 2630
rect 3126 2596 3176 2613
rect 2976 2558 3176 2596
rect 3234 2596 3284 2613
rect 3384 2613 3400 2630
rect 3526 2630 3658 2646
rect 3526 2613 3542 2630
rect 3384 2596 3434 2613
rect 3234 2558 3434 2596
rect 3492 2596 3542 2613
rect 3642 2613 3658 2630
rect 4500 2630 4632 2646
rect 4500 2613 4516 2630
rect 3642 2596 3692 2613
rect 3492 2558 3692 2596
rect 4466 2596 4516 2613
rect 4616 2613 4632 2630
rect 4758 2630 4890 2646
rect 4758 2613 4774 2630
rect 4616 2596 4666 2613
rect 4466 2558 4666 2596
rect 4724 2596 4774 2613
rect 4874 2613 4890 2630
rect 5016 2630 5148 2646
rect 5016 2613 5032 2630
rect 4874 2596 4924 2613
rect 4724 2558 4924 2596
rect 4982 2596 5032 2613
rect 5132 2613 5148 2630
rect 5274 2630 5406 2646
rect 5274 2613 5290 2630
rect 5132 2596 5182 2613
rect 4982 2558 5182 2596
rect 5240 2596 5290 2613
rect 5390 2613 5406 2630
rect 5532 2630 5664 2646
rect 5532 2613 5548 2630
rect 5390 2596 5440 2613
rect 5240 2558 5440 2596
rect 5498 2596 5548 2613
rect 5648 2613 5664 2630
rect 5790 2630 5922 2646
rect 5790 2613 5806 2630
rect 5648 2596 5698 2613
rect 5498 2558 5698 2596
rect 5756 2596 5806 2613
rect 5906 2613 5922 2630
rect 6048 2630 6180 2646
rect 6048 2613 6064 2630
rect 5906 2596 5956 2613
rect 5756 2558 5956 2596
rect 6014 2596 6064 2613
rect 6164 2613 6180 2630
rect 6306 2630 6438 2646
rect 6306 2613 6322 2630
rect 6164 2596 6214 2613
rect 6014 2558 6214 2596
rect 6272 2596 6322 2613
rect 6422 2613 6438 2630
rect 6564 2630 6696 2646
rect 6564 2613 6580 2630
rect 6422 2596 6472 2613
rect 6272 2558 6472 2596
rect 6530 2596 6580 2613
rect 6680 2613 6696 2630
rect 6822 2630 6954 2646
rect 6822 2613 6838 2630
rect 6680 2596 6730 2613
rect 6530 2558 6730 2596
rect 6788 2596 6838 2613
rect 6938 2613 6954 2630
rect 7796 2630 7928 2646
rect 7796 2613 7812 2630
rect 6938 2596 6988 2613
rect 6788 2558 6988 2596
rect 7762 2596 7812 2613
rect 7912 2613 7928 2630
rect 8054 2630 8186 2646
rect 8054 2613 8070 2630
rect 7912 2596 7962 2613
rect 7762 2558 7962 2596
rect 8020 2596 8070 2613
rect 8170 2613 8186 2630
rect 8312 2630 8444 2646
rect 8312 2613 8328 2630
rect 8170 2596 8220 2613
rect 8020 2558 8220 2596
rect 8278 2596 8328 2613
rect 8428 2613 8444 2630
rect 8570 2630 8702 2646
rect 8570 2613 8586 2630
rect 8428 2596 8478 2613
rect 8278 2558 8478 2596
rect 8536 2596 8586 2613
rect 8686 2613 8702 2630
rect 8828 2630 8960 2646
rect 8828 2613 8844 2630
rect 8686 2596 8736 2613
rect 8536 2558 8736 2596
rect 8794 2596 8844 2613
rect 8944 2613 8960 2630
rect 9086 2630 9218 2646
rect 9086 2613 9102 2630
rect 8944 2596 8994 2613
rect 8794 2558 8994 2596
rect 9052 2596 9102 2613
rect 9202 2613 9218 2630
rect 9344 2630 9476 2646
rect 9344 2613 9360 2630
rect 9202 2596 9252 2613
rect 9052 2558 9252 2596
rect 9310 2596 9360 2613
rect 9460 2613 9476 2630
rect 9602 2630 9734 2646
rect 9602 2613 9618 2630
rect 9460 2596 9510 2613
rect 9310 2558 9510 2596
rect 9568 2596 9618 2613
rect 9718 2613 9734 2630
rect 9860 2630 9992 2646
rect 9860 2613 9876 2630
rect 9718 2596 9768 2613
rect 9568 2558 9768 2596
rect 9826 2596 9876 2613
rect 9976 2613 9992 2630
rect 10118 2630 10250 2646
rect 10118 2613 10134 2630
rect 9976 2596 10026 2613
rect 9826 2558 10026 2596
rect 10084 2596 10134 2613
rect 10234 2613 10250 2630
rect 10234 2596 10284 2613
rect 10084 2558 10284 2596
rect 1170 2120 1370 2158
rect 1170 2103 1220 2120
rect 1204 2086 1220 2103
rect 1320 2103 1370 2120
rect 1428 2120 1628 2158
rect 1428 2103 1478 2120
rect 1320 2086 1336 2103
rect 1204 2070 1336 2086
rect 1462 2086 1478 2103
rect 1578 2103 1628 2120
rect 1686 2120 1886 2158
rect 1686 2103 1736 2120
rect 1578 2086 1594 2103
rect 1462 2070 1594 2086
rect 1720 2086 1736 2103
rect 1836 2103 1886 2120
rect 1944 2120 2144 2158
rect 1944 2103 1994 2120
rect 1836 2086 1852 2103
rect 1720 2070 1852 2086
rect 1978 2086 1994 2103
rect 2094 2103 2144 2120
rect 2202 2120 2402 2158
rect 2202 2103 2252 2120
rect 2094 2086 2110 2103
rect 1978 2070 2110 2086
rect 2236 2086 2252 2103
rect 2352 2103 2402 2120
rect 2460 2120 2660 2158
rect 2460 2103 2510 2120
rect 2352 2086 2368 2103
rect 2236 2070 2368 2086
rect 2494 2086 2510 2103
rect 2610 2103 2660 2120
rect 2718 2120 2918 2158
rect 2718 2103 2768 2120
rect 2610 2086 2626 2103
rect 2494 2070 2626 2086
rect 2752 2086 2768 2103
rect 2868 2103 2918 2120
rect 2976 2120 3176 2158
rect 2976 2103 3026 2120
rect 2868 2086 2884 2103
rect 2752 2070 2884 2086
rect 3010 2086 3026 2103
rect 3126 2103 3176 2120
rect 3234 2120 3434 2158
rect 3234 2103 3284 2120
rect 3126 2086 3142 2103
rect 3010 2070 3142 2086
rect 3268 2086 3284 2103
rect 3384 2103 3434 2120
rect 3492 2120 3692 2158
rect 3492 2103 3542 2120
rect 3384 2086 3400 2103
rect 3268 2070 3400 2086
rect 3526 2086 3542 2103
rect 3642 2103 3692 2120
rect 4466 2120 4666 2158
rect 4466 2103 4516 2120
rect 3642 2086 3658 2103
rect 3526 2070 3658 2086
rect 4500 2086 4516 2103
rect 4616 2103 4666 2120
rect 4724 2120 4924 2158
rect 4724 2103 4774 2120
rect 4616 2086 4632 2103
rect 4500 2070 4632 2086
rect 4758 2086 4774 2103
rect 4874 2103 4924 2120
rect 4982 2120 5182 2158
rect 4982 2103 5032 2120
rect 4874 2086 4890 2103
rect 4758 2070 4890 2086
rect 5016 2086 5032 2103
rect 5132 2103 5182 2120
rect 5240 2120 5440 2158
rect 5240 2103 5290 2120
rect 5132 2086 5148 2103
rect 5016 2070 5148 2086
rect 5274 2086 5290 2103
rect 5390 2103 5440 2120
rect 5498 2120 5698 2158
rect 5498 2103 5548 2120
rect 5390 2086 5406 2103
rect 5274 2070 5406 2086
rect 5532 2086 5548 2103
rect 5648 2103 5698 2120
rect 5756 2120 5956 2158
rect 5756 2103 5806 2120
rect 5648 2086 5664 2103
rect 5532 2070 5664 2086
rect 5790 2086 5806 2103
rect 5906 2103 5956 2120
rect 6014 2120 6214 2158
rect 6014 2103 6064 2120
rect 5906 2086 5922 2103
rect 5790 2070 5922 2086
rect 6048 2086 6064 2103
rect 6164 2103 6214 2120
rect 6272 2120 6472 2158
rect 6272 2103 6322 2120
rect 6164 2086 6180 2103
rect 6048 2070 6180 2086
rect 6306 2086 6322 2103
rect 6422 2103 6472 2120
rect 6530 2120 6730 2158
rect 6530 2103 6580 2120
rect 6422 2086 6438 2103
rect 6306 2070 6438 2086
rect 6564 2086 6580 2103
rect 6680 2103 6730 2120
rect 6788 2120 6988 2158
rect 6788 2103 6838 2120
rect 6680 2086 6696 2103
rect 6564 2070 6696 2086
rect 6822 2086 6838 2103
rect 6938 2103 6988 2120
rect 7762 2120 7962 2158
rect 7762 2103 7812 2120
rect 6938 2086 6954 2103
rect 6822 2070 6954 2086
rect 7796 2086 7812 2103
rect 7912 2103 7962 2120
rect 8020 2120 8220 2158
rect 8020 2103 8070 2120
rect 7912 2086 7928 2103
rect 7796 2070 7928 2086
rect 8054 2086 8070 2103
rect 8170 2103 8220 2120
rect 8278 2120 8478 2158
rect 8278 2103 8328 2120
rect 8170 2086 8186 2103
rect 8054 2070 8186 2086
rect 8312 2086 8328 2103
rect 8428 2103 8478 2120
rect 8536 2120 8736 2158
rect 8536 2103 8586 2120
rect 8428 2086 8444 2103
rect 8312 2070 8444 2086
rect 8570 2086 8586 2103
rect 8686 2103 8736 2120
rect 8794 2120 8994 2158
rect 8794 2103 8844 2120
rect 8686 2086 8702 2103
rect 8570 2070 8702 2086
rect 8828 2086 8844 2103
rect 8944 2103 8994 2120
rect 9052 2120 9252 2158
rect 9052 2103 9102 2120
rect 8944 2086 8960 2103
rect 8828 2070 8960 2086
rect 9086 2086 9102 2103
rect 9202 2103 9252 2120
rect 9310 2120 9510 2158
rect 9310 2103 9360 2120
rect 9202 2086 9218 2103
rect 9086 2070 9218 2086
rect 9344 2086 9360 2103
rect 9460 2103 9510 2120
rect 9568 2120 9768 2158
rect 9568 2103 9618 2120
rect 9460 2086 9476 2103
rect 9344 2070 9476 2086
rect 9602 2086 9618 2103
rect 9718 2103 9768 2120
rect 9826 2120 10026 2158
rect 9826 2103 9876 2120
rect 9718 2086 9734 2103
rect 9602 2070 9734 2086
rect 9860 2086 9876 2103
rect 9976 2103 10026 2120
rect 10084 2120 10284 2158
rect 10084 2103 10134 2120
rect 9976 2086 9992 2103
rect 9860 2070 9992 2086
rect 10118 2086 10134 2103
rect 10234 2103 10284 2120
rect 10234 2086 10250 2103
rect 10118 2070 10250 2086
rect 776 1522 1268 1538
rect 776 1505 792 1522
rect 622 1488 792 1505
rect 1252 1505 1268 1522
rect 1634 1522 2126 1538
rect 1634 1505 1650 1522
rect 1252 1488 1422 1505
rect 622 1450 1422 1488
rect 1480 1488 1650 1505
rect 2110 1505 2126 1522
rect 2492 1522 2984 1538
rect 2492 1505 2508 1522
rect 2110 1488 2280 1505
rect 1480 1450 2280 1488
rect 2338 1488 2508 1505
rect 2968 1505 2984 1522
rect 3350 1522 3842 1538
rect 3350 1505 3366 1522
rect 2968 1488 3138 1505
rect 2338 1450 3138 1488
rect 3196 1488 3366 1505
rect 3826 1505 3842 1522
rect 4208 1522 4700 1538
rect 4208 1505 4224 1522
rect 3826 1488 3996 1505
rect 3196 1450 3996 1488
rect 4054 1488 4224 1505
rect 4684 1505 4700 1522
rect 5066 1522 5558 1538
rect 5066 1505 5082 1522
rect 4684 1488 4854 1505
rect 4054 1450 4854 1488
rect 4912 1488 5082 1505
rect 5542 1505 5558 1522
rect 5924 1522 6416 1538
rect 5924 1505 5940 1522
rect 5542 1488 5712 1505
rect 4912 1450 5712 1488
rect 5770 1488 5940 1505
rect 6400 1505 6416 1522
rect 6782 1522 7274 1538
rect 6782 1505 6798 1522
rect 6400 1488 6570 1505
rect 5770 1450 6570 1488
rect 6628 1488 6798 1505
rect 7258 1505 7274 1522
rect 7640 1522 8132 1538
rect 7640 1505 7656 1522
rect 7258 1488 7428 1505
rect 6628 1450 7428 1488
rect 7486 1488 7656 1505
rect 8116 1505 8132 1522
rect 8498 1522 8990 1538
rect 8498 1505 8514 1522
rect 8116 1488 8286 1505
rect 7486 1450 8286 1488
rect 8344 1488 8514 1505
rect 8974 1505 8990 1522
rect 9356 1522 9848 1538
rect 9356 1505 9372 1522
rect 8974 1488 9144 1505
rect 8344 1450 9144 1488
rect 9202 1488 9372 1505
rect 9832 1505 9848 1522
rect 10214 1522 10706 1538
rect 10214 1505 10230 1522
rect 9832 1488 10002 1505
rect 9202 1450 10002 1488
rect 10060 1488 10230 1505
rect 10690 1505 10706 1522
rect 10690 1488 10860 1505
rect 10060 1450 10860 1488
rect 622 1212 1422 1250
rect 622 1195 792 1212
rect 776 1178 792 1195
rect 1252 1195 1422 1212
rect 1480 1212 2280 1250
rect 1480 1195 1650 1212
rect 1252 1178 1268 1195
rect 776 1162 1268 1178
rect 1634 1178 1650 1195
rect 2110 1195 2280 1212
rect 2338 1212 3138 1250
rect 2338 1195 2508 1212
rect 2110 1178 2126 1195
rect 1634 1162 2126 1178
rect 2492 1178 2508 1195
rect 2968 1195 3138 1212
rect 3196 1212 3996 1250
rect 3196 1195 3366 1212
rect 2968 1178 2984 1195
rect 2492 1162 2984 1178
rect 3350 1178 3366 1195
rect 3826 1195 3996 1212
rect 4054 1212 4854 1250
rect 4054 1195 4224 1212
rect 3826 1178 3842 1195
rect 3350 1162 3842 1178
rect 4208 1178 4224 1195
rect 4684 1195 4854 1212
rect 4912 1212 5712 1250
rect 4912 1195 5082 1212
rect 4684 1178 4700 1195
rect 4208 1162 4700 1178
rect 5066 1178 5082 1195
rect 5542 1195 5712 1212
rect 5770 1212 6570 1250
rect 5770 1195 5940 1212
rect 5542 1178 5558 1195
rect 5066 1162 5558 1178
rect 5924 1178 5940 1195
rect 6400 1195 6570 1212
rect 6628 1212 7428 1250
rect 6628 1195 6798 1212
rect 6400 1178 6416 1195
rect 5924 1162 6416 1178
rect 6782 1178 6798 1195
rect 7258 1195 7428 1212
rect 7486 1212 8286 1250
rect 7486 1195 7656 1212
rect 7258 1178 7274 1195
rect 6782 1162 7274 1178
rect 7640 1178 7656 1195
rect 8116 1195 8286 1212
rect 8344 1212 9144 1250
rect 8344 1195 8514 1212
rect 8116 1178 8132 1195
rect 7640 1162 8132 1178
rect 8498 1178 8514 1195
rect 8974 1195 9144 1212
rect 9202 1212 10002 1250
rect 9202 1195 9372 1212
rect 8974 1178 8990 1195
rect 8498 1162 8990 1178
rect 9356 1178 9372 1195
rect 9832 1195 10002 1212
rect 10060 1212 10860 1250
rect 10060 1195 10230 1212
rect 9832 1178 9848 1195
rect 9356 1162 9848 1178
rect 10214 1178 10230 1195
rect 10690 1195 10860 1212
rect 10690 1178 10706 1195
rect 10214 1162 10706 1178
rect 776 982 1268 998
rect 776 965 792 982
rect 622 948 792 965
rect 1252 965 1268 982
rect 1634 982 2126 998
rect 1634 965 1650 982
rect 1252 948 1422 965
rect 622 910 1422 948
rect 1480 948 1650 965
rect 2110 965 2126 982
rect 2492 982 2984 998
rect 2492 965 2508 982
rect 2110 948 2280 965
rect 1480 910 2280 948
rect 2338 948 2508 965
rect 2968 965 2984 982
rect 3350 982 3842 998
rect 3350 965 3366 982
rect 2968 948 3138 965
rect 2338 910 3138 948
rect 3196 948 3366 965
rect 3826 965 3842 982
rect 4208 982 4700 998
rect 4208 965 4224 982
rect 3826 948 3996 965
rect 3196 910 3996 948
rect 4054 948 4224 965
rect 4684 965 4700 982
rect 5066 982 5558 998
rect 5066 965 5082 982
rect 4684 948 4854 965
rect 4054 910 4854 948
rect 4912 948 5082 965
rect 5542 965 5558 982
rect 5924 982 6416 998
rect 5924 965 5940 982
rect 5542 948 5712 965
rect 4912 910 5712 948
rect 5770 948 5940 965
rect 6400 965 6416 982
rect 6782 982 7274 998
rect 6782 965 6798 982
rect 6400 948 6570 965
rect 5770 910 6570 948
rect 6628 948 6798 965
rect 7258 965 7274 982
rect 7640 982 8132 998
rect 7640 965 7656 982
rect 7258 948 7428 965
rect 6628 910 7428 948
rect 7486 948 7656 965
rect 8116 965 8132 982
rect 8498 982 8990 998
rect 8498 965 8514 982
rect 8116 948 8286 965
rect 7486 910 8286 948
rect 8344 948 8514 965
rect 8974 965 8990 982
rect 9356 982 9848 998
rect 9356 965 9372 982
rect 8974 948 9144 965
rect 8344 910 9144 948
rect 9202 948 9372 965
rect 9832 965 9848 982
rect 10214 982 10706 998
rect 10214 965 10230 982
rect 9832 948 10002 965
rect 9202 910 10002 948
rect 10060 948 10230 965
rect 10690 965 10706 982
rect 10690 948 10860 965
rect 10060 910 10860 948
rect 622 672 1422 710
rect 622 655 792 672
rect 776 638 792 655
rect 1252 655 1422 672
rect 1480 672 2280 710
rect 1480 655 1650 672
rect 1252 638 1268 655
rect 776 622 1268 638
rect 1634 638 1650 655
rect 2110 655 2280 672
rect 2338 672 3138 710
rect 2338 655 2508 672
rect 2110 638 2126 655
rect 1634 622 2126 638
rect 2492 638 2508 655
rect 2968 655 3138 672
rect 3196 672 3996 710
rect 3196 655 3366 672
rect 2968 638 2984 655
rect 2492 622 2984 638
rect 3350 638 3366 655
rect 3826 655 3996 672
rect 4054 672 4854 710
rect 4054 655 4224 672
rect 3826 638 3842 655
rect 3350 622 3842 638
rect 4208 638 4224 655
rect 4684 655 4854 672
rect 4912 672 5712 710
rect 4912 655 5082 672
rect 4684 638 4700 655
rect 4208 622 4700 638
rect 5066 638 5082 655
rect 5542 655 5712 672
rect 5770 672 6570 710
rect 5770 655 5940 672
rect 5542 638 5558 655
rect 5066 622 5558 638
rect 5924 638 5940 655
rect 6400 655 6570 672
rect 6628 672 7428 710
rect 6628 655 6798 672
rect 6400 638 6416 655
rect 5924 622 6416 638
rect 6782 638 6798 655
rect 7258 655 7428 672
rect 7486 672 8286 710
rect 7486 655 7656 672
rect 7258 638 7274 655
rect 6782 622 7274 638
rect 7640 638 7656 655
rect 8116 655 8286 672
rect 8344 672 9144 710
rect 8344 655 8514 672
rect 8116 638 8132 655
rect 7640 622 8132 638
rect 8498 638 8514 655
rect 8974 655 9144 672
rect 9202 672 10002 710
rect 9202 655 9372 672
rect 8974 638 8990 655
rect 8498 622 8990 638
rect 9356 638 9372 655
rect 9832 655 10002 672
rect 10060 672 10860 710
rect 10060 655 10230 672
rect 9832 638 9848 655
rect 9356 622 9848 638
rect 10214 638 10230 655
rect 10690 655 10860 672
rect 10690 638 10706 655
rect 10214 622 10706 638
rect 13004 2630 13136 2646
rect 13004 2613 13020 2630
rect 12970 2596 13020 2613
rect 13120 2613 13136 2630
rect 13262 2630 13394 2646
rect 13262 2613 13278 2630
rect 13120 2596 13170 2613
rect 12970 2558 13170 2596
rect 13228 2596 13278 2613
rect 13378 2613 13394 2630
rect 13520 2630 13652 2646
rect 13520 2613 13536 2630
rect 13378 2596 13428 2613
rect 13228 2558 13428 2596
rect 13486 2596 13536 2613
rect 13636 2613 13652 2630
rect 13778 2630 13910 2646
rect 13778 2613 13794 2630
rect 13636 2596 13686 2613
rect 13486 2558 13686 2596
rect 13744 2596 13794 2613
rect 13894 2613 13910 2630
rect 14036 2630 14168 2646
rect 14036 2613 14052 2630
rect 13894 2596 13944 2613
rect 13744 2558 13944 2596
rect 14002 2596 14052 2613
rect 14152 2613 14168 2630
rect 14294 2630 14426 2646
rect 14294 2613 14310 2630
rect 14152 2596 14202 2613
rect 14002 2558 14202 2596
rect 14260 2596 14310 2613
rect 14410 2613 14426 2630
rect 14552 2630 14684 2646
rect 14552 2613 14568 2630
rect 14410 2596 14460 2613
rect 14260 2558 14460 2596
rect 14518 2596 14568 2613
rect 14668 2613 14684 2630
rect 14810 2630 14942 2646
rect 14810 2613 14826 2630
rect 14668 2596 14718 2613
rect 14518 2558 14718 2596
rect 14776 2596 14826 2613
rect 14926 2613 14942 2630
rect 15068 2630 15200 2646
rect 15068 2613 15084 2630
rect 14926 2596 14976 2613
rect 14776 2558 14976 2596
rect 15034 2596 15084 2613
rect 15184 2613 15200 2630
rect 15326 2630 15458 2646
rect 15326 2613 15342 2630
rect 15184 2596 15234 2613
rect 15034 2558 15234 2596
rect 15292 2596 15342 2613
rect 15442 2613 15458 2630
rect 16300 2630 16432 2646
rect 16300 2613 16316 2630
rect 15442 2596 15492 2613
rect 15292 2558 15492 2596
rect 16266 2596 16316 2613
rect 16416 2613 16432 2630
rect 16558 2630 16690 2646
rect 16558 2613 16574 2630
rect 16416 2596 16466 2613
rect 16266 2558 16466 2596
rect 16524 2596 16574 2613
rect 16674 2613 16690 2630
rect 16816 2630 16948 2646
rect 16816 2613 16832 2630
rect 16674 2596 16724 2613
rect 16524 2558 16724 2596
rect 16782 2596 16832 2613
rect 16932 2613 16948 2630
rect 17074 2630 17206 2646
rect 17074 2613 17090 2630
rect 16932 2596 16982 2613
rect 16782 2558 16982 2596
rect 17040 2596 17090 2613
rect 17190 2613 17206 2630
rect 17332 2630 17464 2646
rect 17332 2613 17348 2630
rect 17190 2596 17240 2613
rect 17040 2558 17240 2596
rect 17298 2596 17348 2613
rect 17448 2613 17464 2630
rect 17590 2630 17722 2646
rect 17590 2613 17606 2630
rect 17448 2596 17498 2613
rect 17298 2558 17498 2596
rect 17556 2596 17606 2613
rect 17706 2613 17722 2630
rect 17848 2630 17980 2646
rect 17848 2613 17864 2630
rect 17706 2596 17756 2613
rect 17556 2558 17756 2596
rect 17814 2596 17864 2613
rect 17964 2613 17980 2630
rect 18106 2630 18238 2646
rect 18106 2613 18122 2630
rect 17964 2596 18014 2613
rect 17814 2558 18014 2596
rect 18072 2596 18122 2613
rect 18222 2613 18238 2630
rect 18364 2630 18496 2646
rect 18364 2613 18380 2630
rect 18222 2596 18272 2613
rect 18072 2558 18272 2596
rect 18330 2596 18380 2613
rect 18480 2613 18496 2630
rect 18622 2630 18754 2646
rect 18622 2613 18638 2630
rect 18480 2596 18530 2613
rect 18330 2558 18530 2596
rect 18588 2596 18638 2613
rect 18738 2613 18754 2630
rect 19596 2630 19728 2646
rect 19596 2613 19612 2630
rect 18738 2596 18788 2613
rect 18588 2558 18788 2596
rect 19562 2596 19612 2613
rect 19712 2613 19728 2630
rect 19854 2630 19986 2646
rect 19854 2613 19870 2630
rect 19712 2596 19762 2613
rect 19562 2558 19762 2596
rect 19820 2596 19870 2613
rect 19970 2613 19986 2630
rect 20112 2630 20244 2646
rect 20112 2613 20128 2630
rect 19970 2596 20020 2613
rect 19820 2558 20020 2596
rect 20078 2596 20128 2613
rect 20228 2613 20244 2630
rect 20370 2630 20502 2646
rect 20370 2613 20386 2630
rect 20228 2596 20278 2613
rect 20078 2558 20278 2596
rect 20336 2596 20386 2613
rect 20486 2613 20502 2630
rect 20628 2630 20760 2646
rect 20628 2613 20644 2630
rect 20486 2596 20536 2613
rect 20336 2558 20536 2596
rect 20594 2596 20644 2613
rect 20744 2613 20760 2630
rect 20886 2630 21018 2646
rect 20886 2613 20902 2630
rect 20744 2596 20794 2613
rect 20594 2558 20794 2596
rect 20852 2596 20902 2613
rect 21002 2613 21018 2630
rect 21144 2630 21276 2646
rect 21144 2613 21160 2630
rect 21002 2596 21052 2613
rect 20852 2558 21052 2596
rect 21110 2596 21160 2613
rect 21260 2613 21276 2630
rect 21402 2630 21534 2646
rect 21402 2613 21418 2630
rect 21260 2596 21310 2613
rect 21110 2558 21310 2596
rect 21368 2596 21418 2613
rect 21518 2613 21534 2630
rect 21660 2630 21792 2646
rect 21660 2613 21676 2630
rect 21518 2596 21568 2613
rect 21368 2558 21568 2596
rect 21626 2596 21676 2613
rect 21776 2613 21792 2630
rect 21918 2630 22050 2646
rect 21918 2613 21934 2630
rect 21776 2596 21826 2613
rect 21626 2558 21826 2596
rect 21884 2596 21934 2613
rect 22034 2613 22050 2630
rect 22034 2596 22084 2613
rect 21884 2558 22084 2596
rect 12970 2120 13170 2158
rect 12970 2103 13020 2120
rect 13004 2086 13020 2103
rect 13120 2103 13170 2120
rect 13228 2120 13428 2158
rect 13228 2103 13278 2120
rect 13120 2086 13136 2103
rect 13004 2070 13136 2086
rect 13262 2086 13278 2103
rect 13378 2103 13428 2120
rect 13486 2120 13686 2158
rect 13486 2103 13536 2120
rect 13378 2086 13394 2103
rect 13262 2070 13394 2086
rect 13520 2086 13536 2103
rect 13636 2103 13686 2120
rect 13744 2120 13944 2158
rect 13744 2103 13794 2120
rect 13636 2086 13652 2103
rect 13520 2070 13652 2086
rect 13778 2086 13794 2103
rect 13894 2103 13944 2120
rect 14002 2120 14202 2158
rect 14002 2103 14052 2120
rect 13894 2086 13910 2103
rect 13778 2070 13910 2086
rect 14036 2086 14052 2103
rect 14152 2103 14202 2120
rect 14260 2120 14460 2158
rect 14260 2103 14310 2120
rect 14152 2086 14168 2103
rect 14036 2070 14168 2086
rect 14294 2086 14310 2103
rect 14410 2103 14460 2120
rect 14518 2120 14718 2158
rect 14518 2103 14568 2120
rect 14410 2086 14426 2103
rect 14294 2070 14426 2086
rect 14552 2086 14568 2103
rect 14668 2103 14718 2120
rect 14776 2120 14976 2158
rect 14776 2103 14826 2120
rect 14668 2086 14684 2103
rect 14552 2070 14684 2086
rect 14810 2086 14826 2103
rect 14926 2103 14976 2120
rect 15034 2120 15234 2158
rect 15034 2103 15084 2120
rect 14926 2086 14942 2103
rect 14810 2070 14942 2086
rect 15068 2086 15084 2103
rect 15184 2103 15234 2120
rect 15292 2120 15492 2158
rect 15292 2103 15342 2120
rect 15184 2086 15200 2103
rect 15068 2070 15200 2086
rect 15326 2086 15342 2103
rect 15442 2103 15492 2120
rect 16266 2120 16466 2158
rect 16266 2103 16316 2120
rect 15442 2086 15458 2103
rect 15326 2070 15458 2086
rect 16300 2086 16316 2103
rect 16416 2103 16466 2120
rect 16524 2120 16724 2158
rect 16524 2103 16574 2120
rect 16416 2086 16432 2103
rect 16300 2070 16432 2086
rect 16558 2086 16574 2103
rect 16674 2103 16724 2120
rect 16782 2120 16982 2158
rect 16782 2103 16832 2120
rect 16674 2086 16690 2103
rect 16558 2070 16690 2086
rect 16816 2086 16832 2103
rect 16932 2103 16982 2120
rect 17040 2120 17240 2158
rect 17040 2103 17090 2120
rect 16932 2086 16948 2103
rect 16816 2070 16948 2086
rect 17074 2086 17090 2103
rect 17190 2103 17240 2120
rect 17298 2120 17498 2158
rect 17298 2103 17348 2120
rect 17190 2086 17206 2103
rect 17074 2070 17206 2086
rect 17332 2086 17348 2103
rect 17448 2103 17498 2120
rect 17556 2120 17756 2158
rect 17556 2103 17606 2120
rect 17448 2086 17464 2103
rect 17332 2070 17464 2086
rect 17590 2086 17606 2103
rect 17706 2103 17756 2120
rect 17814 2120 18014 2158
rect 17814 2103 17864 2120
rect 17706 2086 17722 2103
rect 17590 2070 17722 2086
rect 17848 2086 17864 2103
rect 17964 2103 18014 2120
rect 18072 2120 18272 2158
rect 18072 2103 18122 2120
rect 17964 2086 17980 2103
rect 17848 2070 17980 2086
rect 18106 2086 18122 2103
rect 18222 2103 18272 2120
rect 18330 2120 18530 2158
rect 18330 2103 18380 2120
rect 18222 2086 18238 2103
rect 18106 2070 18238 2086
rect 18364 2086 18380 2103
rect 18480 2103 18530 2120
rect 18588 2120 18788 2158
rect 18588 2103 18638 2120
rect 18480 2086 18496 2103
rect 18364 2070 18496 2086
rect 18622 2086 18638 2103
rect 18738 2103 18788 2120
rect 19562 2120 19762 2158
rect 19562 2103 19612 2120
rect 18738 2086 18754 2103
rect 18622 2070 18754 2086
rect 19596 2086 19612 2103
rect 19712 2103 19762 2120
rect 19820 2120 20020 2158
rect 19820 2103 19870 2120
rect 19712 2086 19728 2103
rect 19596 2070 19728 2086
rect 19854 2086 19870 2103
rect 19970 2103 20020 2120
rect 20078 2120 20278 2158
rect 20078 2103 20128 2120
rect 19970 2086 19986 2103
rect 19854 2070 19986 2086
rect 20112 2086 20128 2103
rect 20228 2103 20278 2120
rect 20336 2120 20536 2158
rect 20336 2103 20386 2120
rect 20228 2086 20244 2103
rect 20112 2070 20244 2086
rect 20370 2086 20386 2103
rect 20486 2103 20536 2120
rect 20594 2120 20794 2158
rect 20594 2103 20644 2120
rect 20486 2086 20502 2103
rect 20370 2070 20502 2086
rect 20628 2086 20644 2103
rect 20744 2103 20794 2120
rect 20852 2120 21052 2158
rect 20852 2103 20902 2120
rect 20744 2086 20760 2103
rect 20628 2070 20760 2086
rect 20886 2086 20902 2103
rect 21002 2103 21052 2120
rect 21110 2120 21310 2158
rect 21110 2103 21160 2120
rect 21002 2086 21018 2103
rect 20886 2070 21018 2086
rect 21144 2086 21160 2103
rect 21260 2103 21310 2120
rect 21368 2120 21568 2158
rect 21368 2103 21418 2120
rect 21260 2086 21276 2103
rect 21144 2070 21276 2086
rect 21402 2086 21418 2103
rect 21518 2103 21568 2120
rect 21626 2120 21826 2158
rect 21626 2103 21676 2120
rect 21518 2086 21534 2103
rect 21402 2070 21534 2086
rect 21660 2086 21676 2103
rect 21776 2103 21826 2120
rect 21884 2120 22084 2158
rect 21884 2103 21934 2120
rect 21776 2086 21792 2103
rect 21660 2070 21792 2086
rect 21918 2086 21934 2103
rect 22034 2103 22084 2120
rect 22034 2086 22050 2103
rect 21918 2070 22050 2086
rect 12576 1522 13068 1538
rect 12576 1505 12592 1522
rect 12422 1488 12592 1505
rect 13052 1505 13068 1522
rect 13434 1522 13926 1538
rect 13434 1505 13450 1522
rect 13052 1488 13222 1505
rect 12422 1450 13222 1488
rect 13280 1488 13450 1505
rect 13910 1505 13926 1522
rect 14292 1522 14784 1538
rect 14292 1505 14308 1522
rect 13910 1488 14080 1505
rect 13280 1450 14080 1488
rect 14138 1488 14308 1505
rect 14768 1505 14784 1522
rect 15150 1522 15642 1538
rect 15150 1505 15166 1522
rect 14768 1488 14938 1505
rect 14138 1450 14938 1488
rect 14996 1488 15166 1505
rect 15626 1505 15642 1522
rect 16008 1522 16500 1538
rect 16008 1505 16024 1522
rect 15626 1488 15796 1505
rect 14996 1450 15796 1488
rect 15854 1488 16024 1505
rect 16484 1505 16500 1522
rect 16866 1522 17358 1538
rect 16866 1505 16882 1522
rect 16484 1488 16654 1505
rect 15854 1450 16654 1488
rect 16712 1488 16882 1505
rect 17342 1505 17358 1522
rect 17724 1522 18216 1538
rect 17724 1505 17740 1522
rect 17342 1488 17512 1505
rect 16712 1450 17512 1488
rect 17570 1488 17740 1505
rect 18200 1505 18216 1522
rect 18582 1522 19074 1538
rect 18582 1505 18598 1522
rect 18200 1488 18370 1505
rect 17570 1450 18370 1488
rect 18428 1488 18598 1505
rect 19058 1505 19074 1522
rect 19440 1522 19932 1538
rect 19440 1505 19456 1522
rect 19058 1488 19228 1505
rect 18428 1450 19228 1488
rect 19286 1488 19456 1505
rect 19916 1505 19932 1522
rect 20298 1522 20790 1538
rect 20298 1505 20314 1522
rect 19916 1488 20086 1505
rect 19286 1450 20086 1488
rect 20144 1488 20314 1505
rect 20774 1505 20790 1522
rect 21156 1522 21648 1538
rect 21156 1505 21172 1522
rect 20774 1488 20944 1505
rect 20144 1450 20944 1488
rect 21002 1488 21172 1505
rect 21632 1505 21648 1522
rect 22014 1522 22506 1538
rect 22014 1505 22030 1522
rect 21632 1488 21802 1505
rect 21002 1450 21802 1488
rect 21860 1488 22030 1505
rect 22490 1505 22506 1522
rect 22490 1488 22660 1505
rect 21860 1450 22660 1488
rect 12422 1212 13222 1250
rect 12422 1195 12592 1212
rect 12576 1178 12592 1195
rect 13052 1195 13222 1212
rect 13280 1212 14080 1250
rect 13280 1195 13450 1212
rect 13052 1178 13068 1195
rect 12576 1162 13068 1178
rect 13434 1178 13450 1195
rect 13910 1195 14080 1212
rect 14138 1212 14938 1250
rect 14138 1195 14308 1212
rect 13910 1178 13926 1195
rect 13434 1162 13926 1178
rect 14292 1178 14308 1195
rect 14768 1195 14938 1212
rect 14996 1212 15796 1250
rect 14996 1195 15166 1212
rect 14768 1178 14784 1195
rect 14292 1162 14784 1178
rect 15150 1178 15166 1195
rect 15626 1195 15796 1212
rect 15854 1212 16654 1250
rect 15854 1195 16024 1212
rect 15626 1178 15642 1195
rect 15150 1162 15642 1178
rect 16008 1178 16024 1195
rect 16484 1195 16654 1212
rect 16712 1212 17512 1250
rect 16712 1195 16882 1212
rect 16484 1178 16500 1195
rect 16008 1162 16500 1178
rect 16866 1178 16882 1195
rect 17342 1195 17512 1212
rect 17570 1212 18370 1250
rect 17570 1195 17740 1212
rect 17342 1178 17358 1195
rect 16866 1162 17358 1178
rect 17724 1178 17740 1195
rect 18200 1195 18370 1212
rect 18428 1212 19228 1250
rect 18428 1195 18598 1212
rect 18200 1178 18216 1195
rect 17724 1162 18216 1178
rect 18582 1178 18598 1195
rect 19058 1195 19228 1212
rect 19286 1212 20086 1250
rect 19286 1195 19456 1212
rect 19058 1178 19074 1195
rect 18582 1162 19074 1178
rect 19440 1178 19456 1195
rect 19916 1195 20086 1212
rect 20144 1212 20944 1250
rect 20144 1195 20314 1212
rect 19916 1178 19932 1195
rect 19440 1162 19932 1178
rect 20298 1178 20314 1195
rect 20774 1195 20944 1212
rect 21002 1212 21802 1250
rect 21002 1195 21172 1212
rect 20774 1178 20790 1195
rect 20298 1162 20790 1178
rect 21156 1178 21172 1195
rect 21632 1195 21802 1212
rect 21860 1212 22660 1250
rect 21860 1195 22030 1212
rect 21632 1178 21648 1195
rect 21156 1162 21648 1178
rect 22014 1178 22030 1195
rect 22490 1195 22660 1212
rect 22490 1178 22506 1195
rect 22014 1162 22506 1178
rect 12576 982 13068 998
rect 12576 965 12592 982
rect 12422 948 12592 965
rect 13052 965 13068 982
rect 13434 982 13926 998
rect 13434 965 13450 982
rect 13052 948 13222 965
rect 12422 910 13222 948
rect 13280 948 13450 965
rect 13910 965 13926 982
rect 14292 982 14784 998
rect 14292 965 14308 982
rect 13910 948 14080 965
rect 13280 910 14080 948
rect 14138 948 14308 965
rect 14768 965 14784 982
rect 15150 982 15642 998
rect 15150 965 15166 982
rect 14768 948 14938 965
rect 14138 910 14938 948
rect 14996 948 15166 965
rect 15626 965 15642 982
rect 16008 982 16500 998
rect 16008 965 16024 982
rect 15626 948 15796 965
rect 14996 910 15796 948
rect 15854 948 16024 965
rect 16484 965 16500 982
rect 16866 982 17358 998
rect 16866 965 16882 982
rect 16484 948 16654 965
rect 15854 910 16654 948
rect 16712 948 16882 965
rect 17342 965 17358 982
rect 17724 982 18216 998
rect 17724 965 17740 982
rect 17342 948 17512 965
rect 16712 910 17512 948
rect 17570 948 17740 965
rect 18200 965 18216 982
rect 18582 982 19074 998
rect 18582 965 18598 982
rect 18200 948 18370 965
rect 17570 910 18370 948
rect 18428 948 18598 965
rect 19058 965 19074 982
rect 19440 982 19932 998
rect 19440 965 19456 982
rect 19058 948 19228 965
rect 18428 910 19228 948
rect 19286 948 19456 965
rect 19916 965 19932 982
rect 20298 982 20790 998
rect 20298 965 20314 982
rect 19916 948 20086 965
rect 19286 910 20086 948
rect 20144 948 20314 965
rect 20774 965 20790 982
rect 21156 982 21648 998
rect 21156 965 21172 982
rect 20774 948 20944 965
rect 20144 910 20944 948
rect 21002 948 21172 965
rect 21632 965 21648 982
rect 22014 982 22506 998
rect 22014 965 22030 982
rect 21632 948 21802 965
rect 21002 910 21802 948
rect 21860 948 22030 965
rect 22490 965 22506 982
rect 22490 948 22660 965
rect 21860 910 22660 948
rect 12422 672 13222 710
rect 12422 655 12592 672
rect 12576 638 12592 655
rect 13052 655 13222 672
rect 13280 672 14080 710
rect 13280 655 13450 672
rect 13052 638 13068 655
rect 12576 622 13068 638
rect 13434 638 13450 655
rect 13910 655 14080 672
rect 14138 672 14938 710
rect 14138 655 14308 672
rect 13910 638 13926 655
rect 13434 622 13926 638
rect 14292 638 14308 655
rect 14768 655 14938 672
rect 14996 672 15796 710
rect 14996 655 15166 672
rect 14768 638 14784 655
rect 14292 622 14784 638
rect 15150 638 15166 655
rect 15626 655 15796 672
rect 15854 672 16654 710
rect 15854 655 16024 672
rect 15626 638 15642 655
rect 15150 622 15642 638
rect 16008 638 16024 655
rect 16484 655 16654 672
rect 16712 672 17512 710
rect 16712 655 16882 672
rect 16484 638 16500 655
rect 16008 622 16500 638
rect 16866 638 16882 655
rect 17342 655 17512 672
rect 17570 672 18370 710
rect 17570 655 17740 672
rect 17342 638 17358 655
rect 16866 622 17358 638
rect 17724 638 17740 655
rect 18200 655 18370 672
rect 18428 672 19228 710
rect 18428 655 18598 672
rect 18200 638 18216 655
rect 17724 622 18216 638
rect 18582 638 18598 655
rect 19058 655 19228 672
rect 19286 672 20086 710
rect 19286 655 19456 672
rect 19058 638 19074 655
rect 18582 622 19074 638
rect 19440 638 19456 655
rect 19916 655 20086 672
rect 20144 672 20944 710
rect 20144 655 20314 672
rect 19916 638 19932 655
rect 19440 622 19932 638
rect 20298 638 20314 655
rect 20774 655 20944 672
rect 21002 672 21802 710
rect 21002 655 21172 672
rect 20774 638 20790 655
rect 20298 622 20790 638
rect 21156 638 21172 655
rect 21632 655 21802 672
rect 21860 672 22660 710
rect 21860 655 22030 672
rect 21632 638 21648 655
rect 21156 622 21648 638
rect 22014 638 22030 655
rect 22490 655 22660 672
rect 22490 638 22506 655
rect 22014 622 22506 638
rect 776 -1442 1268 -1426
rect 776 -1459 792 -1442
rect 622 -1476 792 -1459
rect 1252 -1459 1268 -1442
rect 1634 -1442 2126 -1426
rect 1634 -1459 1650 -1442
rect 1252 -1476 1422 -1459
rect 622 -1514 1422 -1476
rect 1480 -1476 1650 -1459
rect 2110 -1459 2126 -1442
rect 2492 -1442 2984 -1426
rect 2492 -1459 2508 -1442
rect 2110 -1476 2280 -1459
rect 1480 -1514 2280 -1476
rect 2338 -1476 2508 -1459
rect 2968 -1459 2984 -1442
rect 3350 -1442 3842 -1426
rect 3350 -1459 3366 -1442
rect 2968 -1476 3138 -1459
rect 2338 -1514 3138 -1476
rect 3196 -1476 3366 -1459
rect 3826 -1459 3842 -1442
rect 4208 -1442 4700 -1426
rect 4208 -1459 4224 -1442
rect 3826 -1476 3996 -1459
rect 3196 -1514 3996 -1476
rect 4054 -1476 4224 -1459
rect 4684 -1459 4700 -1442
rect 5066 -1442 5558 -1426
rect 5066 -1459 5082 -1442
rect 4684 -1476 4854 -1459
rect 4054 -1514 4854 -1476
rect 4912 -1476 5082 -1459
rect 5542 -1459 5558 -1442
rect 5924 -1442 6416 -1426
rect 5924 -1459 5940 -1442
rect 5542 -1476 5712 -1459
rect 4912 -1514 5712 -1476
rect 5770 -1476 5940 -1459
rect 6400 -1459 6416 -1442
rect 6782 -1442 7274 -1426
rect 6782 -1459 6798 -1442
rect 6400 -1476 6570 -1459
rect 5770 -1514 6570 -1476
rect 6628 -1476 6798 -1459
rect 7258 -1459 7274 -1442
rect 7640 -1442 8132 -1426
rect 7640 -1459 7656 -1442
rect 7258 -1476 7428 -1459
rect 6628 -1514 7428 -1476
rect 7486 -1476 7656 -1459
rect 8116 -1459 8132 -1442
rect 8498 -1442 8990 -1426
rect 8498 -1459 8514 -1442
rect 8116 -1476 8286 -1459
rect 7486 -1514 8286 -1476
rect 8344 -1476 8514 -1459
rect 8974 -1459 8990 -1442
rect 9356 -1442 9848 -1426
rect 9356 -1459 9372 -1442
rect 8974 -1476 9144 -1459
rect 8344 -1514 9144 -1476
rect 9202 -1476 9372 -1459
rect 9832 -1459 9848 -1442
rect 10214 -1442 10706 -1426
rect 10214 -1459 10230 -1442
rect 9832 -1476 10002 -1459
rect 9202 -1514 10002 -1476
rect 10060 -1476 10230 -1459
rect 10690 -1459 10706 -1442
rect 10690 -1476 10860 -1459
rect 10060 -1514 10860 -1476
rect 622 -1752 1422 -1714
rect 622 -1769 792 -1752
rect 776 -1786 792 -1769
rect 1252 -1769 1422 -1752
rect 1480 -1752 2280 -1714
rect 1480 -1769 1650 -1752
rect 1252 -1786 1268 -1769
rect 776 -1802 1268 -1786
rect 1634 -1786 1650 -1769
rect 2110 -1769 2280 -1752
rect 2338 -1752 3138 -1714
rect 2338 -1769 2508 -1752
rect 2110 -1786 2126 -1769
rect 1634 -1802 2126 -1786
rect 2492 -1786 2508 -1769
rect 2968 -1769 3138 -1752
rect 3196 -1752 3996 -1714
rect 3196 -1769 3366 -1752
rect 2968 -1786 2984 -1769
rect 2492 -1802 2984 -1786
rect 3350 -1786 3366 -1769
rect 3826 -1769 3996 -1752
rect 4054 -1752 4854 -1714
rect 4054 -1769 4224 -1752
rect 3826 -1786 3842 -1769
rect 3350 -1802 3842 -1786
rect 4208 -1786 4224 -1769
rect 4684 -1769 4854 -1752
rect 4912 -1752 5712 -1714
rect 4912 -1769 5082 -1752
rect 4684 -1786 4700 -1769
rect 4208 -1802 4700 -1786
rect 5066 -1786 5082 -1769
rect 5542 -1769 5712 -1752
rect 5770 -1752 6570 -1714
rect 5770 -1769 5940 -1752
rect 5542 -1786 5558 -1769
rect 5066 -1802 5558 -1786
rect 5924 -1786 5940 -1769
rect 6400 -1769 6570 -1752
rect 6628 -1752 7428 -1714
rect 6628 -1769 6798 -1752
rect 6400 -1786 6416 -1769
rect 5924 -1802 6416 -1786
rect 6782 -1786 6798 -1769
rect 7258 -1769 7428 -1752
rect 7486 -1752 8286 -1714
rect 7486 -1769 7656 -1752
rect 7258 -1786 7274 -1769
rect 6782 -1802 7274 -1786
rect 7640 -1786 7656 -1769
rect 8116 -1769 8286 -1752
rect 8344 -1752 9144 -1714
rect 8344 -1769 8514 -1752
rect 8116 -1786 8132 -1769
rect 7640 -1802 8132 -1786
rect 8498 -1786 8514 -1769
rect 8974 -1769 9144 -1752
rect 9202 -1752 10002 -1714
rect 9202 -1769 9372 -1752
rect 8974 -1786 8990 -1769
rect 8498 -1802 8990 -1786
rect 9356 -1786 9372 -1769
rect 9832 -1769 10002 -1752
rect 10060 -1752 10860 -1714
rect 10060 -1769 10230 -1752
rect 9832 -1786 9848 -1769
rect 9356 -1802 9848 -1786
rect 10214 -1786 10230 -1769
rect 10690 -1769 10860 -1752
rect 10690 -1786 10706 -1769
rect 10214 -1802 10706 -1786
rect 776 -1982 1268 -1966
rect 776 -1999 792 -1982
rect 622 -2016 792 -1999
rect 1252 -1999 1268 -1982
rect 1634 -1982 2126 -1966
rect 1634 -1999 1650 -1982
rect 1252 -2016 1422 -1999
rect 622 -2054 1422 -2016
rect 1480 -2016 1650 -1999
rect 2110 -1999 2126 -1982
rect 2492 -1982 2984 -1966
rect 2492 -1999 2508 -1982
rect 2110 -2016 2280 -1999
rect 1480 -2054 2280 -2016
rect 2338 -2016 2508 -1999
rect 2968 -1999 2984 -1982
rect 3350 -1982 3842 -1966
rect 3350 -1999 3366 -1982
rect 2968 -2016 3138 -1999
rect 2338 -2054 3138 -2016
rect 3196 -2016 3366 -1999
rect 3826 -1999 3842 -1982
rect 4208 -1982 4700 -1966
rect 4208 -1999 4224 -1982
rect 3826 -2016 3996 -1999
rect 3196 -2054 3996 -2016
rect 4054 -2016 4224 -1999
rect 4684 -1999 4700 -1982
rect 5066 -1982 5558 -1966
rect 5066 -1999 5082 -1982
rect 4684 -2016 4854 -1999
rect 4054 -2054 4854 -2016
rect 4912 -2016 5082 -1999
rect 5542 -1999 5558 -1982
rect 5924 -1982 6416 -1966
rect 5924 -1999 5940 -1982
rect 5542 -2016 5712 -1999
rect 4912 -2054 5712 -2016
rect 5770 -2016 5940 -1999
rect 6400 -1999 6416 -1982
rect 6782 -1982 7274 -1966
rect 6782 -1999 6798 -1982
rect 6400 -2016 6570 -1999
rect 5770 -2054 6570 -2016
rect 6628 -2016 6798 -1999
rect 7258 -1999 7274 -1982
rect 7640 -1982 8132 -1966
rect 7640 -1999 7656 -1982
rect 7258 -2016 7428 -1999
rect 6628 -2054 7428 -2016
rect 7486 -2016 7656 -1999
rect 8116 -1999 8132 -1982
rect 8498 -1982 8990 -1966
rect 8498 -1999 8514 -1982
rect 8116 -2016 8286 -1999
rect 7486 -2054 8286 -2016
rect 8344 -2016 8514 -1999
rect 8974 -1999 8990 -1982
rect 9356 -1982 9848 -1966
rect 9356 -1999 9372 -1982
rect 8974 -2016 9144 -1999
rect 8344 -2054 9144 -2016
rect 9202 -2016 9372 -1999
rect 9832 -1999 9848 -1982
rect 10214 -1982 10706 -1966
rect 10214 -1999 10230 -1982
rect 9832 -2016 10002 -1999
rect 9202 -2054 10002 -2016
rect 10060 -2016 10230 -1999
rect 10690 -1999 10706 -1982
rect 10690 -2016 10860 -1999
rect 10060 -2054 10860 -2016
rect 622 -2292 1422 -2254
rect 622 -2309 792 -2292
rect 776 -2326 792 -2309
rect 1252 -2309 1422 -2292
rect 1480 -2292 2280 -2254
rect 1480 -2309 1650 -2292
rect 1252 -2326 1268 -2309
rect 776 -2342 1268 -2326
rect 1634 -2326 1650 -2309
rect 2110 -2309 2280 -2292
rect 2338 -2292 3138 -2254
rect 2338 -2309 2508 -2292
rect 2110 -2326 2126 -2309
rect 1634 -2342 2126 -2326
rect 2492 -2326 2508 -2309
rect 2968 -2309 3138 -2292
rect 3196 -2292 3996 -2254
rect 3196 -2309 3366 -2292
rect 2968 -2326 2984 -2309
rect 2492 -2342 2984 -2326
rect 3350 -2326 3366 -2309
rect 3826 -2309 3996 -2292
rect 4054 -2292 4854 -2254
rect 4054 -2309 4224 -2292
rect 3826 -2326 3842 -2309
rect 3350 -2342 3842 -2326
rect 4208 -2326 4224 -2309
rect 4684 -2309 4854 -2292
rect 4912 -2292 5712 -2254
rect 4912 -2309 5082 -2292
rect 4684 -2326 4700 -2309
rect 4208 -2342 4700 -2326
rect 5066 -2326 5082 -2309
rect 5542 -2309 5712 -2292
rect 5770 -2292 6570 -2254
rect 5770 -2309 5940 -2292
rect 5542 -2326 5558 -2309
rect 5066 -2342 5558 -2326
rect 5924 -2326 5940 -2309
rect 6400 -2309 6570 -2292
rect 6628 -2292 7428 -2254
rect 6628 -2309 6798 -2292
rect 6400 -2326 6416 -2309
rect 5924 -2342 6416 -2326
rect 6782 -2326 6798 -2309
rect 7258 -2309 7428 -2292
rect 7486 -2292 8286 -2254
rect 7486 -2309 7656 -2292
rect 7258 -2326 7274 -2309
rect 6782 -2342 7274 -2326
rect 7640 -2326 7656 -2309
rect 8116 -2309 8286 -2292
rect 8344 -2292 9144 -2254
rect 8344 -2309 8514 -2292
rect 8116 -2326 8132 -2309
rect 7640 -2342 8132 -2326
rect 8498 -2326 8514 -2309
rect 8974 -2309 9144 -2292
rect 9202 -2292 10002 -2254
rect 9202 -2309 9372 -2292
rect 8974 -2326 8990 -2309
rect 8498 -2342 8990 -2326
rect 9356 -2326 9372 -2309
rect 9832 -2309 10002 -2292
rect 10060 -2292 10860 -2254
rect 10060 -2309 10230 -2292
rect 9832 -2326 9848 -2309
rect 9356 -2342 9848 -2326
rect 10214 -2326 10230 -2309
rect 10690 -2309 10860 -2292
rect 10690 -2326 10706 -2309
rect 10214 -2342 10706 -2326
rect 1204 -2890 1336 -2874
rect 1204 -2907 1220 -2890
rect 1170 -2924 1220 -2907
rect 1320 -2907 1336 -2890
rect 1462 -2890 1594 -2874
rect 1462 -2907 1478 -2890
rect 1320 -2924 1370 -2907
rect 1170 -2962 1370 -2924
rect 1428 -2924 1478 -2907
rect 1578 -2907 1594 -2890
rect 1720 -2890 1852 -2874
rect 1720 -2907 1736 -2890
rect 1578 -2924 1628 -2907
rect 1428 -2962 1628 -2924
rect 1686 -2924 1736 -2907
rect 1836 -2907 1852 -2890
rect 1978 -2890 2110 -2874
rect 1978 -2907 1994 -2890
rect 1836 -2924 1886 -2907
rect 1686 -2962 1886 -2924
rect 1944 -2924 1994 -2907
rect 2094 -2907 2110 -2890
rect 2236 -2890 2368 -2874
rect 2236 -2907 2252 -2890
rect 2094 -2924 2144 -2907
rect 1944 -2962 2144 -2924
rect 2202 -2924 2252 -2907
rect 2352 -2907 2368 -2890
rect 2494 -2890 2626 -2874
rect 2494 -2907 2510 -2890
rect 2352 -2924 2402 -2907
rect 2202 -2962 2402 -2924
rect 2460 -2924 2510 -2907
rect 2610 -2907 2626 -2890
rect 2752 -2890 2884 -2874
rect 2752 -2907 2768 -2890
rect 2610 -2924 2660 -2907
rect 2460 -2962 2660 -2924
rect 2718 -2924 2768 -2907
rect 2868 -2907 2884 -2890
rect 3010 -2890 3142 -2874
rect 3010 -2907 3026 -2890
rect 2868 -2924 2918 -2907
rect 2718 -2962 2918 -2924
rect 2976 -2924 3026 -2907
rect 3126 -2907 3142 -2890
rect 3268 -2890 3400 -2874
rect 3268 -2907 3284 -2890
rect 3126 -2924 3176 -2907
rect 2976 -2962 3176 -2924
rect 3234 -2924 3284 -2907
rect 3384 -2907 3400 -2890
rect 3526 -2890 3658 -2874
rect 3526 -2907 3542 -2890
rect 3384 -2924 3434 -2907
rect 3234 -2962 3434 -2924
rect 3492 -2924 3542 -2907
rect 3642 -2907 3658 -2890
rect 4500 -2890 4632 -2874
rect 4500 -2907 4516 -2890
rect 3642 -2924 3692 -2907
rect 3492 -2962 3692 -2924
rect 4466 -2924 4516 -2907
rect 4616 -2907 4632 -2890
rect 4758 -2890 4890 -2874
rect 4758 -2907 4774 -2890
rect 4616 -2924 4666 -2907
rect 4466 -2962 4666 -2924
rect 4724 -2924 4774 -2907
rect 4874 -2907 4890 -2890
rect 5016 -2890 5148 -2874
rect 5016 -2907 5032 -2890
rect 4874 -2924 4924 -2907
rect 4724 -2962 4924 -2924
rect 4982 -2924 5032 -2907
rect 5132 -2907 5148 -2890
rect 5274 -2890 5406 -2874
rect 5274 -2907 5290 -2890
rect 5132 -2924 5182 -2907
rect 4982 -2962 5182 -2924
rect 5240 -2924 5290 -2907
rect 5390 -2907 5406 -2890
rect 5532 -2890 5664 -2874
rect 5532 -2907 5548 -2890
rect 5390 -2924 5440 -2907
rect 5240 -2962 5440 -2924
rect 5498 -2924 5548 -2907
rect 5648 -2907 5664 -2890
rect 5790 -2890 5922 -2874
rect 5790 -2907 5806 -2890
rect 5648 -2924 5698 -2907
rect 5498 -2962 5698 -2924
rect 5756 -2924 5806 -2907
rect 5906 -2907 5922 -2890
rect 6048 -2890 6180 -2874
rect 6048 -2907 6064 -2890
rect 5906 -2924 5956 -2907
rect 5756 -2962 5956 -2924
rect 6014 -2924 6064 -2907
rect 6164 -2907 6180 -2890
rect 6306 -2890 6438 -2874
rect 6306 -2907 6322 -2890
rect 6164 -2924 6214 -2907
rect 6014 -2962 6214 -2924
rect 6272 -2924 6322 -2907
rect 6422 -2907 6438 -2890
rect 6564 -2890 6696 -2874
rect 6564 -2907 6580 -2890
rect 6422 -2924 6472 -2907
rect 6272 -2962 6472 -2924
rect 6530 -2924 6580 -2907
rect 6680 -2907 6696 -2890
rect 6822 -2890 6954 -2874
rect 6822 -2907 6838 -2890
rect 6680 -2924 6730 -2907
rect 6530 -2962 6730 -2924
rect 6788 -2924 6838 -2907
rect 6938 -2907 6954 -2890
rect 7796 -2890 7928 -2874
rect 7796 -2907 7812 -2890
rect 6938 -2924 6988 -2907
rect 6788 -2962 6988 -2924
rect 7762 -2924 7812 -2907
rect 7912 -2907 7928 -2890
rect 8054 -2890 8186 -2874
rect 8054 -2907 8070 -2890
rect 7912 -2924 7962 -2907
rect 7762 -2962 7962 -2924
rect 8020 -2924 8070 -2907
rect 8170 -2907 8186 -2890
rect 8312 -2890 8444 -2874
rect 8312 -2907 8328 -2890
rect 8170 -2924 8220 -2907
rect 8020 -2962 8220 -2924
rect 8278 -2924 8328 -2907
rect 8428 -2907 8444 -2890
rect 8570 -2890 8702 -2874
rect 8570 -2907 8586 -2890
rect 8428 -2924 8478 -2907
rect 8278 -2962 8478 -2924
rect 8536 -2924 8586 -2907
rect 8686 -2907 8702 -2890
rect 8828 -2890 8960 -2874
rect 8828 -2907 8844 -2890
rect 8686 -2924 8736 -2907
rect 8536 -2962 8736 -2924
rect 8794 -2924 8844 -2907
rect 8944 -2907 8960 -2890
rect 9086 -2890 9218 -2874
rect 9086 -2907 9102 -2890
rect 8944 -2924 8994 -2907
rect 8794 -2962 8994 -2924
rect 9052 -2924 9102 -2907
rect 9202 -2907 9218 -2890
rect 9344 -2890 9476 -2874
rect 9344 -2907 9360 -2890
rect 9202 -2924 9252 -2907
rect 9052 -2962 9252 -2924
rect 9310 -2924 9360 -2907
rect 9460 -2907 9476 -2890
rect 9602 -2890 9734 -2874
rect 9602 -2907 9618 -2890
rect 9460 -2924 9510 -2907
rect 9310 -2962 9510 -2924
rect 9568 -2924 9618 -2907
rect 9718 -2907 9734 -2890
rect 9860 -2890 9992 -2874
rect 9860 -2907 9876 -2890
rect 9718 -2924 9768 -2907
rect 9568 -2962 9768 -2924
rect 9826 -2924 9876 -2907
rect 9976 -2907 9992 -2890
rect 10118 -2890 10250 -2874
rect 10118 -2907 10134 -2890
rect 9976 -2924 10026 -2907
rect 9826 -2962 10026 -2924
rect 10084 -2924 10134 -2907
rect 10234 -2907 10250 -2890
rect 10234 -2924 10284 -2907
rect 10084 -2962 10284 -2924
rect 1170 -3400 1370 -3362
rect 1170 -3417 1220 -3400
rect 1204 -3434 1220 -3417
rect 1320 -3417 1370 -3400
rect 1428 -3400 1628 -3362
rect 1428 -3417 1478 -3400
rect 1320 -3434 1336 -3417
rect 1204 -3450 1336 -3434
rect 1462 -3434 1478 -3417
rect 1578 -3417 1628 -3400
rect 1686 -3400 1886 -3362
rect 1686 -3417 1736 -3400
rect 1578 -3434 1594 -3417
rect 1462 -3450 1594 -3434
rect 1720 -3434 1736 -3417
rect 1836 -3417 1886 -3400
rect 1944 -3400 2144 -3362
rect 1944 -3417 1994 -3400
rect 1836 -3434 1852 -3417
rect 1720 -3450 1852 -3434
rect 1978 -3434 1994 -3417
rect 2094 -3417 2144 -3400
rect 2202 -3400 2402 -3362
rect 2202 -3417 2252 -3400
rect 2094 -3434 2110 -3417
rect 1978 -3450 2110 -3434
rect 2236 -3434 2252 -3417
rect 2352 -3417 2402 -3400
rect 2460 -3400 2660 -3362
rect 2460 -3417 2510 -3400
rect 2352 -3434 2368 -3417
rect 2236 -3450 2368 -3434
rect 2494 -3434 2510 -3417
rect 2610 -3417 2660 -3400
rect 2718 -3400 2918 -3362
rect 2718 -3417 2768 -3400
rect 2610 -3434 2626 -3417
rect 2494 -3450 2626 -3434
rect 2752 -3434 2768 -3417
rect 2868 -3417 2918 -3400
rect 2976 -3400 3176 -3362
rect 2976 -3417 3026 -3400
rect 2868 -3434 2884 -3417
rect 2752 -3450 2884 -3434
rect 3010 -3434 3026 -3417
rect 3126 -3417 3176 -3400
rect 3234 -3400 3434 -3362
rect 3234 -3417 3284 -3400
rect 3126 -3434 3142 -3417
rect 3010 -3450 3142 -3434
rect 3268 -3434 3284 -3417
rect 3384 -3417 3434 -3400
rect 3492 -3400 3692 -3362
rect 3492 -3417 3542 -3400
rect 3384 -3434 3400 -3417
rect 3268 -3450 3400 -3434
rect 3526 -3434 3542 -3417
rect 3642 -3417 3692 -3400
rect 4466 -3400 4666 -3362
rect 4466 -3417 4516 -3400
rect 3642 -3434 3658 -3417
rect 3526 -3450 3658 -3434
rect 4500 -3434 4516 -3417
rect 4616 -3417 4666 -3400
rect 4724 -3400 4924 -3362
rect 4724 -3417 4774 -3400
rect 4616 -3434 4632 -3417
rect 4500 -3450 4632 -3434
rect 4758 -3434 4774 -3417
rect 4874 -3417 4924 -3400
rect 4982 -3400 5182 -3362
rect 4982 -3417 5032 -3400
rect 4874 -3434 4890 -3417
rect 4758 -3450 4890 -3434
rect 5016 -3434 5032 -3417
rect 5132 -3417 5182 -3400
rect 5240 -3400 5440 -3362
rect 5240 -3417 5290 -3400
rect 5132 -3434 5148 -3417
rect 5016 -3450 5148 -3434
rect 5274 -3434 5290 -3417
rect 5390 -3417 5440 -3400
rect 5498 -3400 5698 -3362
rect 5498 -3417 5548 -3400
rect 5390 -3434 5406 -3417
rect 5274 -3450 5406 -3434
rect 5532 -3434 5548 -3417
rect 5648 -3417 5698 -3400
rect 5756 -3400 5956 -3362
rect 5756 -3417 5806 -3400
rect 5648 -3434 5664 -3417
rect 5532 -3450 5664 -3434
rect 5790 -3434 5806 -3417
rect 5906 -3417 5956 -3400
rect 6014 -3400 6214 -3362
rect 6014 -3417 6064 -3400
rect 5906 -3434 5922 -3417
rect 5790 -3450 5922 -3434
rect 6048 -3434 6064 -3417
rect 6164 -3417 6214 -3400
rect 6272 -3400 6472 -3362
rect 6272 -3417 6322 -3400
rect 6164 -3434 6180 -3417
rect 6048 -3450 6180 -3434
rect 6306 -3434 6322 -3417
rect 6422 -3417 6472 -3400
rect 6530 -3400 6730 -3362
rect 6530 -3417 6580 -3400
rect 6422 -3434 6438 -3417
rect 6306 -3450 6438 -3434
rect 6564 -3434 6580 -3417
rect 6680 -3417 6730 -3400
rect 6788 -3400 6988 -3362
rect 6788 -3417 6838 -3400
rect 6680 -3434 6696 -3417
rect 6564 -3450 6696 -3434
rect 6822 -3434 6838 -3417
rect 6938 -3417 6988 -3400
rect 7762 -3400 7962 -3362
rect 7762 -3417 7812 -3400
rect 6938 -3434 6954 -3417
rect 6822 -3450 6954 -3434
rect 7796 -3434 7812 -3417
rect 7912 -3417 7962 -3400
rect 8020 -3400 8220 -3362
rect 8020 -3417 8070 -3400
rect 7912 -3434 7928 -3417
rect 7796 -3450 7928 -3434
rect 8054 -3434 8070 -3417
rect 8170 -3417 8220 -3400
rect 8278 -3400 8478 -3362
rect 8278 -3417 8328 -3400
rect 8170 -3434 8186 -3417
rect 8054 -3450 8186 -3434
rect 8312 -3434 8328 -3417
rect 8428 -3417 8478 -3400
rect 8536 -3400 8736 -3362
rect 8536 -3417 8586 -3400
rect 8428 -3434 8444 -3417
rect 8312 -3450 8444 -3434
rect 8570 -3434 8586 -3417
rect 8686 -3417 8736 -3400
rect 8794 -3400 8994 -3362
rect 8794 -3417 8844 -3400
rect 8686 -3434 8702 -3417
rect 8570 -3450 8702 -3434
rect 8828 -3434 8844 -3417
rect 8944 -3417 8994 -3400
rect 9052 -3400 9252 -3362
rect 9052 -3417 9102 -3400
rect 8944 -3434 8960 -3417
rect 8828 -3450 8960 -3434
rect 9086 -3434 9102 -3417
rect 9202 -3417 9252 -3400
rect 9310 -3400 9510 -3362
rect 9310 -3417 9360 -3400
rect 9202 -3434 9218 -3417
rect 9086 -3450 9218 -3434
rect 9344 -3434 9360 -3417
rect 9460 -3417 9510 -3400
rect 9568 -3400 9768 -3362
rect 9568 -3417 9618 -3400
rect 9460 -3434 9476 -3417
rect 9344 -3450 9476 -3434
rect 9602 -3434 9618 -3417
rect 9718 -3417 9768 -3400
rect 9826 -3400 10026 -3362
rect 9826 -3417 9876 -3400
rect 9718 -3434 9734 -3417
rect 9602 -3450 9734 -3434
rect 9860 -3434 9876 -3417
rect 9976 -3417 10026 -3400
rect 10084 -3400 10284 -3362
rect 10084 -3417 10134 -3400
rect 9976 -3434 9992 -3417
rect 9860 -3450 9992 -3434
rect 10118 -3434 10134 -3417
rect 10234 -3417 10284 -3400
rect 10234 -3434 10250 -3417
rect 10118 -3450 10250 -3434
rect 12576 -1442 13068 -1426
rect 12576 -1459 12592 -1442
rect 12422 -1476 12592 -1459
rect 13052 -1459 13068 -1442
rect 13434 -1442 13926 -1426
rect 13434 -1459 13450 -1442
rect 13052 -1476 13222 -1459
rect 12422 -1514 13222 -1476
rect 13280 -1476 13450 -1459
rect 13910 -1459 13926 -1442
rect 14292 -1442 14784 -1426
rect 14292 -1459 14308 -1442
rect 13910 -1476 14080 -1459
rect 13280 -1514 14080 -1476
rect 14138 -1476 14308 -1459
rect 14768 -1459 14784 -1442
rect 15150 -1442 15642 -1426
rect 15150 -1459 15166 -1442
rect 14768 -1476 14938 -1459
rect 14138 -1514 14938 -1476
rect 14996 -1476 15166 -1459
rect 15626 -1459 15642 -1442
rect 16008 -1442 16500 -1426
rect 16008 -1459 16024 -1442
rect 15626 -1476 15796 -1459
rect 14996 -1514 15796 -1476
rect 15854 -1476 16024 -1459
rect 16484 -1459 16500 -1442
rect 16866 -1442 17358 -1426
rect 16866 -1459 16882 -1442
rect 16484 -1476 16654 -1459
rect 15854 -1514 16654 -1476
rect 16712 -1476 16882 -1459
rect 17342 -1459 17358 -1442
rect 17724 -1442 18216 -1426
rect 17724 -1459 17740 -1442
rect 17342 -1476 17512 -1459
rect 16712 -1514 17512 -1476
rect 17570 -1476 17740 -1459
rect 18200 -1459 18216 -1442
rect 18582 -1442 19074 -1426
rect 18582 -1459 18598 -1442
rect 18200 -1476 18370 -1459
rect 17570 -1514 18370 -1476
rect 18428 -1476 18598 -1459
rect 19058 -1459 19074 -1442
rect 19440 -1442 19932 -1426
rect 19440 -1459 19456 -1442
rect 19058 -1476 19228 -1459
rect 18428 -1514 19228 -1476
rect 19286 -1476 19456 -1459
rect 19916 -1459 19932 -1442
rect 20298 -1442 20790 -1426
rect 20298 -1459 20314 -1442
rect 19916 -1476 20086 -1459
rect 19286 -1514 20086 -1476
rect 20144 -1476 20314 -1459
rect 20774 -1459 20790 -1442
rect 21156 -1442 21648 -1426
rect 21156 -1459 21172 -1442
rect 20774 -1476 20944 -1459
rect 20144 -1514 20944 -1476
rect 21002 -1476 21172 -1459
rect 21632 -1459 21648 -1442
rect 22014 -1442 22506 -1426
rect 22014 -1459 22030 -1442
rect 21632 -1476 21802 -1459
rect 21002 -1514 21802 -1476
rect 21860 -1476 22030 -1459
rect 22490 -1459 22506 -1442
rect 22490 -1476 22660 -1459
rect 21860 -1514 22660 -1476
rect 12422 -1752 13222 -1714
rect 12422 -1769 12592 -1752
rect 12576 -1786 12592 -1769
rect 13052 -1769 13222 -1752
rect 13280 -1752 14080 -1714
rect 13280 -1769 13450 -1752
rect 13052 -1786 13068 -1769
rect 12576 -1802 13068 -1786
rect 13434 -1786 13450 -1769
rect 13910 -1769 14080 -1752
rect 14138 -1752 14938 -1714
rect 14138 -1769 14308 -1752
rect 13910 -1786 13926 -1769
rect 13434 -1802 13926 -1786
rect 14292 -1786 14308 -1769
rect 14768 -1769 14938 -1752
rect 14996 -1752 15796 -1714
rect 14996 -1769 15166 -1752
rect 14768 -1786 14784 -1769
rect 14292 -1802 14784 -1786
rect 15150 -1786 15166 -1769
rect 15626 -1769 15796 -1752
rect 15854 -1752 16654 -1714
rect 15854 -1769 16024 -1752
rect 15626 -1786 15642 -1769
rect 15150 -1802 15642 -1786
rect 16008 -1786 16024 -1769
rect 16484 -1769 16654 -1752
rect 16712 -1752 17512 -1714
rect 16712 -1769 16882 -1752
rect 16484 -1786 16500 -1769
rect 16008 -1802 16500 -1786
rect 16866 -1786 16882 -1769
rect 17342 -1769 17512 -1752
rect 17570 -1752 18370 -1714
rect 17570 -1769 17740 -1752
rect 17342 -1786 17358 -1769
rect 16866 -1802 17358 -1786
rect 17724 -1786 17740 -1769
rect 18200 -1769 18370 -1752
rect 18428 -1752 19228 -1714
rect 18428 -1769 18598 -1752
rect 18200 -1786 18216 -1769
rect 17724 -1802 18216 -1786
rect 18582 -1786 18598 -1769
rect 19058 -1769 19228 -1752
rect 19286 -1752 20086 -1714
rect 19286 -1769 19456 -1752
rect 19058 -1786 19074 -1769
rect 18582 -1802 19074 -1786
rect 19440 -1786 19456 -1769
rect 19916 -1769 20086 -1752
rect 20144 -1752 20944 -1714
rect 20144 -1769 20314 -1752
rect 19916 -1786 19932 -1769
rect 19440 -1802 19932 -1786
rect 20298 -1786 20314 -1769
rect 20774 -1769 20944 -1752
rect 21002 -1752 21802 -1714
rect 21002 -1769 21172 -1752
rect 20774 -1786 20790 -1769
rect 20298 -1802 20790 -1786
rect 21156 -1786 21172 -1769
rect 21632 -1769 21802 -1752
rect 21860 -1752 22660 -1714
rect 21860 -1769 22030 -1752
rect 21632 -1786 21648 -1769
rect 21156 -1802 21648 -1786
rect 22014 -1786 22030 -1769
rect 22490 -1769 22660 -1752
rect 22490 -1786 22506 -1769
rect 22014 -1802 22506 -1786
rect 12576 -1982 13068 -1966
rect 12576 -1999 12592 -1982
rect 12422 -2016 12592 -1999
rect 13052 -1999 13068 -1982
rect 13434 -1982 13926 -1966
rect 13434 -1999 13450 -1982
rect 13052 -2016 13222 -1999
rect 12422 -2054 13222 -2016
rect 13280 -2016 13450 -1999
rect 13910 -1999 13926 -1982
rect 14292 -1982 14784 -1966
rect 14292 -1999 14308 -1982
rect 13910 -2016 14080 -1999
rect 13280 -2054 14080 -2016
rect 14138 -2016 14308 -1999
rect 14768 -1999 14784 -1982
rect 15150 -1982 15642 -1966
rect 15150 -1999 15166 -1982
rect 14768 -2016 14938 -1999
rect 14138 -2054 14938 -2016
rect 14996 -2016 15166 -1999
rect 15626 -1999 15642 -1982
rect 16008 -1982 16500 -1966
rect 16008 -1999 16024 -1982
rect 15626 -2016 15796 -1999
rect 14996 -2054 15796 -2016
rect 15854 -2016 16024 -1999
rect 16484 -1999 16500 -1982
rect 16866 -1982 17358 -1966
rect 16866 -1999 16882 -1982
rect 16484 -2016 16654 -1999
rect 15854 -2054 16654 -2016
rect 16712 -2016 16882 -1999
rect 17342 -1999 17358 -1982
rect 17724 -1982 18216 -1966
rect 17724 -1999 17740 -1982
rect 17342 -2016 17512 -1999
rect 16712 -2054 17512 -2016
rect 17570 -2016 17740 -1999
rect 18200 -1999 18216 -1982
rect 18582 -1982 19074 -1966
rect 18582 -1999 18598 -1982
rect 18200 -2016 18370 -1999
rect 17570 -2054 18370 -2016
rect 18428 -2016 18598 -1999
rect 19058 -1999 19074 -1982
rect 19440 -1982 19932 -1966
rect 19440 -1999 19456 -1982
rect 19058 -2016 19228 -1999
rect 18428 -2054 19228 -2016
rect 19286 -2016 19456 -1999
rect 19916 -1999 19932 -1982
rect 20298 -1982 20790 -1966
rect 20298 -1999 20314 -1982
rect 19916 -2016 20086 -1999
rect 19286 -2054 20086 -2016
rect 20144 -2016 20314 -1999
rect 20774 -1999 20790 -1982
rect 21156 -1982 21648 -1966
rect 21156 -1999 21172 -1982
rect 20774 -2016 20944 -1999
rect 20144 -2054 20944 -2016
rect 21002 -2016 21172 -1999
rect 21632 -1999 21648 -1982
rect 22014 -1982 22506 -1966
rect 22014 -1999 22030 -1982
rect 21632 -2016 21802 -1999
rect 21002 -2054 21802 -2016
rect 21860 -2016 22030 -1999
rect 22490 -1999 22506 -1982
rect 22490 -2016 22660 -1999
rect 21860 -2054 22660 -2016
rect 12422 -2292 13222 -2254
rect 12422 -2309 12592 -2292
rect 12576 -2326 12592 -2309
rect 13052 -2309 13222 -2292
rect 13280 -2292 14080 -2254
rect 13280 -2309 13450 -2292
rect 13052 -2326 13068 -2309
rect 12576 -2342 13068 -2326
rect 13434 -2326 13450 -2309
rect 13910 -2309 14080 -2292
rect 14138 -2292 14938 -2254
rect 14138 -2309 14308 -2292
rect 13910 -2326 13926 -2309
rect 13434 -2342 13926 -2326
rect 14292 -2326 14308 -2309
rect 14768 -2309 14938 -2292
rect 14996 -2292 15796 -2254
rect 14996 -2309 15166 -2292
rect 14768 -2326 14784 -2309
rect 14292 -2342 14784 -2326
rect 15150 -2326 15166 -2309
rect 15626 -2309 15796 -2292
rect 15854 -2292 16654 -2254
rect 15854 -2309 16024 -2292
rect 15626 -2326 15642 -2309
rect 15150 -2342 15642 -2326
rect 16008 -2326 16024 -2309
rect 16484 -2309 16654 -2292
rect 16712 -2292 17512 -2254
rect 16712 -2309 16882 -2292
rect 16484 -2326 16500 -2309
rect 16008 -2342 16500 -2326
rect 16866 -2326 16882 -2309
rect 17342 -2309 17512 -2292
rect 17570 -2292 18370 -2254
rect 17570 -2309 17740 -2292
rect 17342 -2326 17358 -2309
rect 16866 -2342 17358 -2326
rect 17724 -2326 17740 -2309
rect 18200 -2309 18370 -2292
rect 18428 -2292 19228 -2254
rect 18428 -2309 18598 -2292
rect 18200 -2326 18216 -2309
rect 17724 -2342 18216 -2326
rect 18582 -2326 18598 -2309
rect 19058 -2309 19228 -2292
rect 19286 -2292 20086 -2254
rect 19286 -2309 19456 -2292
rect 19058 -2326 19074 -2309
rect 18582 -2342 19074 -2326
rect 19440 -2326 19456 -2309
rect 19916 -2309 20086 -2292
rect 20144 -2292 20944 -2254
rect 20144 -2309 20314 -2292
rect 19916 -2326 19932 -2309
rect 19440 -2342 19932 -2326
rect 20298 -2326 20314 -2309
rect 20774 -2309 20944 -2292
rect 21002 -2292 21802 -2254
rect 21002 -2309 21172 -2292
rect 20774 -2326 20790 -2309
rect 20298 -2342 20790 -2326
rect 21156 -2326 21172 -2309
rect 21632 -2309 21802 -2292
rect 21860 -2292 22660 -2254
rect 21860 -2309 22030 -2292
rect 21632 -2326 21648 -2309
rect 21156 -2342 21648 -2326
rect 22014 -2326 22030 -2309
rect 22490 -2309 22660 -2292
rect 22490 -2326 22506 -2309
rect 22014 -2342 22506 -2326
rect 13004 -2890 13136 -2874
rect 13004 -2907 13020 -2890
rect 12970 -2924 13020 -2907
rect 13120 -2907 13136 -2890
rect 13262 -2890 13394 -2874
rect 13262 -2907 13278 -2890
rect 13120 -2924 13170 -2907
rect 12970 -2962 13170 -2924
rect 13228 -2924 13278 -2907
rect 13378 -2907 13394 -2890
rect 13520 -2890 13652 -2874
rect 13520 -2907 13536 -2890
rect 13378 -2924 13428 -2907
rect 13228 -2962 13428 -2924
rect 13486 -2924 13536 -2907
rect 13636 -2907 13652 -2890
rect 13778 -2890 13910 -2874
rect 13778 -2907 13794 -2890
rect 13636 -2924 13686 -2907
rect 13486 -2962 13686 -2924
rect 13744 -2924 13794 -2907
rect 13894 -2907 13910 -2890
rect 14036 -2890 14168 -2874
rect 14036 -2907 14052 -2890
rect 13894 -2924 13944 -2907
rect 13744 -2962 13944 -2924
rect 14002 -2924 14052 -2907
rect 14152 -2907 14168 -2890
rect 14294 -2890 14426 -2874
rect 14294 -2907 14310 -2890
rect 14152 -2924 14202 -2907
rect 14002 -2962 14202 -2924
rect 14260 -2924 14310 -2907
rect 14410 -2907 14426 -2890
rect 14552 -2890 14684 -2874
rect 14552 -2907 14568 -2890
rect 14410 -2924 14460 -2907
rect 14260 -2962 14460 -2924
rect 14518 -2924 14568 -2907
rect 14668 -2907 14684 -2890
rect 14810 -2890 14942 -2874
rect 14810 -2907 14826 -2890
rect 14668 -2924 14718 -2907
rect 14518 -2962 14718 -2924
rect 14776 -2924 14826 -2907
rect 14926 -2907 14942 -2890
rect 15068 -2890 15200 -2874
rect 15068 -2907 15084 -2890
rect 14926 -2924 14976 -2907
rect 14776 -2962 14976 -2924
rect 15034 -2924 15084 -2907
rect 15184 -2907 15200 -2890
rect 15326 -2890 15458 -2874
rect 15326 -2907 15342 -2890
rect 15184 -2924 15234 -2907
rect 15034 -2962 15234 -2924
rect 15292 -2924 15342 -2907
rect 15442 -2907 15458 -2890
rect 16300 -2890 16432 -2874
rect 16300 -2907 16316 -2890
rect 15442 -2924 15492 -2907
rect 15292 -2962 15492 -2924
rect 16266 -2924 16316 -2907
rect 16416 -2907 16432 -2890
rect 16558 -2890 16690 -2874
rect 16558 -2907 16574 -2890
rect 16416 -2924 16466 -2907
rect 16266 -2962 16466 -2924
rect 16524 -2924 16574 -2907
rect 16674 -2907 16690 -2890
rect 16816 -2890 16948 -2874
rect 16816 -2907 16832 -2890
rect 16674 -2924 16724 -2907
rect 16524 -2962 16724 -2924
rect 16782 -2924 16832 -2907
rect 16932 -2907 16948 -2890
rect 17074 -2890 17206 -2874
rect 17074 -2907 17090 -2890
rect 16932 -2924 16982 -2907
rect 16782 -2962 16982 -2924
rect 17040 -2924 17090 -2907
rect 17190 -2907 17206 -2890
rect 17332 -2890 17464 -2874
rect 17332 -2907 17348 -2890
rect 17190 -2924 17240 -2907
rect 17040 -2962 17240 -2924
rect 17298 -2924 17348 -2907
rect 17448 -2907 17464 -2890
rect 17590 -2890 17722 -2874
rect 17590 -2907 17606 -2890
rect 17448 -2924 17498 -2907
rect 17298 -2962 17498 -2924
rect 17556 -2924 17606 -2907
rect 17706 -2907 17722 -2890
rect 17848 -2890 17980 -2874
rect 17848 -2907 17864 -2890
rect 17706 -2924 17756 -2907
rect 17556 -2962 17756 -2924
rect 17814 -2924 17864 -2907
rect 17964 -2907 17980 -2890
rect 18106 -2890 18238 -2874
rect 18106 -2907 18122 -2890
rect 17964 -2924 18014 -2907
rect 17814 -2962 18014 -2924
rect 18072 -2924 18122 -2907
rect 18222 -2907 18238 -2890
rect 18364 -2890 18496 -2874
rect 18364 -2907 18380 -2890
rect 18222 -2924 18272 -2907
rect 18072 -2962 18272 -2924
rect 18330 -2924 18380 -2907
rect 18480 -2907 18496 -2890
rect 18622 -2890 18754 -2874
rect 18622 -2907 18638 -2890
rect 18480 -2924 18530 -2907
rect 18330 -2962 18530 -2924
rect 18588 -2924 18638 -2907
rect 18738 -2907 18754 -2890
rect 19596 -2890 19728 -2874
rect 19596 -2907 19612 -2890
rect 18738 -2924 18788 -2907
rect 18588 -2962 18788 -2924
rect 19562 -2924 19612 -2907
rect 19712 -2907 19728 -2890
rect 19854 -2890 19986 -2874
rect 19854 -2907 19870 -2890
rect 19712 -2924 19762 -2907
rect 19562 -2962 19762 -2924
rect 19820 -2924 19870 -2907
rect 19970 -2907 19986 -2890
rect 20112 -2890 20244 -2874
rect 20112 -2907 20128 -2890
rect 19970 -2924 20020 -2907
rect 19820 -2962 20020 -2924
rect 20078 -2924 20128 -2907
rect 20228 -2907 20244 -2890
rect 20370 -2890 20502 -2874
rect 20370 -2907 20386 -2890
rect 20228 -2924 20278 -2907
rect 20078 -2962 20278 -2924
rect 20336 -2924 20386 -2907
rect 20486 -2907 20502 -2890
rect 20628 -2890 20760 -2874
rect 20628 -2907 20644 -2890
rect 20486 -2924 20536 -2907
rect 20336 -2962 20536 -2924
rect 20594 -2924 20644 -2907
rect 20744 -2907 20760 -2890
rect 20886 -2890 21018 -2874
rect 20886 -2907 20902 -2890
rect 20744 -2924 20794 -2907
rect 20594 -2962 20794 -2924
rect 20852 -2924 20902 -2907
rect 21002 -2907 21018 -2890
rect 21144 -2890 21276 -2874
rect 21144 -2907 21160 -2890
rect 21002 -2924 21052 -2907
rect 20852 -2962 21052 -2924
rect 21110 -2924 21160 -2907
rect 21260 -2907 21276 -2890
rect 21402 -2890 21534 -2874
rect 21402 -2907 21418 -2890
rect 21260 -2924 21310 -2907
rect 21110 -2962 21310 -2924
rect 21368 -2924 21418 -2907
rect 21518 -2907 21534 -2890
rect 21660 -2890 21792 -2874
rect 21660 -2907 21676 -2890
rect 21518 -2924 21568 -2907
rect 21368 -2962 21568 -2924
rect 21626 -2924 21676 -2907
rect 21776 -2907 21792 -2890
rect 21918 -2890 22050 -2874
rect 21918 -2907 21934 -2890
rect 21776 -2924 21826 -2907
rect 21626 -2962 21826 -2924
rect 21884 -2924 21934 -2907
rect 22034 -2907 22050 -2890
rect 22034 -2924 22084 -2907
rect 21884 -2962 22084 -2924
rect 12970 -3400 13170 -3362
rect 12970 -3417 13020 -3400
rect 13004 -3434 13020 -3417
rect 13120 -3417 13170 -3400
rect 13228 -3400 13428 -3362
rect 13228 -3417 13278 -3400
rect 13120 -3434 13136 -3417
rect 13004 -3450 13136 -3434
rect 13262 -3434 13278 -3417
rect 13378 -3417 13428 -3400
rect 13486 -3400 13686 -3362
rect 13486 -3417 13536 -3400
rect 13378 -3434 13394 -3417
rect 13262 -3450 13394 -3434
rect 13520 -3434 13536 -3417
rect 13636 -3417 13686 -3400
rect 13744 -3400 13944 -3362
rect 13744 -3417 13794 -3400
rect 13636 -3434 13652 -3417
rect 13520 -3450 13652 -3434
rect 13778 -3434 13794 -3417
rect 13894 -3417 13944 -3400
rect 14002 -3400 14202 -3362
rect 14002 -3417 14052 -3400
rect 13894 -3434 13910 -3417
rect 13778 -3450 13910 -3434
rect 14036 -3434 14052 -3417
rect 14152 -3417 14202 -3400
rect 14260 -3400 14460 -3362
rect 14260 -3417 14310 -3400
rect 14152 -3434 14168 -3417
rect 14036 -3450 14168 -3434
rect 14294 -3434 14310 -3417
rect 14410 -3417 14460 -3400
rect 14518 -3400 14718 -3362
rect 14518 -3417 14568 -3400
rect 14410 -3434 14426 -3417
rect 14294 -3450 14426 -3434
rect 14552 -3434 14568 -3417
rect 14668 -3417 14718 -3400
rect 14776 -3400 14976 -3362
rect 14776 -3417 14826 -3400
rect 14668 -3434 14684 -3417
rect 14552 -3450 14684 -3434
rect 14810 -3434 14826 -3417
rect 14926 -3417 14976 -3400
rect 15034 -3400 15234 -3362
rect 15034 -3417 15084 -3400
rect 14926 -3434 14942 -3417
rect 14810 -3450 14942 -3434
rect 15068 -3434 15084 -3417
rect 15184 -3417 15234 -3400
rect 15292 -3400 15492 -3362
rect 15292 -3417 15342 -3400
rect 15184 -3434 15200 -3417
rect 15068 -3450 15200 -3434
rect 15326 -3434 15342 -3417
rect 15442 -3417 15492 -3400
rect 16266 -3400 16466 -3362
rect 16266 -3417 16316 -3400
rect 15442 -3434 15458 -3417
rect 15326 -3450 15458 -3434
rect 16300 -3434 16316 -3417
rect 16416 -3417 16466 -3400
rect 16524 -3400 16724 -3362
rect 16524 -3417 16574 -3400
rect 16416 -3434 16432 -3417
rect 16300 -3450 16432 -3434
rect 16558 -3434 16574 -3417
rect 16674 -3417 16724 -3400
rect 16782 -3400 16982 -3362
rect 16782 -3417 16832 -3400
rect 16674 -3434 16690 -3417
rect 16558 -3450 16690 -3434
rect 16816 -3434 16832 -3417
rect 16932 -3417 16982 -3400
rect 17040 -3400 17240 -3362
rect 17040 -3417 17090 -3400
rect 16932 -3434 16948 -3417
rect 16816 -3450 16948 -3434
rect 17074 -3434 17090 -3417
rect 17190 -3417 17240 -3400
rect 17298 -3400 17498 -3362
rect 17298 -3417 17348 -3400
rect 17190 -3434 17206 -3417
rect 17074 -3450 17206 -3434
rect 17332 -3434 17348 -3417
rect 17448 -3417 17498 -3400
rect 17556 -3400 17756 -3362
rect 17556 -3417 17606 -3400
rect 17448 -3434 17464 -3417
rect 17332 -3450 17464 -3434
rect 17590 -3434 17606 -3417
rect 17706 -3417 17756 -3400
rect 17814 -3400 18014 -3362
rect 17814 -3417 17864 -3400
rect 17706 -3434 17722 -3417
rect 17590 -3450 17722 -3434
rect 17848 -3434 17864 -3417
rect 17964 -3417 18014 -3400
rect 18072 -3400 18272 -3362
rect 18072 -3417 18122 -3400
rect 17964 -3434 17980 -3417
rect 17848 -3450 17980 -3434
rect 18106 -3434 18122 -3417
rect 18222 -3417 18272 -3400
rect 18330 -3400 18530 -3362
rect 18330 -3417 18380 -3400
rect 18222 -3434 18238 -3417
rect 18106 -3450 18238 -3434
rect 18364 -3434 18380 -3417
rect 18480 -3417 18530 -3400
rect 18588 -3400 18788 -3362
rect 18588 -3417 18638 -3400
rect 18480 -3434 18496 -3417
rect 18364 -3450 18496 -3434
rect 18622 -3434 18638 -3417
rect 18738 -3417 18788 -3400
rect 19562 -3400 19762 -3362
rect 19562 -3417 19612 -3400
rect 18738 -3434 18754 -3417
rect 18622 -3450 18754 -3434
rect 19596 -3434 19612 -3417
rect 19712 -3417 19762 -3400
rect 19820 -3400 20020 -3362
rect 19820 -3417 19870 -3400
rect 19712 -3434 19728 -3417
rect 19596 -3450 19728 -3434
rect 19854 -3434 19870 -3417
rect 19970 -3417 20020 -3400
rect 20078 -3400 20278 -3362
rect 20078 -3417 20128 -3400
rect 19970 -3434 19986 -3417
rect 19854 -3450 19986 -3434
rect 20112 -3434 20128 -3417
rect 20228 -3417 20278 -3400
rect 20336 -3400 20536 -3362
rect 20336 -3417 20386 -3400
rect 20228 -3434 20244 -3417
rect 20112 -3450 20244 -3434
rect 20370 -3434 20386 -3417
rect 20486 -3417 20536 -3400
rect 20594 -3400 20794 -3362
rect 20594 -3417 20644 -3400
rect 20486 -3434 20502 -3417
rect 20370 -3450 20502 -3434
rect 20628 -3434 20644 -3417
rect 20744 -3417 20794 -3400
rect 20852 -3400 21052 -3362
rect 20852 -3417 20902 -3400
rect 20744 -3434 20760 -3417
rect 20628 -3450 20760 -3434
rect 20886 -3434 20902 -3417
rect 21002 -3417 21052 -3400
rect 21110 -3400 21310 -3362
rect 21110 -3417 21160 -3400
rect 21002 -3434 21018 -3417
rect 20886 -3450 21018 -3434
rect 21144 -3434 21160 -3417
rect 21260 -3417 21310 -3400
rect 21368 -3400 21568 -3362
rect 21368 -3417 21418 -3400
rect 21260 -3434 21276 -3417
rect 21144 -3450 21276 -3434
rect 21402 -3434 21418 -3417
rect 21518 -3417 21568 -3400
rect 21626 -3400 21826 -3362
rect 21626 -3417 21676 -3400
rect 21518 -3434 21534 -3417
rect 21402 -3450 21534 -3434
rect 21660 -3434 21676 -3417
rect 21776 -3417 21826 -3400
rect 21884 -3400 22084 -3362
rect 21884 -3417 21934 -3400
rect 21776 -3434 21792 -3417
rect 21660 -3450 21792 -3434
rect 21918 -3434 21934 -3417
rect 22034 -3417 22084 -3400
rect 22034 -3434 22050 -3417
rect 21918 -3450 22050 -3434
rect 3988 -4549 4120 -4533
rect 3988 -4566 4004 -4549
rect 3954 -4583 4004 -4566
rect 4104 -4566 4120 -4549
rect 4246 -4549 4378 -4533
rect 4246 -4566 4262 -4549
rect 4104 -4583 4154 -4566
rect 3954 -4630 4154 -4583
rect 4212 -4583 4262 -4566
rect 4362 -4566 4378 -4549
rect 4504 -4549 4636 -4533
rect 4504 -4566 4520 -4549
rect 4362 -4583 4412 -4566
rect 4212 -4630 4412 -4583
rect 4470 -4583 4520 -4566
rect 4620 -4566 4636 -4549
rect 4762 -4549 4894 -4533
rect 4762 -4566 4778 -4549
rect 4620 -4583 4670 -4566
rect 4470 -4630 4670 -4583
rect 4728 -4583 4778 -4566
rect 4878 -4566 4894 -4549
rect 5020 -4549 5152 -4533
rect 5020 -4566 5036 -4549
rect 4878 -4583 4928 -4566
rect 4728 -4630 4928 -4583
rect 4986 -4583 5036 -4566
rect 5136 -4566 5152 -4549
rect 5278 -4549 5410 -4533
rect 5278 -4566 5294 -4549
rect 5136 -4583 5186 -4566
rect 4986 -4630 5186 -4583
rect 5244 -4583 5294 -4566
rect 5394 -4566 5410 -4549
rect 5536 -4549 5668 -4533
rect 5536 -4566 5552 -4549
rect 5394 -4583 5444 -4566
rect 5244 -4630 5444 -4583
rect 5502 -4583 5552 -4566
rect 5652 -4566 5668 -4549
rect 5794 -4549 5926 -4533
rect 5794 -4566 5810 -4549
rect 5652 -4583 5702 -4566
rect 5502 -4630 5702 -4583
rect 5760 -4583 5810 -4566
rect 5910 -4566 5926 -4549
rect 6052 -4549 6184 -4533
rect 6052 -4566 6068 -4549
rect 5910 -4583 5960 -4566
rect 5760 -4630 5960 -4583
rect 6018 -4583 6068 -4566
rect 6168 -4566 6184 -4549
rect 6310 -4549 6442 -4533
rect 6310 -4566 6326 -4549
rect 6168 -4583 6218 -4566
rect 6018 -4630 6218 -4583
rect 6276 -4583 6326 -4566
rect 6426 -4566 6442 -4549
rect 6568 -4549 6700 -4533
rect 6568 -4566 6584 -4549
rect 6426 -4583 6476 -4566
rect 6276 -4630 6476 -4583
rect 6534 -4583 6584 -4566
rect 6684 -4566 6700 -4549
rect 6826 -4549 6958 -4533
rect 6826 -4566 6842 -4549
rect 6684 -4583 6734 -4566
rect 6534 -4630 6734 -4583
rect 6792 -4583 6842 -4566
rect 6942 -4566 6958 -4549
rect 7084 -4549 7216 -4533
rect 7084 -4566 7100 -4549
rect 6942 -4583 6992 -4566
rect 6792 -4630 6992 -4583
rect 7050 -4583 7100 -4566
rect 7200 -4566 7216 -4549
rect 7342 -4549 7474 -4533
rect 7342 -4566 7358 -4549
rect 7200 -4583 7250 -4566
rect 7050 -4630 7250 -4583
rect 7308 -4583 7358 -4566
rect 7458 -4566 7474 -4549
rect 7458 -4583 7508 -4566
rect 7308 -4630 7508 -4583
rect 3954 -4877 4154 -4830
rect 3954 -4894 4004 -4877
rect 3988 -4911 4004 -4894
rect 4104 -4894 4154 -4877
rect 4212 -4877 4412 -4830
rect 4212 -4894 4262 -4877
rect 4104 -4911 4120 -4894
rect 3988 -4927 4120 -4911
rect 4246 -4911 4262 -4894
rect 4362 -4894 4412 -4877
rect 4470 -4877 4670 -4830
rect 4470 -4894 4520 -4877
rect 4362 -4911 4378 -4894
rect 4246 -4927 4378 -4911
rect 4504 -4911 4520 -4894
rect 4620 -4894 4670 -4877
rect 4728 -4877 4928 -4830
rect 4728 -4894 4778 -4877
rect 4620 -4911 4636 -4894
rect 4504 -4927 4636 -4911
rect 4762 -4911 4778 -4894
rect 4878 -4894 4928 -4877
rect 4986 -4877 5186 -4830
rect 4986 -4894 5036 -4877
rect 4878 -4911 4894 -4894
rect 4762 -4927 4894 -4911
rect 5020 -4911 5036 -4894
rect 5136 -4894 5186 -4877
rect 5244 -4877 5444 -4830
rect 5244 -4894 5294 -4877
rect 5136 -4911 5152 -4894
rect 5020 -4927 5152 -4911
rect 5278 -4911 5294 -4894
rect 5394 -4894 5444 -4877
rect 5502 -4877 5702 -4830
rect 5502 -4894 5552 -4877
rect 5394 -4911 5410 -4894
rect 5278 -4927 5410 -4911
rect 5536 -4911 5552 -4894
rect 5652 -4894 5702 -4877
rect 5760 -4877 5960 -4830
rect 5760 -4894 5810 -4877
rect 5652 -4911 5668 -4894
rect 5536 -4927 5668 -4911
rect 5794 -4911 5810 -4894
rect 5910 -4894 5960 -4877
rect 6018 -4877 6218 -4830
rect 6018 -4894 6068 -4877
rect 5910 -4911 5926 -4894
rect 5794 -4927 5926 -4911
rect 6052 -4911 6068 -4894
rect 6168 -4894 6218 -4877
rect 6276 -4877 6476 -4830
rect 6276 -4894 6326 -4877
rect 6168 -4911 6184 -4894
rect 6052 -4927 6184 -4911
rect 6310 -4911 6326 -4894
rect 6426 -4894 6476 -4877
rect 6534 -4877 6734 -4830
rect 6534 -4894 6584 -4877
rect 6426 -4911 6442 -4894
rect 6310 -4927 6442 -4911
rect 6568 -4911 6584 -4894
rect 6684 -4894 6734 -4877
rect 6792 -4877 6992 -4830
rect 6792 -4894 6842 -4877
rect 6684 -4911 6700 -4894
rect 6568 -4927 6700 -4911
rect 6826 -4911 6842 -4894
rect 6942 -4894 6992 -4877
rect 7050 -4877 7250 -4830
rect 7050 -4894 7100 -4877
rect 6942 -4911 6958 -4894
rect 6826 -4927 6958 -4911
rect 7084 -4911 7100 -4894
rect 7200 -4894 7250 -4877
rect 7308 -4877 7508 -4830
rect 7308 -4894 7358 -4877
rect 7200 -4911 7216 -4894
rect 7084 -4927 7216 -4911
rect 7342 -4911 7358 -4894
rect 7458 -4894 7508 -4877
rect 7458 -4911 7474 -4894
rect 7342 -4927 7474 -4911
rect 15788 -4549 15920 -4533
rect 15788 -4566 15804 -4549
rect 15754 -4583 15804 -4566
rect 15904 -4566 15920 -4549
rect 16046 -4549 16178 -4533
rect 16046 -4566 16062 -4549
rect 15904 -4583 15954 -4566
rect 15754 -4630 15954 -4583
rect 16012 -4583 16062 -4566
rect 16162 -4566 16178 -4549
rect 16304 -4549 16436 -4533
rect 16304 -4566 16320 -4549
rect 16162 -4583 16212 -4566
rect 16012 -4630 16212 -4583
rect 16270 -4583 16320 -4566
rect 16420 -4566 16436 -4549
rect 16562 -4549 16694 -4533
rect 16562 -4566 16578 -4549
rect 16420 -4583 16470 -4566
rect 16270 -4630 16470 -4583
rect 16528 -4583 16578 -4566
rect 16678 -4566 16694 -4549
rect 16820 -4549 16952 -4533
rect 16820 -4566 16836 -4549
rect 16678 -4583 16728 -4566
rect 16528 -4630 16728 -4583
rect 16786 -4583 16836 -4566
rect 16936 -4566 16952 -4549
rect 17078 -4549 17210 -4533
rect 17078 -4566 17094 -4549
rect 16936 -4583 16986 -4566
rect 16786 -4630 16986 -4583
rect 17044 -4583 17094 -4566
rect 17194 -4566 17210 -4549
rect 17336 -4549 17468 -4533
rect 17336 -4566 17352 -4549
rect 17194 -4583 17244 -4566
rect 17044 -4630 17244 -4583
rect 17302 -4583 17352 -4566
rect 17452 -4566 17468 -4549
rect 17594 -4549 17726 -4533
rect 17594 -4566 17610 -4549
rect 17452 -4583 17502 -4566
rect 17302 -4630 17502 -4583
rect 17560 -4583 17610 -4566
rect 17710 -4566 17726 -4549
rect 17852 -4549 17984 -4533
rect 17852 -4566 17868 -4549
rect 17710 -4583 17760 -4566
rect 17560 -4630 17760 -4583
rect 17818 -4583 17868 -4566
rect 17968 -4566 17984 -4549
rect 18110 -4549 18242 -4533
rect 18110 -4566 18126 -4549
rect 17968 -4583 18018 -4566
rect 17818 -4630 18018 -4583
rect 18076 -4583 18126 -4566
rect 18226 -4566 18242 -4549
rect 18368 -4549 18500 -4533
rect 18368 -4566 18384 -4549
rect 18226 -4583 18276 -4566
rect 18076 -4630 18276 -4583
rect 18334 -4583 18384 -4566
rect 18484 -4566 18500 -4549
rect 18626 -4549 18758 -4533
rect 18626 -4566 18642 -4549
rect 18484 -4583 18534 -4566
rect 18334 -4630 18534 -4583
rect 18592 -4583 18642 -4566
rect 18742 -4566 18758 -4549
rect 18884 -4549 19016 -4533
rect 18884 -4566 18900 -4549
rect 18742 -4583 18792 -4566
rect 18592 -4630 18792 -4583
rect 18850 -4583 18900 -4566
rect 19000 -4566 19016 -4549
rect 19142 -4549 19274 -4533
rect 19142 -4566 19158 -4549
rect 19000 -4583 19050 -4566
rect 18850 -4630 19050 -4583
rect 19108 -4583 19158 -4566
rect 19258 -4566 19274 -4549
rect 19258 -4583 19308 -4566
rect 19108 -4630 19308 -4583
rect 15754 -4877 15954 -4830
rect 15754 -4894 15804 -4877
rect 15788 -4911 15804 -4894
rect 15904 -4894 15954 -4877
rect 16012 -4877 16212 -4830
rect 16012 -4894 16062 -4877
rect 15904 -4911 15920 -4894
rect 15788 -4927 15920 -4911
rect 16046 -4911 16062 -4894
rect 16162 -4894 16212 -4877
rect 16270 -4877 16470 -4830
rect 16270 -4894 16320 -4877
rect 16162 -4911 16178 -4894
rect 16046 -4927 16178 -4911
rect 16304 -4911 16320 -4894
rect 16420 -4894 16470 -4877
rect 16528 -4877 16728 -4830
rect 16528 -4894 16578 -4877
rect 16420 -4911 16436 -4894
rect 16304 -4927 16436 -4911
rect 16562 -4911 16578 -4894
rect 16678 -4894 16728 -4877
rect 16786 -4877 16986 -4830
rect 16786 -4894 16836 -4877
rect 16678 -4911 16694 -4894
rect 16562 -4927 16694 -4911
rect 16820 -4911 16836 -4894
rect 16936 -4894 16986 -4877
rect 17044 -4877 17244 -4830
rect 17044 -4894 17094 -4877
rect 16936 -4911 16952 -4894
rect 16820 -4927 16952 -4911
rect 17078 -4911 17094 -4894
rect 17194 -4894 17244 -4877
rect 17302 -4877 17502 -4830
rect 17302 -4894 17352 -4877
rect 17194 -4911 17210 -4894
rect 17078 -4927 17210 -4911
rect 17336 -4911 17352 -4894
rect 17452 -4894 17502 -4877
rect 17560 -4877 17760 -4830
rect 17560 -4894 17610 -4877
rect 17452 -4911 17468 -4894
rect 17336 -4927 17468 -4911
rect 17594 -4911 17610 -4894
rect 17710 -4894 17760 -4877
rect 17818 -4877 18018 -4830
rect 17818 -4894 17868 -4877
rect 17710 -4911 17726 -4894
rect 17594 -4927 17726 -4911
rect 17852 -4911 17868 -4894
rect 17968 -4894 18018 -4877
rect 18076 -4877 18276 -4830
rect 18076 -4894 18126 -4877
rect 17968 -4911 17984 -4894
rect 17852 -4927 17984 -4911
rect 18110 -4911 18126 -4894
rect 18226 -4894 18276 -4877
rect 18334 -4877 18534 -4830
rect 18334 -4894 18384 -4877
rect 18226 -4911 18242 -4894
rect 18110 -4927 18242 -4911
rect 18368 -4911 18384 -4894
rect 18484 -4894 18534 -4877
rect 18592 -4877 18792 -4830
rect 18592 -4894 18642 -4877
rect 18484 -4911 18500 -4894
rect 18368 -4927 18500 -4911
rect 18626 -4911 18642 -4894
rect 18742 -4894 18792 -4877
rect 18850 -4877 19050 -4830
rect 18850 -4894 18900 -4877
rect 18742 -4911 18758 -4894
rect 18626 -4927 18758 -4911
rect 18884 -4911 18900 -4894
rect 19000 -4894 19050 -4877
rect 19108 -4877 19308 -4830
rect 19108 -4894 19158 -4877
rect 19000 -4911 19016 -4894
rect 18884 -4927 19016 -4911
rect 19142 -4911 19158 -4894
rect 19258 -4894 19308 -4877
rect 19258 -4911 19274 -4894
rect 19142 -4927 19274 -4911
<< polycont >>
rect 4004 4073 4104 4107
rect 4262 4073 4362 4107
rect 4520 4073 4620 4107
rect 4778 4073 4878 4107
rect 5036 4073 5136 4107
rect 5294 4073 5394 4107
rect 5552 4073 5652 4107
rect 5810 4073 5910 4107
rect 6068 4073 6168 4107
rect 6326 4073 6426 4107
rect 6584 4073 6684 4107
rect 6842 4073 6942 4107
rect 7100 4073 7200 4107
rect 7358 4073 7458 4107
rect 4004 3745 4104 3779
rect 4262 3745 4362 3779
rect 4520 3745 4620 3779
rect 4778 3745 4878 3779
rect 5036 3745 5136 3779
rect 5294 3745 5394 3779
rect 5552 3745 5652 3779
rect 5810 3745 5910 3779
rect 6068 3745 6168 3779
rect 6326 3745 6426 3779
rect 6584 3745 6684 3779
rect 6842 3745 6942 3779
rect 7100 3745 7200 3779
rect 7358 3745 7458 3779
rect 15804 4073 15904 4107
rect 16062 4073 16162 4107
rect 16320 4073 16420 4107
rect 16578 4073 16678 4107
rect 16836 4073 16936 4107
rect 17094 4073 17194 4107
rect 17352 4073 17452 4107
rect 17610 4073 17710 4107
rect 17868 4073 17968 4107
rect 18126 4073 18226 4107
rect 18384 4073 18484 4107
rect 18642 4073 18742 4107
rect 18900 4073 19000 4107
rect 19158 4073 19258 4107
rect 15804 3745 15904 3779
rect 16062 3745 16162 3779
rect 16320 3745 16420 3779
rect 16578 3745 16678 3779
rect 16836 3745 16936 3779
rect 17094 3745 17194 3779
rect 17352 3745 17452 3779
rect 17610 3745 17710 3779
rect 17868 3745 17968 3779
rect 18126 3745 18226 3779
rect 18384 3745 18484 3779
rect 18642 3745 18742 3779
rect 18900 3745 19000 3779
rect 19158 3745 19258 3779
rect 1220 2596 1320 2630
rect 1478 2596 1578 2630
rect 1736 2596 1836 2630
rect 1994 2596 2094 2630
rect 2252 2596 2352 2630
rect 2510 2596 2610 2630
rect 2768 2596 2868 2630
rect 3026 2596 3126 2630
rect 3284 2596 3384 2630
rect 3542 2596 3642 2630
rect 4516 2596 4616 2630
rect 4774 2596 4874 2630
rect 5032 2596 5132 2630
rect 5290 2596 5390 2630
rect 5548 2596 5648 2630
rect 5806 2596 5906 2630
rect 6064 2596 6164 2630
rect 6322 2596 6422 2630
rect 6580 2596 6680 2630
rect 6838 2596 6938 2630
rect 7812 2596 7912 2630
rect 8070 2596 8170 2630
rect 8328 2596 8428 2630
rect 8586 2596 8686 2630
rect 8844 2596 8944 2630
rect 9102 2596 9202 2630
rect 9360 2596 9460 2630
rect 9618 2596 9718 2630
rect 9876 2596 9976 2630
rect 10134 2596 10234 2630
rect 1220 2086 1320 2120
rect 1478 2086 1578 2120
rect 1736 2086 1836 2120
rect 1994 2086 2094 2120
rect 2252 2086 2352 2120
rect 2510 2086 2610 2120
rect 2768 2086 2868 2120
rect 3026 2086 3126 2120
rect 3284 2086 3384 2120
rect 3542 2086 3642 2120
rect 4516 2086 4616 2120
rect 4774 2086 4874 2120
rect 5032 2086 5132 2120
rect 5290 2086 5390 2120
rect 5548 2086 5648 2120
rect 5806 2086 5906 2120
rect 6064 2086 6164 2120
rect 6322 2086 6422 2120
rect 6580 2086 6680 2120
rect 6838 2086 6938 2120
rect 7812 2086 7912 2120
rect 8070 2086 8170 2120
rect 8328 2086 8428 2120
rect 8586 2086 8686 2120
rect 8844 2086 8944 2120
rect 9102 2086 9202 2120
rect 9360 2086 9460 2120
rect 9618 2086 9718 2120
rect 9876 2086 9976 2120
rect 10134 2086 10234 2120
rect 792 1488 1252 1522
rect 1650 1488 2110 1522
rect 2508 1488 2968 1522
rect 3366 1488 3826 1522
rect 4224 1488 4684 1522
rect 5082 1488 5542 1522
rect 5940 1488 6400 1522
rect 6798 1488 7258 1522
rect 7656 1488 8116 1522
rect 8514 1488 8974 1522
rect 9372 1488 9832 1522
rect 10230 1488 10690 1522
rect 792 1178 1252 1212
rect 1650 1178 2110 1212
rect 2508 1178 2968 1212
rect 3366 1178 3826 1212
rect 4224 1178 4684 1212
rect 5082 1178 5542 1212
rect 5940 1178 6400 1212
rect 6798 1178 7258 1212
rect 7656 1178 8116 1212
rect 8514 1178 8974 1212
rect 9372 1178 9832 1212
rect 10230 1178 10690 1212
rect 792 948 1252 982
rect 1650 948 2110 982
rect 2508 948 2968 982
rect 3366 948 3826 982
rect 4224 948 4684 982
rect 5082 948 5542 982
rect 5940 948 6400 982
rect 6798 948 7258 982
rect 7656 948 8116 982
rect 8514 948 8974 982
rect 9372 948 9832 982
rect 10230 948 10690 982
rect 792 638 1252 672
rect 1650 638 2110 672
rect 2508 638 2968 672
rect 3366 638 3826 672
rect 4224 638 4684 672
rect 5082 638 5542 672
rect 5940 638 6400 672
rect 6798 638 7258 672
rect 7656 638 8116 672
rect 8514 638 8974 672
rect 9372 638 9832 672
rect 10230 638 10690 672
rect 13020 2596 13120 2630
rect 13278 2596 13378 2630
rect 13536 2596 13636 2630
rect 13794 2596 13894 2630
rect 14052 2596 14152 2630
rect 14310 2596 14410 2630
rect 14568 2596 14668 2630
rect 14826 2596 14926 2630
rect 15084 2596 15184 2630
rect 15342 2596 15442 2630
rect 16316 2596 16416 2630
rect 16574 2596 16674 2630
rect 16832 2596 16932 2630
rect 17090 2596 17190 2630
rect 17348 2596 17448 2630
rect 17606 2596 17706 2630
rect 17864 2596 17964 2630
rect 18122 2596 18222 2630
rect 18380 2596 18480 2630
rect 18638 2596 18738 2630
rect 19612 2596 19712 2630
rect 19870 2596 19970 2630
rect 20128 2596 20228 2630
rect 20386 2596 20486 2630
rect 20644 2596 20744 2630
rect 20902 2596 21002 2630
rect 21160 2596 21260 2630
rect 21418 2596 21518 2630
rect 21676 2596 21776 2630
rect 21934 2596 22034 2630
rect 13020 2086 13120 2120
rect 13278 2086 13378 2120
rect 13536 2086 13636 2120
rect 13794 2086 13894 2120
rect 14052 2086 14152 2120
rect 14310 2086 14410 2120
rect 14568 2086 14668 2120
rect 14826 2086 14926 2120
rect 15084 2086 15184 2120
rect 15342 2086 15442 2120
rect 16316 2086 16416 2120
rect 16574 2086 16674 2120
rect 16832 2086 16932 2120
rect 17090 2086 17190 2120
rect 17348 2086 17448 2120
rect 17606 2086 17706 2120
rect 17864 2086 17964 2120
rect 18122 2086 18222 2120
rect 18380 2086 18480 2120
rect 18638 2086 18738 2120
rect 19612 2086 19712 2120
rect 19870 2086 19970 2120
rect 20128 2086 20228 2120
rect 20386 2086 20486 2120
rect 20644 2086 20744 2120
rect 20902 2086 21002 2120
rect 21160 2086 21260 2120
rect 21418 2086 21518 2120
rect 21676 2086 21776 2120
rect 21934 2086 22034 2120
rect 12592 1488 13052 1522
rect 13450 1488 13910 1522
rect 14308 1488 14768 1522
rect 15166 1488 15626 1522
rect 16024 1488 16484 1522
rect 16882 1488 17342 1522
rect 17740 1488 18200 1522
rect 18598 1488 19058 1522
rect 19456 1488 19916 1522
rect 20314 1488 20774 1522
rect 21172 1488 21632 1522
rect 22030 1488 22490 1522
rect 12592 1178 13052 1212
rect 13450 1178 13910 1212
rect 14308 1178 14768 1212
rect 15166 1178 15626 1212
rect 16024 1178 16484 1212
rect 16882 1178 17342 1212
rect 17740 1178 18200 1212
rect 18598 1178 19058 1212
rect 19456 1178 19916 1212
rect 20314 1178 20774 1212
rect 21172 1178 21632 1212
rect 22030 1178 22490 1212
rect 12592 948 13052 982
rect 13450 948 13910 982
rect 14308 948 14768 982
rect 15166 948 15626 982
rect 16024 948 16484 982
rect 16882 948 17342 982
rect 17740 948 18200 982
rect 18598 948 19058 982
rect 19456 948 19916 982
rect 20314 948 20774 982
rect 21172 948 21632 982
rect 22030 948 22490 982
rect 12592 638 13052 672
rect 13450 638 13910 672
rect 14308 638 14768 672
rect 15166 638 15626 672
rect 16024 638 16484 672
rect 16882 638 17342 672
rect 17740 638 18200 672
rect 18598 638 19058 672
rect 19456 638 19916 672
rect 20314 638 20774 672
rect 21172 638 21632 672
rect 22030 638 22490 672
rect 792 -1476 1252 -1442
rect 1650 -1476 2110 -1442
rect 2508 -1476 2968 -1442
rect 3366 -1476 3826 -1442
rect 4224 -1476 4684 -1442
rect 5082 -1476 5542 -1442
rect 5940 -1476 6400 -1442
rect 6798 -1476 7258 -1442
rect 7656 -1476 8116 -1442
rect 8514 -1476 8974 -1442
rect 9372 -1476 9832 -1442
rect 10230 -1476 10690 -1442
rect 792 -1786 1252 -1752
rect 1650 -1786 2110 -1752
rect 2508 -1786 2968 -1752
rect 3366 -1786 3826 -1752
rect 4224 -1786 4684 -1752
rect 5082 -1786 5542 -1752
rect 5940 -1786 6400 -1752
rect 6798 -1786 7258 -1752
rect 7656 -1786 8116 -1752
rect 8514 -1786 8974 -1752
rect 9372 -1786 9832 -1752
rect 10230 -1786 10690 -1752
rect 792 -2016 1252 -1982
rect 1650 -2016 2110 -1982
rect 2508 -2016 2968 -1982
rect 3366 -2016 3826 -1982
rect 4224 -2016 4684 -1982
rect 5082 -2016 5542 -1982
rect 5940 -2016 6400 -1982
rect 6798 -2016 7258 -1982
rect 7656 -2016 8116 -1982
rect 8514 -2016 8974 -1982
rect 9372 -2016 9832 -1982
rect 10230 -2016 10690 -1982
rect 792 -2326 1252 -2292
rect 1650 -2326 2110 -2292
rect 2508 -2326 2968 -2292
rect 3366 -2326 3826 -2292
rect 4224 -2326 4684 -2292
rect 5082 -2326 5542 -2292
rect 5940 -2326 6400 -2292
rect 6798 -2326 7258 -2292
rect 7656 -2326 8116 -2292
rect 8514 -2326 8974 -2292
rect 9372 -2326 9832 -2292
rect 10230 -2326 10690 -2292
rect 1220 -2924 1320 -2890
rect 1478 -2924 1578 -2890
rect 1736 -2924 1836 -2890
rect 1994 -2924 2094 -2890
rect 2252 -2924 2352 -2890
rect 2510 -2924 2610 -2890
rect 2768 -2924 2868 -2890
rect 3026 -2924 3126 -2890
rect 3284 -2924 3384 -2890
rect 3542 -2924 3642 -2890
rect 4516 -2924 4616 -2890
rect 4774 -2924 4874 -2890
rect 5032 -2924 5132 -2890
rect 5290 -2924 5390 -2890
rect 5548 -2924 5648 -2890
rect 5806 -2924 5906 -2890
rect 6064 -2924 6164 -2890
rect 6322 -2924 6422 -2890
rect 6580 -2924 6680 -2890
rect 6838 -2924 6938 -2890
rect 7812 -2924 7912 -2890
rect 8070 -2924 8170 -2890
rect 8328 -2924 8428 -2890
rect 8586 -2924 8686 -2890
rect 8844 -2924 8944 -2890
rect 9102 -2924 9202 -2890
rect 9360 -2924 9460 -2890
rect 9618 -2924 9718 -2890
rect 9876 -2924 9976 -2890
rect 10134 -2924 10234 -2890
rect 1220 -3434 1320 -3400
rect 1478 -3434 1578 -3400
rect 1736 -3434 1836 -3400
rect 1994 -3434 2094 -3400
rect 2252 -3434 2352 -3400
rect 2510 -3434 2610 -3400
rect 2768 -3434 2868 -3400
rect 3026 -3434 3126 -3400
rect 3284 -3434 3384 -3400
rect 3542 -3434 3642 -3400
rect 4516 -3434 4616 -3400
rect 4774 -3434 4874 -3400
rect 5032 -3434 5132 -3400
rect 5290 -3434 5390 -3400
rect 5548 -3434 5648 -3400
rect 5806 -3434 5906 -3400
rect 6064 -3434 6164 -3400
rect 6322 -3434 6422 -3400
rect 6580 -3434 6680 -3400
rect 6838 -3434 6938 -3400
rect 7812 -3434 7912 -3400
rect 8070 -3434 8170 -3400
rect 8328 -3434 8428 -3400
rect 8586 -3434 8686 -3400
rect 8844 -3434 8944 -3400
rect 9102 -3434 9202 -3400
rect 9360 -3434 9460 -3400
rect 9618 -3434 9718 -3400
rect 9876 -3434 9976 -3400
rect 10134 -3434 10234 -3400
rect 12592 -1476 13052 -1442
rect 13450 -1476 13910 -1442
rect 14308 -1476 14768 -1442
rect 15166 -1476 15626 -1442
rect 16024 -1476 16484 -1442
rect 16882 -1476 17342 -1442
rect 17740 -1476 18200 -1442
rect 18598 -1476 19058 -1442
rect 19456 -1476 19916 -1442
rect 20314 -1476 20774 -1442
rect 21172 -1476 21632 -1442
rect 22030 -1476 22490 -1442
rect 12592 -1786 13052 -1752
rect 13450 -1786 13910 -1752
rect 14308 -1786 14768 -1752
rect 15166 -1786 15626 -1752
rect 16024 -1786 16484 -1752
rect 16882 -1786 17342 -1752
rect 17740 -1786 18200 -1752
rect 18598 -1786 19058 -1752
rect 19456 -1786 19916 -1752
rect 20314 -1786 20774 -1752
rect 21172 -1786 21632 -1752
rect 22030 -1786 22490 -1752
rect 12592 -2016 13052 -1982
rect 13450 -2016 13910 -1982
rect 14308 -2016 14768 -1982
rect 15166 -2016 15626 -1982
rect 16024 -2016 16484 -1982
rect 16882 -2016 17342 -1982
rect 17740 -2016 18200 -1982
rect 18598 -2016 19058 -1982
rect 19456 -2016 19916 -1982
rect 20314 -2016 20774 -1982
rect 21172 -2016 21632 -1982
rect 22030 -2016 22490 -1982
rect 12592 -2326 13052 -2292
rect 13450 -2326 13910 -2292
rect 14308 -2326 14768 -2292
rect 15166 -2326 15626 -2292
rect 16024 -2326 16484 -2292
rect 16882 -2326 17342 -2292
rect 17740 -2326 18200 -2292
rect 18598 -2326 19058 -2292
rect 19456 -2326 19916 -2292
rect 20314 -2326 20774 -2292
rect 21172 -2326 21632 -2292
rect 22030 -2326 22490 -2292
rect 13020 -2924 13120 -2890
rect 13278 -2924 13378 -2890
rect 13536 -2924 13636 -2890
rect 13794 -2924 13894 -2890
rect 14052 -2924 14152 -2890
rect 14310 -2924 14410 -2890
rect 14568 -2924 14668 -2890
rect 14826 -2924 14926 -2890
rect 15084 -2924 15184 -2890
rect 15342 -2924 15442 -2890
rect 16316 -2924 16416 -2890
rect 16574 -2924 16674 -2890
rect 16832 -2924 16932 -2890
rect 17090 -2924 17190 -2890
rect 17348 -2924 17448 -2890
rect 17606 -2924 17706 -2890
rect 17864 -2924 17964 -2890
rect 18122 -2924 18222 -2890
rect 18380 -2924 18480 -2890
rect 18638 -2924 18738 -2890
rect 19612 -2924 19712 -2890
rect 19870 -2924 19970 -2890
rect 20128 -2924 20228 -2890
rect 20386 -2924 20486 -2890
rect 20644 -2924 20744 -2890
rect 20902 -2924 21002 -2890
rect 21160 -2924 21260 -2890
rect 21418 -2924 21518 -2890
rect 21676 -2924 21776 -2890
rect 21934 -2924 22034 -2890
rect 13020 -3434 13120 -3400
rect 13278 -3434 13378 -3400
rect 13536 -3434 13636 -3400
rect 13794 -3434 13894 -3400
rect 14052 -3434 14152 -3400
rect 14310 -3434 14410 -3400
rect 14568 -3434 14668 -3400
rect 14826 -3434 14926 -3400
rect 15084 -3434 15184 -3400
rect 15342 -3434 15442 -3400
rect 16316 -3434 16416 -3400
rect 16574 -3434 16674 -3400
rect 16832 -3434 16932 -3400
rect 17090 -3434 17190 -3400
rect 17348 -3434 17448 -3400
rect 17606 -3434 17706 -3400
rect 17864 -3434 17964 -3400
rect 18122 -3434 18222 -3400
rect 18380 -3434 18480 -3400
rect 18638 -3434 18738 -3400
rect 19612 -3434 19712 -3400
rect 19870 -3434 19970 -3400
rect 20128 -3434 20228 -3400
rect 20386 -3434 20486 -3400
rect 20644 -3434 20744 -3400
rect 20902 -3434 21002 -3400
rect 21160 -3434 21260 -3400
rect 21418 -3434 21518 -3400
rect 21676 -3434 21776 -3400
rect 21934 -3434 22034 -3400
rect 4004 -4583 4104 -4549
rect 4262 -4583 4362 -4549
rect 4520 -4583 4620 -4549
rect 4778 -4583 4878 -4549
rect 5036 -4583 5136 -4549
rect 5294 -4583 5394 -4549
rect 5552 -4583 5652 -4549
rect 5810 -4583 5910 -4549
rect 6068 -4583 6168 -4549
rect 6326 -4583 6426 -4549
rect 6584 -4583 6684 -4549
rect 6842 -4583 6942 -4549
rect 7100 -4583 7200 -4549
rect 7358 -4583 7458 -4549
rect 4004 -4911 4104 -4877
rect 4262 -4911 4362 -4877
rect 4520 -4911 4620 -4877
rect 4778 -4911 4878 -4877
rect 5036 -4911 5136 -4877
rect 5294 -4911 5394 -4877
rect 5552 -4911 5652 -4877
rect 5810 -4911 5910 -4877
rect 6068 -4911 6168 -4877
rect 6326 -4911 6426 -4877
rect 6584 -4911 6684 -4877
rect 6842 -4911 6942 -4877
rect 7100 -4911 7200 -4877
rect 7358 -4911 7458 -4877
rect 15804 -4583 15904 -4549
rect 16062 -4583 16162 -4549
rect 16320 -4583 16420 -4549
rect 16578 -4583 16678 -4549
rect 16836 -4583 16936 -4549
rect 17094 -4583 17194 -4549
rect 17352 -4583 17452 -4549
rect 17610 -4583 17710 -4549
rect 17868 -4583 17968 -4549
rect 18126 -4583 18226 -4549
rect 18384 -4583 18484 -4549
rect 18642 -4583 18742 -4549
rect 18900 -4583 19000 -4549
rect 19158 -4583 19258 -4549
rect 15804 -4911 15904 -4877
rect 16062 -4911 16162 -4877
rect 16320 -4911 16420 -4877
rect 16578 -4911 16678 -4877
rect 16836 -4911 16936 -4877
rect 17094 -4911 17194 -4877
rect 17352 -4911 17452 -4877
rect 17610 -4911 17710 -4877
rect 17868 -4911 17968 -4877
rect 18126 -4911 18226 -4877
rect 18384 -4911 18484 -4877
rect 18642 -4911 18742 -4877
rect 18900 -4911 19000 -4877
rect 19158 -4911 19258 -4877
<< locali >>
rect 66 4978 166 5138
rect 11310 4978 11410 5138
rect 3988 4073 4004 4107
rect 4104 4073 4120 4107
rect 4246 4073 4262 4107
rect 4362 4073 4378 4107
rect 4504 4073 4520 4107
rect 4620 4073 4636 4107
rect 4762 4073 4778 4107
rect 4878 4073 4894 4107
rect 5020 4073 5036 4107
rect 5136 4073 5152 4107
rect 5278 4073 5294 4107
rect 5394 4073 5410 4107
rect 5536 4073 5552 4107
rect 5652 4073 5668 4107
rect 5794 4073 5810 4107
rect 5910 4073 5926 4107
rect 6052 4073 6068 4107
rect 6168 4073 6184 4107
rect 6310 4073 6326 4107
rect 6426 4073 6442 4107
rect 6568 4073 6584 4107
rect 6684 4073 6700 4107
rect 6826 4073 6842 4107
rect 6942 4073 6958 4107
rect 7084 4073 7100 4107
rect 7200 4073 7216 4107
rect 7342 4073 7358 4107
rect 7458 4073 7474 4107
rect 3908 4014 3942 4030
rect 3908 3822 3942 3838
rect 4166 4014 4200 4030
rect 4166 3822 4200 3838
rect 4424 4014 4458 4030
rect 4424 3822 4458 3838
rect 4682 4014 4716 4030
rect 4682 3822 4716 3838
rect 4940 4014 4974 4030
rect 4940 3822 4974 3838
rect 5198 4014 5232 4030
rect 5198 3822 5232 3838
rect 5456 4014 5490 4030
rect 5456 3822 5490 3838
rect 5714 4014 5748 4030
rect 5714 3822 5748 3838
rect 5972 4014 6006 4030
rect 5972 3822 6006 3838
rect 6230 4014 6264 4030
rect 6230 3822 6264 3838
rect 6488 4014 6522 4030
rect 6488 3822 6522 3838
rect 6746 4014 6780 4030
rect 6746 3822 6780 3838
rect 7004 4014 7038 4030
rect 7004 3822 7038 3838
rect 7262 4014 7296 4030
rect 7262 3822 7296 3838
rect 7520 4014 7554 4030
rect 7520 3822 7554 3838
rect 3988 3745 4004 3779
rect 4104 3745 4120 3779
rect 4246 3745 4262 3779
rect 4362 3745 4378 3779
rect 4504 3745 4520 3779
rect 4620 3745 4636 3779
rect 4762 3745 4778 3779
rect 4878 3745 4894 3779
rect 5020 3745 5036 3779
rect 5136 3745 5152 3779
rect 5278 3745 5294 3779
rect 5394 3745 5410 3779
rect 5536 3745 5552 3779
rect 5652 3745 5668 3779
rect 5794 3745 5810 3779
rect 5910 3745 5926 3779
rect 6052 3745 6068 3779
rect 6168 3745 6184 3779
rect 6310 3745 6326 3779
rect 6426 3745 6442 3779
rect 6568 3745 6584 3779
rect 6684 3745 6700 3779
rect 6826 3745 6842 3779
rect 6942 3745 6958 3779
rect 7084 3745 7100 3779
rect 7200 3745 7216 3779
rect 7342 3745 7358 3779
rect 7458 3745 7474 3779
rect 66 3354 166 3514
rect 11310 3354 11410 3514
rect 11866 4978 11966 5138
rect 23110 4978 23210 5138
rect 15788 4073 15804 4107
rect 15904 4073 15920 4107
rect 16046 4073 16062 4107
rect 16162 4073 16178 4107
rect 16304 4073 16320 4107
rect 16420 4073 16436 4107
rect 16562 4073 16578 4107
rect 16678 4073 16694 4107
rect 16820 4073 16836 4107
rect 16936 4073 16952 4107
rect 17078 4073 17094 4107
rect 17194 4073 17210 4107
rect 17336 4073 17352 4107
rect 17452 4073 17468 4107
rect 17594 4073 17610 4107
rect 17710 4073 17726 4107
rect 17852 4073 17868 4107
rect 17968 4073 17984 4107
rect 18110 4073 18126 4107
rect 18226 4073 18242 4107
rect 18368 4073 18384 4107
rect 18484 4073 18500 4107
rect 18626 4073 18642 4107
rect 18742 4073 18758 4107
rect 18884 4073 18900 4107
rect 19000 4073 19016 4107
rect 19142 4073 19158 4107
rect 19258 4073 19274 4107
rect 15708 4014 15742 4030
rect 15708 3822 15742 3838
rect 15966 4014 16000 4030
rect 15966 3822 16000 3838
rect 16224 4014 16258 4030
rect 16224 3822 16258 3838
rect 16482 4014 16516 4030
rect 16482 3822 16516 3838
rect 16740 4014 16774 4030
rect 16740 3822 16774 3838
rect 16998 4014 17032 4030
rect 16998 3822 17032 3838
rect 17256 4014 17290 4030
rect 17256 3822 17290 3838
rect 17514 4014 17548 4030
rect 17514 3822 17548 3838
rect 17772 4014 17806 4030
rect 17772 3822 17806 3838
rect 18030 4014 18064 4030
rect 18030 3822 18064 3838
rect 18288 4014 18322 4030
rect 18288 3822 18322 3838
rect 18546 4014 18580 4030
rect 18546 3822 18580 3838
rect 18804 4014 18838 4030
rect 18804 3822 18838 3838
rect 19062 4014 19096 4030
rect 19062 3822 19096 3838
rect 19320 4014 19354 4030
rect 19320 3822 19354 3838
rect 15788 3745 15804 3779
rect 15904 3745 15920 3779
rect 16046 3745 16062 3779
rect 16162 3745 16178 3779
rect 16304 3745 16320 3779
rect 16420 3745 16436 3779
rect 16562 3745 16578 3779
rect 16678 3745 16694 3779
rect 16820 3745 16836 3779
rect 16936 3745 16952 3779
rect 17078 3745 17094 3779
rect 17194 3745 17210 3779
rect 17336 3745 17352 3779
rect 17452 3745 17468 3779
rect 17594 3745 17610 3779
rect 17710 3745 17726 3779
rect 17852 3745 17868 3779
rect 17968 3745 17984 3779
rect 18110 3745 18126 3779
rect 18226 3745 18242 3779
rect 18368 3745 18384 3779
rect 18484 3745 18500 3779
rect 18626 3745 18642 3779
rect 18742 3745 18758 3779
rect 18884 3745 18900 3779
rect 19000 3745 19016 3779
rect 19142 3745 19158 3779
rect 19258 3745 19274 3779
rect 11866 3354 11966 3514
rect 23110 3354 23210 3514
rect 66 2956 166 3118
rect 11310 2956 11410 3118
rect 1204 2596 1220 2630
rect 1320 2596 1336 2630
rect 1462 2596 1478 2630
rect 1578 2596 1594 2630
rect 1720 2596 1736 2630
rect 1836 2596 1852 2630
rect 1978 2596 1994 2630
rect 2094 2596 2110 2630
rect 2236 2596 2252 2630
rect 2352 2596 2368 2630
rect 2494 2596 2510 2630
rect 2610 2596 2626 2630
rect 2752 2596 2768 2630
rect 2868 2596 2884 2630
rect 3010 2596 3026 2630
rect 3126 2596 3142 2630
rect 3268 2596 3284 2630
rect 3384 2596 3400 2630
rect 3526 2596 3542 2630
rect 3642 2596 3658 2630
rect 4500 2596 4516 2630
rect 4616 2596 4632 2630
rect 4758 2596 4774 2630
rect 4874 2596 4890 2630
rect 5016 2596 5032 2630
rect 5132 2596 5148 2630
rect 5274 2596 5290 2630
rect 5390 2596 5406 2630
rect 5532 2596 5548 2630
rect 5648 2596 5664 2630
rect 5790 2596 5806 2630
rect 5906 2596 5922 2630
rect 6048 2596 6064 2630
rect 6164 2596 6180 2630
rect 6306 2596 6322 2630
rect 6422 2596 6438 2630
rect 6564 2596 6580 2630
rect 6680 2596 6696 2630
rect 6822 2596 6838 2630
rect 6938 2596 6954 2630
rect 7796 2596 7812 2630
rect 7912 2596 7928 2630
rect 8054 2596 8070 2630
rect 8170 2596 8186 2630
rect 8312 2596 8328 2630
rect 8428 2596 8444 2630
rect 8570 2596 8586 2630
rect 8686 2596 8702 2630
rect 8828 2596 8844 2630
rect 8944 2596 8960 2630
rect 9086 2596 9102 2630
rect 9202 2596 9218 2630
rect 9344 2596 9360 2630
rect 9460 2596 9476 2630
rect 9602 2596 9618 2630
rect 9718 2596 9734 2630
rect 9860 2596 9876 2630
rect 9976 2596 9992 2630
rect 10118 2596 10134 2630
rect 10234 2596 10250 2630
rect 1124 2546 1158 2562
rect 1124 2154 1158 2170
rect 1382 2546 1416 2562
rect 1382 2154 1416 2170
rect 1640 2546 1674 2562
rect 1640 2154 1674 2170
rect 1898 2546 1932 2562
rect 1898 2154 1932 2170
rect 2156 2546 2190 2562
rect 2156 2154 2190 2170
rect 2414 2546 2448 2562
rect 2414 2154 2448 2170
rect 2672 2546 2706 2562
rect 2672 2154 2706 2170
rect 2930 2546 2964 2562
rect 2930 2154 2964 2170
rect 3188 2546 3222 2562
rect 3188 2154 3222 2170
rect 3446 2546 3480 2562
rect 3446 2154 3480 2170
rect 3704 2546 3738 2562
rect 3704 2154 3738 2170
rect 4420 2546 4454 2562
rect 4420 2154 4454 2170
rect 4678 2546 4712 2562
rect 4678 2154 4712 2170
rect 4936 2546 4970 2562
rect 4936 2154 4970 2170
rect 5194 2546 5228 2562
rect 5194 2154 5228 2170
rect 5452 2546 5486 2562
rect 5452 2154 5486 2170
rect 5710 2546 5744 2562
rect 5710 2154 5744 2170
rect 5968 2546 6002 2562
rect 5968 2154 6002 2170
rect 6226 2546 6260 2562
rect 6226 2154 6260 2170
rect 6484 2546 6518 2562
rect 6484 2154 6518 2170
rect 6742 2546 6776 2562
rect 6742 2154 6776 2170
rect 7000 2546 7034 2562
rect 7000 2154 7034 2170
rect 7716 2546 7750 2562
rect 7716 2154 7750 2170
rect 7974 2546 8008 2562
rect 7974 2154 8008 2170
rect 8232 2546 8266 2562
rect 8232 2154 8266 2170
rect 8490 2546 8524 2562
rect 8490 2154 8524 2170
rect 8748 2546 8782 2562
rect 8748 2154 8782 2170
rect 9006 2546 9040 2562
rect 9006 2154 9040 2170
rect 9264 2546 9298 2562
rect 9264 2154 9298 2170
rect 9522 2546 9556 2562
rect 9522 2154 9556 2170
rect 9780 2546 9814 2562
rect 9780 2154 9814 2170
rect 10038 2546 10072 2562
rect 10038 2154 10072 2170
rect 10296 2546 10330 2562
rect 10296 2154 10330 2170
rect 1204 2086 1220 2120
rect 1320 2086 1336 2120
rect 1462 2086 1478 2120
rect 1578 2086 1594 2120
rect 1720 2086 1736 2120
rect 1836 2086 1852 2120
rect 1978 2086 1994 2120
rect 2094 2086 2110 2120
rect 2236 2086 2252 2120
rect 2352 2086 2368 2120
rect 2494 2086 2510 2120
rect 2610 2086 2626 2120
rect 2752 2086 2768 2120
rect 2868 2086 2884 2120
rect 3010 2086 3026 2120
rect 3126 2086 3142 2120
rect 3268 2086 3284 2120
rect 3384 2086 3400 2120
rect 3526 2086 3542 2120
rect 3642 2086 3658 2120
rect 4500 2086 4516 2120
rect 4616 2086 4632 2120
rect 4758 2086 4774 2120
rect 4874 2086 4890 2120
rect 5016 2086 5032 2120
rect 5132 2086 5148 2120
rect 5274 2086 5290 2120
rect 5390 2086 5406 2120
rect 5532 2086 5548 2120
rect 5648 2086 5664 2120
rect 5790 2086 5806 2120
rect 5906 2086 5922 2120
rect 6048 2086 6064 2120
rect 6164 2086 6180 2120
rect 6306 2086 6322 2120
rect 6422 2086 6438 2120
rect 6564 2086 6580 2120
rect 6680 2086 6696 2120
rect 6822 2086 6838 2120
rect 6938 2086 6954 2120
rect 7796 2086 7812 2120
rect 7912 2086 7928 2120
rect 8054 2086 8070 2120
rect 8170 2086 8186 2120
rect 8312 2086 8328 2120
rect 8428 2086 8444 2120
rect 8570 2086 8586 2120
rect 8686 2086 8702 2120
rect 8828 2086 8844 2120
rect 8944 2086 8960 2120
rect 9086 2086 9102 2120
rect 9202 2086 9218 2120
rect 9344 2086 9360 2120
rect 9460 2086 9476 2120
rect 9602 2086 9618 2120
rect 9718 2086 9734 2120
rect 9860 2086 9876 2120
rect 9976 2086 9992 2120
rect 10118 2086 10134 2120
rect 10234 2086 10250 2120
rect 776 1488 792 1522
rect 1252 1488 1268 1522
rect 1634 1488 1650 1522
rect 2110 1488 2126 1522
rect 2492 1488 2508 1522
rect 2968 1488 2984 1522
rect 3350 1488 3366 1522
rect 3826 1488 3842 1522
rect 4208 1488 4224 1522
rect 4684 1488 4700 1522
rect 5066 1488 5082 1522
rect 5542 1488 5558 1522
rect 5924 1488 5940 1522
rect 6400 1488 6416 1522
rect 6782 1488 6798 1522
rect 7258 1488 7274 1522
rect 7640 1488 7656 1522
rect 8116 1488 8132 1522
rect 8498 1488 8514 1522
rect 8974 1488 8990 1522
rect 9356 1488 9372 1522
rect 9832 1488 9848 1522
rect 10214 1488 10230 1522
rect 10690 1488 10706 1522
rect 576 1438 610 1454
rect 576 1246 610 1262
rect 1434 1438 1468 1454
rect 1434 1246 1468 1262
rect 2292 1438 2326 1454
rect 2292 1246 2326 1262
rect 3150 1438 3184 1454
rect 3150 1246 3184 1262
rect 4008 1438 4042 1454
rect 4008 1246 4042 1262
rect 4866 1438 4900 1454
rect 4866 1246 4900 1262
rect 5724 1438 5758 1454
rect 5724 1246 5758 1262
rect 6582 1438 6616 1454
rect 6582 1246 6616 1262
rect 7440 1438 7474 1454
rect 7440 1246 7474 1262
rect 8298 1438 8332 1454
rect 8298 1246 8332 1262
rect 9156 1438 9190 1454
rect 9156 1246 9190 1262
rect 10014 1438 10048 1454
rect 10014 1246 10048 1262
rect 10872 1438 10906 1454
rect 10872 1246 10906 1262
rect 776 1178 792 1212
rect 1252 1178 1268 1212
rect 1634 1178 1650 1212
rect 2110 1178 2126 1212
rect 2492 1178 2508 1212
rect 2968 1178 2984 1212
rect 3350 1178 3366 1212
rect 3826 1178 3842 1212
rect 4208 1178 4224 1212
rect 4684 1178 4700 1212
rect 5066 1178 5082 1212
rect 5542 1178 5558 1212
rect 5924 1178 5940 1212
rect 6400 1178 6416 1212
rect 6782 1178 6798 1212
rect 7258 1178 7274 1212
rect 7640 1178 7656 1212
rect 8116 1178 8132 1212
rect 8498 1178 8514 1212
rect 8974 1178 8990 1212
rect 9356 1178 9372 1212
rect 9832 1178 9848 1212
rect 10214 1178 10230 1212
rect 10690 1178 10706 1212
rect 776 948 792 982
rect 1252 948 1268 982
rect 1634 948 1650 982
rect 2110 948 2126 982
rect 2492 948 2508 982
rect 2968 948 2984 982
rect 3350 948 3366 982
rect 3826 948 3842 982
rect 4208 948 4224 982
rect 4684 948 4700 982
rect 5066 948 5082 982
rect 5542 948 5558 982
rect 5924 948 5940 982
rect 6400 948 6416 982
rect 6782 948 6798 982
rect 7258 948 7274 982
rect 7640 948 7656 982
rect 8116 948 8132 982
rect 8498 948 8514 982
rect 8974 948 8990 982
rect 9356 948 9372 982
rect 9832 948 9848 982
rect 10214 948 10230 982
rect 10690 948 10706 982
rect 576 898 610 914
rect 576 706 610 722
rect 1434 898 1468 914
rect 1434 706 1468 722
rect 2292 898 2326 914
rect 2292 706 2326 722
rect 3150 898 3184 914
rect 3150 706 3184 722
rect 4008 898 4042 914
rect 4008 706 4042 722
rect 4866 898 4900 914
rect 4866 706 4900 722
rect 5724 898 5758 914
rect 5724 706 5758 722
rect 6582 898 6616 914
rect 6582 706 6616 722
rect 7440 898 7474 914
rect 7440 706 7474 722
rect 8298 898 8332 914
rect 8298 706 8332 722
rect 9156 898 9190 914
rect 9156 706 9190 722
rect 10014 898 10048 914
rect 10014 706 10048 722
rect 10872 898 10906 914
rect 10872 706 10906 722
rect 776 638 792 672
rect 1252 638 1268 672
rect 1634 638 1650 672
rect 2110 638 2126 672
rect 2492 638 2508 672
rect 2968 638 2984 672
rect 3350 638 3366 672
rect 3826 638 3842 672
rect 4208 638 4224 672
rect 4684 638 4700 672
rect 5066 638 5082 672
rect 5542 638 5558 672
rect 5924 638 5940 672
rect 6400 638 6416 672
rect 6782 638 6798 672
rect 7258 638 7274 672
rect 7640 638 7656 672
rect 8116 638 8132 672
rect 8498 638 8514 672
rect 8974 638 8990 672
rect 9356 638 9372 672
rect 9832 638 9848 672
rect 10214 638 10230 672
rect 10690 638 10706 672
rect 66 -286 166 -124
rect 11310 -286 11410 -124
rect 11866 2956 11966 3118
rect 23110 2956 23210 3118
rect 13004 2596 13020 2630
rect 13120 2596 13136 2630
rect 13262 2596 13278 2630
rect 13378 2596 13394 2630
rect 13520 2596 13536 2630
rect 13636 2596 13652 2630
rect 13778 2596 13794 2630
rect 13894 2596 13910 2630
rect 14036 2596 14052 2630
rect 14152 2596 14168 2630
rect 14294 2596 14310 2630
rect 14410 2596 14426 2630
rect 14552 2596 14568 2630
rect 14668 2596 14684 2630
rect 14810 2596 14826 2630
rect 14926 2596 14942 2630
rect 15068 2596 15084 2630
rect 15184 2596 15200 2630
rect 15326 2596 15342 2630
rect 15442 2596 15458 2630
rect 16300 2596 16316 2630
rect 16416 2596 16432 2630
rect 16558 2596 16574 2630
rect 16674 2596 16690 2630
rect 16816 2596 16832 2630
rect 16932 2596 16948 2630
rect 17074 2596 17090 2630
rect 17190 2596 17206 2630
rect 17332 2596 17348 2630
rect 17448 2596 17464 2630
rect 17590 2596 17606 2630
rect 17706 2596 17722 2630
rect 17848 2596 17864 2630
rect 17964 2596 17980 2630
rect 18106 2596 18122 2630
rect 18222 2596 18238 2630
rect 18364 2596 18380 2630
rect 18480 2596 18496 2630
rect 18622 2596 18638 2630
rect 18738 2596 18754 2630
rect 19596 2596 19612 2630
rect 19712 2596 19728 2630
rect 19854 2596 19870 2630
rect 19970 2596 19986 2630
rect 20112 2596 20128 2630
rect 20228 2596 20244 2630
rect 20370 2596 20386 2630
rect 20486 2596 20502 2630
rect 20628 2596 20644 2630
rect 20744 2596 20760 2630
rect 20886 2596 20902 2630
rect 21002 2596 21018 2630
rect 21144 2596 21160 2630
rect 21260 2596 21276 2630
rect 21402 2596 21418 2630
rect 21518 2596 21534 2630
rect 21660 2596 21676 2630
rect 21776 2596 21792 2630
rect 21918 2596 21934 2630
rect 22034 2596 22050 2630
rect 12924 2546 12958 2562
rect 12924 2154 12958 2170
rect 13182 2546 13216 2562
rect 13182 2154 13216 2170
rect 13440 2546 13474 2562
rect 13440 2154 13474 2170
rect 13698 2546 13732 2562
rect 13698 2154 13732 2170
rect 13956 2546 13990 2562
rect 13956 2154 13990 2170
rect 14214 2546 14248 2562
rect 14214 2154 14248 2170
rect 14472 2546 14506 2562
rect 14472 2154 14506 2170
rect 14730 2546 14764 2562
rect 14730 2154 14764 2170
rect 14988 2546 15022 2562
rect 14988 2154 15022 2170
rect 15246 2546 15280 2562
rect 15246 2154 15280 2170
rect 15504 2546 15538 2562
rect 15504 2154 15538 2170
rect 16220 2546 16254 2562
rect 16220 2154 16254 2170
rect 16478 2546 16512 2562
rect 16478 2154 16512 2170
rect 16736 2546 16770 2562
rect 16736 2154 16770 2170
rect 16994 2546 17028 2562
rect 16994 2154 17028 2170
rect 17252 2546 17286 2562
rect 17252 2154 17286 2170
rect 17510 2546 17544 2562
rect 17510 2154 17544 2170
rect 17768 2546 17802 2562
rect 17768 2154 17802 2170
rect 18026 2546 18060 2562
rect 18026 2154 18060 2170
rect 18284 2546 18318 2562
rect 18284 2154 18318 2170
rect 18542 2546 18576 2562
rect 18542 2154 18576 2170
rect 18800 2546 18834 2562
rect 18800 2154 18834 2170
rect 19516 2546 19550 2562
rect 19516 2154 19550 2170
rect 19774 2546 19808 2562
rect 19774 2154 19808 2170
rect 20032 2546 20066 2562
rect 20032 2154 20066 2170
rect 20290 2546 20324 2562
rect 20290 2154 20324 2170
rect 20548 2546 20582 2562
rect 20548 2154 20582 2170
rect 20806 2546 20840 2562
rect 20806 2154 20840 2170
rect 21064 2546 21098 2562
rect 21064 2154 21098 2170
rect 21322 2546 21356 2562
rect 21322 2154 21356 2170
rect 21580 2546 21614 2562
rect 21580 2154 21614 2170
rect 21838 2546 21872 2562
rect 21838 2154 21872 2170
rect 22096 2546 22130 2562
rect 22096 2154 22130 2170
rect 13004 2086 13020 2120
rect 13120 2086 13136 2120
rect 13262 2086 13278 2120
rect 13378 2086 13394 2120
rect 13520 2086 13536 2120
rect 13636 2086 13652 2120
rect 13778 2086 13794 2120
rect 13894 2086 13910 2120
rect 14036 2086 14052 2120
rect 14152 2086 14168 2120
rect 14294 2086 14310 2120
rect 14410 2086 14426 2120
rect 14552 2086 14568 2120
rect 14668 2086 14684 2120
rect 14810 2086 14826 2120
rect 14926 2086 14942 2120
rect 15068 2086 15084 2120
rect 15184 2086 15200 2120
rect 15326 2086 15342 2120
rect 15442 2086 15458 2120
rect 16300 2086 16316 2120
rect 16416 2086 16432 2120
rect 16558 2086 16574 2120
rect 16674 2086 16690 2120
rect 16816 2086 16832 2120
rect 16932 2086 16948 2120
rect 17074 2086 17090 2120
rect 17190 2086 17206 2120
rect 17332 2086 17348 2120
rect 17448 2086 17464 2120
rect 17590 2086 17606 2120
rect 17706 2086 17722 2120
rect 17848 2086 17864 2120
rect 17964 2086 17980 2120
rect 18106 2086 18122 2120
rect 18222 2086 18238 2120
rect 18364 2086 18380 2120
rect 18480 2086 18496 2120
rect 18622 2086 18638 2120
rect 18738 2086 18754 2120
rect 19596 2086 19612 2120
rect 19712 2086 19728 2120
rect 19854 2086 19870 2120
rect 19970 2086 19986 2120
rect 20112 2086 20128 2120
rect 20228 2086 20244 2120
rect 20370 2086 20386 2120
rect 20486 2086 20502 2120
rect 20628 2086 20644 2120
rect 20744 2086 20760 2120
rect 20886 2086 20902 2120
rect 21002 2086 21018 2120
rect 21144 2086 21160 2120
rect 21260 2086 21276 2120
rect 21402 2086 21418 2120
rect 21518 2086 21534 2120
rect 21660 2086 21676 2120
rect 21776 2086 21792 2120
rect 21918 2086 21934 2120
rect 22034 2086 22050 2120
rect 12576 1488 12592 1522
rect 13052 1488 13068 1522
rect 13434 1488 13450 1522
rect 13910 1488 13926 1522
rect 14292 1488 14308 1522
rect 14768 1488 14784 1522
rect 15150 1488 15166 1522
rect 15626 1488 15642 1522
rect 16008 1488 16024 1522
rect 16484 1488 16500 1522
rect 16866 1488 16882 1522
rect 17342 1488 17358 1522
rect 17724 1488 17740 1522
rect 18200 1488 18216 1522
rect 18582 1488 18598 1522
rect 19058 1488 19074 1522
rect 19440 1488 19456 1522
rect 19916 1488 19932 1522
rect 20298 1488 20314 1522
rect 20774 1488 20790 1522
rect 21156 1488 21172 1522
rect 21632 1488 21648 1522
rect 22014 1488 22030 1522
rect 22490 1488 22506 1522
rect 12376 1438 12410 1454
rect 12376 1246 12410 1262
rect 13234 1438 13268 1454
rect 13234 1246 13268 1262
rect 14092 1438 14126 1454
rect 14092 1246 14126 1262
rect 14950 1438 14984 1454
rect 14950 1246 14984 1262
rect 15808 1438 15842 1454
rect 15808 1246 15842 1262
rect 16666 1438 16700 1454
rect 16666 1246 16700 1262
rect 17524 1438 17558 1454
rect 17524 1246 17558 1262
rect 18382 1438 18416 1454
rect 18382 1246 18416 1262
rect 19240 1438 19274 1454
rect 19240 1246 19274 1262
rect 20098 1438 20132 1454
rect 20098 1246 20132 1262
rect 20956 1438 20990 1454
rect 20956 1246 20990 1262
rect 21814 1438 21848 1454
rect 21814 1246 21848 1262
rect 22672 1438 22706 1454
rect 22672 1246 22706 1262
rect 12576 1178 12592 1212
rect 13052 1178 13068 1212
rect 13434 1178 13450 1212
rect 13910 1178 13926 1212
rect 14292 1178 14308 1212
rect 14768 1178 14784 1212
rect 15150 1178 15166 1212
rect 15626 1178 15642 1212
rect 16008 1178 16024 1212
rect 16484 1178 16500 1212
rect 16866 1178 16882 1212
rect 17342 1178 17358 1212
rect 17724 1178 17740 1212
rect 18200 1178 18216 1212
rect 18582 1178 18598 1212
rect 19058 1178 19074 1212
rect 19440 1178 19456 1212
rect 19916 1178 19932 1212
rect 20298 1178 20314 1212
rect 20774 1178 20790 1212
rect 21156 1178 21172 1212
rect 21632 1178 21648 1212
rect 22014 1178 22030 1212
rect 22490 1178 22506 1212
rect 12576 948 12592 982
rect 13052 948 13068 982
rect 13434 948 13450 982
rect 13910 948 13926 982
rect 14292 948 14308 982
rect 14768 948 14784 982
rect 15150 948 15166 982
rect 15626 948 15642 982
rect 16008 948 16024 982
rect 16484 948 16500 982
rect 16866 948 16882 982
rect 17342 948 17358 982
rect 17724 948 17740 982
rect 18200 948 18216 982
rect 18582 948 18598 982
rect 19058 948 19074 982
rect 19440 948 19456 982
rect 19916 948 19932 982
rect 20298 948 20314 982
rect 20774 948 20790 982
rect 21156 948 21172 982
rect 21632 948 21648 982
rect 22014 948 22030 982
rect 22490 948 22506 982
rect 12376 898 12410 914
rect 12376 706 12410 722
rect 13234 898 13268 914
rect 13234 706 13268 722
rect 14092 898 14126 914
rect 14092 706 14126 722
rect 14950 898 14984 914
rect 14950 706 14984 722
rect 15808 898 15842 914
rect 15808 706 15842 722
rect 16666 898 16700 914
rect 16666 706 16700 722
rect 17524 898 17558 914
rect 17524 706 17558 722
rect 18382 898 18416 914
rect 18382 706 18416 722
rect 19240 898 19274 914
rect 19240 706 19274 722
rect 20098 898 20132 914
rect 20098 706 20132 722
rect 20956 898 20990 914
rect 20956 706 20990 722
rect 21814 898 21848 914
rect 21814 706 21848 722
rect 22672 898 22706 914
rect 22672 706 22706 722
rect 12576 638 12592 672
rect 13052 638 13068 672
rect 13434 638 13450 672
rect 13910 638 13926 672
rect 14292 638 14308 672
rect 14768 638 14784 672
rect 15150 638 15166 672
rect 15626 638 15642 672
rect 16008 638 16024 672
rect 16484 638 16500 672
rect 16866 638 16882 672
rect 17342 638 17358 672
rect 17724 638 17740 672
rect 18200 638 18216 672
rect 18582 638 18598 672
rect 19058 638 19074 672
rect 19440 638 19456 672
rect 19916 638 19932 672
rect 20298 638 20314 672
rect 20774 638 20790 672
rect 21156 638 21172 672
rect 21632 638 21648 672
rect 22014 638 22030 672
rect 22490 638 22506 672
rect 11866 -286 11966 -124
rect 23110 -286 23210 -124
rect 66 -680 166 -518
rect 11310 -680 11410 -518
rect 776 -1476 792 -1442
rect 1252 -1476 1268 -1442
rect 1634 -1476 1650 -1442
rect 2110 -1476 2126 -1442
rect 2492 -1476 2508 -1442
rect 2968 -1476 2984 -1442
rect 3350 -1476 3366 -1442
rect 3826 -1476 3842 -1442
rect 4208 -1476 4224 -1442
rect 4684 -1476 4700 -1442
rect 5066 -1476 5082 -1442
rect 5542 -1476 5558 -1442
rect 5924 -1476 5940 -1442
rect 6400 -1476 6416 -1442
rect 6782 -1476 6798 -1442
rect 7258 -1476 7274 -1442
rect 7640 -1476 7656 -1442
rect 8116 -1476 8132 -1442
rect 8498 -1476 8514 -1442
rect 8974 -1476 8990 -1442
rect 9356 -1476 9372 -1442
rect 9832 -1476 9848 -1442
rect 10214 -1476 10230 -1442
rect 10690 -1476 10706 -1442
rect 576 -1526 610 -1510
rect 576 -1718 610 -1702
rect 1434 -1526 1468 -1510
rect 1434 -1718 1468 -1702
rect 2292 -1526 2326 -1510
rect 2292 -1718 2326 -1702
rect 3150 -1526 3184 -1510
rect 3150 -1718 3184 -1702
rect 4008 -1526 4042 -1510
rect 4008 -1718 4042 -1702
rect 4866 -1526 4900 -1510
rect 4866 -1718 4900 -1702
rect 5724 -1526 5758 -1510
rect 5724 -1718 5758 -1702
rect 6582 -1526 6616 -1510
rect 6582 -1718 6616 -1702
rect 7440 -1526 7474 -1510
rect 7440 -1718 7474 -1702
rect 8298 -1526 8332 -1510
rect 8298 -1718 8332 -1702
rect 9156 -1526 9190 -1510
rect 9156 -1718 9190 -1702
rect 10014 -1526 10048 -1510
rect 10014 -1718 10048 -1702
rect 10872 -1526 10906 -1510
rect 10872 -1718 10906 -1702
rect 776 -1786 792 -1752
rect 1252 -1786 1268 -1752
rect 1634 -1786 1650 -1752
rect 2110 -1786 2126 -1752
rect 2492 -1786 2508 -1752
rect 2968 -1786 2984 -1752
rect 3350 -1786 3366 -1752
rect 3826 -1786 3842 -1752
rect 4208 -1786 4224 -1752
rect 4684 -1786 4700 -1752
rect 5066 -1786 5082 -1752
rect 5542 -1786 5558 -1752
rect 5924 -1786 5940 -1752
rect 6400 -1786 6416 -1752
rect 6782 -1786 6798 -1752
rect 7258 -1786 7274 -1752
rect 7640 -1786 7656 -1752
rect 8116 -1786 8132 -1752
rect 8498 -1786 8514 -1752
rect 8974 -1786 8990 -1752
rect 9356 -1786 9372 -1752
rect 9832 -1786 9848 -1752
rect 10214 -1786 10230 -1752
rect 10690 -1786 10706 -1752
rect 776 -2016 792 -1982
rect 1252 -2016 1268 -1982
rect 1634 -2016 1650 -1982
rect 2110 -2016 2126 -1982
rect 2492 -2016 2508 -1982
rect 2968 -2016 2984 -1982
rect 3350 -2016 3366 -1982
rect 3826 -2016 3842 -1982
rect 4208 -2016 4224 -1982
rect 4684 -2016 4700 -1982
rect 5066 -2016 5082 -1982
rect 5542 -2016 5558 -1982
rect 5924 -2016 5940 -1982
rect 6400 -2016 6416 -1982
rect 6782 -2016 6798 -1982
rect 7258 -2016 7274 -1982
rect 7640 -2016 7656 -1982
rect 8116 -2016 8132 -1982
rect 8498 -2016 8514 -1982
rect 8974 -2016 8990 -1982
rect 9356 -2016 9372 -1982
rect 9832 -2016 9848 -1982
rect 10214 -2016 10230 -1982
rect 10690 -2016 10706 -1982
rect 576 -2066 610 -2050
rect 576 -2258 610 -2242
rect 1434 -2066 1468 -2050
rect 1434 -2258 1468 -2242
rect 2292 -2066 2326 -2050
rect 2292 -2258 2326 -2242
rect 3150 -2066 3184 -2050
rect 3150 -2258 3184 -2242
rect 4008 -2066 4042 -2050
rect 4008 -2258 4042 -2242
rect 4866 -2066 4900 -2050
rect 4866 -2258 4900 -2242
rect 5724 -2066 5758 -2050
rect 5724 -2258 5758 -2242
rect 6582 -2066 6616 -2050
rect 6582 -2258 6616 -2242
rect 7440 -2066 7474 -2050
rect 7440 -2258 7474 -2242
rect 8298 -2066 8332 -2050
rect 8298 -2258 8332 -2242
rect 9156 -2066 9190 -2050
rect 9156 -2258 9190 -2242
rect 10014 -2066 10048 -2050
rect 10014 -2258 10048 -2242
rect 10872 -2066 10906 -2050
rect 10872 -2258 10906 -2242
rect 776 -2326 792 -2292
rect 1252 -2326 1268 -2292
rect 1634 -2326 1650 -2292
rect 2110 -2326 2126 -2292
rect 2492 -2326 2508 -2292
rect 2968 -2326 2984 -2292
rect 3350 -2326 3366 -2292
rect 3826 -2326 3842 -2292
rect 4208 -2326 4224 -2292
rect 4684 -2326 4700 -2292
rect 5066 -2326 5082 -2292
rect 5542 -2326 5558 -2292
rect 5924 -2326 5940 -2292
rect 6400 -2326 6416 -2292
rect 6782 -2326 6798 -2292
rect 7258 -2326 7274 -2292
rect 7640 -2326 7656 -2292
rect 8116 -2326 8132 -2292
rect 8498 -2326 8514 -2292
rect 8974 -2326 8990 -2292
rect 9356 -2326 9372 -2292
rect 9832 -2326 9848 -2292
rect 10214 -2326 10230 -2292
rect 10690 -2326 10706 -2292
rect 1204 -2924 1220 -2890
rect 1320 -2924 1336 -2890
rect 1462 -2924 1478 -2890
rect 1578 -2924 1594 -2890
rect 1720 -2924 1736 -2890
rect 1836 -2924 1852 -2890
rect 1978 -2924 1994 -2890
rect 2094 -2924 2110 -2890
rect 2236 -2924 2252 -2890
rect 2352 -2924 2368 -2890
rect 2494 -2924 2510 -2890
rect 2610 -2924 2626 -2890
rect 2752 -2924 2768 -2890
rect 2868 -2924 2884 -2890
rect 3010 -2924 3026 -2890
rect 3126 -2924 3142 -2890
rect 3268 -2924 3284 -2890
rect 3384 -2924 3400 -2890
rect 3526 -2924 3542 -2890
rect 3642 -2924 3658 -2890
rect 4500 -2924 4516 -2890
rect 4616 -2924 4632 -2890
rect 4758 -2924 4774 -2890
rect 4874 -2924 4890 -2890
rect 5016 -2924 5032 -2890
rect 5132 -2924 5148 -2890
rect 5274 -2924 5290 -2890
rect 5390 -2924 5406 -2890
rect 5532 -2924 5548 -2890
rect 5648 -2924 5664 -2890
rect 5790 -2924 5806 -2890
rect 5906 -2924 5922 -2890
rect 6048 -2924 6064 -2890
rect 6164 -2924 6180 -2890
rect 6306 -2924 6322 -2890
rect 6422 -2924 6438 -2890
rect 6564 -2924 6580 -2890
rect 6680 -2924 6696 -2890
rect 6822 -2924 6838 -2890
rect 6938 -2924 6954 -2890
rect 7796 -2924 7812 -2890
rect 7912 -2924 7928 -2890
rect 8054 -2924 8070 -2890
rect 8170 -2924 8186 -2890
rect 8312 -2924 8328 -2890
rect 8428 -2924 8444 -2890
rect 8570 -2924 8586 -2890
rect 8686 -2924 8702 -2890
rect 8828 -2924 8844 -2890
rect 8944 -2924 8960 -2890
rect 9086 -2924 9102 -2890
rect 9202 -2924 9218 -2890
rect 9344 -2924 9360 -2890
rect 9460 -2924 9476 -2890
rect 9602 -2924 9618 -2890
rect 9718 -2924 9734 -2890
rect 9860 -2924 9876 -2890
rect 9976 -2924 9992 -2890
rect 10118 -2924 10134 -2890
rect 10234 -2924 10250 -2890
rect 1124 -2974 1158 -2958
rect 1124 -3366 1158 -3350
rect 1382 -2974 1416 -2958
rect 1382 -3366 1416 -3350
rect 1640 -2974 1674 -2958
rect 1640 -3366 1674 -3350
rect 1898 -2974 1932 -2958
rect 1898 -3366 1932 -3350
rect 2156 -2974 2190 -2958
rect 2156 -3366 2190 -3350
rect 2414 -2974 2448 -2958
rect 2414 -3366 2448 -3350
rect 2672 -2974 2706 -2958
rect 2672 -3366 2706 -3350
rect 2930 -2974 2964 -2958
rect 2930 -3366 2964 -3350
rect 3188 -2974 3222 -2958
rect 3188 -3366 3222 -3350
rect 3446 -2974 3480 -2958
rect 3446 -3366 3480 -3350
rect 3704 -2974 3738 -2958
rect 3704 -3366 3738 -3350
rect 4420 -2974 4454 -2958
rect 4420 -3366 4454 -3350
rect 4678 -2974 4712 -2958
rect 4678 -3366 4712 -3350
rect 4936 -2974 4970 -2958
rect 4936 -3366 4970 -3350
rect 5194 -2974 5228 -2958
rect 5194 -3366 5228 -3350
rect 5452 -2974 5486 -2958
rect 5452 -3366 5486 -3350
rect 5710 -2974 5744 -2958
rect 5710 -3366 5744 -3350
rect 5968 -2974 6002 -2958
rect 5968 -3366 6002 -3350
rect 6226 -2974 6260 -2958
rect 6226 -3366 6260 -3350
rect 6484 -2974 6518 -2958
rect 6484 -3366 6518 -3350
rect 6742 -2974 6776 -2958
rect 6742 -3366 6776 -3350
rect 7000 -2974 7034 -2958
rect 7000 -3366 7034 -3350
rect 7716 -2974 7750 -2958
rect 7716 -3366 7750 -3350
rect 7974 -2974 8008 -2958
rect 7974 -3366 8008 -3350
rect 8232 -2974 8266 -2958
rect 8232 -3366 8266 -3350
rect 8490 -2974 8524 -2958
rect 8490 -3366 8524 -3350
rect 8748 -2974 8782 -2958
rect 8748 -3366 8782 -3350
rect 9006 -2974 9040 -2958
rect 9006 -3366 9040 -3350
rect 9264 -2974 9298 -2958
rect 9264 -3366 9298 -3350
rect 9522 -2974 9556 -2958
rect 9522 -3366 9556 -3350
rect 9780 -2974 9814 -2958
rect 9780 -3366 9814 -3350
rect 10038 -2974 10072 -2958
rect 10038 -3366 10072 -3350
rect 10296 -2974 10330 -2958
rect 10296 -3366 10330 -3350
rect 1204 -3434 1220 -3400
rect 1320 -3434 1336 -3400
rect 1462 -3434 1478 -3400
rect 1578 -3434 1594 -3400
rect 1720 -3434 1736 -3400
rect 1836 -3434 1852 -3400
rect 1978 -3434 1994 -3400
rect 2094 -3434 2110 -3400
rect 2236 -3434 2252 -3400
rect 2352 -3434 2368 -3400
rect 2494 -3434 2510 -3400
rect 2610 -3434 2626 -3400
rect 2752 -3434 2768 -3400
rect 2868 -3434 2884 -3400
rect 3010 -3434 3026 -3400
rect 3126 -3434 3142 -3400
rect 3268 -3434 3284 -3400
rect 3384 -3434 3400 -3400
rect 3526 -3434 3542 -3400
rect 3642 -3434 3658 -3400
rect 4500 -3434 4516 -3400
rect 4616 -3434 4632 -3400
rect 4758 -3434 4774 -3400
rect 4874 -3434 4890 -3400
rect 5016 -3434 5032 -3400
rect 5132 -3434 5148 -3400
rect 5274 -3434 5290 -3400
rect 5390 -3434 5406 -3400
rect 5532 -3434 5548 -3400
rect 5648 -3434 5664 -3400
rect 5790 -3434 5806 -3400
rect 5906 -3434 5922 -3400
rect 6048 -3434 6064 -3400
rect 6164 -3434 6180 -3400
rect 6306 -3434 6322 -3400
rect 6422 -3434 6438 -3400
rect 6564 -3434 6580 -3400
rect 6680 -3434 6696 -3400
rect 6822 -3434 6838 -3400
rect 6938 -3434 6954 -3400
rect 7796 -3434 7812 -3400
rect 7912 -3434 7928 -3400
rect 8054 -3434 8070 -3400
rect 8170 -3434 8186 -3400
rect 8312 -3434 8328 -3400
rect 8428 -3434 8444 -3400
rect 8570 -3434 8586 -3400
rect 8686 -3434 8702 -3400
rect 8828 -3434 8844 -3400
rect 8944 -3434 8960 -3400
rect 9086 -3434 9102 -3400
rect 9202 -3434 9218 -3400
rect 9344 -3434 9360 -3400
rect 9460 -3434 9476 -3400
rect 9602 -3434 9618 -3400
rect 9718 -3434 9734 -3400
rect 9860 -3434 9876 -3400
rect 9976 -3434 9992 -3400
rect 10118 -3434 10134 -3400
rect 10234 -3434 10250 -3400
rect 66 -3922 166 -3760
rect 11310 -3922 11410 -3760
rect 11866 -680 11966 -518
rect 23110 -680 23210 -518
rect 12576 -1476 12592 -1442
rect 13052 -1476 13068 -1442
rect 13434 -1476 13450 -1442
rect 13910 -1476 13926 -1442
rect 14292 -1476 14308 -1442
rect 14768 -1476 14784 -1442
rect 15150 -1476 15166 -1442
rect 15626 -1476 15642 -1442
rect 16008 -1476 16024 -1442
rect 16484 -1476 16500 -1442
rect 16866 -1476 16882 -1442
rect 17342 -1476 17358 -1442
rect 17724 -1476 17740 -1442
rect 18200 -1476 18216 -1442
rect 18582 -1476 18598 -1442
rect 19058 -1476 19074 -1442
rect 19440 -1476 19456 -1442
rect 19916 -1476 19932 -1442
rect 20298 -1476 20314 -1442
rect 20774 -1476 20790 -1442
rect 21156 -1476 21172 -1442
rect 21632 -1476 21648 -1442
rect 22014 -1476 22030 -1442
rect 22490 -1476 22506 -1442
rect 12376 -1526 12410 -1510
rect 12376 -1718 12410 -1702
rect 13234 -1526 13268 -1510
rect 13234 -1718 13268 -1702
rect 14092 -1526 14126 -1510
rect 14092 -1718 14126 -1702
rect 14950 -1526 14984 -1510
rect 14950 -1718 14984 -1702
rect 15808 -1526 15842 -1510
rect 15808 -1718 15842 -1702
rect 16666 -1526 16700 -1510
rect 16666 -1718 16700 -1702
rect 17524 -1526 17558 -1510
rect 17524 -1718 17558 -1702
rect 18382 -1526 18416 -1510
rect 18382 -1718 18416 -1702
rect 19240 -1526 19274 -1510
rect 19240 -1718 19274 -1702
rect 20098 -1526 20132 -1510
rect 20098 -1718 20132 -1702
rect 20956 -1526 20990 -1510
rect 20956 -1718 20990 -1702
rect 21814 -1526 21848 -1510
rect 21814 -1718 21848 -1702
rect 22672 -1526 22706 -1510
rect 22672 -1718 22706 -1702
rect 12576 -1786 12592 -1752
rect 13052 -1786 13068 -1752
rect 13434 -1786 13450 -1752
rect 13910 -1786 13926 -1752
rect 14292 -1786 14308 -1752
rect 14768 -1786 14784 -1752
rect 15150 -1786 15166 -1752
rect 15626 -1786 15642 -1752
rect 16008 -1786 16024 -1752
rect 16484 -1786 16500 -1752
rect 16866 -1786 16882 -1752
rect 17342 -1786 17358 -1752
rect 17724 -1786 17740 -1752
rect 18200 -1786 18216 -1752
rect 18582 -1786 18598 -1752
rect 19058 -1786 19074 -1752
rect 19440 -1786 19456 -1752
rect 19916 -1786 19932 -1752
rect 20298 -1786 20314 -1752
rect 20774 -1786 20790 -1752
rect 21156 -1786 21172 -1752
rect 21632 -1786 21648 -1752
rect 22014 -1786 22030 -1752
rect 22490 -1786 22506 -1752
rect 12576 -2016 12592 -1982
rect 13052 -2016 13068 -1982
rect 13434 -2016 13450 -1982
rect 13910 -2016 13926 -1982
rect 14292 -2016 14308 -1982
rect 14768 -2016 14784 -1982
rect 15150 -2016 15166 -1982
rect 15626 -2016 15642 -1982
rect 16008 -2016 16024 -1982
rect 16484 -2016 16500 -1982
rect 16866 -2016 16882 -1982
rect 17342 -2016 17358 -1982
rect 17724 -2016 17740 -1982
rect 18200 -2016 18216 -1982
rect 18582 -2016 18598 -1982
rect 19058 -2016 19074 -1982
rect 19440 -2016 19456 -1982
rect 19916 -2016 19932 -1982
rect 20298 -2016 20314 -1982
rect 20774 -2016 20790 -1982
rect 21156 -2016 21172 -1982
rect 21632 -2016 21648 -1982
rect 22014 -2016 22030 -1982
rect 22490 -2016 22506 -1982
rect 12376 -2066 12410 -2050
rect 12376 -2258 12410 -2242
rect 13234 -2066 13268 -2050
rect 13234 -2258 13268 -2242
rect 14092 -2066 14126 -2050
rect 14092 -2258 14126 -2242
rect 14950 -2066 14984 -2050
rect 14950 -2258 14984 -2242
rect 15808 -2066 15842 -2050
rect 15808 -2258 15842 -2242
rect 16666 -2066 16700 -2050
rect 16666 -2258 16700 -2242
rect 17524 -2066 17558 -2050
rect 17524 -2258 17558 -2242
rect 18382 -2066 18416 -2050
rect 18382 -2258 18416 -2242
rect 19240 -2066 19274 -2050
rect 19240 -2258 19274 -2242
rect 20098 -2066 20132 -2050
rect 20098 -2258 20132 -2242
rect 20956 -2066 20990 -2050
rect 20956 -2258 20990 -2242
rect 21814 -2066 21848 -2050
rect 21814 -2258 21848 -2242
rect 22672 -2066 22706 -2050
rect 22672 -2258 22706 -2242
rect 12576 -2326 12592 -2292
rect 13052 -2326 13068 -2292
rect 13434 -2326 13450 -2292
rect 13910 -2326 13926 -2292
rect 14292 -2326 14308 -2292
rect 14768 -2326 14784 -2292
rect 15150 -2326 15166 -2292
rect 15626 -2326 15642 -2292
rect 16008 -2326 16024 -2292
rect 16484 -2326 16500 -2292
rect 16866 -2326 16882 -2292
rect 17342 -2326 17358 -2292
rect 17724 -2326 17740 -2292
rect 18200 -2326 18216 -2292
rect 18582 -2326 18598 -2292
rect 19058 -2326 19074 -2292
rect 19440 -2326 19456 -2292
rect 19916 -2326 19932 -2292
rect 20298 -2326 20314 -2292
rect 20774 -2326 20790 -2292
rect 21156 -2326 21172 -2292
rect 21632 -2326 21648 -2292
rect 22014 -2326 22030 -2292
rect 22490 -2326 22506 -2292
rect 13004 -2924 13020 -2890
rect 13120 -2924 13136 -2890
rect 13262 -2924 13278 -2890
rect 13378 -2924 13394 -2890
rect 13520 -2924 13536 -2890
rect 13636 -2924 13652 -2890
rect 13778 -2924 13794 -2890
rect 13894 -2924 13910 -2890
rect 14036 -2924 14052 -2890
rect 14152 -2924 14168 -2890
rect 14294 -2924 14310 -2890
rect 14410 -2924 14426 -2890
rect 14552 -2924 14568 -2890
rect 14668 -2924 14684 -2890
rect 14810 -2924 14826 -2890
rect 14926 -2924 14942 -2890
rect 15068 -2924 15084 -2890
rect 15184 -2924 15200 -2890
rect 15326 -2924 15342 -2890
rect 15442 -2924 15458 -2890
rect 16300 -2924 16316 -2890
rect 16416 -2924 16432 -2890
rect 16558 -2924 16574 -2890
rect 16674 -2924 16690 -2890
rect 16816 -2924 16832 -2890
rect 16932 -2924 16948 -2890
rect 17074 -2924 17090 -2890
rect 17190 -2924 17206 -2890
rect 17332 -2924 17348 -2890
rect 17448 -2924 17464 -2890
rect 17590 -2924 17606 -2890
rect 17706 -2924 17722 -2890
rect 17848 -2924 17864 -2890
rect 17964 -2924 17980 -2890
rect 18106 -2924 18122 -2890
rect 18222 -2924 18238 -2890
rect 18364 -2924 18380 -2890
rect 18480 -2924 18496 -2890
rect 18622 -2924 18638 -2890
rect 18738 -2924 18754 -2890
rect 19596 -2924 19612 -2890
rect 19712 -2924 19728 -2890
rect 19854 -2924 19870 -2890
rect 19970 -2924 19986 -2890
rect 20112 -2924 20128 -2890
rect 20228 -2924 20244 -2890
rect 20370 -2924 20386 -2890
rect 20486 -2924 20502 -2890
rect 20628 -2924 20644 -2890
rect 20744 -2924 20760 -2890
rect 20886 -2924 20902 -2890
rect 21002 -2924 21018 -2890
rect 21144 -2924 21160 -2890
rect 21260 -2924 21276 -2890
rect 21402 -2924 21418 -2890
rect 21518 -2924 21534 -2890
rect 21660 -2924 21676 -2890
rect 21776 -2924 21792 -2890
rect 21918 -2924 21934 -2890
rect 22034 -2924 22050 -2890
rect 12924 -2974 12958 -2958
rect 12924 -3366 12958 -3350
rect 13182 -2974 13216 -2958
rect 13182 -3366 13216 -3350
rect 13440 -2974 13474 -2958
rect 13440 -3366 13474 -3350
rect 13698 -2974 13732 -2958
rect 13698 -3366 13732 -3350
rect 13956 -2974 13990 -2958
rect 13956 -3366 13990 -3350
rect 14214 -2974 14248 -2958
rect 14214 -3366 14248 -3350
rect 14472 -2974 14506 -2958
rect 14472 -3366 14506 -3350
rect 14730 -2974 14764 -2958
rect 14730 -3366 14764 -3350
rect 14988 -2974 15022 -2958
rect 14988 -3366 15022 -3350
rect 15246 -2974 15280 -2958
rect 15246 -3366 15280 -3350
rect 15504 -2974 15538 -2958
rect 15504 -3366 15538 -3350
rect 16220 -2974 16254 -2958
rect 16220 -3366 16254 -3350
rect 16478 -2974 16512 -2958
rect 16478 -3366 16512 -3350
rect 16736 -2974 16770 -2958
rect 16736 -3366 16770 -3350
rect 16994 -2974 17028 -2958
rect 16994 -3366 17028 -3350
rect 17252 -2974 17286 -2958
rect 17252 -3366 17286 -3350
rect 17510 -2974 17544 -2958
rect 17510 -3366 17544 -3350
rect 17768 -2974 17802 -2958
rect 17768 -3366 17802 -3350
rect 18026 -2974 18060 -2958
rect 18026 -3366 18060 -3350
rect 18284 -2974 18318 -2958
rect 18284 -3366 18318 -3350
rect 18542 -2974 18576 -2958
rect 18542 -3366 18576 -3350
rect 18800 -2974 18834 -2958
rect 18800 -3366 18834 -3350
rect 19516 -2974 19550 -2958
rect 19516 -3366 19550 -3350
rect 19774 -2974 19808 -2958
rect 19774 -3366 19808 -3350
rect 20032 -2974 20066 -2958
rect 20032 -3366 20066 -3350
rect 20290 -2974 20324 -2958
rect 20290 -3366 20324 -3350
rect 20548 -2974 20582 -2958
rect 20548 -3366 20582 -3350
rect 20806 -2974 20840 -2958
rect 20806 -3366 20840 -3350
rect 21064 -2974 21098 -2958
rect 21064 -3366 21098 -3350
rect 21322 -2974 21356 -2958
rect 21322 -3366 21356 -3350
rect 21580 -2974 21614 -2958
rect 21580 -3366 21614 -3350
rect 21838 -2974 21872 -2958
rect 21838 -3366 21872 -3350
rect 22096 -2974 22130 -2958
rect 22096 -3366 22130 -3350
rect 13004 -3434 13020 -3400
rect 13120 -3434 13136 -3400
rect 13262 -3434 13278 -3400
rect 13378 -3434 13394 -3400
rect 13520 -3434 13536 -3400
rect 13636 -3434 13652 -3400
rect 13778 -3434 13794 -3400
rect 13894 -3434 13910 -3400
rect 14036 -3434 14052 -3400
rect 14152 -3434 14168 -3400
rect 14294 -3434 14310 -3400
rect 14410 -3434 14426 -3400
rect 14552 -3434 14568 -3400
rect 14668 -3434 14684 -3400
rect 14810 -3434 14826 -3400
rect 14926 -3434 14942 -3400
rect 15068 -3434 15084 -3400
rect 15184 -3434 15200 -3400
rect 15326 -3434 15342 -3400
rect 15442 -3434 15458 -3400
rect 16300 -3434 16316 -3400
rect 16416 -3434 16432 -3400
rect 16558 -3434 16574 -3400
rect 16674 -3434 16690 -3400
rect 16816 -3434 16832 -3400
rect 16932 -3434 16948 -3400
rect 17074 -3434 17090 -3400
rect 17190 -3434 17206 -3400
rect 17332 -3434 17348 -3400
rect 17448 -3434 17464 -3400
rect 17590 -3434 17606 -3400
rect 17706 -3434 17722 -3400
rect 17848 -3434 17864 -3400
rect 17964 -3434 17980 -3400
rect 18106 -3434 18122 -3400
rect 18222 -3434 18238 -3400
rect 18364 -3434 18380 -3400
rect 18480 -3434 18496 -3400
rect 18622 -3434 18638 -3400
rect 18738 -3434 18754 -3400
rect 19596 -3434 19612 -3400
rect 19712 -3434 19728 -3400
rect 19854 -3434 19870 -3400
rect 19970 -3434 19986 -3400
rect 20112 -3434 20128 -3400
rect 20228 -3434 20244 -3400
rect 20370 -3434 20386 -3400
rect 20486 -3434 20502 -3400
rect 20628 -3434 20644 -3400
rect 20744 -3434 20760 -3400
rect 20886 -3434 20902 -3400
rect 21002 -3434 21018 -3400
rect 21144 -3434 21160 -3400
rect 21260 -3434 21276 -3400
rect 21402 -3434 21418 -3400
rect 21518 -3434 21534 -3400
rect 21660 -3434 21676 -3400
rect 21776 -3434 21792 -3400
rect 21918 -3434 21934 -3400
rect 22034 -3434 22050 -3400
rect 11866 -3922 11966 -3760
rect 23110 -3922 23210 -3760
rect 66 -4318 166 -4158
rect 11310 -4318 11410 -4158
rect 3988 -4583 4004 -4549
rect 4104 -4583 4120 -4549
rect 4246 -4583 4262 -4549
rect 4362 -4583 4378 -4549
rect 4504 -4583 4520 -4549
rect 4620 -4583 4636 -4549
rect 4762 -4583 4778 -4549
rect 4878 -4583 4894 -4549
rect 5020 -4583 5036 -4549
rect 5136 -4583 5152 -4549
rect 5278 -4583 5294 -4549
rect 5394 -4583 5410 -4549
rect 5536 -4583 5552 -4549
rect 5652 -4583 5668 -4549
rect 5794 -4583 5810 -4549
rect 5910 -4583 5926 -4549
rect 6052 -4583 6068 -4549
rect 6168 -4583 6184 -4549
rect 6310 -4583 6326 -4549
rect 6426 -4583 6442 -4549
rect 6568 -4583 6584 -4549
rect 6684 -4583 6700 -4549
rect 6826 -4583 6842 -4549
rect 6942 -4583 6958 -4549
rect 7084 -4583 7100 -4549
rect 7200 -4583 7216 -4549
rect 7342 -4583 7358 -4549
rect 7458 -4583 7474 -4549
rect 3908 -4642 3942 -4626
rect 3908 -4834 3942 -4818
rect 4166 -4642 4200 -4626
rect 4166 -4834 4200 -4818
rect 4424 -4642 4458 -4626
rect 4424 -4834 4458 -4818
rect 4682 -4642 4716 -4626
rect 4682 -4834 4716 -4818
rect 4940 -4642 4974 -4626
rect 4940 -4834 4974 -4818
rect 5198 -4642 5232 -4626
rect 5198 -4834 5232 -4818
rect 5456 -4642 5490 -4626
rect 5456 -4834 5490 -4818
rect 5714 -4642 5748 -4626
rect 5714 -4834 5748 -4818
rect 5972 -4642 6006 -4626
rect 5972 -4834 6006 -4818
rect 6230 -4642 6264 -4626
rect 6230 -4834 6264 -4818
rect 6488 -4642 6522 -4626
rect 6488 -4834 6522 -4818
rect 6746 -4642 6780 -4626
rect 6746 -4834 6780 -4818
rect 7004 -4642 7038 -4626
rect 7004 -4834 7038 -4818
rect 7262 -4642 7296 -4626
rect 7262 -4834 7296 -4818
rect 7520 -4642 7554 -4626
rect 7520 -4834 7554 -4818
rect 3988 -4911 4004 -4877
rect 4104 -4911 4120 -4877
rect 4246 -4911 4262 -4877
rect 4362 -4911 4378 -4877
rect 4504 -4911 4520 -4877
rect 4620 -4911 4636 -4877
rect 4762 -4911 4778 -4877
rect 4878 -4911 4894 -4877
rect 5020 -4911 5036 -4877
rect 5136 -4911 5152 -4877
rect 5278 -4911 5294 -4877
rect 5394 -4911 5410 -4877
rect 5536 -4911 5552 -4877
rect 5652 -4911 5668 -4877
rect 5794 -4911 5810 -4877
rect 5910 -4911 5926 -4877
rect 6052 -4911 6068 -4877
rect 6168 -4911 6184 -4877
rect 6310 -4911 6326 -4877
rect 6426 -4911 6442 -4877
rect 6568 -4911 6584 -4877
rect 6684 -4911 6700 -4877
rect 6826 -4911 6842 -4877
rect 6942 -4911 6958 -4877
rect 7084 -4911 7100 -4877
rect 7200 -4911 7216 -4877
rect 7342 -4911 7358 -4877
rect 7458 -4911 7474 -4877
rect 66 -5942 166 -5782
rect 11310 -5942 11410 -5782
rect 11866 -4318 11966 -4158
rect 23110 -4318 23210 -4158
rect 15788 -4583 15804 -4549
rect 15904 -4583 15920 -4549
rect 16046 -4583 16062 -4549
rect 16162 -4583 16178 -4549
rect 16304 -4583 16320 -4549
rect 16420 -4583 16436 -4549
rect 16562 -4583 16578 -4549
rect 16678 -4583 16694 -4549
rect 16820 -4583 16836 -4549
rect 16936 -4583 16952 -4549
rect 17078 -4583 17094 -4549
rect 17194 -4583 17210 -4549
rect 17336 -4583 17352 -4549
rect 17452 -4583 17468 -4549
rect 17594 -4583 17610 -4549
rect 17710 -4583 17726 -4549
rect 17852 -4583 17868 -4549
rect 17968 -4583 17984 -4549
rect 18110 -4583 18126 -4549
rect 18226 -4583 18242 -4549
rect 18368 -4583 18384 -4549
rect 18484 -4583 18500 -4549
rect 18626 -4583 18642 -4549
rect 18742 -4583 18758 -4549
rect 18884 -4583 18900 -4549
rect 19000 -4583 19016 -4549
rect 19142 -4583 19158 -4549
rect 19258 -4583 19274 -4549
rect 15708 -4642 15742 -4626
rect 15708 -4834 15742 -4818
rect 15966 -4642 16000 -4626
rect 15966 -4834 16000 -4818
rect 16224 -4642 16258 -4626
rect 16224 -4834 16258 -4818
rect 16482 -4642 16516 -4626
rect 16482 -4834 16516 -4818
rect 16740 -4642 16774 -4626
rect 16740 -4834 16774 -4818
rect 16998 -4642 17032 -4626
rect 16998 -4834 17032 -4818
rect 17256 -4642 17290 -4626
rect 17256 -4834 17290 -4818
rect 17514 -4642 17548 -4626
rect 17514 -4834 17548 -4818
rect 17772 -4642 17806 -4626
rect 17772 -4834 17806 -4818
rect 18030 -4642 18064 -4626
rect 18030 -4834 18064 -4818
rect 18288 -4642 18322 -4626
rect 18288 -4834 18322 -4818
rect 18546 -4642 18580 -4626
rect 18546 -4834 18580 -4818
rect 18804 -4642 18838 -4626
rect 18804 -4834 18838 -4818
rect 19062 -4642 19096 -4626
rect 19062 -4834 19096 -4818
rect 19320 -4642 19354 -4626
rect 19320 -4834 19354 -4818
rect 15788 -4911 15804 -4877
rect 15904 -4911 15920 -4877
rect 16046 -4911 16062 -4877
rect 16162 -4911 16178 -4877
rect 16304 -4911 16320 -4877
rect 16420 -4911 16436 -4877
rect 16562 -4911 16578 -4877
rect 16678 -4911 16694 -4877
rect 16820 -4911 16836 -4877
rect 16936 -4911 16952 -4877
rect 17078 -4911 17094 -4877
rect 17194 -4911 17210 -4877
rect 17336 -4911 17352 -4877
rect 17452 -4911 17468 -4877
rect 17594 -4911 17610 -4877
rect 17710 -4911 17726 -4877
rect 17852 -4911 17868 -4877
rect 17968 -4911 17984 -4877
rect 18110 -4911 18126 -4877
rect 18226 -4911 18242 -4877
rect 18368 -4911 18384 -4877
rect 18484 -4911 18500 -4877
rect 18626 -4911 18642 -4877
rect 18742 -4911 18758 -4877
rect 18884 -4911 18900 -4877
rect 19000 -4911 19016 -4877
rect 19142 -4911 19158 -4877
rect 19258 -4911 19274 -4877
rect 11866 -5942 11966 -5782
rect 23110 -5942 23210 -5782
<< viali >>
rect 166 5038 228 5138
rect 228 5038 11248 5138
rect 11248 5038 11310 5138
rect 66 4976 166 4978
rect 66 3516 166 4976
rect 11310 4976 11410 4978
rect 4012 4073 4096 4107
rect 4270 4073 4354 4107
rect 4528 4073 4612 4107
rect 4786 4073 4870 4107
rect 5044 4073 5128 4107
rect 5302 4073 5386 4107
rect 5560 4073 5644 4107
rect 5818 4073 5902 4107
rect 6076 4073 6160 4107
rect 6334 4073 6418 4107
rect 6592 4073 6676 4107
rect 6850 4073 6934 4107
rect 7108 4073 7192 4107
rect 7366 4073 7450 4107
rect 3908 3838 3942 4014
rect 4166 3838 4200 4014
rect 4424 3838 4458 4014
rect 4682 3838 4716 4014
rect 4940 3838 4974 4014
rect 5198 3838 5232 4014
rect 5456 3838 5490 4014
rect 5714 3838 5748 4014
rect 5972 3838 6006 4014
rect 6230 3838 6264 4014
rect 6488 3838 6522 4014
rect 6746 3838 6780 4014
rect 7004 3838 7038 4014
rect 7262 3838 7296 4014
rect 7520 3838 7554 4014
rect 4012 3745 4096 3779
rect 4270 3745 4354 3779
rect 4528 3745 4612 3779
rect 4786 3745 4870 3779
rect 5044 3745 5128 3779
rect 5302 3745 5386 3779
rect 5560 3745 5644 3779
rect 5818 3745 5902 3779
rect 6076 3745 6160 3779
rect 6334 3745 6418 3779
rect 6592 3745 6676 3779
rect 6850 3745 6934 3779
rect 7108 3745 7192 3779
rect 7366 3745 7450 3779
rect 66 3514 166 3516
rect 11310 3516 11410 4976
rect 11310 3514 11410 3516
rect 166 3354 228 3454
rect 228 3354 11248 3454
rect 11248 3354 11310 3454
rect 11966 5038 12028 5138
rect 12028 5038 23048 5138
rect 23048 5038 23110 5138
rect 11866 4976 11966 4978
rect 11866 3516 11966 4976
rect 23110 4976 23210 4978
rect 15812 4073 15896 4107
rect 16070 4073 16154 4107
rect 16328 4073 16412 4107
rect 16586 4073 16670 4107
rect 16844 4073 16928 4107
rect 17102 4073 17186 4107
rect 17360 4073 17444 4107
rect 17618 4073 17702 4107
rect 17876 4073 17960 4107
rect 18134 4073 18218 4107
rect 18392 4073 18476 4107
rect 18650 4073 18734 4107
rect 18908 4073 18992 4107
rect 19166 4073 19250 4107
rect 15708 3838 15742 4014
rect 15966 3838 16000 4014
rect 16224 3838 16258 4014
rect 16482 3838 16516 4014
rect 16740 3838 16774 4014
rect 16998 3838 17032 4014
rect 17256 3838 17290 4014
rect 17514 3838 17548 4014
rect 17772 3838 17806 4014
rect 18030 3838 18064 4014
rect 18288 3838 18322 4014
rect 18546 3838 18580 4014
rect 18804 3838 18838 4014
rect 19062 3838 19096 4014
rect 19320 3838 19354 4014
rect 15812 3745 15896 3779
rect 16070 3745 16154 3779
rect 16328 3745 16412 3779
rect 16586 3745 16670 3779
rect 16844 3745 16928 3779
rect 17102 3745 17186 3779
rect 17360 3745 17444 3779
rect 17618 3745 17702 3779
rect 17876 3745 17960 3779
rect 18134 3745 18218 3779
rect 18392 3745 18476 3779
rect 18650 3745 18734 3779
rect 18908 3745 18992 3779
rect 19166 3745 19250 3779
rect 11866 3514 11966 3516
rect 23110 3516 23210 4976
rect 23110 3514 23210 3516
rect 11966 3354 12028 3454
rect 12028 3354 23048 3454
rect 23048 3354 23110 3454
rect 166 3018 228 3118
rect 228 3018 11248 3118
rect 11248 3018 11310 3118
rect 66 -26 166 2858
rect 1228 2596 1312 2630
rect 1486 2596 1570 2630
rect 1744 2596 1828 2630
rect 2002 2596 2086 2630
rect 2260 2596 2344 2630
rect 2518 2596 2602 2630
rect 2776 2596 2860 2630
rect 3034 2596 3118 2630
rect 3292 2596 3376 2630
rect 3550 2596 3634 2630
rect 4524 2596 4608 2630
rect 4782 2596 4866 2630
rect 5040 2596 5124 2630
rect 5298 2596 5382 2630
rect 5556 2596 5640 2630
rect 5814 2596 5898 2630
rect 6072 2596 6156 2630
rect 6330 2596 6414 2630
rect 6588 2596 6672 2630
rect 6846 2596 6930 2630
rect 7820 2596 7904 2630
rect 8078 2596 8162 2630
rect 8336 2596 8420 2630
rect 8594 2596 8678 2630
rect 8852 2596 8936 2630
rect 9110 2596 9194 2630
rect 9368 2596 9452 2630
rect 9626 2596 9710 2630
rect 9884 2596 9968 2630
rect 10142 2596 10226 2630
rect 1124 2170 1158 2546
rect 1382 2170 1416 2546
rect 1640 2170 1674 2546
rect 1898 2170 1932 2546
rect 2156 2170 2190 2546
rect 2414 2170 2448 2546
rect 2672 2170 2706 2546
rect 2930 2170 2964 2546
rect 3188 2170 3222 2546
rect 3446 2170 3480 2546
rect 3704 2170 3738 2546
rect 4420 2170 4454 2546
rect 4678 2170 4712 2546
rect 4936 2170 4970 2546
rect 5194 2170 5228 2546
rect 5452 2170 5486 2546
rect 5710 2170 5744 2546
rect 5968 2170 6002 2546
rect 6226 2170 6260 2546
rect 6484 2170 6518 2546
rect 6742 2170 6776 2546
rect 7000 2170 7034 2546
rect 7716 2170 7750 2546
rect 7974 2170 8008 2546
rect 8232 2170 8266 2546
rect 8490 2170 8524 2546
rect 8748 2170 8782 2546
rect 9006 2170 9040 2546
rect 9264 2170 9298 2546
rect 9522 2170 9556 2546
rect 9780 2170 9814 2546
rect 10038 2170 10072 2546
rect 10296 2170 10330 2546
rect 1228 2086 1312 2120
rect 1486 2086 1570 2120
rect 1744 2086 1828 2120
rect 2002 2086 2086 2120
rect 2260 2086 2344 2120
rect 2518 2086 2602 2120
rect 2776 2086 2860 2120
rect 3034 2086 3118 2120
rect 3292 2086 3376 2120
rect 3550 2086 3634 2120
rect 4524 2086 4608 2120
rect 4782 2086 4866 2120
rect 5040 2086 5124 2120
rect 5298 2086 5382 2120
rect 5556 2086 5640 2120
rect 5814 2086 5898 2120
rect 6072 2086 6156 2120
rect 6330 2086 6414 2120
rect 6588 2086 6672 2120
rect 6846 2086 6930 2120
rect 7820 2086 7904 2120
rect 8078 2086 8162 2120
rect 8336 2086 8420 2120
rect 8594 2086 8678 2120
rect 8852 2086 8936 2120
rect 9110 2086 9194 2120
rect 9368 2086 9452 2120
rect 9626 2086 9710 2120
rect 9884 2086 9968 2120
rect 10142 2086 10226 2120
rect 830 1488 1214 1522
rect 1688 1488 2072 1522
rect 2546 1488 2930 1522
rect 3404 1488 3788 1522
rect 4262 1488 4646 1522
rect 5120 1488 5504 1522
rect 5978 1488 6362 1522
rect 6836 1488 7220 1522
rect 7694 1488 8078 1522
rect 8552 1488 8936 1522
rect 9410 1488 9794 1522
rect 10268 1488 10652 1522
rect 576 1262 610 1438
rect 1434 1262 1468 1438
rect 2292 1262 2326 1438
rect 3150 1262 3184 1438
rect 4008 1262 4042 1438
rect 4866 1262 4900 1438
rect 5724 1262 5758 1438
rect 6582 1262 6616 1438
rect 7440 1262 7474 1438
rect 8298 1262 8332 1438
rect 9156 1262 9190 1438
rect 10014 1262 10048 1438
rect 10872 1262 10906 1438
rect 830 1178 1214 1212
rect 1688 1178 2072 1212
rect 2546 1178 2930 1212
rect 3404 1178 3788 1212
rect 4262 1178 4646 1212
rect 5120 1178 5504 1212
rect 5978 1178 6362 1212
rect 6836 1178 7220 1212
rect 7694 1178 8078 1212
rect 8552 1178 8936 1212
rect 9410 1178 9794 1212
rect 10268 1178 10652 1212
rect 830 948 1214 982
rect 1688 948 2072 982
rect 2546 948 2930 982
rect 3404 948 3788 982
rect 4262 948 4646 982
rect 5120 948 5504 982
rect 5978 948 6362 982
rect 6836 948 7220 982
rect 7694 948 8078 982
rect 8552 948 8936 982
rect 9410 948 9794 982
rect 10268 948 10652 982
rect 576 722 610 898
rect 1434 722 1468 898
rect 2292 722 2326 898
rect 3150 722 3184 898
rect 4008 722 4042 898
rect 4866 722 4900 898
rect 5724 722 5758 898
rect 6582 722 6616 898
rect 7440 722 7474 898
rect 8298 722 8332 898
rect 9156 722 9190 898
rect 10014 722 10048 898
rect 10872 722 10906 898
rect 830 638 1214 672
rect 1688 638 2072 672
rect 2546 638 2930 672
rect 3404 638 3788 672
rect 4262 638 4646 672
rect 5120 638 5504 672
rect 5978 638 6362 672
rect 6836 638 7220 672
rect 7694 638 8078 672
rect 8552 638 8936 672
rect 9410 638 9794 672
rect 10268 638 10652 672
rect 11310 -26 11410 2858
rect 166 -286 228 -186
rect 228 -286 11248 -186
rect 11248 -286 11310 -186
rect 11966 3018 12028 3118
rect 12028 3018 23048 3118
rect 23048 3018 23110 3118
rect 11866 -26 11966 2858
rect 13028 2596 13112 2630
rect 13286 2596 13370 2630
rect 13544 2596 13628 2630
rect 13802 2596 13886 2630
rect 14060 2596 14144 2630
rect 14318 2596 14402 2630
rect 14576 2596 14660 2630
rect 14834 2596 14918 2630
rect 15092 2596 15176 2630
rect 15350 2596 15434 2630
rect 16324 2596 16408 2630
rect 16582 2596 16666 2630
rect 16840 2596 16924 2630
rect 17098 2596 17182 2630
rect 17356 2596 17440 2630
rect 17614 2596 17698 2630
rect 17872 2596 17956 2630
rect 18130 2596 18214 2630
rect 18388 2596 18472 2630
rect 18646 2596 18730 2630
rect 19620 2596 19704 2630
rect 19878 2596 19962 2630
rect 20136 2596 20220 2630
rect 20394 2596 20478 2630
rect 20652 2596 20736 2630
rect 20910 2596 20994 2630
rect 21168 2596 21252 2630
rect 21426 2596 21510 2630
rect 21684 2596 21768 2630
rect 21942 2596 22026 2630
rect 12924 2170 12958 2546
rect 13182 2170 13216 2546
rect 13440 2170 13474 2546
rect 13698 2170 13732 2546
rect 13956 2170 13990 2546
rect 14214 2170 14248 2546
rect 14472 2170 14506 2546
rect 14730 2170 14764 2546
rect 14988 2170 15022 2546
rect 15246 2170 15280 2546
rect 15504 2170 15538 2546
rect 16220 2170 16254 2546
rect 16478 2170 16512 2546
rect 16736 2170 16770 2546
rect 16994 2170 17028 2546
rect 17252 2170 17286 2546
rect 17510 2170 17544 2546
rect 17768 2170 17802 2546
rect 18026 2170 18060 2546
rect 18284 2170 18318 2546
rect 18542 2170 18576 2546
rect 18800 2170 18834 2546
rect 19516 2170 19550 2546
rect 19774 2170 19808 2546
rect 20032 2170 20066 2546
rect 20290 2170 20324 2546
rect 20548 2170 20582 2546
rect 20806 2170 20840 2546
rect 21064 2170 21098 2546
rect 21322 2170 21356 2546
rect 21580 2170 21614 2546
rect 21838 2170 21872 2546
rect 22096 2170 22130 2546
rect 13028 2086 13112 2120
rect 13286 2086 13370 2120
rect 13544 2086 13628 2120
rect 13802 2086 13886 2120
rect 14060 2086 14144 2120
rect 14318 2086 14402 2120
rect 14576 2086 14660 2120
rect 14834 2086 14918 2120
rect 15092 2086 15176 2120
rect 15350 2086 15434 2120
rect 16324 2086 16408 2120
rect 16582 2086 16666 2120
rect 16840 2086 16924 2120
rect 17098 2086 17182 2120
rect 17356 2086 17440 2120
rect 17614 2086 17698 2120
rect 17872 2086 17956 2120
rect 18130 2086 18214 2120
rect 18388 2086 18472 2120
rect 18646 2086 18730 2120
rect 19620 2086 19704 2120
rect 19878 2086 19962 2120
rect 20136 2086 20220 2120
rect 20394 2086 20478 2120
rect 20652 2086 20736 2120
rect 20910 2086 20994 2120
rect 21168 2086 21252 2120
rect 21426 2086 21510 2120
rect 21684 2086 21768 2120
rect 21942 2086 22026 2120
rect 12630 1488 13014 1522
rect 13488 1488 13872 1522
rect 14346 1488 14730 1522
rect 15204 1488 15588 1522
rect 16062 1488 16446 1522
rect 16920 1488 17304 1522
rect 17778 1488 18162 1522
rect 18636 1488 19020 1522
rect 19494 1488 19878 1522
rect 20352 1488 20736 1522
rect 21210 1488 21594 1522
rect 22068 1488 22452 1522
rect 12376 1262 12410 1438
rect 13234 1262 13268 1438
rect 14092 1262 14126 1438
rect 14950 1262 14984 1438
rect 15808 1262 15842 1438
rect 16666 1262 16700 1438
rect 17524 1262 17558 1438
rect 18382 1262 18416 1438
rect 19240 1262 19274 1438
rect 20098 1262 20132 1438
rect 20956 1262 20990 1438
rect 21814 1262 21848 1438
rect 22672 1262 22706 1438
rect 12630 1178 13014 1212
rect 13488 1178 13872 1212
rect 14346 1178 14730 1212
rect 15204 1178 15588 1212
rect 16062 1178 16446 1212
rect 16920 1178 17304 1212
rect 17778 1178 18162 1212
rect 18636 1178 19020 1212
rect 19494 1178 19878 1212
rect 20352 1178 20736 1212
rect 21210 1178 21594 1212
rect 22068 1178 22452 1212
rect 12630 948 13014 982
rect 13488 948 13872 982
rect 14346 948 14730 982
rect 15204 948 15588 982
rect 16062 948 16446 982
rect 16920 948 17304 982
rect 17778 948 18162 982
rect 18636 948 19020 982
rect 19494 948 19878 982
rect 20352 948 20736 982
rect 21210 948 21594 982
rect 22068 948 22452 982
rect 12376 722 12410 898
rect 13234 722 13268 898
rect 14092 722 14126 898
rect 14950 722 14984 898
rect 15808 722 15842 898
rect 16666 722 16700 898
rect 17524 722 17558 898
rect 18382 722 18416 898
rect 19240 722 19274 898
rect 20098 722 20132 898
rect 20956 722 20990 898
rect 21814 722 21848 898
rect 22672 722 22706 898
rect 12630 638 13014 672
rect 13488 638 13872 672
rect 14346 638 14730 672
rect 15204 638 15588 672
rect 16062 638 16446 672
rect 16920 638 17304 672
rect 17778 638 18162 672
rect 18636 638 19020 672
rect 19494 638 19878 672
rect 20352 638 20736 672
rect 21210 638 21594 672
rect 22068 638 22452 672
rect 23110 -26 23210 2858
rect 11966 -286 12028 -186
rect 12028 -286 23048 -186
rect 23048 -286 23110 -186
rect 166 -618 228 -518
rect 228 -618 11248 -518
rect 11248 -618 11310 -518
rect 66 -3662 166 -778
rect 830 -1476 1214 -1442
rect 1688 -1476 2072 -1442
rect 2546 -1476 2930 -1442
rect 3404 -1476 3788 -1442
rect 4262 -1476 4646 -1442
rect 5120 -1476 5504 -1442
rect 5978 -1476 6362 -1442
rect 6836 -1476 7220 -1442
rect 7694 -1476 8078 -1442
rect 8552 -1476 8936 -1442
rect 9410 -1476 9794 -1442
rect 10268 -1476 10652 -1442
rect 576 -1702 610 -1526
rect 1434 -1702 1468 -1526
rect 2292 -1702 2326 -1526
rect 3150 -1702 3184 -1526
rect 4008 -1702 4042 -1526
rect 4866 -1702 4900 -1526
rect 5724 -1702 5758 -1526
rect 6582 -1702 6616 -1526
rect 7440 -1702 7474 -1526
rect 8298 -1702 8332 -1526
rect 9156 -1702 9190 -1526
rect 10014 -1702 10048 -1526
rect 10872 -1702 10906 -1526
rect 830 -1786 1214 -1752
rect 1688 -1786 2072 -1752
rect 2546 -1786 2930 -1752
rect 3404 -1786 3788 -1752
rect 4262 -1786 4646 -1752
rect 5120 -1786 5504 -1752
rect 5978 -1786 6362 -1752
rect 6836 -1786 7220 -1752
rect 7694 -1786 8078 -1752
rect 8552 -1786 8936 -1752
rect 9410 -1786 9794 -1752
rect 10268 -1786 10652 -1752
rect 830 -2016 1214 -1982
rect 1688 -2016 2072 -1982
rect 2546 -2016 2930 -1982
rect 3404 -2016 3788 -1982
rect 4262 -2016 4646 -1982
rect 5120 -2016 5504 -1982
rect 5978 -2016 6362 -1982
rect 6836 -2016 7220 -1982
rect 7694 -2016 8078 -1982
rect 8552 -2016 8936 -1982
rect 9410 -2016 9794 -1982
rect 10268 -2016 10652 -1982
rect 576 -2242 610 -2066
rect 1434 -2242 1468 -2066
rect 2292 -2242 2326 -2066
rect 3150 -2242 3184 -2066
rect 4008 -2242 4042 -2066
rect 4866 -2242 4900 -2066
rect 5724 -2242 5758 -2066
rect 6582 -2242 6616 -2066
rect 7440 -2242 7474 -2066
rect 8298 -2242 8332 -2066
rect 9156 -2242 9190 -2066
rect 10014 -2242 10048 -2066
rect 10872 -2242 10906 -2066
rect 830 -2326 1214 -2292
rect 1688 -2326 2072 -2292
rect 2546 -2326 2930 -2292
rect 3404 -2326 3788 -2292
rect 4262 -2326 4646 -2292
rect 5120 -2326 5504 -2292
rect 5978 -2326 6362 -2292
rect 6836 -2326 7220 -2292
rect 7694 -2326 8078 -2292
rect 8552 -2326 8936 -2292
rect 9410 -2326 9794 -2292
rect 10268 -2326 10652 -2292
rect 1228 -2924 1312 -2890
rect 1486 -2924 1570 -2890
rect 1744 -2924 1828 -2890
rect 2002 -2924 2086 -2890
rect 2260 -2924 2344 -2890
rect 2518 -2924 2602 -2890
rect 2776 -2924 2860 -2890
rect 3034 -2924 3118 -2890
rect 3292 -2924 3376 -2890
rect 3550 -2924 3634 -2890
rect 4524 -2924 4608 -2890
rect 4782 -2924 4866 -2890
rect 5040 -2924 5124 -2890
rect 5298 -2924 5382 -2890
rect 5556 -2924 5640 -2890
rect 5814 -2924 5898 -2890
rect 6072 -2924 6156 -2890
rect 6330 -2924 6414 -2890
rect 6588 -2924 6672 -2890
rect 6846 -2924 6930 -2890
rect 7820 -2924 7904 -2890
rect 8078 -2924 8162 -2890
rect 8336 -2924 8420 -2890
rect 8594 -2924 8678 -2890
rect 8852 -2924 8936 -2890
rect 9110 -2924 9194 -2890
rect 9368 -2924 9452 -2890
rect 9626 -2924 9710 -2890
rect 9884 -2924 9968 -2890
rect 10142 -2924 10226 -2890
rect 1124 -3350 1158 -2974
rect 1382 -3350 1416 -2974
rect 1640 -3350 1674 -2974
rect 1898 -3350 1932 -2974
rect 2156 -3350 2190 -2974
rect 2414 -3350 2448 -2974
rect 2672 -3350 2706 -2974
rect 2930 -3350 2964 -2974
rect 3188 -3350 3222 -2974
rect 3446 -3350 3480 -2974
rect 3704 -3350 3738 -2974
rect 4420 -3350 4454 -2974
rect 4678 -3350 4712 -2974
rect 4936 -3350 4970 -2974
rect 5194 -3350 5228 -2974
rect 5452 -3350 5486 -2974
rect 5710 -3350 5744 -2974
rect 5968 -3350 6002 -2974
rect 6226 -3350 6260 -2974
rect 6484 -3350 6518 -2974
rect 6742 -3350 6776 -2974
rect 7000 -3350 7034 -2974
rect 7716 -3350 7750 -2974
rect 7974 -3350 8008 -2974
rect 8232 -3350 8266 -2974
rect 8490 -3350 8524 -2974
rect 8748 -3350 8782 -2974
rect 9006 -3350 9040 -2974
rect 9264 -3350 9298 -2974
rect 9522 -3350 9556 -2974
rect 9780 -3350 9814 -2974
rect 10038 -3350 10072 -2974
rect 10296 -3350 10330 -2974
rect 1228 -3434 1312 -3400
rect 1486 -3434 1570 -3400
rect 1744 -3434 1828 -3400
rect 2002 -3434 2086 -3400
rect 2260 -3434 2344 -3400
rect 2518 -3434 2602 -3400
rect 2776 -3434 2860 -3400
rect 3034 -3434 3118 -3400
rect 3292 -3434 3376 -3400
rect 3550 -3434 3634 -3400
rect 4524 -3434 4608 -3400
rect 4782 -3434 4866 -3400
rect 5040 -3434 5124 -3400
rect 5298 -3434 5382 -3400
rect 5556 -3434 5640 -3400
rect 5814 -3434 5898 -3400
rect 6072 -3434 6156 -3400
rect 6330 -3434 6414 -3400
rect 6588 -3434 6672 -3400
rect 6846 -3434 6930 -3400
rect 7820 -3434 7904 -3400
rect 8078 -3434 8162 -3400
rect 8336 -3434 8420 -3400
rect 8594 -3434 8678 -3400
rect 8852 -3434 8936 -3400
rect 9110 -3434 9194 -3400
rect 9368 -3434 9452 -3400
rect 9626 -3434 9710 -3400
rect 9884 -3434 9968 -3400
rect 10142 -3434 10226 -3400
rect 11310 -3662 11410 -778
rect 166 -3922 228 -3822
rect 228 -3922 11248 -3822
rect 11248 -3922 11310 -3822
rect 11966 -618 12028 -518
rect 12028 -618 23048 -518
rect 23048 -618 23110 -518
rect 11866 -3662 11966 -778
rect 12630 -1476 13014 -1442
rect 13488 -1476 13872 -1442
rect 14346 -1476 14730 -1442
rect 15204 -1476 15588 -1442
rect 16062 -1476 16446 -1442
rect 16920 -1476 17304 -1442
rect 17778 -1476 18162 -1442
rect 18636 -1476 19020 -1442
rect 19494 -1476 19878 -1442
rect 20352 -1476 20736 -1442
rect 21210 -1476 21594 -1442
rect 22068 -1476 22452 -1442
rect 12376 -1702 12410 -1526
rect 13234 -1702 13268 -1526
rect 14092 -1702 14126 -1526
rect 14950 -1702 14984 -1526
rect 15808 -1702 15842 -1526
rect 16666 -1702 16700 -1526
rect 17524 -1702 17558 -1526
rect 18382 -1702 18416 -1526
rect 19240 -1702 19274 -1526
rect 20098 -1702 20132 -1526
rect 20956 -1702 20990 -1526
rect 21814 -1702 21848 -1526
rect 22672 -1702 22706 -1526
rect 12630 -1786 13014 -1752
rect 13488 -1786 13872 -1752
rect 14346 -1786 14730 -1752
rect 15204 -1786 15588 -1752
rect 16062 -1786 16446 -1752
rect 16920 -1786 17304 -1752
rect 17778 -1786 18162 -1752
rect 18636 -1786 19020 -1752
rect 19494 -1786 19878 -1752
rect 20352 -1786 20736 -1752
rect 21210 -1786 21594 -1752
rect 22068 -1786 22452 -1752
rect 12630 -2016 13014 -1982
rect 13488 -2016 13872 -1982
rect 14346 -2016 14730 -1982
rect 15204 -2016 15588 -1982
rect 16062 -2016 16446 -1982
rect 16920 -2016 17304 -1982
rect 17778 -2016 18162 -1982
rect 18636 -2016 19020 -1982
rect 19494 -2016 19878 -1982
rect 20352 -2016 20736 -1982
rect 21210 -2016 21594 -1982
rect 22068 -2016 22452 -1982
rect 12376 -2242 12410 -2066
rect 13234 -2242 13268 -2066
rect 14092 -2242 14126 -2066
rect 14950 -2242 14984 -2066
rect 15808 -2242 15842 -2066
rect 16666 -2242 16700 -2066
rect 17524 -2242 17558 -2066
rect 18382 -2242 18416 -2066
rect 19240 -2242 19274 -2066
rect 20098 -2242 20132 -2066
rect 20956 -2242 20990 -2066
rect 21814 -2242 21848 -2066
rect 22672 -2242 22706 -2066
rect 12630 -2326 13014 -2292
rect 13488 -2326 13872 -2292
rect 14346 -2326 14730 -2292
rect 15204 -2326 15588 -2292
rect 16062 -2326 16446 -2292
rect 16920 -2326 17304 -2292
rect 17778 -2326 18162 -2292
rect 18636 -2326 19020 -2292
rect 19494 -2326 19878 -2292
rect 20352 -2326 20736 -2292
rect 21210 -2326 21594 -2292
rect 22068 -2326 22452 -2292
rect 13028 -2924 13112 -2890
rect 13286 -2924 13370 -2890
rect 13544 -2924 13628 -2890
rect 13802 -2924 13886 -2890
rect 14060 -2924 14144 -2890
rect 14318 -2924 14402 -2890
rect 14576 -2924 14660 -2890
rect 14834 -2924 14918 -2890
rect 15092 -2924 15176 -2890
rect 15350 -2924 15434 -2890
rect 16324 -2924 16408 -2890
rect 16582 -2924 16666 -2890
rect 16840 -2924 16924 -2890
rect 17098 -2924 17182 -2890
rect 17356 -2924 17440 -2890
rect 17614 -2924 17698 -2890
rect 17872 -2924 17956 -2890
rect 18130 -2924 18214 -2890
rect 18388 -2924 18472 -2890
rect 18646 -2924 18730 -2890
rect 19620 -2924 19704 -2890
rect 19878 -2924 19962 -2890
rect 20136 -2924 20220 -2890
rect 20394 -2924 20478 -2890
rect 20652 -2924 20736 -2890
rect 20910 -2924 20994 -2890
rect 21168 -2924 21252 -2890
rect 21426 -2924 21510 -2890
rect 21684 -2924 21768 -2890
rect 21942 -2924 22026 -2890
rect 12924 -3350 12958 -2974
rect 13182 -3350 13216 -2974
rect 13440 -3350 13474 -2974
rect 13698 -3350 13732 -2974
rect 13956 -3350 13990 -2974
rect 14214 -3350 14248 -2974
rect 14472 -3350 14506 -2974
rect 14730 -3350 14764 -2974
rect 14988 -3350 15022 -2974
rect 15246 -3350 15280 -2974
rect 15504 -3350 15538 -2974
rect 16220 -3350 16254 -2974
rect 16478 -3350 16512 -2974
rect 16736 -3350 16770 -2974
rect 16994 -3350 17028 -2974
rect 17252 -3350 17286 -2974
rect 17510 -3350 17544 -2974
rect 17768 -3350 17802 -2974
rect 18026 -3350 18060 -2974
rect 18284 -3350 18318 -2974
rect 18542 -3350 18576 -2974
rect 18800 -3350 18834 -2974
rect 19516 -3350 19550 -2974
rect 19774 -3350 19808 -2974
rect 20032 -3350 20066 -2974
rect 20290 -3350 20324 -2974
rect 20548 -3350 20582 -2974
rect 20806 -3350 20840 -2974
rect 21064 -3350 21098 -2974
rect 21322 -3350 21356 -2974
rect 21580 -3350 21614 -2974
rect 21838 -3350 21872 -2974
rect 22096 -3350 22130 -2974
rect 13028 -3434 13112 -3400
rect 13286 -3434 13370 -3400
rect 13544 -3434 13628 -3400
rect 13802 -3434 13886 -3400
rect 14060 -3434 14144 -3400
rect 14318 -3434 14402 -3400
rect 14576 -3434 14660 -3400
rect 14834 -3434 14918 -3400
rect 15092 -3434 15176 -3400
rect 15350 -3434 15434 -3400
rect 16324 -3434 16408 -3400
rect 16582 -3434 16666 -3400
rect 16840 -3434 16924 -3400
rect 17098 -3434 17182 -3400
rect 17356 -3434 17440 -3400
rect 17614 -3434 17698 -3400
rect 17872 -3434 17956 -3400
rect 18130 -3434 18214 -3400
rect 18388 -3434 18472 -3400
rect 18646 -3434 18730 -3400
rect 19620 -3434 19704 -3400
rect 19878 -3434 19962 -3400
rect 20136 -3434 20220 -3400
rect 20394 -3434 20478 -3400
rect 20652 -3434 20736 -3400
rect 20910 -3434 20994 -3400
rect 21168 -3434 21252 -3400
rect 21426 -3434 21510 -3400
rect 21684 -3434 21768 -3400
rect 21942 -3434 22026 -3400
rect 23110 -3662 23210 -778
rect 11966 -3922 12028 -3822
rect 12028 -3922 23048 -3822
rect 23048 -3922 23110 -3822
rect 166 -4258 228 -4158
rect 228 -4258 11248 -4158
rect 11248 -4258 11310 -4158
rect 66 -4320 166 -4318
rect 66 -5780 166 -4320
rect 11310 -4320 11410 -4318
rect 4012 -4583 4096 -4549
rect 4270 -4583 4354 -4549
rect 4528 -4583 4612 -4549
rect 4786 -4583 4870 -4549
rect 5044 -4583 5128 -4549
rect 5302 -4583 5386 -4549
rect 5560 -4583 5644 -4549
rect 5818 -4583 5902 -4549
rect 6076 -4583 6160 -4549
rect 6334 -4583 6418 -4549
rect 6592 -4583 6676 -4549
rect 6850 -4583 6934 -4549
rect 7108 -4583 7192 -4549
rect 7366 -4583 7450 -4549
rect 3908 -4818 3942 -4642
rect 4166 -4818 4200 -4642
rect 4424 -4818 4458 -4642
rect 4682 -4818 4716 -4642
rect 4940 -4818 4974 -4642
rect 5198 -4818 5232 -4642
rect 5456 -4818 5490 -4642
rect 5714 -4818 5748 -4642
rect 5972 -4818 6006 -4642
rect 6230 -4818 6264 -4642
rect 6488 -4818 6522 -4642
rect 6746 -4818 6780 -4642
rect 7004 -4818 7038 -4642
rect 7262 -4818 7296 -4642
rect 7520 -4818 7554 -4642
rect 4012 -4911 4096 -4877
rect 4270 -4911 4354 -4877
rect 4528 -4911 4612 -4877
rect 4786 -4911 4870 -4877
rect 5044 -4911 5128 -4877
rect 5302 -4911 5386 -4877
rect 5560 -4911 5644 -4877
rect 5818 -4911 5902 -4877
rect 6076 -4911 6160 -4877
rect 6334 -4911 6418 -4877
rect 6592 -4911 6676 -4877
rect 6850 -4911 6934 -4877
rect 7108 -4911 7192 -4877
rect 7366 -4911 7450 -4877
rect 66 -5782 166 -5780
rect 11310 -5780 11410 -4320
rect 11310 -5782 11410 -5780
rect 166 -5942 228 -5842
rect 228 -5942 11248 -5842
rect 11248 -5942 11310 -5842
rect 11966 -4258 12028 -4158
rect 12028 -4258 23048 -4158
rect 23048 -4258 23110 -4158
rect 11866 -4320 11966 -4318
rect 11866 -5780 11966 -4320
rect 23110 -4320 23210 -4318
rect 15812 -4583 15896 -4549
rect 16070 -4583 16154 -4549
rect 16328 -4583 16412 -4549
rect 16586 -4583 16670 -4549
rect 16844 -4583 16928 -4549
rect 17102 -4583 17186 -4549
rect 17360 -4583 17444 -4549
rect 17618 -4583 17702 -4549
rect 17876 -4583 17960 -4549
rect 18134 -4583 18218 -4549
rect 18392 -4583 18476 -4549
rect 18650 -4583 18734 -4549
rect 18908 -4583 18992 -4549
rect 19166 -4583 19250 -4549
rect 15708 -4818 15742 -4642
rect 15966 -4818 16000 -4642
rect 16224 -4818 16258 -4642
rect 16482 -4818 16516 -4642
rect 16740 -4818 16774 -4642
rect 16998 -4818 17032 -4642
rect 17256 -4818 17290 -4642
rect 17514 -4818 17548 -4642
rect 17772 -4818 17806 -4642
rect 18030 -4818 18064 -4642
rect 18288 -4818 18322 -4642
rect 18546 -4818 18580 -4642
rect 18804 -4818 18838 -4642
rect 19062 -4818 19096 -4642
rect 19320 -4818 19354 -4642
rect 15812 -4911 15896 -4877
rect 16070 -4911 16154 -4877
rect 16328 -4911 16412 -4877
rect 16586 -4911 16670 -4877
rect 16844 -4911 16928 -4877
rect 17102 -4911 17186 -4877
rect 17360 -4911 17444 -4877
rect 17618 -4911 17702 -4877
rect 17876 -4911 17960 -4877
rect 18134 -4911 18218 -4877
rect 18392 -4911 18476 -4877
rect 18650 -4911 18734 -4877
rect 18908 -4911 18992 -4877
rect 19166 -4911 19250 -4877
rect 11866 -5782 11966 -5780
rect 23110 -5780 23210 -4320
rect 23110 -5782 23210 -5780
rect 11966 -5942 12028 -5842
rect 12028 -5942 23048 -5842
rect 23048 -5942 23110 -5842
<< metal1 >>
rect 60 5138 11416 5144
rect 60 5038 166 5138
rect 11310 5038 11416 5138
rect 60 5032 11416 5038
rect 60 4978 172 5032
rect 60 3514 66 4978
rect 166 3514 172 4978
rect 772 4732 782 5032
rect 10694 4732 10704 5032
rect 11304 4978 11416 5032
rect 3854 4646 7710 4686
rect 3854 4494 3902 4646
rect 7666 4494 7710 4646
rect 3854 4456 7710 4494
rect 60 3460 172 3514
rect 3892 4239 3952 4456
rect 4028 4239 4088 4456
rect 3892 4179 4088 4239
rect 3892 4014 3952 4179
rect 4028 4113 4088 4179
rect 4000 4107 4108 4113
rect 4000 4073 4012 4107
rect 4096 4073 4108 4107
rect 4000 4067 4108 4073
rect 4258 4107 4366 4113
rect 4258 4073 4270 4107
rect 4354 4073 4366 4107
rect 4258 4067 4366 4073
rect 3892 3838 3908 4014
rect 3942 3838 3952 4014
rect 4160 4014 4206 4026
rect 4160 3878 4166 4014
rect 3892 3692 3952 3838
rect 4152 3838 4166 3878
rect 4200 3878 4206 4014
rect 4410 4014 4470 4456
rect 4800 4234 4860 4456
rect 4926 4234 4986 4456
rect 4800 4174 4986 4234
rect 4800 4113 4860 4174
rect 4516 4107 4624 4113
rect 4516 4073 4528 4107
rect 4612 4073 4624 4107
rect 4516 4067 4624 4073
rect 4774 4107 4882 4113
rect 4774 4073 4786 4107
rect 4870 4073 4882 4107
rect 4774 4067 4882 4073
rect 4410 3984 4424 4014
rect 4200 3838 4212 3878
rect 4000 3779 4108 3785
rect 4000 3745 4012 3779
rect 4096 3745 4108 3779
rect 4000 3739 4108 3745
rect 4024 3692 4084 3739
rect 3892 3632 4084 3692
rect 3892 3460 3952 3632
rect 4024 3460 4084 3632
rect 4152 3688 4212 3838
rect 4418 3838 4424 3984
rect 4458 3984 4470 4014
rect 4676 4014 4722 4026
rect 4458 3838 4464 3984
rect 4676 3861 4682 4014
rect 4418 3826 4464 3838
rect 4668 3838 4682 3861
rect 4716 3861 4722 4014
rect 4926 4014 4986 4174
rect 5314 4239 5374 4456
rect 5442 4239 5502 4456
rect 5566 4239 5626 4456
rect 5690 4292 5696 4352
rect 5756 4292 5762 4352
rect 5314 4179 5626 4239
rect 5314 4113 5374 4179
rect 5032 4107 5140 4113
rect 5032 4073 5044 4107
rect 5128 4073 5140 4107
rect 5032 4067 5140 4073
rect 5290 4107 5398 4113
rect 5290 4073 5302 4107
rect 5386 4073 5398 4107
rect 5290 4067 5398 4073
rect 4716 3838 4728 3861
rect 4258 3779 4366 3785
rect 4258 3745 4270 3779
rect 4354 3745 4366 3779
rect 4258 3739 4366 3745
rect 4516 3779 4624 3785
rect 4516 3745 4528 3779
rect 4612 3745 4624 3779
rect 4516 3739 4624 3745
rect 4284 3688 4344 3739
rect 4540 3688 4600 3739
rect 4152 3628 4540 3688
rect 4600 3628 4606 3688
rect 4668 3578 4728 3838
rect 4926 3838 4940 4014
rect 4974 3838 4986 4014
rect 5192 4014 5238 4026
rect 5192 3893 5198 4014
rect 4774 3779 4882 3785
rect 4774 3745 4786 3779
rect 4870 3745 4882 3779
rect 4774 3739 4882 3745
rect 4668 3512 4728 3518
rect 4926 3460 4986 3838
rect 5182 3838 5198 3893
rect 5232 3893 5238 4014
rect 5442 4014 5502 4179
rect 5566 4113 5626 4179
rect 5548 4107 5656 4113
rect 5548 4073 5560 4107
rect 5644 4073 5656 4107
rect 5548 4067 5656 4073
rect 5232 3838 5242 3893
rect 5032 3779 5140 3785
rect 5032 3745 5044 3779
rect 5128 3745 5140 3779
rect 5032 3739 5140 3745
rect 5056 3688 5116 3739
rect 5050 3628 5056 3688
rect 5116 3628 5122 3688
rect 5182 3576 5242 3838
rect 5442 3838 5456 4014
rect 5490 3838 5502 4014
rect 5696 4014 5756 4292
rect 5806 4107 5914 4113
rect 5806 4073 5818 4107
rect 5902 4073 5914 4107
rect 5806 4067 5914 4073
rect 5696 3974 5714 4014
rect 5290 3779 5398 3785
rect 5290 3745 5302 3779
rect 5386 3745 5398 3779
rect 5290 3739 5398 3745
rect 5182 3510 5242 3516
rect 5314 3692 5374 3739
rect 5442 3692 5502 3838
rect 5708 3838 5714 3974
rect 5748 3974 5756 4014
rect 5956 4014 6016 4456
rect 6346 4233 6406 4456
rect 6474 4233 6534 4456
rect 6606 4233 6666 4456
rect 6346 4173 6666 4233
rect 6346 4113 6406 4173
rect 6064 4107 6172 4113
rect 6064 4073 6076 4107
rect 6160 4073 6172 4107
rect 6064 4067 6172 4073
rect 6322 4107 6430 4113
rect 6322 4073 6334 4107
rect 6418 4073 6430 4107
rect 6322 4067 6430 4073
rect 5956 3984 5972 4014
rect 5748 3838 5754 3974
rect 5708 3826 5754 3838
rect 5966 3838 5972 3984
rect 6006 3984 6016 4014
rect 6224 4014 6270 4026
rect 6006 3838 6012 3984
rect 6224 3876 6230 4014
rect 5966 3826 6012 3838
rect 6214 3838 6230 3876
rect 6264 3876 6270 4014
rect 6474 4014 6534 4173
rect 6606 4113 6666 4173
rect 6728 4170 6734 4230
rect 6794 4170 6800 4230
rect 6580 4107 6688 4113
rect 6580 4073 6592 4107
rect 6676 4073 6688 4107
rect 6580 4067 6688 4073
rect 6264 3838 6274 3876
rect 5548 3779 5656 3785
rect 5548 3745 5560 3779
rect 5644 3745 5656 3779
rect 5548 3739 5656 3745
rect 5806 3779 5914 3785
rect 5806 3745 5818 3779
rect 5902 3745 5914 3779
rect 5806 3739 5914 3745
rect 6064 3779 6172 3785
rect 6064 3745 6076 3779
rect 6160 3745 6172 3779
rect 6064 3739 6172 3745
rect 5570 3692 5630 3739
rect 5314 3632 5630 3692
rect 5314 3460 5374 3632
rect 5442 3460 5502 3632
rect 5570 3460 5630 3632
rect 5828 3686 5888 3739
rect 6088 3686 6148 3739
rect 6214 3686 6274 3838
rect 6474 3838 6488 4014
rect 6522 3838 6534 4014
rect 6322 3779 6430 3785
rect 6322 3745 6334 3779
rect 6418 3745 6430 3779
rect 6322 3739 6430 3745
rect 5828 3626 6274 3686
rect 6344 3686 6404 3739
rect 6474 3686 6534 3838
rect 6734 4014 6794 4170
rect 6838 4107 6946 4113
rect 6838 4073 6850 4107
rect 6934 4073 6946 4107
rect 6838 4067 6946 4073
rect 6734 3838 6746 4014
rect 6780 3838 6794 4014
rect 6580 3779 6688 3785
rect 6580 3745 6592 3779
rect 6676 3745 6688 3779
rect 6580 3739 6688 3745
rect 6598 3686 6658 3739
rect 6344 3626 6658 3686
rect 6088 3574 6148 3626
rect 6088 3508 6148 3514
rect 6344 3460 6404 3626
rect 6474 3460 6534 3626
rect 6598 3460 6658 3626
rect 6734 3684 6794 3838
rect 6990 4014 7050 4456
rect 7376 4232 7436 4456
rect 7506 4232 7566 4456
rect 7376 4172 7566 4232
rect 7376 4113 7436 4172
rect 7096 4107 7204 4113
rect 7096 4073 7108 4107
rect 7192 4073 7204 4107
rect 7096 4067 7204 4073
rect 7354 4107 7462 4113
rect 7354 4073 7366 4107
rect 7450 4073 7462 4107
rect 7354 4067 7462 4073
rect 6990 3838 7004 4014
rect 7038 3838 7050 4014
rect 7256 4014 7302 4026
rect 7256 3884 7262 4014
rect 6838 3779 6946 3785
rect 6838 3745 6850 3779
rect 6934 3745 6946 3779
rect 6838 3739 6946 3745
rect 6860 3684 6920 3739
rect 6734 3624 6920 3684
rect 6990 3460 7050 3838
rect 7252 3838 7262 3884
rect 7296 3884 7302 4014
rect 7506 4014 7566 4172
rect 7296 3838 7312 3884
rect 7096 3779 7204 3785
rect 7096 3745 7108 3779
rect 7192 3745 7204 3779
rect 7096 3739 7204 3745
rect 7124 3684 7184 3739
rect 7252 3684 7312 3838
rect 7506 3838 7520 4014
rect 7554 3838 7566 4014
rect 7354 3779 7462 3785
rect 7354 3745 7366 3779
rect 7450 3745 7462 3779
rect 7354 3739 7462 3745
rect 7124 3624 7312 3684
rect 7252 3572 7312 3624
rect 7376 3688 7436 3739
rect 7506 3688 7566 3838
rect 7376 3628 7566 3688
rect 7246 3512 7252 3572
rect 7312 3512 7318 3572
rect 7376 3460 7436 3628
rect 7506 3460 7566 3628
rect 11304 3514 11310 4978
rect 11410 3514 11416 4978
rect 11304 3460 11416 3514
rect 60 3454 11416 3460
rect 60 3354 166 3454
rect 11310 3354 11416 3454
rect 60 3348 11416 3354
rect 11860 5138 23216 5144
rect 11860 5038 11966 5138
rect 23110 5038 23216 5138
rect 11860 5032 23216 5038
rect 11860 4978 11972 5032
rect 11860 3514 11866 4978
rect 11966 3514 11972 4978
rect 12572 4732 12582 5032
rect 22494 4732 22504 5032
rect 23104 4978 23216 5032
rect 15654 4646 19510 4686
rect 15654 4494 15702 4646
rect 19466 4494 19510 4646
rect 15654 4456 19510 4494
rect 11860 3460 11972 3514
rect 15692 4239 15752 4456
rect 15828 4239 15888 4456
rect 15692 4179 15888 4239
rect 15692 4014 15752 4179
rect 15828 4113 15888 4179
rect 15800 4107 15908 4113
rect 15800 4073 15812 4107
rect 15896 4073 15908 4107
rect 15800 4067 15908 4073
rect 16058 4107 16166 4113
rect 16058 4073 16070 4107
rect 16154 4073 16166 4107
rect 16058 4067 16166 4073
rect 15692 3838 15708 4014
rect 15742 3838 15752 4014
rect 15960 4014 16006 4026
rect 15960 3878 15966 4014
rect 15692 3692 15752 3838
rect 15952 3838 15966 3878
rect 16000 3878 16006 4014
rect 16210 4014 16270 4456
rect 16600 4234 16660 4456
rect 16726 4234 16786 4456
rect 16600 4174 16786 4234
rect 16600 4113 16660 4174
rect 16316 4107 16424 4113
rect 16316 4073 16328 4107
rect 16412 4073 16424 4107
rect 16316 4067 16424 4073
rect 16574 4107 16682 4113
rect 16574 4073 16586 4107
rect 16670 4073 16682 4107
rect 16574 4067 16682 4073
rect 16210 3984 16224 4014
rect 16000 3838 16012 3878
rect 15800 3779 15908 3785
rect 15800 3745 15812 3779
rect 15896 3745 15908 3779
rect 15800 3739 15908 3745
rect 15824 3692 15884 3739
rect 15692 3632 15884 3692
rect 15692 3460 15752 3632
rect 15824 3460 15884 3632
rect 15952 3688 16012 3838
rect 16218 3838 16224 3984
rect 16258 3984 16270 4014
rect 16476 4014 16522 4026
rect 16258 3838 16264 3984
rect 16476 3861 16482 4014
rect 16218 3826 16264 3838
rect 16468 3838 16482 3861
rect 16516 3861 16522 4014
rect 16726 4014 16786 4174
rect 17114 4239 17174 4456
rect 17242 4239 17302 4456
rect 17366 4239 17426 4456
rect 17490 4292 17496 4352
rect 17556 4292 17562 4352
rect 17114 4179 17426 4239
rect 17114 4113 17174 4179
rect 16832 4107 16940 4113
rect 16832 4073 16844 4107
rect 16928 4073 16940 4107
rect 16832 4067 16940 4073
rect 17090 4107 17198 4113
rect 17090 4073 17102 4107
rect 17186 4073 17198 4107
rect 17090 4067 17198 4073
rect 16516 3838 16528 3861
rect 16058 3779 16166 3785
rect 16058 3745 16070 3779
rect 16154 3745 16166 3779
rect 16058 3739 16166 3745
rect 16316 3779 16424 3785
rect 16316 3745 16328 3779
rect 16412 3745 16424 3779
rect 16316 3739 16424 3745
rect 16084 3688 16144 3739
rect 16340 3688 16400 3739
rect 15952 3628 16340 3688
rect 16400 3628 16406 3688
rect 16468 3578 16528 3838
rect 16726 3838 16740 4014
rect 16774 3838 16786 4014
rect 16992 4014 17038 4026
rect 16992 3893 16998 4014
rect 16574 3779 16682 3785
rect 16574 3745 16586 3779
rect 16670 3745 16682 3779
rect 16574 3739 16682 3745
rect 16468 3512 16528 3518
rect 16726 3460 16786 3838
rect 16982 3838 16998 3893
rect 17032 3893 17038 4014
rect 17242 4014 17302 4179
rect 17366 4113 17426 4179
rect 17348 4107 17456 4113
rect 17348 4073 17360 4107
rect 17444 4073 17456 4107
rect 17348 4067 17456 4073
rect 17032 3838 17042 3893
rect 16832 3779 16940 3785
rect 16832 3745 16844 3779
rect 16928 3745 16940 3779
rect 16832 3739 16940 3745
rect 16856 3688 16916 3739
rect 16850 3628 16856 3688
rect 16916 3628 16922 3688
rect 16982 3576 17042 3838
rect 17242 3838 17256 4014
rect 17290 3838 17302 4014
rect 17496 4014 17556 4292
rect 17606 4107 17714 4113
rect 17606 4073 17618 4107
rect 17702 4073 17714 4107
rect 17606 4067 17714 4073
rect 17496 3974 17514 4014
rect 17090 3779 17198 3785
rect 17090 3745 17102 3779
rect 17186 3745 17198 3779
rect 17090 3739 17198 3745
rect 16982 3510 17042 3516
rect 17114 3692 17174 3739
rect 17242 3692 17302 3838
rect 17508 3838 17514 3974
rect 17548 3974 17556 4014
rect 17756 4014 17816 4456
rect 18146 4233 18206 4456
rect 18274 4233 18334 4456
rect 18406 4233 18466 4456
rect 18146 4173 18466 4233
rect 18146 4113 18206 4173
rect 17864 4107 17972 4113
rect 17864 4073 17876 4107
rect 17960 4073 17972 4107
rect 17864 4067 17972 4073
rect 18122 4107 18230 4113
rect 18122 4073 18134 4107
rect 18218 4073 18230 4107
rect 18122 4067 18230 4073
rect 17756 3984 17772 4014
rect 17548 3838 17554 3974
rect 17508 3826 17554 3838
rect 17766 3838 17772 3984
rect 17806 3984 17816 4014
rect 18024 4014 18070 4026
rect 17806 3838 17812 3984
rect 18024 3876 18030 4014
rect 17766 3826 17812 3838
rect 18014 3838 18030 3876
rect 18064 3876 18070 4014
rect 18274 4014 18334 4173
rect 18406 4113 18466 4173
rect 18528 4170 18534 4230
rect 18594 4170 18600 4230
rect 18380 4107 18488 4113
rect 18380 4073 18392 4107
rect 18476 4073 18488 4107
rect 18380 4067 18488 4073
rect 18064 3838 18074 3876
rect 17348 3779 17456 3785
rect 17348 3745 17360 3779
rect 17444 3745 17456 3779
rect 17348 3739 17456 3745
rect 17606 3779 17714 3785
rect 17606 3745 17618 3779
rect 17702 3745 17714 3779
rect 17606 3739 17714 3745
rect 17864 3779 17972 3785
rect 17864 3745 17876 3779
rect 17960 3745 17972 3779
rect 17864 3739 17972 3745
rect 17370 3692 17430 3739
rect 17114 3632 17430 3692
rect 17114 3460 17174 3632
rect 17242 3460 17302 3632
rect 17370 3460 17430 3632
rect 17628 3686 17688 3739
rect 17888 3686 17948 3739
rect 18014 3686 18074 3838
rect 18274 3838 18288 4014
rect 18322 3838 18334 4014
rect 18122 3779 18230 3785
rect 18122 3745 18134 3779
rect 18218 3745 18230 3779
rect 18122 3739 18230 3745
rect 17628 3626 18074 3686
rect 18144 3686 18204 3739
rect 18274 3686 18334 3838
rect 18534 4014 18594 4170
rect 18638 4107 18746 4113
rect 18638 4073 18650 4107
rect 18734 4073 18746 4107
rect 18638 4067 18746 4073
rect 18534 3838 18546 4014
rect 18580 3838 18594 4014
rect 18380 3779 18488 3785
rect 18380 3745 18392 3779
rect 18476 3745 18488 3779
rect 18380 3739 18488 3745
rect 18398 3686 18458 3739
rect 18144 3626 18458 3686
rect 17888 3574 17948 3626
rect 17888 3508 17948 3514
rect 18144 3460 18204 3626
rect 18274 3460 18334 3626
rect 18398 3460 18458 3626
rect 18534 3684 18594 3838
rect 18790 4014 18850 4456
rect 19176 4232 19236 4456
rect 19306 4232 19366 4456
rect 19176 4172 19366 4232
rect 19176 4113 19236 4172
rect 18896 4107 19004 4113
rect 18896 4073 18908 4107
rect 18992 4073 19004 4107
rect 18896 4067 19004 4073
rect 19154 4107 19262 4113
rect 19154 4073 19166 4107
rect 19250 4073 19262 4107
rect 19154 4067 19262 4073
rect 18790 3838 18804 4014
rect 18838 3838 18850 4014
rect 19056 4014 19102 4026
rect 19056 3884 19062 4014
rect 18638 3779 18746 3785
rect 18638 3745 18650 3779
rect 18734 3745 18746 3779
rect 18638 3739 18746 3745
rect 18660 3684 18720 3739
rect 18534 3624 18720 3684
rect 18790 3460 18850 3838
rect 19052 3838 19062 3884
rect 19096 3884 19102 4014
rect 19306 4014 19366 4172
rect 19096 3838 19112 3884
rect 18896 3779 19004 3785
rect 18896 3745 18908 3779
rect 18992 3745 19004 3779
rect 18896 3739 19004 3745
rect 18924 3684 18984 3739
rect 19052 3684 19112 3838
rect 19306 3838 19320 4014
rect 19354 3838 19366 4014
rect 19154 3779 19262 3785
rect 19154 3745 19166 3779
rect 19250 3745 19262 3779
rect 19154 3739 19262 3745
rect 18924 3624 19112 3684
rect 19052 3572 19112 3624
rect 19176 3688 19236 3739
rect 19306 3688 19366 3838
rect 19176 3628 19366 3688
rect 19046 3512 19052 3572
rect 19112 3512 19118 3572
rect 19176 3460 19236 3628
rect 19306 3460 19366 3628
rect 23104 3514 23110 4978
rect 23210 3514 23216 4978
rect 23104 3460 23216 3514
rect 11860 3454 23216 3460
rect 11860 3354 11966 3454
rect 23110 3354 23216 3454
rect 11860 3348 23216 3354
rect 3440 3260 3500 3266
rect 6088 3260 6148 3266
rect 8476 3260 8536 3266
rect 3500 3200 6088 3260
rect 6148 3200 8476 3260
rect 3440 3194 3500 3200
rect 6088 3194 6148 3200
rect 8476 3194 8536 3200
rect 15240 3260 15300 3266
rect 17888 3260 17948 3266
rect 20276 3260 20336 3266
rect 15300 3200 17888 3260
rect 17948 3200 20276 3260
rect 15240 3194 15300 3200
rect 17888 3194 17948 3200
rect 20276 3194 20336 3200
rect 60 3118 11416 3124
rect 60 3018 166 3118
rect 11310 3018 11416 3118
rect 60 3012 11416 3018
rect 60 2858 172 3012
rect 60 -26 66 2858
rect 166 2740 172 2858
rect 1114 2740 1174 3012
rect 1240 2740 1300 3012
rect 1876 2906 1882 2966
rect 1942 2906 1948 2966
rect 2912 2906 2918 2966
rect 2978 2906 2984 2966
rect 1362 2790 1368 2850
rect 1428 2790 1434 2850
rect 166 2680 1300 2740
rect 166 2008 172 2680
rect 1114 2546 1174 2680
rect 1240 2636 1300 2680
rect 1216 2630 1324 2636
rect 1216 2596 1228 2630
rect 1312 2596 1324 2630
rect 1216 2590 1324 2596
rect 1114 2170 1124 2546
rect 1158 2170 1174 2546
rect 1368 2546 1428 2790
rect 1752 2680 1758 2740
rect 1818 2680 1824 2740
rect 1758 2636 1818 2680
rect 1474 2630 1582 2636
rect 1474 2596 1486 2630
rect 1570 2596 1582 2630
rect 1474 2590 1582 2596
rect 1732 2630 1840 2636
rect 1732 2596 1744 2630
rect 1828 2596 1840 2630
rect 1732 2590 1840 2596
rect 1368 2496 1382 2546
rect 1114 2008 1174 2170
rect 1376 2170 1382 2496
rect 1416 2496 1428 2546
rect 1634 2546 1680 2558
rect 1416 2170 1422 2496
rect 1634 2190 1640 2546
rect 1376 2158 1422 2170
rect 1628 2170 1640 2190
rect 1674 2190 1680 2546
rect 1882 2546 1942 2906
rect 2394 2790 2400 2850
rect 2460 2790 2466 2850
rect 2006 2680 2012 2740
rect 2072 2680 2078 2740
rect 2012 2636 2072 2680
rect 1990 2630 2098 2636
rect 1990 2596 2002 2630
rect 2086 2596 2098 2630
rect 1990 2590 2098 2596
rect 2248 2630 2356 2636
rect 2248 2596 2260 2630
rect 2344 2596 2356 2630
rect 2248 2590 2356 2596
rect 1882 2500 1898 2546
rect 1674 2170 1688 2190
rect 1216 2120 1324 2126
rect 1216 2086 1228 2120
rect 1312 2086 1324 2120
rect 1216 2080 1324 2086
rect 1474 2120 1582 2126
rect 1474 2086 1486 2120
rect 1570 2086 1582 2120
rect 1474 2080 1582 2086
rect 1240 2008 1300 2080
rect 1498 2010 1558 2080
rect 166 1948 1300 2008
rect 1492 1950 1498 2010
rect 1558 1950 1564 2010
rect 166 -26 172 1948
rect 414 1840 420 1900
rect 480 1840 486 1900
rect 420 566 480 1840
rect 560 1654 620 1948
rect 1628 1900 1688 2170
rect 1892 2170 1898 2500
rect 1932 2500 1942 2546
rect 2150 2546 2196 2558
rect 1932 2170 1938 2500
rect 2150 2190 2156 2546
rect 1892 2158 1938 2170
rect 2140 2170 2156 2190
rect 2190 2190 2196 2546
rect 2400 2546 2460 2790
rect 2778 2680 2784 2740
rect 2844 2680 2850 2740
rect 2784 2636 2844 2680
rect 2506 2630 2614 2636
rect 2506 2596 2518 2630
rect 2602 2596 2614 2630
rect 2506 2590 2614 2596
rect 2764 2630 2872 2636
rect 2764 2596 2776 2630
rect 2860 2596 2872 2630
rect 2764 2590 2872 2596
rect 2784 2586 2844 2590
rect 2400 2486 2414 2546
rect 2190 2170 2200 2190
rect 1732 2120 1840 2126
rect 1732 2086 1744 2120
rect 1828 2086 1840 2120
rect 1732 2080 1840 2086
rect 1990 2120 2098 2126
rect 1990 2086 2002 2120
rect 2086 2086 2098 2120
rect 1990 2080 2098 2086
rect 2140 1900 2200 2170
rect 2408 2170 2414 2486
rect 2448 2486 2460 2546
rect 2666 2546 2712 2558
rect 2448 2170 2454 2486
rect 2666 2194 2672 2546
rect 2408 2158 2454 2170
rect 2660 2170 2672 2194
rect 2706 2194 2712 2546
rect 2918 2546 2978 2906
rect 3430 2790 3436 2850
rect 3496 2790 3502 2850
rect 3040 2680 3046 2740
rect 3106 2680 3112 2740
rect 3046 2636 3106 2680
rect 3022 2630 3130 2636
rect 3022 2596 3034 2630
rect 3118 2596 3130 2630
rect 3022 2590 3130 2596
rect 3280 2630 3388 2636
rect 3280 2596 3292 2630
rect 3376 2596 3388 2630
rect 3280 2590 3388 2596
rect 2918 2496 2930 2546
rect 2706 2170 2720 2194
rect 2248 2120 2356 2126
rect 2248 2086 2260 2120
rect 2344 2086 2356 2120
rect 2248 2080 2356 2086
rect 2506 2120 2614 2126
rect 2506 2086 2518 2120
rect 2602 2086 2614 2120
rect 2506 2080 2614 2086
rect 2274 2010 2334 2080
rect 2528 2010 2588 2080
rect 2268 1950 2274 2010
rect 2334 1950 2340 2010
rect 2522 1950 2528 2010
rect 2588 1950 2594 2010
rect 2660 1900 2720 2170
rect 2924 2170 2930 2496
rect 2964 2496 2978 2546
rect 3182 2546 3228 2558
rect 2964 2170 2970 2496
rect 3182 2194 3188 2546
rect 2924 2158 2970 2170
rect 3176 2170 3188 2194
rect 3222 2194 3228 2546
rect 3436 2546 3496 2790
rect 3560 2740 3620 3012
rect 3694 2740 3754 3012
rect 4410 2740 4470 3012
rect 4534 2740 4594 3012
rect 5172 2912 5178 2972
rect 5238 2912 5244 2972
rect 6208 2912 6214 2972
rect 6274 2912 6280 2972
rect 4658 2796 4664 2856
rect 4724 2796 4730 2856
rect 3560 2680 4594 2740
rect 3560 2636 3620 2680
rect 3538 2630 3646 2636
rect 3538 2596 3550 2630
rect 3634 2596 3646 2630
rect 3538 2590 3646 2596
rect 3436 2490 3446 2546
rect 3222 2170 3236 2194
rect 2764 2120 2872 2126
rect 2764 2086 2776 2120
rect 2860 2086 2872 2120
rect 2764 2080 2872 2086
rect 3022 2120 3130 2126
rect 3022 2086 3034 2120
rect 3118 2086 3130 2120
rect 3022 2080 3130 2086
rect 3176 1900 3236 2170
rect 3440 2170 3446 2490
rect 3480 2490 3496 2546
rect 3694 2546 3754 2680
rect 3480 2170 3486 2490
rect 3440 2158 3486 2170
rect 3694 2170 3704 2546
rect 3738 2170 3754 2546
rect 3280 2120 3388 2126
rect 3280 2086 3292 2120
rect 3376 2086 3388 2120
rect 3280 2080 3388 2086
rect 3538 2120 3646 2126
rect 3538 2086 3550 2120
rect 3634 2086 3646 2120
rect 3538 2080 3646 2086
rect 3306 2010 3366 2080
rect 3300 1950 3306 2010
rect 3366 1950 3372 2010
rect 3560 2008 3620 2080
rect 3694 2008 3754 2170
rect 4410 2546 4470 2680
rect 4534 2636 4594 2680
rect 4512 2630 4620 2636
rect 4512 2596 4524 2630
rect 4608 2596 4620 2630
rect 4512 2590 4620 2596
rect 4410 2170 4420 2546
rect 4454 2170 4470 2546
rect 4664 2546 4724 2796
rect 5048 2686 5054 2746
rect 5114 2686 5120 2746
rect 5054 2636 5114 2686
rect 4770 2630 4878 2636
rect 4770 2596 4782 2630
rect 4866 2596 4878 2630
rect 4770 2590 4878 2596
rect 5028 2630 5136 2636
rect 5028 2596 5040 2630
rect 5124 2596 5136 2630
rect 5028 2590 5136 2596
rect 4664 2502 4678 2546
rect 4410 2008 4470 2170
rect 4672 2170 4678 2502
rect 4712 2502 4724 2546
rect 4930 2546 4976 2558
rect 4712 2170 4718 2502
rect 4930 2196 4936 2546
rect 4672 2158 4718 2170
rect 4924 2170 4936 2196
rect 4970 2196 4976 2546
rect 5178 2546 5238 2912
rect 5690 2796 5696 2856
rect 5756 2796 5762 2856
rect 5302 2686 5308 2746
rect 5368 2686 5374 2746
rect 5308 2636 5368 2686
rect 5286 2630 5394 2636
rect 5286 2596 5298 2630
rect 5382 2596 5394 2630
rect 5286 2590 5394 2596
rect 5544 2630 5652 2636
rect 5544 2596 5556 2630
rect 5640 2596 5652 2630
rect 5544 2590 5652 2596
rect 5178 2506 5194 2546
rect 5188 2258 5194 2506
rect 4970 2170 4984 2196
rect 4512 2120 4620 2126
rect 4512 2086 4524 2120
rect 4608 2086 4620 2120
rect 4512 2080 4620 2086
rect 4770 2120 4878 2126
rect 4770 2086 4782 2120
rect 4866 2086 4878 2120
rect 4770 2080 4878 2086
rect 4536 2008 4596 2080
rect 4794 2016 4854 2080
rect 2134 1840 2140 1900
rect 2200 1840 2206 1900
rect 2654 1840 2660 1900
rect 2720 1840 2726 1900
rect 3170 1840 3176 1900
rect 3236 1840 3242 1900
rect 1628 1834 1688 1840
rect 3306 1778 3366 1950
rect 3560 1948 4596 2008
rect 4788 1956 4794 2016
rect 4854 1956 4860 2016
rect 3300 1718 3306 1778
rect 3366 1718 3372 1778
rect 560 1594 1042 1654
rect 1412 1594 1418 1654
rect 1478 1594 1484 1654
rect 560 1438 620 1594
rect 982 1528 1042 1594
rect 818 1522 1226 1528
rect 818 1488 830 1522
rect 1214 1488 1226 1522
rect 818 1482 1226 1488
rect 560 1262 576 1438
rect 610 1262 620 1438
rect 1418 1438 1478 1594
rect 1676 1522 2084 1528
rect 1676 1488 1688 1522
rect 2072 1488 2084 1522
rect 1676 1482 2084 1488
rect 2534 1522 2942 1528
rect 2534 1488 2546 1522
rect 2930 1488 2942 1522
rect 2534 1482 2942 1488
rect 3392 1522 3800 1528
rect 3392 1488 3404 1522
rect 3788 1488 3800 1522
rect 3392 1482 3800 1488
rect 1418 1400 1434 1438
rect 560 1104 620 1262
rect 1428 1262 1434 1400
rect 1468 1400 1478 1438
rect 2286 1438 2332 1450
rect 1468 1262 1474 1400
rect 2286 1342 2292 1438
rect 1428 1250 1474 1262
rect 2278 1262 2292 1342
rect 2326 1342 2332 1438
rect 3144 1438 3190 1450
rect 2326 1262 2338 1342
rect 3144 1312 3150 1438
rect 818 1212 1226 1218
rect 818 1178 830 1212
rect 1214 1178 1226 1212
rect 818 1172 1226 1178
rect 1676 1212 2084 1218
rect 1676 1178 1688 1212
rect 2072 1178 2084 1212
rect 1676 1172 2084 1178
rect 984 1104 1044 1172
rect 1844 1110 1904 1172
rect 560 1044 1044 1104
rect 1414 1050 1420 1110
rect 1480 1050 1904 1110
rect 560 898 620 1044
rect 984 988 1044 1044
rect 818 982 1226 988
rect 818 948 830 982
rect 1214 948 1226 982
rect 818 942 1226 948
rect 560 722 576 898
rect 610 722 620 898
rect 1420 898 1480 1050
rect 1844 988 1904 1050
rect 1676 982 2084 988
rect 1676 948 1688 982
rect 2072 948 2084 982
rect 1676 942 2084 948
rect 1420 846 1434 898
rect 560 574 620 722
rect 1428 722 1434 846
rect 1468 846 1480 898
rect 2278 898 2338 1262
rect 3136 1262 3150 1312
rect 3184 1312 3190 1438
rect 3994 1438 4054 1948
rect 4924 1906 4984 2170
rect 5186 2170 5194 2258
rect 5228 2506 5238 2546
rect 5446 2546 5492 2558
rect 5228 2258 5234 2506
rect 5228 2170 5246 2258
rect 5446 2196 5452 2546
rect 5028 2120 5136 2126
rect 5028 2086 5040 2120
rect 5124 2086 5136 2120
rect 5028 2080 5136 2086
rect 4924 1654 4984 1846
rect 5186 1778 5246 2170
rect 5436 2170 5452 2196
rect 5486 2196 5492 2546
rect 5696 2546 5756 2796
rect 6074 2686 6080 2746
rect 6140 2686 6146 2746
rect 6080 2636 6140 2686
rect 5802 2630 5910 2636
rect 5802 2596 5814 2630
rect 5898 2596 5910 2630
rect 5802 2590 5910 2596
rect 6060 2630 6168 2636
rect 6060 2596 6072 2630
rect 6156 2596 6168 2630
rect 6060 2590 6168 2596
rect 5696 2492 5710 2546
rect 5486 2170 5496 2196
rect 5286 2120 5394 2126
rect 5286 2086 5298 2120
rect 5382 2086 5394 2120
rect 5286 2080 5394 2086
rect 5436 1906 5496 2170
rect 5704 2170 5710 2492
rect 5744 2492 5756 2546
rect 5962 2546 6008 2558
rect 5744 2170 5750 2492
rect 5962 2200 5968 2546
rect 5704 2158 5750 2170
rect 5956 2170 5968 2200
rect 6002 2200 6008 2546
rect 6214 2546 6274 2912
rect 6726 2796 6732 2856
rect 6792 2796 6798 2856
rect 6336 2686 6342 2746
rect 6402 2686 6408 2746
rect 6342 2636 6402 2686
rect 6318 2630 6426 2636
rect 6318 2596 6330 2630
rect 6414 2596 6426 2630
rect 6318 2590 6426 2596
rect 6576 2630 6684 2636
rect 6576 2596 6588 2630
rect 6672 2596 6684 2630
rect 6576 2590 6684 2596
rect 6214 2502 6226 2546
rect 6002 2170 6016 2200
rect 5544 2120 5652 2126
rect 5544 2086 5556 2120
rect 5640 2086 5652 2120
rect 5544 2080 5652 2086
rect 5802 2120 5910 2126
rect 5802 2086 5814 2120
rect 5898 2086 5910 2120
rect 5802 2080 5910 2086
rect 5570 2016 5630 2080
rect 5824 2016 5884 2080
rect 5564 1956 5570 2016
rect 5630 1956 5636 2016
rect 5818 1956 5824 2016
rect 5884 1956 5890 2016
rect 5956 1906 6016 2170
rect 6220 2170 6226 2502
rect 6260 2502 6274 2546
rect 6478 2546 6524 2558
rect 6260 2170 6266 2502
rect 6478 2200 6484 2546
rect 6220 2158 6266 2170
rect 6472 2170 6484 2200
rect 6518 2200 6524 2546
rect 6732 2546 6792 2796
rect 6858 2746 6918 3012
rect 6990 2746 7050 3012
rect 7706 2746 7766 3012
rect 7830 2746 7890 3012
rect 8468 2906 8474 2966
rect 8534 2906 8540 2966
rect 9504 2906 9510 2966
rect 9570 2906 9576 2966
rect 7954 2790 7960 2850
rect 8020 2790 8026 2850
rect 6858 2686 7890 2746
rect 6858 2636 6918 2686
rect 6834 2630 6942 2636
rect 6834 2596 6846 2630
rect 6930 2596 6942 2630
rect 6834 2590 6942 2596
rect 6732 2496 6742 2546
rect 6518 2170 6532 2200
rect 6060 2120 6168 2126
rect 6060 2086 6072 2120
rect 6156 2086 6168 2120
rect 6060 2080 6168 2086
rect 6318 2120 6426 2126
rect 6318 2086 6330 2120
rect 6414 2086 6426 2120
rect 6318 2080 6426 2086
rect 6472 1906 6532 2170
rect 6736 2170 6742 2496
rect 6776 2496 6792 2546
rect 6990 2546 7050 2686
rect 6776 2170 6782 2496
rect 6736 2158 6782 2170
rect 6990 2170 7000 2546
rect 7034 2170 7050 2546
rect 6576 2120 6684 2126
rect 6576 2086 6588 2120
rect 6672 2086 6684 2120
rect 6576 2080 6684 2086
rect 6834 2120 6942 2126
rect 6834 2086 6846 2120
rect 6930 2086 6942 2120
rect 6834 2080 6942 2086
rect 6602 2016 6662 2080
rect 6596 1956 6602 2016
rect 6662 1956 6668 2016
rect 6856 2014 6916 2080
rect 6990 2014 7050 2170
rect 7706 2546 7766 2686
rect 7830 2636 7890 2686
rect 7808 2630 7916 2636
rect 7808 2596 7820 2630
rect 7904 2596 7916 2630
rect 7808 2590 7916 2596
rect 7706 2170 7716 2546
rect 7750 2170 7766 2546
rect 7960 2546 8020 2790
rect 8344 2680 8350 2740
rect 8410 2680 8416 2740
rect 8350 2636 8410 2680
rect 8066 2630 8174 2636
rect 8066 2596 8078 2630
rect 8162 2596 8174 2630
rect 8066 2590 8174 2596
rect 8324 2630 8432 2636
rect 8324 2596 8336 2630
rect 8420 2596 8432 2630
rect 8324 2590 8432 2596
rect 7960 2496 7974 2546
rect 7706 2014 7766 2170
rect 7968 2170 7974 2496
rect 8008 2496 8020 2546
rect 8226 2546 8272 2558
rect 8008 2170 8014 2496
rect 8226 2190 8232 2546
rect 7968 2158 8014 2170
rect 8220 2170 8232 2190
rect 8266 2190 8272 2546
rect 8474 2546 8534 2906
rect 8986 2790 8992 2850
rect 9052 2790 9058 2850
rect 8598 2680 8604 2740
rect 8664 2680 8670 2740
rect 8604 2636 8664 2680
rect 8582 2630 8690 2636
rect 8582 2596 8594 2630
rect 8678 2596 8690 2630
rect 8582 2590 8690 2596
rect 8840 2630 8948 2636
rect 8840 2596 8852 2630
rect 8936 2596 8948 2630
rect 8840 2590 8948 2596
rect 8474 2500 8490 2546
rect 8266 2170 8280 2190
rect 7808 2120 7916 2126
rect 7808 2086 7820 2120
rect 7904 2086 7916 2120
rect 7808 2080 7916 2086
rect 8066 2120 8174 2126
rect 8066 2086 8078 2120
rect 8162 2086 8174 2120
rect 8066 2080 8174 2086
rect 7832 2014 7892 2080
rect 6856 1954 7892 2014
rect 8090 2010 8150 2080
rect 5430 1846 5436 1906
rect 5496 1846 5502 1906
rect 5950 1846 5956 1906
rect 6016 1846 6022 1906
rect 6466 1846 6472 1906
rect 6532 1846 6538 1906
rect 5180 1718 5186 1778
rect 5246 1718 5252 1778
rect 4846 1594 4852 1654
rect 4912 1594 4984 1654
rect 5282 1596 6206 1656
rect 4250 1522 4658 1528
rect 4250 1488 4262 1522
rect 4646 1488 4658 1522
rect 4250 1482 4658 1488
rect 3184 1262 3196 1312
rect 2534 1212 2942 1218
rect 2534 1178 2546 1212
rect 2930 1178 2942 1212
rect 2534 1172 2942 1178
rect 2702 1110 2762 1172
rect 3136 1110 3196 1262
rect 3994 1262 4008 1438
rect 4042 1262 4054 1438
rect 4852 1438 4912 1594
rect 5282 1528 5342 1596
rect 5108 1522 5516 1528
rect 5108 1488 5120 1522
rect 5504 1488 5516 1522
rect 5108 1482 5516 1488
rect 4852 1396 4866 1438
rect 3392 1212 3800 1218
rect 3392 1178 3404 1212
rect 3788 1178 3800 1212
rect 3392 1172 3800 1178
rect 3566 1110 3626 1172
rect 2696 1054 2702 1110
rect 2762 1054 2768 1110
rect 2696 1050 2768 1054
rect 3130 1050 3136 1110
rect 3196 1050 3202 1110
rect 2702 988 2762 1050
rect 2534 982 2942 988
rect 2534 948 2546 982
rect 2930 948 2942 982
rect 2534 942 2942 948
rect 1468 722 1474 846
rect 1428 710 1474 722
rect 2278 722 2292 898
rect 2326 722 2338 898
rect 3136 898 3196 1050
rect 3566 988 3626 1054
rect 3392 982 3800 988
rect 3392 948 3404 982
rect 3788 948 3800 982
rect 3392 942 3800 948
rect 3136 870 3150 898
rect 818 672 1226 678
rect 818 638 830 672
rect 1214 638 1226 672
rect 818 632 1226 638
rect 1676 672 2084 678
rect 1676 638 1688 672
rect 2072 638 2084 672
rect 1676 632 2084 638
rect 980 574 1040 632
rect 414 506 420 566
rect 480 506 486 566
rect 560 514 1040 574
rect 560 400 620 514
rect 980 400 1040 514
rect 2278 400 2338 722
rect 3144 722 3150 870
rect 3184 870 3196 898
rect 3994 898 4054 1262
rect 4860 1262 4866 1396
rect 4900 1396 4912 1438
rect 5708 1438 5768 1596
rect 6146 1528 6206 1596
rect 5966 1522 6374 1528
rect 5966 1488 5978 1522
rect 6362 1488 6374 1522
rect 5966 1482 6374 1488
rect 6824 1522 7232 1528
rect 6824 1488 6836 1522
rect 7220 1488 7232 1522
rect 6824 1482 7232 1488
rect 4900 1262 4906 1396
rect 4860 1250 4906 1262
rect 5708 1262 5724 1438
rect 5758 1262 5768 1438
rect 6576 1438 6622 1450
rect 6576 1310 6582 1438
rect 4250 1212 4658 1218
rect 4250 1178 4262 1212
rect 4646 1178 4658 1212
rect 4250 1172 4658 1178
rect 5108 1212 5516 1218
rect 5108 1178 5120 1212
rect 5504 1178 5516 1212
rect 5108 1172 5516 1178
rect 4426 1110 4486 1172
rect 5284 1112 5344 1172
rect 5708 1112 5768 1262
rect 6572 1262 6582 1310
rect 6616 1310 6622 1438
rect 7426 1438 7486 1954
rect 8084 1950 8090 2010
rect 8150 1950 8156 2010
rect 8220 1900 8280 2170
rect 8484 2170 8490 2500
rect 8524 2500 8534 2546
rect 8742 2546 8788 2558
rect 8524 2170 8530 2500
rect 8742 2190 8748 2546
rect 8484 2158 8530 2170
rect 8732 2170 8748 2190
rect 8782 2190 8788 2546
rect 8992 2546 9052 2790
rect 9370 2680 9376 2740
rect 9436 2680 9442 2740
rect 9376 2636 9436 2680
rect 9098 2630 9206 2636
rect 9098 2596 9110 2630
rect 9194 2596 9206 2630
rect 9098 2590 9206 2596
rect 9356 2630 9464 2636
rect 9356 2596 9368 2630
rect 9452 2596 9464 2630
rect 9356 2590 9464 2596
rect 9376 2586 9436 2590
rect 8992 2486 9006 2546
rect 8782 2170 8792 2190
rect 8324 2120 8432 2126
rect 8324 2086 8336 2120
rect 8420 2086 8432 2120
rect 8324 2080 8432 2086
rect 8582 2120 8690 2126
rect 8582 2086 8594 2120
rect 8678 2086 8690 2120
rect 8582 2080 8690 2086
rect 8732 1900 8792 2170
rect 9000 2170 9006 2486
rect 9040 2486 9052 2546
rect 9258 2546 9304 2558
rect 9040 2170 9046 2486
rect 9258 2194 9264 2546
rect 9000 2158 9046 2170
rect 9252 2170 9264 2194
rect 9298 2194 9304 2546
rect 9510 2546 9570 2906
rect 10022 2790 10028 2850
rect 10088 2790 10094 2850
rect 9632 2680 9638 2740
rect 9698 2680 9704 2740
rect 9638 2636 9698 2680
rect 9614 2630 9722 2636
rect 9614 2596 9626 2630
rect 9710 2596 9722 2630
rect 9614 2590 9722 2596
rect 9872 2630 9980 2636
rect 9872 2596 9884 2630
rect 9968 2596 9980 2630
rect 9872 2590 9980 2596
rect 9510 2496 9522 2546
rect 9298 2170 9312 2194
rect 8840 2120 8948 2126
rect 8840 2086 8852 2120
rect 8936 2086 8948 2120
rect 8840 2080 8948 2086
rect 9098 2120 9206 2126
rect 9098 2086 9110 2120
rect 9194 2086 9206 2120
rect 9098 2080 9206 2086
rect 8866 2010 8926 2080
rect 9120 2010 9180 2080
rect 8860 1950 8866 2010
rect 8926 1950 8932 2010
rect 9114 1950 9120 2010
rect 9180 1950 9186 2010
rect 9252 1900 9312 2170
rect 9516 2170 9522 2496
rect 9556 2496 9570 2546
rect 9774 2546 9820 2558
rect 9556 2170 9562 2496
rect 9774 2194 9780 2546
rect 9516 2158 9562 2170
rect 9768 2170 9780 2194
rect 9814 2194 9820 2546
rect 10028 2546 10088 2790
rect 10154 2738 10214 3012
rect 10286 2738 10346 3012
rect 11304 2858 11416 3012
rect 11304 2738 11310 2858
rect 10154 2678 11310 2738
rect 10154 2636 10214 2678
rect 10130 2630 10238 2636
rect 10130 2596 10142 2630
rect 10226 2596 10238 2630
rect 10130 2590 10238 2596
rect 10028 2490 10038 2546
rect 9814 2170 9828 2194
rect 9356 2120 9464 2126
rect 9356 2086 9368 2120
rect 9452 2086 9464 2120
rect 9356 2080 9464 2086
rect 9614 2120 9722 2126
rect 9614 2086 9626 2120
rect 9710 2086 9722 2120
rect 9614 2080 9722 2086
rect 9768 1900 9828 2170
rect 10032 2170 10038 2490
rect 10072 2490 10088 2546
rect 10286 2546 10346 2678
rect 10072 2170 10078 2490
rect 10032 2158 10078 2170
rect 10286 2170 10296 2546
rect 10330 2170 10346 2546
rect 9872 2120 9980 2126
rect 9872 2086 9884 2120
rect 9968 2086 9980 2120
rect 9872 2080 9980 2086
rect 10130 2120 10238 2126
rect 10130 2086 10142 2120
rect 10226 2086 10238 2120
rect 10130 2080 10238 2086
rect 9898 2010 9958 2080
rect 9892 1950 9898 2010
rect 9958 1950 9964 2010
rect 10152 2008 10212 2080
rect 10286 2008 10346 2170
rect 11304 2008 11310 2678
rect 10152 1948 11310 2008
rect 8214 1840 8220 1900
rect 8280 1840 8286 1900
rect 8726 1840 8732 1900
rect 8792 1840 8798 1900
rect 9246 1840 9252 1900
rect 9312 1840 9318 1900
rect 9762 1840 9768 1900
rect 9828 1840 9834 1900
rect 9996 1710 10002 1770
rect 10062 1710 10068 1770
rect 7682 1522 8090 1528
rect 7682 1488 7694 1522
rect 8078 1488 8090 1522
rect 7682 1482 8090 1488
rect 8540 1522 8948 1528
rect 8540 1488 8552 1522
rect 8936 1488 8948 1522
rect 8540 1482 8948 1488
rect 9398 1522 9806 1528
rect 9398 1488 9410 1522
rect 9794 1488 9806 1522
rect 9398 1482 9806 1488
rect 6616 1262 6632 1310
rect 5966 1212 6374 1218
rect 5966 1178 5978 1212
rect 6362 1178 6374 1212
rect 5966 1172 6374 1178
rect 6144 1112 6204 1172
rect 4426 988 4486 1054
rect 4850 1050 4856 1110
rect 4916 1050 4922 1110
rect 5284 1052 6204 1112
rect 6572 1110 6632 1262
rect 7426 1262 7440 1438
rect 7474 1262 7486 1438
rect 8292 1438 8338 1450
rect 8292 1326 8298 1438
rect 6824 1212 7232 1218
rect 6824 1178 6836 1212
rect 7220 1178 7232 1212
rect 6824 1172 7232 1178
rect 6998 1110 7058 1172
rect 4250 982 4658 988
rect 4250 948 4262 982
rect 4646 948 4658 982
rect 4250 942 4658 948
rect 3184 722 3190 870
rect 3144 710 3190 722
rect 3994 722 4008 898
rect 4042 722 4054 898
rect 4856 898 4916 1050
rect 5284 988 5344 1052
rect 5108 982 5516 988
rect 5108 948 5120 982
rect 5504 948 5516 982
rect 5108 942 5516 948
rect 4856 846 4866 898
rect 2534 672 2942 678
rect 2534 638 2546 672
rect 2930 638 2942 672
rect 2534 632 2942 638
rect 3392 672 3800 678
rect 3392 638 3404 672
rect 3788 638 3800 672
rect 3392 632 3800 638
rect 3994 400 4054 722
rect 4860 722 4866 846
rect 4900 846 4916 898
rect 5708 898 5768 1052
rect 6144 988 6204 1052
rect 6566 1050 6572 1110
rect 6632 1050 6638 1110
rect 6992 1054 6998 1110
rect 7058 1054 7064 1110
rect 6992 1050 7064 1054
rect 6998 988 7058 1050
rect 5966 982 6374 988
rect 5966 948 5978 982
rect 6362 948 6374 982
rect 5966 942 6374 948
rect 6824 982 7232 988
rect 6824 948 6836 982
rect 7220 948 7232 982
rect 6824 942 7232 948
rect 4900 722 4906 846
rect 4860 710 4906 722
rect 5708 722 5724 898
rect 5758 722 5768 898
rect 6576 898 6622 910
rect 6576 752 6582 898
rect 4250 672 4658 678
rect 4250 638 4262 672
rect 4646 638 4658 672
rect 4250 632 4658 638
rect 5108 672 5516 678
rect 5108 638 5120 672
rect 5504 638 5516 672
rect 5108 632 5516 638
rect 5282 568 5342 632
rect 5708 568 5768 722
rect 6568 722 6582 752
rect 6616 752 6622 898
rect 7426 898 7486 1262
rect 8284 1262 8298 1326
rect 8332 1326 8338 1438
rect 9150 1438 9196 1450
rect 8332 1262 8344 1326
rect 9150 1318 9156 1438
rect 7682 1212 8090 1218
rect 7682 1178 7694 1212
rect 8078 1178 8090 1212
rect 7682 1172 8090 1178
rect 7856 1110 7916 1172
rect 8284 1110 8344 1262
rect 9144 1262 9156 1318
rect 9190 1318 9196 1438
rect 10002 1438 10062 1710
rect 10432 1640 10492 1948
rect 10856 1640 10916 1948
rect 10982 1840 10988 1900
rect 11048 1840 11054 1900
rect 10432 1580 10916 1640
rect 10432 1528 10492 1580
rect 10256 1522 10664 1528
rect 10256 1488 10268 1522
rect 10652 1488 10664 1522
rect 10256 1482 10664 1488
rect 10002 1404 10014 1438
rect 9190 1262 9204 1318
rect 8540 1212 8948 1218
rect 8540 1178 8552 1212
rect 8936 1178 8948 1212
rect 8540 1172 8948 1178
rect 8710 1110 8770 1172
rect 7856 988 7916 1054
rect 8278 1050 8284 1110
rect 8344 1050 8350 1110
rect 7682 982 8090 988
rect 7682 948 7694 982
rect 8078 948 8090 982
rect 7682 942 8090 948
rect 6616 722 6628 752
rect 5966 672 6374 678
rect 5966 638 5978 672
rect 6362 638 6374 672
rect 5966 632 6374 638
rect 6144 568 6204 632
rect 5282 508 6204 568
rect 6568 566 6628 722
rect 7426 722 7440 898
rect 7474 722 7486 898
rect 8284 898 8344 1050
rect 8710 988 8770 1054
rect 8540 982 8948 988
rect 8540 948 8552 982
rect 8936 948 8948 982
rect 8540 942 8948 948
rect 8284 856 8298 898
rect 6824 672 7232 678
rect 6824 638 6836 672
rect 7220 638 7232 672
rect 6824 632 7232 638
rect 5282 400 5342 508
rect 5708 400 5768 508
rect 6144 400 6204 508
rect 6562 506 6568 566
rect 6628 506 6634 566
rect 7426 400 7486 722
rect 8292 722 8298 856
rect 8332 856 8344 898
rect 9144 898 9204 1262
rect 10008 1262 10014 1404
rect 10048 1404 10062 1438
rect 10856 1438 10916 1580
rect 10048 1262 10054 1404
rect 10008 1250 10054 1262
rect 10856 1262 10872 1438
rect 10906 1262 10916 1438
rect 9398 1212 9806 1218
rect 9398 1178 9410 1212
rect 9794 1178 9806 1212
rect 9398 1172 9806 1178
rect 10256 1212 10664 1218
rect 10256 1178 10268 1212
rect 10652 1178 10664 1212
rect 10256 1172 10664 1178
rect 9574 1116 9634 1172
rect 9574 1110 9636 1116
rect 9574 1050 9576 1110
rect 9574 1044 9636 1050
rect 10430 1106 10490 1172
rect 10856 1106 10916 1262
rect 10430 1046 10916 1106
rect 9574 988 9634 1044
rect 10430 988 10490 1046
rect 9398 982 9806 988
rect 9398 948 9410 982
rect 9794 948 9806 982
rect 9398 942 9806 948
rect 10256 982 10664 988
rect 10256 948 10268 982
rect 10652 948 10664 982
rect 10256 942 10664 948
rect 8332 722 8338 856
rect 8292 710 8338 722
rect 9144 722 9156 898
rect 9190 722 9204 898
rect 10008 898 10054 910
rect 10008 754 10014 898
rect 7682 672 8090 678
rect 7682 638 7694 672
rect 8078 638 8090 672
rect 7682 632 8090 638
rect 8540 672 8948 678
rect 8540 638 8552 672
rect 8936 638 8948 672
rect 8540 632 8948 638
rect 9144 400 9204 722
rect 10000 722 10014 754
rect 10048 754 10054 898
rect 10856 898 10916 1046
rect 10048 722 10060 754
rect 9398 672 9806 678
rect 9398 638 9410 672
rect 9794 638 9806 672
rect 9398 632 9806 638
rect 10000 572 10060 722
rect 10856 722 10872 898
rect 10906 722 10916 898
rect 10256 672 10664 678
rect 10256 638 10268 672
rect 10652 638 10664 672
rect 10256 632 10664 638
rect 10432 572 10492 632
rect 10856 572 10916 722
rect 10988 572 11048 1840
rect 9994 512 10000 572
rect 10060 512 10066 572
rect 10432 512 10916 572
rect 10982 512 10988 572
rect 11048 512 11054 572
rect 10432 400 10492 512
rect 10856 400 10916 512
rect 322 352 11096 400
rect 322 242 384 352
rect 11040 242 11096 352
rect 322 186 11096 242
rect 60 -180 172 -26
rect 772 -180 782 120
rect 10694 -180 10704 120
rect 11304 -26 11310 1948
rect 11410 -26 11416 2858
rect 11304 -180 11416 -26
rect 60 -186 11416 -180
rect 60 -286 166 -186
rect 11310 -286 11416 -186
rect 60 -292 11416 -286
rect 11860 3118 23216 3124
rect 11860 3018 11966 3118
rect 23110 3018 23216 3118
rect 11860 3012 23216 3018
rect 11860 2858 11972 3012
rect 11860 -26 11866 2858
rect 11966 2740 11972 2858
rect 12914 2740 12974 3012
rect 13040 2740 13100 3012
rect 13676 2906 13682 2966
rect 13742 2906 13748 2966
rect 14712 2906 14718 2966
rect 14778 2906 14784 2966
rect 13162 2790 13168 2850
rect 13228 2790 13234 2850
rect 11966 2680 13100 2740
rect 11966 2008 11972 2680
rect 12914 2546 12974 2680
rect 13040 2636 13100 2680
rect 13016 2630 13124 2636
rect 13016 2596 13028 2630
rect 13112 2596 13124 2630
rect 13016 2590 13124 2596
rect 12914 2170 12924 2546
rect 12958 2170 12974 2546
rect 13168 2546 13228 2790
rect 13552 2680 13558 2740
rect 13618 2680 13624 2740
rect 13558 2636 13618 2680
rect 13274 2630 13382 2636
rect 13274 2596 13286 2630
rect 13370 2596 13382 2630
rect 13274 2590 13382 2596
rect 13532 2630 13640 2636
rect 13532 2596 13544 2630
rect 13628 2596 13640 2630
rect 13532 2590 13640 2596
rect 13168 2496 13182 2546
rect 12914 2008 12974 2170
rect 13176 2170 13182 2496
rect 13216 2496 13228 2546
rect 13434 2546 13480 2558
rect 13216 2170 13222 2496
rect 13434 2190 13440 2546
rect 13176 2158 13222 2170
rect 13428 2170 13440 2190
rect 13474 2190 13480 2546
rect 13682 2546 13742 2906
rect 14194 2790 14200 2850
rect 14260 2790 14266 2850
rect 13806 2680 13812 2740
rect 13872 2680 13878 2740
rect 13812 2636 13872 2680
rect 13790 2630 13898 2636
rect 13790 2596 13802 2630
rect 13886 2596 13898 2630
rect 13790 2590 13898 2596
rect 14048 2630 14156 2636
rect 14048 2596 14060 2630
rect 14144 2596 14156 2630
rect 14048 2590 14156 2596
rect 13682 2500 13698 2546
rect 13474 2170 13488 2190
rect 13016 2120 13124 2126
rect 13016 2086 13028 2120
rect 13112 2086 13124 2120
rect 13016 2080 13124 2086
rect 13274 2120 13382 2126
rect 13274 2086 13286 2120
rect 13370 2086 13382 2120
rect 13274 2080 13382 2086
rect 13040 2008 13100 2080
rect 13298 2010 13358 2080
rect 11966 1948 13100 2008
rect 13292 1950 13298 2010
rect 13358 1950 13364 2010
rect 11966 -26 11972 1948
rect 12214 1840 12220 1900
rect 12280 1840 12286 1900
rect 12220 566 12280 1840
rect 12360 1654 12420 1948
rect 13428 1900 13488 2170
rect 13692 2170 13698 2500
rect 13732 2500 13742 2546
rect 13950 2546 13996 2558
rect 13732 2170 13738 2500
rect 13950 2190 13956 2546
rect 13692 2158 13738 2170
rect 13940 2170 13956 2190
rect 13990 2190 13996 2546
rect 14200 2546 14260 2790
rect 14578 2680 14584 2740
rect 14644 2680 14650 2740
rect 14584 2636 14644 2680
rect 14306 2630 14414 2636
rect 14306 2596 14318 2630
rect 14402 2596 14414 2630
rect 14306 2590 14414 2596
rect 14564 2630 14672 2636
rect 14564 2596 14576 2630
rect 14660 2596 14672 2630
rect 14564 2590 14672 2596
rect 14584 2586 14644 2590
rect 14200 2486 14214 2546
rect 13990 2170 14000 2190
rect 13532 2120 13640 2126
rect 13532 2086 13544 2120
rect 13628 2086 13640 2120
rect 13532 2080 13640 2086
rect 13790 2120 13898 2126
rect 13790 2086 13802 2120
rect 13886 2086 13898 2120
rect 13790 2080 13898 2086
rect 13940 1900 14000 2170
rect 14208 2170 14214 2486
rect 14248 2486 14260 2546
rect 14466 2546 14512 2558
rect 14248 2170 14254 2486
rect 14466 2194 14472 2546
rect 14208 2158 14254 2170
rect 14460 2170 14472 2194
rect 14506 2194 14512 2546
rect 14718 2546 14778 2906
rect 15230 2790 15236 2850
rect 15296 2790 15302 2850
rect 14840 2680 14846 2740
rect 14906 2680 14912 2740
rect 14846 2636 14906 2680
rect 14822 2630 14930 2636
rect 14822 2596 14834 2630
rect 14918 2596 14930 2630
rect 14822 2590 14930 2596
rect 15080 2630 15188 2636
rect 15080 2596 15092 2630
rect 15176 2596 15188 2630
rect 15080 2590 15188 2596
rect 14718 2496 14730 2546
rect 14506 2170 14520 2194
rect 14048 2120 14156 2126
rect 14048 2086 14060 2120
rect 14144 2086 14156 2120
rect 14048 2080 14156 2086
rect 14306 2120 14414 2126
rect 14306 2086 14318 2120
rect 14402 2086 14414 2120
rect 14306 2080 14414 2086
rect 14074 2010 14134 2080
rect 14328 2010 14388 2080
rect 14068 1950 14074 2010
rect 14134 1950 14140 2010
rect 14322 1950 14328 2010
rect 14388 1950 14394 2010
rect 14460 1900 14520 2170
rect 14724 2170 14730 2496
rect 14764 2496 14778 2546
rect 14982 2546 15028 2558
rect 14764 2170 14770 2496
rect 14982 2194 14988 2546
rect 14724 2158 14770 2170
rect 14976 2170 14988 2194
rect 15022 2194 15028 2546
rect 15236 2546 15296 2790
rect 15360 2740 15420 3012
rect 15494 2740 15554 3012
rect 16210 2740 16270 3012
rect 16334 2740 16394 3012
rect 16972 2912 16978 2972
rect 17038 2912 17044 2972
rect 18008 2912 18014 2972
rect 18074 2912 18080 2972
rect 16458 2796 16464 2856
rect 16524 2796 16530 2856
rect 15360 2680 16394 2740
rect 15360 2636 15420 2680
rect 15338 2630 15446 2636
rect 15338 2596 15350 2630
rect 15434 2596 15446 2630
rect 15338 2590 15446 2596
rect 15236 2490 15246 2546
rect 15022 2170 15036 2194
rect 14564 2120 14672 2126
rect 14564 2086 14576 2120
rect 14660 2086 14672 2120
rect 14564 2080 14672 2086
rect 14822 2120 14930 2126
rect 14822 2086 14834 2120
rect 14918 2086 14930 2120
rect 14822 2080 14930 2086
rect 14976 1900 15036 2170
rect 15240 2170 15246 2490
rect 15280 2490 15296 2546
rect 15494 2546 15554 2680
rect 15280 2170 15286 2490
rect 15240 2158 15286 2170
rect 15494 2170 15504 2546
rect 15538 2170 15554 2546
rect 15080 2120 15188 2126
rect 15080 2086 15092 2120
rect 15176 2086 15188 2120
rect 15080 2080 15188 2086
rect 15338 2120 15446 2126
rect 15338 2086 15350 2120
rect 15434 2086 15446 2120
rect 15338 2080 15446 2086
rect 15106 2010 15166 2080
rect 15100 1950 15106 2010
rect 15166 1950 15172 2010
rect 15360 2008 15420 2080
rect 15494 2008 15554 2170
rect 16210 2546 16270 2680
rect 16334 2636 16394 2680
rect 16312 2630 16420 2636
rect 16312 2596 16324 2630
rect 16408 2596 16420 2630
rect 16312 2590 16420 2596
rect 16210 2170 16220 2546
rect 16254 2170 16270 2546
rect 16464 2546 16524 2796
rect 16848 2686 16854 2746
rect 16914 2686 16920 2746
rect 16854 2636 16914 2686
rect 16570 2630 16678 2636
rect 16570 2596 16582 2630
rect 16666 2596 16678 2630
rect 16570 2590 16678 2596
rect 16828 2630 16936 2636
rect 16828 2596 16840 2630
rect 16924 2596 16936 2630
rect 16828 2590 16936 2596
rect 16464 2502 16478 2546
rect 16210 2008 16270 2170
rect 16472 2170 16478 2502
rect 16512 2502 16524 2546
rect 16730 2546 16776 2558
rect 16512 2170 16518 2502
rect 16730 2196 16736 2546
rect 16472 2158 16518 2170
rect 16724 2170 16736 2196
rect 16770 2196 16776 2546
rect 16978 2546 17038 2912
rect 17490 2796 17496 2856
rect 17556 2796 17562 2856
rect 17102 2686 17108 2746
rect 17168 2686 17174 2746
rect 17108 2636 17168 2686
rect 17086 2630 17194 2636
rect 17086 2596 17098 2630
rect 17182 2596 17194 2630
rect 17086 2590 17194 2596
rect 17344 2630 17452 2636
rect 17344 2596 17356 2630
rect 17440 2596 17452 2630
rect 17344 2590 17452 2596
rect 16978 2506 16994 2546
rect 16988 2258 16994 2506
rect 16770 2170 16784 2196
rect 16312 2120 16420 2126
rect 16312 2086 16324 2120
rect 16408 2086 16420 2120
rect 16312 2080 16420 2086
rect 16570 2120 16678 2126
rect 16570 2086 16582 2120
rect 16666 2086 16678 2120
rect 16570 2080 16678 2086
rect 16336 2008 16396 2080
rect 16594 2016 16654 2080
rect 13934 1840 13940 1900
rect 14000 1840 14006 1900
rect 14454 1840 14460 1900
rect 14520 1840 14526 1900
rect 14970 1840 14976 1900
rect 15036 1840 15042 1900
rect 13428 1834 13488 1840
rect 15106 1778 15166 1950
rect 15360 1948 16396 2008
rect 16588 1956 16594 2016
rect 16654 1956 16660 2016
rect 15100 1718 15106 1778
rect 15166 1718 15172 1778
rect 12360 1594 12842 1654
rect 13212 1594 13218 1654
rect 13278 1594 13284 1654
rect 12360 1438 12420 1594
rect 12782 1528 12842 1594
rect 12618 1522 13026 1528
rect 12618 1488 12630 1522
rect 13014 1488 13026 1522
rect 12618 1482 13026 1488
rect 12360 1262 12376 1438
rect 12410 1262 12420 1438
rect 13218 1438 13278 1594
rect 13476 1522 13884 1528
rect 13476 1488 13488 1522
rect 13872 1488 13884 1522
rect 13476 1482 13884 1488
rect 14334 1522 14742 1528
rect 14334 1488 14346 1522
rect 14730 1488 14742 1522
rect 14334 1482 14742 1488
rect 15192 1522 15600 1528
rect 15192 1488 15204 1522
rect 15588 1488 15600 1522
rect 15192 1482 15600 1488
rect 13218 1400 13234 1438
rect 12360 1104 12420 1262
rect 13228 1262 13234 1400
rect 13268 1400 13278 1438
rect 14086 1438 14132 1450
rect 13268 1262 13274 1400
rect 14086 1342 14092 1438
rect 13228 1250 13274 1262
rect 14078 1262 14092 1342
rect 14126 1342 14132 1438
rect 14944 1438 14990 1450
rect 14126 1262 14138 1342
rect 14944 1312 14950 1438
rect 12618 1212 13026 1218
rect 12618 1178 12630 1212
rect 13014 1178 13026 1212
rect 12618 1172 13026 1178
rect 13476 1212 13884 1218
rect 13476 1178 13488 1212
rect 13872 1178 13884 1212
rect 13476 1172 13884 1178
rect 12784 1104 12844 1172
rect 13644 1110 13704 1172
rect 12360 1044 12844 1104
rect 13214 1050 13220 1110
rect 13280 1050 13704 1110
rect 12360 898 12420 1044
rect 12784 988 12844 1044
rect 12618 982 13026 988
rect 12618 948 12630 982
rect 13014 948 13026 982
rect 12618 942 13026 948
rect 12360 722 12376 898
rect 12410 722 12420 898
rect 13220 898 13280 1050
rect 13644 988 13704 1050
rect 13476 982 13884 988
rect 13476 948 13488 982
rect 13872 948 13884 982
rect 13476 942 13884 948
rect 13220 846 13234 898
rect 12360 574 12420 722
rect 13228 722 13234 846
rect 13268 846 13280 898
rect 14078 898 14138 1262
rect 14936 1262 14950 1312
rect 14984 1312 14990 1438
rect 15794 1438 15854 1948
rect 16724 1906 16784 2170
rect 16986 2170 16994 2258
rect 17028 2506 17038 2546
rect 17246 2546 17292 2558
rect 17028 2258 17034 2506
rect 17028 2170 17046 2258
rect 17246 2196 17252 2546
rect 16828 2120 16936 2126
rect 16828 2086 16840 2120
rect 16924 2086 16936 2120
rect 16828 2080 16936 2086
rect 16724 1654 16784 1846
rect 16986 1778 17046 2170
rect 17236 2170 17252 2196
rect 17286 2196 17292 2546
rect 17496 2546 17556 2796
rect 17874 2686 17880 2746
rect 17940 2686 17946 2746
rect 17880 2636 17940 2686
rect 17602 2630 17710 2636
rect 17602 2596 17614 2630
rect 17698 2596 17710 2630
rect 17602 2590 17710 2596
rect 17860 2630 17968 2636
rect 17860 2596 17872 2630
rect 17956 2596 17968 2630
rect 17860 2590 17968 2596
rect 17496 2492 17510 2546
rect 17286 2170 17296 2196
rect 17086 2120 17194 2126
rect 17086 2086 17098 2120
rect 17182 2086 17194 2120
rect 17086 2080 17194 2086
rect 17236 1906 17296 2170
rect 17504 2170 17510 2492
rect 17544 2492 17556 2546
rect 17762 2546 17808 2558
rect 17544 2170 17550 2492
rect 17762 2200 17768 2546
rect 17504 2158 17550 2170
rect 17756 2170 17768 2200
rect 17802 2200 17808 2546
rect 18014 2546 18074 2912
rect 18526 2796 18532 2856
rect 18592 2796 18598 2856
rect 18136 2686 18142 2746
rect 18202 2686 18208 2746
rect 18142 2636 18202 2686
rect 18118 2630 18226 2636
rect 18118 2596 18130 2630
rect 18214 2596 18226 2630
rect 18118 2590 18226 2596
rect 18376 2630 18484 2636
rect 18376 2596 18388 2630
rect 18472 2596 18484 2630
rect 18376 2590 18484 2596
rect 18014 2502 18026 2546
rect 17802 2170 17816 2200
rect 17344 2120 17452 2126
rect 17344 2086 17356 2120
rect 17440 2086 17452 2120
rect 17344 2080 17452 2086
rect 17602 2120 17710 2126
rect 17602 2086 17614 2120
rect 17698 2086 17710 2120
rect 17602 2080 17710 2086
rect 17370 2016 17430 2080
rect 17624 2016 17684 2080
rect 17364 1956 17370 2016
rect 17430 1956 17436 2016
rect 17618 1956 17624 2016
rect 17684 1956 17690 2016
rect 17756 1906 17816 2170
rect 18020 2170 18026 2502
rect 18060 2502 18074 2546
rect 18278 2546 18324 2558
rect 18060 2170 18066 2502
rect 18278 2200 18284 2546
rect 18020 2158 18066 2170
rect 18272 2170 18284 2200
rect 18318 2200 18324 2546
rect 18532 2546 18592 2796
rect 18658 2746 18718 3012
rect 18790 2746 18850 3012
rect 19506 2746 19566 3012
rect 19630 2746 19690 3012
rect 20268 2906 20274 2966
rect 20334 2906 20340 2966
rect 21304 2906 21310 2966
rect 21370 2906 21376 2966
rect 19754 2790 19760 2850
rect 19820 2790 19826 2850
rect 18658 2686 19690 2746
rect 18658 2636 18718 2686
rect 18634 2630 18742 2636
rect 18634 2596 18646 2630
rect 18730 2596 18742 2630
rect 18634 2590 18742 2596
rect 18532 2496 18542 2546
rect 18318 2170 18332 2200
rect 17860 2120 17968 2126
rect 17860 2086 17872 2120
rect 17956 2086 17968 2120
rect 17860 2080 17968 2086
rect 18118 2120 18226 2126
rect 18118 2086 18130 2120
rect 18214 2086 18226 2120
rect 18118 2080 18226 2086
rect 18272 1906 18332 2170
rect 18536 2170 18542 2496
rect 18576 2496 18592 2546
rect 18790 2546 18850 2686
rect 18576 2170 18582 2496
rect 18536 2158 18582 2170
rect 18790 2170 18800 2546
rect 18834 2170 18850 2546
rect 18376 2120 18484 2126
rect 18376 2086 18388 2120
rect 18472 2086 18484 2120
rect 18376 2080 18484 2086
rect 18634 2120 18742 2126
rect 18634 2086 18646 2120
rect 18730 2086 18742 2120
rect 18634 2080 18742 2086
rect 18402 2016 18462 2080
rect 18396 1956 18402 2016
rect 18462 1956 18468 2016
rect 18656 2014 18716 2080
rect 18790 2014 18850 2170
rect 19506 2546 19566 2686
rect 19630 2636 19690 2686
rect 19608 2630 19716 2636
rect 19608 2596 19620 2630
rect 19704 2596 19716 2630
rect 19608 2590 19716 2596
rect 19506 2170 19516 2546
rect 19550 2170 19566 2546
rect 19760 2546 19820 2790
rect 20144 2680 20150 2740
rect 20210 2680 20216 2740
rect 20150 2636 20210 2680
rect 19866 2630 19974 2636
rect 19866 2596 19878 2630
rect 19962 2596 19974 2630
rect 19866 2590 19974 2596
rect 20124 2630 20232 2636
rect 20124 2596 20136 2630
rect 20220 2596 20232 2630
rect 20124 2590 20232 2596
rect 19760 2496 19774 2546
rect 19506 2014 19566 2170
rect 19768 2170 19774 2496
rect 19808 2496 19820 2546
rect 20026 2546 20072 2558
rect 19808 2170 19814 2496
rect 20026 2190 20032 2546
rect 19768 2158 19814 2170
rect 20020 2170 20032 2190
rect 20066 2190 20072 2546
rect 20274 2546 20334 2906
rect 20786 2790 20792 2850
rect 20852 2790 20858 2850
rect 20398 2680 20404 2740
rect 20464 2680 20470 2740
rect 20404 2636 20464 2680
rect 20382 2630 20490 2636
rect 20382 2596 20394 2630
rect 20478 2596 20490 2630
rect 20382 2590 20490 2596
rect 20640 2630 20748 2636
rect 20640 2596 20652 2630
rect 20736 2596 20748 2630
rect 20640 2590 20748 2596
rect 20274 2500 20290 2546
rect 20066 2170 20080 2190
rect 19608 2120 19716 2126
rect 19608 2086 19620 2120
rect 19704 2086 19716 2120
rect 19608 2080 19716 2086
rect 19866 2120 19974 2126
rect 19866 2086 19878 2120
rect 19962 2086 19974 2120
rect 19866 2080 19974 2086
rect 19632 2014 19692 2080
rect 18656 1954 19692 2014
rect 19890 2010 19950 2080
rect 17230 1846 17236 1906
rect 17296 1846 17302 1906
rect 17750 1846 17756 1906
rect 17816 1846 17822 1906
rect 18266 1846 18272 1906
rect 18332 1846 18338 1906
rect 16980 1718 16986 1778
rect 17046 1718 17052 1778
rect 16646 1594 16652 1654
rect 16712 1594 16784 1654
rect 17082 1596 18006 1656
rect 16050 1522 16458 1528
rect 16050 1488 16062 1522
rect 16446 1488 16458 1522
rect 16050 1482 16458 1488
rect 14984 1262 14996 1312
rect 14334 1212 14742 1218
rect 14334 1178 14346 1212
rect 14730 1178 14742 1212
rect 14334 1172 14742 1178
rect 14502 1110 14562 1172
rect 14936 1110 14996 1262
rect 15794 1262 15808 1438
rect 15842 1262 15854 1438
rect 16652 1438 16712 1594
rect 17082 1528 17142 1596
rect 16908 1522 17316 1528
rect 16908 1488 16920 1522
rect 17304 1488 17316 1522
rect 16908 1482 17316 1488
rect 16652 1396 16666 1438
rect 15192 1212 15600 1218
rect 15192 1178 15204 1212
rect 15588 1178 15600 1212
rect 15192 1172 15600 1178
rect 15366 1110 15426 1172
rect 14496 1054 14502 1110
rect 14562 1054 14568 1110
rect 14496 1050 14568 1054
rect 14930 1050 14936 1110
rect 14996 1050 15002 1110
rect 14502 988 14562 1050
rect 14334 982 14742 988
rect 14334 948 14346 982
rect 14730 948 14742 982
rect 14334 942 14742 948
rect 13268 722 13274 846
rect 13228 710 13274 722
rect 14078 722 14092 898
rect 14126 722 14138 898
rect 14936 898 14996 1050
rect 15366 988 15426 1054
rect 15192 982 15600 988
rect 15192 948 15204 982
rect 15588 948 15600 982
rect 15192 942 15600 948
rect 14936 870 14950 898
rect 12618 672 13026 678
rect 12618 638 12630 672
rect 13014 638 13026 672
rect 12618 632 13026 638
rect 13476 672 13884 678
rect 13476 638 13488 672
rect 13872 638 13884 672
rect 13476 632 13884 638
rect 12780 574 12840 632
rect 12214 506 12220 566
rect 12280 506 12286 566
rect 12360 514 12840 574
rect 12360 400 12420 514
rect 12780 400 12840 514
rect 14078 400 14138 722
rect 14944 722 14950 870
rect 14984 870 14996 898
rect 15794 898 15854 1262
rect 16660 1262 16666 1396
rect 16700 1396 16712 1438
rect 17508 1438 17568 1596
rect 17946 1528 18006 1596
rect 17766 1522 18174 1528
rect 17766 1488 17778 1522
rect 18162 1488 18174 1522
rect 17766 1482 18174 1488
rect 18624 1522 19032 1528
rect 18624 1488 18636 1522
rect 19020 1488 19032 1522
rect 18624 1482 19032 1488
rect 16700 1262 16706 1396
rect 16660 1250 16706 1262
rect 17508 1262 17524 1438
rect 17558 1262 17568 1438
rect 18376 1438 18422 1450
rect 18376 1310 18382 1438
rect 16050 1212 16458 1218
rect 16050 1178 16062 1212
rect 16446 1178 16458 1212
rect 16050 1172 16458 1178
rect 16908 1212 17316 1218
rect 16908 1178 16920 1212
rect 17304 1178 17316 1212
rect 16908 1172 17316 1178
rect 16226 1110 16286 1172
rect 17084 1112 17144 1172
rect 17508 1112 17568 1262
rect 18372 1262 18382 1310
rect 18416 1310 18422 1438
rect 19226 1438 19286 1954
rect 19884 1950 19890 2010
rect 19950 1950 19956 2010
rect 20020 1900 20080 2170
rect 20284 2170 20290 2500
rect 20324 2500 20334 2546
rect 20542 2546 20588 2558
rect 20324 2170 20330 2500
rect 20542 2190 20548 2546
rect 20284 2158 20330 2170
rect 20532 2170 20548 2190
rect 20582 2190 20588 2546
rect 20792 2546 20852 2790
rect 21170 2680 21176 2740
rect 21236 2680 21242 2740
rect 21176 2636 21236 2680
rect 20898 2630 21006 2636
rect 20898 2596 20910 2630
rect 20994 2596 21006 2630
rect 20898 2590 21006 2596
rect 21156 2630 21264 2636
rect 21156 2596 21168 2630
rect 21252 2596 21264 2630
rect 21156 2590 21264 2596
rect 21176 2586 21236 2590
rect 20792 2486 20806 2546
rect 20582 2170 20592 2190
rect 20124 2120 20232 2126
rect 20124 2086 20136 2120
rect 20220 2086 20232 2120
rect 20124 2080 20232 2086
rect 20382 2120 20490 2126
rect 20382 2086 20394 2120
rect 20478 2086 20490 2120
rect 20382 2080 20490 2086
rect 20532 1900 20592 2170
rect 20800 2170 20806 2486
rect 20840 2486 20852 2546
rect 21058 2546 21104 2558
rect 20840 2170 20846 2486
rect 21058 2194 21064 2546
rect 20800 2158 20846 2170
rect 21052 2170 21064 2194
rect 21098 2194 21104 2546
rect 21310 2546 21370 2906
rect 21822 2790 21828 2850
rect 21888 2790 21894 2850
rect 21432 2680 21438 2740
rect 21498 2680 21504 2740
rect 21438 2636 21498 2680
rect 21414 2630 21522 2636
rect 21414 2596 21426 2630
rect 21510 2596 21522 2630
rect 21414 2590 21522 2596
rect 21672 2630 21780 2636
rect 21672 2596 21684 2630
rect 21768 2596 21780 2630
rect 21672 2590 21780 2596
rect 21310 2496 21322 2546
rect 21098 2170 21112 2194
rect 20640 2120 20748 2126
rect 20640 2086 20652 2120
rect 20736 2086 20748 2120
rect 20640 2080 20748 2086
rect 20898 2120 21006 2126
rect 20898 2086 20910 2120
rect 20994 2086 21006 2120
rect 20898 2080 21006 2086
rect 20666 2010 20726 2080
rect 20920 2010 20980 2080
rect 20660 1950 20666 2010
rect 20726 1950 20732 2010
rect 20914 1950 20920 2010
rect 20980 1950 20986 2010
rect 21052 1900 21112 2170
rect 21316 2170 21322 2496
rect 21356 2496 21370 2546
rect 21574 2546 21620 2558
rect 21356 2170 21362 2496
rect 21574 2194 21580 2546
rect 21316 2158 21362 2170
rect 21568 2170 21580 2194
rect 21614 2194 21620 2546
rect 21828 2546 21888 2790
rect 21954 2738 22014 3012
rect 22086 2738 22146 3012
rect 23104 2858 23216 3012
rect 23104 2738 23110 2858
rect 21954 2678 23110 2738
rect 21954 2636 22014 2678
rect 21930 2630 22038 2636
rect 21930 2596 21942 2630
rect 22026 2596 22038 2630
rect 21930 2590 22038 2596
rect 21828 2490 21838 2546
rect 21614 2170 21628 2194
rect 21156 2120 21264 2126
rect 21156 2086 21168 2120
rect 21252 2086 21264 2120
rect 21156 2080 21264 2086
rect 21414 2120 21522 2126
rect 21414 2086 21426 2120
rect 21510 2086 21522 2120
rect 21414 2080 21522 2086
rect 21568 1900 21628 2170
rect 21832 2170 21838 2490
rect 21872 2490 21888 2546
rect 22086 2546 22146 2678
rect 21872 2170 21878 2490
rect 21832 2158 21878 2170
rect 22086 2170 22096 2546
rect 22130 2170 22146 2546
rect 21672 2120 21780 2126
rect 21672 2086 21684 2120
rect 21768 2086 21780 2120
rect 21672 2080 21780 2086
rect 21930 2120 22038 2126
rect 21930 2086 21942 2120
rect 22026 2086 22038 2120
rect 21930 2080 22038 2086
rect 21698 2010 21758 2080
rect 21692 1950 21698 2010
rect 21758 1950 21764 2010
rect 21952 2008 22012 2080
rect 22086 2008 22146 2170
rect 23104 2008 23110 2678
rect 21952 1948 23110 2008
rect 20014 1840 20020 1900
rect 20080 1840 20086 1900
rect 20526 1840 20532 1900
rect 20592 1840 20598 1900
rect 21046 1840 21052 1900
rect 21112 1840 21118 1900
rect 21562 1840 21568 1900
rect 21628 1840 21634 1900
rect 21796 1710 21802 1770
rect 21862 1710 21868 1770
rect 19482 1522 19890 1528
rect 19482 1488 19494 1522
rect 19878 1488 19890 1522
rect 19482 1482 19890 1488
rect 20340 1522 20748 1528
rect 20340 1488 20352 1522
rect 20736 1488 20748 1522
rect 20340 1482 20748 1488
rect 21198 1522 21606 1528
rect 21198 1488 21210 1522
rect 21594 1488 21606 1522
rect 21198 1482 21606 1488
rect 18416 1262 18432 1310
rect 17766 1212 18174 1218
rect 17766 1178 17778 1212
rect 18162 1178 18174 1212
rect 17766 1172 18174 1178
rect 17944 1112 18004 1172
rect 16226 988 16286 1054
rect 16650 1050 16656 1110
rect 16716 1050 16722 1110
rect 17084 1052 18004 1112
rect 18372 1110 18432 1262
rect 19226 1262 19240 1438
rect 19274 1262 19286 1438
rect 20092 1438 20138 1450
rect 20092 1326 20098 1438
rect 18624 1212 19032 1218
rect 18624 1178 18636 1212
rect 19020 1178 19032 1212
rect 18624 1172 19032 1178
rect 18798 1110 18858 1172
rect 16050 982 16458 988
rect 16050 948 16062 982
rect 16446 948 16458 982
rect 16050 942 16458 948
rect 14984 722 14990 870
rect 14944 710 14990 722
rect 15794 722 15808 898
rect 15842 722 15854 898
rect 16656 898 16716 1050
rect 17084 988 17144 1052
rect 16908 982 17316 988
rect 16908 948 16920 982
rect 17304 948 17316 982
rect 16908 942 17316 948
rect 16656 846 16666 898
rect 14334 672 14742 678
rect 14334 638 14346 672
rect 14730 638 14742 672
rect 14334 632 14742 638
rect 15192 672 15600 678
rect 15192 638 15204 672
rect 15588 638 15600 672
rect 15192 632 15600 638
rect 15794 400 15854 722
rect 16660 722 16666 846
rect 16700 846 16716 898
rect 17508 898 17568 1052
rect 17944 988 18004 1052
rect 18366 1050 18372 1110
rect 18432 1050 18438 1110
rect 18792 1054 18798 1110
rect 18858 1054 18864 1110
rect 18792 1050 18864 1054
rect 18798 988 18858 1050
rect 17766 982 18174 988
rect 17766 948 17778 982
rect 18162 948 18174 982
rect 17766 942 18174 948
rect 18624 982 19032 988
rect 18624 948 18636 982
rect 19020 948 19032 982
rect 18624 942 19032 948
rect 16700 722 16706 846
rect 16660 710 16706 722
rect 17508 722 17524 898
rect 17558 722 17568 898
rect 18376 898 18422 910
rect 18376 752 18382 898
rect 16050 672 16458 678
rect 16050 638 16062 672
rect 16446 638 16458 672
rect 16050 632 16458 638
rect 16908 672 17316 678
rect 16908 638 16920 672
rect 17304 638 17316 672
rect 16908 632 17316 638
rect 17082 568 17142 632
rect 17508 568 17568 722
rect 18368 722 18382 752
rect 18416 752 18422 898
rect 19226 898 19286 1262
rect 20084 1262 20098 1326
rect 20132 1326 20138 1438
rect 20950 1438 20996 1450
rect 20132 1262 20144 1326
rect 20950 1318 20956 1438
rect 19482 1212 19890 1218
rect 19482 1178 19494 1212
rect 19878 1178 19890 1212
rect 19482 1172 19890 1178
rect 19656 1110 19716 1172
rect 20084 1110 20144 1262
rect 20944 1262 20956 1318
rect 20990 1318 20996 1438
rect 21802 1438 21862 1710
rect 22232 1640 22292 1948
rect 22656 1640 22716 1948
rect 22782 1840 22788 1900
rect 22848 1840 22854 1900
rect 22232 1580 22716 1640
rect 22232 1528 22292 1580
rect 22056 1522 22464 1528
rect 22056 1488 22068 1522
rect 22452 1488 22464 1522
rect 22056 1482 22464 1488
rect 21802 1404 21814 1438
rect 20990 1262 21004 1318
rect 20340 1212 20748 1218
rect 20340 1178 20352 1212
rect 20736 1178 20748 1212
rect 20340 1172 20748 1178
rect 20510 1110 20570 1172
rect 19656 988 19716 1054
rect 20078 1050 20084 1110
rect 20144 1050 20150 1110
rect 19482 982 19890 988
rect 19482 948 19494 982
rect 19878 948 19890 982
rect 19482 942 19890 948
rect 18416 722 18428 752
rect 17766 672 18174 678
rect 17766 638 17778 672
rect 18162 638 18174 672
rect 17766 632 18174 638
rect 17944 568 18004 632
rect 17082 508 18004 568
rect 18368 566 18428 722
rect 19226 722 19240 898
rect 19274 722 19286 898
rect 20084 898 20144 1050
rect 20510 988 20570 1054
rect 20340 982 20748 988
rect 20340 948 20352 982
rect 20736 948 20748 982
rect 20340 942 20748 948
rect 20084 856 20098 898
rect 18624 672 19032 678
rect 18624 638 18636 672
rect 19020 638 19032 672
rect 18624 632 19032 638
rect 17082 400 17142 508
rect 17508 400 17568 508
rect 17944 400 18004 508
rect 18362 506 18368 566
rect 18428 506 18434 566
rect 19226 400 19286 722
rect 20092 722 20098 856
rect 20132 856 20144 898
rect 20944 898 21004 1262
rect 21808 1262 21814 1404
rect 21848 1404 21862 1438
rect 22656 1438 22716 1580
rect 21848 1262 21854 1404
rect 21808 1250 21854 1262
rect 22656 1262 22672 1438
rect 22706 1262 22716 1438
rect 21198 1212 21606 1218
rect 21198 1178 21210 1212
rect 21594 1178 21606 1212
rect 21198 1172 21606 1178
rect 22056 1212 22464 1218
rect 22056 1178 22068 1212
rect 22452 1178 22464 1212
rect 22056 1172 22464 1178
rect 21374 1116 21434 1172
rect 21374 1110 21436 1116
rect 21374 1050 21376 1110
rect 21374 1044 21436 1050
rect 22230 1106 22290 1172
rect 22656 1106 22716 1262
rect 22230 1046 22716 1106
rect 21374 988 21434 1044
rect 22230 988 22290 1046
rect 21198 982 21606 988
rect 21198 948 21210 982
rect 21594 948 21606 982
rect 21198 942 21606 948
rect 22056 982 22464 988
rect 22056 948 22068 982
rect 22452 948 22464 982
rect 22056 942 22464 948
rect 20132 722 20138 856
rect 20092 710 20138 722
rect 20944 722 20956 898
rect 20990 722 21004 898
rect 21808 898 21854 910
rect 21808 754 21814 898
rect 19482 672 19890 678
rect 19482 638 19494 672
rect 19878 638 19890 672
rect 19482 632 19890 638
rect 20340 672 20748 678
rect 20340 638 20352 672
rect 20736 638 20748 672
rect 20340 632 20748 638
rect 20944 400 21004 722
rect 21800 722 21814 754
rect 21848 754 21854 898
rect 22656 898 22716 1046
rect 21848 722 21860 754
rect 21198 672 21606 678
rect 21198 638 21210 672
rect 21594 638 21606 672
rect 21198 632 21606 638
rect 21800 572 21860 722
rect 22656 722 22672 898
rect 22706 722 22716 898
rect 22056 672 22464 678
rect 22056 638 22068 672
rect 22452 638 22464 672
rect 22056 632 22464 638
rect 22232 572 22292 632
rect 22656 572 22716 722
rect 22788 572 22848 1840
rect 21794 512 21800 572
rect 21860 512 21866 572
rect 22232 512 22716 572
rect 22782 512 22788 572
rect 22848 512 22854 572
rect 22232 400 22292 512
rect 22656 400 22716 512
rect 12122 352 22896 400
rect 12122 242 12184 352
rect 22840 242 22896 352
rect 12122 186 22896 242
rect 11860 -180 11972 -26
rect 12572 -180 12582 120
rect 22494 -180 22504 120
rect 23104 -26 23110 1948
rect 23210 -26 23216 2858
rect 23104 -180 23216 -26
rect 11860 -186 23216 -180
rect 11860 -286 11966 -186
rect 23110 -286 23216 -186
rect 11860 -292 23216 -286
rect 60 -518 11416 -512
rect 60 -618 166 -518
rect 11310 -618 11416 -518
rect 60 -624 11416 -618
rect 60 -778 172 -624
rect 60 -3662 66 -778
rect 166 -2752 172 -778
rect 772 -924 782 -624
rect 10694 -924 10704 -624
rect 11304 -778 11416 -624
rect 322 -1046 11096 -990
rect 322 -1156 384 -1046
rect 11040 -1156 11096 -1046
rect 322 -1204 11096 -1156
rect 414 -1370 420 -1310
rect 480 -1370 486 -1310
rect 560 -1318 620 -1204
rect 980 -1318 1040 -1204
rect 420 -2644 480 -1370
rect 560 -1378 1040 -1318
rect 560 -1526 620 -1378
rect 980 -1436 1040 -1378
rect 818 -1442 1226 -1436
rect 818 -1476 830 -1442
rect 1214 -1476 1226 -1442
rect 818 -1482 1226 -1476
rect 1676 -1442 2084 -1436
rect 1676 -1476 1688 -1442
rect 2072 -1476 2084 -1442
rect 1676 -1482 2084 -1476
rect 560 -1702 576 -1526
rect 610 -1702 620 -1526
rect 1428 -1526 1474 -1514
rect 1428 -1650 1434 -1526
rect 560 -1848 620 -1702
rect 1420 -1702 1434 -1650
rect 1468 -1650 1474 -1526
rect 2278 -1526 2338 -1204
rect 2534 -1442 2942 -1436
rect 2534 -1476 2546 -1442
rect 2930 -1476 2942 -1442
rect 2534 -1482 2942 -1476
rect 3392 -1442 3800 -1436
rect 3392 -1476 3404 -1442
rect 3788 -1476 3800 -1442
rect 3392 -1482 3800 -1476
rect 1468 -1702 1480 -1650
rect 818 -1752 1226 -1746
rect 818 -1786 830 -1752
rect 1214 -1786 1226 -1752
rect 818 -1792 1226 -1786
rect 984 -1848 1044 -1792
rect 560 -1908 1044 -1848
rect 1420 -1854 1480 -1702
rect 2278 -1702 2292 -1526
rect 2326 -1702 2338 -1526
rect 3144 -1526 3190 -1514
rect 3144 -1674 3150 -1526
rect 1676 -1752 2084 -1746
rect 1676 -1786 1688 -1752
rect 2072 -1786 2084 -1752
rect 1676 -1792 2084 -1786
rect 1844 -1854 1904 -1792
rect 560 -2066 620 -1908
rect 984 -1976 1044 -1908
rect 1414 -1914 1420 -1854
rect 1480 -1914 1904 -1854
rect 1844 -1976 1904 -1914
rect 818 -1982 1226 -1976
rect 818 -2016 830 -1982
rect 1214 -2016 1226 -1982
rect 818 -2022 1226 -2016
rect 1676 -1982 2084 -1976
rect 1676 -2016 1688 -1982
rect 2072 -2016 2084 -1982
rect 1676 -2022 2084 -2016
rect 560 -2242 576 -2066
rect 610 -2242 620 -2066
rect 1428 -2066 1474 -2054
rect 1428 -2204 1434 -2066
rect 560 -2398 620 -2242
rect 1418 -2242 1434 -2204
rect 1468 -2204 1474 -2066
rect 2278 -2066 2338 -1702
rect 3136 -1702 3150 -1674
rect 3184 -1674 3190 -1526
rect 3994 -1526 4054 -1204
rect 5282 -1312 5342 -1204
rect 5708 -1312 5768 -1204
rect 6144 -1312 6204 -1204
rect 5282 -1372 6204 -1312
rect 6562 -1370 6568 -1310
rect 6628 -1370 6634 -1310
rect 5282 -1436 5342 -1372
rect 4250 -1442 4658 -1436
rect 4250 -1476 4262 -1442
rect 4646 -1476 4658 -1442
rect 4250 -1482 4658 -1476
rect 5108 -1442 5516 -1436
rect 5108 -1476 5120 -1442
rect 5504 -1476 5516 -1442
rect 5108 -1482 5516 -1476
rect 3184 -1702 3196 -1674
rect 2534 -1752 2942 -1746
rect 2534 -1786 2546 -1752
rect 2930 -1786 2942 -1752
rect 2534 -1792 2942 -1786
rect 2702 -1854 2762 -1792
rect 3136 -1854 3196 -1702
rect 3994 -1702 4008 -1526
rect 4042 -1702 4054 -1526
rect 4860 -1526 4906 -1514
rect 4860 -1650 4866 -1526
rect 3392 -1752 3800 -1746
rect 3392 -1786 3404 -1752
rect 3788 -1786 3800 -1752
rect 3392 -1792 3800 -1786
rect 2696 -1858 2768 -1854
rect 2696 -1914 2702 -1858
rect 2762 -1914 2768 -1858
rect 3130 -1914 3136 -1854
rect 3196 -1914 3202 -1854
rect 3566 -1858 3626 -1792
rect 2702 -1976 2762 -1914
rect 2534 -1982 2942 -1976
rect 2534 -2016 2546 -1982
rect 2930 -2016 2942 -1982
rect 2534 -2022 2942 -2016
rect 2278 -2146 2292 -2066
rect 1468 -2242 1478 -2204
rect 818 -2292 1226 -2286
rect 818 -2326 830 -2292
rect 1214 -2326 1226 -2292
rect 818 -2332 1226 -2326
rect 982 -2398 1042 -2332
rect 1418 -2398 1478 -2242
rect 2286 -2242 2292 -2146
rect 2326 -2146 2338 -2066
rect 3136 -2066 3196 -1914
rect 3566 -1976 3626 -1914
rect 3392 -1982 3800 -1976
rect 3392 -2016 3404 -1982
rect 3788 -2016 3800 -1982
rect 3392 -2022 3800 -2016
rect 3136 -2116 3150 -2066
rect 2326 -2242 2332 -2146
rect 2286 -2254 2332 -2242
rect 3144 -2242 3150 -2116
rect 3184 -2116 3196 -2066
rect 3994 -2066 4054 -1702
rect 4856 -1702 4866 -1650
rect 4900 -1650 4906 -1526
rect 5708 -1526 5768 -1372
rect 6144 -1436 6204 -1372
rect 5966 -1442 6374 -1436
rect 5966 -1476 5978 -1442
rect 6362 -1476 6374 -1442
rect 5966 -1482 6374 -1476
rect 4900 -1702 4916 -1650
rect 4250 -1752 4658 -1746
rect 4250 -1786 4262 -1752
rect 4646 -1786 4658 -1752
rect 4250 -1792 4658 -1786
rect 4426 -1858 4486 -1792
rect 4856 -1854 4916 -1702
rect 5708 -1702 5724 -1526
rect 5758 -1702 5768 -1526
rect 6568 -1526 6628 -1370
rect 6824 -1442 7232 -1436
rect 6824 -1476 6836 -1442
rect 7220 -1476 7232 -1442
rect 6824 -1482 7232 -1476
rect 6568 -1556 6582 -1526
rect 5108 -1752 5516 -1746
rect 5108 -1786 5120 -1752
rect 5504 -1786 5516 -1752
rect 5108 -1792 5516 -1786
rect 4850 -1914 4856 -1854
rect 4916 -1914 4922 -1854
rect 5284 -1856 5344 -1792
rect 5708 -1856 5768 -1702
rect 6576 -1702 6582 -1556
rect 6616 -1556 6628 -1526
rect 7426 -1526 7486 -1204
rect 7682 -1442 8090 -1436
rect 7682 -1476 7694 -1442
rect 8078 -1476 8090 -1442
rect 7682 -1482 8090 -1476
rect 8540 -1442 8948 -1436
rect 8540 -1476 8552 -1442
rect 8936 -1476 8948 -1442
rect 8540 -1482 8948 -1476
rect 6616 -1702 6622 -1556
rect 6576 -1714 6622 -1702
rect 7426 -1702 7440 -1526
rect 7474 -1702 7486 -1526
rect 8292 -1526 8338 -1514
rect 8292 -1660 8298 -1526
rect 5966 -1752 6374 -1746
rect 5966 -1786 5978 -1752
rect 6362 -1786 6374 -1752
rect 5966 -1792 6374 -1786
rect 6824 -1752 7232 -1746
rect 6824 -1786 6836 -1752
rect 7220 -1786 7232 -1752
rect 6824 -1792 7232 -1786
rect 6144 -1856 6204 -1792
rect 6998 -1854 7058 -1792
rect 4426 -1976 4486 -1914
rect 5284 -1916 6204 -1856
rect 6566 -1914 6572 -1854
rect 6632 -1914 6638 -1854
rect 6992 -1858 7064 -1854
rect 6992 -1914 6998 -1858
rect 7058 -1914 7064 -1858
rect 5284 -1976 5344 -1916
rect 4250 -1982 4658 -1976
rect 4250 -2016 4262 -1982
rect 4646 -2016 4658 -1982
rect 4250 -2022 4658 -2016
rect 5108 -1982 5516 -1976
rect 5108 -2016 5120 -1982
rect 5504 -2016 5516 -1982
rect 5108 -2022 5516 -2016
rect 3184 -2242 3190 -2116
rect 3144 -2254 3190 -2242
rect 3994 -2242 4008 -2066
rect 4042 -2242 4054 -2066
rect 4860 -2066 4906 -2054
rect 4860 -2200 4866 -2066
rect 1676 -2292 2084 -2286
rect 1676 -2326 1688 -2292
rect 2072 -2326 2084 -2292
rect 1676 -2332 2084 -2326
rect 2534 -2292 2942 -2286
rect 2534 -2326 2546 -2292
rect 2930 -2326 2942 -2292
rect 2534 -2332 2942 -2326
rect 3392 -2292 3800 -2286
rect 3392 -2326 3404 -2292
rect 3788 -2326 3800 -2292
rect 3392 -2332 3800 -2326
rect 560 -2458 1042 -2398
rect 1412 -2458 1418 -2398
rect 1478 -2458 1484 -2398
rect 414 -2704 420 -2644
rect 480 -2704 486 -2644
rect 560 -2752 620 -2458
rect 3300 -2582 3306 -2522
rect 3366 -2582 3372 -2522
rect 1628 -2644 1688 -2638
rect 2134 -2704 2140 -2644
rect 2200 -2704 2206 -2644
rect 2654 -2704 2660 -2644
rect 2720 -2704 2726 -2644
rect 3170 -2704 3176 -2644
rect 3236 -2704 3242 -2644
rect 166 -2812 1300 -2752
rect 166 -3484 172 -2812
rect 1114 -2974 1174 -2812
rect 1240 -2884 1300 -2812
rect 1492 -2814 1498 -2754
rect 1558 -2814 1564 -2754
rect 1498 -2884 1558 -2814
rect 1216 -2890 1324 -2884
rect 1216 -2924 1228 -2890
rect 1312 -2924 1324 -2890
rect 1216 -2930 1324 -2924
rect 1474 -2890 1582 -2884
rect 1474 -2924 1486 -2890
rect 1570 -2924 1582 -2890
rect 1474 -2930 1582 -2924
rect 1114 -3350 1124 -2974
rect 1158 -3350 1174 -2974
rect 1376 -2974 1422 -2962
rect 1376 -3300 1382 -2974
rect 1114 -3484 1174 -3350
rect 1368 -3350 1382 -3300
rect 1416 -3300 1422 -2974
rect 1628 -2974 1688 -2704
rect 1732 -2890 1840 -2884
rect 1732 -2924 1744 -2890
rect 1828 -2924 1840 -2890
rect 1732 -2930 1840 -2924
rect 1990 -2890 2098 -2884
rect 1990 -2924 2002 -2890
rect 2086 -2924 2098 -2890
rect 1990 -2930 2098 -2924
rect 1628 -2994 1640 -2974
rect 1416 -3350 1428 -3300
rect 1216 -3400 1324 -3394
rect 1216 -3434 1228 -3400
rect 1312 -3434 1324 -3400
rect 1216 -3440 1324 -3434
rect 1240 -3484 1300 -3440
rect 166 -3544 1300 -3484
rect 166 -3662 172 -3544
rect 60 -3816 172 -3662
rect 1114 -3816 1174 -3544
rect 1240 -3816 1300 -3544
rect 1368 -3594 1428 -3350
rect 1634 -3350 1640 -2994
rect 1674 -2994 1688 -2974
rect 1892 -2974 1938 -2962
rect 1674 -3350 1680 -2994
rect 1892 -3304 1898 -2974
rect 1634 -3362 1680 -3350
rect 1882 -3350 1898 -3304
rect 1932 -3304 1938 -2974
rect 2140 -2974 2200 -2704
rect 2268 -2814 2274 -2754
rect 2334 -2814 2340 -2754
rect 2522 -2814 2528 -2754
rect 2588 -2814 2594 -2754
rect 2274 -2884 2334 -2814
rect 2528 -2884 2588 -2814
rect 2248 -2890 2356 -2884
rect 2248 -2924 2260 -2890
rect 2344 -2924 2356 -2890
rect 2248 -2930 2356 -2924
rect 2506 -2890 2614 -2884
rect 2506 -2924 2518 -2890
rect 2602 -2924 2614 -2890
rect 2506 -2930 2614 -2924
rect 2140 -2994 2156 -2974
rect 1932 -3350 1942 -3304
rect 1474 -3400 1582 -3394
rect 1474 -3434 1486 -3400
rect 1570 -3434 1582 -3400
rect 1474 -3440 1582 -3434
rect 1732 -3400 1840 -3394
rect 1732 -3434 1744 -3400
rect 1828 -3434 1840 -3400
rect 1732 -3440 1840 -3434
rect 1758 -3484 1818 -3440
rect 1752 -3544 1758 -3484
rect 1818 -3544 1824 -3484
rect 1362 -3654 1368 -3594
rect 1428 -3654 1434 -3594
rect 1882 -3710 1942 -3350
rect 2150 -3350 2156 -2994
rect 2190 -2994 2200 -2974
rect 2408 -2974 2454 -2962
rect 2190 -3350 2196 -2994
rect 2408 -3290 2414 -2974
rect 2150 -3362 2196 -3350
rect 2400 -3350 2414 -3290
rect 2448 -3290 2454 -2974
rect 2660 -2974 2720 -2704
rect 2764 -2890 2872 -2884
rect 2764 -2924 2776 -2890
rect 2860 -2924 2872 -2890
rect 2764 -2930 2872 -2924
rect 3022 -2890 3130 -2884
rect 3022 -2924 3034 -2890
rect 3118 -2924 3130 -2890
rect 3022 -2930 3130 -2924
rect 2660 -2998 2672 -2974
rect 2448 -3350 2460 -3290
rect 1990 -3400 2098 -3394
rect 1990 -3434 2002 -3400
rect 2086 -3434 2098 -3400
rect 1990 -3440 2098 -3434
rect 2248 -3400 2356 -3394
rect 2248 -3434 2260 -3400
rect 2344 -3434 2356 -3400
rect 2248 -3440 2356 -3434
rect 2012 -3484 2072 -3440
rect 2006 -3544 2012 -3484
rect 2072 -3544 2078 -3484
rect 2400 -3594 2460 -3350
rect 2666 -3350 2672 -2998
rect 2706 -2998 2720 -2974
rect 2924 -2974 2970 -2962
rect 2706 -3350 2712 -2998
rect 2924 -3300 2930 -2974
rect 2666 -3362 2712 -3350
rect 2918 -3350 2930 -3300
rect 2964 -3300 2970 -2974
rect 3176 -2974 3236 -2704
rect 3306 -2754 3366 -2582
rect 3994 -2752 4054 -2242
rect 4852 -2242 4866 -2200
rect 4900 -2200 4906 -2066
rect 5708 -2066 5768 -1916
rect 6144 -1976 6204 -1916
rect 5966 -1982 6374 -1976
rect 5966 -2016 5978 -1982
rect 6362 -2016 6374 -1982
rect 5966 -2022 6374 -2016
rect 4900 -2242 4912 -2200
rect 4250 -2292 4658 -2286
rect 4250 -2326 4262 -2292
rect 4646 -2326 4658 -2292
rect 4250 -2332 4658 -2326
rect 4852 -2398 4912 -2242
rect 5708 -2242 5724 -2066
rect 5758 -2242 5768 -2066
rect 6572 -2066 6632 -1914
rect 6998 -1976 7058 -1914
rect 6824 -1982 7232 -1976
rect 6824 -2016 6836 -1982
rect 7220 -2016 7232 -1982
rect 6824 -2022 7232 -2016
rect 6572 -2114 6582 -2066
rect 5108 -2292 5516 -2286
rect 5108 -2326 5120 -2292
rect 5504 -2326 5516 -2292
rect 5108 -2332 5516 -2326
rect 4846 -2458 4852 -2398
rect 4912 -2458 4984 -2398
rect 4924 -2650 4984 -2458
rect 5282 -2400 5342 -2332
rect 5708 -2400 5768 -2242
rect 6576 -2242 6582 -2114
rect 6616 -2114 6632 -2066
rect 7426 -2066 7486 -1702
rect 8284 -1702 8298 -1660
rect 8332 -1660 8338 -1526
rect 9144 -1526 9204 -1204
rect 10432 -1316 10492 -1204
rect 10856 -1316 10916 -1204
rect 9994 -1376 10000 -1316
rect 10060 -1376 10066 -1316
rect 10432 -1376 10916 -1316
rect 10982 -1376 10988 -1316
rect 11048 -1376 11054 -1316
rect 9398 -1442 9806 -1436
rect 9398 -1476 9410 -1442
rect 9794 -1476 9806 -1442
rect 9398 -1482 9806 -1476
rect 8332 -1702 8344 -1660
rect 7682 -1752 8090 -1746
rect 7682 -1786 7694 -1752
rect 8078 -1786 8090 -1752
rect 7682 -1792 8090 -1786
rect 7856 -1858 7916 -1792
rect 8284 -1854 8344 -1702
rect 9144 -1702 9156 -1526
rect 9190 -1702 9204 -1526
rect 10000 -1526 10060 -1376
rect 10432 -1436 10492 -1376
rect 10256 -1442 10664 -1436
rect 10256 -1476 10268 -1442
rect 10652 -1476 10664 -1442
rect 10256 -1482 10664 -1476
rect 10000 -1558 10014 -1526
rect 8540 -1752 8948 -1746
rect 8540 -1786 8552 -1752
rect 8936 -1786 8948 -1752
rect 8540 -1792 8948 -1786
rect 8278 -1914 8284 -1854
rect 8344 -1914 8350 -1854
rect 8710 -1858 8770 -1792
rect 7856 -1976 7916 -1914
rect 7682 -1982 8090 -1976
rect 7682 -2016 7694 -1982
rect 8078 -2016 8090 -1982
rect 7682 -2022 8090 -2016
rect 6616 -2242 6622 -2114
rect 6576 -2254 6622 -2242
rect 7426 -2242 7440 -2066
rect 7474 -2242 7486 -2066
rect 8284 -2066 8344 -1914
rect 8710 -1976 8770 -1914
rect 8540 -1982 8948 -1976
rect 8540 -2016 8552 -1982
rect 8936 -2016 8948 -1982
rect 8540 -2022 8948 -2016
rect 8284 -2130 8298 -2066
rect 5966 -2292 6374 -2286
rect 5966 -2326 5978 -2292
rect 6362 -2326 6374 -2292
rect 5966 -2332 6374 -2326
rect 6824 -2292 7232 -2286
rect 6824 -2326 6836 -2292
rect 7220 -2326 7232 -2292
rect 6824 -2332 7232 -2326
rect 6146 -2400 6206 -2332
rect 5282 -2460 6206 -2400
rect 5180 -2582 5186 -2522
rect 5246 -2582 5252 -2522
rect 3300 -2814 3306 -2754
rect 3366 -2814 3372 -2754
rect 3560 -2812 4596 -2752
rect 3306 -2884 3366 -2814
rect 3560 -2884 3620 -2812
rect 3280 -2890 3388 -2884
rect 3280 -2924 3292 -2890
rect 3376 -2924 3388 -2890
rect 3280 -2930 3388 -2924
rect 3538 -2890 3646 -2884
rect 3538 -2924 3550 -2890
rect 3634 -2924 3646 -2890
rect 3538 -2930 3646 -2924
rect 3176 -2998 3188 -2974
rect 2964 -3350 2978 -3300
rect 2784 -3394 2844 -3390
rect 2506 -3400 2614 -3394
rect 2506 -3434 2518 -3400
rect 2602 -3434 2614 -3400
rect 2506 -3440 2614 -3434
rect 2764 -3400 2872 -3394
rect 2764 -3434 2776 -3400
rect 2860 -3434 2872 -3400
rect 2764 -3440 2872 -3434
rect 2784 -3484 2844 -3440
rect 2778 -3544 2784 -3484
rect 2844 -3544 2850 -3484
rect 2394 -3654 2400 -3594
rect 2460 -3654 2466 -3594
rect 2918 -3710 2978 -3350
rect 3182 -3350 3188 -2998
rect 3222 -2998 3236 -2974
rect 3440 -2974 3486 -2962
rect 3222 -3350 3228 -2998
rect 3440 -3294 3446 -2974
rect 3182 -3362 3228 -3350
rect 3436 -3350 3446 -3294
rect 3480 -3294 3486 -2974
rect 3694 -2974 3754 -2812
rect 3480 -3350 3496 -3294
rect 3022 -3400 3130 -3394
rect 3022 -3434 3034 -3400
rect 3118 -3434 3130 -3400
rect 3022 -3440 3130 -3434
rect 3280 -3400 3388 -3394
rect 3280 -3434 3292 -3400
rect 3376 -3434 3388 -3400
rect 3280 -3440 3388 -3434
rect 3046 -3484 3106 -3440
rect 3040 -3544 3046 -3484
rect 3106 -3544 3112 -3484
rect 3436 -3594 3496 -3350
rect 3694 -3350 3704 -2974
rect 3738 -3350 3754 -2974
rect 3538 -3400 3646 -3394
rect 3538 -3434 3550 -3400
rect 3634 -3434 3646 -3400
rect 3538 -3440 3646 -3434
rect 3560 -3484 3620 -3440
rect 3694 -3484 3754 -3350
rect 4410 -2974 4470 -2812
rect 4536 -2884 4596 -2812
rect 4664 -2760 4724 -2754
rect 4788 -2820 4794 -2760
rect 4854 -2820 4860 -2760
rect 4512 -2890 4620 -2884
rect 4512 -2924 4524 -2890
rect 4608 -2924 4620 -2890
rect 4512 -2930 4620 -2924
rect 4410 -3350 4420 -2974
rect 4454 -3350 4470 -2974
rect 4410 -3484 4470 -3350
rect 4664 -2974 4724 -2820
rect 4794 -2884 4854 -2820
rect 4770 -2890 4878 -2884
rect 4770 -2924 4782 -2890
rect 4866 -2924 4878 -2890
rect 4770 -2930 4878 -2924
rect 4664 -3350 4678 -2974
rect 4712 -3350 4724 -2974
rect 4924 -2974 4984 -2710
rect 5028 -2890 5136 -2884
rect 5028 -2924 5040 -2890
rect 5124 -2924 5136 -2890
rect 5028 -2930 5136 -2924
rect 4924 -3000 4936 -2974
rect 4512 -3400 4620 -3394
rect 4512 -3434 4524 -3400
rect 4608 -3434 4620 -3400
rect 4512 -3440 4620 -3434
rect 4534 -3484 4594 -3440
rect 3560 -3544 4594 -3484
rect 3430 -3654 3436 -3594
rect 3496 -3654 3502 -3594
rect 1876 -3770 1882 -3710
rect 1942 -3770 1948 -3710
rect 2912 -3770 2918 -3710
rect 2978 -3770 2984 -3710
rect 3560 -3816 3620 -3544
rect 3694 -3816 3754 -3544
rect 4410 -3816 4470 -3544
rect 4534 -3816 4594 -3544
rect 4664 -3600 4724 -3350
rect 4930 -3350 4936 -3000
rect 4970 -3000 4984 -2974
rect 5186 -2974 5246 -2582
rect 5430 -2710 5436 -2650
rect 5496 -2710 5502 -2650
rect 5950 -2710 5956 -2650
rect 6016 -2710 6022 -2650
rect 6466 -2710 6472 -2650
rect 6532 -2710 6538 -2650
rect 5286 -2890 5394 -2884
rect 5286 -2924 5298 -2890
rect 5382 -2924 5394 -2890
rect 5286 -2930 5394 -2924
rect 4970 -3350 4976 -3000
rect 5186 -3062 5194 -2974
rect 5188 -3310 5194 -3062
rect 4930 -3362 4976 -3350
rect 5178 -3350 5194 -3310
rect 5228 -3062 5246 -2974
rect 5436 -2974 5496 -2710
rect 5564 -2820 5570 -2760
rect 5630 -2820 5636 -2760
rect 5570 -2884 5630 -2820
rect 5690 -2822 5696 -2762
rect 5756 -2822 5762 -2762
rect 5818 -2820 5824 -2760
rect 5884 -2820 5890 -2760
rect 5544 -2890 5652 -2884
rect 5544 -2924 5556 -2890
rect 5640 -2924 5652 -2890
rect 5544 -2930 5652 -2924
rect 5436 -3000 5452 -2974
rect 5228 -3310 5234 -3062
rect 5228 -3350 5238 -3310
rect 4770 -3400 4878 -3394
rect 4770 -3434 4782 -3400
rect 4866 -3434 4878 -3400
rect 4770 -3440 4878 -3434
rect 5028 -3400 5136 -3394
rect 5028 -3434 5040 -3400
rect 5124 -3434 5136 -3400
rect 5028 -3440 5136 -3434
rect 5052 -3490 5114 -3440
rect 5048 -3550 5054 -3490
rect 5114 -3550 5120 -3490
rect 4658 -3660 4664 -3600
rect 4724 -3660 4730 -3600
rect 5052 -3716 5112 -3550
rect 5178 -3716 5238 -3350
rect 5446 -3350 5452 -3000
rect 5486 -3000 5496 -2974
rect 5696 -2974 5756 -2822
rect 5824 -2884 5884 -2820
rect 5802 -2890 5910 -2884
rect 5802 -2924 5814 -2890
rect 5898 -2924 5910 -2890
rect 5802 -2930 5910 -2924
rect 5486 -3350 5492 -3000
rect 5446 -3362 5492 -3350
rect 5696 -3350 5710 -2974
rect 5744 -3350 5756 -2974
rect 5956 -2974 6016 -2710
rect 6060 -2890 6168 -2884
rect 6060 -2924 6072 -2890
rect 6156 -2924 6168 -2890
rect 6060 -2930 6168 -2924
rect 6318 -2890 6426 -2884
rect 6318 -2924 6330 -2890
rect 6414 -2924 6426 -2890
rect 6318 -2930 6426 -2924
rect 5956 -3004 5968 -2974
rect 5286 -3400 5394 -3394
rect 5286 -3434 5298 -3400
rect 5382 -3434 5394 -3400
rect 5286 -3440 5394 -3434
rect 5544 -3400 5652 -3394
rect 5544 -3434 5556 -3400
rect 5640 -3434 5652 -3400
rect 5544 -3440 5652 -3434
rect 5308 -3490 5368 -3440
rect 5302 -3550 5308 -3490
rect 5368 -3550 5374 -3490
rect 5308 -3716 5368 -3550
rect 5696 -3600 5756 -3350
rect 5962 -3350 5968 -3004
rect 6002 -3004 6016 -2974
rect 6220 -2974 6266 -2962
rect 6002 -3350 6008 -3004
rect 6220 -3306 6226 -2974
rect 5962 -3362 6008 -3350
rect 6214 -3350 6226 -3306
rect 6260 -3306 6266 -2974
rect 6472 -2974 6532 -2710
rect 7426 -2758 7486 -2242
rect 8292 -2242 8298 -2130
rect 8332 -2130 8344 -2066
rect 9144 -2066 9204 -1702
rect 10008 -1702 10014 -1558
rect 10048 -1558 10060 -1526
rect 10856 -1526 10916 -1376
rect 10048 -1702 10054 -1558
rect 10008 -1714 10054 -1702
rect 10856 -1702 10872 -1526
rect 10906 -1702 10916 -1526
rect 9398 -1752 9806 -1746
rect 9398 -1786 9410 -1752
rect 9794 -1786 9806 -1752
rect 9398 -1792 9806 -1786
rect 10256 -1752 10664 -1746
rect 10256 -1786 10268 -1752
rect 10652 -1786 10664 -1752
rect 10256 -1792 10664 -1786
rect 9574 -1848 9634 -1792
rect 9574 -1854 9636 -1848
rect 9574 -1914 9576 -1854
rect 9574 -1920 9636 -1914
rect 10430 -1850 10490 -1792
rect 10856 -1850 10916 -1702
rect 10430 -1910 10916 -1850
rect 9574 -1976 9634 -1920
rect 10430 -1976 10490 -1910
rect 9398 -1982 9806 -1976
rect 9398 -2016 9410 -1982
rect 9794 -2016 9806 -1982
rect 9398 -2022 9806 -2016
rect 10256 -1982 10664 -1976
rect 10256 -2016 10268 -1982
rect 10652 -2016 10664 -1982
rect 10256 -2022 10664 -2016
rect 9144 -2122 9156 -2066
rect 8332 -2242 8338 -2130
rect 8292 -2254 8338 -2242
rect 9150 -2242 9156 -2122
rect 9190 -2122 9204 -2066
rect 10008 -2066 10054 -2054
rect 9190 -2242 9196 -2122
rect 10008 -2208 10014 -2066
rect 9150 -2254 9196 -2242
rect 10002 -2242 10014 -2208
rect 10048 -2208 10054 -2066
rect 10856 -2066 10916 -1910
rect 10048 -2242 10062 -2208
rect 7682 -2292 8090 -2286
rect 7682 -2326 7694 -2292
rect 8078 -2326 8090 -2292
rect 7682 -2332 8090 -2326
rect 8540 -2292 8948 -2286
rect 8540 -2326 8552 -2292
rect 8936 -2326 8948 -2292
rect 8540 -2332 8948 -2326
rect 9398 -2292 9806 -2286
rect 9398 -2326 9410 -2292
rect 9794 -2326 9806 -2292
rect 9398 -2332 9806 -2326
rect 10002 -2514 10062 -2242
rect 10856 -2242 10872 -2066
rect 10906 -2242 10916 -2066
rect 10256 -2292 10664 -2286
rect 10256 -2326 10268 -2292
rect 10652 -2326 10664 -2292
rect 10256 -2332 10664 -2326
rect 10432 -2384 10492 -2332
rect 10856 -2384 10916 -2242
rect 10432 -2444 10916 -2384
rect 9996 -2574 10002 -2514
rect 10062 -2574 10068 -2514
rect 8214 -2704 8220 -2644
rect 8280 -2704 8286 -2644
rect 8726 -2704 8732 -2644
rect 8792 -2704 8798 -2644
rect 9246 -2704 9252 -2644
rect 9312 -2704 9318 -2644
rect 9762 -2704 9768 -2644
rect 9828 -2704 9834 -2644
rect 6596 -2820 6602 -2760
rect 6662 -2762 6668 -2760
rect 6662 -2820 6792 -2762
rect 6602 -2822 6792 -2820
rect 6602 -2884 6662 -2822
rect 6576 -2890 6684 -2884
rect 6576 -2924 6588 -2890
rect 6672 -2924 6684 -2890
rect 6576 -2930 6684 -2924
rect 6472 -3004 6484 -2974
rect 6260 -3350 6274 -3306
rect 5802 -3400 5910 -3394
rect 5802 -3434 5814 -3400
rect 5898 -3434 5910 -3400
rect 5802 -3440 5910 -3434
rect 6060 -3400 6168 -3394
rect 6060 -3434 6072 -3400
rect 6156 -3434 6168 -3400
rect 6060 -3440 6168 -3434
rect 6080 -3490 6140 -3440
rect 6074 -3550 6080 -3490
rect 6140 -3550 6146 -3490
rect 5690 -3660 5696 -3600
rect 5756 -3660 5762 -3600
rect 6080 -3716 6140 -3550
rect 6214 -3716 6274 -3350
rect 6478 -3350 6484 -3004
rect 6518 -3004 6532 -2974
rect 6732 -2974 6792 -2822
rect 6856 -2818 7892 -2758
rect 8084 -2814 8090 -2754
rect 8150 -2814 8156 -2754
rect 6856 -2884 6916 -2818
rect 6834 -2890 6942 -2884
rect 6834 -2924 6846 -2890
rect 6930 -2924 6942 -2890
rect 6834 -2930 6942 -2924
rect 6518 -3350 6524 -3004
rect 6478 -3362 6524 -3350
rect 6732 -3350 6742 -2974
rect 6776 -3350 6792 -2974
rect 6318 -3400 6426 -3394
rect 6318 -3434 6330 -3400
rect 6414 -3434 6426 -3400
rect 6318 -3440 6426 -3434
rect 6576 -3400 6684 -3394
rect 6576 -3434 6588 -3400
rect 6672 -3434 6684 -3400
rect 6576 -3440 6684 -3434
rect 6342 -3490 6402 -3440
rect 6336 -3550 6342 -3490
rect 6402 -3550 6408 -3490
rect 6342 -3716 6402 -3550
rect 6732 -3600 6792 -3350
rect 6990 -2974 7050 -2818
rect 6990 -3350 7000 -2974
rect 7034 -3350 7050 -2974
rect 6834 -3400 6942 -3394
rect 6834 -3434 6846 -3400
rect 6930 -3434 6942 -3400
rect 6834 -3440 6942 -3434
rect 6858 -3490 6918 -3440
rect 6990 -3490 7050 -3350
rect 7706 -2974 7766 -2818
rect 7832 -2884 7892 -2818
rect 8090 -2884 8150 -2814
rect 7808 -2890 7916 -2884
rect 7808 -2924 7820 -2890
rect 7904 -2924 7916 -2890
rect 7808 -2930 7916 -2924
rect 8066 -2890 8174 -2884
rect 8066 -2924 8078 -2890
rect 8162 -2924 8174 -2890
rect 8066 -2930 8174 -2924
rect 7706 -3350 7716 -2974
rect 7750 -3350 7766 -2974
rect 7968 -2974 8014 -2962
rect 7968 -3300 7974 -2974
rect 7706 -3490 7766 -3350
rect 7960 -3350 7974 -3300
rect 8008 -3300 8014 -2974
rect 8220 -2974 8280 -2704
rect 8324 -2890 8432 -2884
rect 8324 -2924 8336 -2890
rect 8420 -2924 8432 -2890
rect 8324 -2930 8432 -2924
rect 8582 -2890 8690 -2884
rect 8582 -2924 8594 -2890
rect 8678 -2924 8690 -2890
rect 8582 -2930 8690 -2924
rect 8220 -2994 8232 -2974
rect 8008 -3350 8020 -3300
rect 7808 -3400 7916 -3394
rect 7808 -3434 7820 -3400
rect 7904 -3434 7916 -3400
rect 7808 -3440 7916 -3434
rect 7830 -3490 7890 -3440
rect 6858 -3550 7890 -3490
rect 6726 -3660 6732 -3600
rect 6792 -3660 6798 -3600
rect 5046 -3776 5052 -3716
rect 5112 -3776 5118 -3716
rect 5172 -3776 5178 -3716
rect 5238 -3776 5244 -3716
rect 5302 -3776 5308 -3716
rect 5368 -3776 5374 -3716
rect 6074 -3776 6080 -3716
rect 6140 -3776 6146 -3716
rect 6208 -3776 6214 -3716
rect 6274 -3776 6280 -3716
rect 6336 -3776 6342 -3716
rect 6402 -3776 6408 -3716
rect 6858 -3816 6918 -3550
rect 6990 -3816 7050 -3550
rect 7706 -3816 7766 -3550
rect 7830 -3816 7890 -3550
rect 7960 -3594 8020 -3350
rect 8226 -3350 8232 -2994
rect 8266 -2994 8280 -2974
rect 8484 -2974 8530 -2962
rect 8266 -3350 8272 -2994
rect 8484 -3304 8490 -2974
rect 8226 -3362 8272 -3350
rect 8474 -3350 8490 -3304
rect 8524 -3304 8530 -2974
rect 8732 -2974 8792 -2704
rect 8860 -2814 8866 -2754
rect 8926 -2814 8932 -2754
rect 9114 -2814 9120 -2754
rect 9180 -2814 9186 -2754
rect 8866 -2884 8926 -2814
rect 9120 -2884 9180 -2814
rect 8840 -2890 8948 -2884
rect 8840 -2924 8852 -2890
rect 8936 -2924 8948 -2890
rect 8840 -2930 8948 -2924
rect 9098 -2890 9206 -2884
rect 9098 -2924 9110 -2890
rect 9194 -2924 9206 -2890
rect 9098 -2930 9206 -2924
rect 8732 -2994 8748 -2974
rect 8524 -3350 8534 -3304
rect 8066 -3400 8174 -3394
rect 8066 -3434 8078 -3400
rect 8162 -3434 8174 -3400
rect 8066 -3440 8174 -3434
rect 8324 -3400 8432 -3394
rect 8324 -3434 8336 -3400
rect 8420 -3434 8432 -3400
rect 8324 -3440 8432 -3434
rect 8350 -3484 8410 -3440
rect 8344 -3544 8350 -3484
rect 8410 -3544 8416 -3484
rect 7954 -3654 7960 -3594
rect 8020 -3654 8026 -3594
rect 8474 -3710 8534 -3350
rect 8742 -3350 8748 -2994
rect 8782 -2994 8792 -2974
rect 9000 -2974 9046 -2962
rect 8782 -3350 8788 -2994
rect 9000 -3290 9006 -2974
rect 8742 -3362 8788 -3350
rect 8992 -3350 9006 -3290
rect 9040 -3290 9046 -2974
rect 9252 -2974 9312 -2704
rect 9356 -2890 9464 -2884
rect 9356 -2924 9368 -2890
rect 9452 -2924 9464 -2890
rect 9356 -2930 9464 -2924
rect 9614 -2890 9722 -2884
rect 9614 -2924 9626 -2890
rect 9710 -2924 9722 -2890
rect 9614 -2930 9722 -2924
rect 9252 -2998 9264 -2974
rect 9040 -3350 9052 -3290
rect 8582 -3400 8690 -3394
rect 8582 -3434 8594 -3400
rect 8678 -3434 8690 -3400
rect 8582 -3440 8690 -3434
rect 8840 -3400 8948 -3394
rect 8840 -3434 8852 -3400
rect 8936 -3434 8948 -3400
rect 8840 -3440 8948 -3434
rect 8604 -3484 8664 -3440
rect 8598 -3544 8604 -3484
rect 8664 -3544 8670 -3484
rect 8992 -3594 9052 -3350
rect 9258 -3350 9264 -2998
rect 9298 -2998 9312 -2974
rect 9516 -2974 9562 -2962
rect 9298 -3350 9304 -2998
rect 9516 -3300 9522 -2974
rect 9258 -3362 9304 -3350
rect 9510 -3350 9522 -3300
rect 9556 -3300 9562 -2974
rect 9768 -2974 9828 -2704
rect 10432 -2752 10492 -2444
rect 10856 -2752 10916 -2444
rect 10988 -2644 11048 -1376
rect 10982 -2704 10988 -2644
rect 11048 -2704 11054 -2644
rect 11304 -2752 11310 -778
rect 9892 -2814 9898 -2754
rect 9958 -2814 9964 -2754
rect 10152 -2812 11310 -2752
rect 9898 -2884 9958 -2814
rect 10152 -2884 10212 -2812
rect 9872 -2890 9980 -2884
rect 9872 -2924 9884 -2890
rect 9968 -2924 9980 -2890
rect 9872 -2930 9980 -2924
rect 10130 -2890 10238 -2884
rect 10130 -2924 10142 -2890
rect 10226 -2924 10238 -2890
rect 10130 -2930 10238 -2924
rect 9768 -2998 9780 -2974
rect 9556 -3350 9570 -3300
rect 9376 -3394 9436 -3390
rect 9098 -3400 9206 -3394
rect 9098 -3434 9110 -3400
rect 9194 -3434 9206 -3400
rect 9098 -3440 9206 -3434
rect 9356 -3400 9464 -3394
rect 9356 -3434 9368 -3400
rect 9452 -3434 9464 -3400
rect 9356 -3440 9464 -3434
rect 9376 -3484 9436 -3440
rect 9370 -3544 9376 -3484
rect 9436 -3544 9442 -3484
rect 8986 -3654 8992 -3594
rect 9052 -3654 9058 -3594
rect 9510 -3710 9570 -3350
rect 9774 -3350 9780 -2998
rect 9814 -2998 9828 -2974
rect 10032 -2974 10078 -2962
rect 9814 -3350 9820 -2998
rect 10032 -3294 10038 -2974
rect 9774 -3362 9820 -3350
rect 10028 -3350 10038 -3294
rect 10072 -3294 10078 -2974
rect 10286 -2974 10346 -2812
rect 10072 -3350 10088 -3294
rect 9614 -3400 9722 -3394
rect 9614 -3434 9626 -3400
rect 9710 -3434 9722 -3400
rect 9614 -3440 9722 -3434
rect 9872 -3400 9980 -3394
rect 9872 -3434 9884 -3400
rect 9968 -3434 9980 -3400
rect 9872 -3440 9980 -3434
rect 9638 -3484 9698 -3440
rect 9632 -3544 9638 -3484
rect 9698 -3544 9704 -3484
rect 10028 -3594 10088 -3350
rect 10286 -3350 10296 -2974
rect 10330 -3350 10346 -2974
rect 10130 -3400 10238 -3394
rect 10130 -3434 10142 -3400
rect 10226 -3434 10238 -3400
rect 10130 -3440 10238 -3434
rect 10154 -3482 10214 -3440
rect 10286 -3482 10346 -3350
rect 11304 -3482 11310 -2812
rect 10154 -3542 11310 -3482
rect 10022 -3654 10028 -3594
rect 10088 -3654 10094 -3594
rect 8468 -3770 8474 -3710
rect 8534 -3770 8540 -3710
rect 9504 -3770 9510 -3710
rect 9570 -3770 9576 -3710
rect 10154 -3816 10214 -3542
rect 10286 -3816 10346 -3542
rect 11304 -3662 11310 -3542
rect 11410 -3662 11416 -778
rect 11304 -3816 11416 -3662
rect 60 -3822 11416 -3816
rect 60 -3922 166 -3822
rect 11310 -3922 11416 -3822
rect 60 -3928 11416 -3922
rect 11860 -518 23216 -512
rect 11860 -618 11966 -518
rect 23110 -618 23216 -518
rect 11860 -624 23216 -618
rect 11860 -778 11972 -624
rect 11860 -3662 11866 -778
rect 11966 -2752 11972 -778
rect 12572 -924 12582 -624
rect 22494 -924 22504 -624
rect 23104 -778 23216 -624
rect 12122 -1046 22896 -990
rect 12122 -1156 12184 -1046
rect 22840 -1156 22896 -1046
rect 12122 -1204 22896 -1156
rect 12214 -1370 12220 -1310
rect 12280 -1370 12286 -1310
rect 12360 -1318 12420 -1204
rect 12780 -1318 12840 -1204
rect 12220 -2644 12280 -1370
rect 12360 -1378 12840 -1318
rect 12360 -1526 12420 -1378
rect 12780 -1436 12840 -1378
rect 12618 -1442 13026 -1436
rect 12618 -1476 12630 -1442
rect 13014 -1476 13026 -1442
rect 12618 -1482 13026 -1476
rect 13476 -1442 13884 -1436
rect 13476 -1476 13488 -1442
rect 13872 -1476 13884 -1442
rect 13476 -1482 13884 -1476
rect 12360 -1702 12376 -1526
rect 12410 -1702 12420 -1526
rect 13228 -1526 13274 -1514
rect 13228 -1650 13234 -1526
rect 12360 -1848 12420 -1702
rect 13220 -1702 13234 -1650
rect 13268 -1650 13274 -1526
rect 14078 -1526 14138 -1204
rect 14334 -1442 14742 -1436
rect 14334 -1476 14346 -1442
rect 14730 -1476 14742 -1442
rect 14334 -1482 14742 -1476
rect 15192 -1442 15600 -1436
rect 15192 -1476 15204 -1442
rect 15588 -1476 15600 -1442
rect 15192 -1482 15600 -1476
rect 13268 -1702 13280 -1650
rect 12618 -1752 13026 -1746
rect 12618 -1786 12630 -1752
rect 13014 -1786 13026 -1752
rect 12618 -1792 13026 -1786
rect 12784 -1848 12844 -1792
rect 12360 -1908 12844 -1848
rect 13220 -1854 13280 -1702
rect 14078 -1702 14092 -1526
rect 14126 -1702 14138 -1526
rect 14944 -1526 14990 -1514
rect 14944 -1674 14950 -1526
rect 13476 -1752 13884 -1746
rect 13476 -1786 13488 -1752
rect 13872 -1786 13884 -1752
rect 13476 -1792 13884 -1786
rect 13644 -1854 13704 -1792
rect 12360 -2066 12420 -1908
rect 12784 -1976 12844 -1908
rect 13214 -1914 13220 -1854
rect 13280 -1914 13704 -1854
rect 13644 -1976 13704 -1914
rect 12618 -1982 13026 -1976
rect 12618 -2016 12630 -1982
rect 13014 -2016 13026 -1982
rect 12618 -2022 13026 -2016
rect 13476 -1982 13884 -1976
rect 13476 -2016 13488 -1982
rect 13872 -2016 13884 -1982
rect 13476 -2022 13884 -2016
rect 12360 -2242 12376 -2066
rect 12410 -2242 12420 -2066
rect 13228 -2066 13274 -2054
rect 13228 -2204 13234 -2066
rect 12360 -2398 12420 -2242
rect 13218 -2242 13234 -2204
rect 13268 -2204 13274 -2066
rect 14078 -2066 14138 -1702
rect 14936 -1702 14950 -1674
rect 14984 -1674 14990 -1526
rect 15794 -1526 15854 -1204
rect 17082 -1312 17142 -1204
rect 17508 -1312 17568 -1204
rect 17944 -1312 18004 -1204
rect 17082 -1372 18004 -1312
rect 18362 -1370 18368 -1310
rect 18428 -1370 18434 -1310
rect 17082 -1436 17142 -1372
rect 16050 -1442 16458 -1436
rect 16050 -1476 16062 -1442
rect 16446 -1476 16458 -1442
rect 16050 -1482 16458 -1476
rect 16908 -1442 17316 -1436
rect 16908 -1476 16920 -1442
rect 17304 -1476 17316 -1442
rect 16908 -1482 17316 -1476
rect 14984 -1702 14996 -1674
rect 14334 -1752 14742 -1746
rect 14334 -1786 14346 -1752
rect 14730 -1786 14742 -1752
rect 14334 -1792 14742 -1786
rect 14502 -1854 14562 -1792
rect 14936 -1854 14996 -1702
rect 15794 -1702 15808 -1526
rect 15842 -1702 15854 -1526
rect 16660 -1526 16706 -1514
rect 16660 -1650 16666 -1526
rect 15192 -1752 15600 -1746
rect 15192 -1786 15204 -1752
rect 15588 -1786 15600 -1752
rect 15192 -1792 15600 -1786
rect 14496 -1858 14568 -1854
rect 14496 -1914 14502 -1858
rect 14562 -1914 14568 -1858
rect 14930 -1914 14936 -1854
rect 14996 -1914 15002 -1854
rect 15366 -1858 15426 -1792
rect 14502 -1976 14562 -1914
rect 14334 -1982 14742 -1976
rect 14334 -2016 14346 -1982
rect 14730 -2016 14742 -1982
rect 14334 -2022 14742 -2016
rect 14078 -2146 14092 -2066
rect 13268 -2242 13278 -2204
rect 12618 -2292 13026 -2286
rect 12618 -2326 12630 -2292
rect 13014 -2326 13026 -2292
rect 12618 -2332 13026 -2326
rect 12782 -2398 12842 -2332
rect 13218 -2398 13278 -2242
rect 14086 -2242 14092 -2146
rect 14126 -2146 14138 -2066
rect 14936 -2066 14996 -1914
rect 15366 -1976 15426 -1914
rect 15192 -1982 15600 -1976
rect 15192 -2016 15204 -1982
rect 15588 -2016 15600 -1982
rect 15192 -2022 15600 -2016
rect 14936 -2116 14950 -2066
rect 14126 -2242 14132 -2146
rect 14086 -2254 14132 -2242
rect 14944 -2242 14950 -2116
rect 14984 -2116 14996 -2066
rect 15794 -2066 15854 -1702
rect 16656 -1702 16666 -1650
rect 16700 -1650 16706 -1526
rect 17508 -1526 17568 -1372
rect 17944 -1436 18004 -1372
rect 17766 -1442 18174 -1436
rect 17766 -1476 17778 -1442
rect 18162 -1476 18174 -1442
rect 17766 -1482 18174 -1476
rect 16700 -1702 16716 -1650
rect 16050 -1752 16458 -1746
rect 16050 -1786 16062 -1752
rect 16446 -1786 16458 -1752
rect 16050 -1792 16458 -1786
rect 16226 -1858 16286 -1792
rect 16656 -1854 16716 -1702
rect 17508 -1702 17524 -1526
rect 17558 -1702 17568 -1526
rect 18368 -1526 18428 -1370
rect 18624 -1442 19032 -1436
rect 18624 -1476 18636 -1442
rect 19020 -1476 19032 -1442
rect 18624 -1482 19032 -1476
rect 18368 -1556 18382 -1526
rect 16908 -1752 17316 -1746
rect 16908 -1786 16920 -1752
rect 17304 -1786 17316 -1752
rect 16908 -1792 17316 -1786
rect 16650 -1914 16656 -1854
rect 16716 -1914 16722 -1854
rect 17084 -1856 17144 -1792
rect 17508 -1856 17568 -1702
rect 18376 -1702 18382 -1556
rect 18416 -1556 18428 -1526
rect 19226 -1526 19286 -1204
rect 19482 -1442 19890 -1436
rect 19482 -1476 19494 -1442
rect 19878 -1476 19890 -1442
rect 19482 -1482 19890 -1476
rect 20340 -1442 20748 -1436
rect 20340 -1476 20352 -1442
rect 20736 -1476 20748 -1442
rect 20340 -1482 20748 -1476
rect 18416 -1702 18422 -1556
rect 18376 -1714 18422 -1702
rect 19226 -1702 19240 -1526
rect 19274 -1702 19286 -1526
rect 20092 -1526 20138 -1514
rect 20092 -1660 20098 -1526
rect 17766 -1752 18174 -1746
rect 17766 -1786 17778 -1752
rect 18162 -1786 18174 -1752
rect 17766 -1792 18174 -1786
rect 18624 -1752 19032 -1746
rect 18624 -1786 18636 -1752
rect 19020 -1786 19032 -1752
rect 18624 -1792 19032 -1786
rect 17944 -1856 18004 -1792
rect 18798 -1854 18858 -1792
rect 16226 -1976 16286 -1914
rect 17084 -1916 18004 -1856
rect 18366 -1914 18372 -1854
rect 18432 -1914 18438 -1854
rect 18792 -1858 18864 -1854
rect 18792 -1914 18798 -1858
rect 18858 -1914 18864 -1858
rect 17084 -1976 17144 -1916
rect 16050 -1982 16458 -1976
rect 16050 -2016 16062 -1982
rect 16446 -2016 16458 -1982
rect 16050 -2022 16458 -2016
rect 16908 -1982 17316 -1976
rect 16908 -2016 16920 -1982
rect 17304 -2016 17316 -1982
rect 16908 -2022 17316 -2016
rect 14984 -2242 14990 -2116
rect 14944 -2254 14990 -2242
rect 15794 -2242 15808 -2066
rect 15842 -2242 15854 -2066
rect 16660 -2066 16706 -2054
rect 16660 -2200 16666 -2066
rect 13476 -2292 13884 -2286
rect 13476 -2326 13488 -2292
rect 13872 -2326 13884 -2292
rect 13476 -2332 13884 -2326
rect 14334 -2292 14742 -2286
rect 14334 -2326 14346 -2292
rect 14730 -2326 14742 -2292
rect 14334 -2332 14742 -2326
rect 15192 -2292 15600 -2286
rect 15192 -2326 15204 -2292
rect 15588 -2326 15600 -2292
rect 15192 -2332 15600 -2326
rect 12360 -2458 12842 -2398
rect 13212 -2458 13218 -2398
rect 13278 -2458 13284 -2398
rect 12214 -2704 12220 -2644
rect 12280 -2704 12286 -2644
rect 12360 -2752 12420 -2458
rect 15100 -2582 15106 -2522
rect 15166 -2582 15172 -2522
rect 13428 -2644 13488 -2638
rect 13934 -2704 13940 -2644
rect 14000 -2704 14006 -2644
rect 14454 -2704 14460 -2644
rect 14520 -2704 14526 -2644
rect 14970 -2704 14976 -2644
rect 15036 -2704 15042 -2644
rect 11966 -2812 13100 -2752
rect 11966 -3484 11972 -2812
rect 12914 -2974 12974 -2812
rect 13040 -2884 13100 -2812
rect 13292 -2814 13298 -2754
rect 13358 -2814 13364 -2754
rect 13298 -2884 13358 -2814
rect 13016 -2890 13124 -2884
rect 13016 -2924 13028 -2890
rect 13112 -2924 13124 -2890
rect 13016 -2930 13124 -2924
rect 13274 -2890 13382 -2884
rect 13274 -2924 13286 -2890
rect 13370 -2924 13382 -2890
rect 13274 -2930 13382 -2924
rect 12914 -3350 12924 -2974
rect 12958 -3350 12974 -2974
rect 13176 -2974 13222 -2962
rect 13176 -3300 13182 -2974
rect 12914 -3484 12974 -3350
rect 13168 -3350 13182 -3300
rect 13216 -3300 13222 -2974
rect 13428 -2974 13488 -2704
rect 13532 -2890 13640 -2884
rect 13532 -2924 13544 -2890
rect 13628 -2924 13640 -2890
rect 13532 -2930 13640 -2924
rect 13790 -2890 13898 -2884
rect 13790 -2924 13802 -2890
rect 13886 -2924 13898 -2890
rect 13790 -2930 13898 -2924
rect 13428 -2994 13440 -2974
rect 13216 -3350 13228 -3300
rect 13016 -3400 13124 -3394
rect 13016 -3434 13028 -3400
rect 13112 -3434 13124 -3400
rect 13016 -3440 13124 -3434
rect 13040 -3484 13100 -3440
rect 11966 -3544 13100 -3484
rect 11966 -3662 11972 -3544
rect 11860 -3816 11972 -3662
rect 12914 -3816 12974 -3544
rect 13040 -3816 13100 -3544
rect 13168 -3594 13228 -3350
rect 13434 -3350 13440 -2994
rect 13474 -2994 13488 -2974
rect 13692 -2974 13738 -2962
rect 13474 -3350 13480 -2994
rect 13692 -3304 13698 -2974
rect 13434 -3362 13480 -3350
rect 13682 -3350 13698 -3304
rect 13732 -3304 13738 -2974
rect 13940 -2974 14000 -2704
rect 14068 -2814 14074 -2754
rect 14134 -2814 14140 -2754
rect 14322 -2814 14328 -2754
rect 14388 -2814 14394 -2754
rect 14074 -2884 14134 -2814
rect 14328 -2884 14388 -2814
rect 14048 -2890 14156 -2884
rect 14048 -2924 14060 -2890
rect 14144 -2924 14156 -2890
rect 14048 -2930 14156 -2924
rect 14306 -2890 14414 -2884
rect 14306 -2924 14318 -2890
rect 14402 -2924 14414 -2890
rect 14306 -2930 14414 -2924
rect 13940 -2994 13956 -2974
rect 13732 -3350 13742 -3304
rect 13274 -3400 13382 -3394
rect 13274 -3434 13286 -3400
rect 13370 -3434 13382 -3400
rect 13274 -3440 13382 -3434
rect 13532 -3400 13640 -3394
rect 13532 -3434 13544 -3400
rect 13628 -3434 13640 -3400
rect 13532 -3440 13640 -3434
rect 13558 -3484 13618 -3440
rect 13552 -3544 13558 -3484
rect 13618 -3544 13624 -3484
rect 13162 -3654 13168 -3594
rect 13228 -3654 13234 -3594
rect 13682 -3710 13742 -3350
rect 13950 -3350 13956 -2994
rect 13990 -2994 14000 -2974
rect 14208 -2974 14254 -2962
rect 13990 -3350 13996 -2994
rect 14208 -3290 14214 -2974
rect 13950 -3362 13996 -3350
rect 14200 -3350 14214 -3290
rect 14248 -3290 14254 -2974
rect 14460 -2974 14520 -2704
rect 14564 -2890 14672 -2884
rect 14564 -2924 14576 -2890
rect 14660 -2924 14672 -2890
rect 14564 -2930 14672 -2924
rect 14822 -2890 14930 -2884
rect 14822 -2924 14834 -2890
rect 14918 -2924 14930 -2890
rect 14822 -2930 14930 -2924
rect 14460 -2998 14472 -2974
rect 14248 -3350 14260 -3290
rect 13790 -3400 13898 -3394
rect 13790 -3434 13802 -3400
rect 13886 -3434 13898 -3400
rect 13790 -3440 13898 -3434
rect 14048 -3400 14156 -3394
rect 14048 -3434 14060 -3400
rect 14144 -3434 14156 -3400
rect 14048 -3440 14156 -3434
rect 13812 -3484 13872 -3440
rect 13806 -3544 13812 -3484
rect 13872 -3544 13878 -3484
rect 14200 -3594 14260 -3350
rect 14466 -3350 14472 -2998
rect 14506 -2998 14520 -2974
rect 14724 -2974 14770 -2962
rect 14506 -3350 14512 -2998
rect 14724 -3300 14730 -2974
rect 14466 -3362 14512 -3350
rect 14718 -3350 14730 -3300
rect 14764 -3300 14770 -2974
rect 14976 -2974 15036 -2704
rect 15106 -2754 15166 -2582
rect 15794 -2752 15854 -2242
rect 16652 -2242 16666 -2200
rect 16700 -2200 16706 -2066
rect 17508 -2066 17568 -1916
rect 17944 -1976 18004 -1916
rect 17766 -1982 18174 -1976
rect 17766 -2016 17778 -1982
rect 18162 -2016 18174 -1982
rect 17766 -2022 18174 -2016
rect 16700 -2242 16712 -2200
rect 16050 -2292 16458 -2286
rect 16050 -2326 16062 -2292
rect 16446 -2326 16458 -2292
rect 16050 -2332 16458 -2326
rect 16652 -2398 16712 -2242
rect 17508 -2242 17524 -2066
rect 17558 -2242 17568 -2066
rect 18372 -2066 18432 -1914
rect 18798 -1976 18858 -1914
rect 18624 -1982 19032 -1976
rect 18624 -2016 18636 -1982
rect 19020 -2016 19032 -1982
rect 18624 -2022 19032 -2016
rect 18372 -2114 18382 -2066
rect 16908 -2292 17316 -2286
rect 16908 -2326 16920 -2292
rect 17304 -2326 17316 -2292
rect 16908 -2332 17316 -2326
rect 16646 -2458 16652 -2398
rect 16712 -2458 16784 -2398
rect 16724 -2650 16784 -2458
rect 17082 -2400 17142 -2332
rect 17508 -2400 17568 -2242
rect 18376 -2242 18382 -2114
rect 18416 -2114 18432 -2066
rect 19226 -2066 19286 -1702
rect 20084 -1702 20098 -1660
rect 20132 -1660 20138 -1526
rect 20944 -1526 21004 -1204
rect 22232 -1316 22292 -1204
rect 22656 -1316 22716 -1204
rect 21794 -1376 21800 -1316
rect 21860 -1376 21866 -1316
rect 22232 -1376 22716 -1316
rect 22782 -1376 22788 -1316
rect 22848 -1376 22854 -1316
rect 21198 -1442 21606 -1436
rect 21198 -1476 21210 -1442
rect 21594 -1476 21606 -1442
rect 21198 -1482 21606 -1476
rect 20132 -1702 20144 -1660
rect 19482 -1752 19890 -1746
rect 19482 -1786 19494 -1752
rect 19878 -1786 19890 -1752
rect 19482 -1792 19890 -1786
rect 19656 -1858 19716 -1792
rect 20084 -1854 20144 -1702
rect 20944 -1702 20956 -1526
rect 20990 -1702 21004 -1526
rect 21800 -1526 21860 -1376
rect 22232 -1436 22292 -1376
rect 22056 -1442 22464 -1436
rect 22056 -1476 22068 -1442
rect 22452 -1476 22464 -1442
rect 22056 -1482 22464 -1476
rect 21800 -1558 21814 -1526
rect 20340 -1752 20748 -1746
rect 20340 -1786 20352 -1752
rect 20736 -1786 20748 -1752
rect 20340 -1792 20748 -1786
rect 20078 -1914 20084 -1854
rect 20144 -1914 20150 -1854
rect 20510 -1858 20570 -1792
rect 19656 -1976 19716 -1914
rect 19482 -1982 19890 -1976
rect 19482 -2016 19494 -1982
rect 19878 -2016 19890 -1982
rect 19482 -2022 19890 -2016
rect 18416 -2242 18422 -2114
rect 18376 -2254 18422 -2242
rect 19226 -2242 19240 -2066
rect 19274 -2242 19286 -2066
rect 20084 -2066 20144 -1914
rect 20510 -1976 20570 -1914
rect 20340 -1982 20748 -1976
rect 20340 -2016 20352 -1982
rect 20736 -2016 20748 -1982
rect 20340 -2022 20748 -2016
rect 20084 -2130 20098 -2066
rect 17766 -2292 18174 -2286
rect 17766 -2326 17778 -2292
rect 18162 -2326 18174 -2292
rect 17766 -2332 18174 -2326
rect 18624 -2292 19032 -2286
rect 18624 -2326 18636 -2292
rect 19020 -2326 19032 -2292
rect 18624 -2332 19032 -2326
rect 17946 -2400 18006 -2332
rect 17082 -2460 18006 -2400
rect 16980 -2582 16986 -2522
rect 17046 -2582 17052 -2522
rect 15100 -2814 15106 -2754
rect 15166 -2814 15172 -2754
rect 15360 -2812 16396 -2752
rect 15106 -2884 15166 -2814
rect 15360 -2884 15420 -2812
rect 15080 -2890 15188 -2884
rect 15080 -2924 15092 -2890
rect 15176 -2924 15188 -2890
rect 15080 -2930 15188 -2924
rect 15338 -2890 15446 -2884
rect 15338 -2924 15350 -2890
rect 15434 -2924 15446 -2890
rect 15338 -2930 15446 -2924
rect 14976 -2998 14988 -2974
rect 14764 -3350 14778 -3300
rect 14584 -3394 14644 -3390
rect 14306 -3400 14414 -3394
rect 14306 -3434 14318 -3400
rect 14402 -3434 14414 -3400
rect 14306 -3440 14414 -3434
rect 14564 -3400 14672 -3394
rect 14564 -3434 14576 -3400
rect 14660 -3434 14672 -3400
rect 14564 -3440 14672 -3434
rect 14584 -3484 14644 -3440
rect 14578 -3544 14584 -3484
rect 14644 -3544 14650 -3484
rect 14194 -3654 14200 -3594
rect 14260 -3654 14266 -3594
rect 14718 -3710 14778 -3350
rect 14982 -3350 14988 -2998
rect 15022 -2998 15036 -2974
rect 15240 -2974 15286 -2962
rect 15022 -3350 15028 -2998
rect 15240 -3294 15246 -2974
rect 14982 -3362 15028 -3350
rect 15236 -3350 15246 -3294
rect 15280 -3294 15286 -2974
rect 15494 -2974 15554 -2812
rect 15280 -3350 15296 -3294
rect 14822 -3400 14930 -3394
rect 14822 -3434 14834 -3400
rect 14918 -3434 14930 -3400
rect 14822 -3440 14930 -3434
rect 15080 -3400 15188 -3394
rect 15080 -3434 15092 -3400
rect 15176 -3434 15188 -3400
rect 15080 -3440 15188 -3434
rect 14846 -3484 14906 -3440
rect 14840 -3544 14846 -3484
rect 14906 -3544 14912 -3484
rect 15236 -3594 15296 -3350
rect 15494 -3350 15504 -2974
rect 15538 -3350 15554 -2974
rect 15338 -3400 15446 -3394
rect 15338 -3434 15350 -3400
rect 15434 -3434 15446 -3400
rect 15338 -3440 15446 -3434
rect 15360 -3484 15420 -3440
rect 15494 -3484 15554 -3350
rect 16210 -2974 16270 -2812
rect 16336 -2884 16396 -2812
rect 16588 -2820 16594 -2760
rect 16654 -2820 16660 -2760
rect 16594 -2884 16654 -2820
rect 16312 -2890 16420 -2884
rect 16312 -2924 16324 -2890
rect 16408 -2924 16420 -2890
rect 16312 -2930 16420 -2924
rect 16570 -2890 16678 -2884
rect 16570 -2924 16582 -2890
rect 16666 -2924 16678 -2890
rect 16570 -2930 16678 -2924
rect 16210 -3350 16220 -2974
rect 16254 -3350 16270 -2974
rect 16472 -2974 16518 -2962
rect 16472 -3306 16478 -2974
rect 16210 -3484 16270 -3350
rect 16464 -3350 16478 -3306
rect 16512 -3306 16518 -2974
rect 16724 -2974 16784 -2710
rect 16828 -2890 16936 -2884
rect 16828 -2924 16840 -2890
rect 16924 -2924 16936 -2890
rect 16828 -2930 16936 -2924
rect 16724 -3000 16736 -2974
rect 16512 -3350 16524 -3306
rect 16312 -3400 16420 -3394
rect 16312 -3434 16324 -3400
rect 16408 -3434 16420 -3400
rect 16312 -3440 16420 -3434
rect 16334 -3484 16394 -3440
rect 15360 -3544 16394 -3484
rect 15230 -3654 15236 -3594
rect 15296 -3654 15302 -3594
rect 13676 -3770 13682 -3710
rect 13742 -3770 13748 -3710
rect 14712 -3770 14718 -3710
rect 14778 -3770 14784 -3710
rect 15360 -3816 15420 -3544
rect 15494 -3816 15554 -3544
rect 16210 -3816 16270 -3544
rect 16334 -3816 16394 -3544
rect 16464 -3600 16524 -3350
rect 16730 -3350 16736 -3000
rect 16770 -3000 16784 -2974
rect 16986 -2974 17046 -2582
rect 17230 -2710 17236 -2650
rect 17296 -2710 17302 -2650
rect 17750 -2710 17756 -2650
rect 17816 -2710 17822 -2650
rect 18266 -2710 18272 -2650
rect 18332 -2710 18338 -2650
rect 17086 -2890 17194 -2884
rect 17086 -2924 17098 -2890
rect 17182 -2924 17194 -2890
rect 17086 -2930 17194 -2924
rect 16770 -3350 16776 -3000
rect 16986 -3062 16994 -2974
rect 16988 -3310 16994 -3062
rect 16730 -3362 16776 -3350
rect 16978 -3350 16994 -3310
rect 17028 -3062 17046 -2974
rect 17236 -2974 17296 -2710
rect 17364 -2820 17370 -2760
rect 17430 -2820 17436 -2760
rect 17618 -2820 17624 -2760
rect 17684 -2820 17690 -2760
rect 17370 -2884 17430 -2820
rect 17624 -2884 17684 -2820
rect 17344 -2890 17452 -2884
rect 17344 -2924 17356 -2890
rect 17440 -2924 17452 -2890
rect 17344 -2930 17452 -2924
rect 17602 -2890 17710 -2884
rect 17602 -2924 17614 -2890
rect 17698 -2924 17710 -2890
rect 17602 -2930 17710 -2924
rect 17236 -3000 17252 -2974
rect 17028 -3310 17034 -3062
rect 17028 -3350 17038 -3310
rect 16570 -3400 16678 -3394
rect 16570 -3434 16582 -3400
rect 16666 -3434 16678 -3400
rect 16570 -3440 16678 -3434
rect 16828 -3400 16936 -3394
rect 16828 -3434 16840 -3400
rect 16924 -3434 16936 -3400
rect 16828 -3440 16936 -3434
rect 16854 -3490 16914 -3440
rect 16848 -3550 16854 -3490
rect 16914 -3550 16920 -3490
rect 16458 -3660 16464 -3600
rect 16524 -3660 16530 -3600
rect 16854 -3712 16914 -3550
rect 16848 -3772 16854 -3712
rect 16914 -3772 16920 -3712
rect 16978 -3716 17038 -3350
rect 17246 -3350 17252 -3000
rect 17286 -3000 17296 -2974
rect 17504 -2974 17550 -2962
rect 17286 -3350 17292 -3000
rect 17504 -3296 17510 -2974
rect 17246 -3362 17292 -3350
rect 17496 -3350 17510 -3296
rect 17544 -3296 17550 -2974
rect 17756 -2974 17816 -2710
rect 17860 -2890 17968 -2884
rect 17860 -2924 17872 -2890
rect 17956 -2924 17968 -2890
rect 17860 -2930 17968 -2924
rect 18118 -2890 18226 -2884
rect 18118 -2924 18130 -2890
rect 18214 -2924 18226 -2890
rect 18118 -2930 18226 -2924
rect 17756 -3004 17768 -2974
rect 17544 -3350 17556 -3296
rect 17086 -3400 17194 -3394
rect 17086 -3434 17098 -3400
rect 17182 -3434 17194 -3400
rect 17086 -3440 17194 -3434
rect 17344 -3400 17452 -3394
rect 17344 -3434 17356 -3400
rect 17440 -3434 17452 -3400
rect 17344 -3440 17452 -3434
rect 17108 -3490 17168 -3440
rect 17102 -3550 17108 -3490
rect 17168 -3550 17174 -3490
rect 17496 -3600 17556 -3350
rect 17762 -3350 17768 -3004
rect 17802 -3004 17816 -2974
rect 18020 -2974 18066 -2962
rect 17802 -3350 17808 -3004
rect 18020 -3306 18026 -2974
rect 17762 -3362 17808 -3350
rect 18014 -3350 18026 -3306
rect 18060 -3306 18066 -2974
rect 18272 -2974 18332 -2710
rect 19226 -2758 19286 -2242
rect 20092 -2242 20098 -2130
rect 20132 -2130 20144 -2066
rect 20944 -2066 21004 -1702
rect 21808 -1702 21814 -1558
rect 21848 -1558 21860 -1526
rect 22656 -1526 22716 -1376
rect 21848 -1702 21854 -1558
rect 21808 -1714 21854 -1702
rect 22656 -1702 22672 -1526
rect 22706 -1702 22716 -1526
rect 21198 -1752 21606 -1746
rect 21198 -1786 21210 -1752
rect 21594 -1786 21606 -1752
rect 21198 -1792 21606 -1786
rect 22056 -1752 22464 -1746
rect 22056 -1786 22068 -1752
rect 22452 -1786 22464 -1752
rect 22056 -1792 22464 -1786
rect 21374 -1848 21434 -1792
rect 21374 -1854 21436 -1848
rect 21374 -1914 21376 -1854
rect 21374 -1920 21436 -1914
rect 22230 -1850 22290 -1792
rect 22656 -1850 22716 -1702
rect 22230 -1910 22716 -1850
rect 21374 -1976 21434 -1920
rect 22230 -1976 22290 -1910
rect 21198 -1982 21606 -1976
rect 21198 -2016 21210 -1982
rect 21594 -2016 21606 -1982
rect 21198 -2022 21606 -2016
rect 22056 -1982 22464 -1976
rect 22056 -2016 22068 -1982
rect 22452 -2016 22464 -1982
rect 22056 -2022 22464 -2016
rect 20944 -2122 20956 -2066
rect 20132 -2242 20138 -2130
rect 20092 -2254 20138 -2242
rect 20950 -2242 20956 -2122
rect 20990 -2122 21004 -2066
rect 21808 -2066 21854 -2054
rect 20990 -2242 20996 -2122
rect 21808 -2208 21814 -2066
rect 20950 -2254 20996 -2242
rect 21802 -2242 21814 -2208
rect 21848 -2208 21854 -2066
rect 22656 -2066 22716 -1910
rect 21848 -2242 21862 -2208
rect 19482 -2292 19890 -2286
rect 19482 -2326 19494 -2292
rect 19878 -2326 19890 -2292
rect 19482 -2332 19890 -2326
rect 20340 -2292 20748 -2286
rect 20340 -2326 20352 -2292
rect 20736 -2326 20748 -2292
rect 20340 -2332 20748 -2326
rect 21198 -2292 21606 -2286
rect 21198 -2326 21210 -2292
rect 21594 -2326 21606 -2292
rect 21198 -2332 21606 -2326
rect 21802 -2514 21862 -2242
rect 22656 -2242 22672 -2066
rect 22706 -2242 22716 -2066
rect 22056 -2292 22464 -2286
rect 22056 -2326 22068 -2292
rect 22452 -2326 22464 -2292
rect 22056 -2332 22464 -2326
rect 22232 -2384 22292 -2332
rect 22656 -2384 22716 -2242
rect 22232 -2444 22716 -2384
rect 21796 -2574 21802 -2514
rect 21862 -2574 21868 -2514
rect 20014 -2704 20020 -2644
rect 20080 -2704 20086 -2644
rect 20526 -2704 20532 -2644
rect 20592 -2704 20598 -2644
rect 21046 -2704 21052 -2644
rect 21112 -2704 21118 -2644
rect 21562 -2704 21568 -2644
rect 21628 -2704 21634 -2644
rect 18396 -2820 18402 -2760
rect 18462 -2820 18468 -2760
rect 18656 -2818 19692 -2758
rect 19884 -2814 19890 -2754
rect 19950 -2814 19956 -2754
rect 18402 -2884 18462 -2820
rect 18656 -2884 18716 -2818
rect 18376 -2890 18484 -2884
rect 18376 -2924 18388 -2890
rect 18472 -2924 18484 -2890
rect 18376 -2930 18484 -2924
rect 18634 -2890 18742 -2884
rect 18634 -2924 18646 -2890
rect 18730 -2924 18742 -2890
rect 18634 -2930 18742 -2924
rect 18272 -3004 18284 -2974
rect 18060 -3350 18074 -3306
rect 17602 -3400 17710 -3394
rect 17602 -3434 17614 -3400
rect 17698 -3434 17710 -3400
rect 17602 -3440 17710 -3434
rect 17860 -3400 17968 -3394
rect 17860 -3434 17872 -3400
rect 17956 -3434 17968 -3400
rect 17860 -3440 17968 -3434
rect 17880 -3490 17940 -3440
rect 17874 -3550 17880 -3490
rect 17940 -3550 17946 -3490
rect 17490 -3660 17496 -3600
rect 17556 -3660 17562 -3600
rect 18014 -3716 18074 -3350
rect 18278 -3350 18284 -3004
rect 18318 -3004 18332 -2974
rect 18536 -2974 18582 -2962
rect 18318 -3350 18324 -3004
rect 18536 -3300 18542 -2974
rect 18278 -3362 18324 -3350
rect 18532 -3350 18542 -3300
rect 18576 -3300 18582 -2974
rect 18790 -2974 18850 -2818
rect 18576 -3350 18592 -3300
rect 18118 -3400 18226 -3394
rect 18118 -3434 18130 -3400
rect 18214 -3434 18226 -3400
rect 18118 -3440 18226 -3434
rect 18376 -3400 18484 -3394
rect 18376 -3434 18388 -3400
rect 18472 -3434 18484 -3400
rect 18376 -3440 18484 -3434
rect 18142 -3490 18202 -3440
rect 18136 -3550 18142 -3490
rect 18202 -3550 18208 -3490
rect 18532 -3600 18592 -3350
rect 18790 -3350 18800 -2974
rect 18834 -3350 18850 -2974
rect 18634 -3400 18742 -3394
rect 18634 -3434 18646 -3400
rect 18730 -3434 18742 -3400
rect 18634 -3440 18742 -3434
rect 18658 -3490 18718 -3440
rect 18790 -3490 18850 -3350
rect 19506 -2974 19566 -2818
rect 19632 -2884 19692 -2818
rect 19890 -2884 19950 -2814
rect 19608 -2890 19716 -2884
rect 19608 -2924 19620 -2890
rect 19704 -2924 19716 -2890
rect 19608 -2930 19716 -2924
rect 19866 -2890 19974 -2884
rect 19866 -2924 19878 -2890
rect 19962 -2924 19974 -2890
rect 19866 -2930 19974 -2924
rect 19506 -3350 19516 -2974
rect 19550 -3350 19566 -2974
rect 19768 -2974 19814 -2962
rect 19768 -3300 19774 -2974
rect 19506 -3490 19566 -3350
rect 19760 -3350 19774 -3300
rect 19808 -3300 19814 -2974
rect 20020 -2974 20080 -2704
rect 20124 -2890 20232 -2884
rect 20124 -2924 20136 -2890
rect 20220 -2924 20232 -2890
rect 20124 -2930 20232 -2924
rect 20382 -2890 20490 -2884
rect 20382 -2924 20394 -2890
rect 20478 -2924 20490 -2890
rect 20382 -2930 20490 -2924
rect 20020 -2994 20032 -2974
rect 19808 -3350 19820 -3300
rect 19608 -3400 19716 -3394
rect 19608 -3434 19620 -3400
rect 19704 -3434 19716 -3400
rect 19608 -3440 19716 -3434
rect 19630 -3490 19690 -3440
rect 18658 -3550 19690 -3490
rect 18526 -3660 18532 -3600
rect 18592 -3660 18598 -3600
rect 16972 -3776 16978 -3716
rect 17038 -3776 17044 -3716
rect 18008 -3776 18014 -3716
rect 18074 -3776 18080 -3716
rect 18658 -3816 18718 -3550
rect 18790 -3816 18850 -3550
rect 19506 -3816 19566 -3550
rect 19630 -3816 19690 -3550
rect 19760 -3594 19820 -3350
rect 20026 -3350 20032 -2994
rect 20066 -2994 20080 -2974
rect 20284 -2974 20330 -2962
rect 20066 -3350 20072 -2994
rect 20284 -3304 20290 -2974
rect 20026 -3362 20072 -3350
rect 20274 -3350 20290 -3304
rect 20324 -3304 20330 -2974
rect 20532 -2974 20592 -2704
rect 20660 -2814 20666 -2754
rect 20726 -2814 20732 -2754
rect 20914 -2814 20920 -2754
rect 20980 -2814 20986 -2754
rect 20666 -2884 20726 -2814
rect 20920 -2884 20980 -2814
rect 20640 -2890 20748 -2884
rect 20640 -2924 20652 -2890
rect 20736 -2924 20748 -2890
rect 20640 -2930 20748 -2924
rect 20898 -2890 21006 -2884
rect 20898 -2924 20910 -2890
rect 20994 -2924 21006 -2890
rect 20898 -2930 21006 -2924
rect 20532 -2994 20548 -2974
rect 20324 -3350 20334 -3304
rect 19866 -3400 19974 -3394
rect 19866 -3434 19878 -3400
rect 19962 -3434 19974 -3400
rect 19866 -3440 19974 -3434
rect 20124 -3400 20232 -3394
rect 20124 -3434 20136 -3400
rect 20220 -3434 20232 -3400
rect 20124 -3440 20232 -3434
rect 20150 -3484 20210 -3440
rect 20144 -3544 20150 -3484
rect 20210 -3544 20216 -3484
rect 19754 -3654 19760 -3594
rect 19820 -3654 19826 -3594
rect 20274 -3710 20334 -3350
rect 20542 -3350 20548 -2994
rect 20582 -2994 20592 -2974
rect 20800 -2974 20846 -2962
rect 20582 -3350 20588 -2994
rect 20800 -3290 20806 -2974
rect 20542 -3362 20588 -3350
rect 20792 -3350 20806 -3290
rect 20840 -3290 20846 -2974
rect 21052 -2974 21112 -2704
rect 21156 -2890 21264 -2884
rect 21156 -2924 21168 -2890
rect 21252 -2924 21264 -2890
rect 21156 -2930 21264 -2924
rect 21414 -2890 21522 -2884
rect 21414 -2924 21426 -2890
rect 21510 -2924 21522 -2890
rect 21414 -2930 21522 -2924
rect 21052 -2998 21064 -2974
rect 20840 -3350 20852 -3290
rect 20382 -3400 20490 -3394
rect 20382 -3434 20394 -3400
rect 20478 -3434 20490 -3400
rect 20382 -3440 20490 -3434
rect 20640 -3400 20748 -3394
rect 20640 -3434 20652 -3400
rect 20736 -3434 20748 -3400
rect 20640 -3440 20748 -3434
rect 20404 -3484 20464 -3440
rect 20398 -3544 20404 -3484
rect 20464 -3544 20470 -3484
rect 20792 -3594 20852 -3350
rect 21058 -3350 21064 -2998
rect 21098 -2998 21112 -2974
rect 21316 -2974 21362 -2962
rect 21098 -3350 21104 -2998
rect 21316 -3300 21322 -2974
rect 21058 -3362 21104 -3350
rect 21310 -3350 21322 -3300
rect 21356 -3300 21362 -2974
rect 21568 -2974 21628 -2704
rect 22232 -2752 22292 -2444
rect 22656 -2752 22716 -2444
rect 22788 -2644 22848 -1376
rect 22782 -2704 22788 -2644
rect 22848 -2704 22854 -2644
rect 23104 -2752 23110 -778
rect 21692 -2814 21698 -2754
rect 21758 -2814 21764 -2754
rect 21952 -2812 23110 -2752
rect 21698 -2884 21758 -2814
rect 21952 -2884 22012 -2812
rect 21672 -2890 21780 -2884
rect 21672 -2924 21684 -2890
rect 21768 -2924 21780 -2890
rect 21672 -2930 21780 -2924
rect 21930 -2890 22038 -2884
rect 21930 -2924 21942 -2890
rect 22026 -2924 22038 -2890
rect 21930 -2930 22038 -2924
rect 21568 -2998 21580 -2974
rect 21356 -3350 21370 -3300
rect 21176 -3394 21236 -3390
rect 20898 -3400 21006 -3394
rect 20898 -3434 20910 -3400
rect 20994 -3434 21006 -3400
rect 20898 -3440 21006 -3434
rect 21156 -3400 21264 -3394
rect 21156 -3434 21168 -3400
rect 21252 -3434 21264 -3400
rect 21156 -3440 21264 -3434
rect 21176 -3484 21236 -3440
rect 21170 -3544 21176 -3484
rect 21236 -3544 21242 -3484
rect 20786 -3654 20792 -3594
rect 20852 -3654 20858 -3594
rect 21310 -3710 21370 -3350
rect 21574 -3350 21580 -2998
rect 21614 -2998 21628 -2974
rect 21832 -2974 21878 -2962
rect 21614 -3350 21620 -2998
rect 21832 -3294 21838 -2974
rect 21574 -3362 21620 -3350
rect 21828 -3350 21838 -3294
rect 21872 -3294 21878 -2974
rect 22086 -2974 22146 -2812
rect 21872 -3350 21888 -3294
rect 21414 -3400 21522 -3394
rect 21414 -3434 21426 -3400
rect 21510 -3434 21522 -3400
rect 21414 -3440 21522 -3434
rect 21672 -3400 21780 -3394
rect 21672 -3434 21684 -3400
rect 21768 -3434 21780 -3400
rect 21672 -3440 21780 -3434
rect 21438 -3484 21498 -3440
rect 21432 -3544 21438 -3484
rect 21498 -3544 21504 -3484
rect 21828 -3594 21888 -3350
rect 22086 -3350 22096 -2974
rect 22130 -3350 22146 -2974
rect 21930 -3400 22038 -3394
rect 21930 -3434 21942 -3400
rect 22026 -3434 22038 -3400
rect 21930 -3440 22038 -3434
rect 21954 -3482 22014 -3440
rect 22086 -3482 22146 -3350
rect 23104 -3482 23110 -2812
rect 21954 -3542 23110 -3482
rect 21822 -3654 21828 -3594
rect 21888 -3654 21894 -3594
rect 20268 -3770 20274 -3710
rect 20334 -3770 20340 -3710
rect 21304 -3770 21310 -3710
rect 21370 -3770 21376 -3710
rect 21954 -3816 22014 -3542
rect 22086 -3816 22146 -3542
rect 23104 -3662 23110 -3542
rect 23210 -3662 23216 -778
rect 23104 -3816 23216 -3662
rect 11860 -3822 23216 -3816
rect 11860 -3922 11966 -3822
rect 23110 -3922 23216 -3822
rect 11860 -3928 23216 -3922
rect 3440 -4004 3500 -3998
rect 6088 -4004 6148 -3998
rect 8476 -4004 8536 -3998
rect 3500 -4064 6088 -4004
rect 6148 -4064 8476 -4004
rect 3440 -4070 3500 -4064
rect 6088 -4070 6148 -4064
rect 8476 -4070 8536 -4064
rect 15240 -4004 15300 -3998
rect 17888 -4004 17948 -3998
rect 20276 -4004 20336 -3998
rect 15300 -4064 17888 -4004
rect 17948 -4064 20276 -4004
rect 15240 -4070 15300 -4064
rect 17888 -4070 17948 -4064
rect 20276 -4070 20336 -4064
rect 60 -4158 11416 -4152
rect 60 -4258 166 -4158
rect 11310 -4258 11416 -4158
rect 60 -4264 11416 -4258
rect 60 -4318 172 -4264
rect 60 -5782 66 -4318
rect 166 -5782 172 -4318
rect 3892 -4436 3952 -4264
rect 4024 -4436 4084 -4264
rect 4668 -4322 4728 -4316
rect 3892 -4496 4084 -4436
rect 3892 -4642 3952 -4496
rect 4024 -4543 4084 -4496
rect 4152 -4492 4540 -4432
rect 4600 -4492 4606 -4432
rect 4000 -4549 4108 -4543
rect 4000 -4583 4012 -4549
rect 4096 -4583 4108 -4549
rect 4000 -4589 4108 -4583
rect 3892 -4818 3908 -4642
rect 3942 -4818 3952 -4642
rect 4152 -4642 4212 -4492
rect 4284 -4543 4344 -4492
rect 4540 -4543 4600 -4492
rect 4258 -4549 4366 -4543
rect 4258 -4583 4270 -4549
rect 4354 -4583 4366 -4549
rect 4258 -4589 4366 -4583
rect 4516 -4549 4624 -4543
rect 4516 -4583 4528 -4549
rect 4612 -4583 4624 -4549
rect 4516 -4589 4624 -4583
rect 4152 -4682 4166 -4642
rect 3892 -4983 3952 -4818
rect 4160 -4818 4166 -4682
rect 4200 -4682 4212 -4642
rect 4418 -4642 4464 -4630
rect 4200 -4818 4206 -4682
rect 4418 -4788 4424 -4642
rect 4160 -4830 4206 -4818
rect 4410 -4818 4424 -4788
rect 4458 -4788 4464 -4642
rect 4668 -4642 4728 -4382
rect 4774 -4549 4882 -4543
rect 4774 -4583 4786 -4549
rect 4870 -4583 4882 -4549
rect 4774 -4589 4882 -4583
rect 4668 -4665 4682 -4642
rect 4458 -4818 4470 -4788
rect 4000 -4877 4108 -4871
rect 4000 -4911 4012 -4877
rect 4096 -4911 4108 -4877
rect 4000 -4917 4108 -4911
rect 4258 -4877 4366 -4871
rect 4258 -4911 4270 -4877
rect 4354 -4911 4366 -4877
rect 4258 -4917 4366 -4911
rect 4028 -4983 4088 -4917
rect 3892 -5043 4088 -4983
rect 3892 -5260 3952 -5043
rect 4028 -5260 4088 -5043
rect 4410 -5260 4470 -4818
rect 4676 -4818 4682 -4665
rect 4716 -4665 4728 -4642
rect 4926 -4642 4986 -4264
rect 5182 -4320 5242 -4314
rect 5050 -4492 5056 -4432
rect 5116 -4492 5122 -4432
rect 5056 -4543 5116 -4492
rect 5032 -4549 5140 -4543
rect 5032 -4583 5044 -4549
rect 5128 -4583 5140 -4549
rect 5032 -4589 5140 -4583
rect 4716 -4818 4722 -4665
rect 4676 -4830 4722 -4818
rect 4926 -4818 4940 -4642
rect 4974 -4818 4986 -4642
rect 5182 -4642 5242 -4380
rect 5314 -4436 5374 -4264
rect 5442 -4436 5502 -4264
rect 5570 -4436 5630 -4264
rect 6088 -4318 6148 -4312
rect 6088 -4430 6148 -4378
rect 6344 -4430 6404 -4264
rect 6474 -4430 6534 -4264
rect 6598 -4430 6658 -4264
rect 5314 -4496 5630 -4436
rect 5314 -4543 5374 -4496
rect 5290 -4549 5398 -4543
rect 5290 -4583 5302 -4549
rect 5386 -4583 5398 -4549
rect 5290 -4589 5398 -4583
rect 5182 -4697 5198 -4642
rect 4516 -4877 4624 -4871
rect 4516 -4911 4528 -4877
rect 4612 -4911 4624 -4877
rect 4516 -4917 4624 -4911
rect 4774 -4877 4882 -4871
rect 4774 -4911 4786 -4877
rect 4870 -4911 4882 -4877
rect 4774 -4917 4882 -4911
rect 4800 -4978 4860 -4917
rect 4926 -4978 4986 -4818
rect 5192 -4818 5198 -4697
rect 5232 -4697 5242 -4642
rect 5442 -4642 5502 -4496
rect 5570 -4543 5630 -4496
rect 5828 -4490 6274 -4430
rect 5828 -4543 5888 -4490
rect 6088 -4543 6148 -4490
rect 5548 -4549 5656 -4543
rect 5548 -4583 5560 -4549
rect 5644 -4583 5656 -4549
rect 5548 -4589 5656 -4583
rect 5806 -4549 5914 -4543
rect 5806 -4583 5818 -4549
rect 5902 -4583 5914 -4549
rect 5806 -4589 5914 -4583
rect 6064 -4549 6172 -4543
rect 6064 -4583 6076 -4549
rect 6160 -4583 6172 -4549
rect 6064 -4589 6172 -4583
rect 5232 -4818 5238 -4697
rect 5192 -4830 5238 -4818
rect 5442 -4818 5456 -4642
rect 5490 -4818 5502 -4642
rect 5708 -4642 5754 -4630
rect 5708 -4778 5714 -4642
rect 5032 -4877 5140 -4871
rect 5032 -4911 5044 -4877
rect 5128 -4911 5140 -4877
rect 5032 -4917 5140 -4911
rect 5290 -4877 5398 -4871
rect 5290 -4911 5302 -4877
rect 5386 -4911 5398 -4877
rect 5290 -4917 5398 -4911
rect 4800 -5038 4986 -4978
rect 4800 -5260 4860 -5038
rect 4926 -5260 4986 -5038
rect 5314 -4983 5374 -4917
rect 5442 -4983 5502 -4818
rect 5696 -4818 5714 -4778
rect 5748 -4778 5754 -4642
rect 5966 -4642 6012 -4630
rect 5748 -4818 5756 -4778
rect 5966 -4788 5972 -4642
rect 5548 -4877 5656 -4871
rect 5548 -4911 5560 -4877
rect 5644 -4911 5656 -4877
rect 5548 -4917 5656 -4911
rect 5566 -4983 5626 -4917
rect 5314 -5043 5626 -4983
rect 5314 -5260 5374 -5043
rect 5442 -5260 5502 -5043
rect 5566 -5260 5626 -5043
rect 5696 -5096 5756 -4818
rect 5956 -4818 5972 -4788
rect 6006 -4788 6012 -4642
rect 6214 -4642 6274 -4490
rect 6344 -4490 6658 -4430
rect 6344 -4543 6404 -4490
rect 6322 -4549 6430 -4543
rect 6322 -4583 6334 -4549
rect 6418 -4583 6430 -4549
rect 6322 -4589 6430 -4583
rect 6214 -4680 6230 -4642
rect 6006 -4818 6016 -4788
rect 5806 -4877 5914 -4871
rect 5806 -4911 5818 -4877
rect 5902 -4911 5914 -4877
rect 5806 -4917 5914 -4911
rect 5690 -5156 5696 -5096
rect 5756 -5156 5762 -5096
rect 5956 -5260 6016 -4818
rect 6224 -4818 6230 -4680
rect 6264 -4680 6274 -4642
rect 6474 -4642 6534 -4490
rect 6598 -4543 6658 -4490
rect 6734 -4488 6920 -4428
rect 6580 -4549 6688 -4543
rect 6580 -4583 6592 -4549
rect 6676 -4583 6688 -4549
rect 6580 -4589 6688 -4583
rect 6264 -4818 6270 -4680
rect 6224 -4830 6270 -4818
rect 6474 -4818 6488 -4642
rect 6522 -4818 6534 -4642
rect 6064 -4877 6172 -4871
rect 6064 -4911 6076 -4877
rect 6160 -4911 6172 -4877
rect 6064 -4917 6172 -4911
rect 6322 -4877 6430 -4871
rect 6322 -4911 6334 -4877
rect 6418 -4911 6430 -4877
rect 6322 -4917 6430 -4911
rect 6346 -4977 6406 -4917
rect 6474 -4977 6534 -4818
rect 6734 -4642 6794 -4488
rect 6860 -4543 6920 -4488
rect 6838 -4549 6946 -4543
rect 6838 -4583 6850 -4549
rect 6934 -4583 6946 -4549
rect 6838 -4589 6946 -4583
rect 6734 -4818 6746 -4642
rect 6780 -4818 6794 -4642
rect 6580 -4877 6688 -4871
rect 6580 -4911 6592 -4877
rect 6676 -4911 6688 -4877
rect 6580 -4917 6688 -4911
rect 6606 -4977 6666 -4917
rect 6734 -4974 6794 -4818
rect 6990 -4642 7050 -4264
rect 7246 -4376 7252 -4316
rect 7312 -4376 7318 -4316
rect 7252 -4428 7312 -4376
rect 7124 -4488 7312 -4428
rect 7124 -4543 7184 -4488
rect 7096 -4549 7204 -4543
rect 7096 -4583 7108 -4549
rect 7192 -4583 7204 -4549
rect 7096 -4589 7204 -4583
rect 6990 -4818 7004 -4642
rect 7038 -4818 7050 -4642
rect 7252 -4642 7312 -4488
rect 7376 -4432 7436 -4264
rect 7506 -4432 7566 -4264
rect 7376 -4492 7566 -4432
rect 7376 -4543 7436 -4492
rect 7354 -4549 7462 -4543
rect 7354 -4583 7366 -4549
rect 7450 -4583 7462 -4549
rect 7354 -4589 7462 -4583
rect 7252 -4688 7262 -4642
rect 6838 -4877 6946 -4871
rect 6838 -4911 6850 -4877
rect 6934 -4911 6946 -4877
rect 6838 -4917 6946 -4911
rect 6346 -5037 6666 -4977
rect 6728 -5034 6734 -4974
rect 6794 -5034 6800 -4974
rect 6346 -5260 6406 -5037
rect 6474 -5260 6534 -5037
rect 6606 -5260 6666 -5037
rect 6990 -5260 7050 -4818
rect 7256 -4818 7262 -4688
rect 7296 -4688 7312 -4642
rect 7506 -4642 7566 -4492
rect 7296 -4818 7302 -4688
rect 7256 -4830 7302 -4818
rect 7506 -4818 7520 -4642
rect 7554 -4818 7566 -4642
rect 7096 -4877 7204 -4871
rect 7096 -4911 7108 -4877
rect 7192 -4911 7204 -4877
rect 7096 -4917 7204 -4911
rect 7354 -4877 7462 -4871
rect 7354 -4911 7366 -4877
rect 7450 -4911 7462 -4877
rect 7354 -4917 7462 -4911
rect 7376 -4976 7436 -4917
rect 7506 -4976 7566 -4818
rect 7376 -5036 7566 -4976
rect 7376 -5260 7436 -5036
rect 7506 -5260 7566 -5036
rect 11304 -4318 11416 -4264
rect 3854 -5298 7710 -5260
rect 3854 -5450 3902 -5298
rect 7666 -5450 7710 -5298
rect 3854 -5490 7710 -5450
rect 60 -5836 172 -5782
rect 772 -5836 782 -5536
rect 10694 -5836 10704 -5536
rect 11304 -5782 11310 -4318
rect 11410 -5782 11416 -4318
rect 11304 -5836 11416 -5782
rect 60 -5842 11416 -5836
rect 60 -5942 166 -5842
rect 11310 -5942 11416 -5842
rect 60 -5948 11416 -5942
rect 11860 -4158 23216 -4152
rect 11860 -4258 11966 -4158
rect 23110 -4258 23216 -4158
rect 11860 -4264 23216 -4258
rect 11860 -4318 11972 -4264
rect 11860 -5782 11866 -4318
rect 11966 -5782 11972 -4318
rect 15692 -4436 15752 -4264
rect 15824 -4436 15884 -4264
rect 16468 -4322 16528 -4316
rect 15692 -4496 15884 -4436
rect 15692 -4642 15752 -4496
rect 15824 -4543 15884 -4496
rect 15952 -4492 16340 -4432
rect 16400 -4492 16406 -4432
rect 15800 -4549 15908 -4543
rect 15800 -4583 15812 -4549
rect 15896 -4583 15908 -4549
rect 15800 -4589 15908 -4583
rect 15692 -4818 15708 -4642
rect 15742 -4818 15752 -4642
rect 15952 -4642 16012 -4492
rect 16084 -4543 16144 -4492
rect 16340 -4543 16400 -4492
rect 16058 -4549 16166 -4543
rect 16058 -4583 16070 -4549
rect 16154 -4583 16166 -4549
rect 16058 -4589 16166 -4583
rect 16316 -4549 16424 -4543
rect 16316 -4583 16328 -4549
rect 16412 -4583 16424 -4549
rect 16316 -4589 16424 -4583
rect 15952 -4682 15966 -4642
rect 15692 -4983 15752 -4818
rect 15960 -4818 15966 -4682
rect 16000 -4682 16012 -4642
rect 16218 -4642 16264 -4630
rect 16000 -4818 16006 -4682
rect 16218 -4788 16224 -4642
rect 15960 -4830 16006 -4818
rect 16210 -4818 16224 -4788
rect 16258 -4788 16264 -4642
rect 16468 -4642 16528 -4382
rect 16574 -4549 16682 -4543
rect 16574 -4583 16586 -4549
rect 16670 -4583 16682 -4549
rect 16574 -4589 16682 -4583
rect 16468 -4665 16482 -4642
rect 16258 -4818 16270 -4788
rect 15800 -4877 15908 -4871
rect 15800 -4911 15812 -4877
rect 15896 -4911 15908 -4877
rect 15800 -4917 15908 -4911
rect 16058 -4877 16166 -4871
rect 16058 -4911 16070 -4877
rect 16154 -4911 16166 -4877
rect 16058 -4917 16166 -4911
rect 15828 -4983 15888 -4917
rect 15692 -5043 15888 -4983
rect 15692 -5260 15752 -5043
rect 15828 -5260 15888 -5043
rect 16210 -5260 16270 -4818
rect 16476 -4818 16482 -4665
rect 16516 -4665 16528 -4642
rect 16726 -4642 16786 -4264
rect 16982 -4320 17042 -4314
rect 16850 -4492 16856 -4432
rect 16916 -4492 16922 -4432
rect 16856 -4543 16916 -4492
rect 16832 -4549 16940 -4543
rect 16832 -4583 16844 -4549
rect 16928 -4583 16940 -4549
rect 16832 -4589 16940 -4583
rect 16516 -4818 16522 -4665
rect 16476 -4830 16522 -4818
rect 16726 -4818 16740 -4642
rect 16774 -4818 16786 -4642
rect 16982 -4642 17042 -4380
rect 17114 -4436 17174 -4264
rect 17242 -4436 17302 -4264
rect 17370 -4436 17430 -4264
rect 17888 -4318 17948 -4312
rect 17888 -4430 17948 -4378
rect 18144 -4430 18204 -4264
rect 18274 -4430 18334 -4264
rect 18398 -4430 18458 -4264
rect 17114 -4496 17430 -4436
rect 17114 -4543 17174 -4496
rect 17090 -4549 17198 -4543
rect 17090 -4583 17102 -4549
rect 17186 -4583 17198 -4549
rect 17090 -4589 17198 -4583
rect 16982 -4697 16998 -4642
rect 16316 -4877 16424 -4871
rect 16316 -4911 16328 -4877
rect 16412 -4911 16424 -4877
rect 16316 -4917 16424 -4911
rect 16574 -4877 16682 -4871
rect 16574 -4911 16586 -4877
rect 16670 -4911 16682 -4877
rect 16574 -4917 16682 -4911
rect 16600 -4978 16660 -4917
rect 16726 -4978 16786 -4818
rect 16992 -4818 16998 -4697
rect 17032 -4697 17042 -4642
rect 17242 -4642 17302 -4496
rect 17370 -4543 17430 -4496
rect 17628 -4490 18074 -4430
rect 17628 -4543 17688 -4490
rect 17888 -4543 17948 -4490
rect 17348 -4549 17456 -4543
rect 17348 -4583 17360 -4549
rect 17444 -4583 17456 -4549
rect 17348 -4589 17456 -4583
rect 17606 -4549 17714 -4543
rect 17606 -4583 17618 -4549
rect 17702 -4583 17714 -4549
rect 17606 -4589 17714 -4583
rect 17864 -4549 17972 -4543
rect 17864 -4583 17876 -4549
rect 17960 -4583 17972 -4549
rect 17864 -4589 17972 -4583
rect 17032 -4818 17038 -4697
rect 16992 -4830 17038 -4818
rect 17242 -4818 17256 -4642
rect 17290 -4818 17302 -4642
rect 17508 -4642 17554 -4630
rect 17508 -4778 17514 -4642
rect 16832 -4877 16940 -4871
rect 16832 -4911 16844 -4877
rect 16928 -4911 16940 -4877
rect 16832 -4917 16940 -4911
rect 17090 -4877 17198 -4871
rect 17090 -4911 17102 -4877
rect 17186 -4911 17198 -4877
rect 17090 -4917 17198 -4911
rect 16600 -5038 16786 -4978
rect 16600 -5260 16660 -5038
rect 16726 -5260 16786 -5038
rect 17114 -4983 17174 -4917
rect 17242 -4983 17302 -4818
rect 17496 -4818 17514 -4778
rect 17548 -4778 17554 -4642
rect 17766 -4642 17812 -4630
rect 17548 -4818 17556 -4778
rect 17766 -4788 17772 -4642
rect 17348 -4877 17456 -4871
rect 17348 -4911 17360 -4877
rect 17444 -4911 17456 -4877
rect 17348 -4917 17456 -4911
rect 17366 -4983 17426 -4917
rect 17114 -5043 17426 -4983
rect 17114 -5260 17174 -5043
rect 17242 -5260 17302 -5043
rect 17366 -5260 17426 -5043
rect 17496 -5096 17556 -4818
rect 17756 -4818 17772 -4788
rect 17806 -4788 17812 -4642
rect 18014 -4642 18074 -4490
rect 18144 -4490 18458 -4430
rect 18144 -4543 18204 -4490
rect 18122 -4549 18230 -4543
rect 18122 -4583 18134 -4549
rect 18218 -4583 18230 -4549
rect 18122 -4589 18230 -4583
rect 18014 -4680 18030 -4642
rect 17806 -4818 17816 -4788
rect 17606 -4877 17714 -4871
rect 17606 -4911 17618 -4877
rect 17702 -4911 17714 -4877
rect 17606 -4917 17714 -4911
rect 17490 -5156 17496 -5096
rect 17556 -5156 17562 -5096
rect 17756 -5260 17816 -4818
rect 18024 -4818 18030 -4680
rect 18064 -4680 18074 -4642
rect 18274 -4642 18334 -4490
rect 18398 -4543 18458 -4490
rect 18534 -4488 18720 -4428
rect 18380 -4549 18488 -4543
rect 18380 -4583 18392 -4549
rect 18476 -4583 18488 -4549
rect 18380 -4589 18488 -4583
rect 18064 -4818 18070 -4680
rect 18024 -4830 18070 -4818
rect 18274 -4818 18288 -4642
rect 18322 -4818 18334 -4642
rect 17864 -4877 17972 -4871
rect 17864 -4911 17876 -4877
rect 17960 -4911 17972 -4877
rect 17864 -4917 17972 -4911
rect 18122 -4877 18230 -4871
rect 18122 -4911 18134 -4877
rect 18218 -4911 18230 -4877
rect 18122 -4917 18230 -4911
rect 18146 -4977 18206 -4917
rect 18274 -4977 18334 -4818
rect 18534 -4642 18594 -4488
rect 18660 -4543 18720 -4488
rect 18638 -4549 18746 -4543
rect 18638 -4583 18650 -4549
rect 18734 -4583 18746 -4549
rect 18638 -4589 18746 -4583
rect 18534 -4818 18546 -4642
rect 18580 -4818 18594 -4642
rect 18380 -4877 18488 -4871
rect 18380 -4911 18392 -4877
rect 18476 -4911 18488 -4877
rect 18380 -4917 18488 -4911
rect 18406 -4977 18466 -4917
rect 18534 -4974 18594 -4818
rect 18790 -4642 18850 -4264
rect 19046 -4376 19052 -4316
rect 19112 -4376 19118 -4316
rect 19052 -4428 19112 -4376
rect 18924 -4488 19112 -4428
rect 18924 -4543 18984 -4488
rect 18896 -4549 19004 -4543
rect 18896 -4583 18908 -4549
rect 18992 -4583 19004 -4549
rect 18896 -4589 19004 -4583
rect 18790 -4818 18804 -4642
rect 18838 -4818 18850 -4642
rect 19052 -4642 19112 -4488
rect 19176 -4432 19236 -4264
rect 19306 -4432 19366 -4264
rect 19176 -4492 19366 -4432
rect 19176 -4543 19236 -4492
rect 19154 -4549 19262 -4543
rect 19154 -4583 19166 -4549
rect 19250 -4583 19262 -4549
rect 19154 -4589 19262 -4583
rect 19052 -4688 19062 -4642
rect 18638 -4877 18746 -4871
rect 18638 -4911 18650 -4877
rect 18734 -4911 18746 -4877
rect 18638 -4917 18746 -4911
rect 18146 -5037 18466 -4977
rect 18528 -5034 18534 -4974
rect 18594 -5034 18600 -4974
rect 18146 -5260 18206 -5037
rect 18274 -5260 18334 -5037
rect 18406 -5260 18466 -5037
rect 18790 -5260 18850 -4818
rect 19056 -4818 19062 -4688
rect 19096 -4688 19112 -4642
rect 19306 -4642 19366 -4492
rect 19096 -4818 19102 -4688
rect 19056 -4830 19102 -4818
rect 19306 -4818 19320 -4642
rect 19354 -4818 19366 -4642
rect 18896 -4877 19004 -4871
rect 18896 -4911 18908 -4877
rect 18992 -4911 19004 -4877
rect 18896 -4917 19004 -4911
rect 19154 -4877 19262 -4871
rect 19154 -4911 19166 -4877
rect 19250 -4911 19262 -4877
rect 19154 -4917 19262 -4911
rect 19176 -4976 19236 -4917
rect 19306 -4976 19366 -4818
rect 19176 -5036 19366 -4976
rect 19176 -5260 19236 -5036
rect 19306 -5260 19366 -5036
rect 23104 -4318 23216 -4264
rect 15654 -5298 19510 -5260
rect 15654 -5450 15702 -5298
rect 19466 -5450 19510 -5298
rect 15654 -5490 19510 -5450
rect 11860 -5836 11972 -5782
rect 12572 -5836 12582 -5536
rect 22494 -5836 22504 -5536
rect 23104 -5782 23110 -4318
rect 23210 -5782 23216 -4318
rect 23104 -5836 23216 -5782
rect 11860 -5842 23216 -5836
rect 11860 -5942 11966 -5842
rect 23110 -5942 23216 -5842
rect 11860 -5948 23216 -5942
<< via1 >>
rect 172 4732 772 5032
rect 10704 4732 11304 5032
rect 3902 4494 7666 4646
rect 5696 4292 5756 4352
rect 4540 3628 4600 3688
rect 4668 3518 4728 3578
rect 5056 3628 5116 3688
rect 5182 3516 5242 3576
rect 6734 4170 6794 4230
rect 6088 3514 6148 3574
rect 7252 3512 7312 3572
rect 11972 4732 12572 5032
rect 22504 4732 23104 5032
rect 15702 4494 19466 4646
rect 17496 4292 17556 4352
rect 16340 3628 16400 3688
rect 16468 3518 16528 3578
rect 16856 3628 16916 3688
rect 16982 3516 17042 3576
rect 18534 4170 18594 4230
rect 17888 3514 17948 3574
rect 19052 3512 19112 3572
rect 3440 3200 3500 3260
rect 6088 3200 6148 3260
rect 8476 3200 8536 3260
rect 15240 3200 15300 3260
rect 17888 3200 17948 3260
rect 20276 3200 20336 3260
rect 1882 2906 1942 2966
rect 2918 2906 2978 2966
rect 1368 2790 1428 2850
rect 1758 2680 1818 2740
rect 2400 2790 2460 2850
rect 2012 2680 2072 2740
rect 1498 1950 1558 2010
rect 420 1840 480 1900
rect 2784 2680 2844 2740
rect 3436 2790 3496 2850
rect 3046 2680 3106 2740
rect 2274 1950 2334 2010
rect 2528 1950 2588 2010
rect 5178 2912 5238 2972
rect 6214 2912 6274 2972
rect 4664 2796 4724 2856
rect 3306 1950 3366 2010
rect 5054 2686 5114 2746
rect 5696 2796 5756 2856
rect 5308 2686 5368 2746
rect 1628 1840 1688 1900
rect 2140 1840 2200 1900
rect 2660 1840 2720 1900
rect 3176 1840 3236 1900
rect 4794 1956 4854 2016
rect 3306 1718 3366 1778
rect 1418 1594 1478 1654
rect 1420 1050 1480 1110
rect 4924 1846 4984 1906
rect 6080 2686 6140 2746
rect 6732 2796 6792 2856
rect 6342 2686 6402 2746
rect 5570 1956 5630 2016
rect 5824 1956 5884 2016
rect 8474 2906 8534 2966
rect 9510 2906 9570 2966
rect 7960 2790 8020 2850
rect 6602 1956 6662 2016
rect 8350 2680 8410 2740
rect 8992 2790 9052 2850
rect 8604 2680 8664 2740
rect 5436 1846 5496 1906
rect 5956 1846 6016 1906
rect 6472 1846 6532 1906
rect 5186 1718 5246 1778
rect 4852 1594 4912 1654
rect 2702 1054 2762 1110
rect 3136 1050 3196 1110
rect 3566 1054 3626 1110
rect 420 506 480 566
rect 8090 1950 8150 2010
rect 9376 2680 9436 2740
rect 10028 2790 10088 2850
rect 9638 2680 9698 2740
rect 8866 1950 8926 2010
rect 9120 1950 9180 2010
rect 9898 1950 9958 2010
rect 8220 1840 8280 1900
rect 8732 1840 8792 1900
rect 9252 1840 9312 1900
rect 9768 1840 9828 1900
rect 10002 1710 10062 1770
rect 4426 1054 4486 1110
rect 4856 1050 4916 1110
rect 6572 1050 6632 1110
rect 6998 1054 7058 1110
rect 10988 1840 11048 1900
rect 7856 1054 7916 1110
rect 8284 1050 8344 1110
rect 8710 1054 8770 1110
rect 6568 506 6628 566
rect 9576 1050 9636 1110
rect 10000 512 10060 572
rect 10988 512 11048 572
rect 384 242 11040 352
rect 172 -180 772 120
rect 10704 -180 11304 120
rect 13682 2906 13742 2966
rect 14718 2906 14778 2966
rect 13168 2790 13228 2850
rect 13558 2680 13618 2740
rect 14200 2790 14260 2850
rect 13812 2680 13872 2740
rect 13298 1950 13358 2010
rect 12220 1840 12280 1900
rect 14584 2680 14644 2740
rect 15236 2790 15296 2850
rect 14846 2680 14906 2740
rect 14074 1950 14134 2010
rect 14328 1950 14388 2010
rect 16978 2912 17038 2972
rect 18014 2912 18074 2972
rect 16464 2796 16524 2856
rect 15106 1950 15166 2010
rect 16854 2686 16914 2746
rect 17496 2796 17556 2856
rect 17108 2686 17168 2746
rect 13428 1840 13488 1900
rect 13940 1840 14000 1900
rect 14460 1840 14520 1900
rect 14976 1840 15036 1900
rect 16594 1956 16654 2016
rect 15106 1718 15166 1778
rect 13218 1594 13278 1654
rect 13220 1050 13280 1110
rect 16724 1846 16784 1906
rect 17880 2686 17940 2746
rect 18532 2796 18592 2856
rect 18142 2686 18202 2746
rect 17370 1956 17430 2016
rect 17624 1956 17684 2016
rect 20274 2906 20334 2966
rect 21310 2906 21370 2966
rect 19760 2790 19820 2850
rect 18402 1956 18462 2016
rect 20150 2680 20210 2740
rect 20792 2790 20852 2850
rect 20404 2680 20464 2740
rect 17236 1846 17296 1906
rect 17756 1846 17816 1906
rect 18272 1846 18332 1906
rect 16986 1718 17046 1778
rect 16652 1594 16712 1654
rect 14502 1054 14562 1110
rect 14936 1050 14996 1110
rect 15366 1054 15426 1110
rect 12220 506 12280 566
rect 19890 1950 19950 2010
rect 21176 2680 21236 2740
rect 21828 2790 21888 2850
rect 21438 2680 21498 2740
rect 20666 1950 20726 2010
rect 20920 1950 20980 2010
rect 21698 1950 21758 2010
rect 20020 1840 20080 1900
rect 20532 1840 20592 1900
rect 21052 1840 21112 1900
rect 21568 1840 21628 1900
rect 21802 1710 21862 1770
rect 16226 1054 16286 1110
rect 16656 1050 16716 1110
rect 18372 1050 18432 1110
rect 18798 1054 18858 1110
rect 22788 1840 22848 1900
rect 19656 1054 19716 1110
rect 20084 1050 20144 1110
rect 20510 1054 20570 1110
rect 18368 506 18428 566
rect 21376 1050 21436 1110
rect 21800 512 21860 572
rect 22788 512 22848 572
rect 12184 242 22840 352
rect 11972 -180 12572 120
rect 22504 -180 23104 120
rect 172 -924 772 -624
rect 10704 -924 11304 -624
rect 384 -1156 11040 -1046
rect 420 -1370 480 -1310
rect 1420 -1914 1480 -1854
rect 6568 -1370 6628 -1310
rect 2702 -1914 2762 -1858
rect 3136 -1914 3196 -1854
rect 3566 -1914 3626 -1858
rect 4426 -1914 4486 -1858
rect 4856 -1914 4916 -1854
rect 6572 -1914 6632 -1854
rect 6998 -1914 7058 -1858
rect 1418 -2458 1478 -2398
rect 420 -2704 480 -2644
rect 3306 -2582 3366 -2522
rect 1628 -2704 1688 -2644
rect 2140 -2704 2200 -2644
rect 2660 -2704 2720 -2644
rect 3176 -2704 3236 -2644
rect 1498 -2814 1558 -2754
rect 2274 -2814 2334 -2754
rect 2528 -2814 2588 -2754
rect 1758 -3544 1818 -3484
rect 1368 -3654 1428 -3594
rect 2012 -3544 2072 -3484
rect 4852 -2458 4912 -2398
rect 10000 -1376 10060 -1316
rect 10988 -1376 11048 -1316
rect 7856 -1914 7916 -1858
rect 8284 -1914 8344 -1854
rect 8710 -1914 8770 -1858
rect 5186 -2582 5246 -2522
rect 4924 -2710 4984 -2650
rect 3306 -2814 3366 -2754
rect 2784 -3544 2844 -3484
rect 2400 -3654 2460 -3594
rect 3046 -3544 3106 -3484
rect 4664 -2820 4724 -2760
rect 4794 -2820 4854 -2760
rect 3436 -3654 3496 -3594
rect 1882 -3770 1942 -3710
rect 2918 -3770 2978 -3710
rect 5436 -2710 5496 -2650
rect 5956 -2710 6016 -2650
rect 6472 -2710 6532 -2650
rect 5570 -2820 5630 -2760
rect 5696 -2822 5756 -2762
rect 5824 -2820 5884 -2760
rect 5054 -3550 5114 -3490
rect 4664 -3660 4724 -3600
rect 5308 -3550 5368 -3490
rect 9576 -1914 9636 -1854
rect 10002 -2574 10062 -2514
rect 8220 -2704 8280 -2644
rect 8732 -2704 8792 -2644
rect 9252 -2704 9312 -2644
rect 9768 -2704 9828 -2644
rect 6602 -2820 6662 -2760
rect 6080 -3550 6140 -3490
rect 5696 -3660 5756 -3600
rect 8090 -2814 8150 -2754
rect 6342 -3550 6402 -3490
rect 6732 -3660 6792 -3600
rect 5052 -3776 5112 -3716
rect 5178 -3776 5238 -3716
rect 5308 -3776 5368 -3716
rect 6080 -3776 6140 -3716
rect 6214 -3776 6274 -3716
rect 6342 -3776 6402 -3716
rect 8866 -2814 8926 -2754
rect 9120 -2814 9180 -2754
rect 8350 -3544 8410 -3484
rect 7960 -3654 8020 -3594
rect 8604 -3544 8664 -3484
rect 10988 -2704 11048 -2644
rect 9898 -2814 9958 -2754
rect 9376 -3544 9436 -3484
rect 8992 -3654 9052 -3594
rect 9638 -3544 9698 -3484
rect 10028 -3654 10088 -3594
rect 8474 -3770 8534 -3710
rect 9510 -3770 9570 -3710
rect 11972 -924 12572 -624
rect 22504 -924 23104 -624
rect 12184 -1156 22840 -1046
rect 12220 -1370 12280 -1310
rect 13220 -1914 13280 -1854
rect 18368 -1370 18428 -1310
rect 14502 -1914 14562 -1858
rect 14936 -1914 14996 -1854
rect 15366 -1914 15426 -1858
rect 16226 -1914 16286 -1858
rect 16656 -1914 16716 -1854
rect 18372 -1914 18432 -1854
rect 18798 -1914 18858 -1858
rect 13218 -2458 13278 -2398
rect 12220 -2704 12280 -2644
rect 15106 -2582 15166 -2522
rect 13428 -2704 13488 -2644
rect 13940 -2704 14000 -2644
rect 14460 -2704 14520 -2644
rect 14976 -2704 15036 -2644
rect 13298 -2814 13358 -2754
rect 14074 -2814 14134 -2754
rect 14328 -2814 14388 -2754
rect 13558 -3544 13618 -3484
rect 13168 -3654 13228 -3594
rect 13812 -3544 13872 -3484
rect 16652 -2458 16712 -2398
rect 21800 -1376 21860 -1316
rect 22788 -1376 22848 -1316
rect 19656 -1914 19716 -1858
rect 20084 -1914 20144 -1854
rect 20510 -1914 20570 -1858
rect 16986 -2582 17046 -2522
rect 16724 -2710 16784 -2650
rect 15106 -2814 15166 -2754
rect 14584 -3544 14644 -3484
rect 14200 -3654 14260 -3594
rect 14846 -3544 14906 -3484
rect 16594 -2820 16654 -2760
rect 15236 -3654 15296 -3594
rect 13682 -3770 13742 -3710
rect 14718 -3770 14778 -3710
rect 17236 -2710 17296 -2650
rect 17756 -2710 17816 -2650
rect 18272 -2710 18332 -2650
rect 17370 -2820 17430 -2760
rect 17624 -2820 17684 -2760
rect 16854 -3550 16914 -3490
rect 16464 -3660 16524 -3600
rect 16854 -3772 16914 -3712
rect 17108 -3550 17168 -3490
rect 21376 -1914 21436 -1854
rect 21802 -2574 21862 -2514
rect 20020 -2704 20080 -2644
rect 20532 -2704 20592 -2644
rect 21052 -2704 21112 -2644
rect 21568 -2704 21628 -2644
rect 18402 -2820 18462 -2760
rect 19890 -2814 19950 -2754
rect 17880 -3550 17940 -3490
rect 17496 -3660 17556 -3600
rect 18142 -3550 18202 -3490
rect 18532 -3660 18592 -3600
rect 16978 -3776 17038 -3716
rect 18014 -3776 18074 -3716
rect 20666 -2814 20726 -2754
rect 20920 -2814 20980 -2754
rect 20150 -3544 20210 -3484
rect 19760 -3654 19820 -3594
rect 20404 -3544 20464 -3484
rect 22788 -2704 22848 -2644
rect 21698 -2814 21758 -2754
rect 21176 -3544 21236 -3484
rect 20792 -3654 20852 -3594
rect 21438 -3544 21498 -3484
rect 21828 -3654 21888 -3594
rect 20274 -3770 20334 -3710
rect 21310 -3770 21370 -3710
rect 3440 -4064 3500 -4004
rect 6088 -4064 6148 -4004
rect 8476 -4064 8536 -4004
rect 15240 -4064 15300 -4004
rect 17888 -4064 17948 -4004
rect 20276 -4064 20336 -4004
rect 4668 -4382 4728 -4322
rect 4540 -4492 4600 -4432
rect 5182 -4380 5242 -4320
rect 5056 -4492 5116 -4432
rect 6088 -4378 6148 -4318
rect 5696 -5156 5756 -5096
rect 7252 -4376 7312 -4316
rect 6734 -5034 6794 -4974
rect 3902 -5450 7666 -5298
rect 172 -5836 772 -5536
rect 10704 -5836 11304 -5536
rect 16468 -4382 16528 -4322
rect 16340 -4492 16400 -4432
rect 16982 -4380 17042 -4320
rect 16856 -4492 16916 -4432
rect 17888 -4378 17948 -4318
rect 17496 -5156 17556 -5096
rect 19052 -4376 19112 -4316
rect 18534 -5034 18594 -4974
rect 15702 -5450 19466 -5298
rect 11972 -5836 12572 -5536
rect 22504 -5836 23104 -5536
<< metal2 >>
rect 172 5032 772 5042
rect 172 4722 772 4732
rect 10704 5032 11304 5042
rect 10704 4722 11304 4732
rect 11972 5032 12572 5042
rect 11972 4722 12572 4732
rect 22504 5032 23104 5042
rect 22504 4722 23104 4732
rect 3854 4646 7710 4686
rect 3854 4494 3902 4646
rect 7666 4494 7710 4646
rect 3854 4456 7710 4494
rect 15654 4646 19510 4686
rect 15654 4494 15702 4646
rect 19466 4494 19510 4646
rect 15654 4456 19510 4494
rect 5696 4352 5756 4358
rect 17496 4352 17556 4358
rect 990 4292 5696 4352
rect 990 2904 1050 4292
rect 5696 4286 5756 4292
rect 12790 4292 17496 4352
rect 6734 4230 6794 4236
rect 2920 4170 6734 4230
rect 2920 2972 2980 4170
rect 6734 4164 6794 4170
rect 4540 3688 4600 3694
rect 5056 3688 5116 3694
rect 4600 3628 5056 3688
rect 5116 3628 11180 3688
rect 4540 3622 4600 3628
rect 5056 3622 5116 3628
rect 4662 3518 4668 3578
rect 4728 3518 4734 3578
rect 3434 3200 3440 3260
rect 3500 3200 3506 3260
rect 304 2844 1050 2904
rect 1882 2966 1942 2972
rect 2918 2966 2980 2972
rect 1942 2906 2918 2966
rect 2978 2906 2980 2966
rect 1882 2900 1942 2906
rect 2918 2900 2978 2906
rect 3440 2856 3500 3200
rect 4668 2988 4728 3518
rect 5176 3516 5182 3576
rect 5242 3516 5248 3576
rect 4659 2928 4668 2988
rect 4728 2928 4737 2988
rect 5182 2978 5242 3516
rect 6082 3514 6088 3574
rect 6148 3514 6154 3574
rect 7252 3572 7312 3578
rect 6088 3260 6148 3514
rect 7312 3512 8020 3572
rect 7252 3506 7312 3512
rect 6082 3200 6088 3260
rect 6148 3200 6154 3260
rect 5178 2972 5242 2978
rect 6214 2972 6274 2978
rect 4668 2862 4728 2928
rect 5238 2912 6214 2972
rect 5178 2906 5238 2912
rect 6214 2906 6274 2912
rect 1368 2850 1428 2856
rect 2400 2850 2460 2856
rect 3436 2850 3500 2856
rect 304 1110 364 2844
rect 1428 2790 2400 2850
rect 2460 2790 3436 2850
rect 3496 2790 3500 2850
rect 4664 2856 4728 2862
rect 5696 2856 5756 2862
rect 6732 2856 6792 2862
rect 4724 2796 5696 2856
rect 5756 2796 6732 2856
rect 6792 2796 7650 2856
rect 4664 2790 4724 2796
rect 5696 2790 5756 2796
rect 6732 2790 6792 2796
rect 1368 2784 1428 2790
rect 2400 2784 2460 2790
rect 3436 2784 3496 2790
rect 5054 2746 5114 2752
rect 5308 2746 5368 2752
rect 6080 2746 6140 2752
rect 6342 2746 6402 2752
rect 1758 2740 1818 2746
rect 2012 2740 2072 2746
rect 2784 2740 2844 2746
rect 3046 2740 3106 2746
rect 1818 2680 2012 2740
rect 2072 2680 2784 2740
rect 2844 2680 3046 2740
rect 3106 2680 4104 2740
rect 4998 2686 5054 2746
rect 5114 2686 5308 2746
rect 5368 2686 6080 2746
rect 6140 2686 6342 2746
rect 5054 2680 5114 2686
rect 5308 2680 5368 2686
rect 6080 2680 6140 2686
rect 6342 2680 6402 2686
rect 7590 2740 7650 2796
rect 7960 2850 8020 3512
rect 8470 3200 8476 3260
rect 8536 3200 8542 3260
rect 8476 2972 8536 3200
rect 8474 2966 8536 2972
rect 9510 2966 9570 2972
rect 8534 2906 9510 2966
rect 8474 2900 8534 2906
rect 9510 2900 9570 2906
rect 8992 2850 9052 2856
rect 10028 2850 10088 2856
rect 8020 2790 8992 2850
rect 9052 2790 10028 2850
rect 7960 2784 8020 2790
rect 8992 2784 9052 2790
rect 10028 2784 10088 2790
rect 9642 2746 9702 2749
rect 8350 2740 8410 2746
rect 8604 2740 8664 2746
rect 9376 2740 9436 2746
rect 9638 2740 9702 2746
rect 7590 2680 8350 2740
rect 8410 2680 8604 2740
rect 8664 2680 9376 2740
rect 9436 2680 9638 2740
rect 1758 2674 1818 2680
rect 2012 2674 2072 2680
rect 2784 2674 2844 2680
rect 3046 2674 3106 2680
rect 1498 2010 1558 2016
rect 2274 2010 2334 2016
rect 2528 2010 2588 2016
rect 3306 2010 3366 2016
rect 1489 1950 1498 2010
rect 1558 1950 2274 2010
rect 2334 1950 2528 2010
rect 2588 1950 3306 2010
rect 1498 1944 1558 1950
rect 2274 1944 2334 1950
rect 2528 1944 2588 1950
rect 3306 1944 3366 1950
rect 420 1900 480 1906
rect 2140 1900 2200 1906
rect 2660 1900 2720 1906
rect 3176 1900 3236 1906
rect 480 1840 1628 1900
rect 1688 1840 2140 1900
rect 2200 1840 2660 1900
rect 2720 1840 3176 1900
rect 4044 1898 4104 2680
rect 8350 2674 8410 2680
rect 8604 2674 8664 2680
rect 9376 2674 9436 2680
rect 9638 2674 9702 2680
rect 9642 2671 9702 2674
rect 4794 2016 4854 2022
rect 5570 2016 5630 2022
rect 5824 2016 5884 2022
rect 6602 2016 6662 2022
rect 4732 1956 4794 2016
rect 4854 1956 5570 2016
rect 5630 1956 5824 2016
rect 5884 1956 6602 2016
rect 4794 1950 4854 1956
rect 5570 1950 5630 1956
rect 5824 1950 5884 1956
rect 6602 1950 6662 1956
rect 8090 2010 8150 2016
rect 8866 2010 8926 2016
rect 9120 2010 9180 2016
rect 9898 2010 9958 2016
rect 8150 1950 8866 2010
rect 8926 1950 9120 2010
rect 9180 1950 9898 2010
rect 8090 1944 8152 1950
rect 8866 1944 8926 1950
rect 9120 1944 9180 1950
rect 9898 1944 9958 1950
rect 5436 1906 5496 1912
rect 5956 1906 6016 1912
rect 6472 1906 6532 1912
rect 420 1834 480 1840
rect 2140 1834 2200 1840
rect 2660 1834 2720 1840
rect 3176 1834 3236 1840
rect 4035 1838 4044 1898
rect 4104 1838 4113 1898
rect 4918 1846 4924 1906
rect 4984 1846 5436 1906
rect 5496 1846 5956 1906
rect 6016 1846 6472 1906
rect 8092 1896 8152 1944
rect 8220 1900 8280 1906
rect 8732 1900 8792 1906
rect 9252 1900 9312 1906
rect 9768 1900 9828 1906
rect 10988 1900 11048 1906
rect 5436 1840 5496 1846
rect 5956 1840 6016 1846
rect 6472 1840 6532 1846
rect 8085 1840 8094 1896
rect 8150 1840 8159 1896
rect 8280 1840 8732 1900
rect 8792 1840 9252 1900
rect 9312 1840 9768 1900
rect 9828 1840 10988 1900
rect 8092 1838 8152 1840
rect 8220 1834 8280 1840
rect 8732 1834 8792 1840
rect 9252 1834 9312 1840
rect 9768 1834 9828 1840
rect 10988 1834 11048 1840
rect 3306 1778 3366 1784
rect 5186 1778 5246 1784
rect 3366 1718 5186 1778
rect 3306 1712 3366 1718
rect 5186 1712 5246 1718
rect 10002 1770 10062 1776
rect 11120 1770 11180 3628
rect 12790 2904 12850 4292
rect 17496 4286 17556 4292
rect 18534 4230 18594 4236
rect 14720 4170 18534 4230
rect 14720 2972 14780 4170
rect 18534 4164 18594 4170
rect 16340 3688 16400 3694
rect 16856 3688 16916 3694
rect 16400 3628 16856 3688
rect 16916 3628 22980 3688
rect 16340 3622 16400 3628
rect 16856 3622 16916 3628
rect 16462 3518 16468 3578
rect 16528 3518 16534 3578
rect 15234 3200 15240 3260
rect 15300 3200 15306 3260
rect 11488 2871 11588 2876
rect 11484 2781 11493 2871
rect 11583 2781 11592 2871
rect 12104 2844 12850 2904
rect 13682 2966 13742 2972
rect 14718 2966 14780 2972
rect 13742 2906 14718 2966
rect 14778 2906 14780 2966
rect 13682 2900 13742 2906
rect 14718 2900 14778 2906
rect 15240 2856 15300 3200
rect 16468 2862 16528 3518
rect 16976 3516 16982 3576
rect 17042 3516 17048 3576
rect 16982 3264 17042 3516
rect 17882 3514 17888 3574
rect 17948 3514 17954 3574
rect 19052 3572 19112 3578
rect 16973 3204 16982 3264
rect 17042 3204 17051 3264
rect 17888 3260 17948 3514
rect 19112 3512 19820 3572
rect 19052 3506 19112 3512
rect 16982 2978 17042 3204
rect 17882 3200 17888 3260
rect 17948 3200 17954 3260
rect 16978 2972 17042 2978
rect 18014 2972 18074 2978
rect 17038 2912 18014 2972
rect 16978 2906 17038 2912
rect 18014 2906 18074 2912
rect 16464 2856 16528 2862
rect 17496 2856 17556 2862
rect 18532 2856 18592 2862
rect 13168 2850 13228 2856
rect 14200 2850 14260 2856
rect 15236 2850 15300 2856
rect 10062 1710 11180 1770
rect 10002 1704 10062 1710
rect 1418 1654 1478 1660
rect 4852 1654 4912 1660
rect 1478 1594 4852 1654
rect 1418 1588 1478 1594
rect 4852 1588 4912 1594
rect 1420 1110 1480 1116
rect 304 1050 1420 1110
rect 1420 1044 1480 1050
rect 2702 1110 2762 1116
rect 3136 1110 3196 1116
rect 4856 1110 4916 1116
rect 6572 1110 6632 1116
rect 6998 1110 7058 1116
rect 8284 1110 8344 1116
rect 2762 1054 3136 1110
rect 2702 1050 3136 1054
rect 3196 1054 3566 1110
rect 3626 1054 4426 1110
rect 4486 1054 4856 1110
rect 3196 1050 4856 1054
rect 4916 1050 6572 1110
rect 6632 1054 6998 1110
rect 7058 1054 7856 1110
rect 7916 1054 8284 1110
rect 6632 1050 8284 1054
rect 8344 1054 8710 1110
rect 8770 1054 9576 1110
rect 8344 1050 9576 1054
rect 9636 1050 9642 1110
rect 2702 1044 2762 1050
rect 3136 1044 3196 1050
rect 4856 1044 4916 1050
rect 6572 1044 6632 1050
rect 6998 1044 7058 1050
rect 8284 1044 8344 1050
rect 10000 572 10060 578
rect 10988 572 11048 578
rect 420 566 480 572
rect 6568 566 6628 572
rect 480 506 6568 566
rect 10060 512 10988 572
rect 10000 506 10060 512
rect 10988 506 11048 512
rect 420 500 480 506
rect 6568 500 6628 506
rect 322 352 11096 400
rect 322 242 384 352
rect 11040 242 11096 352
rect 322 186 11096 242
rect 172 120 772 130
rect 172 -190 772 -180
rect 10704 120 11304 130
rect 10704 -190 11304 -180
rect 172 -624 772 -614
rect 172 -934 772 -924
rect 10704 -624 11304 -614
rect 10704 -934 11304 -924
rect 322 -1046 11096 -990
rect 322 -1156 384 -1046
rect 11040 -1156 11096 -1046
rect 322 -1204 11096 -1156
rect 420 -1310 480 -1304
rect 6568 -1310 6628 -1304
rect 480 -1370 6568 -1310
rect 420 -1376 480 -1370
rect 6568 -1376 6628 -1370
rect 10000 -1316 10060 -1310
rect 10988 -1316 11048 -1310
rect 10060 -1376 10988 -1316
rect 10000 -1382 10060 -1376
rect 10988 -1382 11048 -1376
rect 1420 -1854 1480 -1848
rect 304 -1914 1420 -1854
rect 304 -3648 364 -1914
rect 1420 -1920 1480 -1914
rect 2702 -1854 2762 -1848
rect 3136 -1854 3196 -1848
rect 4856 -1854 4916 -1848
rect 6572 -1854 6632 -1848
rect 6998 -1854 7058 -1848
rect 8284 -1854 8344 -1848
rect 2702 -1858 3136 -1854
rect 2762 -1914 3136 -1858
rect 3196 -1858 4856 -1854
rect 3196 -1914 3566 -1858
rect 3626 -1914 4426 -1858
rect 4486 -1914 4856 -1858
rect 4916 -1914 6572 -1854
rect 6632 -1858 8284 -1854
rect 6632 -1914 6998 -1858
rect 7058 -1914 7856 -1858
rect 7916 -1914 8284 -1858
rect 8344 -1858 9576 -1854
rect 8344 -1914 8710 -1858
rect 8770 -1914 9576 -1858
rect 9636 -1914 9642 -1854
rect 2702 -1920 2762 -1914
rect 3136 -1920 3196 -1914
rect 4856 -1920 4916 -1914
rect 6572 -1920 6632 -1914
rect 6998 -1920 7058 -1914
rect 8284 -1920 8344 -1914
rect 1418 -2398 1478 -2392
rect 4852 -2398 4912 -2392
rect 1478 -2458 4852 -2398
rect 1418 -2464 1478 -2458
rect 4852 -2464 4912 -2458
rect 10002 -2514 10062 -2508
rect 3306 -2522 3366 -2516
rect 5186 -2522 5246 -2516
rect 3366 -2582 5186 -2522
rect 10062 -2574 11180 -2514
rect 10002 -2580 10062 -2574
rect 3306 -2588 3366 -2582
rect 5186 -2588 5246 -2582
rect 420 -2644 480 -2638
rect 2140 -2644 2200 -2638
rect 2660 -2644 2720 -2638
rect 3176 -2644 3236 -2638
rect 480 -2704 1628 -2644
rect 1688 -2704 2140 -2644
rect 2200 -2704 2660 -2644
rect 2720 -2704 3176 -2644
rect 4035 -2702 4044 -2642
rect 4104 -2702 4113 -2642
rect 8092 -2644 8152 -2642
rect 8220 -2644 8280 -2638
rect 8732 -2644 8792 -2638
rect 9252 -2644 9312 -2638
rect 9768 -2644 9828 -2638
rect 10988 -2644 11048 -2638
rect 5436 -2650 5496 -2644
rect 5956 -2650 6016 -2644
rect 6472 -2650 6532 -2644
rect 420 -2710 480 -2704
rect 2140 -2710 2200 -2704
rect 2660 -2710 2720 -2704
rect 3176 -2710 3236 -2704
rect 1498 -2754 1558 -2748
rect 2274 -2754 2334 -2748
rect 2528 -2754 2588 -2748
rect 3306 -2754 3366 -2748
rect 1558 -2814 2274 -2754
rect 2334 -2814 2528 -2754
rect 2588 -2814 3306 -2754
rect 1498 -2820 1558 -2814
rect 2274 -2820 2334 -2814
rect 2528 -2820 2588 -2814
rect 3306 -2820 3366 -2814
rect 1758 -3484 1818 -3478
rect 2012 -3484 2072 -3478
rect 2784 -3484 2844 -3478
rect 3046 -3484 3106 -3478
rect 4044 -3484 4104 -2702
rect 4918 -2710 4924 -2650
rect 4984 -2710 5436 -2650
rect 5496 -2710 5956 -2650
rect 6016 -2710 6472 -2650
rect 8085 -2700 8094 -2644
rect 8150 -2700 8159 -2644
rect 5436 -2716 5496 -2710
rect 5956 -2716 6016 -2710
rect 6472 -2716 6532 -2710
rect 8092 -2748 8152 -2700
rect 8280 -2704 8732 -2644
rect 8792 -2704 9252 -2644
rect 9312 -2704 9768 -2644
rect 9828 -2704 10988 -2644
rect 8220 -2710 8280 -2704
rect 8732 -2710 8792 -2704
rect 9252 -2710 9312 -2704
rect 9768 -2710 9828 -2704
rect 10988 -2710 11048 -2704
rect 8090 -2754 8152 -2748
rect 8866 -2754 8926 -2748
rect 9120 -2754 9180 -2748
rect 9898 -2754 9958 -2748
rect 4794 -2760 4854 -2754
rect 5570 -2760 5630 -2754
rect 5696 -2760 5756 -2756
rect 5824 -2760 5884 -2754
rect 6602 -2760 6662 -2754
rect 4268 -2820 4664 -2760
rect 4724 -2820 4794 -2760
rect 4854 -2820 5570 -2760
rect 5630 -2762 5824 -2760
rect 5630 -2820 5696 -2762
rect 4268 -2916 4328 -2820
rect 4794 -2826 4854 -2820
rect 5570 -2826 5630 -2820
rect 5756 -2820 5824 -2762
rect 5884 -2820 6602 -2760
rect 8150 -2814 8866 -2754
rect 8926 -2814 9120 -2754
rect 9180 -2814 9898 -2754
rect 8090 -2820 8150 -2814
rect 8866 -2820 8926 -2814
rect 9120 -2820 9180 -2814
rect 9898 -2820 9958 -2814
rect 5696 -2828 5756 -2822
rect 5824 -2826 5884 -2820
rect 6602 -2826 6662 -2820
rect 4259 -2976 4268 -2916
rect 4328 -2976 4337 -2916
rect 8350 -3484 8410 -3478
rect 8604 -3484 8664 -3478
rect 9376 -3484 9436 -3478
rect 9638 -3484 9698 -3478
rect 1818 -3544 2012 -3484
rect 2072 -3544 2784 -3484
rect 2844 -3544 3046 -3484
rect 3106 -3544 4104 -3484
rect 5054 -3490 5114 -3484
rect 5308 -3490 5368 -3484
rect 6080 -3490 6140 -3484
rect 6342 -3490 6402 -3484
rect 1758 -3550 1818 -3544
rect 2012 -3550 2072 -3544
rect 2784 -3550 2844 -3544
rect 3046 -3550 3106 -3544
rect 5045 -3550 5054 -3490
rect 5114 -3550 5308 -3490
rect 5368 -3550 6080 -3490
rect 6140 -3550 6342 -3490
rect 5054 -3556 5114 -3550
rect 5308 -3556 5368 -3550
rect 6080 -3556 6140 -3550
rect 6342 -3556 6402 -3550
rect 7590 -3544 8350 -3484
rect 8410 -3544 8604 -3484
rect 8664 -3544 9376 -3484
rect 9436 -3544 9638 -3484
rect 9698 -3544 9707 -3484
rect 1368 -3594 1428 -3588
rect 2400 -3594 2460 -3588
rect 3436 -3594 3496 -3588
rect 304 -3708 1050 -3648
rect 1428 -3654 2400 -3594
rect 2460 -3654 3436 -3594
rect 3496 -3654 3500 -3594
rect 1368 -3660 1428 -3654
rect 2400 -3660 2460 -3654
rect 3436 -3660 3500 -3654
rect 990 -5096 1050 -3708
rect 1882 -3710 1942 -3704
rect 2918 -3710 2978 -3704
rect 1942 -3770 2918 -3710
rect 2978 -3770 2980 -3710
rect 1882 -3776 1942 -3770
rect 2918 -3776 2980 -3770
rect 2920 -4974 2980 -3776
rect 3440 -4004 3500 -3660
rect 4664 -3600 4724 -3594
rect 5696 -3600 5756 -3594
rect 6732 -3600 6792 -3594
rect 7590 -3600 7650 -3544
rect 8350 -3550 8410 -3544
rect 8604 -3550 8664 -3544
rect 9376 -3550 9436 -3544
rect 9638 -3550 9698 -3544
rect 4724 -3660 5696 -3600
rect 5756 -3660 6732 -3600
rect 6792 -3660 7650 -3600
rect 7960 -3594 8020 -3588
rect 8992 -3594 9052 -3588
rect 10028 -3594 10088 -3588
rect 8020 -3654 8992 -3594
rect 9052 -3654 10028 -3594
rect 4664 -3666 4728 -3660
rect 5696 -3666 5756 -3660
rect 6732 -3666 6792 -3660
rect 3434 -4064 3440 -4004
rect 3500 -4064 3506 -4004
rect 4668 -4322 4728 -3666
rect 5052 -3716 5112 -3710
rect 5178 -3716 5238 -3710
rect 5308 -3716 5368 -3710
rect 6080 -3716 6140 -3710
rect 6214 -3716 6274 -3710
rect 6342 -3716 6402 -3710
rect 5112 -3776 5178 -3716
rect 5238 -3776 5308 -3716
rect 5368 -3776 6080 -3716
rect 6140 -3776 6214 -3716
rect 6274 -3776 6342 -3716
rect 6402 -3776 6411 -3716
rect 5052 -3782 5112 -3776
rect 5178 -3782 5242 -3776
rect 5308 -3782 5368 -3776
rect 6080 -3782 6140 -3776
rect 6214 -3782 6274 -3776
rect 6342 -3782 6402 -3776
rect 5182 -4320 5242 -3782
rect 6082 -4064 6088 -4004
rect 6148 -4064 6154 -4004
rect 6088 -4318 6148 -4064
rect 7252 -4316 7312 -4310
rect 7960 -4316 8020 -3654
rect 8992 -3660 9052 -3654
rect 10028 -3660 10088 -3654
rect 8474 -3710 8534 -3704
rect 9510 -3710 9570 -3704
rect 8534 -3770 9510 -3710
rect 8474 -3776 8536 -3770
rect 9510 -3776 9570 -3770
rect 8476 -4004 8536 -3776
rect 8470 -4064 8476 -4004
rect 8536 -4064 8542 -4004
rect 4662 -4382 4668 -4322
rect 4728 -4382 4734 -4322
rect 5176 -4380 5182 -4320
rect 5242 -4380 5248 -4320
rect 6082 -4378 6088 -4318
rect 6148 -4378 6154 -4318
rect 7312 -4376 8020 -4316
rect 7252 -4382 7312 -4376
rect 4540 -4432 4600 -4426
rect 5056 -4432 5116 -4426
rect 11120 -4432 11180 -2574
rect 11488 -3464 11588 2781
rect 11691 1816 11700 1916
rect 11800 1816 11809 1916
rect 11700 -2625 11800 1816
rect 12104 1110 12164 2844
rect 13228 2790 14200 2850
rect 14260 2790 15236 2850
rect 15296 2790 15300 2850
rect 16459 2796 16464 2856
rect 16528 2796 17496 2856
rect 17556 2796 18532 2856
rect 18592 2796 19450 2856
rect 16464 2790 16524 2796
rect 17496 2790 17556 2796
rect 18532 2790 18592 2796
rect 13168 2784 13228 2790
rect 14200 2784 14260 2790
rect 15236 2784 15296 2790
rect 16854 2746 16914 2752
rect 17108 2746 17168 2752
rect 17880 2746 17940 2752
rect 18142 2746 18202 2752
rect 13558 2740 13618 2746
rect 13812 2740 13872 2746
rect 14584 2740 14644 2746
rect 14846 2740 14906 2746
rect 13618 2680 13812 2740
rect 13872 2680 14584 2740
rect 14644 2680 14846 2740
rect 14906 2680 15904 2740
rect 16914 2686 17108 2746
rect 17168 2686 17880 2746
rect 17940 2686 18142 2746
rect 18204 2686 18213 2746
rect 19390 2740 19450 2796
rect 19760 2850 19820 3512
rect 20270 3200 20276 3260
rect 20336 3200 20342 3260
rect 20276 2972 20336 3200
rect 20274 2966 20336 2972
rect 21310 2966 21370 2972
rect 20334 2906 21310 2966
rect 20274 2900 20334 2906
rect 21310 2900 21370 2906
rect 20792 2850 20852 2856
rect 21828 2850 21888 2856
rect 19820 2790 20792 2850
rect 20852 2790 21828 2850
rect 19760 2784 19820 2790
rect 20792 2784 20852 2790
rect 21828 2784 21888 2790
rect 20150 2740 20210 2746
rect 20404 2740 20464 2746
rect 21176 2740 21236 2746
rect 21438 2740 21498 2746
rect 16854 2680 16914 2686
rect 17108 2680 17168 2686
rect 17880 2680 17940 2686
rect 18142 2680 18202 2686
rect 19390 2680 20150 2740
rect 20210 2680 20404 2740
rect 20464 2680 21176 2740
rect 21236 2680 21438 2740
rect 13558 2674 13618 2680
rect 13812 2674 13872 2680
rect 14584 2674 14644 2680
rect 14846 2674 14906 2680
rect 13298 2010 13358 2016
rect 14074 2010 14134 2016
rect 14328 2010 14388 2016
rect 15106 2010 15166 2016
rect 13358 1950 14074 2010
rect 14134 1950 14328 2010
rect 14388 1950 15106 2010
rect 13298 1944 13358 1950
rect 14074 1944 14134 1950
rect 14328 1944 14388 1950
rect 15106 1944 15166 1950
rect 12220 1900 12280 1906
rect 13940 1900 14000 1906
rect 14460 1900 14520 1906
rect 14976 1900 15036 1906
rect 12280 1840 13428 1900
rect 13488 1840 13940 1900
rect 14000 1840 14460 1900
rect 14520 1840 14976 1900
rect 15844 1898 15904 2680
rect 20150 2674 20210 2680
rect 20404 2674 20464 2680
rect 21176 2674 21236 2680
rect 21438 2674 21498 2680
rect 16594 2016 16654 2022
rect 17370 2016 17430 2022
rect 17624 2016 17684 2022
rect 18402 2016 18462 2022
rect 16654 1956 17370 2016
rect 17430 1956 17624 2016
rect 17684 1956 18402 2016
rect 18462 1956 18980 2016
rect 16594 1950 16654 1956
rect 17370 1950 17430 1956
rect 17624 1950 17684 1956
rect 18402 1950 18462 1956
rect 17236 1906 17296 1912
rect 17756 1906 17816 1912
rect 18272 1906 18332 1912
rect 12220 1834 12280 1840
rect 13940 1834 14000 1840
rect 14460 1834 14520 1840
rect 14976 1834 15036 1840
rect 15835 1838 15844 1898
rect 15904 1838 15913 1898
rect 16718 1846 16724 1906
rect 16784 1846 17236 1906
rect 17296 1846 17756 1906
rect 17816 1846 18272 1906
rect 17236 1840 17296 1846
rect 17756 1840 17816 1846
rect 18272 1840 18332 1846
rect 15106 1778 15166 1784
rect 16986 1778 17046 1784
rect 15166 1718 16986 1778
rect 15106 1712 15166 1718
rect 16986 1712 17046 1718
rect 18920 1684 18980 1956
rect 19890 2010 19950 2016
rect 20666 2010 20726 2016
rect 20920 2010 20980 2016
rect 21698 2010 21758 2016
rect 19950 1950 20666 2010
rect 20726 1950 20920 2010
rect 20980 1950 21698 2010
rect 19890 1944 19952 1950
rect 20666 1944 20726 1950
rect 20920 1944 20980 1950
rect 21698 1944 21758 1950
rect 19892 1896 19952 1944
rect 20020 1900 20080 1906
rect 20532 1900 20592 1906
rect 21052 1900 21112 1906
rect 21568 1900 21628 1906
rect 22788 1900 22848 1906
rect 19885 1840 19894 1896
rect 19950 1840 19959 1896
rect 20080 1840 20532 1900
rect 20592 1840 21052 1900
rect 21112 1840 21568 1900
rect 21628 1840 22788 1900
rect 19892 1838 19952 1840
rect 20020 1834 20080 1840
rect 20532 1834 20592 1840
rect 21052 1834 21112 1840
rect 21568 1834 21628 1840
rect 22788 1834 22848 1840
rect 21802 1770 21862 1776
rect 22920 1770 22980 3628
rect 21862 1710 22980 1770
rect 21802 1704 21862 1710
rect 13218 1654 13278 1660
rect 16652 1654 16712 1660
rect 13278 1594 16652 1654
rect 18911 1624 18920 1684
rect 18980 1624 18989 1684
rect 13218 1588 13278 1594
rect 16652 1588 16712 1594
rect 13220 1110 13280 1116
rect 12104 1050 13220 1110
rect 13220 1044 13280 1050
rect 14502 1110 14562 1116
rect 14936 1110 14996 1116
rect 16656 1110 16716 1116
rect 18372 1110 18432 1116
rect 18798 1110 18858 1116
rect 20084 1110 20144 1116
rect 14562 1054 14936 1110
rect 14502 1050 14936 1054
rect 14996 1054 15366 1110
rect 15426 1054 16226 1110
rect 16286 1054 16656 1110
rect 14996 1050 16656 1054
rect 16716 1050 18372 1110
rect 18432 1054 18798 1110
rect 18858 1054 19656 1110
rect 19716 1054 20084 1110
rect 18432 1050 20084 1054
rect 20144 1054 20510 1110
rect 20570 1054 21376 1110
rect 20144 1050 21376 1054
rect 21436 1050 21442 1110
rect 14502 1044 14562 1050
rect 14936 1044 14996 1050
rect 16656 1044 16716 1050
rect 18372 1044 18432 1050
rect 18798 1044 18858 1050
rect 20084 1044 20144 1050
rect 21800 572 21860 578
rect 22788 572 22848 578
rect 12220 566 12280 572
rect 18368 566 18428 572
rect 12280 506 18368 566
rect 21860 512 22788 572
rect 21800 506 21860 512
rect 22788 506 22848 512
rect 12220 500 12280 506
rect 18368 500 18428 506
rect 12122 352 22896 400
rect 12122 242 12184 352
rect 22840 242 22896 352
rect 12122 186 22896 242
rect 11972 120 12572 130
rect 11972 -190 12572 -180
rect 22504 120 23104 130
rect 22504 -190 23104 -180
rect 11972 -624 12572 -614
rect 11972 -934 12572 -924
rect 22504 -624 23104 -614
rect 22504 -934 23104 -924
rect 12122 -1046 22896 -990
rect 12122 -1156 12184 -1046
rect 22840 -1156 22896 -1046
rect 12122 -1204 22896 -1156
rect 12220 -1310 12280 -1304
rect 18368 -1310 18428 -1304
rect 12280 -1370 18368 -1310
rect 12220 -1376 12280 -1370
rect 18368 -1376 18428 -1370
rect 21800 -1316 21860 -1310
rect 22788 -1316 22848 -1310
rect 21860 -1376 22788 -1316
rect 21800 -1382 21860 -1376
rect 22788 -1382 22848 -1376
rect 13220 -1854 13280 -1848
rect 12104 -1914 13220 -1854
rect 11696 -2715 11705 -2625
rect 11795 -2715 11804 -2625
rect 11700 -2720 11800 -2715
rect 11479 -3564 11488 -3464
rect 11588 -3564 11597 -3464
rect 12104 -3648 12164 -1914
rect 13220 -1920 13280 -1914
rect 14502 -1854 14562 -1848
rect 14936 -1854 14996 -1848
rect 16656 -1854 16716 -1848
rect 18372 -1854 18432 -1848
rect 18798 -1854 18858 -1848
rect 20084 -1854 20144 -1848
rect 14502 -1858 14936 -1854
rect 14562 -1914 14936 -1858
rect 14996 -1858 16656 -1854
rect 14996 -1914 15366 -1858
rect 15426 -1914 16226 -1858
rect 16286 -1914 16656 -1858
rect 16716 -1914 18372 -1854
rect 18432 -1858 20084 -1854
rect 18432 -1914 18798 -1858
rect 18858 -1914 19656 -1858
rect 19716 -1914 20084 -1858
rect 20144 -1858 21376 -1854
rect 20144 -1914 20510 -1858
rect 20570 -1914 21376 -1858
rect 21436 -1914 21442 -1854
rect 14502 -1920 14562 -1914
rect 14936 -1920 14996 -1914
rect 16656 -1920 16716 -1914
rect 18372 -1920 18432 -1914
rect 18798 -1920 18858 -1914
rect 20084 -1920 20144 -1914
rect 13218 -2398 13278 -2392
rect 16652 -2398 16712 -2392
rect 13278 -2458 16652 -2398
rect 13218 -2464 13278 -2458
rect 16652 -2464 16712 -2458
rect 16979 -2462 16988 -2402
rect 17048 -2462 17057 -2402
rect 16988 -2516 17048 -2462
rect 15106 -2522 15166 -2516
rect 16986 -2522 17048 -2516
rect 15166 -2582 16986 -2522
rect 17046 -2582 17048 -2522
rect 21802 -2514 21862 -2508
rect 21862 -2574 22980 -2514
rect 21802 -2580 21862 -2574
rect 15106 -2588 15166 -2582
rect 16986 -2588 17046 -2582
rect 12220 -2644 12280 -2638
rect 13940 -2644 14000 -2638
rect 14460 -2644 14520 -2638
rect 14976 -2644 15036 -2638
rect 12280 -2704 13428 -2644
rect 13488 -2704 13940 -2644
rect 14000 -2704 14460 -2644
rect 14520 -2704 14976 -2644
rect 15835 -2702 15844 -2642
rect 15904 -2702 15913 -2642
rect 19892 -2644 19952 -2642
rect 20020 -2644 20080 -2638
rect 20532 -2644 20592 -2638
rect 21052 -2644 21112 -2638
rect 21568 -2644 21628 -2638
rect 22788 -2644 22848 -2638
rect 17236 -2650 17296 -2644
rect 17756 -2650 17816 -2644
rect 18272 -2650 18332 -2644
rect 12220 -2710 12280 -2704
rect 13940 -2710 14000 -2704
rect 14460 -2710 14520 -2704
rect 14976 -2710 15036 -2704
rect 13298 -2754 13358 -2748
rect 14074 -2754 14134 -2748
rect 14328 -2754 14388 -2748
rect 15106 -2754 15166 -2748
rect 13358 -2814 14074 -2754
rect 14134 -2814 14328 -2754
rect 14388 -2814 15106 -2754
rect 13298 -2820 13358 -2814
rect 14074 -2820 14134 -2814
rect 14328 -2820 14388 -2814
rect 15106 -2820 15166 -2814
rect 13558 -3484 13618 -3478
rect 13812 -3484 13872 -3478
rect 14584 -3484 14644 -3478
rect 14846 -3484 14906 -3478
rect 15844 -3484 15904 -2702
rect 16718 -2710 16724 -2650
rect 16784 -2710 17236 -2650
rect 17296 -2710 17756 -2650
rect 17816 -2710 18272 -2650
rect 19885 -2700 19894 -2644
rect 19950 -2700 19959 -2644
rect 17236 -2716 17296 -2710
rect 17756 -2716 17816 -2710
rect 18272 -2716 18332 -2710
rect 19892 -2748 19952 -2700
rect 20080 -2704 20532 -2644
rect 20592 -2704 21052 -2644
rect 21112 -2704 21568 -2644
rect 21628 -2704 22788 -2644
rect 20020 -2710 20080 -2704
rect 20532 -2710 20592 -2704
rect 21052 -2710 21112 -2704
rect 21568 -2710 21628 -2704
rect 22788 -2710 22848 -2704
rect 19890 -2754 19952 -2748
rect 20666 -2754 20726 -2748
rect 20920 -2754 20980 -2748
rect 21698 -2754 21758 -2748
rect 16594 -2760 16654 -2754
rect 17370 -2760 17430 -2754
rect 17624 -2760 17684 -2754
rect 18402 -2760 18462 -2754
rect 16070 -2820 16594 -2760
rect 16654 -2820 17370 -2760
rect 17430 -2820 17624 -2760
rect 17684 -2820 18402 -2760
rect 19950 -2814 20666 -2754
rect 20726 -2814 20920 -2754
rect 20980 -2814 21698 -2754
rect 19890 -2820 19950 -2814
rect 20666 -2820 20726 -2814
rect 20920 -2820 20980 -2814
rect 21698 -2820 21758 -2814
rect 16070 -3480 16130 -2820
rect 16594 -2826 16654 -2820
rect 17370 -2826 17430 -2820
rect 17624 -2826 17684 -2820
rect 18402 -2826 18462 -2820
rect 13618 -3544 13812 -3484
rect 13872 -3544 14584 -3484
rect 14644 -3544 14846 -3484
rect 14906 -3544 15904 -3484
rect 16061 -3540 16070 -3480
rect 16130 -3540 16139 -3480
rect 20150 -3484 20210 -3478
rect 20404 -3484 20464 -3478
rect 21176 -3484 21236 -3478
rect 21438 -3484 21498 -3478
rect 16854 -3490 16914 -3484
rect 17108 -3490 17168 -3484
rect 17880 -3490 17940 -3484
rect 18142 -3490 18202 -3484
rect 13558 -3550 13618 -3544
rect 13812 -3550 13872 -3544
rect 14584 -3550 14644 -3544
rect 14846 -3550 14906 -3544
rect 16914 -3550 17108 -3490
rect 17168 -3550 17880 -3490
rect 17940 -3550 18142 -3490
rect 16854 -3556 16914 -3550
rect 17108 -3556 17168 -3550
rect 17880 -3556 17940 -3550
rect 18142 -3556 18202 -3550
rect 19390 -3544 20150 -3484
rect 20210 -3544 20404 -3484
rect 20464 -3544 21176 -3484
rect 21236 -3544 21438 -3484
rect 21500 -3544 21509 -3484
rect 13168 -3594 13228 -3588
rect 14200 -3594 14260 -3588
rect 15236 -3594 15296 -3588
rect 12104 -3708 12850 -3648
rect 13228 -3654 14200 -3594
rect 14260 -3654 15236 -3594
rect 15296 -3654 15300 -3594
rect 13168 -3660 13228 -3654
rect 14200 -3660 14260 -3654
rect 15236 -3660 15300 -3654
rect 4600 -4492 5056 -4432
rect 5116 -4492 11180 -4432
rect 4540 -4498 4600 -4492
rect 5056 -4498 5116 -4492
rect 6734 -4974 6794 -4968
rect 2920 -5034 6734 -4974
rect 6734 -5040 6794 -5034
rect 5696 -5096 5756 -5090
rect 990 -5156 5696 -5096
rect 12790 -5096 12850 -3708
rect 13682 -3710 13742 -3704
rect 14718 -3710 14778 -3704
rect 13742 -3770 14718 -3710
rect 14778 -3770 14780 -3710
rect 13682 -3776 13742 -3770
rect 14718 -3776 14780 -3770
rect 14720 -4974 14780 -3776
rect 15240 -4004 15300 -3660
rect 16464 -3600 16524 -3594
rect 17496 -3600 17556 -3594
rect 18532 -3600 18592 -3594
rect 19390 -3600 19450 -3544
rect 20150 -3550 20210 -3544
rect 20404 -3550 20464 -3544
rect 21176 -3550 21236 -3544
rect 21438 -3550 21498 -3544
rect 16524 -3660 17496 -3600
rect 17556 -3660 18532 -3600
rect 18592 -3660 19450 -3600
rect 19760 -3594 19820 -3588
rect 20792 -3594 20852 -3588
rect 21828 -3594 21888 -3588
rect 19820 -3654 20792 -3594
rect 20852 -3654 21828 -3594
rect 16464 -3666 16528 -3660
rect 17496 -3666 17556 -3660
rect 18532 -3666 18592 -3660
rect 15234 -4064 15240 -4004
rect 15300 -4064 15306 -4004
rect 16468 -4322 16528 -3666
rect 16854 -3712 16914 -3706
rect 16845 -3772 16854 -3712
rect 16914 -3772 16923 -3712
rect 16978 -3716 17038 -3710
rect 18014 -3716 18074 -3710
rect 16854 -3778 16914 -3772
rect 17038 -3776 18014 -3716
rect 16978 -3782 17042 -3776
rect 18014 -3782 18074 -3776
rect 16982 -4320 17042 -3782
rect 17882 -4064 17888 -4004
rect 17948 -4064 17954 -4004
rect 17888 -4318 17948 -4064
rect 19052 -4316 19112 -4310
rect 19760 -4316 19820 -3654
rect 20792 -3660 20852 -3654
rect 21828 -3660 21888 -3654
rect 20274 -3710 20334 -3704
rect 21310 -3710 21370 -3704
rect 20334 -3770 21310 -3710
rect 20274 -3776 20336 -3770
rect 21310 -3776 21370 -3770
rect 20276 -4004 20336 -3776
rect 20270 -4064 20276 -4004
rect 20336 -4064 20342 -4004
rect 16462 -4382 16468 -4322
rect 16528 -4382 16534 -4322
rect 16976 -4380 16982 -4320
rect 17042 -4380 17048 -4320
rect 17882 -4378 17888 -4318
rect 17948 -4378 17954 -4318
rect 19112 -4376 19820 -4316
rect 19052 -4382 19112 -4376
rect 16340 -4432 16400 -4426
rect 16856 -4432 16916 -4426
rect 22920 -4432 22980 -2574
rect 16400 -4492 16856 -4432
rect 16916 -4492 22980 -4432
rect 16340 -4498 16400 -4492
rect 16856 -4498 16916 -4492
rect 18534 -4974 18594 -4968
rect 14720 -5034 18534 -4974
rect 18534 -5040 18594 -5034
rect 17496 -5096 17556 -5090
rect 12790 -5156 17496 -5096
rect 5696 -5162 5756 -5156
rect 17496 -5162 17556 -5156
rect 3854 -5298 7710 -5260
rect 3854 -5450 3902 -5298
rect 7666 -5450 7710 -5298
rect 3854 -5490 7710 -5450
rect 15654 -5298 19510 -5260
rect 15654 -5450 15702 -5298
rect 19466 -5450 19510 -5298
rect 15654 -5490 19510 -5450
rect 172 -5536 772 -5526
rect 172 -5846 772 -5836
rect 10704 -5536 11304 -5526
rect 10704 -5846 11304 -5836
rect 11972 -5536 12572 -5526
rect 11972 -5846 12572 -5836
rect 22504 -5536 23104 -5526
rect 22504 -5846 23104 -5836
<< via2 >>
rect 172 4732 772 5032
rect 10704 4732 11304 5032
rect 11972 4732 12572 5032
rect 22504 4732 23104 5032
rect 3902 4494 7666 4646
rect 15702 4494 19466 4646
rect 4668 2928 4728 2988
rect 9642 2680 9698 2740
rect 9698 2680 9702 2740
rect 1498 1950 1558 2010
rect 4044 1838 4104 1898
rect 8094 1840 8150 1896
rect 11493 2781 11583 2871
rect 16982 3204 17042 3264
rect 384 242 11040 352
rect 172 -180 772 120
rect 10704 -180 11304 120
rect 172 -924 772 -624
rect 10704 -924 11304 -624
rect 384 -1156 11040 -1046
rect 4044 -2702 4104 -2642
rect 8094 -2700 8150 -2644
rect 4268 -2976 4328 -2916
rect 5054 -3550 5114 -3490
rect 9638 -3544 9698 -3484
rect 6342 -3776 6402 -3716
rect 11700 1816 11800 1916
rect 16468 2796 16524 2856
rect 16524 2796 16528 2856
rect 18144 2686 18202 2746
rect 18202 2686 18204 2746
rect 15844 1838 15904 1898
rect 19894 1840 19950 1896
rect 18920 1624 18980 1684
rect 12184 242 22840 352
rect 11972 -180 12572 120
rect 22504 -180 23104 120
rect 11972 -924 12572 -624
rect 22504 -924 23104 -624
rect 12184 -1156 22840 -1046
rect 11705 -2715 11795 -2625
rect 11488 -3564 11588 -3464
rect 16988 -2462 17048 -2402
rect 15844 -2702 15904 -2642
rect 19894 -2700 19950 -2644
rect 16070 -3540 16130 -3480
rect 21440 -3544 21498 -3484
rect 21498 -3544 21500 -3484
rect 16854 -3772 16914 -3712
rect 3902 -5450 7666 -5298
rect 15702 -5450 19466 -5298
rect 172 -5836 772 -5536
rect 10704 -5836 11304 -5536
rect 11972 -5836 12572 -5536
rect 22504 -5836 23104 -5536
<< metal3 >>
rect 162 5032 782 5037
rect 162 4732 172 5032
rect 772 4732 782 5032
rect 162 4727 782 4732
rect 10694 5032 11314 5037
rect 10694 4732 10704 5032
rect 11304 4732 11314 5032
rect 10694 4727 11314 4732
rect 11962 5032 12582 5037
rect 11962 4732 11972 5032
rect 12572 4732 12582 5032
rect 11962 4727 12582 4732
rect 22494 5032 23114 5037
rect 22494 4732 22504 5032
rect 23104 4732 23114 5032
rect 22494 4727 23114 4732
rect 3854 4646 7710 4686
rect 3854 4494 3902 4646
rect 7666 4494 7710 4646
rect 3854 4456 7710 4494
rect 15654 4646 19510 4686
rect 15654 4494 15702 4646
rect 19466 4494 19510 4646
rect 15654 4456 19510 4494
rect 9620 3264 17070 3284
rect 9620 3204 16982 3264
rect 17042 3204 17070 3264
rect 9620 3184 17070 3204
rect -592 2988 4752 3008
rect -592 2928 4668 2988
rect 4728 2928 4752 2988
rect -592 2908 4752 2928
rect -592 -3466 -492 2908
rect 9620 2740 9720 3184
rect 11488 2871 16550 2876
rect 11488 2781 11493 2871
rect 11583 2856 16550 2871
rect 11583 2796 16468 2856
rect 16528 2796 16550 2856
rect 11583 2781 16550 2796
rect 11488 2776 16550 2781
rect 9620 2680 9642 2740
rect 9702 2680 9720 2740
rect 9620 2660 9720 2680
rect 18128 2746 23682 2764
rect 18128 2686 18144 2746
rect 18204 2686 23682 2746
rect 18128 2664 23682 2686
rect -330 2010 1580 2030
rect -330 1950 1498 2010
rect 1558 1950 1580 2010
rect -330 1930 1580 1950
rect -330 -2450 -230 1930
rect 11695 1916 11805 1921
rect 4016 1898 11700 1916
rect 4016 1838 4044 1898
rect 4104 1896 11700 1898
rect 4104 1840 8094 1896
rect 8150 1840 11700 1896
rect 4104 1838 11700 1840
rect 4016 1816 11700 1838
rect 11800 1898 19974 1916
rect 11800 1838 15844 1898
rect 15904 1896 19974 1898
rect 15904 1840 19894 1896
rect 19950 1840 19974 1896
rect 15904 1838 19974 1840
rect 11800 1816 19974 1838
rect 11695 1811 11805 1816
rect 18890 1684 23412 1706
rect 18890 1624 18920 1684
rect 18980 1624 23412 1684
rect 18890 1606 23412 1624
rect 322 352 11096 400
rect 322 242 384 352
rect 11040 242 11096 352
rect 322 186 11096 242
rect 12122 352 22896 400
rect 12122 242 12184 352
rect 22840 242 22896 352
rect 12122 186 22896 242
rect 162 120 782 125
rect 162 -180 172 120
rect 772 -180 782 120
rect 162 -185 782 -180
rect 10694 120 11314 125
rect 10694 -180 10704 120
rect 11304 -180 11314 120
rect 10694 -185 11314 -180
rect 11962 120 12582 125
rect 11962 -180 11972 120
rect 12572 -180 12582 120
rect 11962 -185 12582 -180
rect 22494 120 23114 125
rect 22494 -180 22504 120
rect 23104 -180 23114 120
rect 22494 -185 23114 -180
rect 162 -624 782 -619
rect 162 -924 172 -624
rect 772 -924 782 -624
rect 162 -929 782 -924
rect 10694 -624 11314 -619
rect 10694 -924 10704 -624
rect 11304 -924 11314 -624
rect 10694 -929 11314 -924
rect 11962 -624 12582 -619
rect 11962 -924 11972 -624
rect 12572 -924 12582 -624
rect 11962 -929 12582 -924
rect 22494 -624 23114 -619
rect 22494 -924 22504 -624
rect 23104 -924 23114 -624
rect 22494 -929 23114 -924
rect 322 -1046 11096 -990
rect 322 -1156 384 -1046
rect 11040 -1156 11096 -1046
rect 322 -1204 11096 -1156
rect 12122 -1046 22896 -990
rect 12122 -1156 12184 -1046
rect 22840 -1156 22896 -1046
rect 12122 -1204 22896 -1156
rect 23312 -2384 23412 1606
rect 16958 -2402 23412 -2384
rect -330 -2550 3908 -2450
rect 16958 -2462 16988 -2402
rect 17048 -2462 23412 -2402
rect 16958 -2484 23412 -2462
rect 3808 -2896 3908 -2550
rect 4016 -2625 19974 -2620
rect 4016 -2642 11705 -2625
rect 4016 -2702 4044 -2642
rect 4104 -2644 11705 -2642
rect 4104 -2700 8094 -2644
rect 8150 -2700 11705 -2644
rect 4104 -2702 11705 -2700
rect 4016 -2715 11705 -2702
rect 11795 -2642 19974 -2625
rect 11795 -2702 15844 -2642
rect 15904 -2644 19974 -2642
rect 15904 -2700 19894 -2644
rect 19950 -2700 19974 -2644
rect 15904 -2702 19974 -2700
rect 11795 -2715 19974 -2702
rect 4016 -2720 19974 -2715
rect 3808 -2916 4358 -2896
rect 3808 -2976 4268 -2916
rect 4328 -2976 4358 -2916
rect 3808 -2996 4358 -2976
rect 11483 -3464 11593 -3459
rect -592 -3490 5138 -3466
rect -592 -3550 5054 -3490
rect 5114 -3550 5138 -3490
rect -592 -3566 5138 -3550
rect 9614 -3484 11488 -3464
rect 9614 -3544 9638 -3484
rect 9698 -3544 11488 -3484
rect 9614 -3564 11488 -3544
rect 11588 -3480 16158 -3464
rect 23582 -3466 23682 2664
rect 11588 -3540 16070 -3480
rect 16130 -3540 16158 -3480
rect 11588 -3564 16158 -3540
rect 21422 -3484 23682 -3466
rect 21422 -3544 21440 -3484
rect 21500 -3544 23682 -3484
rect 11483 -3569 11593 -3564
rect 21422 -3566 23682 -3544
rect 6324 -3712 16934 -3696
rect 6324 -3716 16854 -3712
rect 6324 -3776 6342 -3716
rect 6402 -3772 16854 -3716
rect 16914 -3772 16934 -3712
rect 6402 -3776 16934 -3772
rect 6324 -3796 16934 -3776
rect 3854 -5298 7710 -5260
rect 3854 -5450 3902 -5298
rect 7666 -5450 7710 -5298
rect 3854 -5490 7710 -5450
rect 15654 -5298 19510 -5260
rect 15654 -5450 15702 -5298
rect 19466 -5450 19510 -5298
rect 15654 -5490 19510 -5450
rect 162 -5536 782 -5531
rect 162 -5836 172 -5536
rect 772 -5836 782 -5536
rect 162 -5841 782 -5836
rect 10694 -5536 11314 -5531
rect 10694 -5836 10704 -5536
rect 11304 -5836 11314 -5536
rect 10694 -5841 11314 -5836
rect 11962 -5536 12582 -5531
rect 11962 -5836 11972 -5536
rect 12572 -5836 12582 -5536
rect 11962 -5841 12582 -5836
rect 22494 -5536 23114 -5531
rect 22494 -5836 22504 -5536
rect 23104 -5836 23114 -5536
rect 22494 -5841 23114 -5836
<< via3 >>
rect 172 4732 772 5032
rect 10704 4732 11304 5032
rect 11972 4732 12572 5032
rect 22504 4732 23104 5032
rect 3902 4494 7666 4646
rect 15702 4494 19466 4646
rect 384 242 11040 352
rect 12184 242 22840 352
rect 172 -180 772 120
rect 10704 -180 11304 120
rect 11972 -180 12572 120
rect 22504 -180 23104 120
rect 172 -924 772 -624
rect 10704 -924 11304 -624
rect 11972 -924 12572 -624
rect 22504 -924 23104 -624
rect 384 -1156 11040 -1046
rect 12184 -1156 22840 -1046
rect 3902 -5450 7666 -5298
rect 15702 -5450 19466 -5298
rect 172 -5836 772 -5536
rect 10704 -5836 11304 -5536
rect 11972 -5836 12572 -5536
rect 22504 -5836 23104 -5536
<< metal4 >>
rect -728 5032 23288 5216
rect -728 4732 172 5032
rect 772 4732 10704 5032
rect 11304 4732 11972 5032
rect 12572 4732 22504 5032
rect 23104 4732 23288 5032
rect -728 4646 23288 4732
rect -728 4494 3902 4646
rect 7666 4494 15702 4646
rect 19466 4494 23288 4646
rect -728 4416 23288 4494
rect -12 434 11488 436
rect 11788 434 23288 436
rect -12 352 23288 434
rect -12 242 384 352
rect 11040 242 12184 352
rect 22840 242 23288 352
rect -12 120 23288 242
rect -12 -180 172 120
rect 772 -180 10704 120
rect 11304 -180 11972 120
rect 12572 -180 22504 120
rect 23104 -180 23288 120
rect -12 -624 23288 -180
rect -12 -924 172 -624
rect 772 -924 10704 -624
rect 11304 -924 11972 -624
rect 12572 -924 22504 -624
rect 23104 -924 23288 -624
rect -12 -1046 23288 -924
rect -12 -1156 384 -1046
rect 11040 -1156 12184 -1046
rect 22840 -1156 23288 -1046
rect -12 -1240 23288 -1156
rect 11292 -1242 12036 -1240
rect -1528 -5246 23288 -5220
rect -1528 -5998 -1504 -5246
rect -752 -5298 23288 -5246
rect -752 -5450 3902 -5298
rect 7666 -5450 15702 -5298
rect 19466 -5450 23288 -5298
rect -752 -5536 23288 -5450
rect -752 -5836 172 -5536
rect 772 -5836 10704 -5536
rect 11304 -5836 11972 -5536
rect 12572 -5836 22504 -5536
rect 23104 -5836 23288 -5536
rect -752 -5998 23288 -5836
rect -1528 -6020 23288 -5998
<< via4 >>
rect -1528 4416 -728 5216
rect -1504 -5998 -752 -5246
<< metal5 >>
rect -1552 5216 -704 5240
rect -1552 4416 -1528 5216
rect -728 4416 -704 5216
rect -1552 4392 -704 4416
rect -1528 -5246 -728 4392
rect -1528 -5998 -1504 -5246
rect -752 -5998 -728 -5246
rect -1528 -6022 -728 -5998
<< labels >>
flabel metal2 4746 1978 4762 1992 1 FreeSans 480 0 0 0 vip
port 3 n
flabel metal2 5012 2710 5020 2724 1 FreeSans 480 0 0 0 vim
port 4 n
flabel metal3 11604 1874 11614 1882 1 FreeSans 480 0 0 0 vocm
port 6 n
flabel metal4 11516 5188 11546 5206 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel metal4 11416 -406 11440 -390 1 FreeSans 480 0 0 0 VSS
port 2 n ground bidirectional
flabel metal3 23620 1100 23640 1116 1 FreeSans 480 0 0 0 vfiltm
port 8 n
flabel metal3 23360 1060 23382 1076 1 FreeSans 480 0 0 0 vfiltp
port 7 n
flabel metal3 -562 1138 -542 1158 1 FreeSans 480 0 0 0 vintp
port 9 n
flabel metal3 -290 1124 -268 1144 1 FreeSans 480 0 0 0 vintm
port 10 n
flabel metal2 6858 1072 6874 1080 1 FreeSans 480 0 0 0 ibiasn1
port 5 n
flabel metal2 6844 -1890 6870 -1878 1 FreeSans 480 0 0 0 ibiasn2
port 11 n
flabel metal2 18656 -1896 18670 -1880 1 FreeSans 480 0 0 0 ibiasn3
port 12 n
flabel metal2 18640 1074 18656 1084 1 FreeSans 480 0 0 0 ibiasn4
port 13 n
flabel metal1 1432 1572 1450 1584 1 FreeSans 480 0 0 0 gm_c_stage_0/vtail_diff
flabel metal1 10022 1604 10038 1620 1 FreeSans 480 0 0 0 gm_c_stage_0/vbiasp
flabel metal1 10016 604 10032 614 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmn_tail2
flabel metal1 6590 590 6602 602 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmn_tail1
flabel metal1 1650 1074 1658 1082 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmc
flabel metal2 7266 1074 7280 1084 1 FreeSans 480 0 0 0 gm_c_stage_0/ibiasn
flabel metal2 9028 1864 9038 1878 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmn_tail2
flabel metal2 8816 2706 8828 2722 1 FreeSans 480 0 0 0 gm_c_stage_0/vom
flabel metal2 8470 1968 8492 1986 1 FreeSans 480 0 0 0 gm_c_stage_0/vocm
flabel metal2 8204 2820 8216 2830 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmcn2
flabel metal2 9026 2932 9036 2944 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmcn
flabel metal2 4756 3654 4762 3666 1 FreeSans 480 0 0 0 gm_c_stage_0/vbiasp
flabel metal2 5722 1860 5740 1876 1 FreeSans 480 0 0 0 gm_c_stage_0/vtail_diff
flabel metal2 5542 2708 5560 2724 1 FreeSans 480 0 0 0 gm_c_stage_0/vim
flabel metal2 4874 2820 4894 2832 1 FreeSans 480 0 0 0 gm_c_stage_0/vom
flabel metal2 5698 2934 5718 2950 1 FreeSans 480 0 0 0 gm_c_stage_0/vop
flabel metal2 2420 2926 2438 2946 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmcn1
flabel metal2 1524 2808 1544 2822 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmcn
flabel metal2 2244 2694 2266 2706 1 FreeSans 480 0 0 0 gm_c_stage_0/vocm
flabel metal2 1880 1976 1898 1988 1 FreeSans 480 0 0 0 gm_c_stage_0/vop
flabel metal2 2418 1862 2438 1878 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmn_tail1
flabel metal2 5072 1982 5080 1988 1 FreeSans 480 0 0 0 gm_c_stage_0/vip
flabel metal1 5716 4058 5734 4074 1 FreeSans 480 0 0 0 gm_c_stage_0/vcmc
flabel metal2 4694 3290 4700 3294 1 FreeSans 480 0 0 0 gm_c_stage_0/vom
flabel metal2 5206 3288 5212 3294 1 FreeSans 480 0 0 0 gm_c_stage_0/vop
flabel metal4 322 5192 334 5206 1 FreeSans 480 0 0 0 gm_c_stage_0/VDD
flabel metal4 560 -352 574 -338 1 FreeSans 480 0 0 0 gm_c_stage_0/VSS
flabel metal1 1432 -2388 1450 -2376 5 FreeSans 480 0 0 0 gm_c_stage_1/vtail_diff
flabel metal1 10022 -2424 10038 -2408 5 FreeSans 480 0 0 0 gm_c_stage_1/vbiasp
flabel metal1 10016 -1418 10032 -1408 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmn_tail2
flabel metal1 6590 -1406 6602 -1394 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmn_tail1
flabel metal1 1650 -1886 1658 -1878 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmc
flabel metal2 7266 -1888 7280 -1878 5 FreeSans 480 0 0 0 gm_c_stage_1/ibiasn
flabel metal2 9028 -2682 9038 -2668 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmn_tail2
flabel metal2 8816 -3526 8828 -3510 5 FreeSans 480 0 0 0 gm_c_stage_1/vom
flabel metal2 8470 -2790 8492 -2772 5 FreeSans 480 0 0 0 gm_c_stage_1/vocm
flabel metal2 8204 -3634 8216 -3624 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmcn2
flabel metal2 9026 -3748 9036 -3736 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmcn
flabel metal2 4756 -4470 4762 -4458 5 FreeSans 480 0 0 0 gm_c_stage_1/vbiasp
flabel metal2 5722 -2680 5740 -2664 5 FreeSans 480 0 0 0 gm_c_stage_1/vtail_diff
flabel metal2 5542 -3528 5560 -3512 5 FreeSans 480 0 0 0 gm_c_stage_1/vim
flabel metal2 4874 -3636 4894 -3624 5 FreeSans 480 0 0 0 gm_c_stage_1/vom
flabel metal2 5698 -3754 5718 -3738 5 FreeSans 480 0 0 0 gm_c_stage_1/vop
flabel metal2 2420 -3750 2438 -3730 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmcn1
flabel metal2 1524 -3626 1544 -3612 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmcn
flabel metal2 2244 -3510 2266 -3498 5 FreeSans 480 0 0 0 gm_c_stage_1/vocm
flabel metal2 1880 -2792 1898 -2780 5 FreeSans 480 0 0 0 gm_c_stage_1/vop
flabel metal2 2418 -2682 2438 -2666 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmn_tail1
flabel metal2 5072 -2792 5080 -2786 5 FreeSans 480 0 0 0 gm_c_stage_1/vip
flabel metal1 5716 -4878 5734 -4862 5 FreeSans 480 0 0 0 gm_c_stage_1/vcmc
flabel metal2 4694 -4098 4700 -4094 5 FreeSans 480 0 0 0 gm_c_stage_1/vom
flabel metal2 5206 -4098 5212 -4092 5 FreeSans 480 0 0 0 gm_c_stage_1/vop
flabel metal4 322 -6010 334 -5996 5 FreeSans 480 0 0 0 gm_c_stage_1/VDD
flabel metal4 560 -466 574 -452 5 FreeSans 480 0 0 0 gm_c_stage_1/VSS
flabel metal1 13232 -2388 13250 -2376 5 FreeSans 480 0 0 0 gm_c_stage_3/vtail_diff
flabel metal1 21822 -2424 21838 -2408 5 FreeSans 480 0 0 0 gm_c_stage_3/vbiasp
flabel metal1 21816 -1418 21832 -1408 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmn_tail2
flabel metal1 18390 -1406 18402 -1394 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmn_tail1
flabel metal1 13450 -1886 13458 -1878 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmc
flabel metal2 19066 -1888 19080 -1878 5 FreeSans 480 0 0 0 gm_c_stage_3/ibiasn
flabel metal2 20828 -2682 20838 -2668 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmn_tail2
flabel metal2 20616 -3526 20628 -3510 5 FreeSans 480 0 0 0 gm_c_stage_3/vom
flabel metal2 20270 -2790 20292 -2772 5 FreeSans 480 0 0 0 gm_c_stage_3/vocm
flabel metal2 20004 -3634 20016 -3624 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmcn2
flabel metal2 20826 -3748 20836 -3736 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmcn
flabel metal2 16556 -4470 16562 -4458 5 FreeSans 480 0 0 0 gm_c_stage_3/vbiasp
flabel metal2 17522 -2680 17540 -2664 5 FreeSans 480 0 0 0 gm_c_stage_3/vtail_diff
flabel metal2 17342 -3528 17360 -3512 5 FreeSans 480 0 0 0 gm_c_stage_3/vim
flabel metal2 16674 -3636 16694 -3624 5 FreeSans 480 0 0 0 gm_c_stage_3/vom
flabel metal2 17498 -3754 17518 -3738 5 FreeSans 480 0 0 0 gm_c_stage_3/vop
flabel metal2 14220 -3750 14238 -3730 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmcn1
flabel metal2 13324 -3626 13344 -3612 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmcn
flabel metal2 14044 -3510 14066 -3498 5 FreeSans 480 0 0 0 gm_c_stage_3/vocm
flabel metal2 13680 -2792 13698 -2780 5 FreeSans 480 0 0 0 gm_c_stage_3/vop
flabel metal2 14218 -2682 14238 -2666 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmn_tail1
flabel metal2 16872 -2792 16880 -2786 5 FreeSans 480 0 0 0 gm_c_stage_3/vip
flabel metal1 17516 -4878 17534 -4862 5 FreeSans 480 0 0 0 gm_c_stage_3/vcmc
flabel metal2 16494 -4098 16500 -4094 5 FreeSans 480 0 0 0 gm_c_stage_3/vom
flabel metal2 17006 -4098 17012 -4092 5 FreeSans 480 0 0 0 gm_c_stage_3/vop
flabel metal4 12122 -6010 12134 -5996 5 FreeSans 480 0 0 0 gm_c_stage_3/VDD
flabel metal4 12360 -466 12374 -452 5 FreeSans 480 0 0 0 gm_c_stage_3/VSS
flabel metal1 13232 1572 13250 1584 1 FreeSans 480 0 0 0 gm_c_stage_2/vtail_diff
flabel metal1 21822 1604 21838 1620 1 FreeSans 480 0 0 0 gm_c_stage_2/vbiasp
flabel metal1 21816 604 21832 614 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmn_tail2
flabel metal1 18390 590 18402 602 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmn_tail1
flabel metal1 13450 1074 13458 1082 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmc
flabel metal2 19066 1074 19080 1084 1 FreeSans 480 0 0 0 gm_c_stage_2/ibiasn
flabel metal2 20828 1864 20838 1878 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmn_tail2
flabel metal2 20616 2706 20628 2722 1 FreeSans 480 0 0 0 gm_c_stage_2/vom
flabel metal2 20270 1968 20292 1986 1 FreeSans 480 0 0 0 gm_c_stage_2/vocm
flabel metal2 20004 2820 20016 2830 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmcn2
flabel metal2 20826 2932 20836 2944 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmcn
flabel metal2 16556 3654 16562 3666 1 FreeSans 480 0 0 0 gm_c_stage_2/vbiasp
flabel metal2 17522 1860 17540 1876 1 FreeSans 480 0 0 0 gm_c_stage_2/vtail_diff
flabel metal2 17342 2708 17360 2724 1 FreeSans 480 0 0 0 gm_c_stage_2/vim
flabel metal2 16674 2820 16694 2832 1 FreeSans 480 0 0 0 gm_c_stage_2/vom
flabel metal2 17498 2934 17518 2950 1 FreeSans 480 0 0 0 gm_c_stage_2/vop
flabel metal2 14220 2926 14238 2946 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmcn1
flabel metal2 13324 2808 13344 2822 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmcn
flabel metal2 14044 2694 14066 2706 1 FreeSans 480 0 0 0 gm_c_stage_2/vocm
flabel metal2 13680 1976 13698 1988 1 FreeSans 480 0 0 0 gm_c_stage_2/vop
flabel metal2 14218 1862 14238 1878 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmn_tail1
flabel metal2 16872 1982 16880 1988 1 FreeSans 480 0 0 0 gm_c_stage_2/vip
flabel metal1 17516 4058 17534 4074 1 FreeSans 480 0 0 0 gm_c_stage_2/vcmc
flabel metal2 16494 3290 16500 3294 1 FreeSans 480 0 0 0 gm_c_stage_2/vom
flabel metal2 17006 3288 17012 3294 1 FreeSans 480 0 0 0 gm_c_stage_2/vop
flabel metal4 12122 5192 12134 5206 1 FreeSans 480 0 0 0 gm_c_stage_2/VDD
flabel metal4 12360 -352 12374 -338 1 FreeSans 480 0 0 0 gm_c_stage_2/VSS
<< end >>
