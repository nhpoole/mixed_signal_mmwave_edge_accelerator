magic
tech sky130A
magscale 1 2
timestamp 1622230533
<< nwell >>
rect -354 333 1930 654
<< pwell >>
rect -313 110 -227 267
rect 679 229 865 273
rect 1409 229 1880 275
rect -223 93 1880 229
rect -195 55 -161 93
<< scnmos >>
rect -145 119 -115 203
rect -61 119 -31 203
rect 194 119 224 203
rect 289 119 319 191
rect 385 119 415 191
rect 551 119 581 203
rect 623 119 653 203
rect 755 119 785 247
rect 854 119 884 191
rect 963 119 993 191
rect 1059 119 1089 203
rect 1208 119 1238 203
rect 1299 119 1329 203
rect 1487 119 1517 249
rect 1675 119 1705 203
rect 1772 119 1802 249
<< scpmoshvt >>
rect -145 435 -115 563
rect -61 435 -31 563
rect 206 485 236 569
rect 298 485 328 569
rect 397 485 427 569
rect 537 485 567 569
rect 634 485 664 569
rect 831 401 861 569
rect 930 485 960 569
rect 1016 485 1046 569
rect 1100 485 1130 569
rect 1208 485 1238 569
rect 1292 485 1322 569
rect 1456 369 1486 569
rect 1675 441 1705 569
rect 1772 369 1802 569
<< ndiff >>
rect -197 191 -145 203
rect -197 157 -189 191
rect -155 157 -145 191
rect -197 119 -145 157
rect -115 165 -61 203
rect -115 131 -105 165
rect -71 131 -61 165
rect -115 119 -61 131
rect -31 191 21 203
rect -31 157 -21 191
rect 13 157 21 191
rect -31 119 21 157
rect 89 161 194 203
rect 89 127 101 161
rect 135 127 194 161
rect 89 119 194 127
rect 224 191 274 203
rect 705 203 755 247
rect 433 191 551 203
rect 224 167 289 191
rect 224 133 234 167
rect 268 133 289 167
rect 224 119 289 133
rect 319 167 385 191
rect 319 133 341 167
rect 375 133 385 167
rect 319 119 385 133
rect 415 119 551 191
rect 581 119 623 203
rect 653 165 755 203
rect 653 131 687 165
rect 721 131 755 165
rect 653 119 755 131
rect 785 191 839 247
rect 1435 204 1487 249
rect 1009 191 1059 203
rect 785 161 854 191
rect 785 127 799 161
rect 833 127 854 161
rect 785 119 854 127
rect 884 165 963 191
rect 884 131 909 165
rect 943 131 963 165
rect 884 119 963 131
rect 993 119 1059 191
rect 1089 161 1208 203
rect 1089 127 1121 161
rect 1155 127 1208 161
rect 1089 119 1208 127
rect 1238 119 1299 203
rect 1329 181 1381 203
rect 1329 147 1339 181
rect 1373 147 1381 181
rect 1329 119 1381 147
rect 1435 170 1443 204
rect 1477 170 1487 204
rect 1435 119 1487 170
rect 1517 237 1569 249
rect 1517 203 1527 237
rect 1561 203 1569 237
rect 1720 203 1772 249
rect 1517 169 1569 203
rect 1517 135 1527 169
rect 1561 135 1569 169
rect 1517 119 1569 135
rect 1623 191 1675 203
rect 1623 157 1631 191
rect 1665 157 1675 191
rect 1623 119 1675 157
rect 1705 185 1772 203
rect 1705 151 1728 185
rect 1762 151 1772 185
rect 1705 119 1772 151
rect 1802 215 1854 249
rect 1802 181 1812 215
rect 1846 181 1854 215
rect 1802 119 1854 181
<< pdiff >>
rect -197 549 -145 563
rect -197 515 -189 549
rect -155 515 -145 549
rect -197 481 -145 515
rect -197 447 -189 481
rect -155 447 -145 481
rect -197 435 -145 447
rect -115 533 -61 563
rect -115 499 -105 533
rect -71 499 -61 533
rect -115 435 -61 499
rect -31 549 21 563
rect -31 515 -21 549
rect 13 515 21 549
rect -31 481 21 515
rect 154 557 206 569
rect 154 523 162 557
rect 196 523 206 557
rect 154 485 206 523
rect 236 549 298 569
rect 236 515 246 549
rect 280 515 298 549
rect 236 485 298 515
rect 328 555 397 569
rect 328 521 339 555
rect 373 521 397 555
rect 328 485 397 521
rect 427 531 537 569
rect 427 497 493 531
rect 527 497 537 531
rect 427 485 537 497
rect 567 547 634 569
rect 567 513 590 547
rect 624 513 634 547
rect 567 485 634 513
rect 664 531 716 569
rect 664 497 674 531
rect 708 497 716 531
rect 664 485 716 497
rect 779 557 831 569
rect 779 523 787 557
rect 821 523 831 557
rect -31 447 -21 481
rect 13 447 21 481
rect -31 435 21 447
rect 779 401 831 523
rect 861 549 930 569
rect 861 515 875 549
rect 909 515 930 549
rect 861 485 930 515
rect 960 556 1016 569
rect 960 522 972 556
rect 1006 522 1016 556
rect 960 485 1016 522
rect 1046 485 1100 569
rect 1130 557 1208 569
rect 1130 523 1164 557
rect 1198 523 1208 557
rect 1130 485 1208 523
rect 1238 531 1292 569
rect 1238 497 1248 531
rect 1282 497 1292 531
rect 1238 485 1292 497
rect 1322 557 1456 569
rect 1322 523 1334 557
rect 1368 523 1412 557
rect 1446 523 1456 557
rect 1322 485 1456 523
rect 861 401 915 485
rect 1406 369 1456 485
rect 1486 549 1542 569
rect 1486 515 1496 549
rect 1530 515 1542 549
rect 1486 481 1542 515
rect 1486 447 1496 481
rect 1530 447 1542 481
rect 1486 413 1542 447
rect 1623 557 1675 569
rect 1623 523 1631 557
rect 1665 523 1675 557
rect 1623 489 1675 523
rect 1623 455 1631 489
rect 1665 455 1675 489
rect 1623 441 1675 455
rect 1705 557 1772 569
rect 1705 523 1728 557
rect 1762 523 1772 557
rect 1705 489 1772 523
rect 1705 455 1728 489
rect 1762 455 1772 489
rect 1705 441 1772 455
rect 1486 379 1496 413
rect 1530 379 1542 413
rect 1486 369 1542 379
rect 1720 421 1772 441
rect 1720 387 1728 421
rect 1762 387 1772 421
rect 1720 369 1772 387
rect 1802 521 1854 569
rect 1802 487 1812 521
rect 1846 487 1854 521
rect 1802 453 1854 487
rect 1802 419 1812 453
rect 1846 419 1854 453
rect 1802 369 1854 419
<< ndiffc >>
rect -189 157 -155 191
rect -105 131 -71 165
rect -21 157 13 191
rect 101 127 135 161
rect 234 133 268 167
rect 341 133 375 167
rect 687 131 721 165
rect 799 127 833 161
rect 909 131 943 165
rect 1121 127 1155 161
rect 1339 147 1373 181
rect 1443 170 1477 204
rect 1527 203 1561 237
rect 1527 135 1561 169
rect 1631 157 1665 191
rect 1728 151 1762 185
rect 1812 181 1846 215
<< pdiffc >>
rect -189 515 -155 549
rect -189 447 -155 481
rect -105 499 -71 533
rect -21 515 13 549
rect 162 523 196 557
rect 246 515 280 549
rect 339 521 373 555
rect 493 497 527 531
rect 590 513 624 547
rect 674 497 708 531
rect 787 523 821 557
rect -21 447 13 481
rect 875 515 909 549
rect 972 522 1006 556
rect 1164 523 1198 557
rect 1248 497 1282 531
rect 1334 523 1368 557
rect 1412 523 1446 557
rect 1496 515 1530 549
rect 1496 447 1530 481
rect 1631 523 1665 557
rect 1631 455 1665 489
rect 1728 523 1762 557
rect 1728 455 1762 489
rect 1496 379 1530 413
rect 1728 387 1762 421
rect 1812 487 1846 521
rect 1812 419 1846 453
<< psubdiff >>
rect -287 217 -253 241
rect -287 136 -253 183
<< nsubdiff >>
rect -287 528 -253 552
rect -287 435 -253 494
rect -287 377 -253 401
<< psubdiffcont >>
rect -287 183 -253 217
<< nsubdiffcont >>
rect -287 494 -253 528
rect -287 401 -253 435
<< poly >>
rect -145 563 -115 589
rect -61 563 -31 589
rect 206 569 236 595
rect 298 569 328 595
rect 397 569 427 595
rect 537 569 567 595
rect 634 569 664 595
rect 831 569 861 595
rect 930 569 960 595
rect 1016 569 1046 595
rect 1100 569 1130 595
rect 1208 569 1238 595
rect 1292 569 1322 595
rect 1456 569 1486 595
rect 1675 569 1705 595
rect 1772 569 1802 595
rect -145 420 -115 435
rect -178 390 -115 420
rect -178 337 -148 390
rect -61 346 -31 435
rect 206 398 236 485
rect 298 447 328 485
rect -202 321 -148 337
rect -202 287 -192 321
rect -158 287 -148 321
rect -106 336 -31 346
rect -106 302 -90 336
rect -56 302 -31 336
rect 107 382 236 398
rect 282 437 348 447
rect 282 403 298 437
rect 332 403 348 437
rect 282 393 348 403
rect 107 348 117 382
rect 151 368 236 382
rect 151 348 224 368
rect 397 351 427 485
rect 537 427 567 485
rect 537 411 592 427
rect 537 377 547 411
rect 581 377 592 411
rect 537 361 592 377
rect 107 332 224 348
rect -106 292 -31 302
rect -202 271 -148 287
rect -178 248 -148 271
rect -178 218 -115 248
rect -145 203 -115 218
rect -61 203 -31 292
rect 194 203 224 332
rect 289 321 427 351
rect 289 291 320 321
rect 266 275 320 291
rect 266 241 276 275
rect 310 241 320 275
rect 266 225 320 241
rect 362 269 428 279
rect 362 235 378 269
rect 412 235 428 269
rect 362 225 428 235
rect 289 191 319 225
rect 385 191 415 225
rect 551 203 581 361
rect 634 291 664 485
rect 831 386 861 401
rect 755 356 861 386
rect 755 339 785 356
rect 719 323 785 339
rect 623 275 677 291
rect 623 241 633 275
rect 667 241 677 275
rect 719 289 729 323
rect 763 289 785 323
rect 930 351 960 485
rect 1016 453 1046 485
rect 1002 437 1056 453
rect 1002 403 1012 437
rect 1046 403 1056 437
rect 1002 387 1056 403
rect 930 339 980 351
rect 930 327 993 339
rect 930 321 1017 327
rect 951 311 1017 321
rect 951 309 973 311
rect 719 273 785 289
rect 755 247 785 273
rect 854 263 921 279
rect 623 225 677 241
rect 623 203 653 225
rect 854 229 877 263
rect 911 229 921 263
rect 854 213 921 229
rect 963 277 973 309
rect 1007 277 1017 311
rect 963 261 1017 277
rect 1100 301 1130 485
rect 1208 329 1238 485
rect 1292 437 1322 485
rect 1280 421 1334 437
rect 1280 387 1290 421
rect 1324 387 1334 421
rect 1280 371 1334 387
rect 1203 313 1257 329
rect 1100 285 1161 301
rect 1100 265 1117 285
rect 854 191 884 213
rect 963 191 993 261
rect 1059 251 1117 265
rect 1151 251 1161 285
rect 1203 279 1213 313
rect 1247 279 1257 313
rect 1203 263 1257 279
rect 1059 235 1161 251
rect 1059 203 1089 235
rect 1208 203 1238 263
rect 1299 203 1329 371
rect 1675 405 1705 441
rect 1664 375 1705 405
rect 1456 337 1486 369
rect 1664 337 1694 375
rect 1772 337 1802 369
rect 1385 321 1694 337
rect 1385 287 1413 321
rect 1447 287 1694 321
rect 1385 271 1694 287
rect 1743 321 1802 337
rect 1743 287 1753 321
rect 1787 287 1802 321
rect 1743 271 1802 287
rect 1487 249 1517 271
rect 1664 248 1694 271
rect 1772 249 1802 271
rect 1664 218 1705 248
rect 1675 203 1705 218
rect -145 93 -115 119
rect -61 93 -31 119
rect 194 93 224 119
rect 289 93 319 119
rect 385 93 415 119
rect 551 93 581 119
rect 623 93 653 119
rect 755 93 785 119
rect 854 93 884 119
rect 963 93 993 119
rect 1059 93 1089 119
rect 1208 93 1238 119
rect 1299 93 1329 119
rect 1487 93 1517 119
rect 1675 93 1705 119
rect 1772 93 1802 119
<< polycont >>
rect -192 287 -158 321
rect -90 302 -56 336
rect 298 403 332 437
rect 117 348 151 382
rect 547 377 581 411
rect 276 241 310 275
rect 378 235 412 269
rect 633 241 667 275
rect 729 289 763 323
rect 1012 403 1046 437
rect 877 229 911 263
rect 973 277 1007 311
rect 1290 387 1324 421
rect 1117 251 1151 285
rect 1213 279 1247 313
rect 1413 287 1447 321
rect 1753 287 1787 321
<< locali >>
rect -316 599 -287 633
rect -253 599 -195 633
rect -161 599 -103 633
rect -69 599 -11 633
rect 23 599 81 633
rect 115 599 173 633
rect 207 599 265 633
rect 299 599 357 633
rect 391 599 449 633
rect 483 599 541 633
rect 575 599 633 633
rect 667 599 725 633
rect 759 599 817 633
rect 851 599 909 633
rect 943 599 1001 633
rect 1035 599 1093 633
rect 1127 599 1185 633
rect 1219 599 1277 633
rect 1311 599 1369 633
rect 1403 599 1461 633
rect 1495 599 1553 633
rect 1587 599 1645 633
rect 1679 599 1737 633
rect 1771 599 1829 633
rect 1863 599 1892 633
rect -299 528 -241 599
rect -299 494 -287 528
rect -253 494 -241 528
rect -299 435 -241 494
rect -299 401 -287 435
rect -253 401 -241 435
rect -206 549 -155 565
rect -206 515 -189 549
rect -206 481 -155 515
rect -121 533 -55 599
rect -121 499 -105 533
rect -71 499 -55 533
rect -21 549 13 565
rect -206 447 -189 481
rect -21 481 13 515
rect -155 447 -56 465
rect -206 431 -56 447
rect -299 366 -241 401
rect -206 338 -136 397
rect -206 290 -202 338
rect -154 290 -136 338
rect -206 287 -192 290
rect -158 287 -136 290
rect -206 267 -136 287
rect -102 336 -56 431
rect -102 327 -90 336
rect -68 293 -56 302
rect -299 217 -241 234
rect -102 233 -56 293
rect -299 183 -287 217
rect -253 183 -241 217
rect -299 89 -241 183
rect -206 199 -56 233
rect -206 191 -155 199
rect -206 157 -189 191
rect -21 191 13 429
rect 47 531 112 562
rect 47 497 73 531
rect 107 497 112 531
rect 146 557 196 599
rect 146 523 162 557
rect 146 507 196 523
rect 230 549 280 565
rect 230 515 246 549
rect 47 405 112 497
rect 230 499 280 515
rect 323 555 459 565
rect 323 521 339 555
rect 373 521 459 555
rect 574 547 640 599
rect 767 557 841 599
rect 323 499 459 521
rect 230 473 264 499
rect 185 439 264 473
rect 298 463 391 465
rect 59 382 151 405
rect 59 348 117 382
rect 59 195 151 348
rect -206 141 -155 157
rect -121 131 -105 165
rect -71 131 -55 165
rect 185 167 219 439
rect 298 437 357 463
rect 332 429 357 437
rect 332 403 391 429
rect 298 387 391 403
rect 253 327 323 349
rect 253 293 265 327
rect 299 293 323 327
rect 253 275 323 293
rect 253 241 276 275
rect 310 241 323 275
rect 253 225 323 241
rect 357 269 391 387
rect 425 343 459 499
rect 493 531 527 547
rect 574 513 590 547
rect 624 513 640 547
rect 674 531 708 547
rect 493 479 527 497
rect 767 523 787 557
rect 821 523 841 557
rect 767 507 841 523
rect 875 549 909 565
rect 674 479 708 497
rect 493 445 708 479
rect 875 473 909 515
rect 956 556 1130 565
rect 956 522 972 556
rect 1006 522 1130 556
rect 956 497 1130 522
rect 1164 557 1214 599
rect 1198 523 1214 557
rect 1318 557 1462 599
rect 1164 507 1214 523
rect 1248 531 1282 547
rect 797 439 909 473
rect 797 411 831 439
rect 531 377 547 411
rect 581 377 831 411
rect 970 429 981 463
rect 1015 437 1062 463
rect 970 405 1012 429
rect 425 323 763 343
rect 425 309 729 323
rect 357 235 378 269
rect 412 235 428 269
rect 357 225 428 235
rect 462 167 496 309
rect 537 259 633 275
rect 571 225 609 259
rect 667 241 695 275
rect 729 273 763 289
rect 643 225 695 241
rect 797 239 831 377
rect -21 141 13 157
rect -121 89 -55 131
rect 85 127 101 161
rect 135 127 151 161
rect 185 133 234 167
rect 268 133 284 167
rect 325 133 341 167
rect 375 133 496 167
rect 671 165 737 181
rect 85 89 151 127
rect 671 131 687 165
rect 721 131 737 165
rect 671 89 737 131
rect 779 161 831 239
rect 869 403 1012 405
rect 1046 403 1062 437
rect 1096 421 1130 497
rect 1318 523 1334 557
rect 1368 523 1412 557
rect 1446 523 1462 557
rect 1496 549 1577 565
rect 1728 557 1762 599
rect 1248 489 1282 497
rect 1530 515 1577 549
rect 1248 455 1408 489
rect 869 371 1004 403
rect 1096 387 1290 421
rect 1324 387 1340 421
rect 869 263 911 371
rect 1096 369 1130 387
rect 869 229 877 263
rect 869 213 911 229
rect 945 327 1015 337
rect 945 311 981 327
rect 945 277 973 311
rect 1007 277 1015 293
rect 945 213 1015 277
rect 1049 335 1130 369
rect 1049 179 1083 335
rect 1197 322 1305 353
rect 1374 337 1408 455
rect 1496 481 1577 515
rect 1530 456 1577 481
rect 1496 414 1519 447
rect 1561 414 1577 456
rect 1496 413 1577 414
rect 1530 379 1577 413
rect 1496 363 1577 379
rect 1374 331 1463 337
rect 1231 313 1305 322
rect 1117 285 1161 301
rect 1151 251 1161 285
rect 1197 279 1213 288
rect 1247 279 1305 313
rect 1117 245 1161 251
rect 1257 259 1305 279
rect 1117 211 1223 245
rect 893 165 1083 179
rect 779 127 799 161
rect 833 127 849 161
rect 893 131 909 165
rect 943 131 1083 165
rect 893 123 1083 131
rect 1117 161 1155 177
rect 1117 127 1121 161
rect 1189 165 1223 211
rect 1291 225 1305 259
rect 1257 199 1305 225
rect 1339 321 1463 331
rect 1339 287 1413 321
rect 1447 287 1463 321
rect 1339 271 1463 287
rect 1339 236 1404 271
rect 1511 237 1577 363
rect 1339 181 1403 236
rect 1189 147 1339 165
rect 1373 147 1403 181
rect 1189 131 1403 147
rect 1443 204 1477 226
rect 1117 89 1155 127
rect 1443 89 1477 170
rect 1511 203 1527 237
rect 1561 203 1577 237
rect 1511 169 1577 203
rect 1511 135 1527 169
rect 1561 135 1577 169
rect 1615 523 1631 557
rect 1665 523 1681 557
rect 1615 489 1681 523
rect 1615 455 1631 489
rect 1665 455 1681 489
rect 1615 337 1681 455
rect 1728 489 1762 523
rect 1728 421 1762 455
rect 1728 371 1762 387
rect 1812 521 1863 537
rect 1846 487 1863 521
rect 1812 453 1863 487
rect 1846 419 1863 453
rect 1812 361 1863 419
rect 1615 321 1787 337
rect 1615 287 1753 321
rect 1615 271 1787 287
rect 1821 317 1863 361
rect 1821 283 1835 317
rect 1615 191 1665 271
rect 1821 231 1863 283
rect 1812 215 1863 231
rect 1615 157 1631 191
rect 1615 141 1665 157
rect 1728 185 1762 208
rect 1511 127 1577 135
rect 1728 89 1762 151
rect 1846 181 1863 215
rect 1812 125 1863 181
rect -316 55 -287 89
rect -253 55 -195 89
rect -161 55 -103 89
rect -69 55 -11 89
rect 23 55 81 89
rect 115 55 173 89
rect 207 55 265 89
rect 299 55 357 89
rect 391 55 449 89
rect 483 55 541 89
rect 575 55 633 89
rect 667 55 725 89
rect 759 55 817 89
rect 851 55 909 89
rect 943 55 1001 89
rect 1035 55 1093 89
rect 1127 55 1185 89
rect 1219 55 1277 89
rect 1311 55 1369 89
rect 1403 55 1461 89
rect 1495 55 1553 89
rect 1587 55 1645 89
rect 1679 55 1737 89
rect 1771 55 1829 89
rect 1863 55 1892 89
<< viali >>
rect -287 599 -253 633
rect -195 599 -161 633
rect -103 599 -69 633
rect -11 599 23 633
rect 81 599 115 633
rect 173 599 207 633
rect 265 599 299 633
rect 357 599 391 633
rect 449 599 483 633
rect 541 599 575 633
rect 633 599 667 633
rect 725 599 759 633
rect 817 599 851 633
rect 909 599 943 633
rect 1001 599 1035 633
rect 1093 599 1127 633
rect 1185 599 1219 633
rect 1277 599 1311 633
rect 1369 599 1403 633
rect 1461 599 1495 633
rect 1553 599 1587 633
rect 1645 599 1679 633
rect 1737 599 1771 633
rect 1829 599 1863 633
rect -202 321 -154 338
rect -202 290 -192 321
rect -192 290 -158 321
rect -158 290 -154 321
rect -102 302 -90 327
rect -90 302 -68 327
rect -102 293 -68 302
rect -21 447 13 463
rect -21 429 13 447
rect 73 497 107 531
rect 357 429 391 463
rect 265 293 299 327
rect 981 437 1015 463
rect 981 429 1012 437
rect 1012 429 1015 437
rect 537 225 571 259
rect 609 241 633 259
rect 633 241 643 259
rect 609 225 643 241
rect 981 311 1015 327
rect 981 293 1007 311
rect 1007 293 1015 311
rect 1519 447 1530 456
rect 1530 447 1561 456
rect 1519 414 1561 447
rect 1197 313 1231 322
rect 1197 288 1213 313
rect 1213 288 1231 313
rect 1257 225 1291 259
rect 1835 283 1869 317
rect -287 55 -253 89
rect -195 55 -161 89
rect -103 55 -69 89
rect -11 55 23 89
rect 81 55 115 89
rect 173 55 207 89
rect 265 55 299 89
rect 357 55 391 89
rect 449 55 483 89
rect 541 55 575 89
rect 633 55 667 89
rect 725 55 759 89
rect 817 55 851 89
rect 909 55 943 89
rect 1001 55 1035 89
rect 1093 55 1127 89
rect 1185 55 1219 89
rect 1277 55 1311 89
rect 1369 55 1403 89
rect 1461 55 1495 89
rect 1553 55 1587 89
rect 1645 55 1679 89
rect 1737 55 1771 89
rect 1829 55 1863 89
<< metal1 >>
rect 1698 664 2104 668
rect -316 633 2104 664
rect -316 599 -287 633
rect -253 599 -195 633
rect -161 599 -103 633
rect -69 599 -11 633
rect 23 599 81 633
rect 115 599 173 633
rect 207 599 265 633
rect 299 599 357 633
rect 391 599 449 633
rect 483 599 541 633
rect 575 599 633 633
rect 667 599 725 633
rect 759 599 817 633
rect 851 599 909 633
rect 943 599 1001 633
rect 1035 599 1093 633
rect 1127 599 1185 633
rect 1219 599 1277 633
rect 1311 599 1369 633
rect 1403 599 1461 633
rect 1495 599 1553 633
rect 1587 599 1645 633
rect 1679 599 1737 633
rect 1771 599 1829 633
rect 1863 599 2104 633
rect -316 570 2104 599
rect -316 568 1892 570
rect 61 531 119 537
rect 61 530 73 531
rect -366 498 73 530
rect 61 497 73 498
rect 107 497 119 531
rect 61 491 119 497
rect -33 463 25 469
rect -33 429 -21 463
rect 13 460 25 463
rect 345 463 403 469
rect 345 460 357 463
rect 13 432 357 460
rect 13 429 25 432
rect -33 423 25 429
rect 345 429 357 432
rect 391 460 403 463
rect 969 463 1027 469
rect 969 460 981 463
rect 391 432 981 460
rect 391 429 403 432
rect 345 423 403 429
rect 969 429 981 432
rect 1015 429 1027 463
rect 969 423 1027 429
rect 1507 456 1980 462
rect 1507 414 1519 456
rect 1561 414 1980 456
rect 1507 408 1980 414
rect -342 338 -142 344
rect -342 290 -202 338
rect -154 290 -142 338
rect -342 284 -142 290
rect -114 327 -56 333
rect -114 293 -102 327
rect -68 324 -56 327
rect 253 327 311 333
rect 253 324 265 327
rect -68 296 265 324
rect -68 293 -56 296
rect -114 287 -56 293
rect 253 293 265 296
rect 299 324 311 327
rect 969 327 1027 333
rect 1186 328 1192 378
rect 969 324 981 327
rect 299 296 981 324
rect 299 293 311 296
rect 253 287 311 293
rect 969 293 981 296
rect 1015 293 1027 327
rect 969 287 1027 293
rect 1185 314 1192 328
rect 1256 314 1262 378
rect 1823 322 1881 323
rect 1823 317 2062 322
rect 1185 288 1197 314
rect 1231 288 1243 314
rect 1185 265 1243 288
rect 1823 283 1835 317
rect 1869 283 2062 317
rect 1823 278 2062 283
rect 1823 277 1881 278
rect 525 259 655 265
rect 525 225 537 259
rect 571 225 609 259
rect 643 256 655 259
rect 1185 259 1303 265
rect 1185 256 1257 259
rect 643 228 1257 256
rect 643 225 655 228
rect 525 219 655 225
rect 1245 225 1257 228
rect 1291 225 1303 259
rect 1245 219 1303 225
rect -316 118 1892 120
rect -316 89 2116 118
rect -316 55 -287 89
rect -253 55 -195 89
rect -161 55 -103 89
rect -69 55 -11 89
rect 23 55 81 89
rect 115 55 173 89
rect 207 55 265 89
rect 299 55 357 89
rect 391 55 449 89
rect 483 55 541 89
rect 575 55 633 89
rect 667 55 725 89
rect 759 55 817 89
rect 851 55 909 89
rect 943 55 1001 89
rect 1035 55 1093 89
rect 1127 55 1185 89
rect 1219 55 1277 89
rect 1311 55 1369 89
rect 1403 55 1461 89
rect 1495 55 1553 89
rect 1587 55 1645 89
rect 1679 55 1737 89
rect 1771 55 1829 89
rect 1863 55 2116 89
rect -316 24 2116 55
rect 1858 22 2116 24
<< via1 >>
rect 1192 322 1256 378
rect 1192 314 1197 322
rect 1197 314 1231 322
rect 1231 314 1256 322
<< metal2 >>
rect 1192 378 1256 384
rect 1256 314 1460 378
rect 1192 308 1256 314
rect 1396 -118 1460 314
<< labels >>
flabel metal1 -300 312 -294 320 1 FreeSans 480 0 0 0 CLK
port 2 n
flabel metal1 -320 512 -312 516 1 FreeSans 480 0 0 0 D
port 1 n
flabel metal2 1414 -50 1424 -42 1 FreeSans 480 0 0 0 RN
port 5 n
flabel metal1 1948 434 1956 440 1 FreeSans 480 0 0 0 Q
port 3 n
flabel metal1 2002 298 2010 304 1 FreeSans 480 0 0 0 QB
port 4 n
flabel metal1 2052 604 2060 610 1 FreeSans 480 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 2048 68 2066 76 1 FreeSans 480 0 0 0 VSS
port 7 n ground bidirectional
flabel locali 1530 290 1559 325 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/Q
flabel locali 1832 293 1854 326 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/Q_N
flabel locali 1257 225 1291 259 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 81 361 115 395 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/D
flabel locali -194 361 -160 395 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali -194 293 -160 327 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 1257 293 1291 327 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel metal1 -195 55 -161 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VGND
flabel metal1 -195 599 -161 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VPWR
flabel nwell -195 599 -161 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VPB
flabel pwell -195 55 -161 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VNB
rlabel comment -224 72 -224 72 4 sky130_fd_sc_hd__dfrbp_1_0/dfrbp_1
rlabel viali 1257 225 1291 259 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel viali 1197 288 1231 322 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 1257 199 1305 279 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 1197 279 1305 353 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1245 219 1303 228 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1185 265 1243 328 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1185 256 1303 265 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 525 256 655 265 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 525 228 1303 256 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 525 219 655 228 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel metal1 -294 596 -241 625 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -295 54 -244 92 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment -316 72 -316 72 4 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
<< end >>
