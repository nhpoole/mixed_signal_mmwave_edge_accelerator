magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< nwell >>
rect -3358 582 3358 3158
<< pwell >>
rect -3358 -3558 3358 418
<< psubdiff >>
rect -3322 282 -3160 382
rect 3160 282 3322 382
rect -3322 220 -3222 282
rect 3222 220 3322 282
rect -3122 82 -2960 182
rect -240 82 -78 182
rect -3122 20 -3022 82
rect -3122 -1002 -3022 -940
rect -178 20 -78 82
rect -178 -1002 -78 -940
rect -3122 -1102 -2960 -1002
rect -240 -1102 -78 -1002
rect -3122 -1318 -2960 -1218
rect 2960 -1318 3122 -1218
rect -3122 -1380 -3022 -1318
rect -3122 -2642 -3022 -2580
rect 3022 -1380 3122 -1318
rect 3022 -2642 3122 -2580
rect -3122 -2742 -2960 -2642
rect 2960 -2742 3122 -2642
rect -3322 -3422 -3222 -3360
rect 3222 -3422 3322 -3360
rect -3322 -3522 -3160 -3422
rect 3160 -3522 3322 -3422
<< nsubdiff >>
rect -3322 3022 -3160 3122
rect 3160 3022 3322 3122
rect -3322 2960 -3222 3022
rect -3322 718 -3222 780
rect 3222 2960 3322 3022
rect 3222 718 3322 780
rect -3322 618 -3160 718
rect 3160 618 3322 718
<< psubdiffcont >>
rect -3160 282 3160 382
rect -3322 -3360 -3222 220
rect -2960 82 -240 182
rect -3122 -940 -3022 20
rect -178 -940 -78 20
rect -2960 -1102 -240 -1002
rect -2960 -1318 2960 -1218
rect -3122 -2580 -3022 -1380
rect 3022 -2580 3122 -1380
rect -2960 -2742 2960 -2642
rect 3222 -3360 3322 220
rect -3160 -3522 3160 -3422
<< nsubdiffcont >>
rect -3160 3022 3160 3122
rect -3322 780 -3222 2960
rect 3222 780 3322 2960
rect -3160 618 3160 718
<< locali >>
rect -3322 2960 -3222 3122
rect -3322 618 -3222 780
rect 3222 2960 3322 3122
rect 3222 618 3322 780
rect -3322 220 -3222 382
rect 3222 220 3322 382
rect -3122 28 -3022 182
rect -3122 -1102 -3022 -948
rect -178 28 -78 182
rect -178 -1102 -78 -948
rect -3122 -1380 -3022 -1218
rect -3122 -2742 -3022 -2580
rect 3022 -1380 3122 -1218
rect 3022 -2742 3122 -2580
rect -3322 -3522 -3222 -3360
rect 3222 -3522 3322 -3360
<< viali >>
rect -3222 3022 -3160 3122
rect -3160 3022 3160 3122
rect 3160 3022 3222 3122
rect -3322 833 -3222 2907
rect 3222 833 3322 2907
rect -3222 618 -3160 718
rect -3160 618 3160 718
rect 3160 618 3222 718
rect -3222 282 -3160 382
rect -3160 282 3160 382
rect 3160 282 3222 382
rect -3322 -3237 -3222 97
rect -3022 82 -2960 182
rect -2960 82 -240 182
rect -240 82 -178 182
rect -3122 20 -3022 28
rect -3122 -940 -3022 20
rect -3122 -948 -3022 -940
rect -178 20 -78 28
rect -178 -940 -78 20
rect -178 -948 -78 -940
rect -3022 -1102 -2960 -1002
rect -2960 -1102 -240 -1002
rect -240 -1102 -178 -1002
rect -3022 -1318 -2960 -1218
rect -2960 -1318 2960 -1218
rect 2960 -1318 3022 -1218
rect -3122 -2576 -3022 -1384
rect 3022 -2576 3122 -1384
rect -3022 -2742 -2960 -2642
rect -2960 -2742 2960 -2642
rect 2960 -2742 3022 -2642
rect 3222 -3237 3322 97
rect -3222 -3522 -3160 -3422
rect -3160 -3522 3160 -3422
rect 3160 -3522 3222 -3422
<< metal1 >>
rect -3328 3122 3328 3128
rect -3328 3022 -3222 3122
rect 3222 3022 3328 3122
rect -3328 3016 3328 3022
rect -3328 2907 -3216 3016
rect -3328 833 -3322 2907
rect -3222 833 -3216 2907
rect -2616 2716 -2606 3016
rect 2606 2716 2616 3016
rect 3216 2907 3328 3016
rect -2674 2528 2566 2562
rect -2674 2456 -2646 2528
rect 2544 2456 2566 2528
rect -2674 2430 2566 2456
rect -2782 2146 -2776 2206
rect -2716 2146 -2710 2206
rect -2776 978 -2716 2146
rect -2654 1602 -2594 2430
rect -2528 1602 -2468 1764
rect -2400 1602 -2340 2430
rect -2272 2146 -2266 2206
rect -2206 2146 -2200 2206
rect -2266 2056 -2206 2146
rect -2270 1664 -2210 1766
rect -2276 1604 -2270 1664
rect -2210 1604 -2204 1664
rect -2654 1542 -2340 1602
rect -2654 1318 -2594 1542
rect -2528 1390 -2468 1542
rect -2400 1284 -2340 1542
rect -2270 1388 -2210 1604
rect -2138 1530 -2078 1890
rect -2008 1530 -1948 1768
rect -2144 1470 -2138 1530
rect -2078 1470 -2072 1530
rect -2014 1470 -2008 1530
rect -1948 1470 -1942 1530
rect -2008 1392 -1948 1470
rect -1880 1292 -1820 2430
rect -1628 2146 -1622 2206
rect -1562 2146 -1556 2206
rect -1502 2146 -1496 2206
rect -1436 2146 -1430 2206
rect -1622 1966 -1562 2146
rect -1496 2060 -1436 2146
rect -1750 1530 -1690 1770
rect -1494 1664 -1434 1766
rect -1500 1604 -1494 1664
rect -1434 1604 -1428 1664
rect -1756 1470 -1750 1530
rect -1690 1470 -1684 1530
rect -1634 1470 -1628 1530
rect -1568 1470 -1562 1530
rect -1750 1386 -1690 1470
rect -1628 1280 -1568 1470
rect -1494 1388 -1434 1604
rect -1366 1298 -1306 2430
rect -1238 2146 -1232 2206
rect -1172 2146 -1166 2206
rect -1232 2060 -1172 2146
rect -1240 1664 -1180 1766
rect -1246 1604 -1240 1664
rect -1180 1604 -1174 1664
rect -1240 1392 -1180 1604
rect -1112 1530 -1052 1872
rect -980 1530 -920 1770
rect -1118 1470 -1112 1530
rect -1052 1470 -1046 1530
rect -986 1470 -980 1530
rect -920 1470 -914 1530
rect -980 1386 -920 1470
rect -846 1284 -786 2430
rect -602 2146 -596 2206
rect -536 2146 -530 2206
rect -470 2146 -464 2206
rect -404 2146 -398 2206
rect -596 1940 -536 2146
rect -464 2056 -404 2146
rect -720 1530 -660 1766
rect -464 1664 -404 1766
rect -470 1604 -464 1664
rect -404 1604 -398 1664
rect -726 1470 -720 1530
rect -660 1470 -654 1530
rect -602 1470 -596 1530
rect -536 1470 -530 1530
rect -720 1388 -660 1470
rect -596 1272 -536 1470
rect -464 1388 -404 1604
rect -334 1598 -274 2430
rect -210 1598 -150 1768
rect -76 1598 -16 2430
rect 210 2258 216 2318
rect 276 2258 282 2318
rect 594 2258 600 2318
rect 660 2258 666 2318
rect -334 1538 -16 1598
rect -334 1276 -274 1538
rect -210 1390 -150 1538
rect -76 1302 -16 1538
rect -2274 978 -2214 1088
rect -2142 978 -2082 1198
rect -2782 918 -2776 978
rect -2716 918 -2710 978
rect -2280 918 -2274 978
rect -2214 918 -2208 978
rect -2148 918 -2142 978
rect -2082 918 -2076 978
rect -2014 874 -1954 1090
rect -1500 978 -1440 1094
rect -1240 978 -1180 1092
rect -1108 978 -1048 1190
rect -1506 918 -1500 978
rect -1440 918 -1434 978
rect -1246 918 -1240 978
rect -1180 918 -1174 978
rect -1114 918 -1108 978
rect -1048 918 -1042 978
rect -3328 724 -3216 833
rect -2020 814 -2014 874
rect -1954 814 -1948 874
rect -724 866 -664 1088
rect -464 978 -404 1088
rect -470 918 -464 978
rect -404 918 -398 978
rect 216 874 276 2258
rect 344 1664 404 1858
rect 474 1664 534 1764
rect 600 1664 660 2258
rect 344 1604 660 1664
rect 730 1662 790 1764
rect 724 1602 730 1662
rect 790 1602 796 1662
rect 592 1478 598 1538
rect 658 1478 664 1538
rect 342 988 402 1192
rect 474 988 534 1088
rect 598 988 658 1478
rect 856 1292 916 2430
rect 982 2146 988 2206
rect 1048 2146 1054 2206
rect 1238 2146 1244 2206
rect 1304 2146 1310 2206
rect 988 2060 1048 2146
rect 1244 2060 1304 2146
rect 982 1602 988 1662
rect 1048 1602 1054 1662
rect 988 1386 1048 1602
rect 1116 1538 1176 1854
rect 1240 1602 1246 1662
rect 1306 1602 1312 1662
rect 1110 1478 1116 1538
rect 1176 1478 1182 1538
rect 1246 1386 1306 1602
rect 1374 1310 1434 2430
rect 1626 2258 1632 2318
rect 1692 2258 1698 2318
rect 1500 1662 1560 1764
rect 1632 1662 1692 2258
rect 1996 2146 2002 2206
rect 2062 2146 2068 2206
rect 1762 1662 1822 1764
rect 1892 1662 1952 1872
rect 1494 1602 1500 1662
rect 1560 1602 1566 1662
rect 1632 1602 1952 1662
rect 1624 1478 1630 1538
rect 1690 1478 1950 1538
rect 1630 1300 1690 1478
rect 1762 1390 1822 1478
rect 1890 1288 1950 1478
rect 342 928 658 988
rect 728 986 788 1088
rect 722 926 728 986
rect 788 926 794 986
rect 1114 874 1174 1186
rect 1502 986 1562 1088
rect 2002 986 2062 2146
rect 2304 1888 2364 2430
rect 2426 2094 2432 2154
rect 2492 2094 2498 2154
rect 2432 1982 2492 2094
rect 1496 926 1502 986
rect 1562 926 1568 986
rect 1996 926 2002 986
rect 2062 926 2068 986
rect 2432 984 2492 1092
rect 2556 976 2616 1196
rect 2432 918 2492 924
rect 2550 916 2556 976
rect 2616 916 2622 976
rect 210 814 216 874
rect 276 814 282 874
rect 1108 814 1114 874
rect 1174 814 1180 874
rect 3216 833 3222 2907
rect 3322 833 3328 2907
rect -724 800 -664 806
rect 3216 724 3328 833
rect -3328 718 3328 724
rect -3328 618 -3222 718
rect 3222 618 3328 718
rect -3328 612 3328 618
rect -3328 382 3328 388
rect -3328 282 -3222 382
rect 3222 282 3328 382
rect -3328 276 3328 282
rect -3328 97 -3216 276
rect -3328 -3237 -3322 97
rect -3222 -3237 -3216 97
rect -3128 182 -72 188
rect -3128 82 -3022 182
rect -178 82 -72 182
rect -3128 76 -72 82
rect -3128 28 -3016 76
rect -3128 -948 -3122 28
rect -3022 -948 -3016 28
rect -184 28 -72 76
rect -2112 -46 -2106 14
rect -2046 -46 -2040 14
rect -1078 -46 -1072 14
rect -1012 -46 -1006 14
rect -2628 -162 -2622 -102
rect -2562 -162 -2556 -102
rect -2622 -220 -2562 -162
rect -2876 -280 -2562 -220
rect -2496 -280 -2490 -220
rect -2430 -280 -2424 -220
rect -2876 -462 -2816 -280
rect -2750 -382 -2690 -280
rect -2622 -486 -2562 -280
rect -2490 -386 -2430 -280
rect -2106 -474 -2046 -46
rect -1592 -162 -1586 -102
rect -1526 -162 -1520 -102
rect -1720 -280 -1714 -220
rect -1654 -280 -1648 -220
rect -1714 -382 -1654 -280
rect -1586 -474 -1526 -162
rect -1466 -280 -1460 -220
rect -1400 -280 -1394 -220
rect -1460 -386 -1400 -280
rect -1072 -472 -1012 -46
rect -562 -162 -556 -102
rect -496 -162 -490 -102
rect -556 -220 -496 -162
rect -686 -280 -680 -220
rect -620 -280 -614 -220
rect -556 -280 -236 -220
rect -680 -386 -620 -280
rect -556 -480 -496 -280
rect -426 -382 -366 -280
rect -296 -480 -236 -280
rect -2362 -874 -2302 -580
rect -2230 -756 -2170 -658
rect -1974 -756 -1914 -660
rect -2236 -816 -2230 -756
rect -2170 -816 -2164 -756
rect -1980 -816 -1974 -756
rect -1914 -816 -1908 -756
rect -1846 -874 -1786 -570
rect -1326 -874 -1266 -580
rect -1200 -756 -1140 -656
rect -942 -756 -882 -656
rect -1206 -816 -1200 -756
rect -1140 -816 -1134 -756
rect -948 -816 -942 -756
rect -882 -816 -876 -756
rect -814 -874 -754 -576
rect -2368 -934 -2362 -874
rect -2302 -934 -2296 -874
rect -1852 -934 -1846 -874
rect -1786 -934 -1780 -874
rect -1332 -934 -1326 -874
rect -1266 -934 -1260 -874
rect -820 -934 -814 -874
rect -754 -934 -748 -874
rect -3128 -996 -3016 -948
rect -184 -948 -178 28
rect -78 -948 -72 28
rect 3216 97 3328 276
rect 1114 -66 1174 -60
rect 2426 -124 2432 -64
rect 2492 -124 2498 -64
rect 2556 -72 2616 -66
rect 1114 -182 1174 -126
rect 726 -242 1560 -182
rect 726 -346 786 -242
rect 988 -344 1048 -242
rect 344 -702 404 -542
rect 470 -702 530 -620
rect 596 -702 656 -524
rect 344 -762 596 -702
rect 656 -762 662 -702
rect -184 -996 -72 -948
rect -3128 -1002 -72 -996
rect -3128 -1102 -3022 -1002
rect -178 -1102 -72 -1002
rect -3128 -1108 -72 -1102
rect 854 -850 914 -526
rect 1114 -558 1174 -242
rect 1242 -346 1302 -242
rect 1500 -346 1560 -242
rect 2432 -322 2492 -124
rect 2556 -422 2616 -132
rect 1370 -850 1430 -526
rect 1630 -702 1690 -530
rect 1760 -702 1820 -622
rect 1888 -702 1948 -546
rect 1624 -762 1630 -702
rect 1690 -762 1948 -702
rect 2296 -850 2356 -690
rect 854 -910 2356 -850
rect 2432 -888 2492 -796
rect 854 -1212 914 -910
rect 2296 -1212 2356 -910
rect 2426 -948 2432 -888
rect 2492 -948 2498 -888
rect -3128 -1218 3128 -1212
rect -3128 -1318 -3022 -1218
rect 3022 -1318 3128 -1218
rect -3128 -1324 3128 -1318
rect -3128 -1384 -3016 -1324
rect -3128 -2576 -3122 -1384
rect -3022 -2576 -3016 -1384
rect -2728 -1468 -2722 -1408
rect -2662 -1468 -2656 -1408
rect -2722 -2356 -2662 -1468
rect -2576 -1489 -1660 -1429
rect -1302 -1468 -1296 -1408
rect -1236 -1468 -1230 -1408
rect -434 -1468 -428 -1408
rect -368 -1468 -362 -1408
rect -8 -1468 -2 -1408
rect 58 -1468 64 -1408
rect 418 -1468 424 -1408
rect 484 -1468 490 -1408
rect -2576 -1672 -2516 -1489
rect -2138 -1576 -2078 -1489
rect -1720 -1676 -1660 -1489
rect -1296 -1588 -1236 -1468
rect -428 -1582 -368 -1468
rect -2 -1674 58 -1468
rect 424 -1586 484 -1468
rect 854 -1680 914 -1324
rect 3016 -1384 3128 -1324
rect 1290 -1468 1296 -1408
rect 1356 -1468 1362 -1408
rect 1296 -1582 1356 -1468
rect 1712 -1489 2768 -1429
rect 1712 -1660 1772 -1489
rect 2132 -1576 2192 -1489
rect 2568 -1694 2628 -1489
rect -2582 -1892 -2522 -1742
rect -2588 -1952 -2582 -1892
rect -2522 -1952 -2516 -1892
rect -1286 -1998 -1226 -1851
rect -2576 -2356 -2516 -2160
rect -2138 -2356 -2078 -2269
rect -1720 -2356 -1660 -2166
rect -2722 -2416 -1660 -2356
rect -860 -2372 -800 -1765
rect -424 -1998 -364 -1851
rect 432 -1998 492 -1851
rect 852 -2088 912 -1761
rect 1284 -2002 1344 -1855
rect 2562 -1958 2568 -1898
rect 2628 -1958 2634 -1898
rect -866 -2432 -860 -2372
rect -800 -2432 -794 -2372
rect -3128 -2636 -3016 -2576
rect -860 -2636 -800 -2432
rect -2 -2486 58 -2178
rect 850 -2372 910 -2162
rect 1712 -2356 1772 -2160
rect 2150 -2356 2210 -2269
rect 2568 -2356 2628 -1958
rect 844 -2432 850 -2372
rect 910 -2432 916 -2372
rect 1712 -2416 2628 -2356
rect -8 -2546 -2 -2486
rect 58 -2546 64 -2486
rect 850 -2636 910 -2432
rect 2708 -2486 2768 -1489
rect 2702 -2546 2708 -2486
rect 2768 -2546 2774 -2486
rect 3016 -2576 3022 -1384
rect 3122 -2576 3128 -1384
rect 3016 -2636 3128 -2576
rect -3128 -2642 3128 -2636
rect -3128 -2742 -3022 -2642
rect 3022 -2742 3128 -2642
rect -3128 -2748 3128 -2742
rect -860 -2836 -800 -2748
rect 850 -2836 910 -2748
rect -928 -2864 970 -2836
rect -928 -2974 -898 -2864
rect 942 -2974 970 -2864
rect -928 -3002 970 -2974
rect -3328 -3416 -3216 -3237
rect -2616 -3416 -2606 -3116
rect 2606 -3416 2616 -3116
rect 3216 -3237 3222 97
rect 3322 -3237 3328 97
rect 3216 -3416 3328 -3237
rect -3328 -3422 3328 -3416
rect -3328 -3522 -3222 -3422
rect 3222 -3522 3328 -3422
rect -3328 -3528 3328 -3522
<< via1 >>
rect -3216 2716 -2616 3016
rect 2616 2716 3216 3016
rect -2646 2456 2544 2528
rect -2776 2146 -2716 2206
rect -2266 2146 -2206 2206
rect -2270 1604 -2210 1664
rect -2138 1470 -2078 1530
rect -2008 1470 -1948 1530
rect -1622 2146 -1562 2206
rect -1496 2146 -1436 2206
rect -1494 1604 -1434 1664
rect -1750 1470 -1690 1530
rect -1628 1470 -1568 1530
rect -1232 2146 -1172 2206
rect -1240 1604 -1180 1664
rect -1112 1470 -1052 1530
rect -980 1470 -920 1530
rect -596 2146 -536 2206
rect -464 2146 -404 2206
rect -464 1604 -404 1664
rect -720 1470 -660 1530
rect -596 1470 -536 1530
rect 216 2258 276 2318
rect 600 2258 660 2318
rect -2776 918 -2716 978
rect -2274 918 -2214 978
rect -2142 918 -2082 978
rect -1500 918 -1440 978
rect -1240 918 -1180 978
rect -1108 918 -1048 978
rect -2014 814 -1954 874
rect -464 918 -404 978
rect 730 1602 790 1662
rect 598 1478 658 1538
rect 988 2146 1048 2206
rect 1244 2146 1304 2206
rect 988 1602 1048 1662
rect 1246 1602 1306 1662
rect 1116 1478 1176 1538
rect 1632 2258 1692 2318
rect 2002 2146 2062 2206
rect 1500 1602 1560 1662
rect 1630 1478 1690 1538
rect 728 926 788 986
rect 2432 2094 2492 2154
rect 1502 926 1562 986
rect 2002 926 2062 986
rect 2432 924 2492 984
rect 2556 916 2616 976
rect -724 806 -664 866
rect 216 814 276 874
rect 1114 814 1174 874
rect -2106 -46 -2046 14
rect -1072 -46 -1012 14
rect -2622 -162 -2562 -102
rect -2490 -280 -2430 -220
rect -1586 -162 -1526 -102
rect -1714 -280 -1654 -220
rect -1460 -280 -1400 -220
rect -556 -162 -496 -102
rect -680 -280 -620 -220
rect -2230 -816 -2170 -756
rect -1974 -816 -1914 -756
rect -1200 -816 -1140 -756
rect -942 -816 -882 -756
rect -2362 -934 -2302 -874
rect -1846 -934 -1786 -874
rect -1326 -934 -1266 -874
rect -814 -934 -754 -874
rect 1114 -126 1174 -66
rect 2432 -124 2492 -64
rect 596 -762 656 -702
rect 2556 -132 2616 -72
rect 1630 -762 1690 -702
rect 2432 -948 2492 -888
rect -2722 -1468 -2662 -1408
rect -1296 -1468 -1236 -1408
rect -428 -1468 -368 -1408
rect -2 -1468 58 -1408
rect 424 -1468 484 -1408
rect 1296 -1468 1356 -1408
rect -2582 -1952 -2522 -1892
rect 2568 -1958 2628 -1898
rect -860 -2432 -800 -2372
rect 850 -2432 910 -2372
rect -2 -2546 58 -2486
rect 2708 -2546 2768 -2486
rect -898 -2974 942 -2864
rect -3216 -3416 -2616 -3116
rect 2616 -3416 3216 -3116
<< metal2 >>
rect -3216 3016 -2616 3026
rect -3216 2706 -2616 2716
rect 2616 3016 3216 3026
rect 2616 2706 3216 2716
rect -2674 2528 2566 2562
rect -2674 2456 -2646 2528
rect 2544 2456 2566 2528
rect -2674 2430 2566 2456
rect 216 2318 276 2324
rect 600 2318 660 2324
rect 1632 2318 1692 2324
rect 276 2258 600 2318
rect 660 2258 1632 2318
rect 216 2252 276 2258
rect 600 2252 660 2258
rect 1632 2252 1692 2258
rect -2776 2206 -2716 2212
rect -2266 2206 -2206 2212
rect -1622 2206 -1562 2212
rect -1496 2206 -1436 2212
rect -1232 2206 -1172 2212
rect -596 2206 -536 2212
rect -464 2206 -404 2212
rect 988 2206 1048 2212
rect 1244 2206 1304 2212
rect 2002 2206 2062 2212
rect -2716 2146 -2266 2206
rect -2206 2146 -1622 2206
rect -1562 2146 -1496 2206
rect -1436 2146 -1232 2206
rect -1172 2146 -596 2206
rect -536 2146 -464 2206
rect -404 2146 988 2206
rect 1048 2146 1244 2206
rect 1304 2146 2002 2206
rect 2432 2154 2492 2160
rect -2776 2140 -2716 2146
rect -2266 2140 -2206 2146
rect -1622 2140 -1562 2146
rect -1496 2140 -1436 2146
rect -1232 2140 -1172 2146
rect -596 2140 -536 2146
rect -464 2140 -404 2146
rect 988 2140 1048 2146
rect 1244 2140 1304 2146
rect 2002 2140 2062 2146
rect 2132 2094 2432 2154
rect -2270 1664 -2210 1670
rect -1494 1664 -1434 1670
rect -1240 1664 -1180 1670
rect -464 1664 -404 1670
rect -2210 1604 -1494 1664
rect -1434 1604 -1240 1664
rect -1180 1604 -464 1664
rect 730 1662 790 1668
rect 988 1662 1048 1668
rect 1246 1662 1306 1668
rect 1500 1662 1560 1668
rect -2270 1598 -2210 1604
rect -1494 1598 -1434 1604
rect -1240 1598 -1180 1604
rect -464 1598 -404 1604
rect 72 1602 730 1662
rect 790 1602 988 1662
rect 1048 1602 1246 1662
rect 1306 1602 1500 1662
rect -2138 1530 -2078 1536
rect -2008 1530 -1948 1536
rect -1750 1530 -1690 1536
rect -1628 1530 -1568 1536
rect -1112 1530 -1052 1536
rect -980 1530 -920 1536
rect -720 1530 -660 1536
rect -596 1530 -536 1536
rect 72 1530 132 1602
rect 730 1596 790 1602
rect 988 1596 1048 1602
rect 1246 1596 1306 1602
rect 1500 1596 1560 1602
rect -2078 1470 -2008 1530
rect -1948 1470 -1750 1530
rect -1690 1470 -1628 1530
rect -1568 1470 -1112 1530
rect -1052 1470 -980 1530
rect -920 1470 -720 1530
rect -660 1470 -596 1530
rect -536 1470 132 1530
rect 598 1538 658 1544
rect 1116 1538 1176 1544
rect 1630 1538 1690 1544
rect 2132 1538 2192 2094
rect 2432 2088 2492 2094
rect 658 1478 1116 1538
rect 1176 1478 1630 1538
rect 1690 1478 2192 1538
rect 598 1472 658 1478
rect 1116 1472 1176 1478
rect 1630 1472 1690 1478
rect -2138 1464 -2078 1470
rect -2008 1464 -1948 1470
rect -1750 1464 -1690 1470
rect -1628 1464 -1568 1470
rect -1112 1464 -1052 1470
rect -980 1464 -920 1470
rect -720 1464 -660 1470
rect -596 1464 -536 1470
rect 728 986 788 992
rect 1502 986 1562 992
rect 2002 986 2062 992
rect -2776 978 -2716 984
rect -2274 978 -2214 984
rect -2142 978 -2082 984
rect -1500 978 -1440 984
rect -1240 978 -1180 984
rect -1108 978 -1048 984
rect -464 978 -404 984
rect -2716 918 -2274 978
rect -2214 918 -2142 978
rect -2082 918 -1500 978
rect -1440 918 -1240 978
rect -1180 918 -1108 978
rect -1048 918 -464 978
rect 788 926 1502 986
rect 1562 926 2002 986
rect 728 920 788 926
rect 1502 920 1562 926
rect 2002 920 2062 926
rect -2776 912 -2716 918
rect -2274 912 -2214 918
rect -2142 912 -2082 918
rect -2014 874 -1954 880
rect -2014 534 -1954 814
rect -2234 474 -1954 534
rect -2622 -102 -2562 -96
rect -2234 -102 -2174 474
rect -2106 14 -2046 20
rect -1748 14 -1688 918
rect -1500 912 -1440 918
rect -1370 14 -1310 918
rect -1240 912 -1180 918
rect -1108 912 -1048 918
rect -464 912 -404 918
rect 216 874 276 880
rect 1114 874 1174 880
rect -730 806 -724 866
rect -664 806 -658 866
rect 276 814 1114 874
rect 216 808 276 814
rect -1072 14 -1012 20
rect -2046 -46 -1072 14
rect -2106 -52 -2046 -46
rect -1072 -52 -1012 -46
rect -1586 -102 -1526 -96
rect -724 -102 -664 806
rect 1114 -66 1174 814
rect 2132 254 2192 1478
rect 2426 924 2432 984
rect 2492 924 2498 984
rect 2556 976 2616 982
rect 2432 254 2492 924
rect 2132 194 2492 254
rect -556 -102 -496 -96
rect -2562 -162 -1586 -102
rect -1526 -162 -556 -102
rect 1108 -126 1114 -66
rect 1174 -126 1180 -66
rect -2622 -168 -2562 -162
rect -1586 -168 -1526 -162
rect -556 -168 -496 -162
rect -2490 -220 -2430 -214
rect -1714 -220 -1654 -214
rect -1460 -220 -1400 -214
rect -680 -220 -620 -214
rect -2430 -280 -1714 -220
rect -1654 -280 -1460 -220
rect -1400 -280 -680 -220
rect -2490 -286 -2430 -280
rect -1714 -286 -1654 -280
rect -1460 -286 -1400 -280
rect -680 -286 -620 -280
rect 596 -702 656 -696
rect 1630 -702 1690 -696
rect 2132 -702 2192 194
rect 2432 -64 2492 194
rect 2556 -72 2616 916
rect 2432 -130 2492 -124
rect 2550 -132 2556 -72
rect 2616 -132 2622 -72
rect -2230 -756 -2170 -750
rect -1974 -756 -1914 -750
rect -1200 -756 -1140 -750
rect -942 -756 -882 -750
rect -2170 -816 -1974 -756
rect -1914 -816 -1200 -756
rect -1140 -816 -942 -756
rect 656 -762 1630 -702
rect 1690 -762 2192 -702
rect 596 -768 656 -762
rect 1630 -768 1690 -762
rect -2230 -822 -2170 -816
rect -1974 -822 -1914 -816
rect -1200 -822 -1140 -816
rect -942 -822 -882 -816
rect -2362 -874 -2302 -868
rect -1846 -874 -1786 -868
rect -1326 -874 -1266 -868
rect -814 -874 -754 -868
rect -2852 -934 -2362 -874
rect -2302 -934 -1846 -874
rect -1786 -934 -1326 -874
rect -1266 -934 -814 -874
rect -2852 -1892 -2792 -934
rect -2362 -940 -2302 -934
rect -1846 -940 -1786 -934
rect -1326 -940 -1266 -934
rect -814 -940 -754 -934
rect 2132 -888 2192 -762
rect 2432 -888 2492 -882
rect 2132 -948 2432 -888
rect 2432 -954 2492 -948
rect -2722 -1408 -2662 -1402
rect -1296 -1408 -1236 -1402
rect -428 -1408 -368 -1402
rect -2 -1408 58 -1402
rect 424 -1408 484 -1402
rect 1296 -1408 1356 -1402
rect -2662 -1468 -1296 -1408
rect -1236 -1468 -428 -1408
rect -368 -1468 -2 -1408
rect 58 -1468 424 -1408
rect 484 -1468 1296 -1408
rect 1356 -1468 2908 -1408
rect -2722 -1474 -2662 -1468
rect -1296 -1474 -1236 -1468
rect -428 -1474 -368 -1468
rect -2 -1474 58 -1468
rect 424 -1474 484 -1468
rect 1296 -1474 1356 -1468
rect -2582 -1892 -2522 -1886
rect -2852 -1952 -2582 -1892
rect -2852 -2486 -2792 -1952
rect -2582 -1958 -2522 -1952
rect 2568 -1898 2628 -1892
rect 2848 -1898 2908 -1468
rect 2628 -1958 2908 -1898
rect 2568 -1964 2628 -1958
rect -860 -2372 -800 -2366
rect 850 -2372 910 -2366
rect -800 -2432 850 -2372
rect -860 -2438 -800 -2432
rect 850 -2438 910 -2432
rect -2 -2486 58 -2480
rect 2708 -2486 2768 -2480
rect -2852 -2546 -2 -2486
rect 58 -2546 2708 -2486
rect -2 -2552 58 -2546
rect 2708 -2552 2768 -2546
rect -928 -2864 970 -2836
rect -928 -2974 -898 -2864
rect 942 -2974 970 -2864
rect -928 -3002 970 -2974
rect -3216 -3116 -2616 -3106
rect -3216 -3426 -2616 -3416
rect 2616 -3116 3216 -3106
rect 2616 -3426 3216 -3416
<< via2 >>
rect -3216 2716 -2616 3016
rect 2616 2716 3216 3016
rect -2646 2456 2544 2528
rect -898 -2974 942 -2864
rect -3216 -3416 -2616 -3116
rect 2616 -3416 3216 -3116
<< metal3 >>
rect -3226 3016 -2606 3021
rect -3226 2716 -3216 3016
rect -2616 2716 -2606 3016
rect -3226 2711 -2606 2716
rect 2606 3016 3226 3021
rect 2606 2716 2616 3016
rect 3216 2716 3226 3016
rect 2606 2711 3226 2716
rect -2674 2528 2566 2562
rect -2674 2456 -2646 2528
rect 2544 2456 2566 2528
rect -2674 2430 2566 2456
rect -928 -2864 970 -2836
rect -928 -2974 -898 -2864
rect 942 -2974 970 -2864
rect -928 -3002 970 -2974
rect -3226 -3116 -2606 -3111
rect -3226 -3416 -3216 -3116
rect -2616 -3416 -2606 -3116
rect -3226 -3421 -2606 -3416
rect 2606 -3116 3226 -3111
rect 2606 -3416 2616 -3116
rect 3216 -3416 3226 -3116
rect 2606 -3421 3226 -3416
<< via3 >>
rect -3216 2716 -2616 3016
rect 2616 2716 3216 3016
rect -2646 2456 2544 2528
rect -898 -2974 942 -2864
rect -3216 -3416 -2616 -3116
rect 2616 -3416 3216 -3116
<< metal4 >>
rect -3400 3016 3400 3200
rect -3400 2716 -3216 3016
rect -2616 2716 2616 3016
rect 3216 2716 3400 3016
rect -3400 2528 3400 2716
rect -3400 2456 -2646 2528
rect 2544 2456 3400 2528
rect -3400 2400 3400 2456
rect -3400 -2864 3400 -2800
rect -3400 -2974 -898 -2864
rect 942 -2974 3400 -2864
rect -3400 -3116 3400 -2974
rect -3400 -3416 -3216 -3116
rect -2616 -3416 2616 -3116
rect 3216 -3416 3400 -3116
rect -3400 -3600 3400 -3416
use sky130_fd_pr__nfet_01v8_lvt_G98Z6N  sky130_fd_pr__nfet_01v8_lvt_G98Z6N_0
timestamp 1624477805
transform 1 0 -1557 0 1 -522
box -1319 -188 1319 188
use sky130_fd_pr__nfet_01v8_JP3XZJ  sky130_fd_pr__nfet_01v8_JP3XZJ_0
timestamp 1624477805
transform 1 0 28 0 1 -1924
box -2603 -397 2603 397
use sky130_fd_pr__nfet_01v8_V7Q58M  sky130_fd_pr__nfet_01v8_V7Q58M_0
timestamp 1624477805
transform 1 0 2462 0 1 -558
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_8B5GXQ  sky130_fd_pr__nfet_01v8_8B5GXQ_0
timestamp 1624477805
transform 1 0 1145 0 1 -484
box -803 -188 803 188
use sky130_fd_pr__pfet_01v8_H2H4BB  sky130_fd_pr__pfet_01v8_H2H4BB_1
timestamp 1624477805
transform 1 0 -1336 0 1 1239
box -1355 -200 1355 200
use sky130_fd_pr__pfet_01v8_H2H4BB  sky130_fd_pr__pfet_01v8_H2H4BB_0
timestamp 1624477805
transform 1 0 -1336 0 1 1913
box -1355 -200 1355 200
use sky130_fd_pr__pfet_01v8_hvt_ATGTW6  sky130_fd_pr__pfet_01v8_hvt_ATGTW6_0
timestamp 1624477805
transform 1 0 2462 0 1 1538
box -194 -500 194 500
use sky130_fd_pr__pfet_01v8_RC2RSP  sky130_fd_pr__pfet_01v8_RC2RSP_0
timestamp 1624477805
transform 1 0 1147 0 1 1912
box -839 -200 839 200
use sky130_fd_pr__pfet_01v8_RC2RSP  sky130_fd_pr__pfet_01v8_RC2RSP_1
timestamp 1624477805
transform 1 0 1147 0 1 1238
box -839 -200 839 200
<< labels >>
flabel metal1 886 -216 900 -202 1 FreeSans 480 0 0 0 vmirror
flabel metal1 436 -744 448 -730 1 FreeSans 480 0 0 0 vo1
flabel metal1 2726 -2168 2748 -2144 1 FreeSans 480 0 0 0 vtail
flabel metal2 -820 -1444 -780 -1426 1 FreeSans 480 0 0 0 ibiasn
flabel metal2 -452 -2416 -440 -2394 1 FreeSans 480 0 0 0 VSS
flabel metal1 -2766 -264 -2732 -234 1 FreeSans 480 0 0 0 vcompm
flabel metal2 -2292 -262 -2260 -238 1 FreeSans 480 0 0 0 vip
flabel metal2 -1592 -802 -1560 -774 1 FreeSans 480 0 0 0 vim
flabel metal2 -1592 -914 -1566 -890 1 FreeSans 480 0 0 0 vtail
flabel metal2 -1654 -28 -1634 -4 1 FreeSans 480 0 0 0 vcompp
flabel metal1 2026 1582 2042 1600 1 FreeSans 480 0 0 0 vcompp
flabel metal1 1522 1686 1534 1696 1 FreeSans 480 0 0 0 vcompm
flabel metal2 1500 1502 1516 1514 1 FreeSans 480 0 0 0 vo1
flabel metal2 824 832 836 848 1 FreeSans 480 0 0 0 vmirror
flabel metal1 -2122 1544 -2104 1566 1 FreeSans 480 0 0 0 vcompm
flabel metal2 2586 472 2596 480 1 FreeSans 480 0 0 0 vo
flabel metal2 -720 2168 -702 2188 1 FreeSans 480 0 0 0 vcompp
flabel metal4 -1674 2724 -1612 2786 1 FreeSans 480 0 0 0 VDD
<< properties >>
string FIXED_BBOX -3272 -3472 3272 332
<< end >>
