magic
tech sky130A
magscale 1 2
timestamp 1624234649
<< nwell >>
rect 11292 17622 35808 28298
rect 47228 24930 49137 25448
rect 47228 24609 49462 24930
rect 47228 24608 49137 24609
rect 47228 22930 49137 23448
rect 47228 22609 49462 22930
rect 47228 22608 49137 22609
rect 65292 17622 89808 28298
rect -13130 15800 -8621 16318
rect -13130 15479 -7796 15800
rect -13130 15478 -8621 15479
rect 48654 7966 50563 8484
rect 48654 7645 50888 7966
rect 48654 7644 50563 7645
rect 48654 6002 50563 6520
rect 48654 5681 50888 6002
rect 48654 5680 50563 5681
rect 48654 4002 50563 4520
rect 48654 3681 50888 4002
rect 48654 3680 50563 3681
rect 48654 1912 50563 2430
rect 48654 1591 50888 1912
rect 48654 1590 50563 1591
<< pwell >>
rect 49086 24550 49116 24552
rect 49086 24514 49137 24550
rect 47228 23894 49137 24514
rect 49196 24369 49382 24551
rect 49361 24365 49382 24369
rect 49361 24331 49395 24365
rect 49086 22550 49116 22552
rect 49086 22514 49137 22550
rect 47228 21894 49137 22514
rect 49196 22369 49382 22551
rect 49361 22365 49382 22369
rect 49361 22331 49395 22365
rect -11272 15420 -11242 15422
rect -11272 15384 -11221 15420
rect -11162 15384 -10976 15421
rect -8672 15420 -8642 15422
rect -8672 15384 -8621 15420
rect -13130 14764 -8621 15384
rect -8562 15406 -8084 15421
rect -8062 15406 -7876 15421
rect -8562 15239 -7876 15406
rect -8397 15235 -8376 15239
rect -7897 15235 -7876 15239
rect -8397 15201 -8363 15235
rect -7897 15201 -7863 15235
rect -1408 -718 35908 15398
rect 50512 7586 50542 7588
rect 50512 7550 50563 7586
rect 48654 6930 50563 7550
rect 50622 7405 50808 7587
rect 50787 7401 50808 7405
rect 50787 7367 50821 7401
rect 50512 5622 50542 5624
rect 50512 5586 50563 5622
rect 48654 4966 50563 5586
rect 50622 5441 50808 5623
rect 50787 5437 50808 5441
rect 50787 5403 50821 5437
rect 50512 3622 50542 3624
rect 50512 3586 50563 3622
rect 48654 2966 50563 3586
rect 50622 3441 50808 3623
rect 50787 3437 50808 3441
rect 50787 3403 50821 3437
rect 50512 1532 50542 1534
rect 50512 1496 50563 1532
rect 48654 876 50563 1496
rect 50622 1351 50808 1533
rect 50787 1347 50808 1351
rect 50787 1313 50821 1347
rect 52592 -718 89908 15398
<< nmos >>
rect 47424 24104 47624 24304
rect 47682 24104 47882 24304
rect 47940 24104 48140 24304
rect 48198 24104 48398 24304
rect 48456 24104 48656 24304
rect 48714 24104 48914 24304
rect 47424 22104 47624 22304
rect 47682 22104 47882 22304
rect 47940 22104 48140 22304
rect 48198 22104 48398 22304
rect 48456 22104 48656 22304
rect 48714 22104 48914 22304
rect -12934 14974 -12734 15174
rect -12676 14974 -12476 15174
rect -12418 14974 -12218 15174
rect -12160 14974 -11960 15174
rect -11902 14974 -11702 15174
rect -11644 14974 -11444 15174
rect -10334 14974 -10134 15174
rect -10076 14974 -9876 15174
rect -9818 14974 -9618 15174
rect -9560 14974 -9360 15174
rect -9302 14974 -9102 15174
rect -9044 14974 -8844 15174
rect 13578 14222 14538 14822
rect 14596 14222 15556 14822
rect 15614 14222 16574 14822
rect 16632 14222 17592 14822
rect 17650 14222 18610 14822
rect 18668 14222 19628 14822
rect 19686 14222 20646 14822
rect 20704 14222 21664 14822
rect 21722 14222 22682 14822
rect 22740 14222 23700 14822
rect 23758 14222 24718 14822
rect 24776 14222 25736 14822
rect 25794 14222 26754 14822
rect 26812 14222 27772 14822
rect 27830 14222 28790 14822
rect 28848 14222 29808 14822
rect 29866 14222 30826 14822
rect 30884 14222 31844 14822
rect 31902 14222 32862 14822
rect 32920 14222 33880 14822
rect 13578 12988 14538 13588
rect 14596 12988 15556 13588
rect 15614 12988 16574 13588
rect 16632 12988 17592 13588
rect 17650 12988 18610 13588
rect 18668 12988 19628 13588
rect 19686 12988 20646 13588
rect 20704 12988 21664 13588
rect 21722 12988 22682 13588
rect 22740 12988 23700 13588
rect 23758 12988 24718 13588
rect 24776 12988 25736 13588
rect 25794 12988 26754 13588
rect 26812 12988 27772 13588
rect 27830 12988 28790 13588
rect 28848 12988 29808 13588
rect 29866 12988 30826 13588
rect 30884 12988 31844 13588
rect 31902 12988 32862 13588
rect 32920 12988 33880 13588
rect 13578 11756 14538 12356
rect 14596 11756 15556 12356
rect 15614 11756 16574 12356
rect 16632 11756 17592 12356
rect 17650 11756 18610 12356
rect 18668 11756 19628 12356
rect 19686 11756 20646 12356
rect 20704 11756 21664 12356
rect 21722 11756 22682 12356
rect 22740 11756 23700 12356
rect 23758 11756 24718 12356
rect 24776 11756 25736 12356
rect 25794 11756 26754 12356
rect 26812 11756 27772 12356
rect 27830 11756 28790 12356
rect 28848 11756 29808 12356
rect 29866 11756 30826 12356
rect 30884 11756 31844 12356
rect 31902 11756 32862 12356
rect 32920 11756 33880 12356
rect 13576 10522 14536 11122
rect 14594 10522 15554 11122
rect 15612 10522 16572 11122
rect 16630 10522 17590 11122
rect 17648 10522 18608 11122
rect 18666 10522 19626 11122
rect 19684 10522 20644 11122
rect 20702 10522 21662 11122
rect 21720 10522 22680 11122
rect 22738 10522 23698 11122
rect 23756 10522 24716 11122
rect 24774 10522 25734 11122
rect 25792 10522 26752 11122
rect 26810 10522 27770 11122
rect 27828 10522 28788 11122
rect 28846 10522 29806 11122
rect 29864 10522 30824 11122
rect 30882 10522 31842 11122
rect 31900 10522 32860 11122
rect 32918 10522 33878 11122
rect 13576 9288 14536 9888
rect 14594 9288 15554 9888
rect 15612 9288 16572 9888
rect 16630 9288 17590 9888
rect 17648 9288 18608 9888
rect 18666 9288 19626 9888
rect 19684 9288 20644 9888
rect 20702 9288 21662 9888
rect 21720 9288 22680 9888
rect 22738 9288 23698 9888
rect 23756 9288 24716 9888
rect 24774 9288 25734 9888
rect 25792 9288 26752 9888
rect 26810 9288 27770 9888
rect 27828 9288 28788 9888
rect 28846 9288 29806 9888
rect 29864 9288 30824 9888
rect 30882 9288 31842 9888
rect 31900 9288 32860 9888
rect 32918 9288 33878 9888
rect 13576 8056 14536 8656
rect 14594 8056 15554 8656
rect 15612 8056 16572 8656
rect 16630 8056 17590 8656
rect 17648 8056 18608 8656
rect 18666 8056 19626 8656
rect 19684 8056 20644 8656
rect 20702 8056 21662 8656
rect 21720 8056 22680 8656
rect 22738 8056 23698 8656
rect 23756 8056 24716 8656
rect 24774 8056 25734 8656
rect 25792 8056 26752 8656
rect 26810 8056 27770 8656
rect 27828 8056 28788 8656
rect 28846 8056 29806 8656
rect 29864 8056 30824 8656
rect 30882 8056 31842 8656
rect 31900 8056 32860 8656
rect 32918 8056 33878 8656
rect 13576 6822 14536 7422
rect 14594 6822 15554 7422
rect 15612 6822 16572 7422
rect 16630 6822 17590 7422
rect 17648 6822 18608 7422
rect 18666 6822 19626 7422
rect 19684 6822 20644 7422
rect 20702 6822 21662 7422
rect 21720 6822 22680 7422
rect 22738 6822 23698 7422
rect 23756 6822 24716 7422
rect 24774 6822 25734 7422
rect 25792 6822 26752 7422
rect 26810 6822 27770 7422
rect 27828 6822 28788 7422
rect 28846 6822 29806 7422
rect 29864 6822 30824 7422
rect 30882 6822 31842 7422
rect 31900 6822 32860 7422
rect 32918 6822 33878 7422
rect 13576 5588 14536 6188
rect 14594 5588 15554 6188
rect 15612 5588 16572 6188
rect 16630 5588 17590 6188
rect 17648 5588 18608 6188
rect 18666 5588 19626 6188
rect 19684 5588 20644 6188
rect 20702 5588 21662 6188
rect 21720 5588 22680 6188
rect 22738 5588 23698 6188
rect 23756 5588 24716 6188
rect 24774 5588 25734 6188
rect 25792 5588 26752 6188
rect 26810 5588 27770 6188
rect 27828 5588 28788 6188
rect 28846 5588 29806 6188
rect 29864 5588 30824 6188
rect 30882 5588 31842 6188
rect 31900 5588 32860 6188
rect 32918 5588 33878 6188
rect 1591 4159 2551 4759
rect 2609 4159 3569 4759
rect 3627 4159 4587 4759
rect 4645 4159 5605 4759
rect 5663 4159 6623 4759
rect 6681 4159 7641 4759
rect 13576 4356 14536 4956
rect 14594 4356 15554 4956
rect 15612 4356 16572 4956
rect 16630 4356 17590 4956
rect 17648 4356 18608 4956
rect 18666 4356 19626 4956
rect 19684 4356 20644 4956
rect 20702 4356 21662 4956
rect 21720 4356 22680 4956
rect 22738 4356 23698 4956
rect 23756 4356 24716 4956
rect 24774 4356 25734 4956
rect 25792 4356 26752 4956
rect 26810 4356 27770 4956
rect 27828 4356 28788 4956
rect 28846 4356 29806 4956
rect 29864 4356 30824 4956
rect 30882 4356 31842 4956
rect 31900 4356 32860 4956
rect 32918 4356 33878 4956
rect 1590 3046 2550 3646
rect 2608 3046 3568 3646
rect 3626 3046 4586 3646
rect 4644 3046 5604 3646
rect 5662 3046 6622 3646
rect 6680 3046 7640 3646
rect 13576 3122 14536 3722
rect 14594 3122 15554 3722
rect 15612 3122 16572 3722
rect 16630 3122 17590 3722
rect 17648 3122 18608 3722
rect 18666 3122 19626 3722
rect 19684 3122 20644 3722
rect 20702 3122 21662 3722
rect 21720 3122 22680 3722
rect 22738 3122 23698 3722
rect 23756 3122 24716 3722
rect 24774 3122 25734 3722
rect 25792 3122 26752 3722
rect 26810 3122 27770 3722
rect 27828 3122 28788 3722
rect 28846 3122 29806 3722
rect 29864 3122 30824 3722
rect 30882 3122 31842 3722
rect 31900 3122 32860 3722
rect 32918 3122 33878 3722
rect 1591 1935 2551 2535
rect 2609 1935 3569 2535
rect 3627 1935 4587 2535
rect 4645 1935 5605 2535
rect 5663 1935 6623 2535
rect 6681 1935 7641 2535
rect 13576 1888 14536 2488
rect 14594 1888 15554 2488
rect 15612 1888 16572 2488
rect 16630 1888 17590 2488
rect 17648 1888 18608 2488
rect 18666 1888 19626 2488
rect 19684 1888 20644 2488
rect 20702 1888 21662 2488
rect 21720 1888 22680 2488
rect 22738 1888 23698 2488
rect 23756 1888 24716 2488
rect 24774 1888 25734 2488
rect 25792 1888 26752 2488
rect 26810 1888 27770 2488
rect 27828 1888 28788 2488
rect 28846 1888 29806 2488
rect 29864 1888 30824 2488
rect 30882 1888 31842 2488
rect 31900 1888 32860 2488
rect 32918 1888 33878 2488
rect 1590 822 2550 1422
rect 2608 822 3568 1422
rect 3626 822 4586 1422
rect 4644 822 5604 1422
rect 5662 822 6622 1422
rect 6680 822 7640 1422
rect 13576 656 14536 1256
rect 14594 656 15554 1256
rect 15612 656 16572 1256
rect 16630 656 17590 1256
rect 17648 656 18608 1256
rect 18666 656 19626 1256
rect 19684 656 20644 1256
rect 20702 656 21662 1256
rect 21720 656 22680 1256
rect 22738 656 23698 1256
rect 23756 656 24716 1256
rect 24774 656 25734 1256
rect 25792 656 26752 1256
rect 26810 656 27770 1256
rect 27828 656 28788 1256
rect 28846 656 29806 1256
rect 29864 656 30824 1256
rect 30882 656 31842 1256
rect 31900 656 32860 1256
rect 32918 656 33878 1256
rect 48850 7140 49050 7340
rect 49108 7140 49308 7340
rect 49366 7140 49566 7340
rect 49624 7140 49824 7340
rect 49882 7140 50082 7340
rect 50140 7140 50340 7340
rect 48850 5176 49050 5376
rect 49108 5176 49308 5376
rect 49366 5176 49566 5376
rect 49624 5176 49824 5376
rect 49882 5176 50082 5376
rect 50140 5176 50340 5376
rect 48850 3176 49050 3376
rect 49108 3176 49308 3376
rect 49366 3176 49566 3376
rect 49624 3176 49824 3376
rect 49882 3176 50082 3376
rect 50140 3176 50340 3376
rect 48850 1086 49050 1286
rect 49108 1086 49308 1286
rect 49366 1086 49566 1286
rect 49624 1086 49824 1286
rect 49882 1086 50082 1286
rect 50140 1086 50340 1286
rect 67578 14222 68538 14822
rect 68596 14222 69556 14822
rect 69614 14222 70574 14822
rect 70632 14222 71592 14822
rect 71650 14222 72610 14822
rect 72668 14222 73628 14822
rect 73686 14222 74646 14822
rect 74704 14222 75664 14822
rect 75722 14222 76682 14822
rect 76740 14222 77700 14822
rect 77758 14222 78718 14822
rect 78776 14222 79736 14822
rect 79794 14222 80754 14822
rect 80812 14222 81772 14822
rect 81830 14222 82790 14822
rect 82848 14222 83808 14822
rect 83866 14222 84826 14822
rect 84884 14222 85844 14822
rect 85902 14222 86862 14822
rect 86920 14222 87880 14822
rect 67578 12988 68538 13588
rect 68596 12988 69556 13588
rect 69614 12988 70574 13588
rect 70632 12988 71592 13588
rect 71650 12988 72610 13588
rect 72668 12988 73628 13588
rect 73686 12988 74646 13588
rect 74704 12988 75664 13588
rect 75722 12988 76682 13588
rect 76740 12988 77700 13588
rect 77758 12988 78718 13588
rect 78776 12988 79736 13588
rect 79794 12988 80754 13588
rect 80812 12988 81772 13588
rect 81830 12988 82790 13588
rect 82848 12988 83808 13588
rect 83866 12988 84826 13588
rect 84884 12988 85844 13588
rect 85902 12988 86862 13588
rect 86920 12988 87880 13588
rect 67578 11756 68538 12356
rect 68596 11756 69556 12356
rect 69614 11756 70574 12356
rect 70632 11756 71592 12356
rect 71650 11756 72610 12356
rect 72668 11756 73628 12356
rect 73686 11756 74646 12356
rect 74704 11756 75664 12356
rect 75722 11756 76682 12356
rect 76740 11756 77700 12356
rect 77758 11756 78718 12356
rect 78776 11756 79736 12356
rect 79794 11756 80754 12356
rect 80812 11756 81772 12356
rect 81830 11756 82790 12356
rect 82848 11756 83808 12356
rect 83866 11756 84826 12356
rect 84884 11756 85844 12356
rect 85902 11756 86862 12356
rect 86920 11756 87880 12356
rect 67576 10522 68536 11122
rect 68594 10522 69554 11122
rect 69612 10522 70572 11122
rect 70630 10522 71590 11122
rect 71648 10522 72608 11122
rect 72666 10522 73626 11122
rect 73684 10522 74644 11122
rect 74702 10522 75662 11122
rect 75720 10522 76680 11122
rect 76738 10522 77698 11122
rect 77756 10522 78716 11122
rect 78774 10522 79734 11122
rect 79792 10522 80752 11122
rect 80810 10522 81770 11122
rect 81828 10522 82788 11122
rect 82846 10522 83806 11122
rect 83864 10522 84824 11122
rect 84882 10522 85842 11122
rect 85900 10522 86860 11122
rect 86918 10522 87878 11122
rect 67576 9288 68536 9888
rect 68594 9288 69554 9888
rect 69612 9288 70572 9888
rect 70630 9288 71590 9888
rect 71648 9288 72608 9888
rect 72666 9288 73626 9888
rect 73684 9288 74644 9888
rect 74702 9288 75662 9888
rect 75720 9288 76680 9888
rect 76738 9288 77698 9888
rect 77756 9288 78716 9888
rect 78774 9288 79734 9888
rect 79792 9288 80752 9888
rect 80810 9288 81770 9888
rect 81828 9288 82788 9888
rect 82846 9288 83806 9888
rect 83864 9288 84824 9888
rect 84882 9288 85842 9888
rect 85900 9288 86860 9888
rect 86918 9288 87878 9888
rect 67576 8056 68536 8656
rect 68594 8056 69554 8656
rect 69612 8056 70572 8656
rect 70630 8056 71590 8656
rect 71648 8056 72608 8656
rect 72666 8056 73626 8656
rect 73684 8056 74644 8656
rect 74702 8056 75662 8656
rect 75720 8056 76680 8656
rect 76738 8056 77698 8656
rect 77756 8056 78716 8656
rect 78774 8056 79734 8656
rect 79792 8056 80752 8656
rect 80810 8056 81770 8656
rect 81828 8056 82788 8656
rect 82846 8056 83806 8656
rect 83864 8056 84824 8656
rect 84882 8056 85842 8656
rect 85900 8056 86860 8656
rect 86918 8056 87878 8656
rect 67576 6822 68536 7422
rect 68594 6822 69554 7422
rect 69612 6822 70572 7422
rect 70630 6822 71590 7422
rect 71648 6822 72608 7422
rect 72666 6822 73626 7422
rect 73684 6822 74644 7422
rect 74702 6822 75662 7422
rect 75720 6822 76680 7422
rect 76738 6822 77698 7422
rect 77756 6822 78716 7422
rect 78774 6822 79734 7422
rect 79792 6822 80752 7422
rect 80810 6822 81770 7422
rect 81828 6822 82788 7422
rect 82846 6822 83806 7422
rect 83864 6822 84824 7422
rect 84882 6822 85842 7422
rect 85900 6822 86860 7422
rect 86918 6822 87878 7422
rect 67576 5588 68536 6188
rect 68594 5588 69554 6188
rect 69612 5588 70572 6188
rect 70630 5588 71590 6188
rect 71648 5588 72608 6188
rect 72666 5588 73626 6188
rect 73684 5588 74644 6188
rect 74702 5588 75662 6188
rect 75720 5588 76680 6188
rect 76738 5588 77698 6188
rect 77756 5588 78716 6188
rect 78774 5588 79734 6188
rect 79792 5588 80752 6188
rect 80810 5588 81770 6188
rect 81828 5588 82788 6188
rect 82846 5588 83806 6188
rect 83864 5588 84824 6188
rect 84882 5588 85842 6188
rect 85900 5588 86860 6188
rect 86918 5588 87878 6188
rect 55591 4159 56551 4759
rect 56609 4159 57569 4759
rect 57627 4159 58587 4759
rect 58645 4159 59605 4759
rect 59663 4159 60623 4759
rect 60681 4159 61641 4759
rect 67576 4356 68536 4956
rect 68594 4356 69554 4956
rect 69612 4356 70572 4956
rect 70630 4356 71590 4956
rect 71648 4356 72608 4956
rect 72666 4356 73626 4956
rect 73684 4356 74644 4956
rect 74702 4356 75662 4956
rect 75720 4356 76680 4956
rect 76738 4356 77698 4956
rect 77756 4356 78716 4956
rect 78774 4356 79734 4956
rect 79792 4356 80752 4956
rect 80810 4356 81770 4956
rect 81828 4356 82788 4956
rect 82846 4356 83806 4956
rect 83864 4356 84824 4956
rect 84882 4356 85842 4956
rect 85900 4356 86860 4956
rect 86918 4356 87878 4956
rect 55590 3046 56550 3646
rect 56608 3046 57568 3646
rect 57626 3046 58586 3646
rect 58644 3046 59604 3646
rect 59662 3046 60622 3646
rect 60680 3046 61640 3646
rect 67576 3122 68536 3722
rect 68594 3122 69554 3722
rect 69612 3122 70572 3722
rect 70630 3122 71590 3722
rect 71648 3122 72608 3722
rect 72666 3122 73626 3722
rect 73684 3122 74644 3722
rect 74702 3122 75662 3722
rect 75720 3122 76680 3722
rect 76738 3122 77698 3722
rect 77756 3122 78716 3722
rect 78774 3122 79734 3722
rect 79792 3122 80752 3722
rect 80810 3122 81770 3722
rect 81828 3122 82788 3722
rect 82846 3122 83806 3722
rect 83864 3122 84824 3722
rect 84882 3122 85842 3722
rect 85900 3122 86860 3722
rect 86918 3122 87878 3722
rect 55591 1935 56551 2535
rect 56609 1935 57569 2535
rect 57627 1935 58587 2535
rect 58645 1935 59605 2535
rect 59663 1935 60623 2535
rect 60681 1935 61641 2535
rect 67576 1888 68536 2488
rect 68594 1888 69554 2488
rect 69612 1888 70572 2488
rect 70630 1888 71590 2488
rect 71648 1888 72608 2488
rect 72666 1888 73626 2488
rect 73684 1888 74644 2488
rect 74702 1888 75662 2488
rect 75720 1888 76680 2488
rect 76738 1888 77698 2488
rect 77756 1888 78716 2488
rect 78774 1888 79734 2488
rect 79792 1888 80752 2488
rect 80810 1888 81770 2488
rect 81828 1888 82788 2488
rect 82846 1888 83806 2488
rect 83864 1888 84824 2488
rect 84882 1888 85842 2488
rect 85900 1888 86860 2488
rect 86918 1888 87878 2488
rect 55590 822 56550 1422
rect 56608 822 57568 1422
rect 57626 822 58586 1422
rect 58644 822 59604 1422
rect 59662 822 60622 1422
rect 60680 822 61640 1422
rect 67576 656 68536 1256
rect 68594 656 69554 1256
rect 69612 656 70572 1256
rect 70630 656 71590 1256
rect 71648 656 72608 1256
rect 72666 656 73626 1256
rect 73684 656 74644 1256
rect 74702 656 75662 1256
rect 75720 656 76680 1256
rect 76738 656 77698 1256
rect 77756 656 78716 1256
rect 78774 656 79734 1256
rect 79792 656 80752 1256
rect 80810 656 81770 1256
rect 81828 656 82788 1256
rect 82846 656 83806 1256
rect 83864 656 84824 1256
rect 84882 656 85842 1256
rect 85900 656 86860 1256
rect 86918 656 87878 1256
<< scnmos >>
rect 49274 24395 49304 24525
rect 49274 22395 49304 22525
rect -11084 15265 -11054 15395
rect -8484 15265 -8454 15395
rect -7984 15265 -7954 15395
rect 50700 7431 50730 7561
rect 50700 5467 50730 5597
rect 50700 3467 50730 3597
rect 50700 1377 50730 1507
<< pmos >>
rect 18470 22334 19430 22934
rect 19488 22334 20448 22934
rect 20506 22334 21466 22934
rect 21524 22334 22484 22934
rect 22542 22334 23502 22934
rect 23560 22334 24520 22934
rect 24578 22334 25538 22934
rect 25596 22334 26556 22934
rect 26614 22334 27574 22934
rect 27632 22334 28592 22934
rect 28650 22334 29610 22934
rect 29668 22334 30628 22934
rect 30686 22334 31646 22934
rect 31704 22334 32664 22934
rect 32722 22334 33682 22934
rect 14622 21450 14782 21850
rect 14840 21450 15000 21850
rect 15058 21450 15218 21850
rect 15276 21450 15436 21850
rect 15494 21450 15654 21850
rect 15712 21450 15872 21850
rect 15930 21450 16090 21850
rect 16148 21450 16308 21850
rect 16366 21450 16526 21850
rect 16584 21450 16744 21850
rect 18470 21078 19430 21678
rect 19488 21078 20448 21678
rect 20506 21078 21466 21678
rect 21524 21078 22484 21678
rect 22542 21078 23502 21678
rect 23560 21078 24520 21678
rect 24578 21078 25538 21678
rect 25596 21078 26556 21678
rect 26614 21078 27574 21678
rect 27632 21078 28592 21678
rect 28650 21078 29610 21678
rect 29668 21078 30628 21678
rect 30686 21078 31646 21678
rect 31704 21078 32664 21678
rect 32722 21078 33682 21678
rect 14622 20512 14782 20912
rect 14840 20512 15000 20912
rect 15058 20512 15218 20912
rect 15276 20512 15436 20912
rect 15494 20512 15654 20912
rect 15712 20512 15872 20912
rect 15930 20512 16090 20912
rect 16148 20512 16308 20912
rect 16366 20512 16526 20912
rect 16584 20512 16744 20912
rect 14622 19574 14782 19974
rect 14840 19574 15000 19974
rect 15058 19574 15218 19974
rect 15276 19574 15436 19974
rect 15494 19574 15654 19974
rect 15712 19574 15872 19974
rect 15930 19574 16090 19974
rect 16148 19574 16308 19974
rect 16366 19574 16526 19974
rect 16584 19574 16744 19974
rect 18470 19822 19430 20422
rect 19488 19822 20448 20422
rect 20506 19822 21466 20422
rect 21524 19822 22484 20422
rect 22542 19822 23502 20422
rect 23560 19822 24520 20422
rect 24578 19822 25538 20422
rect 25596 19822 26556 20422
rect 26614 19822 27574 20422
rect 27632 19822 28592 20422
rect 28650 19822 29610 20422
rect 29668 19822 30628 20422
rect 30686 19822 31646 20422
rect 31704 19822 32664 20422
rect 32722 19822 33682 20422
rect 14622 18636 14782 19036
rect 14840 18636 15000 19036
rect 15058 18636 15218 19036
rect 15276 18636 15436 19036
rect 15494 18636 15654 19036
rect 15712 18636 15872 19036
rect 15930 18636 16090 19036
rect 16148 18636 16308 19036
rect 16366 18636 16526 19036
rect 16584 18636 16744 19036
rect 18470 18566 19430 19166
rect 19488 18566 20448 19166
rect 20506 18566 21466 19166
rect 21524 18566 22484 19166
rect 22542 18566 23502 19166
rect 23560 18566 24520 19166
rect 24578 18566 25538 19166
rect 25596 18566 26556 19166
rect 26614 18566 27574 19166
rect 27632 18566 28592 19166
rect 28650 18566 29610 19166
rect 29668 18566 30628 19166
rect 30686 18566 31646 19166
rect 31704 18566 32664 19166
rect 32722 18566 33682 19166
rect 72470 22334 73430 22934
rect 73488 22334 74448 22934
rect 74506 22334 75466 22934
rect 75524 22334 76484 22934
rect 76542 22334 77502 22934
rect 77560 22334 78520 22934
rect 78578 22334 79538 22934
rect 79596 22334 80556 22934
rect 80614 22334 81574 22934
rect 81632 22334 82592 22934
rect 82650 22334 83610 22934
rect 83668 22334 84628 22934
rect 84686 22334 85646 22934
rect 85704 22334 86664 22934
rect 86722 22334 87682 22934
rect 68622 21450 68782 21850
rect 68840 21450 69000 21850
rect 69058 21450 69218 21850
rect 69276 21450 69436 21850
rect 69494 21450 69654 21850
rect 69712 21450 69872 21850
rect 69930 21450 70090 21850
rect 70148 21450 70308 21850
rect 70366 21450 70526 21850
rect 70584 21450 70744 21850
rect 72470 21078 73430 21678
rect 73488 21078 74448 21678
rect 74506 21078 75466 21678
rect 75524 21078 76484 21678
rect 76542 21078 77502 21678
rect 77560 21078 78520 21678
rect 78578 21078 79538 21678
rect 79596 21078 80556 21678
rect 80614 21078 81574 21678
rect 81632 21078 82592 21678
rect 82650 21078 83610 21678
rect 83668 21078 84628 21678
rect 84686 21078 85646 21678
rect 85704 21078 86664 21678
rect 86722 21078 87682 21678
rect 68622 20512 68782 20912
rect 68840 20512 69000 20912
rect 69058 20512 69218 20912
rect 69276 20512 69436 20912
rect 69494 20512 69654 20912
rect 69712 20512 69872 20912
rect 69930 20512 70090 20912
rect 70148 20512 70308 20912
rect 70366 20512 70526 20912
rect 70584 20512 70744 20912
rect 68622 19574 68782 19974
rect 68840 19574 69000 19974
rect 69058 19574 69218 19974
rect 69276 19574 69436 19974
rect 69494 19574 69654 19974
rect 69712 19574 69872 19974
rect 69930 19574 70090 19974
rect 70148 19574 70308 19974
rect 70366 19574 70526 19974
rect 70584 19574 70744 19974
rect 72470 19822 73430 20422
rect 73488 19822 74448 20422
rect 74506 19822 75466 20422
rect 75524 19822 76484 20422
rect 76542 19822 77502 20422
rect 77560 19822 78520 20422
rect 78578 19822 79538 20422
rect 79596 19822 80556 20422
rect 80614 19822 81574 20422
rect 81632 19822 82592 20422
rect 82650 19822 83610 20422
rect 83668 19822 84628 20422
rect 84686 19822 85646 20422
rect 85704 19822 86664 20422
rect 86722 19822 87682 20422
rect 68622 18636 68782 19036
rect 68840 18636 69000 19036
rect 69058 18636 69218 19036
rect 69276 18636 69436 19036
rect 69494 18636 69654 19036
rect 69712 18636 69872 19036
rect 69930 18636 70090 19036
rect 70148 18636 70308 19036
rect 70366 18636 70526 19036
rect 70584 18636 70744 19036
rect 72470 18566 73430 19166
rect 73488 18566 74448 19166
rect 74506 18566 75466 19166
rect 75524 18566 76484 19166
rect 76542 18566 77502 19166
rect 77560 18566 78520 19166
rect 78578 18566 79538 19166
rect 79596 18566 80556 19166
rect 80614 18566 81574 19166
rect 81632 18566 82592 19166
rect 82650 18566 83610 19166
rect 83668 18566 84628 19166
rect 84686 18566 85646 19166
rect 85704 18566 86664 19166
rect 86722 18566 87682 19166
<< scpmoshvt >>
rect 49274 24645 49304 24845
rect 49274 22645 49304 22845
rect -11084 15515 -11054 15715
rect -8484 15515 -8454 15715
rect -7984 15515 -7954 15715
rect 50700 7681 50730 7881
rect 50700 5717 50730 5917
rect 50700 3717 50730 3917
rect 50700 1627 50730 1827
<< pmoslvt >>
rect 17484 26380 18444 26980
rect 18502 26380 19462 26980
rect 19520 26380 20480 26980
rect 20538 26380 21498 26980
rect 21556 26380 22516 26980
rect 22574 26380 23534 26980
rect 23592 26380 24552 26980
rect 24610 26380 25570 26980
rect 25628 26380 26588 26980
rect 26646 26380 27606 26980
rect 27664 26380 28624 26980
rect 28682 26380 29642 26980
rect 29700 26380 30660 26980
rect 30718 26380 31678 26980
rect 31736 26380 32696 26980
rect 32754 26380 33714 26980
rect 17484 25244 18444 25844
rect 18502 25244 19462 25844
rect 19520 25244 20480 25844
rect 20538 25244 21498 25844
rect 21556 25244 22516 25844
rect 22574 25244 23534 25844
rect 23592 25244 24552 25844
rect 24610 25244 25570 25844
rect 25628 25244 26588 25844
rect 26646 25244 27606 25844
rect 27664 25244 28624 25844
rect 28682 25244 29642 25844
rect 29700 25244 30660 25844
rect 30718 25244 31678 25844
rect 31736 25244 32696 25844
rect 32754 25244 33714 25844
rect 17484 24108 18444 24708
rect 18502 24108 19462 24708
rect 19520 24108 20480 24708
rect 20538 24108 21498 24708
rect 21556 24108 22516 24708
rect 22574 24108 23534 24708
rect 23592 24108 24552 24708
rect 24610 24108 25570 24708
rect 25628 24108 26588 24708
rect 26646 24108 27606 24708
rect 27664 24108 28624 24708
rect 28682 24108 29642 24708
rect 29700 24108 30660 24708
rect 30718 24108 31678 24708
rect 31736 24108 32696 24708
rect 32754 24108 33714 24708
rect 71484 26380 72444 26980
rect 72502 26380 73462 26980
rect 73520 26380 74480 26980
rect 74538 26380 75498 26980
rect 75556 26380 76516 26980
rect 76574 26380 77534 26980
rect 77592 26380 78552 26980
rect 78610 26380 79570 26980
rect 79628 26380 80588 26980
rect 80646 26380 81606 26980
rect 81664 26380 82624 26980
rect 82682 26380 83642 26980
rect 83700 26380 84660 26980
rect 84718 26380 85678 26980
rect 85736 26380 86696 26980
rect 86754 26380 87714 26980
rect 71484 25244 72444 25844
rect 72502 25244 73462 25844
rect 73520 25244 74480 25844
rect 74538 25244 75498 25844
rect 75556 25244 76516 25844
rect 76574 25244 77534 25844
rect 77592 25244 78552 25844
rect 78610 25244 79570 25844
rect 79628 25244 80588 25844
rect 80646 25244 81606 25844
rect 81664 25244 82624 25844
rect 82682 25244 83642 25844
rect 83700 25244 84660 25844
rect 84718 25244 85678 25844
rect 85736 25244 86696 25844
rect 86754 25244 87714 25844
rect 71484 24108 72444 24708
rect 72502 24108 73462 24708
rect 73520 24108 74480 24708
rect 74538 24108 75498 24708
rect 75556 24108 76516 24708
rect 76574 24108 77534 24708
rect 77592 24108 78552 24708
rect 78610 24108 79570 24708
rect 79628 24108 80588 24708
rect 80646 24108 81606 24708
rect 81664 24108 82624 24708
rect 82682 24108 83642 24708
rect 83700 24108 84660 24708
rect 84718 24108 85678 24708
rect 85736 24108 86696 24708
rect 86754 24108 87714 24708
<< pmoshvt >>
rect 47424 24828 47624 25228
rect 47682 24828 47882 25228
rect 47940 24828 48140 25228
rect 48198 24828 48398 25228
rect 48456 24828 48656 25228
rect 48714 24828 48914 25228
rect 47424 22828 47624 23228
rect 47682 22828 47882 23228
rect 47940 22828 48140 23228
rect 48198 22828 48398 23228
rect 48456 22828 48656 23228
rect 48714 22828 48914 23228
rect -12934 15698 -12734 16098
rect -12676 15698 -12476 16098
rect -12418 15698 -12218 16098
rect -12160 15698 -11960 16098
rect -11902 15698 -11702 16098
rect -11644 15698 -11444 16098
rect -10334 15698 -10134 16098
rect -10076 15698 -9876 16098
rect -9818 15698 -9618 16098
rect -9560 15698 -9360 16098
rect -9302 15698 -9102 16098
rect -9044 15698 -8844 16098
rect 48850 7864 49050 8264
rect 49108 7864 49308 8264
rect 49366 7864 49566 8264
rect 49624 7864 49824 8264
rect 49882 7864 50082 8264
rect 50140 7864 50340 8264
rect 48850 5900 49050 6300
rect 49108 5900 49308 6300
rect 49366 5900 49566 6300
rect 49624 5900 49824 6300
rect 49882 5900 50082 6300
rect 50140 5900 50340 6300
rect 48850 3900 49050 4300
rect 49108 3900 49308 4300
rect 49366 3900 49566 4300
rect 49624 3900 49824 4300
rect 49882 3900 50082 4300
rect 50140 3900 50340 4300
rect 48850 1810 49050 2210
rect 49108 1810 49308 2210
rect 49366 1810 49566 2210
rect 49624 1810 49824 2210
rect 49882 1810 50082 2210
rect 50140 1810 50340 2210
<< nmoslvt >>
rect 1812 13428 2772 14028
rect 2830 13428 3790 14028
rect 3848 13428 4808 14028
rect 4866 13428 5826 14028
rect 5884 13428 6844 14028
rect 6902 13428 7862 14028
rect 7920 13428 8880 14028
rect 8938 13428 9898 14028
rect 9956 13428 10916 14028
rect 1812 12610 2772 13210
rect 2830 12610 3790 13210
rect 3848 12610 4808 13210
rect 4866 12610 5826 13210
rect 5884 12610 6844 13210
rect 6902 12610 7862 13210
rect 7920 12610 8880 13210
rect 8938 12610 9898 13210
rect 9956 12610 10916 13210
rect 1812 11792 2772 12392
rect 2830 11792 3790 12392
rect 3848 11792 4808 12392
rect 4866 11792 5826 12392
rect 5884 11792 6844 12392
rect 6902 11792 7862 12392
rect 7920 11792 8880 12392
rect 8938 11792 9898 12392
rect 9956 11792 10916 12392
rect 1812 10974 2772 11574
rect 2830 10974 3790 11574
rect 3848 10974 4808 11574
rect 4866 10974 5826 11574
rect 5884 10974 6844 11574
rect 6902 10974 7862 11574
rect 7920 10974 8880 11574
rect 8938 10974 9898 11574
rect 9956 10974 10916 11574
rect 1812 10156 2772 10756
rect 2830 10156 3790 10756
rect 3848 10156 4808 10756
rect 4866 10156 5826 10756
rect 5884 10156 6844 10756
rect 6902 10156 7862 10756
rect 7920 10156 8880 10756
rect 8938 10156 9898 10756
rect 9956 10156 10916 10756
rect 1812 9338 2772 9938
rect 2830 9338 3790 9938
rect 3848 9338 4808 9938
rect 4866 9338 5826 9938
rect 5884 9338 6844 9938
rect 6902 9338 7862 9938
rect 7920 9338 8880 9938
rect 8938 9338 9898 9938
rect 9956 9338 10916 9938
rect 1812 8520 2772 9120
rect 2830 8520 3790 9120
rect 3848 8520 4808 9120
rect 4866 8520 5826 9120
rect 5884 8520 6844 9120
rect 6902 8520 7862 9120
rect 7920 8520 8880 9120
rect 8938 8520 9898 9120
rect 9956 8520 10916 9120
rect 1812 7702 2772 8302
rect 2830 7702 3790 8302
rect 3848 7702 4808 8302
rect 4866 7702 5826 8302
rect 5884 7702 6844 8302
rect 6902 7702 7862 8302
rect 7920 7702 8880 8302
rect 8938 7702 9898 8302
rect 9956 7702 10916 8302
rect 8672 6718 8832 6918
rect 8890 6718 9050 6918
rect 9108 6718 9268 6918
rect 9326 6718 9486 6918
rect 9544 6718 9704 6918
rect 9762 6718 9922 6918
rect 9980 6718 10140 6918
rect 10198 6718 10358 6918
rect 10416 6718 10576 6918
rect 10634 6718 10794 6918
rect 8672 5886 8832 6086
rect 8890 5886 9050 6086
rect 9108 5886 9268 6086
rect 9326 5886 9486 6086
rect 9544 5886 9704 6086
rect 9762 5886 9922 6086
rect 9980 5886 10140 6086
rect 10198 5886 10358 6086
rect 10416 5886 10576 6086
rect 10634 5886 10794 6086
rect 8586 4160 8826 4760
rect 8884 4160 9124 4760
rect 9182 4160 9422 4760
rect 9480 4160 9720 4760
rect 9778 4160 10018 4760
rect 10076 4160 10316 4760
rect 10374 4160 10614 4760
rect 10672 4160 10912 4760
rect 10970 4160 11210 4760
rect 11268 4160 11508 4760
rect 11566 4160 11806 4760
rect 8586 3048 8826 3648
rect 8884 3048 9124 3648
rect 9182 3048 9422 3648
rect 9480 3048 9720 3648
rect 9778 3048 10018 3648
rect 10076 3048 10316 3648
rect 10374 3048 10614 3648
rect 10672 3048 10912 3648
rect 10970 3048 11210 3648
rect 11268 3048 11508 3648
rect 11566 3048 11806 3648
rect 8584 1936 8824 2536
rect 8882 1936 9122 2536
rect 9180 1936 9420 2536
rect 9478 1936 9718 2536
rect 9776 1936 10016 2536
rect 10074 1936 10314 2536
rect 10372 1936 10612 2536
rect 10670 1936 10910 2536
rect 10968 1936 11208 2536
rect 11266 1936 11506 2536
rect 11564 1936 11804 2536
rect 8584 826 8824 1426
rect 8882 826 9122 1426
rect 9180 826 9420 1426
rect 9478 826 9718 1426
rect 9776 826 10016 1426
rect 10074 826 10314 1426
rect 10372 826 10612 1426
rect 10670 826 10910 1426
rect 10968 826 11208 1426
rect 11266 826 11506 1426
rect 11564 826 11804 1426
rect 55812 13428 56772 14028
rect 56830 13428 57790 14028
rect 57848 13428 58808 14028
rect 58866 13428 59826 14028
rect 59884 13428 60844 14028
rect 60902 13428 61862 14028
rect 61920 13428 62880 14028
rect 62938 13428 63898 14028
rect 63956 13428 64916 14028
rect 55812 12610 56772 13210
rect 56830 12610 57790 13210
rect 57848 12610 58808 13210
rect 58866 12610 59826 13210
rect 59884 12610 60844 13210
rect 60902 12610 61862 13210
rect 61920 12610 62880 13210
rect 62938 12610 63898 13210
rect 63956 12610 64916 13210
rect 55812 11792 56772 12392
rect 56830 11792 57790 12392
rect 57848 11792 58808 12392
rect 58866 11792 59826 12392
rect 59884 11792 60844 12392
rect 60902 11792 61862 12392
rect 61920 11792 62880 12392
rect 62938 11792 63898 12392
rect 63956 11792 64916 12392
rect 55812 10974 56772 11574
rect 56830 10974 57790 11574
rect 57848 10974 58808 11574
rect 58866 10974 59826 11574
rect 59884 10974 60844 11574
rect 60902 10974 61862 11574
rect 61920 10974 62880 11574
rect 62938 10974 63898 11574
rect 63956 10974 64916 11574
rect 55812 10156 56772 10756
rect 56830 10156 57790 10756
rect 57848 10156 58808 10756
rect 58866 10156 59826 10756
rect 59884 10156 60844 10756
rect 60902 10156 61862 10756
rect 61920 10156 62880 10756
rect 62938 10156 63898 10756
rect 63956 10156 64916 10756
rect 55812 9338 56772 9938
rect 56830 9338 57790 9938
rect 57848 9338 58808 9938
rect 58866 9338 59826 9938
rect 59884 9338 60844 9938
rect 60902 9338 61862 9938
rect 61920 9338 62880 9938
rect 62938 9338 63898 9938
rect 63956 9338 64916 9938
rect 55812 8520 56772 9120
rect 56830 8520 57790 9120
rect 57848 8520 58808 9120
rect 58866 8520 59826 9120
rect 59884 8520 60844 9120
rect 60902 8520 61862 9120
rect 61920 8520 62880 9120
rect 62938 8520 63898 9120
rect 63956 8520 64916 9120
rect 55812 7702 56772 8302
rect 56830 7702 57790 8302
rect 57848 7702 58808 8302
rect 58866 7702 59826 8302
rect 59884 7702 60844 8302
rect 60902 7702 61862 8302
rect 61920 7702 62880 8302
rect 62938 7702 63898 8302
rect 63956 7702 64916 8302
rect 62672 6718 62832 6918
rect 62890 6718 63050 6918
rect 63108 6718 63268 6918
rect 63326 6718 63486 6918
rect 63544 6718 63704 6918
rect 63762 6718 63922 6918
rect 63980 6718 64140 6918
rect 64198 6718 64358 6918
rect 64416 6718 64576 6918
rect 64634 6718 64794 6918
rect 62672 5886 62832 6086
rect 62890 5886 63050 6086
rect 63108 5886 63268 6086
rect 63326 5886 63486 6086
rect 63544 5886 63704 6086
rect 63762 5886 63922 6086
rect 63980 5886 64140 6086
rect 64198 5886 64358 6086
rect 64416 5886 64576 6086
rect 64634 5886 64794 6086
rect 62586 4160 62826 4760
rect 62884 4160 63124 4760
rect 63182 4160 63422 4760
rect 63480 4160 63720 4760
rect 63778 4160 64018 4760
rect 64076 4160 64316 4760
rect 64374 4160 64614 4760
rect 64672 4160 64912 4760
rect 64970 4160 65210 4760
rect 65268 4160 65508 4760
rect 65566 4160 65806 4760
rect 62586 3048 62826 3648
rect 62884 3048 63124 3648
rect 63182 3048 63422 3648
rect 63480 3048 63720 3648
rect 63778 3048 64018 3648
rect 64076 3048 64316 3648
rect 64374 3048 64614 3648
rect 64672 3048 64912 3648
rect 64970 3048 65210 3648
rect 65268 3048 65508 3648
rect 65566 3048 65806 3648
rect 62584 1936 62824 2536
rect 62882 1936 63122 2536
rect 63180 1936 63420 2536
rect 63478 1936 63718 2536
rect 63776 1936 64016 2536
rect 64074 1936 64314 2536
rect 64372 1936 64612 2536
rect 64670 1936 64910 2536
rect 64968 1936 65208 2536
rect 65266 1936 65506 2536
rect 65564 1936 65804 2536
rect 62584 826 62824 1426
rect 62882 826 63122 1426
rect 63180 826 63420 1426
rect 63478 826 63718 1426
rect 63776 826 64016 1426
rect 64074 826 64314 1426
rect 64372 826 64612 1426
rect 64670 826 64910 1426
rect 64968 826 65208 1426
rect 65266 826 65506 1426
rect 65564 826 65804 1426
<< ndiff >>
rect 49222 24513 49274 24525
rect 49222 24479 49230 24513
rect 49264 24479 49274 24513
rect 49222 24445 49274 24479
rect 49222 24411 49230 24445
rect 49264 24411 49274 24445
rect 49222 24395 49274 24411
rect 49304 24513 49356 24525
rect 49304 24479 49314 24513
rect 49348 24479 49356 24513
rect 49304 24445 49356 24479
rect 49304 24411 49314 24445
rect 49348 24411 49356 24445
rect 49304 24395 49356 24411
rect 47366 24292 47424 24304
rect 47366 24116 47378 24292
rect 47412 24116 47424 24292
rect 47366 24104 47424 24116
rect 47624 24292 47682 24304
rect 47624 24116 47636 24292
rect 47670 24116 47682 24292
rect 47624 24104 47682 24116
rect 47882 24292 47940 24304
rect 47882 24116 47894 24292
rect 47928 24116 47940 24292
rect 47882 24104 47940 24116
rect 48140 24292 48198 24304
rect 48140 24116 48152 24292
rect 48186 24116 48198 24292
rect 48140 24104 48198 24116
rect 48398 24292 48456 24304
rect 48398 24116 48410 24292
rect 48444 24116 48456 24292
rect 48398 24104 48456 24116
rect 48656 24292 48714 24304
rect 48656 24116 48668 24292
rect 48702 24116 48714 24292
rect 48656 24104 48714 24116
rect 48914 24292 48972 24304
rect 48914 24116 48926 24292
rect 48960 24116 48972 24292
rect 48914 24104 48972 24116
rect 49222 22513 49274 22525
rect 49222 22479 49230 22513
rect 49264 22479 49274 22513
rect 49222 22445 49274 22479
rect 49222 22411 49230 22445
rect 49264 22411 49274 22445
rect 49222 22395 49274 22411
rect 49304 22513 49356 22525
rect 49304 22479 49314 22513
rect 49348 22479 49356 22513
rect 49304 22445 49356 22479
rect 49304 22411 49314 22445
rect 49348 22411 49356 22445
rect 49304 22395 49356 22411
rect 47366 22292 47424 22304
rect 47366 22116 47378 22292
rect 47412 22116 47424 22292
rect 47366 22104 47424 22116
rect 47624 22292 47682 22304
rect 47624 22116 47636 22292
rect 47670 22116 47682 22292
rect 47624 22104 47682 22116
rect 47882 22292 47940 22304
rect 47882 22116 47894 22292
rect 47928 22116 47940 22292
rect 47882 22104 47940 22116
rect 48140 22292 48198 22304
rect 48140 22116 48152 22292
rect 48186 22116 48198 22292
rect 48140 22104 48198 22116
rect 48398 22292 48456 22304
rect 48398 22116 48410 22292
rect 48444 22116 48456 22292
rect 48398 22104 48456 22116
rect 48656 22292 48714 22304
rect 48656 22116 48668 22292
rect 48702 22116 48714 22292
rect 48656 22104 48714 22116
rect 48914 22292 48972 22304
rect 48914 22116 48926 22292
rect 48960 22116 48972 22292
rect 48914 22104 48972 22116
rect -11136 15383 -11084 15395
rect -11136 15349 -11128 15383
rect -11094 15349 -11084 15383
rect -11136 15315 -11084 15349
rect -11136 15281 -11128 15315
rect -11094 15281 -11084 15315
rect -11136 15265 -11084 15281
rect -11054 15383 -11002 15395
rect -11054 15349 -11044 15383
rect -11010 15349 -11002 15383
rect -11054 15315 -11002 15349
rect -8536 15383 -8484 15395
rect -8536 15349 -8528 15383
rect -8494 15349 -8484 15383
rect -11054 15281 -11044 15315
rect -11010 15281 -11002 15315
rect -11054 15265 -11002 15281
rect -12992 15162 -12934 15174
rect -12992 14986 -12980 15162
rect -12946 14986 -12934 15162
rect -12992 14974 -12934 14986
rect -12734 15162 -12676 15174
rect -12734 14986 -12722 15162
rect -12688 14986 -12676 15162
rect -12734 14974 -12676 14986
rect -12476 15162 -12418 15174
rect -12476 14986 -12464 15162
rect -12430 14986 -12418 15162
rect -12476 14974 -12418 14986
rect -12218 15162 -12160 15174
rect -12218 14986 -12206 15162
rect -12172 14986 -12160 15162
rect -12218 14974 -12160 14986
rect -11960 15162 -11902 15174
rect -11960 14986 -11948 15162
rect -11914 14986 -11902 15162
rect -11960 14974 -11902 14986
rect -11702 15162 -11644 15174
rect -11702 14986 -11690 15162
rect -11656 14986 -11644 15162
rect -11702 14974 -11644 14986
rect -11444 15162 -11386 15174
rect -11444 14986 -11432 15162
rect -11398 14986 -11386 15162
rect -11444 14974 -11386 14986
rect -8536 15315 -8484 15349
rect -8536 15281 -8528 15315
rect -8494 15281 -8484 15315
rect -8536 15265 -8484 15281
rect -8454 15383 -8402 15395
rect -8454 15349 -8444 15383
rect -8410 15349 -8402 15383
rect -8454 15315 -8402 15349
rect -8454 15281 -8444 15315
rect -8410 15281 -8402 15315
rect -8454 15265 -8402 15281
rect -8036 15383 -7984 15395
rect -8036 15349 -8028 15383
rect -7994 15349 -7984 15383
rect -8036 15315 -7984 15349
rect -8036 15281 -8028 15315
rect -7994 15281 -7984 15315
rect -8036 15265 -7984 15281
rect -7954 15383 -7902 15395
rect -7954 15349 -7944 15383
rect -7910 15349 -7902 15383
rect -7954 15315 -7902 15349
rect -7954 15281 -7944 15315
rect -7910 15281 -7902 15315
rect -7954 15265 -7902 15281
rect -10392 15162 -10334 15174
rect -10392 14986 -10380 15162
rect -10346 14986 -10334 15162
rect -10392 14974 -10334 14986
rect -10134 15162 -10076 15174
rect -10134 14986 -10122 15162
rect -10088 14986 -10076 15162
rect -10134 14974 -10076 14986
rect -9876 15162 -9818 15174
rect -9876 14986 -9864 15162
rect -9830 14986 -9818 15162
rect -9876 14974 -9818 14986
rect -9618 15162 -9560 15174
rect -9618 14986 -9606 15162
rect -9572 14986 -9560 15162
rect -9618 14974 -9560 14986
rect -9360 15162 -9302 15174
rect -9360 14986 -9348 15162
rect -9314 14986 -9302 15162
rect -9360 14974 -9302 14986
rect -9102 15162 -9044 15174
rect -9102 14986 -9090 15162
rect -9056 14986 -9044 15162
rect -9102 14974 -9044 14986
rect -8844 15162 -8786 15174
rect -8844 14986 -8832 15162
rect -8798 14986 -8786 15162
rect -8844 14974 -8786 14986
rect 13520 14810 13578 14822
rect 13520 14234 13532 14810
rect 13566 14234 13578 14810
rect 13520 14222 13578 14234
rect 14538 14810 14596 14822
rect 14538 14234 14550 14810
rect 14584 14234 14596 14810
rect 14538 14222 14596 14234
rect 15556 14810 15614 14822
rect 15556 14234 15568 14810
rect 15602 14234 15614 14810
rect 15556 14222 15614 14234
rect 16574 14810 16632 14822
rect 16574 14234 16586 14810
rect 16620 14234 16632 14810
rect 16574 14222 16632 14234
rect 17592 14810 17650 14822
rect 17592 14234 17604 14810
rect 17638 14234 17650 14810
rect 17592 14222 17650 14234
rect 18610 14810 18668 14822
rect 18610 14234 18622 14810
rect 18656 14234 18668 14810
rect 18610 14222 18668 14234
rect 19628 14810 19686 14822
rect 19628 14234 19640 14810
rect 19674 14234 19686 14810
rect 19628 14222 19686 14234
rect 20646 14810 20704 14822
rect 20646 14234 20658 14810
rect 20692 14234 20704 14810
rect 20646 14222 20704 14234
rect 21664 14810 21722 14822
rect 21664 14234 21676 14810
rect 21710 14234 21722 14810
rect 21664 14222 21722 14234
rect 22682 14810 22740 14822
rect 22682 14234 22694 14810
rect 22728 14234 22740 14810
rect 22682 14222 22740 14234
rect 23700 14810 23758 14822
rect 23700 14234 23712 14810
rect 23746 14234 23758 14810
rect 23700 14222 23758 14234
rect 24718 14810 24776 14822
rect 24718 14234 24730 14810
rect 24764 14234 24776 14810
rect 24718 14222 24776 14234
rect 25736 14810 25794 14822
rect 25736 14234 25748 14810
rect 25782 14234 25794 14810
rect 25736 14222 25794 14234
rect 26754 14810 26812 14822
rect 26754 14234 26766 14810
rect 26800 14234 26812 14810
rect 26754 14222 26812 14234
rect 27772 14810 27830 14822
rect 27772 14234 27784 14810
rect 27818 14234 27830 14810
rect 27772 14222 27830 14234
rect 28790 14810 28848 14822
rect 28790 14234 28802 14810
rect 28836 14234 28848 14810
rect 28790 14222 28848 14234
rect 29808 14810 29866 14822
rect 29808 14234 29820 14810
rect 29854 14234 29866 14810
rect 29808 14222 29866 14234
rect 30826 14810 30884 14822
rect 30826 14234 30838 14810
rect 30872 14234 30884 14810
rect 30826 14222 30884 14234
rect 31844 14810 31902 14822
rect 31844 14234 31856 14810
rect 31890 14234 31902 14810
rect 31844 14222 31902 14234
rect 32862 14810 32920 14822
rect 32862 14234 32874 14810
rect 32908 14234 32920 14810
rect 32862 14222 32920 14234
rect 33880 14810 33938 14822
rect 33880 14234 33892 14810
rect 33926 14234 33938 14810
rect 33880 14222 33938 14234
rect 1754 14016 1812 14028
rect 1754 13440 1766 14016
rect 1800 13440 1812 14016
rect 1754 13428 1812 13440
rect 2772 14016 2830 14028
rect 2772 13440 2784 14016
rect 2818 13440 2830 14016
rect 2772 13428 2830 13440
rect 3790 14016 3848 14028
rect 3790 13440 3802 14016
rect 3836 13440 3848 14016
rect 3790 13428 3848 13440
rect 4808 14016 4866 14028
rect 4808 13440 4820 14016
rect 4854 13440 4866 14016
rect 4808 13428 4866 13440
rect 5826 14016 5884 14028
rect 5826 13440 5838 14016
rect 5872 13440 5884 14016
rect 5826 13428 5884 13440
rect 6844 14016 6902 14028
rect 6844 13440 6856 14016
rect 6890 13440 6902 14016
rect 6844 13428 6902 13440
rect 7862 14016 7920 14028
rect 7862 13440 7874 14016
rect 7908 13440 7920 14016
rect 7862 13428 7920 13440
rect 8880 14016 8938 14028
rect 8880 13440 8892 14016
rect 8926 13440 8938 14016
rect 8880 13428 8938 13440
rect 9898 14016 9956 14028
rect 9898 13440 9910 14016
rect 9944 13440 9956 14016
rect 9898 13428 9956 13440
rect 10916 14016 10974 14028
rect 10916 13440 10928 14016
rect 10962 13440 10974 14016
rect 10916 13428 10974 13440
rect 13520 13576 13578 13588
rect 1754 13198 1812 13210
rect 1754 12622 1766 13198
rect 1800 12622 1812 13198
rect 1754 12610 1812 12622
rect 2772 13198 2830 13210
rect 2772 12622 2784 13198
rect 2818 12622 2830 13198
rect 2772 12610 2830 12622
rect 3790 13198 3848 13210
rect 3790 12622 3802 13198
rect 3836 12622 3848 13198
rect 3790 12610 3848 12622
rect 4808 13198 4866 13210
rect 4808 12622 4820 13198
rect 4854 12622 4866 13198
rect 4808 12610 4866 12622
rect 5826 13198 5884 13210
rect 5826 12622 5838 13198
rect 5872 12622 5884 13198
rect 5826 12610 5884 12622
rect 6844 13198 6902 13210
rect 6844 12622 6856 13198
rect 6890 12622 6902 13198
rect 6844 12610 6902 12622
rect 7862 13198 7920 13210
rect 7862 12622 7874 13198
rect 7908 12622 7920 13198
rect 7862 12610 7920 12622
rect 8880 13198 8938 13210
rect 8880 12622 8892 13198
rect 8926 12622 8938 13198
rect 8880 12610 8938 12622
rect 9898 13198 9956 13210
rect 9898 12622 9910 13198
rect 9944 12622 9956 13198
rect 9898 12610 9956 12622
rect 10916 13198 10974 13210
rect 10916 12622 10928 13198
rect 10962 12622 10974 13198
rect 13520 13000 13532 13576
rect 13566 13000 13578 13576
rect 13520 12988 13578 13000
rect 14538 13576 14596 13588
rect 14538 13000 14550 13576
rect 14584 13000 14596 13576
rect 14538 12988 14596 13000
rect 15556 13576 15614 13588
rect 15556 13000 15568 13576
rect 15602 13000 15614 13576
rect 15556 12988 15614 13000
rect 16574 13576 16632 13588
rect 16574 13000 16586 13576
rect 16620 13000 16632 13576
rect 16574 12988 16632 13000
rect 17592 13576 17650 13588
rect 17592 13000 17604 13576
rect 17638 13000 17650 13576
rect 17592 12988 17650 13000
rect 18610 13576 18668 13588
rect 18610 13000 18622 13576
rect 18656 13000 18668 13576
rect 18610 12988 18668 13000
rect 19628 13576 19686 13588
rect 19628 13000 19640 13576
rect 19674 13000 19686 13576
rect 19628 12988 19686 13000
rect 20646 13576 20704 13588
rect 20646 13000 20658 13576
rect 20692 13000 20704 13576
rect 20646 12988 20704 13000
rect 21664 13576 21722 13588
rect 21664 13000 21676 13576
rect 21710 13000 21722 13576
rect 21664 12988 21722 13000
rect 22682 13576 22740 13588
rect 22682 13000 22694 13576
rect 22728 13000 22740 13576
rect 22682 12988 22740 13000
rect 23700 13576 23758 13588
rect 23700 13000 23712 13576
rect 23746 13000 23758 13576
rect 23700 12988 23758 13000
rect 24718 13576 24776 13588
rect 24718 13000 24730 13576
rect 24764 13000 24776 13576
rect 24718 12988 24776 13000
rect 25736 13576 25794 13588
rect 25736 13000 25748 13576
rect 25782 13000 25794 13576
rect 25736 12988 25794 13000
rect 26754 13576 26812 13588
rect 26754 13000 26766 13576
rect 26800 13000 26812 13576
rect 26754 12988 26812 13000
rect 27772 13576 27830 13588
rect 27772 13000 27784 13576
rect 27818 13000 27830 13576
rect 27772 12988 27830 13000
rect 28790 13576 28848 13588
rect 28790 13000 28802 13576
rect 28836 13000 28848 13576
rect 28790 12988 28848 13000
rect 29808 13576 29866 13588
rect 29808 13000 29820 13576
rect 29854 13000 29866 13576
rect 29808 12988 29866 13000
rect 30826 13576 30884 13588
rect 30826 13000 30838 13576
rect 30872 13000 30884 13576
rect 30826 12988 30884 13000
rect 31844 13576 31902 13588
rect 31844 13000 31856 13576
rect 31890 13000 31902 13576
rect 31844 12988 31902 13000
rect 32862 13576 32920 13588
rect 32862 13000 32874 13576
rect 32908 13000 32920 13576
rect 32862 12988 32920 13000
rect 33880 13576 33938 13588
rect 33880 13000 33892 13576
rect 33926 13000 33938 13576
rect 33880 12988 33938 13000
rect 10916 12610 10974 12622
rect 1754 12380 1812 12392
rect 1754 11804 1766 12380
rect 1800 11804 1812 12380
rect 1754 11792 1812 11804
rect 2772 12380 2830 12392
rect 2772 11804 2784 12380
rect 2818 11804 2830 12380
rect 2772 11792 2830 11804
rect 3790 12380 3848 12392
rect 3790 11804 3802 12380
rect 3836 11804 3848 12380
rect 3790 11792 3848 11804
rect 4808 12380 4866 12392
rect 4808 11804 4820 12380
rect 4854 11804 4866 12380
rect 4808 11792 4866 11804
rect 5826 12380 5884 12392
rect 5826 11804 5838 12380
rect 5872 11804 5884 12380
rect 5826 11792 5884 11804
rect 6844 12380 6902 12392
rect 6844 11804 6856 12380
rect 6890 11804 6902 12380
rect 6844 11792 6902 11804
rect 7862 12380 7920 12392
rect 7862 11804 7874 12380
rect 7908 11804 7920 12380
rect 7862 11792 7920 11804
rect 8880 12380 8938 12392
rect 8880 11804 8892 12380
rect 8926 11804 8938 12380
rect 8880 11792 8938 11804
rect 9898 12380 9956 12392
rect 9898 11804 9910 12380
rect 9944 11804 9956 12380
rect 9898 11792 9956 11804
rect 10916 12380 10974 12392
rect 10916 11804 10928 12380
rect 10962 11804 10974 12380
rect 10916 11792 10974 11804
rect 13520 12344 13578 12356
rect 13520 11768 13532 12344
rect 13566 11768 13578 12344
rect 13520 11756 13578 11768
rect 14538 12344 14596 12356
rect 14538 11768 14550 12344
rect 14584 11768 14596 12344
rect 14538 11756 14596 11768
rect 15556 12344 15614 12356
rect 15556 11768 15568 12344
rect 15602 11768 15614 12344
rect 15556 11756 15614 11768
rect 16574 12344 16632 12356
rect 16574 11768 16586 12344
rect 16620 11768 16632 12344
rect 16574 11756 16632 11768
rect 17592 12344 17650 12356
rect 17592 11768 17604 12344
rect 17638 11768 17650 12344
rect 17592 11756 17650 11768
rect 18610 12344 18668 12356
rect 18610 11768 18622 12344
rect 18656 11768 18668 12344
rect 18610 11756 18668 11768
rect 19628 12344 19686 12356
rect 19628 11768 19640 12344
rect 19674 11768 19686 12344
rect 19628 11756 19686 11768
rect 20646 12344 20704 12356
rect 20646 11768 20658 12344
rect 20692 11768 20704 12344
rect 20646 11756 20704 11768
rect 21664 12344 21722 12356
rect 21664 11768 21676 12344
rect 21710 11768 21722 12344
rect 21664 11756 21722 11768
rect 22682 12344 22740 12356
rect 22682 11768 22694 12344
rect 22728 11768 22740 12344
rect 22682 11756 22740 11768
rect 23700 12344 23758 12356
rect 23700 11768 23712 12344
rect 23746 11768 23758 12344
rect 23700 11756 23758 11768
rect 24718 12344 24776 12356
rect 24718 11768 24730 12344
rect 24764 11768 24776 12344
rect 24718 11756 24776 11768
rect 25736 12344 25794 12356
rect 25736 11768 25748 12344
rect 25782 11768 25794 12344
rect 25736 11756 25794 11768
rect 26754 12344 26812 12356
rect 26754 11768 26766 12344
rect 26800 11768 26812 12344
rect 26754 11756 26812 11768
rect 27772 12344 27830 12356
rect 27772 11768 27784 12344
rect 27818 11768 27830 12344
rect 27772 11756 27830 11768
rect 28790 12344 28848 12356
rect 28790 11768 28802 12344
rect 28836 11768 28848 12344
rect 28790 11756 28848 11768
rect 29808 12344 29866 12356
rect 29808 11768 29820 12344
rect 29854 11768 29866 12344
rect 29808 11756 29866 11768
rect 30826 12344 30884 12356
rect 30826 11768 30838 12344
rect 30872 11768 30884 12344
rect 30826 11756 30884 11768
rect 31844 12344 31902 12356
rect 31844 11768 31856 12344
rect 31890 11768 31902 12344
rect 31844 11756 31902 11768
rect 32862 12344 32920 12356
rect 32862 11768 32874 12344
rect 32908 11768 32920 12344
rect 32862 11756 32920 11768
rect 33880 12344 33938 12356
rect 33880 11768 33892 12344
rect 33926 11768 33938 12344
rect 33880 11756 33938 11768
rect 1754 11562 1812 11574
rect 1754 10986 1766 11562
rect 1800 10986 1812 11562
rect 1754 10974 1812 10986
rect 2772 11562 2830 11574
rect 2772 10986 2784 11562
rect 2818 10986 2830 11562
rect 2772 10974 2830 10986
rect 3790 11562 3848 11574
rect 3790 10986 3802 11562
rect 3836 10986 3848 11562
rect 3790 10974 3848 10986
rect 4808 11562 4866 11574
rect 4808 10986 4820 11562
rect 4854 10986 4866 11562
rect 4808 10974 4866 10986
rect 5826 11562 5884 11574
rect 5826 10986 5838 11562
rect 5872 10986 5884 11562
rect 5826 10974 5884 10986
rect 6844 11562 6902 11574
rect 6844 10986 6856 11562
rect 6890 10986 6902 11562
rect 6844 10974 6902 10986
rect 7862 11562 7920 11574
rect 7862 10986 7874 11562
rect 7908 10986 7920 11562
rect 7862 10974 7920 10986
rect 8880 11562 8938 11574
rect 8880 10986 8892 11562
rect 8926 10986 8938 11562
rect 8880 10974 8938 10986
rect 9898 11562 9956 11574
rect 9898 10986 9910 11562
rect 9944 10986 9956 11562
rect 9898 10974 9956 10986
rect 10916 11562 10974 11574
rect 10916 10986 10928 11562
rect 10962 10986 10974 11562
rect 10916 10974 10974 10986
rect 13518 11110 13576 11122
rect 1754 10744 1812 10756
rect 1754 10168 1766 10744
rect 1800 10168 1812 10744
rect 1754 10156 1812 10168
rect 2772 10744 2830 10756
rect 2772 10168 2784 10744
rect 2818 10168 2830 10744
rect 2772 10156 2830 10168
rect 3790 10744 3848 10756
rect 3790 10168 3802 10744
rect 3836 10168 3848 10744
rect 3790 10156 3848 10168
rect 4808 10744 4866 10756
rect 4808 10168 4820 10744
rect 4854 10168 4866 10744
rect 4808 10156 4866 10168
rect 5826 10744 5884 10756
rect 5826 10168 5838 10744
rect 5872 10168 5884 10744
rect 5826 10156 5884 10168
rect 6844 10744 6902 10756
rect 6844 10168 6856 10744
rect 6890 10168 6902 10744
rect 6844 10156 6902 10168
rect 7862 10744 7920 10756
rect 7862 10168 7874 10744
rect 7908 10168 7920 10744
rect 7862 10156 7920 10168
rect 8880 10744 8938 10756
rect 8880 10168 8892 10744
rect 8926 10168 8938 10744
rect 8880 10156 8938 10168
rect 9898 10744 9956 10756
rect 9898 10168 9910 10744
rect 9944 10168 9956 10744
rect 9898 10156 9956 10168
rect 10916 10744 10974 10756
rect 10916 10168 10928 10744
rect 10962 10168 10974 10744
rect 13518 10534 13530 11110
rect 13564 10534 13576 11110
rect 13518 10522 13576 10534
rect 14536 11110 14594 11122
rect 14536 10534 14548 11110
rect 14582 10534 14594 11110
rect 14536 10522 14594 10534
rect 15554 11110 15612 11122
rect 15554 10534 15566 11110
rect 15600 10534 15612 11110
rect 15554 10522 15612 10534
rect 16572 11110 16630 11122
rect 16572 10534 16584 11110
rect 16618 10534 16630 11110
rect 16572 10522 16630 10534
rect 17590 11110 17648 11122
rect 17590 10534 17602 11110
rect 17636 10534 17648 11110
rect 17590 10522 17648 10534
rect 18608 11110 18666 11122
rect 18608 10534 18620 11110
rect 18654 10534 18666 11110
rect 18608 10522 18666 10534
rect 19626 11110 19684 11122
rect 19626 10534 19638 11110
rect 19672 10534 19684 11110
rect 19626 10522 19684 10534
rect 20644 11110 20702 11122
rect 20644 10534 20656 11110
rect 20690 10534 20702 11110
rect 20644 10522 20702 10534
rect 21662 11110 21720 11122
rect 21662 10534 21674 11110
rect 21708 10534 21720 11110
rect 21662 10522 21720 10534
rect 22680 11110 22738 11122
rect 22680 10534 22692 11110
rect 22726 10534 22738 11110
rect 22680 10522 22738 10534
rect 23698 11110 23756 11122
rect 23698 10534 23710 11110
rect 23744 10534 23756 11110
rect 23698 10522 23756 10534
rect 24716 11110 24774 11122
rect 24716 10534 24728 11110
rect 24762 10534 24774 11110
rect 24716 10522 24774 10534
rect 25734 11110 25792 11122
rect 25734 10534 25746 11110
rect 25780 10534 25792 11110
rect 25734 10522 25792 10534
rect 26752 11110 26810 11122
rect 26752 10534 26764 11110
rect 26798 10534 26810 11110
rect 26752 10522 26810 10534
rect 27770 11110 27828 11122
rect 27770 10534 27782 11110
rect 27816 10534 27828 11110
rect 27770 10522 27828 10534
rect 28788 11110 28846 11122
rect 28788 10534 28800 11110
rect 28834 10534 28846 11110
rect 28788 10522 28846 10534
rect 29806 11110 29864 11122
rect 29806 10534 29818 11110
rect 29852 10534 29864 11110
rect 29806 10522 29864 10534
rect 30824 11110 30882 11122
rect 30824 10534 30836 11110
rect 30870 10534 30882 11110
rect 30824 10522 30882 10534
rect 31842 11110 31900 11122
rect 31842 10534 31854 11110
rect 31888 10534 31900 11110
rect 31842 10522 31900 10534
rect 32860 11110 32918 11122
rect 32860 10534 32872 11110
rect 32906 10534 32918 11110
rect 32860 10522 32918 10534
rect 33878 11110 33936 11122
rect 33878 10534 33890 11110
rect 33924 10534 33936 11110
rect 33878 10522 33936 10534
rect 10916 10156 10974 10168
rect 1754 9926 1812 9938
rect 1754 9350 1766 9926
rect 1800 9350 1812 9926
rect 1754 9338 1812 9350
rect 2772 9926 2830 9938
rect 2772 9350 2784 9926
rect 2818 9350 2830 9926
rect 2772 9338 2830 9350
rect 3790 9926 3848 9938
rect 3790 9350 3802 9926
rect 3836 9350 3848 9926
rect 3790 9338 3848 9350
rect 4808 9926 4866 9938
rect 4808 9350 4820 9926
rect 4854 9350 4866 9926
rect 4808 9338 4866 9350
rect 5826 9926 5884 9938
rect 5826 9350 5838 9926
rect 5872 9350 5884 9926
rect 5826 9338 5884 9350
rect 6844 9926 6902 9938
rect 6844 9350 6856 9926
rect 6890 9350 6902 9926
rect 6844 9338 6902 9350
rect 7862 9926 7920 9938
rect 7862 9350 7874 9926
rect 7908 9350 7920 9926
rect 7862 9338 7920 9350
rect 8880 9926 8938 9938
rect 8880 9350 8892 9926
rect 8926 9350 8938 9926
rect 8880 9338 8938 9350
rect 9898 9926 9956 9938
rect 9898 9350 9910 9926
rect 9944 9350 9956 9926
rect 9898 9338 9956 9350
rect 10916 9926 10974 9938
rect 10916 9350 10928 9926
rect 10962 9350 10974 9926
rect 10916 9338 10974 9350
rect 13518 9876 13576 9888
rect 13518 9300 13530 9876
rect 13564 9300 13576 9876
rect 13518 9288 13576 9300
rect 14536 9876 14594 9888
rect 14536 9300 14548 9876
rect 14582 9300 14594 9876
rect 14536 9288 14594 9300
rect 15554 9876 15612 9888
rect 15554 9300 15566 9876
rect 15600 9300 15612 9876
rect 15554 9288 15612 9300
rect 16572 9876 16630 9888
rect 16572 9300 16584 9876
rect 16618 9300 16630 9876
rect 16572 9288 16630 9300
rect 17590 9876 17648 9888
rect 17590 9300 17602 9876
rect 17636 9300 17648 9876
rect 17590 9288 17648 9300
rect 18608 9876 18666 9888
rect 18608 9300 18620 9876
rect 18654 9300 18666 9876
rect 18608 9288 18666 9300
rect 19626 9876 19684 9888
rect 19626 9300 19638 9876
rect 19672 9300 19684 9876
rect 19626 9288 19684 9300
rect 20644 9876 20702 9888
rect 20644 9300 20656 9876
rect 20690 9300 20702 9876
rect 20644 9288 20702 9300
rect 21662 9876 21720 9888
rect 21662 9300 21674 9876
rect 21708 9300 21720 9876
rect 21662 9288 21720 9300
rect 22680 9876 22738 9888
rect 22680 9300 22692 9876
rect 22726 9300 22738 9876
rect 22680 9288 22738 9300
rect 23698 9876 23756 9888
rect 23698 9300 23710 9876
rect 23744 9300 23756 9876
rect 23698 9288 23756 9300
rect 24716 9876 24774 9888
rect 24716 9300 24728 9876
rect 24762 9300 24774 9876
rect 24716 9288 24774 9300
rect 25734 9876 25792 9888
rect 25734 9300 25746 9876
rect 25780 9300 25792 9876
rect 25734 9288 25792 9300
rect 26752 9876 26810 9888
rect 26752 9300 26764 9876
rect 26798 9300 26810 9876
rect 26752 9288 26810 9300
rect 27770 9876 27828 9888
rect 27770 9300 27782 9876
rect 27816 9300 27828 9876
rect 27770 9288 27828 9300
rect 28788 9876 28846 9888
rect 28788 9300 28800 9876
rect 28834 9300 28846 9876
rect 28788 9288 28846 9300
rect 29806 9876 29864 9888
rect 29806 9300 29818 9876
rect 29852 9300 29864 9876
rect 29806 9288 29864 9300
rect 30824 9876 30882 9888
rect 30824 9300 30836 9876
rect 30870 9300 30882 9876
rect 30824 9288 30882 9300
rect 31842 9876 31900 9888
rect 31842 9300 31854 9876
rect 31888 9300 31900 9876
rect 31842 9288 31900 9300
rect 32860 9876 32918 9888
rect 32860 9300 32872 9876
rect 32906 9300 32918 9876
rect 32860 9288 32918 9300
rect 33878 9876 33936 9888
rect 33878 9300 33890 9876
rect 33924 9300 33936 9876
rect 33878 9288 33936 9300
rect 1754 9108 1812 9120
rect 1754 8532 1766 9108
rect 1800 8532 1812 9108
rect 1754 8520 1812 8532
rect 2772 9108 2830 9120
rect 2772 8532 2784 9108
rect 2818 8532 2830 9108
rect 2772 8520 2830 8532
rect 3790 9108 3848 9120
rect 3790 8532 3802 9108
rect 3836 8532 3848 9108
rect 3790 8520 3848 8532
rect 4808 9108 4866 9120
rect 4808 8532 4820 9108
rect 4854 8532 4866 9108
rect 4808 8520 4866 8532
rect 5826 9108 5884 9120
rect 5826 8532 5838 9108
rect 5872 8532 5884 9108
rect 5826 8520 5884 8532
rect 6844 9108 6902 9120
rect 6844 8532 6856 9108
rect 6890 8532 6902 9108
rect 6844 8520 6902 8532
rect 7862 9108 7920 9120
rect 7862 8532 7874 9108
rect 7908 8532 7920 9108
rect 7862 8520 7920 8532
rect 8880 9108 8938 9120
rect 8880 8532 8892 9108
rect 8926 8532 8938 9108
rect 8880 8520 8938 8532
rect 9898 9108 9956 9120
rect 9898 8532 9910 9108
rect 9944 8532 9956 9108
rect 9898 8520 9956 8532
rect 10916 9108 10974 9120
rect 10916 8532 10928 9108
rect 10962 8532 10974 9108
rect 10916 8520 10974 8532
rect 13518 8644 13576 8656
rect 1754 8290 1812 8302
rect 1754 7714 1766 8290
rect 1800 7714 1812 8290
rect 1754 7702 1812 7714
rect 2772 8290 2830 8302
rect 2772 7714 2784 8290
rect 2818 7714 2830 8290
rect 2772 7702 2830 7714
rect 3790 8290 3848 8302
rect 3790 7714 3802 8290
rect 3836 7714 3848 8290
rect 3790 7702 3848 7714
rect 4808 8290 4866 8302
rect 4808 7714 4820 8290
rect 4854 7714 4866 8290
rect 4808 7702 4866 7714
rect 5826 8290 5884 8302
rect 5826 7714 5838 8290
rect 5872 7714 5884 8290
rect 5826 7702 5884 7714
rect 6844 8290 6902 8302
rect 6844 7714 6856 8290
rect 6890 7714 6902 8290
rect 6844 7702 6902 7714
rect 7862 8290 7920 8302
rect 7862 7714 7874 8290
rect 7908 7714 7920 8290
rect 7862 7702 7920 7714
rect 8880 8290 8938 8302
rect 8880 7714 8892 8290
rect 8926 7714 8938 8290
rect 8880 7702 8938 7714
rect 9898 8290 9956 8302
rect 9898 7714 9910 8290
rect 9944 7714 9956 8290
rect 9898 7702 9956 7714
rect 10916 8290 10974 8302
rect 10916 7714 10928 8290
rect 10962 7714 10974 8290
rect 13518 8068 13530 8644
rect 13564 8068 13576 8644
rect 13518 8056 13576 8068
rect 14536 8644 14594 8656
rect 14536 8068 14548 8644
rect 14582 8068 14594 8644
rect 14536 8056 14594 8068
rect 15554 8644 15612 8656
rect 15554 8068 15566 8644
rect 15600 8068 15612 8644
rect 15554 8056 15612 8068
rect 16572 8644 16630 8656
rect 16572 8068 16584 8644
rect 16618 8068 16630 8644
rect 16572 8056 16630 8068
rect 17590 8644 17648 8656
rect 17590 8068 17602 8644
rect 17636 8068 17648 8644
rect 17590 8056 17648 8068
rect 18608 8644 18666 8656
rect 18608 8068 18620 8644
rect 18654 8068 18666 8644
rect 18608 8056 18666 8068
rect 19626 8644 19684 8656
rect 19626 8068 19638 8644
rect 19672 8068 19684 8644
rect 19626 8056 19684 8068
rect 20644 8644 20702 8656
rect 20644 8068 20656 8644
rect 20690 8068 20702 8644
rect 20644 8056 20702 8068
rect 21662 8644 21720 8656
rect 21662 8068 21674 8644
rect 21708 8068 21720 8644
rect 21662 8056 21720 8068
rect 22680 8644 22738 8656
rect 22680 8068 22692 8644
rect 22726 8068 22738 8644
rect 22680 8056 22738 8068
rect 23698 8644 23756 8656
rect 23698 8068 23710 8644
rect 23744 8068 23756 8644
rect 23698 8056 23756 8068
rect 24716 8644 24774 8656
rect 24716 8068 24728 8644
rect 24762 8068 24774 8644
rect 24716 8056 24774 8068
rect 25734 8644 25792 8656
rect 25734 8068 25746 8644
rect 25780 8068 25792 8644
rect 25734 8056 25792 8068
rect 26752 8644 26810 8656
rect 26752 8068 26764 8644
rect 26798 8068 26810 8644
rect 26752 8056 26810 8068
rect 27770 8644 27828 8656
rect 27770 8068 27782 8644
rect 27816 8068 27828 8644
rect 27770 8056 27828 8068
rect 28788 8644 28846 8656
rect 28788 8068 28800 8644
rect 28834 8068 28846 8644
rect 28788 8056 28846 8068
rect 29806 8644 29864 8656
rect 29806 8068 29818 8644
rect 29852 8068 29864 8644
rect 29806 8056 29864 8068
rect 30824 8644 30882 8656
rect 30824 8068 30836 8644
rect 30870 8068 30882 8644
rect 30824 8056 30882 8068
rect 31842 8644 31900 8656
rect 31842 8068 31854 8644
rect 31888 8068 31900 8644
rect 31842 8056 31900 8068
rect 32860 8644 32918 8656
rect 32860 8068 32872 8644
rect 32906 8068 32918 8644
rect 32860 8056 32918 8068
rect 33878 8644 33936 8656
rect 33878 8068 33890 8644
rect 33924 8068 33936 8644
rect 33878 8056 33936 8068
rect 10916 7702 10974 7714
rect 13518 7410 13576 7422
rect 8614 6906 8672 6918
rect 8614 6730 8626 6906
rect 8660 6730 8672 6906
rect 8614 6718 8672 6730
rect 8832 6906 8890 6918
rect 8832 6730 8844 6906
rect 8878 6730 8890 6906
rect 8832 6718 8890 6730
rect 9050 6906 9108 6918
rect 9050 6730 9062 6906
rect 9096 6730 9108 6906
rect 9050 6718 9108 6730
rect 9268 6906 9326 6918
rect 9268 6730 9280 6906
rect 9314 6730 9326 6906
rect 9268 6718 9326 6730
rect 9486 6906 9544 6918
rect 9486 6730 9498 6906
rect 9532 6730 9544 6906
rect 9486 6718 9544 6730
rect 9704 6906 9762 6918
rect 9704 6730 9716 6906
rect 9750 6730 9762 6906
rect 9704 6718 9762 6730
rect 9922 6906 9980 6918
rect 9922 6730 9934 6906
rect 9968 6730 9980 6906
rect 9922 6718 9980 6730
rect 10140 6906 10198 6918
rect 10140 6730 10152 6906
rect 10186 6730 10198 6906
rect 10140 6718 10198 6730
rect 10358 6906 10416 6918
rect 10358 6730 10370 6906
rect 10404 6730 10416 6906
rect 10358 6718 10416 6730
rect 10576 6906 10634 6918
rect 10576 6730 10588 6906
rect 10622 6730 10634 6906
rect 10576 6718 10634 6730
rect 10794 6906 10852 6918
rect 10794 6730 10806 6906
rect 10840 6730 10852 6906
rect 13518 6834 13530 7410
rect 13564 6834 13576 7410
rect 13518 6822 13576 6834
rect 14536 7410 14594 7422
rect 14536 6834 14548 7410
rect 14582 6834 14594 7410
rect 14536 6822 14594 6834
rect 15554 7410 15612 7422
rect 15554 6834 15566 7410
rect 15600 6834 15612 7410
rect 15554 6822 15612 6834
rect 16572 7410 16630 7422
rect 16572 6834 16584 7410
rect 16618 6834 16630 7410
rect 16572 6822 16630 6834
rect 17590 7410 17648 7422
rect 17590 6834 17602 7410
rect 17636 6834 17648 7410
rect 17590 6822 17648 6834
rect 18608 7410 18666 7422
rect 18608 6834 18620 7410
rect 18654 6834 18666 7410
rect 18608 6822 18666 6834
rect 19626 7410 19684 7422
rect 19626 6834 19638 7410
rect 19672 6834 19684 7410
rect 19626 6822 19684 6834
rect 20644 7410 20702 7422
rect 20644 6834 20656 7410
rect 20690 6834 20702 7410
rect 20644 6822 20702 6834
rect 21662 7410 21720 7422
rect 21662 6834 21674 7410
rect 21708 6834 21720 7410
rect 21662 6822 21720 6834
rect 22680 7410 22738 7422
rect 22680 6834 22692 7410
rect 22726 6834 22738 7410
rect 22680 6822 22738 6834
rect 23698 7410 23756 7422
rect 23698 6834 23710 7410
rect 23744 6834 23756 7410
rect 23698 6822 23756 6834
rect 24716 7410 24774 7422
rect 24716 6834 24728 7410
rect 24762 6834 24774 7410
rect 24716 6822 24774 6834
rect 25734 7410 25792 7422
rect 25734 6834 25746 7410
rect 25780 6834 25792 7410
rect 25734 6822 25792 6834
rect 26752 7410 26810 7422
rect 26752 6834 26764 7410
rect 26798 6834 26810 7410
rect 26752 6822 26810 6834
rect 27770 7410 27828 7422
rect 27770 6834 27782 7410
rect 27816 6834 27828 7410
rect 27770 6822 27828 6834
rect 28788 7410 28846 7422
rect 28788 6834 28800 7410
rect 28834 6834 28846 7410
rect 28788 6822 28846 6834
rect 29806 7410 29864 7422
rect 29806 6834 29818 7410
rect 29852 6834 29864 7410
rect 29806 6822 29864 6834
rect 30824 7410 30882 7422
rect 30824 6834 30836 7410
rect 30870 6834 30882 7410
rect 30824 6822 30882 6834
rect 31842 7410 31900 7422
rect 31842 6834 31854 7410
rect 31888 6834 31900 7410
rect 31842 6822 31900 6834
rect 32860 7410 32918 7422
rect 32860 6834 32872 7410
rect 32906 6834 32918 7410
rect 32860 6822 32918 6834
rect 33878 7410 33936 7422
rect 33878 6834 33890 7410
rect 33924 6834 33936 7410
rect 33878 6822 33936 6834
rect 10794 6718 10852 6730
rect 13518 6176 13576 6188
rect 8614 6074 8672 6086
rect 8614 5898 8626 6074
rect 8660 5898 8672 6074
rect 8614 5886 8672 5898
rect 8832 6074 8890 6086
rect 8832 5898 8844 6074
rect 8878 5898 8890 6074
rect 8832 5886 8890 5898
rect 9050 6074 9108 6086
rect 9050 5898 9062 6074
rect 9096 5898 9108 6074
rect 9050 5886 9108 5898
rect 9268 6074 9326 6086
rect 9268 5898 9280 6074
rect 9314 5898 9326 6074
rect 9268 5886 9326 5898
rect 9486 6074 9544 6086
rect 9486 5898 9498 6074
rect 9532 5898 9544 6074
rect 9486 5886 9544 5898
rect 9704 6074 9762 6086
rect 9704 5898 9716 6074
rect 9750 5898 9762 6074
rect 9704 5886 9762 5898
rect 9922 6074 9980 6086
rect 9922 5898 9934 6074
rect 9968 5898 9980 6074
rect 9922 5886 9980 5898
rect 10140 6074 10198 6086
rect 10140 5898 10152 6074
rect 10186 5898 10198 6074
rect 10140 5886 10198 5898
rect 10358 6074 10416 6086
rect 10358 5898 10370 6074
rect 10404 5898 10416 6074
rect 10358 5886 10416 5898
rect 10576 6074 10634 6086
rect 10576 5898 10588 6074
rect 10622 5898 10634 6074
rect 10576 5886 10634 5898
rect 10794 6074 10852 6086
rect 10794 5898 10806 6074
rect 10840 5898 10852 6074
rect 10794 5886 10852 5898
rect 13518 5600 13530 6176
rect 13564 5600 13576 6176
rect 13518 5588 13576 5600
rect 14536 6176 14594 6188
rect 14536 5600 14548 6176
rect 14582 5600 14594 6176
rect 14536 5588 14594 5600
rect 15554 6176 15612 6188
rect 15554 5600 15566 6176
rect 15600 5600 15612 6176
rect 15554 5588 15612 5600
rect 16572 6176 16630 6188
rect 16572 5600 16584 6176
rect 16618 5600 16630 6176
rect 16572 5588 16630 5600
rect 17590 6176 17648 6188
rect 17590 5600 17602 6176
rect 17636 5600 17648 6176
rect 17590 5588 17648 5600
rect 18608 6176 18666 6188
rect 18608 5600 18620 6176
rect 18654 5600 18666 6176
rect 18608 5588 18666 5600
rect 19626 6176 19684 6188
rect 19626 5600 19638 6176
rect 19672 5600 19684 6176
rect 19626 5588 19684 5600
rect 20644 6176 20702 6188
rect 20644 5600 20656 6176
rect 20690 5600 20702 6176
rect 20644 5588 20702 5600
rect 21662 6176 21720 6188
rect 21662 5600 21674 6176
rect 21708 5600 21720 6176
rect 21662 5588 21720 5600
rect 22680 6176 22738 6188
rect 22680 5600 22692 6176
rect 22726 5600 22738 6176
rect 22680 5588 22738 5600
rect 23698 6176 23756 6188
rect 23698 5600 23710 6176
rect 23744 5600 23756 6176
rect 23698 5588 23756 5600
rect 24716 6176 24774 6188
rect 24716 5600 24728 6176
rect 24762 5600 24774 6176
rect 24716 5588 24774 5600
rect 25734 6176 25792 6188
rect 25734 5600 25746 6176
rect 25780 5600 25792 6176
rect 25734 5588 25792 5600
rect 26752 6176 26810 6188
rect 26752 5600 26764 6176
rect 26798 5600 26810 6176
rect 26752 5588 26810 5600
rect 27770 6176 27828 6188
rect 27770 5600 27782 6176
rect 27816 5600 27828 6176
rect 27770 5588 27828 5600
rect 28788 6176 28846 6188
rect 28788 5600 28800 6176
rect 28834 5600 28846 6176
rect 28788 5588 28846 5600
rect 29806 6176 29864 6188
rect 29806 5600 29818 6176
rect 29852 5600 29864 6176
rect 29806 5588 29864 5600
rect 30824 6176 30882 6188
rect 30824 5600 30836 6176
rect 30870 5600 30882 6176
rect 30824 5588 30882 5600
rect 31842 6176 31900 6188
rect 31842 5600 31854 6176
rect 31888 5600 31900 6176
rect 31842 5588 31900 5600
rect 32860 6176 32918 6188
rect 32860 5600 32872 6176
rect 32906 5600 32918 6176
rect 32860 5588 32918 5600
rect 33878 6176 33936 6188
rect 33878 5600 33890 6176
rect 33924 5600 33936 6176
rect 33878 5588 33936 5600
rect 13518 4944 13576 4956
rect 1533 4747 1591 4759
rect 1533 4171 1545 4747
rect 1579 4171 1591 4747
rect 1533 4159 1591 4171
rect 2551 4747 2609 4759
rect 2551 4171 2563 4747
rect 2597 4171 2609 4747
rect 2551 4159 2609 4171
rect 3569 4747 3627 4759
rect 3569 4171 3581 4747
rect 3615 4171 3627 4747
rect 3569 4159 3627 4171
rect 4587 4747 4645 4759
rect 4587 4171 4599 4747
rect 4633 4171 4645 4747
rect 4587 4159 4645 4171
rect 5605 4747 5663 4759
rect 5605 4171 5617 4747
rect 5651 4171 5663 4747
rect 5605 4159 5663 4171
rect 6623 4747 6681 4759
rect 6623 4171 6635 4747
rect 6669 4171 6681 4747
rect 6623 4159 6681 4171
rect 7641 4747 7699 4759
rect 7641 4171 7653 4747
rect 7687 4171 7699 4747
rect 7641 4159 7699 4171
rect 8528 4748 8586 4760
rect 8528 4172 8540 4748
rect 8574 4172 8586 4748
rect 8528 4160 8586 4172
rect 8826 4748 8884 4760
rect 8826 4172 8838 4748
rect 8872 4172 8884 4748
rect 8826 4160 8884 4172
rect 9124 4748 9182 4760
rect 9124 4172 9136 4748
rect 9170 4172 9182 4748
rect 9124 4160 9182 4172
rect 9422 4748 9480 4760
rect 9422 4172 9434 4748
rect 9468 4172 9480 4748
rect 9422 4160 9480 4172
rect 9720 4748 9778 4760
rect 9720 4172 9732 4748
rect 9766 4172 9778 4748
rect 9720 4160 9778 4172
rect 10018 4748 10076 4760
rect 10018 4172 10030 4748
rect 10064 4172 10076 4748
rect 10018 4160 10076 4172
rect 10316 4748 10374 4760
rect 10316 4172 10328 4748
rect 10362 4172 10374 4748
rect 10316 4160 10374 4172
rect 10614 4748 10672 4760
rect 10614 4172 10626 4748
rect 10660 4172 10672 4748
rect 10614 4160 10672 4172
rect 10912 4748 10970 4760
rect 10912 4172 10924 4748
rect 10958 4172 10970 4748
rect 10912 4160 10970 4172
rect 11210 4748 11268 4760
rect 11210 4172 11222 4748
rect 11256 4172 11268 4748
rect 11210 4160 11268 4172
rect 11508 4748 11566 4760
rect 11508 4172 11520 4748
rect 11554 4172 11566 4748
rect 11508 4160 11566 4172
rect 11806 4748 11864 4760
rect 11806 4172 11818 4748
rect 11852 4172 11864 4748
rect 13518 4368 13530 4944
rect 13564 4368 13576 4944
rect 13518 4356 13576 4368
rect 14536 4944 14594 4956
rect 14536 4368 14548 4944
rect 14582 4368 14594 4944
rect 14536 4356 14594 4368
rect 15554 4944 15612 4956
rect 15554 4368 15566 4944
rect 15600 4368 15612 4944
rect 15554 4356 15612 4368
rect 16572 4944 16630 4956
rect 16572 4368 16584 4944
rect 16618 4368 16630 4944
rect 16572 4356 16630 4368
rect 17590 4944 17648 4956
rect 17590 4368 17602 4944
rect 17636 4368 17648 4944
rect 17590 4356 17648 4368
rect 18608 4944 18666 4956
rect 18608 4368 18620 4944
rect 18654 4368 18666 4944
rect 18608 4356 18666 4368
rect 19626 4944 19684 4956
rect 19626 4368 19638 4944
rect 19672 4368 19684 4944
rect 19626 4356 19684 4368
rect 20644 4944 20702 4956
rect 20644 4368 20656 4944
rect 20690 4368 20702 4944
rect 20644 4356 20702 4368
rect 21662 4944 21720 4956
rect 21662 4368 21674 4944
rect 21708 4368 21720 4944
rect 21662 4356 21720 4368
rect 22680 4944 22738 4956
rect 22680 4368 22692 4944
rect 22726 4368 22738 4944
rect 22680 4356 22738 4368
rect 23698 4944 23756 4956
rect 23698 4368 23710 4944
rect 23744 4368 23756 4944
rect 23698 4356 23756 4368
rect 24716 4944 24774 4956
rect 24716 4368 24728 4944
rect 24762 4368 24774 4944
rect 24716 4356 24774 4368
rect 25734 4944 25792 4956
rect 25734 4368 25746 4944
rect 25780 4368 25792 4944
rect 25734 4356 25792 4368
rect 26752 4944 26810 4956
rect 26752 4368 26764 4944
rect 26798 4368 26810 4944
rect 26752 4356 26810 4368
rect 27770 4944 27828 4956
rect 27770 4368 27782 4944
rect 27816 4368 27828 4944
rect 27770 4356 27828 4368
rect 28788 4944 28846 4956
rect 28788 4368 28800 4944
rect 28834 4368 28846 4944
rect 28788 4356 28846 4368
rect 29806 4944 29864 4956
rect 29806 4368 29818 4944
rect 29852 4368 29864 4944
rect 29806 4356 29864 4368
rect 30824 4944 30882 4956
rect 30824 4368 30836 4944
rect 30870 4368 30882 4944
rect 30824 4356 30882 4368
rect 31842 4944 31900 4956
rect 31842 4368 31854 4944
rect 31888 4368 31900 4944
rect 31842 4356 31900 4368
rect 32860 4944 32918 4956
rect 32860 4368 32872 4944
rect 32906 4368 32918 4944
rect 32860 4356 32918 4368
rect 33878 4944 33936 4956
rect 33878 4368 33890 4944
rect 33924 4368 33936 4944
rect 33878 4356 33936 4368
rect 11806 4160 11864 4172
rect 13518 3710 13576 3722
rect 1532 3634 1590 3646
rect 1532 3058 1544 3634
rect 1578 3058 1590 3634
rect 1532 3046 1590 3058
rect 2550 3634 2608 3646
rect 2550 3058 2562 3634
rect 2596 3058 2608 3634
rect 2550 3046 2608 3058
rect 3568 3634 3626 3646
rect 3568 3058 3580 3634
rect 3614 3058 3626 3634
rect 3568 3046 3626 3058
rect 4586 3634 4644 3646
rect 4586 3058 4598 3634
rect 4632 3058 4644 3634
rect 4586 3046 4644 3058
rect 5604 3634 5662 3646
rect 5604 3058 5616 3634
rect 5650 3058 5662 3634
rect 5604 3046 5662 3058
rect 6622 3634 6680 3646
rect 6622 3058 6634 3634
rect 6668 3058 6680 3634
rect 6622 3046 6680 3058
rect 7640 3634 7698 3646
rect 7640 3058 7652 3634
rect 7686 3058 7698 3634
rect 7640 3046 7698 3058
rect 8528 3636 8586 3648
rect 8528 3060 8540 3636
rect 8574 3060 8586 3636
rect 8528 3048 8586 3060
rect 8826 3636 8884 3648
rect 8826 3060 8838 3636
rect 8872 3060 8884 3636
rect 8826 3048 8884 3060
rect 9124 3636 9182 3648
rect 9124 3060 9136 3636
rect 9170 3060 9182 3636
rect 9124 3048 9182 3060
rect 9422 3636 9480 3648
rect 9422 3060 9434 3636
rect 9468 3060 9480 3636
rect 9422 3048 9480 3060
rect 9720 3636 9778 3648
rect 9720 3060 9732 3636
rect 9766 3060 9778 3636
rect 9720 3048 9778 3060
rect 10018 3636 10076 3648
rect 10018 3060 10030 3636
rect 10064 3060 10076 3636
rect 10018 3048 10076 3060
rect 10316 3636 10374 3648
rect 10316 3060 10328 3636
rect 10362 3060 10374 3636
rect 10316 3048 10374 3060
rect 10614 3636 10672 3648
rect 10614 3060 10626 3636
rect 10660 3060 10672 3636
rect 10614 3048 10672 3060
rect 10912 3636 10970 3648
rect 10912 3060 10924 3636
rect 10958 3060 10970 3636
rect 10912 3048 10970 3060
rect 11210 3636 11268 3648
rect 11210 3060 11222 3636
rect 11256 3060 11268 3636
rect 11210 3048 11268 3060
rect 11508 3636 11566 3648
rect 11508 3060 11520 3636
rect 11554 3060 11566 3636
rect 11508 3048 11566 3060
rect 11806 3636 11864 3648
rect 11806 3060 11818 3636
rect 11852 3060 11864 3636
rect 13518 3134 13530 3710
rect 13564 3134 13576 3710
rect 13518 3122 13576 3134
rect 14536 3710 14594 3722
rect 14536 3134 14548 3710
rect 14582 3134 14594 3710
rect 14536 3122 14594 3134
rect 15554 3710 15612 3722
rect 15554 3134 15566 3710
rect 15600 3134 15612 3710
rect 15554 3122 15612 3134
rect 16572 3710 16630 3722
rect 16572 3134 16584 3710
rect 16618 3134 16630 3710
rect 16572 3122 16630 3134
rect 17590 3710 17648 3722
rect 17590 3134 17602 3710
rect 17636 3134 17648 3710
rect 17590 3122 17648 3134
rect 18608 3710 18666 3722
rect 18608 3134 18620 3710
rect 18654 3134 18666 3710
rect 18608 3122 18666 3134
rect 19626 3710 19684 3722
rect 19626 3134 19638 3710
rect 19672 3134 19684 3710
rect 19626 3122 19684 3134
rect 20644 3710 20702 3722
rect 20644 3134 20656 3710
rect 20690 3134 20702 3710
rect 20644 3122 20702 3134
rect 21662 3710 21720 3722
rect 21662 3134 21674 3710
rect 21708 3134 21720 3710
rect 21662 3122 21720 3134
rect 22680 3710 22738 3722
rect 22680 3134 22692 3710
rect 22726 3134 22738 3710
rect 22680 3122 22738 3134
rect 23698 3710 23756 3722
rect 23698 3134 23710 3710
rect 23744 3134 23756 3710
rect 23698 3122 23756 3134
rect 24716 3710 24774 3722
rect 24716 3134 24728 3710
rect 24762 3134 24774 3710
rect 24716 3122 24774 3134
rect 25734 3710 25792 3722
rect 25734 3134 25746 3710
rect 25780 3134 25792 3710
rect 25734 3122 25792 3134
rect 26752 3710 26810 3722
rect 26752 3134 26764 3710
rect 26798 3134 26810 3710
rect 26752 3122 26810 3134
rect 27770 3710 27828 3722
rect 27770 3134 27782 3710
rect 27816 3134 27828 3710
rect 27770 3122 27828 3134
rect 28788 3710 28846 3722
rect 28788 3134 28800 3710
rect 28834 3134 28846 3710
rect 28788 3122 28846 3134
rect 29806 3710 29864 3722
rect 29806 3134 29818 3710
rect 29852 3134 29864 3710
rect 29806 3122 29864 3134
rect 30824 3710 30882 3722
rect 30824 3134 30836 3710
rect 30870 3134 30882 3710
rect 30824 3122 30882 3134
rect 31842 3710 31900 3722
rect 31842 3134 31854 3710
rect 31888 3134 31900 3710
rect 31842 3122 31900 3134
rect 32860 3710 32918 3722
rect 32860 3134 32872 3710
rect 32906 3134 32918 3710
rect 32860 3122 32918 3134
rect 33878 3710 33936 3722
rect 33878 3134 33890 3710
rect 33924 3134 33936 3710
rect 33878 3122 33936 3134
rect 11806 3048 11864 3060
rect 1533 2523 1591 2535
rect 1533 1947 1545 2523
rect 1579 1947 1591 2523
rect 1533 1935 1591 1947
rect 2551 2523 2609 2535
rect 2551 1947 2563 2523
rect 2597 1947 2609 2523
rect 2551 1935 2609 1947
rect 3569 2523 3627 2535
rect 3569 1947 3581 2523
rect 3615 1947 3627 2523
rect 3569 1935 3627 1947
rect 4587 2523 4645 2535
rect 4587 1947 4599 2523
rect 4633 1947 4645 2523
rect 4587 1935 4645 1947
rect 5605 2523 5663 2535
rect 5605 1947 5617 2523
rect 5651 1947 5663 2523
rect 5605 1935 5663 1947
rect 6623 2523 6681 2535
rect 6623 1947 6635 2523
rect 6669 1947 6681 2523
rect 6623 1935 6681 1947
rect 7641 2523 7699 2535
rect 7641 1947 7653 2523
rect 7687 1947 7699 2523
rect 7641 1935 7699 1947
rect 8526 2524 8584 2536
rect 8526 1948 8538 2524
rect 8572 1948 8584 2524
rect 8526 1936 8584 1948
rect 8824 2524 8882 2536
rect 8824 1948 8836 2524
rect 8870 1948 8882 2524
rect 8824 1936 8882 1948
rect 9122 2524 9180 2536
rect 9122 1948 9134 2524
rect 9168 1948 9180 2524
rect 9122 1936 9180 1948
rect 9420 2524 9478 2536
rect 9420 1948 9432 2524
rect 9466 1948 9478 2524
rect 9420 1936 9478 1948
rect 9718 2524 9776 2536
rect 9718 1948 9730 2524
rect 9764 1948 9776 2524
rect 9718 1936 9776 1948
rect 10016 2524 10074 2536
rect 10016 1948 10028 2524
rect 10062 1948 10074 2524
rect 10016 1936 10074 1948
rect 10314 2524 10372 2536
rect 10314 1948 10326 2524
rect 10360 1948 10372 2524
rect 10314 1936 10372 1948
rect 10612 2524 10670 2536
rect 10612 1948 10624 2524
rect 10658 1948 10670 2524
rect 10612 1936 10670 1948
rect 10910 2524 10968 2536
rect 10910 1948 10922 2524
rect 10956 1948 10968 2524
rect 10910 1936 10968 1948
rect 11208 2524 11266 2536
rect 11208 1948 11220 2524
rect 11254 1948 11266 2524
rect 11208 1936 11266 1948
rect 11506 2524 11564 2536
rect 11506 1948 11518 2524
rect 11552 1948 11564 2524
rect 11506 1936 11564 1948
rect 11804 2524 11862 2536
rect 11804 1948 11816 2524
rect 11850 1948 11862 2524
rect 11804 1936 11862 1948
rect 13518 2476 13576 2488
rect 13518 1900 13530 2476
rect 13564 1900 13576 2476
rect 13518 1888 13576 1900
rect 14536 2476 14594 2488
rect 14536 1900 14548 2476
rect 14582 1900 14594 2476
rect 14536 1888 14594 1900
rect 15554 2476 15612 2488
rect 15554 1900 15566 2476
rect 15600 1900 15612 2476
rect 15554 1888 15612 1900
rect 16572 2476 16630 2488
rect 16572 1900 16584 2476
rect 16618 1900 16630 2476
rect 16572 1888 16630 1900
rect 17590 2476 17648 2488
rect 17590 1900 17602 2476
rect 17636 1900 17648 2476
rect 17590 1888 17648 1900
rect 18608 2476 18666 2488
rect 18608 1900 18620 2476
rect 18654 1900 18666 2476
rect 18608 1888 18666 1900
rect 19626 2476 19684 2488
rect 19626 1900 19638 2476
rect 19672 1900 19684 2476
rect 19626 1888 19684 1900
rect 20644 2476 20702 2488
rect 20644 1900 20656 2476
rect 20690 1900 20702 2476
rect 20644 1888 20702 1900
rect 21662 2476 21720 2488
rect 21662 1900 21674 2476
rect 21708 1900 21720 2476
rect 21662 1888 21720 1900
rect 22680 2476 22738 2488
rect 22680 1900 22692 2476
rect 22726 1900 22738 2476
rect 22680 1888 22738 1900
rect 23698 2476 23756 2488
rect 23698 1900 23710 2476
rect 23744 1900 23756 2476
rect 23698 1888 23756 1900
rect 24716 2476 24774 2488
rect 24716 1900 24728 2476
rect 24762 1900 24774 2476
rect 24716 1888 24774 1900
rect 25734 2476 25792 2488
rect 25734 1900 25746 2476
rect 25780 1900 25792 2476
rect 25734 1888 25792 1900
rect 26752 2476 26810 2488
rect 26752 1900 26764 2476
rect 26798 1900 26810 2476
rect 26752 1888 26810 1900
rect 27770 2476 27828 2488
rect 27770 1900 27782 2476
rect 27816 1900 27828 2476
rect 27770 1888 27828 1900
rect 28788 2476 28846 2488
rect 28788 1900 28800 2476
rect 28834 1900 28846 2476
rect 28788 1888 28846 1900
rect 29806 2476 29864 2488
rect 29806 1900 29818 2476
rect 29852 1900 29864 2476
rect 29806 1888 29864 1900
rect 30824 2476 30882 2488
rect 30824 1900 30836 2476
rect 30870 1900 30882 2476
rect 30824 1888 30882 1900
rect 31842 2476 31900 2488
rect 31842 1900 31854 2476
rect 31888 1900 31900 2476
rect 31842 1888 31900 1900
rect 32860 2476 32918 2488
rect 32860 1900 32872 2476
rect 32906 1900 32918 2476
rect 32860 1888 32918 1900
rect 33878 2476 33936 2488
rect 33878 1900 33890 2476
rect 33924 1900 33936 2476
rect 33878 1888 33936 1900
rect 1532 1410 1590 1422
rect 1532 834 1544 1410
rect 1578 834 1590 1410
rect 1532 822 1590 834
rect 2550 1410 2608 1422
rect 2550 834 2562 1410
rect 2596 834 2608 1410
rect 2550 822 2608 834
rect 3568 1410 3626 1422
rect 3568 834 3580 1410
rect 3614 834 3626 1410
rect 3568 822 3626 834
rect 4586 1410 4644 1422
rect 4586 834 4598 1410
rect 4632 834 4644 1410
rect 4586 822 4644 834
rect 5604 1410 5662 1422
rect 5604 834 5616 1410
rect 5650 834 5662 1410
rect 5604 822 5662 834
rect 6622 1410 6680 1422
rect 6622 834 6634 1410
rect 6668 834 6680 1410
rect 6622 822 6680 834
rect 7640 1410 7698 1422
rect 7640 834 7652 1410
rect 7686 834 7698 1410
rect 7640 822 7698 834
rect 8526 1414 8584 1426
rect 8526 838 8538 1414
rect 8572 838 8584 1414
rect 8526 826 8584 838
rect 8824 1414 8882 1426
rect 8824 838 8836 1414
rect 8870 838 8882 1414
rect 8824 826 8882 838
rect 9122 1414 9180 1426
rect 9122 838 9134 1414
rect 9168 838 9180 1414
rect 9122 826 9180 838
rect 9420 1414 9478 1426
rect 9420 838 9432 1414
rect 9466 838 9478 1414
rect 9420 826 9478 838
rect 9718 1414 9776 1426
rect 9718 838 9730 1414
rect 9764 838 9776 1414
rect 9718 826 9776 838
rect 10016 1414 10074 1426
rect 10016 838 10028 1414
rect 10062 838 10074 1414
rect 10016 826 10074 838
rect 10314 1414 10372 1426
rect 10314 838 10326 1414
rect 10360 838 10372 1414
rect 10314 826 10372 838
rect 10612 1414 10670 1426
rect 10612 838 10624 1414
rect 10658 838 10670 1414
rect 10612 826 10670 838
rect 10910 1414 10968 1426
rect 10910 838 10922 1414
rect 10956 838 10968 1414
rect 10910 826 10968 838
rect 11208 1414 11266 1426
rect 11208 838 11220 1414
rect 11254 838 11266 1414
rect 11208 826 11266 838
rect 11506 1414 11564 1426
rect 11506 838 11518 1414
rect 11552 838 11564 1414
rect 11506 826 11564 838
rect 11804 1414 11862 1426
rect 11804 838 11816 1414
rect 11850 838 11862 1414
rect 11804 826 11862 838
rect 13518 1244 13576 1256
rect 13518 668 13530 1244
rect 13564 668 13576 1244
rect 13518 656 13576 668
rect 14536 1244 14594 1256
rect 14536 668 14548 1244
rect 14582 668 14594 1244
rect 14536 656 14594 668
rect 15554 1244 15612 1256
rect 15554 668 15566 1244
rect 15600 668 15612 1244
rect 15554 656 15612 668
rect 16572 1244 16630 1256
rect 16572 668 16584 1244
rect 16618 668 16630 1244
rect 16572 656 16630 668
rect 17590 1244 17648 1256
rect 17590 668 17602 1244
rect 17636 668 17648 1244
rect 17590 656 17648 668
rect 18608 1244 18666 1256
rect 18608 668 18620 1244
rect 18654 668 18666 1244
rect 18608 656 18666 668
rect 19626 1244 19684 1256
rect 19626 668 19638 1244
rect 19672 668 19684 1244
rect 19626 656 19684 668
rect 20644 1244 20702 1256
rect 20644 668 20656 1244
rect 20690 668 20702 1244
rect 20644 656 20702 668
rect 21662 1244 21720 1256
rect 21662 668 21674 1244
rect 21708 668 21720 1244
rect 21662 656 21720 668
rect 22680 1244 22738 1256
rect 22680 668 22692 1244
rect 22726 668 22738 1244
rect 22680 656 22738 668
rect 23698 1244 23756 1256
rect 23698 668 23710 1244
rect 23744 668 23756 1244
rect 23698 656 23756 668
rect 24716 1244 24774 1256
rect 24716 668 24728 1244
rect 24762 668 24774 1244
rect 24716 656 24774 668
rect 25734 1244 25792 1256
rect 25734 668 25746 1244
rect 25780 668 25792 1244
rect 25734 656 25792 668
rect 26752 1244 26810 1256
rect 26752 668 26764 1244
rect 26798 668 26810 1244
rect 26752 656 26810 668
rect 27770 1244 27828 1256
rect 27770 668 27782 1244
rect 27816 668 27828 1244
rect 27770 656 27828 668
rect 28788 1244 28846 1256
rect 28788 668 28800 1244
rect 28834 668 28846 1244
rect 28788 656 28846 668
rect 29806 1244 29864 1256
rect 29806 668 29818 1244
rect 29852 668 29864 1244
rect 29806 656 29864 668
rect 30824 1244 30882 1256
rect 30824 668 30836 1244
rect 30870 668 30882 1244
rect 30824 656 30882 668
rect 31842 1244 31900 1256
rect 31842 668 31854 1244
rect 31888 668 31900 1244
rect 31842 656 31900 668
rect 32860 1244 32918 1256
rect 32860 668 32872 1244
rect 32906 668 32918 1244
rect 32860 656 32918 668
rect 33878 1244 33936 1256
rect 33878 668 33890 1244
rect 33924 668 33936 1244
rect 33878 656 33936 668
rect 50648 7549 50700 7561
rect 50648 7515 50656 7549
rect 50690 7515 50700 7549
rect 50648 7481 50700 7515
rect 50648 7447 50656 7481
rect 50690 7447 50700 7481
rect 50648 7431 50700 7447
rect 50730 7549 50782 7561
rect 50730 7515 50740 7549
rect 50774 7515 50782 7549
rect 50730 7481 50782 7515
rect 50730 7447 50740 7481
rect 50774 7447 50782 7481
rect 50730 7431 50782 7447
rect 48792 7328 48850 7340
rect 48792 7152 48804 7328
rect 48838 7152 48850 7328
rect 48792 7140 48850 7152
rect 49050 7328 49108 7340
rect 49050 7152 49062 7328
rect 49096 7152 49108 7328
rect 49050 7140 49108 7152
rect 49308 7328 49366 7340
rect 49308 7152 49320 7328
rect 49354 7152 49366 7328
rect 49308 7140 49366 7152
rect 49566 7328 49624 7340
rect 49566 7152 49578 7328
rect 49612 7152 49624 7328
rect 49566 7140 49624 7152
rect 49824 7328 49882 7340
rect 49824 7152 49836 7328
rect 49870 7152 49882 7328
rect 49824 7140 49882 7152
rect 50082 7328 50140 7340
rect 50082 7152 50094 7328
rect 50128 7152 50140 7328
rect 50082 7140 50140 7152
rect 50340 7328 50398 7340
rect 50340 7152 50352 7328
rect 50386 7152 50398 7328
rect 50340 7140 50398 7152
rect 50648 5585 50700 5597
rect 50648 5551 50656 5585
rect 50690 5551 50700 5585
rect 50648 5517 50700 5551
rect 50648 5483 50656 5517
rect 50690 5483 50700 5517
rect 50648 5467 50700 5483
rect 50730 5585 50782 5597
rect 50730 5551 50740 5585
rect 50774 5551 50782 5585
rect 50730 5517 50782 5551
rect 50730 5483 50740 5517
rect 50774 5483 50782 5517
rect 50730 5467 50782 5483
rect 48792 5364 48850 5376
rect 48792 5188 48804 5364
rect 48838 5188 48850 5364
rect 48792 5176 48850 5188
rect 49050 5364 49108 5376
rect 49050 5188 49062 5364
rect 49096 5188 49108 5364
rect 49050 5176 49108 5188
rect 49308 5364 49366 5376
rect 49308 5188 49320 5364
rect 49354 5188 49366 5364
rect 49308 5176 49366 5188
rect 49566 5364 49624 5376
rect 49566 5188 49578 5364
rect 49612 5188 49624 5364
rect 49566 5176 49624 5188
rect 49824 5364 49882 5376
rect 49824 5188 49836 5364
rect 49870 5188 49882 5364
rect 49824 5176 49882 5188
rect 50082 5364 50140 5376
rect 50082 5188 50094 5364
rect 50128 5188 50140 5364
rect 50082 5176 50140 5188
rect 50340 5364 50398 5376
rect 50340 5188 50352 5364
rect 50386 5188 50398 5364
rect 50340 5176 50398 5188
rect 50648 3585 50700 3597
rect 50648 3551 50656 3585
rect 50690 3551 50700 3585
rect 50648 3517 50700 3551
rect 50648 3483 50656 3517
rect 50690 3483 50700 3517
rect 50648 3467 50700 3483
rect 50730 3585 50782 3597
rect 50730 3551 50740 3585
rect 50774 3551 50782 3585
rect 50730 3517 50782 3551
rect 50730 3483 50740 3517
rect 50774 3483 50782 3517
rect 50730 3467 50782 3483
rect 48792 3364 48850 3376
rect 48792 3188 48804 3364
rect 48838 3188 48850 3364
rect 48792 3176 48850 3188
rect 49050 3364 49108 3376
rect 49050 3188 49062 3364
rect 49096 3188 49108 3364
rect 49050 3176 49108 3188
rect 49308 3364 49366 3376
rect 49308 3188 49320 3364
rect 49354 3188 49366 3364
rect 49308 3176 49366 3188
rect 49566 3364 49624 3376
rect 49566 3188 49578 3364
rect 49612 3188 49624 3364
rect 49566 3176 49624 3188
rect 49824 3364 49882 3376
rect 49824 3188 49836 3364
rect 49870 3188 49882 3364
rect 49824 3176 49882 3188
rect 50082 3364 50140 3376
rect 50082 3188 50094 3364
rect 50128 3188 50140 3364
rect 50082 3176 50140 3188
rect 50340 3364 50398 3376
rect 50340 3188 50352 3364
rect 50386 3188 50398 3364
rect 50340 3176 50398 3188
rect 50648 1495 50700 1507
rect 50648 1461 50656 1495
rect 50690 1461 50700 1495
rect 50648 1427 50700 1461
rect 50648 1393 50656 1427
rect 50690 1393 50700 1427
rect 50648 1377 50700 1393
rect 50730 1495 50782 1507
rect 50730 1461 50740 1495
rect 50774 1461 50782 1495
rect 50730 1427 50782 1461
rect 50730 1393 50740 1427
rect 50774 1393 50782 1427
rect 50730 1377 50782 1393
rect 48792 1274 48850 1286
rect 48792 1098 48804 1274
rect 48838 1098 48850 1274
rect 48792 1086 48850 1098
rect 49050 1274 49108 1286
rect 49050 1098 49062 1274
rect 49096 1098 49108 1274
rect 49050 1086 49108 1098
rect 49308 1274 49366 1286
rect 49308 1098 49320 1274
rect 49354 1098 49366 1274
rect 49308 1086 49366 1098
rect 49566 1274 49624 1286
rect 49566 1098 49578 1274
rect 49612 1098 49624 1274
rect 49566 1086 49624 1098
rect 49824 1274 49882 1286
rect 49824 1098 49836 1274
rect 49870 1098 49882 1274
rect 49824 1086 49882 1098
rect 50082 1274 50140 1286
rect 50082 1098 50094 1274
rect 50128 1098 50140 1274
rect 50082 1086 50140 1098
rect 50340 1274 50398 1286
rect 50340 1098 50352 1274
rect 50386 1098 50398 1274
rect 50340 1086 50398 1098
rect 67520 14810 67578 14822
rect 67520 14234 67532 14810
rect 67566 14234 67578 14810
rect 67520 14222 67578 14234
rect 68538 14810 68596 14822
rect 68538 14234 68550 14810
rect 68584 14234 68596 14810
rect 68538 14222 68596 14234
rect 69556 14810 69614 14822
rect 69556 14234 69568 14810
rect 69602 14234 69614 14810
rect 69556 14222 69614 14234
rect 70574 14810 70632 14822
rect 70574 14234 70586 14810
rect 70620 14234 70632 14810
rect 70574 14222 70632 14234
rect 71592 14810 71650 14822
rect 71592 14234 71604 14810
rect 71638 14234 71650 14810
rect 71592 14222 71650 14234
rect 72610 14810 72668 14822
rect 72610 14234 72622 14810
rect 72656 14234 72668 14810
rect 72610 14222 72668 14234
rect 73628 14810 73686 14822
rect 73628 14234 73640 14810
rect 73674 14234 73686 14810
rect 73628 14222 73686 14234
rect 74646 14810 74704 14822
rect 74646 14234 74658 14810
rect 74692 14234 74704 14810
rect 74646 14222 74704 14234
rect 75664 14810 75722 14822
rect 75664 14234 75676 14810
rect 75710 14234 75722 14810
rect 75664 14222 75722 14234
rect 76682 14810 76740 14822
rect 76682 14234 76694 14810
rect 76728 14234 76740 14810
rect 76682 14222 76740 14234
rect 77700 14810 77758 14822
rect 77700 14234 77712 14810
rect 77746 14234 77758 14810
rect 77700 14222 77758 14234
rect 78718 14810 78776 14822
rect 78718 14234 78730 14810
rect 78764 14234 78776 14810
rect 78718 14222 78776 14234
rect 79736 14810 79794 14822
rect 79736 14234 79748 14810
rect 79782 14234 79794 14810
rect 79736 14222 79794 14234
rect 80754 14810 80812 14822
rect 80754 14234 80766 14810
rect 80800 14234 80812 14810
rect 80754 14222 80812 14234
rect 81772 14810 81830 14822
rect 81772 14234 81784 14810
rect 81818 14234 81830 14810
rect 81772 14222 81830 14234
rect 82790 14810 82848 14822
rect 82790 14234 82802 14810
rect 82836 14234 82848 14810
rect 82790 14222 82848 14234
rect 83808 14810 83866 14822
rect 83808 14234 83820 14810
rect 83854 14234 83866 14810
rect 83808 14222 83866 14234
rect 84826 14810 84884 14822
rect 84826 14234 84838 14810
rect 84872 14234 84884 14810
rect 84826 14222 84884 14234
rect 85844 14810 85902 14822
rect 85844 14234 85856 14810
rect 85890 14234 85902 14810
rect 85844 14222 85902 14234
rect 86862 14810 86920 14822
rect 86862 14234 86874 14810
rect 86908 14234 86920 14810
rect 86862 14222 86920 14234
rect 87880 14810 87938 14822
rect 87880 14234 87892 14810
rect 87926 14234 87938 14810
rect 87880 14222 87938 14234
rect 55754 14016 55812 14028
rect 55754 13440 55766 14016
rect 55800 13440 55812 14016
rect 55754 13428 55812 13440
rect 56772 14016 56830 14028
rect 56772 13440 56784 14016
rect 56818 13440 56830 14016
rect 56772 13428 56830 13440
rect 57790 14016 57848 14028
rect 57790 13440 57802 14016
rect 57836 13440 57848 14016
rect 57790 13428 57848 13440
rect 58808 14016 58866 14028
rect 58808 13440 58820 14016
rect 58854 13440 58866 14016
rect 58808 13428 58866 13440
rect 59826 14016 59884 14028
rect 59826 13440 59838 14016
rect 59872 13440 59884 14016
rect 59826 13428 59884 13440
rect 60844 14016 60902 14028
rect 60844 13440 60856 14016
rect 60890 13440 60902 14016
rect 60844 13428 60902 13440
rect 61862 14016 61920 14028
rect 61862 13440 61874 14016
rect 61908 13440 61920 14016
rect 61862 13428 61920 13440
rect 62880 14016 62938 14028
rect 62880 13440 62892 14016
rect 62926 13440 62938 14016
rect 62880 13428 62938 13440
rect 63898 14016 63956 14028
rect 63898 13440 63910 14016
rect 63944 13440 63956 14016
rect 63898 13428 63956 13440
rect 64916 14016 64974 14028
rect 64916 13440 64928 14016
rect 64962 13440 64974 14016
rect 64916 13428 64974 13440
rect 67520 13576 67578 13588
rect 55754 13198 55812 13210
rect 55754 12622 55766 13198
rect 55800 12622 55812 13198
rect 55754 12610 55812 12622
rect 56772 13198 56830 13210
rect 56772 12622 56784 13198
rect 56818 12622 56830 13198
rect 56772 12610 56830 12622
rect 57790 13198 57848 13210
rect 57790 12622 57802 13198
rect 57836 12622 57848 13198
rect 57790 12610 57848 12622
rect 58808 13198 58866 13210
rect 58808 12622 58820 13198
rect 58854 12622 58866 13198
rect 58808 12610 58866 12622
rect 59826 13198 59884 13210
rect 59826 12622 59838 13198
rect 59872 12622 59884 13198
rect 59826 12610 59884 12622
rect 60844 13198 60902 13210
rect 60844 12622 60856 13198
rect 60890 12622 60902 13198
rect 60844 12610 60902 12622
rect 61862 13198 61920 13210
rect 61862 12622 61874 13198
rect 61908 12622 61920 13198
rect 61862 12610 61920 12622
rect 62880 13198 62938 13210
rect 62880 12622 62892 13198
rect 62926 12622 62938 13198
rect 62880 12610 62938 12622
rect 63898 13198 63956 13210
rect 63898 12622 63910 13198
rect 63944 12622 63956 13198
rect 63898 12610 63956 12622
rect 64916 13198 64974 13210
rect 64916 12622 64928 13198
rect 64962 12622 64974 13198
rect 67520 13000 67532 13576
rect 67566 13000 67578 13576
rect 67520 12988 67578 13000
rect 68538 13576 68596 13588
rect 68538 13000 68550 13576
rect 68584 13000 68596 13576
rect 68538 12988 68596 13000
rect 69556 13576 69614 13588
rect 69556 13000 69568 13576
rect 69602 13000 69614 13576
rect 69556 12988 69614 13000
rect 70574 13576 70632 13588
rect 70574 13000 70586 13576
rect 70620 13000 70632 13576
rect 70574 12988 70632 13000
rect 71592 13576 71650 13588
rect 71592 13000 71604 13576
rect 71638 13000 71650 13576
rect 71592 12988 71650 13000
rect 72610 13576 72668 13588
rect 72610 13000 72622 13576
rect 72656 13000 72668 13576
rect 72610 12988 72668 13000
rect 73628 13576 73686 13588
rect 73628 13000 73640 13576
rect 73674 13000 73686 13576
rect 73628 12988 73686 13000
rect 74646 13576 74704 13588
rect 74646 13000 74658 13576
rect 74692 13000 74704 13576
rect 74646 12988 74704 13000
rect 75664 13576 75722 13588
rect 75664 13000 75676 13576
rect 75710 13000 75722 13576
rect 75664 12988 75722 13000
rect 76682 13576 76740 13588
rect 76682 13000 76694 13576
rect 76728 13000 76740 13576
rect 76682 12988 76740 13000
rect 77700 13576 77758 13588
rect 77700 13000 77712 13576
rect 77746 13000 77758 13576
rect 77700 12988 77758 13000
rect 78718 13576 78776 13588
rect 78718 13000 78730 13576
rect 78764 13000 78776 13576
rect 78718 12988 78776 13000
rect 79736 13576 79794 13588
rect 79736 13000 79748 13576
rect 79782 13000 79794 13576
rect 79736 12988 79794 13000
rect 80754 13576 80812 13588
rect 80754 13000 80766 13576
rect 80800 13000 80812 13576
rect 80754 12988 80812 13000
rect 81772 13576 81830 13588
rect 81772 13000 81784 13576
rect 81818 13000 81830 13576
rect 81772 12988 81830 13000
rect 82790 13576 82848 13588
rect 82790 13000 82802 13576
rect 82836 13000 82848 13576
rect 82790 12988 82848 13000
rect 83808 13576 83866 13588
rect 83808 13000 83820 13576
rect 83854 13000 83866 13576
rect 83808 12988 83866 13000
rect 84826 13576 84884 13588
rect 84826 13000 84838 13576
rect 84872 13000 84884 13576
rect 84826 12988 84884 13000
rect 85844 13576 85902 13588
rect 85844 13000 85856 13576
rect 85890 13000 85902 13576
rect 85844 12988 85902 13000
rect 86862 13576 86920 13588
rect 86862 13000 86874 13576
rect 86908 13000 86920 13576
rect 86862 12988 86920 13000
rect 87880 13576 87938 13588
rect 87880 13000 87892 13576
rect 87926 13000 87938 13576
rect 87880 12988 87938 13000
rect 64916 12610 64974 12622
rect 55754 12380 55812 12392
rect 55754 11804 55766 12380
rect 55800 11804 55812 12380
rect 55754 11792 55812 11804
rect 56772 12380 56830 12392
rect 56772 11804 56784 12380
rect 56818 11804 56830 12380
rect 56772 11792 56830 11804
rect 57790 12380 57848 12392
rect 57790 11804 57802 12380
rect 57836 11804 57848 12380
rect 57790 11792 57848 11804
rect 58808 12380 58866 12392
rect 58808 11804 58820 12380
rect 58854 11804 58866 12380
rect 58808 11792 58866 11804
rect 59826 12380 59884 12392
rect 59826 11804 59838 12380
rect 59872 11804 59884 12380
rect 59826 11792 59884 11804
rect 60844 12380 60902 12392
rect 60844 11804 60856 12380
rect 60890 11804 60902 12380
rect 60844 11792 60902 11804
rect 61862 12380 61920 12392
rect 61862 11804 61874 12380
rect 61908 11804 61920 12380
rect 61862 11792 61920 11804
rect 62880 12380 62938 12392
rect 62880 11804 62892 12380
rect 62926 11804 62938 12380
rect 62880 11792 62938 11804
rect 63898 12380 63956 12392
rect 63898 11804 63910 12380
rect 63944 11804 63956 12380
rect 63898 11792 63956 11804
rect 64916 12380 64974 12392
rect 64916 11804 64928 12380
rect 64962 11804 64974 12380
rect 64916 11792 64974 11804
rect 67520 12344 67578 12356
rect 67520 11768 67532 12344
rect 67566 11768 67578 12344
rect 67520 11756 67578 11768
rect 68538 12344 68596 12356
rect 68538 11768 68550 12344
rect 68584 11768 68596 12344
rect 68538 11756 68596 11768
rect 69556 12344 69614 12356
rect 69556 11768 69568 12344
rect 69602 11768 69614 12344
rect 69556 11756 69614 11768
rect 70574 12344 70632 12356
rect 70574 11768 70586 12344
rect 70620 11768 70632 12344
rect 70574 11756 70632 11768
rect 71592 12344 71650 12356
rect 71592 11768 71604 12344
rect 71638 11768 71650 12344
rect 71592 11756 71650 11768
rect 72610 12344 72668 12356
rect 72610 11768 72622 12344
rect 72656 11768 72668 12344
rect 72610 11756 72668 11768
rect 73628 12344 73686 12356
rect 73628 11768 73640 12344
rect 73674 11768 73686 12344
rect 73628 11756 73686 11768
rect 74646 12344 74704 12356
rect 74646 11768 74658 12344
rect 74692 11768 74704 12344
rect 74646 11756 74704 11768
rect 75664 12344 75722 12356
rect 75664 11768 75676 12344
rect 75710 11768 75722 12344
rect 75664 11756 75722 11768
rect 76682 12344 76740 12356
rect 76682 11768 76694 12344
rect 76728 11768 76740 12344
rect 76682 11756 76740 11768
rect 77700 12344 77758 12356
rect 77700 11768 77712 12344
rect 77746 11768 77758 12344
rect 77700 11756 77758 11768
rect 78718 12344 78776 12356
rect 78718 11768 78730 12344
rect 78764 11768 78776 12344
rect 78718 11756 78776 11768
rect 79736 12344 79794 12356
rect 79736 11768 79748 12344
rect 79782 11768 79794 12344
rect 79736 11756 79794 11768
rect 80754 12344 80812 12356
rect 80754 11768 80766 12344
rect 80800 11768 80812 12344
rect 80754 11756 80812 11768
rect 81772 12344 81830 12356
rect 81772 11768 81784 12344
rect 81818 11768 81830 12344
rect 81772 11756 81830 11768
rect 82790 12344 82848 12356
rect 82790 11768 82802 12344
rect 82836 11768 82848 12344
rect 82790 11756 82848 11768
rect 83808 12344 83866 12356
rect 83808 11768 83820 12344
rect 83854 11768 83866 12344
rect 83808 11756 83866 11768
rect 84826 12344 84884 12356
rect 84826 11768 84838 12344
rect 84872 11768 84884 12344
rect 84826 11756 84884 11768
rect 85844 12344 85902 12356
rect 85844 11768 85856 12344
rect 85890 11768 85902 12344
rect 85844 11756 85902 11768
rect 86862 12344 86920 12356
rect 86862 11768 86874 12344
rect 86908 11768 86920 12344
rect 86862 11756 86920 11768
rect 87880 12344 87938 12356
rect 87880 11768 87892 12344
rect 87926 11768 87938 12344
rect 87880 11756 87938 11768
rect 55754 11562 55812 11574
rect 55754 10986 55766 11562
rect 55800 10986 55812 11562
rect 55754 10974 55812 10986
rect 56772 11562 56830 11574
rect 56772 10986 56784 11562
rect 56818 10986 56830 11562
rect 56772 10974 56830 10986
rect 57790 11562 57848 11574
rect 57790 10986 57802 11562
rect 57836 10986 57848 11562
rect 57790 10974 57848 10986
rect 58808 11562 58866 11574
rect 58808 10986 58820 11562
rect 58854 10986 58866 11562
rect 58808 10974 58866 10986
rect 59826 11562 59884 11574
rect 59826 10986 59838 11562
rect 59872 10986 59884 11562
rect 59826 10974 59884 10986
rect 60844 11562 60902 11574
rect 60844 10986 60856 11562
rect 60890 10986 60902 11562
rect 60844 10974 60902 10986
rect 61862 11562 61920 11574
rect 61862 10986 61874 11562
rect 61908 10986 61920 11562
rect 61862 10974 61920 10986
rect 62880 11562 62938 11574
rect 62880 10986 62892 11562
rect 62926 10986 62938 11562
rect 62880 10974 62938 10986
rect 63898 11562 63956 11574
rect 63898 10986 63910 11562
rect 63944 10986 63956 11562
rect 63898 10974 63956 10986
rect 64916 11562 64974 11574
rect 64916 10986 64928 11562
rect 64962 10986 64974 11562
rect 64916 10974 64974 10986
rect 67518 11110 67576 11122
rect 55754 10744 55812 10756
rect 55754 10168 55766 10744
rect 55800 10168 55812 10744
rect 55754 10156 55812 10168
rect 56772 10744 56830 10756
rect 56772 10168 56784 10744
rect 56818 10168 56830 10744
rect 56772 10156 56830 10168
rect 57790 10744 57848 10756
rect 57790 10168 57802 10744
rect 57836 10168 57848 10744
rect 57790 10156 57848 10168
rect 58808 10744 58866 10756
rect 58808 10168 58820 10744
rect 58854 10168 58866 10744
rect 58808 10156 58866 10168
rect 59826 10744 59884 10756
rect 59826 10168 59838 10744
rect 59872 10168 59884 10744
rect 59826 10156 59884 10168
rect 60844 10744 60902 10756
rect 60844 10168 60856 10744
rect 60890 10168 60902 10744
rect 60844 10156 60902 10168
rect 61862 10744 61920 10756
rect 61862 10168 61874 10744
rect 61908 10168 61920 10744
rect 61862 10156 61920 10168
rect 62880 10744 62938 10756
rect 62880 10168 62892 10744
rect 62926 10168 62938 10744
rect 62880 10156 62938 10168
rect 63898 10744 63956 10756
rect 63898 10168 63910 10744
rect 63944 10168 63956 10744
rect 63898 10156 63956 10168
rect 64916 10744 64974 10756
rect 64916 10168 64928 10744
rect 64962 10168 64974 10744
rect 67518 10534 67530 11110
rect 67564 10534 67576 11110
rect 67518 10522 67576 10534
rect 68536 11110 68594 11122
rect 68536 10534 68548 11110
rect 68582 10534 68594 11110
rect 68536 10522 68594 10534
rect 69554 11110 69612 11122
rect 69554 10534 69566 11110
rect 69600 10534 69612 11110
rect 69554 10522 69612 10534
rect 70572 11110 70630 11122
rect 70572 10534 70584 11110
rect 70618 10534 70630 11110
rect 70572 10522 70630 10534
rect 71590 11110 71648 11122
rect 71590 10534 71602 11110
rect 71636 10534 71648 11110
rect 71590 10522 71648 10534
rect 72608 11110 72666 11122
rect 72608 10534 72620 11110
rect 72654 10534 72666 11110
rect 72608 10522 72666 10534
rect 73626 11110 73684 11122
rect 73626 10534 73638 11110
rect 73672 10534 73684 11110
rect 73626 10522 73684 10534
rect 74644 11110 74702 11122
rect 74644 10534 74656 11110
rect 74690 10534 74702 11110
rect 74644 10522 74702 10534
rect 75662 11110 75720 11122
rect 75662 10534 75674 11110
rect 75708 10534 75720 11110
rect 75662 10522 75720 10534
rect 76680 11110 76738 11122
rect 76680 10534 76692 11110
rect 76726 10534 76738 11110
rect 76680 10522 76738 10534
rect 77698 11110 77756 11122
rect 77698 10534 77710 11110
rect 77744 10534 77756 11110
rect 77698 10522 77756 10534
rect 78716 11110 78774 11122
rect 78716 10534 78728 11110
rect 78762 10534 78774 11110
rect 78716 10522 78774 10534
rect 79734 11110 79792 11122
rect 79734 10534 79746 11110
rect 79780 10534 79792 11110
rect 79734 10522 79792 10534
rect 80752 11110 80810 11122
rect 80752 10534 80764 11110
rect 80798 10534 80810 11110
rect 80752 10522 80810 10534
rect 81770 11110 81828 11122
rect 81770 10534 81782 11110
rect 81816 10534 81828 11110
rect 81770 10522 81828 10534
rect 82788 11110 82846 11122
rect 82788 10534 82800 11110
rect 82834 10534 82846 11110
rect 82788 10522 82846 10534
rect 83806 11110 83864 11122
rect 83806 10534 83818 11110
rect 83852 10534 83864 11110
rect 83806 10522 83864 10534
rect 84824 11110 84882 11122
rect 84824 10534 84836 11110
rect 84870 10534 84882 11110
rect 84824 10522 84882 10534
rect 85842 11110 85900 11122
rect 85842 10534 85854 11110
rect 85888 10534 85900 11110
rect 85842 10522 85900 10534
rect 86860 11110 86918 11122
rect 86860 10534 86872 11110
rect 86906 10534 86918 11110
rect 86860 10522 86918 10534
rect 87878 11110 87936 11122
rect 87878 10534 87890 11110
rect 87924 10534 87936 11110
rect 87878 10522 87936 10534
rect 64916 10156 64974 10168
rect 55754 9926 55812 9938
rect 55754 9350 55766 9926
rect 55800 9350 55812 9926
rect 55754 9338 55812 9350
rect 56772 9926 56830 9938
rect 56772 9350 56784 9926
rect 56818 9350 56830 9926
rect 56772 9338 56830 9350
rect 57790 9926 57848 9938
rect 57790 9350 57802 9926
rect 57836 9350 57848 9926
rect 57790 9338 57848 9350
rect 58808 9926 58866 9938
rect 58808 9350 58820 9926
rect 58854 9350 58866 9926
rect 58808 9338 58866 9350
rect 59826 9926 59884 9938
rect 59826 9350 59838 9926
rect 59872 9350 59884 9926
rect 59826 9338 59884 9350
rect 60844 9926 60902 9938
rect 60844 9350 60856 9926
rect 60890 9350 60902 9926
rect 60844 9338 60902 9350
rect 61862 9926 61920 9938
rect 61862 9350 61874 9926
rect 61908 9350 61920 9926
rect 61862 9338 61920 9350
rect 62880 9926 62938 9938
rect 62880 9350 62892 9926
rect 62926 9350 62938 9926
rect 62880 9338 62938 9350
rect 63898 9926 63956 9938
rect 63898 9350 63910 9926
rect 63944 9350 63956 9926
rect 63898 9338 63956 9350
rect 64916 9926 64974 9938
rect 64916 9350 64928 9926
rect 64962 9350 64974 9926
rect 64916 9338 64974 9350
rect 67518 9876 67576 9888
rect 67518 9300 67530 9876
rect 67564 9300 67576 9876
rect 67518 9288 67576 9300
rect 68536 9876 68594 9888
rect 68536 9300 68548 9876
rect 68582 9300 68594 9876
rect 68536 9288 68594 9300
rect 69554 9876 69612 9888
rect 69554 9300 69566 9876
rect 69600 9300 69612 9876
rect 69554 9288 69612 9300
rect 70572 9876 70630 9888
rect 70572 9300 70584 9876
rect 70618 9300 70630 9876
rect 70572 9288 70630 9300
rect 71590 9876 71648 9888
rect 71590 9300 71602 9876
rect 71636 9300 71648 9876
rect 71590 9288 71648 9300
rect 72608 9876 72666 9888
rect 72608 9300 72620 9876
rect 72654 9300 72666 9876
rect 72608 9288 72666 9300
rect 73626 9876 73684 9888
rect 73626 9300 73638 9876
rect 73672 9300 73684 9876
rect 73626 9288 73684 9300
rect 74644 9876 74702 9888
rect 74644 9300 74656 9876
rect 74690 9300 74702 9876
rect 74644 9288 74702 9300
rect 75662 9876 75720 9888
rect 75662 9300 75674 9876
rect 75708 9300 75720 9876
rect 75662 9288 75720 9300
rect 76680 9876 76738 9888
rect 76680 9300 76692 9876
rect 76726 9300 76738 9876
rect 76680 9288 76738 9300
rect 77698 9876 77756 9888
rect 77698 9300 77710 9876
rect 77744 9300 77756 9876
rect 77698 9288 77756 9300
rect 78716 9876 78774 9888
rect 78716 9300 78728 9876
rect 78762 9300 78774 9876
rect 78716 9288 78774 9300
rect 79734 9876 79792 9888
rect 79734 9300 79746 9876
rect 79780 9300 79792 9876
rect 79734 9288 79792 9300
rect 80752 9876 80810 9888
rect 80752 9300 80764 9876
rect 80798 9300 80810 9876
rect 80752 9288 80810 9300
rect 81770 9876 81828 9888
rect 81770 9300 81782 9876
rect 81816 9300 81828 9876
rect 81770 9288 81828 9300
rect 82788 9876 82846 9888
rect 82788 9300 82800 9876
rect 82834 9300 82846 9876
rect 82788 9288 82846 9300
rect 83806 9876 83864 9888
rect 83806 9300 83818 9876
rect 83852 9300 83864 9876
rect 83806 9288 83864 9300
rect 84824 9876 84882 9888
rect 84824 9300 84836 9876
rect 84870 9300 84882 9876
rect 84824 9288 84882 9300
rect 85842 9876 85900 9888
rect 85842 9300 85854 9876
rect 85888 9300 85900 9876
rect 85842 9288 85900 9300
rect 86860 9876 86918 9888
rect 86860 9300 86872 9876
rect 86906 9300 86918 9876
rect 86860 9288 86918 9300
rect 87878 9876 87936 9888
rect 87878 9300 87890 9876
rect 87924 9300 87936 9876
rect 87878 9288 87936 9300
rect 55754 9108 55812 9120
rect 55754 8532 55766 9108
rect 55800 8532 55812 9108
rect 55754 8520 55812 8532
rect 56772 9108 56830 9120
rect 56772 8532 56784 9108
rect 56818 8532 56830 9108
rect 56772 8520 56830 8532
rect 57790 9108 57848 9120
rect 57790 8532 57802 9108
rect 57836 8532 57848 9108
rect 57790 8520 57848 8532
rect 58808 9108 58866 9120
rect 58808 8532 58820 9108
rect 58854 8532 58866 9108
rect 58808 8520 58866 8532
rect 59826 9108 59884 9120
rect 59826 8532 59838 9108
rect 59872 8532 59884 9108
rect 59826 8520 59884 8532
rect 60844 9108 60902 9120
rect 60844 8532 60856 9108
rect 60890 8532 60902 9108
rect 60844 8520 60902 8532
rect 61862 9108 61920 9120
rect 61862 8532 61874 9108
rect 61908 8532 61920 9108
rect 61862 8520 61920 8532
rect 62880 9108 62938 9120
rect 62880 8532 62892 9108
rect 62926 8532 62938 9108
rect 62880 8520 62938 8532
rect 63898 9108 63956 9120
rect 63898 8532 63910 9108
rect 63944 8532 63956 9108
rect 63898 8520 63956 8532
rect 64916 9108 64974 9120
rect 64916 8532 64928 9108
rect 64962 8532 64974 9108
rect 64916 8520 64974 8532
rect 67518 8644 67576 8656
rect 55754 8290 55812 8302
rect 55754 7714 55766 8290
rect 55800 7714 55812 8290
rect 55754 7702 55812 7714
rect 56772 8290 56830 8302
rect 56772 7714 56784 8290
rect 56818 7714 56830 8290
rect 56772 7702 56830 7714
rect 57790 8290 57848 8302
rect 57790 7714 57802 8290
rect 57836 7714 57848 8290
rect 57790 7702 57848 7714
rect 58808 8290 58866 8302
rect 58808 7714 58820 8290
rect 58854 7714 58866 8290
rect 58808 7702 58866 7714
rect 59826 8290 59884 8302
rect 59826 7714 59838 8290
rect 59872 7714 59884 8290
rect 59826 7702 59884 7714
rect 60844 8290 60902 8302
rect 60844 7714 60856 8290
rect 60890 7714 60902 8290
rect 60844 7702 60902 7714
rect 61862 8290 61920 8302
rect 61862 7714 61874 8290
rect 61908 7714 61920 8290
rect 61862 7702 61920 7714
rect 62880 8290 62938 8302
rect 62880 7714 62892 8290
rect 62926 7714 62938 8290
rect 62880 7702 62938 7714
rect 63898 8290 63956 8302
rect 63898 7714 63910 8290
rect 63944 7714 63956 8290
rect 63898 7702 63956 7714
rect 64916 8290 64974 8302
rect 64916 7714 64928 8290
rect 64962 7714 64974 8290
rect 67518 8068 67530 8644
rect 67564 8068 67576 8644
rect 67518 8056 67576 8068
rect 68536 8644 68594 8656
rect 68536 8068 68548 8644
rect 68582 8068 68594 8644
rect 68536 8056 68594 8068
rect 69554 8644 69612 8656
rect 69554 8068 69566 8644
rect 69600 8068 69612 8644
rect 69554 8056 69612 8068
rect 70572 8644 70630 8656
rect 70572 8068 70584 8644
rect 70618 8068 70630 8644
rect 70572 8056 70630 8068
rect 71590 8644 71648 8656
rect 71590 8068 71602 8644
rect 71636 8068 71648 8644
rect 71590 8056 71648 8068
rect 72608 8644 72666 8656
rect 72608 8068 72620 8644
rect 72654 8068 72666 8644
rect 72608 8056 72666 8068
rect 73626 8644 73684 8656
rect 73626 8068 73638 8644
rect 73672 8068 73684 8644
rect 73626 8056 73684 8068
rect 74644 8644 74702 8656
rect 74644 8068 74656 8644
rect 74690 8068 74702 8644
rect 74644 8056 74702 8068
rect 75662 8644 75720 8656
rect 75662 8068 75674 8644
rect 75708 8068 75720 8644
rect 75662 8056 75720 8068
rect 76680 8644 76738 8656
rect 76680 8068 76692 8644
rect 76726 8068 76738 8644
rect 76680 8056 76738 8068
rect 77698 8644 77756 8656
rect 77698 8068 77710 8644
rect 77744 8068 77756 8644
rect 77698 8056 77756 8068
rect 78716 8644 78774 8656
rect 78716 8068 78728 8644
rect 78762 8068 78774 8644
rect 78716 8056 78774 8068
rect 79734 8644 79792 8656
rect 79734 8068 79746 8644
rect 79780 8068 79792 8644
rect 79734 8056 79792 8068
rect 80752 8644 80810 8656
rect 80752 8068 80764 8644
rect 80798 8068 80810 8644
rect 80752 8056 80810 8068
rect 81770 8644 81828 8656
rect 81770 8068 81782 8644
rect 81816 8068 81828 8644
rect 81770 8056 81828 8068
rect 82788 8644 82846 8656
rect 82788 8068 82800 8644
rect 82834 8068 82846 8644
rect 82788 8056 82846 8068
rect 83806 8644 83864 8656
rect 83806 8068 83818 8644
rect 83852 8068 83864 8644
rect 83806 8056 83864 8068
rect 84824 8644 84882 8656
rect 84824 8068 84836 8644
rect 84870 8068 84882 8644
rect 84824 8056 84882 8068
rect 85842 8644 85900 8656
rect 85842 8068 85854 8644
rect 85888 8068 85900 8644
rect 85842 8056 85900 8068
rect 86860 8644 86918 8656
rect 86860 8068 86872 8644
rect 86906 8068 86918 8644
rect 86860 8056 86918 8068
rect 87878 8644 87936 8656
rect 87878 8068 87890 8644
rect 87924 8068 87936 8644
rect 87878 8056 87936 8068
rect 64916 7702 64974 7714
rect 67518 7410 67576 7422
rect 62614 6906 62672 6918
rect 62614 6730 62626 6906
rect 62660 6730 62672 6906
rect 62614 6718 62672 6730
rect 62832 6906 62890 6918
rect 62832 6730 62844 6906
rect 62878 6730 62890 6906
rect 62832 6718 62890 6730
rect 63050 6906 63108 6918
rect 63050 6730 63062 6906
rect 63096 6730 63108 6906
rect 63050 6718 63108 6730
rect 63268 6906 63326 6918
rect 63268 6730 63280 6906
rect 63314 6730 63326 6906
rect 63268 6718 63326 6730
rect 63486 6906 63544 6918
rect 63486 6730 63498 6906
rect 63532 6730 63544 6906
rect 63486 6718 63544 6730
rect 63704 6906 63762 6918
rect 63704 6730 63716 6906
rect 63750 6730 63762 6906
rect 63704 6718 63762 6730
rect 63922 6906 63980 6918
rect 63922 6730 63934 6906
rect 63968 6730 63980 6906
rect 63922 6718 63980 6730
rect 64140 6906 64198 6918
rect 64140 6730 64152 6906
rect 64186 6730 64198 6906
rect 64140 6718 64198 6730
rect 64358 6906 64416 6918
rect 64358 6730 64370 6906
rect 64404 6730 64416 6906
rect 64358 6718 64416 6730
rect 64576 6906 64634 6918
rect 64576 6730 64588 6906
rect 64622 6730 64634 6906
rect 64576 6718 64634 6730
rect 64794 6906 64852 6918
rect 64794 6730 64806 6906
rect 64840 6730 64852 6906
rect 67518 6834 67530 7410
rect 67564 6834 67576 7410
rect 67518 6822 67576 6834
rect 68536 7410 68594 7422
rect 68536 6834 68548 7410
rect 68582 6834 68594 7410
rect 68536 6822 68594 6834
rect 69554 7410 69612 7422
rect 69554 6834 69566 7410
rect 69600 6834 69612 7410
rect 69554 6822 69612 6834
rect 70572 7410 70630 7422
rect 70572 6834 70584 7410
rect 70618 6834 70630 7410
rect 70572 6822 70630 6834
rect 71590 7410 71648 7422
rect 71590 6834 71602 7410
rect 71636 6834 71648 7410
rect 71590 6822 71648 6834
rect 72608 7410 72666 7422
rect 72608 6834 72620 7410
rect 72654 6834 72666 7410
rect 72608 6822 72666 6834
rect 73626 7410 73684 7422
rect 73626 6834 73638 7410
rect 73672 6834 73684 7410
rect 73626 6822 73684 6834
rect 74644 7410 74702 7422
rect 74644 6834 74656 7410
rect 74690 6834 74702 7410
rect 74644 6822 74702 6834
rect 75662 7410 75720 7422
rect 75662 6834 75674 7410
rect 75708 6834 75720 7410
rect 75662 6822 75720 6834
rect 76680 7410 76738 7422
rect 76680 6834 76692 7410
rect 76726 6834 76738 7410
rect 76680 6822 76738 6834
rect 77698 7410 77756 7422
rect 77698 6834 77710 7410
rect 77744 6834 77756 7410
rect 77698 6822 77756 6834
rect 78716 7410 78774 7422
rect 78716 6834 78728 7410
rect 78762 6834 78774 7410
rect 78716 6822 78774 6834
rect 79734 7410 79792 7422
rect 79734 6834 79746 7410
rect 79780 6834 79792 7410
rect 79734 6822 79792 6834
rect 80752 7410 80810 7422
rect 80752 6834 80764 7410
rect 80798 6834 80810 7410
rect 80752 6822 80810 6834
rect 81770 7410 81828 7422
rect 81770 6834 81782 7410
rect 81816 6834 81828 7410
rect 81770 6822 81828 6834
rect 82788 7410 82846 7422
rect 82788 6834 82800 7410
rect 82834 6834 82846 7410
rect 82788 6822 82846 6834
rect 83806 7410 83864 7422
rect 83806 6834 83818 7410
rect 83852 6834 83864 7410
rect 83806 6822 83864 6834
rect 84824 7410 84882 7422
rect 84824 6834 84836 7410
rect 84870 6834 84882 7410
rect 84824 6822 84882 6834
rect 85842 7410 85900 7422
rect 85842 6834 85854 7410
rect 85888 6834 85900 7410
rect 85842 6822 85900 6834
rect 86860 7410 86918 7422
rect 86860 6834 86872 7410
rect 86906 6834 86918 7410
rect 86860 6822 86918 6834
rect 87878 7410 87936 7422
rect 87878 6834 87890 7410
rect 87924 6834 87936 7410
rect 87878 6822 87936 6834
rect 64794 6718 64852 6730
rect 67518 6176 67576 6188
rect 62614 6074 62672 6086
rect 62614 5898 62626 6074
rect 62660 5898 62672 6074
rect 62614 5886 62672 5898
rect 62832 6074 62890 6086
rect 62832 5898 62844 6074
rect 62878 5898 62890 6074
rect 62832 5886 62890 5898
rect 63050 6074 63108 6086
rect 63050 5898 63062 6074
rect 63096 5898 63108 6074
rect 63050 5886 63108 5898
rect 63268 6074 63326 6086
rect 63268 5898 63280 6074
rect 63314 5898 63326 6074
rect 63268 5886 63326 5898
rect 63486 6074 63544 6086
rect 63486 5898 63498 6074
rect 63532 5898 63544 6074
rect 63486 5886 63544 5898
rect 63704 6074 63762 6086
rect 63704 5898 63716 6074
rect 63750 5898 63762 6074
rect 63704 5886 63762 5898
rect 63922 6074 63980 6086
rect 63922 5898 63934 6074
rect 63968 5898 63980 6074
rect 63922 5886 63980 5898
rect 64140 6074 64198 6086
rect 64140 5898 64152 6074
rect 64186 5898 64198 6074
rect 64140 5886 64198 5898
rect 64358 6074 64416 6086
rect 64358 5898 64370 6074
rect 64404 5898 64416 6074
rect 64358 5886 64416 5898
rect 64576 6074 64634 6086
rect 64576 5898 64588 6074
rect 64622 5898 64634 6074
rect 64576 5886 64634 5898
rect 64794 6074 64852 6086
rect 64794 5898 64806 6074
rect 64840 5898 64852 6074
rect 64794 5886 64852 5898
rect 67518 5600 67530 6176
rect 67564 5600 67576 6176
rect 67518 5588 67576 5600
rect 68536 6176 68594 6188
rect 68536 5600 68548 6176
rect 68582 5600 68594 6176
rect 68536 5588 68594 5600
rect 69554 6176 69612 6188
rect 69554 5600 69566 6176
rect 69600 5600 69612 6176
rect 69554 5588 69612 5600
rect 70572 6176 70630 6188
rect 70572 5600 70584 6176
rect 70618 5600 70630 6176
rect 70572 5588 70630 5600
rect 71590 6176 71648 6188
rect 71590 5600 71602 6176
rect 71636 5600 71648 6176
rect 71590 5588 71648 5600
rect 72608 6176 72666 6188
rect 72608 5600 72620 6176
rect 72654 5600 72666 6176
rect 72608 5588 72666 5600
rect 73626 6176 73684 6188
rect 73626 5600 73638 6176
rect 73672 5600 73684 6176
rect 73626 5588 73684 5600
rect 74644 6176 74702 6188
rect 74644 5600 74656 6176
rect 74690 5600 74702 6176
rect 74644 5588 74702 5600
rect 75662 6176 75720 6188
rect 75662 5600 75674 6176
rect 75708 5600 75720 6176
rect 75662 5588 75720 5600
rect 76680 6176 76738 6188
rect 76680 5600 76692 6176
rect 76726 5600 76738 6176
rect 76680 5588 76738 5600
rect 77698 6176 77756 6188
rect 77698 5600 77710 6176
rect 77744 5600 77756 6176
rect 77698 5588 77756 5600
rect 78716 6176 78774 6188
rect 78716 5600 78728 6176
rect 78762 5600 78774 6176
rect 78716 5588 78774 5600
rect 79734 6176 79792 6188
rect 79734 5600 79746 6176
rect 79780 5600 79792 6176
rect 79734 5588 79792 5600
rect 80752 6176 80810 6188
rect 80752 5600 80764 6176
rect 80798 5600 80810 6176
rect 80752 5588 80810 5600
rect 81770 6176 81828 6188
rect 81770 5600 81782 6176
rect 81816 5600 81828 6176
rect 81770 5588 81828 5600
rect 82788 6176 82846 6188
rect 82788 5600 82800 6176
rect 82834 5600 82846 6176
rect 82788 5588 82846 5600
rect 83806 6176 83864 6188
rect 83806 5600 83818 6176
rect 83852 5600 83864 6176
rect 83806 5588 83864 5600
rect 84824 6176 84882 6188
rect 84824 5600 84836 6176
rect 84870 5600 84882 6176
rect 84824 5588 84882 5600
rect 85842 6176 85900 6188
rect 85842 5600 85854 6176
rect 85888 5600 85900 6176
rect 85842 5588 85900 5600
rect 86860 6176 86918 6188
rect 86860 5600 86872 6176
rect 86906 5600 86918 6176
rect 86860 5588 86918 5600
rect 87878 6176 87936 6188
rect 87878 5600 87890 6176
rect 87924 5600 87936 6176
rect 87878 5588 87936 5600
rect 67518 4944 67576 4956
rect 55533 4747 55591 4759
rect 55533 4171 55545 4747
rect 55579 4171 55591 4747
rect 55533 4159 55591 4171
rect 56551 4747 56609 4759
rect 56551 4171 56563 4747
rect 56597 4171 56609 4747
rect 56551 4159 56609 4171
rect 57569 4747 57627 4759
rect 57569 4171 57581 4747
rect 57615 4171 57627 4747
rect 57569 4159 57627 4171
rect 58587 4747 58645 4759
rect 58587 4171 58599 4747
rect 58633 4171 58645 4747
rect 58587 4159 58645 4171
rect 59605 4747 59663 4759
rect 59605 4171 59617 4747
rect 59651 4171 59663 4747
rect 59605 4159 59663 4171
rect 60623 4747 60681 4759
rect 60623 4171 60635 4747
rect 60669 4171 60681 4747
rect 60623 4159 60681 4171
rect 61641 4747 61699 4759
rect 61641 4171 61653 4747
rect 61687 4171 61699 4747
rect 61641 4159 61699 4171
rect 62528 4748 62586 4760
rect 62528 4172 62540 4748
rect 62574 4172 62586 4748
rect 62528 4160 62586 4172
rect 62826 4748 62884 4760
rect 62826 4172 62838 4748
rect 62872 4172 62884 4748
rect 62826 4160 62884 4172
rect 63124 4748 63182 4760
rect 63124 4172 63136 4748
rect 63170 4172 63182 4748
rect 63124 4160 63182 4172
rect 63422 4748 63480 4760
rect 63422 4172 63434 4748
rect 63468 4172 63480 4748
rect 63422 4160 63480 4172
rect 63720 4748 63778 4760
rect 63720 4172 63732 4748
rect 63766 4172 63778 4748
rect 63720 4160 63778 4172
rect 64018 4748 64076 4760
rect 64018 4172 64030 4748
rect 64064 4172 64076 4748
rect 64018 4160 64076 4172
rect 64316 4748 64374 4760
rect 64316 4172 64328 4748
rect 64362 4172 64374 4748
rect 64316 4160 64374 4172
rect 64614 4748 64672 4760
rect 64614 4172 64626 4748
rect 64660 4172 64672 4748
rect 64614 4160 64672 4172
rect 64912 4748 64970 4760
rect 64912 4172 64924 4748
rect 64958 4172 64970 4748
rect 64912 4160 64970 4172
rect 65210 4748 65268 4760
rect 65210 4172 65222 4748
rect 65256 4172 65268 4748
rect 65210 4160 65268 4172
rect 65508 4748 65566 4760
rect 65508 4172 65520 4748
rect 65554 4172 65566 4748
rect 65508 4160 65566 4172
rect 65806 4748 65864 4760
rect 65806 4172 65818 4748
rect 65852 4172 65864 4748
rect 67518 4368 67530 4944
rect 67564 4368 67576 4944
rect 67518 4356 67576 4368
rect 68536 4944 68594 4956
rect 68536 4368 68548 4944
rect 68582 4368 68594 4944
rect 68536 4356 68594 4368
rect 69554 4944 69612 4956
rect 69554 4368 69566 4944
rect 69600 4368 69612 4944
rect 69554 4356 69612 4368
rect 70572 4944 70630 4956
rect 70572 4368 70584 4944
rect 70618 4368 70630 4944
rect 70572 4356 70630 4368
rect 71590 4944 71648 4956
rect 71590 4368 71602 4944
rect 71636 4368 71648 4944
rect 71590 4356 71648 4368
rect 72608 4944 72666 4956
rect 72608 4368 72620 4944
rect 72654 4368 72666 4944
rect 72608 4356 72666 4368
rect 73626 4944 73684 4956
rect 73626 4368 73638 4944
rect 73672 4368 73684 4944
rect 73626 4356 73684 4368
rect 74644 4944 74702 4956
rect 74644 4368 74656 4944
rect 74690 4368 74702 4944
rect 74644 4356 74702 4368
rect 75662 4944 75720 4956
rect 75662 4368 75674 4944
rect 75708 4368 75720 4944
rect 75662 4356 75720 4368
rect 76680 4944 76738 4956
rect 76680 4368 76692 4944
rect 76726 4368 76738 4944
rect 76680 4356 76738 4368
rect 77698 4944 77756 4956
rect 77698 4368 77710 4944
rect 77744 4368 77756 4944
rect 77698 4356 77756 4368
rect 78716 4944 78774 4956
rect 78716 4368 78728 4944
rect 78762 4368 78774 4944
rect 78716 4356 78774 4368
rect 79734 4944 79792 4956
rect 79734 4368 79746 4944
rect 79780 4368 79792 4944
rect 79734 4356 79792 4368
rect 80752 4944 80810 4956
rect 80752 4368 80764 4944
rect 80798 4368 80810 4944
rect 80752 4356 80810 4368
rect 81770 4944 81828 4956
rect 81770 4368 81782 4944
rect 81816 4368 81828 4944
rect 81770 4356 81828 4368
rect 82788 4944 82846 4956
rect 82788 4368 82800 4944
rect 82834 4368 82846 4944
rect 82788 4356 82846 4368
rect 83806 4944 83864 4956
rect 83806 4368 83818 4944
rect 83852 4368 83864 4944
rect 83806 4356 83864 4368
rect 84824 4944 84882 4956
rect 84824 4368 84836 4944
rect 84870 4368 84882 4944
rect 84824 4356 84882 4368
rect 85842 4944 85900 4956
rect 85842 4368 85854 4944
rect 85888 4368 85900 4944
rect 85842 4356 85900 4368
rect 86860 4944 86918 4956
rect 86860 4368 86872 4944
rect 86906 4368 86918 4944
rect 86860 4356 86918 4368
rect 87878 4944 87936 4956
rect 87878 4368 87890 4944
rect 87924 4368 87936 4944
rect 87878 4356 87936 4368
rect 65806 4160 65864 4172
rect 67518 3710 67576 3722
rect 55532 3634 55590 3646
rect 55532 3058 55544 3634
rect 55578 3058 55590 3634
rect 55532 3046 55590 3058
rect 56550 3634 56608 3646
rect 56550 3058 56562 3634
rect 56596 3058 56608 3634
rect 56550 3046 56608 3058
rect 57568 3634 57626 3646
rect 57568 3058 57580 3634
rect 57614 3058 57626 3634
rect 57568 3046 57626 3058
rect 58586 3634 58644 3646
rect 58586 3058 58598 3634
rect 58632 3058 58644 3634
rect 58586 3046 58644 3058
rect 59604 3634 59662 3646
rect 59604 3058 59616 3634
rect 59650 3058 59662 3634
rect 59604 3046 59662 3058
rect 60622 3634 60680 3646
rect 60622 3058 60634 3634
rect 60668 3058 60680 3634
rect 60622 3046 60680 3058
rect 61640 3634 61698 3646
rect 61640 3058 61652 3634
rect 61686 3058 61698 3634
rect 61640 3046 61698 3058
rect 62528 3636 62586 3648
rect 62528 3060 62540 3636
rect 62574 3060 62586 3636
rect 62528 3048 62586 3060
rect 62826 3636 62884 3648
rect 62826 3060 62838 3636
rect 62872 3060 62884 3636
rect 62826 3048 62884 3060
rect 63124 3636 63182 3648
rect 63124 3060 63136 3636
rect 63170 3060 63182 3636
rect 63124 3048 63182 3060
rect 63422 3636 63480 3648
rect 63422 3060 63434 3636
rect 63468 3060 63480 3636
rect 63422 3048 63480 3060
rect 63720 3636 63778 3648
rect 63720 3060 63732 3636
rect 63766 3060 63778 3636
rect 63720 3048 63778 3060
rect 64018 3636 64076 3648
rect 64018 3060 64030 3636
rect 64064 3060 64076 3636
rect 64018 3048 64076 3060
rect 64316 3636 64374 3648
rect 64316 3060 64328 3636
rect 64362 3060 64374 3636
rect 64316 3048 64374 3060
rect 64614 3636 64672 3648
rect 64614 3060 64626 3636
rect 64660 3060 64672 3636
rect 64614 3048 64672 3060
rect 64912 3636 64970 3648
rect 64912 3060 64924 3636
rect 64958 3060 64970 3636
rect 64912 3048 64970 3060
rect 65210 3636 65268 3648
rect 65210 3060 65222 3636
rect 65256 3060 65268 3636
rect 65210 3048 65268 3060
rect 65508 3636 65566 3648
rect 65508 3060 65520 3636
rect 65554 3060 65566 3636
rect 65508 3048 65566 3060
rect 65806 3636 65864 3648
rect 65806 3060 65818 3636
rect 65852 3060 65864 3636
rect 67518 3134 67530 3710
rect 67564 3134 67576 3710
rect 67518 3122 67576 3134
rect 68536 3710 68594 3722
rect 68536 3134 68548 3710
rect 68582 3134 68594 3710
rect 68536 3122 68594 3134
rect 69554 3710 69612 3722
rect 69554 3134 69566 3710
rect 69600 3134 69612 3710
rect 69554 3122 69612 3134
rect 70572 3710 70630 3722
rect 70572 3134 70584 3710
rect 70618 3134 70630 3710
rect 70572 3122 70630 3134
rect 71590 3710 71648 3722
rect 71590 3134 71602 3710
rect 71636 3134 71648 3710
rect 71590 3122 71648 3134
rect 72608 3710 72666 3722
rect 72608 3134 72620 3710
rect 72654 3134 72666 3710
rect 72608 3122 72666 3134
rect 73626 3710 73684 3722
rect 73626 3134 73638 3710
rect 73672 3134 73684 3710
rect 73626 3122 73684 3134
rect 74644 3710 74702 3722
rect 74644 3134 74656 3710
rect 74690 3134 74702 3710
rect 74644 3122 74702 3134
rect 75662 3710 75720 3722
rect 75662 3134 75674 3710
rect 75708 3134 75720 3710
rect 75662 3122 75720 3134
rect 76680 3710 76738 3722
rect 76680 3134 76692 3710
rect 76726 3134 76738 3710
rect 76680 3122 76738 3134
rect 77698 3710 77756 3722
rect 77698 3134 77710 3710
rect 77744 3134 77756 3710
rect 77698 3122 77756 3134
rect 78716 3710 78774 3722
rect 78716 3134 78728 3710
rect 78762 3134 78774 3710
rect 78716 3122 78774 3134
rect 79734 3710 79792 3722
rect 79734 3134 79746 3710
rect 79780 3134 79792 3710
rect 79734 3122 79792 3134
rect 80752 3710 80810 3722
rect 80752 3134 80764 3710
rect 80798 3134 80810 3710
rect 80752 3122 80810 3134
rect 81770 3710 81828 3722
rect 81770 3134 81782 3710
rect 81816 3134 81828 3710
rect 81770 3122 81828 3134
rect 82788 3710 82846 3722
rect 82788 3134 82800 3710
rect 82834 3134 82846 3710
rect 82788 3122 82846 3134
rect 83806 3710 83864 3722
rect 83806 3134 83818 3710
rect 83852 3134 83864 3710
rect 83806 3122 83864 3134
rect 84824 3710 84882 3722
rect 84824 3134 84836 3710
rect 84870 3134 84882 3710
rect 84824 3122 84882 3134
rect 85842 3710 85900 3722
rect 85842 3134 85854 3710
rect 85888 3134 85900 3710
rect 85842 3122 85900 3134
rect 86860 3710 86918 3722
rect 86860 3134 86872 3710
rect 86906 3134 86918 3710
rect 86860 3122 86918 3134
rect 87878 3710 87936 3722
rect 87878 3134 87890 3710
rect 87924 3134 87936 3710
rect 87878 3122 87936 3134
rect 65806 3048 65864 3060
rect 55533 2523 55591 2535
rect 55533 1947 55545 2523
rect 55579 1947 55591 2523
rect 55533 1935 55591 1947
rect 56551 2523 56609 2535
rect 56551 1947 56563 2523
rect 56597 1947 56609 2523
rect 56551 1935 56609 1947
rect 57569 2523 57627 2535
rect 57569 1947 57581 2523
rect 57615 1947 57627 2523
rect 57569 1935 57627 1947
rect 58587 2523 58645 2535
rect 58587 1947 58599 2523
rect 58633 1947 58645 2523
rect 58587 1935 58645 1947
rect 59605 2523 59663 2535
rect 59605 1947 59617 2523
rect 59651 1947 59663 2523
rect 59605 1935 59663 1947
rect 60623 2523 60681 2535
rect 60623 1947 60635 2523
rect 60669 1947 60681 2523
rect 60623 1935 60681 1947
rect 61641 2523 61699 2535
rect 61641 1947 61653 2523
rect 61687 1947 61699 2523
rect 61641 1935 61699 1947
rect 62526 2524 62584 2536
rect 62526 1948 62538 2524
rect 62572 1948 62584 2524
rect 62526 1936 62584 1948
rect 62824 2524 62882 2536
rect 62824 1948 62836 2524
rect 62870 1948 62882 2524
rect 62824 1936 62882 1948
rect 63122 2524 63180 2536
rect 63122 1948 63134 2524
rect 63168 1948 63180 2524
rect 63122 1936 63180 1948
rect 63420 2524 63478 2536
rect 63420 1948 63432 2524
rect 63466 1948 63478 2524
rect 63420 1936 63478 1948
rect 63718 2524 63776 2536
rect 63718 1948 63730 2524
rect 63764 1948 63776 2524
rect 63718 1936 63776 1948
rect 64016 2524 64074 2536
rect 64016 1948 64028 2524
rect 64062 1948 64074 2524
rect 64016 1936 64074 1948
rect 64314 2524 64372 2536
rect 64314 1948 64326 2524
rect 64360 1948 64372 2524
rect 64314 1936 64372 1948
rect 64612 2524 64670 2536
rect 64612 1948 64624 2524
rect 64658 1948 64670 2524
rect 64612 1936 64670 1948
rect 64910 2524 64968 2536
rect 64910 1948 64922 2524
rect 64956 1948 64968 2524
rect 64910 1936 64968 1948
rect 65208 2524 65266 2536
rect 65208 1948 65220 2524
rect 65254 1948 65266 2524
rect 65208 1936 65266 1948
rect 65506 2524 65564 2536
rect 65506 1948 65518 2524
rect 65552 1948 65564 2524
rect 65506 1936 65564 1948
rect 65804 2524 65862 2536
rect 65804 1948 65816 2524
rect 65850 1948 65862 2524
rect 65804 1936 65862 1948
rect 67518 2476 67576 2488
rect 67518 1900 67530 2476
rect 67564 1900 67576 2476
rect 67518 1888 67576 1900
rect 68536 2476 68594 2488
rect 68536 1900 68548 2476
rect 68582 1900 68594 2476
rect 68536 1888 68594 1900
rect 69554 2476 69612 2488
rect 69554 1900 69566 2476
rect 69600 1900 69612 2476
rect 69554 1888 69612 1900
rect 70572 2476 70630 2488
rect 70572 1900 70584 2476
rect 70618 1900 70630 2476
rect 70572 1888 70630 1900
rect 71590 2476 71648 2488
rect 71590 1900 71602 2476
rect 71636 1900 71648 2476
rect 71590 1888 71648 1900
rect 72608 2476 72666 2488
rect 72608 1900 72620 2476
rect 72654 1900 72666 2476
rect 72608 1888 72666 1900
rect 73626 2476 73684 2488
rect 73626 1900 73638 2476
rect 73672 1900 73684 2476
rect 73626 1888 73684 1900
rect 74644 2476 74702 2488
rect 74644 1900 74656 2476
rect 74690 1900 74702 2476
rect 74644 1888 74702 1900
rect 75662 2476 75720 2488
rect 75662 1900 75674 2476
rect 75708 1900 75720 2476
rect 75662 1888 75720 1900
rect 76680 2476 76738 2488
rect 76680 1900 76692 2476
rect 76726 1900 76738 2476
rect 76680 1888 76738 1900
rect 77698 2476 77756 2488
rect 77698 1900 77710 2476
rect 77744 1900 77756 2476
rect 77698 1888 77756 1900
rect 78716 2476 78774 2488
rect 78716 1900 78728 2476
rect 78762 1900 78774 2476
rect 78716 1888 78774 1900
rect 79734 2476 79792 2488
rect 79734 1900 79746 2476
rect 79780 1900 79792 2476
rect 79734 1888 79792 1900
rect 80752 2476 80810 2488
rect 80752 1900 80764 2476
rect 80798 1900 80810 2476
rect 80752 1888 80810 1900
rect 81770 2476 81828 2488
rect 81770 1900 81782 2476
rect 81816 1900 81828 2476
rect 81770 1888 81828 1900
rect 82788 2476 82846 2488
rect 82788 1900 82800 2476
rect 82834 1900 82846 2476
rect 82788 1888 82846 1900
rect 83806 2476 83864 2488
rect 83806 1900 83818 2476
rect 83852 1900 83864 2476
rect 83806 1888 83864 1900
rect 84824 2476 84882 2488
rect 84824 1900 84836 2476
rect 84870 1900 84882 2476
rect 84824 1888 84882 1900
rect 85842 2476 85900 2488
rect 85842 1900 85854 2476
rect 85888 1900 85900 2476
rect 85842 1888 85900 1900
rect 86860 2476 86918 2488
rect 86860 1900 86872 2476
rect 86906 1900 86918 2476
rect 86860 1888 86918 1900
rect 87878 2476 87936 2488
rect 87878 1900 87890 2476
rect 87924 1900 87936 2476
rect 87878 1888 87936 1900
rect 55532 1410 55590 1422
rect 55532 834 55544 1410
rect 55578 834 55590 1410
rect 55532 822 55590 834
rect 56550 1410 56608 1422
rect 56550 834 56562 1410
rect 56596 834 56608 1410
rect 56550 822 56608 834
rect 57568 1410 57626 1422
rect 57568 834 57580 1410
rect 57614 834 57626 1410
rect 57568 822 57626 834
rect 58586 1410 58644 1422
rect 58586 834 58598 1410
rect 58632 834 58644 1410
rect 58586 822 58644 834
rect 59604 1410 59662 1422
rect 59604 834 59616 1410
rect 59650 834 59662 1410
rect 59604 822 59662 834
rect 60622 1410 60680 1422
rect 60622 834 60634 1410
rect 60668 834 60680 1410
rect 60622 822 60680 834
rect 61640 1410 61698 1422
rect 61640 834 61652 1410
rect 61686 834 61698 1410
rect 61640 822 61698 834
rect 62526 1414 62584 1426
rect 62526 838 62538 1414
rect 62572 838 62584 1414
rect 62526 826 62584 838
rect 62824 1414 62882 1426
rect 62824 838 62836 1414
rect 62870 838 62882 1414
rect 62824 826 62882 838
rect 63122 1414 63180 1426
rect 63122 838 63134 1414
rect 63168 838 63180 1414
rect 63122 826 63180 838
rect 63420 1414 63478 1426
rect 63420 838 63432 1414
rect 63466 838 63478 1414
rect 63420 826 63478 838
rect 63718 1414 63776 1426
rect 63718 838 63730 1414
rect 63764 838 63776 1414
rect 63718 826 63776 838
rect 64016 1414 64074 1426
rect 64016 838 64028 1414
rect 64062 838 64074 1414
rect 64016 826 64074 838
rect 64314 1414 64372 1426
rect 64314 838 64326 1414
rect 64360 838 64372 1414
rect 64314 826 64372 838
rect 64612 1414 64670 1426
rect 64612 838 64624 1414
rect 64658 838 64670 1414
rect 64612 826 64670 838
rect 64910 1414 64968 1426
rect 64910 838 64922 1414
rect 64956 838 64968 1414
rect 64910 826 64968 838
rect 65208 1414 65266 1426
rect 65208 838 65220 1414
rect 65254 838 65266 1414
rect 65208 826 65266 838
rect 65506 1414 65564 1426
rect 65506 838 65518 1414
rect 65552 838 65564 1414
rect 65506 826 65564 838
rect 65804 1414 65862 1426
rect 65804 838 65816 1414
rect 65850 838 65862 1414
rect 65804 826 65862 838
rect 67518 1244 67576 1256
rect 67518 668 67530 1244
rect 67564 668 67576 1244
rect 67518 656 67576 668
rect 68536 1244 68594 1256
rect 68536 668 68548 1244
rect 68582 668 68594 1244
rect 68536 656 68594 668
rect 69554 1244 69612 1256
rect 69554 668 69566 1244
rect 69600 668 69612 1244
rect 69554 656 69612 668
rect 70572 1244 70630 1256
rect 70572 668 70584 1244
rect 70618 668 70630 1244
rect 70572 656 70630 668
rect 71590 1244 71648 1256
rect 71590 668 71602 1244
rect 71636 668 71648 1244
rect 71590 656 71648 668
rect 72608 1244 72666 1256
rect 72608 668 72620 1244
rect 72654 668 72666 1244
rect 72608 656 72666 668
rect 73626 1244 73684 1256
rect 73626 668 73638 1244
rect 73672 668 73684 1244
rect 73626 656 73684 668
rect 74644 1244 74702 1256
rect 74644 668 74656 1244
rect 74690 668 74702 1244
rect 74644 656 74702 668
rect 75662 1244 75720 1256
rect 75662 668 75674 1244
rect 75708 668 75720 1244
rect 75662 656 75720 668
rect 76680 1244 76738 1256
rect 76680 668 76692 1244
rect 76726 668 76738 1244
rect 76680 656 76738 668
rect 77698 1244 77756 1256
rect 77698 668 77710 1244
rect 77744 668 77756 1244
rect 77698 656 77756 668
rect 78716 1244 78774 1256
rect 78716 668 78728 1244
rect 78762 668 78774 1244
rect 78716 656 78774 668
rect 79734 1244 79792 1256
rect 79734 668 79746 1244
rect 79780 668 79792 1244
rect 79734 656 79792 668
rect 80752 1244 80810 1256
rect 80752 668 80764 1244
rect 80798 668 80810 1244
rect 80752 656 80810 668
rect 81770 1244 81828 1256
rect 81770 668 81782 1244
rect 81816 668 81828 1244
rect 81770 656 81828 668
rect 82788 1244 82846 1256
rect 82788 668 82800 1244
rect 82834 668 82846 1244
rect 82788 656 82846 668
rect 83806 1244 83864 1256
rect 83806 668 83818 1244
rect 83852 668 83864 1244
rect 83806 656 83864 668
rect 84824 1244 84882 1256
rect 84824 668 84836 1244
rect 84870 668 84882 1244
rect 84824 656 84882 668
rect 85842 1244 85900 1256
rect 85842 668 85854 1244
rect 85888 668 85900 1244
rect 85842 656 85900 668
rect 86860 1244 86918 1256
rect 86860 668 86872 1244
rect 86906 668 86918 1244
rect 86860 656 86918 668
rect 87878 1244 87936 1256
rect 87878 668 87890 1244
rect 87924 668 87936 1244
rect 87878 656 87936 668
<< pdiff >>
rect 17426 26968 17484 26980
rect 17426 26392 17438 26968
rect 17472 26392 17484 26968
rect 17426 26380 17484 26392
rect 18444 26968 18502 26980
rect 18444 26392 18456 26968
rect 18490 26392 18502 26968
rect 18444 26380 18502 26392
rect 19462 26968 19520 26980
rect 19462 26392 19474 26968
rect 19508 26392 19520 26968
rect 19462 26380 19520 26392
rect 20480 26968 20538 26980
rect 20480 26392 20492 26968
rect 20526 26392 20538 26968
rect 20480 26380 20538 26392
rect 21498 26968 21556 26980
rect 21498 26392 21510 26968
rect 21544 26392 21556 26968
rect 21498 26380 21556 26392
rect 22516 26968 22574 26980
rect 22516 26392 22528 26968
rect 22562 26392 22574 26968
rect 22516 26380 22574 26392
rect 23534 26968 23592 26980
rect 23534 26392 23546 26968
rect 23580 26392 23592 26968
rect 23534 26380 23592 26392
rect 24552 26968 24610 26980
rect 24552 26392 24564 26968
rect 24598 26392 24610 26968
rect 24552 26380 24610 26392
rect 25570 26968 25628 26980
rect 25570 26392 25582 26968
rect 25616 26392 25628 26968
rect 25570 26380 25628 26392
rect 26588 26968 26646 26980
rect 26588 26392 26600 26968
rect 26634 26392 26646 26968
rect 26588 26380 26646 26392
rect 27606 26968 27664 26980
rect 27606 26392 27618 26968
rect 27652 26392 27664 26968
rect 27606 26380 27664 26392
rect 28624 26968 28682 26980
rect 28624 26392 28636 26968
rect 28670 26392 28682 26968
rect 28624 26380 28682 26392
rect 29642 26968 29700 26980
rect 29642 26392 29654 26968
rect 29688 26392 29700 26968
rect 29642 26380 29700 26392
rect 30660 26968 30718 26980
rect 30660 26392 30672 26968
rect 30706 26392 30718 26968
rect 30660 26380 30718 26392
rect 31678 26968 31736 26980
rect 31678 26392 31690 26968
rect 31724 26392 31736 26968
rect 31678 26380 31736 26392
rect 32696 26968 32754 26980
rect 32696 26392 32708 26968
rect 32742 26392 32754 26968
rect 32696 26380 32754 26392
rect 33714 26968 33772 26980
rect 33714 26392 33726 26968
rect 33760 26392 33772 26968
rect 33714 26380 33772 26392
rect 17426 25832 17484 25844
rect 17426 25256 17438 25832
rect 17472 25256 17484 25832
rect 17426 25244 17484 25256
rect 18444 25832 18502 25844
rect 18444 25256 18456 25832
rect 18490 25256 18502 25832
rect 18444 25244 18502 25256
rect 19462 25832 19520 25844
rect 19462 25256 19474 25832
rect 19508 25256 19520 25832
rect 19462 25244 19520 25256
rect 20480 25832 20538 25844
rect 20480 25256 20492 25832
rect 20526 25256 20538 25832
rect 20480 25244 20538 25256
rect 21498 25832 21556 25844
rect 21498 25256 21510 25832
rect 21544 25256 21556 25832
rect 21498 25244 21556 25256
rect 22516 25832 22574 25844
rect 22516 25256 22528 25832
rect 22562 25256 22574 25832
rect 22516 25244 22574 25256
rect 23534 25832 23592 25844
rect 23534 25256 23546 25832
rect 23580 25256 23592 25832
rect 23534 25244 23592 25256
rect 24552 25832 24610 25844
rect 24552 25256 24564 25832
rect 24598 25256 24610 25832
rect 24552 25244 24610 25256
rect 25570 25832 25628 25844
rect 25570 25256 25582 25832
rect 25616 25256 25628 25832
rect 25570 25244 25628 25256
rect 26588 25832 26646 25844
rect 26588 25256 26600 25832
rect 26634 25256 26646 25832
rect 26588 25244 26646 25256
rect 27606 25832 27664 25844
rect 27606 25256 27618 25832
rect 27652 25256 27664 25832
rect 27606 25244 27664 25256
rect 28624 25832 28682 25844
rect 28624 25256 28636 25832
rect 28670 25256 28682 25832
rect 28624 25244 28682 25256
rect 29642 25832 29700 25844
rect 29642 25256 29654 25832
rect 29688 25256 29700 25832
rect 29642 25244 29700 25256
rect 30660 25832 30718 25844
rect 30660 25256 30672 25832
rect 30706 25256 30718 25832
rect 30660 25244 30718 25256
rect 31678 25832 31736 25844
rect 31678 25256 31690 25832
rect 31724 25256 31736 25832
rect 31678 25244 31736 25256
rect 32696 25832 32754 25844
rect 32696 25256 32708 25832
rect 32742 25256 32754 25832
rect 32696 25244 32754 25256
rect 33714 25832 33772 25844
rect 33714 25256 33726 25832
rect 33760 25256 33772 25832
rect 33714 25244 33772 25256
rect 17426 24696 17484 24708
rect 17426 24120 17438 24696
rect 17472 24120 17484 24696
rect 17426 24108 17484 24120
rect 18444 24696 18502 24708
rect 18444 24120 18456 24696
rect 18490 24120 18502 24696
rect 18444 24108 18502 24120
rect 19462 24696 19520 24708
rect 19462 24120 19474 24696
rect 19508 24120 19520 24696
rect 19462 24108 19520 24120
rect 20480 24696 20538 24708
rect 20480 24120 20492 24696
rect 20526 24120 20538 24696
rect 20480 24108 20538 24120
rect 21498 24696 21556 24708
rect 21498 24120 21510 24696
rect 21544 24120 21556 24696
rect 21498 24108 21556 24120
rect 22516 24696 22574 24708
rect 22516 24120 22528 24696
rect 22562 24120 22574 24696
rect 22516 24108 22574 24120
rect 23534 24696 23592 24708
rect 23534 24120 23546 24696
rect 23580 24120 23592 24696
rect 23534 24108 23592 24120
rect 24552 24696 24610 24708
rect 24552 24120 24564 24696
rect 24598 24120 24610 24696
rect 24552 24108 24610 24120
rect 25570 24696 25628 24708
rect 25570 24120 25582 24696
rect 25616 24120 25628 24696
rect 25570 24108 25628 24120
rect 26588 24696 26646 24708
rect 26588 24120 26600 24696
rect 26634 24120 26646 24696
rect 26588 24108 26646 24120
rect 27606 24696 27664 24708
rect 27606 24120 27618 24696
rect 27652 24120 27664 24696
rect 27606 24108 27664 24120
rect 28624 24696 28682 24708
rect 28624 24120 28636 24696
rect 28670 24120 28682 24696
rect 28624 24108 28682 24120
rect 29642 24696 29700 24708
rect 29642 24120 29654 24696
rect 29688 24120 29700 24696
rect 29642 24108 29700 24120
rect 30660 24696 30718 24708
rect 30660 24120 30672 24696
rect 30706 24120 30718 24696
rect 30660 24108 30718 24120
rect 31678 24696 31736 24708
rect 31678 24120 31690 24696
rect 31724 24120 31736 24696
rect 31678 24108 31736 24120
rect 32696 24696 32754 24708
rect 32696 24120 32708 24696
rect 32742 24120 32754 24696
rect 32696 24108 32754 24120
rect 33714 24696 33772 24708
rect 33714 24120 33726 24696
rect 33760 24120 33772 24696
rect 33714 24108 33772 24120
rect 18412 22922 18470 22934
rect 18412 22346 18424 22922
rect 18458 22346 18470 22922
rect 18412 22334 18470 22346
rect 19430 22922 19488 22934
rect 19430 22346 19442 22922
rect 19476 22346 19488 22922
rect 19430 22334 19488 22346
rect 20448 22922 20506 22934
rect 20448 22346 20460 22922
rect 20494 22346 20506 22922
rect 20448 22334 20506 22346
rect 21466 22922 21524 22934
rect 21466 22346 21478 22922
rect 21512 22346 21524 22922
rect 21466 22334 21524 22346
rect 22484 22922 22542 22934
rect 22484 22346 22496 22922
rect 22530 22346 22542 22922
rect 22484 22334 22542 22346
rect 23502 22922 23560 22934
rect 23502 22346 23514 22922
rect 23548 22346 23560 22922
rect 23502 22334 23560 22346
rect 24520 22922 24578 22934
rect 24520 22346 24532 22922
rect 24566 22346 24578 22922
rect 24520 22334 24578 22346
rect 25538 22922 25596 22934
rect 25538 22346 25550 22922
rect 25584 22346 25596 22922
rect 25538 22334 25596 22346
rect 26556 22922 26614 22934
rect 26556 22346 26568 22922
rect 26602 22346 26614 22922
rect 26556 22334 26614 22346
rect 27574 22922 27632 22934
rect 27574 22346 27586 22922
rect 27620 22346 27632 22922
rect 27574 22334 27632 22346
rect 28592 22922 28650 22934
rect 28592 22346 28604 22922
rect 28638 22346 28650 22922
rect 28592 22334 28650 22346
rect 29610 22922 29668 22934
rect 29610 22346 29622 22922
rect 29656 22346 29668 22922
rect 29610 22334 29668 22346
rect 30628 22922 30686 22934
rect 30628 22346 30640 22922
rect 30674 22346 30686 22922
rect 30628 22334 30686 22346
rect 31646 22922 31704 22934
rect 31646 22346 31658 22922
rect 31692 22346 31704 22922
rect 31646 22334 31704 22346
rect 32664 22922 32722 22934
rect 32664 22346 32676 22922
rect 32710 22346 32722 22922
rect 32664 22334 32722 22346
rect 33682 22922 33740 22934
rect 33682 22346 33694 22922
rect 33728 22346 33740 22922
rect 33682 22334 33740 22346
rect 14564 21838 14622 21850
rect 14564 21462 14576 21838
rect 14610 21462 14622 21838
rect 14564 21450 14622 21462
rect 14782 21838 14840 21850
rect 14782 21462 14794 21838
rect 14828 21462 14840 21838
rect 14782 21450 14840 21462
rect 15000 21838 15058 21850
rect 15000 21462 15012 21838
rect 15046 21462 15058 21838
rect 15000 21450 15058 21462
rect 15218 21838 15276 21850
rect 15218 21462 15230 21838
rect 15264 21462 15276 21838
rect 15218 21450 15276 21462
rect 15436 21838 15494 21850
rect 15436 21462 15448 21838
rect 15482 21462 15494 21838
rect 15436 21450 15494 21462
rect 15654 21838 15712 21850
rect 15654 21462 15666 21838
rect 15700 21462 15712 21838
rect 15654 21450 15712 21462
rect 15872 21838 15930 21850
rect 15872 21462 15884 21838
rect 15918 21462 15930 21838
rect 15872 21450 15930 21462
rect 16090 21838 16148 21850
rect 16090 21462 16102 21838
rect 16136 21462 16148 21838
rect 16090 21450 16148 21462
rect 16308 21838 16366 21850
rect 16308 21462 16320 21838
rect 16354 21462 16366 21838
rect 16308 21450 16366 21462
rect 16526 21838 16584 21850
rect 16526 21462 16538 21838
rect 16572 21462 16584 21838
rect 16526 21450 16584 21462
rect 16744 21838 16802 21850
rect 16744 21462 16756 21838
rect 16790 21462 16802 21838
rect 16744 21450 16802 21462
rect 18412 21666 18470 21678
rect 18412 21090 18424 21666
rect 18458 21090 18470 21666
rect 18412 21078 18470 21090
rect 19430 21666 19488 21678
rect 19430 21090 19442 21666
rect 19476 21090 19488 21666
rect 19430 21078 19488 21090
rect 20448 21666 20506 21678
rect 20448 21090 20460 21666
rect 20494 21090 20506 21666
rect 20448 21078 20506 21090
rect 21466 21666 21524 21678
rect 21466 21090 21478 21666
rect 21512 21090 21524 21666
rect 21466 21078 21524 21090
rect 22484 21666 22542 21678
rect 22484 21090 22496 21666
rect 22530 21090 22542 21666
rect 22484 21078 22542 21090
rect 23502 21666 23560 21678
rect 23502 21090 23514 21666
rect 23548 21090 23560 21666
rect 23502 21078 23560 21090
rect 24520 21666 24578 21678
rect 24520 21090 24532 21666
rect 24566 21090 24578 21666
rect 24520 21078 24578 21090
rect 25538 21666 25596 21678
rect 25538 21090 25550 21666
rect 25584 21090 25596 21666
rect 25538 21078 25596 21090
rect 26556 21666 26614 21678
rect 26556 21090 26568 21666
rect 26602 21090 26614 21666
rect 26556 21078 26614 21090
rect 27574 21666 27632 21678
rect 27574 21090 27586 21666
rect 27620 21090 27632 21666
rect 27574 21078 27632 21090
rect 28592 21666 28650 21678
rect 28592 21090 28604 21666
rect 28638 21090 28650 21666
rect 28592 21078 28650 21090
rect 29610 21666 29668 21678
rect 29610 21090 29622 21666
rect 29656 21090 29668 21666
rect 29610 21078 29668 21090
rect 30628 21666 30686 21678
rect 30628 21090 30640 21666
rect 30674 21090 30686 21666
rect 30628 21078 30686 21090
rect 31646 21666 31704 21678
rect 31646 21090 31658 21666
rect 31692 21090 31704 21666
rect 31646 21078 31704 21090
rect 32664 21666 32722 21678
rect 32664 21090 32676 21666
rect 32710 21090 32722 21666
rect 32664 21078 32722 21090
rect 33682 21666 33740 21678
rect 33682 21090 33694 21666
rect 33728 21090 33740 21666
rect 33682 21078 33740 21090
rect 14564 20900 14622 20912
rect 14564 20524 14576 20900
rect 14610 20524 14622 20900
rect 14564 20512 14622 20524
rect 14782 20900 14840 20912
rect 14782 20524 14794 20900
rect 14828 20524 14840 20900
rect 14782 20512 14840 20524
rect 15000 20900 15058 20912
rect 15000 20524 15012 20900
rect 15046 20524 15058 20900
rect 15000 20512 15058 20524
rect 15218 20900 15276 20912
rect 15218 20524 15230 20900
rect 15264 20524 15276 20900
rect 15218 20512 15276 20524
rect 15436 20900 15494 20912
rect 15436 20524 15448 20900
rect 15482 20524 15494 20900
rect 15436 20512 15494 20524
rect 15654 20900 15712 20912
rect 15654 20524 15666 20900
rect 15700 20524 15712 20900
rect 15654 20512 15712 20524
rect 15872 20900 15930 20912
rect 15872 20524 15884 20900
rect 15918 20524 15930 20900
rect 15872 20512 15930 20524
rect 16090 20900 16148 20912
rect 16090 20524 16102 20900
rect 16136 20524 16148 20900
rect 16090 20512 16148 20524
rect 16308 20900 16366 20912
rect 16308 20524 16320 20900
rect 16354 20524 16366 20900
rect 16308 20512 16366 20524
rect 16526 20900 16584 20912
rect 16526 20524 16538 20900
rect 16572 20524 16584 20900
rect 16526 20512 16584 20524
rect 16744 20900 16802 20912
rect 16744 20524 16756 20900
rect 16790 20524 16802 20900
rect 16744 20512 16802 20524
rect 18412 20410 18470 20422
rect 14564 19962 14622 19974
rect 14564 19586 14576 19962
rect 14610 19586 14622 19962
rect 14564 19574 14622 19586
rect 14782 19962 14840 19974
rect 14782 19586 14794 19962
rect 14828 19586 14840 19962
rect 14782 19574 14840 19586
rect 15000 19962 15058 19974
rect 15000 19586 15012 19962
rect 15046 19586 15058 19962
rect 15000 19574 15058 19586
rect 15218 19962 15276 19974
rect 15218 19586 15230 19962
rect 15264 19586 15276 19962
rect 15218 19574 15276 19586
rect 15436 19962 15494 19974
rect 15436 19586 15448 19962
rect 15482 19586 15494 19962
rect 15436 19574 15494 19586
rect 15654 19962 15712 19974
rect 15654 19586 15666 19962
rect 15700 19586 15712 19962
rect 15654 19574 15712 19586
rect 15872 19962 15930 19974
rect 15872 19586 15884 19962
rect 15918 19586 15930 19962
rect 15872 19574 15930 19586
rect 16090 19962 16148 19974
rect 16090 19586 16102 19962
rect 16136 19586 16148 19962
rect 16090 19574 16148 19586
rect 16308 19962 16366 19974
rect 16308 19586 16320 19962
rect 16354 19586 16366 19962
rect 16308 19574 16366 19586
rect 16526 19962 16584 19974
rect 16526 19586 16538 19962
rect 16572 19586 16584 19962
rect 16526 19574 16584 19586
rect 16744 19962 16802 19974
rect 16744 19586 16756 19962
rect 16790 19586 16802 19962
rect 18412 19834 18424 20410
rect 18458 19834 18470 20410
rect 18412 19822 18470 19834
rect 19430 20410 19488 20422
rect 19430 19834 19442 20410
rect 19476 19834 19488 20410
rect 19430 19822 19488 19834
rect 20448 20410 20506 20422
rect 20448 19834 20460 20410
rect 20494 19834 20506 20410
rect 20448 19822 20506 19834
rect 21466 20410 21524 20422
rect 21466 19834 21478 20410
rect 21512 19834 21524 20410
rect 21466 19822 21524 19834
rect 22484 20410 22542 20422
rect 22484 19834 22496 20410
rect 22530 19834 22542 20410
rect 22484 19822 22542 19834
rect 23502 20410 23560 20422
rect 23502 19834 23514 20410
rect 23548 19834 23560 20410
rect 23502 19822 23560 19834
rect 24520 20410 24578 20422
rect 24520 19834 24532 20410
rect 24566 19834 24578 20410
rect 24520 19822 24578 19834
rect 25538 20410 25596 20422
rect 25538 19834 25550 20410
rect 25584 19834 25596 20410
rect 25538 19822 25596 19834
rect 26556 20410 26614 20422
rect 26556 19834 26568 20410
rect 26602 19834 26614 20410
rect 26556 19822 26614 19834
rect 27574 20410 27632 20422
rect 27574 19834 27586 20410
rect 27620 19834 27632 20410
rect 27574 19822 27632 19834
rect 28592 20410 28650 20422
rect 28592 19834 28604 20410
rect 28638 19834 28650 20410
rect 28592 19822 28650 19834
rect 29610 20410 29668 20422
rect 29610 19834 29622 20410
rect 29656 19834 29668 20410
rect 29610 19822 29668 19834
rect 30628 20410 30686 20422
rect 30628 19834 30640 20410
rect 30674 19834 30686 20410
rect 30628 19822 30686 19834
rect 31646 20410 31704 20422
rect 31646 19834 31658 20410
rect 31692 19834 31704 20410
rect 31646 19822 31704 19834
rect 32664 20410 32722 20422
rect 32664 19834 32676 20410
rect 32710 19834 32722 20410
rect 32664 19822 32722 19834
rect 33682 20410 33740 20422
rect 33682 19834 33694 20410
rect 33728 19834 33740 20410
rect 33682 19822 33740 19834
rect 16744 19574 16802 19586
rect 18412 19154 18470 19166
rect 14564 19024 14622 19036
rect 14564 18648 14576 19024
rect 14610 18648 14622 19024
rect 14564 18636 14622 18648
rect 14782 19024 14840 19036
rect 14782 18648 14794 19024
rect 14828 18648 14840 19024
rect 14782 18636 14840 18648
rect 15000 19024 15058 19036
rect 15000 18648 15012 19024
rect 15046 18648 15058 19024
rect 15000 18636 15058 18648
rect 15218 19024 15276 19036
rect 15218 18648 15230 19024
rect 15264 18648 15276 19024
rect 15218 18636 15276 18648
rect 15436 19024 15494 19036
rect 15436 18648 15448 19024
rect 15482 18648 15494 19024
rect 15436 18636 15494 18648
rect 15654 19024 15712 19036
rect 15654 18648 15666 19024
rect 15700 18648 15712 19024
rect 15654 18636 15712 18648
rect 15872 19024 15930 19036
rect 15872 18648 15884 19024
rect 15918 18648 15930 19024
rect 15872 18636 15930 18648
rect 16090 19024 16148 19036
rect 16090 18648 16102 19024
rect 16136 18648 16148 19024
rect 16090 18636 16148 18648
rect 16308 19024 16366 19036
rect 16308 18648 16320 19024
rect 16354 18648 16366 19024
rect 16308 18636 16366 18648
rect 16526 19024 16584 19036
rect 16526 18648 16538 19024
rect 16572 18648 16584 19024
rect 16526 18636 16584 18648
rect 16744 19024 16802 19036
rect 16744 18648 16756 19024
rect 16790 18648 16802 19024
rect 16744 18636 16802 18648
rect 18412 18578 18424 19154
rect 18458 18578 18470 19154
rect 18412 18566 18470 18578
rect 19430 19154 19488 19166
rect 19430 18578 19442 19154
rect 19476 18578 19488 19154
rect 19430 18566 19488 18578
rect 20448 19154 20506 19166
rect 20448 18578 20460 19154
rect 20494 18578 20506 19154
rect 20448 18566 20506 18578
rect 21466 19154 21524 19166
rect 21466 18578 21478 19154
rect 21512 18578 21524 19154
rect 21466 18566 21524 18578
rect 22484 19154 22542 19166
rect 22484 18578 22496 19154
rect 22530 18578 22542 19154
rect 22484 18566 22542 18578
rect 23502 19154 23560 19166
rect 23502 18578 23514 19154
rect 23548 18578 23560 19154
rect 23502 18566 23560 18578
rect 24520 19154 24578 19166
rect 24520 18578 24532 19154
rect 24566 18578 24578 19154
rect 24520 18566 24578 18578
rect 25538 19154 25596 19166
rect 25538 18578 25550 19154
rect 25584 18578 25596 19154
rect 25538 18566 25596 18578
rect 26556 19154 26614 19166
rect 26556 18578 26568 19154
rect 26602 18578 26614 19154
rect 26556 18566 26614 18578
rect 27574 19154 27632 19166
rect 27574 18578 27586 19154
rect 27620 18578 27632 19154
rect 27574 18566 27632 18578
rect 28592 19154 28650 19166
rect 28592 18578 28604 19154
rect 28638 18578 28650 19154
rect 28592 18566 28650 18578
rect 29610 19154 29668 19166
rect 29610 18578 29622 19154
rect 29656 18578 29668 19154
rect 29610 18566 29668 18578
rect 30628 19154 30686 19166
rect 30628 18578 30640 19154
rect 30674 18578 30686 19154
rect 30628 18566 30686 18578
rect 31646 19154 31704 19166
rect 31646 18578 31658 19154
rect 31692 18578 31704 19154
rect 31646 18566 31704 18578
rect 32664 19154 32722 19166
rect 32664 18578 32676 19154
rect 32710 18578 32722 19154
rect 32664 18566 32722 18578
rect 33682 19154 33740 19166
rect 33682 18578 33694 19154
rect 33728 18578 33740 19154
rect 33682 18566 33740 18578
rect 47366 25216 47424 25228
rect 47366 24840 47378 25216
rect 47412 24840 47424 25216
rect 47366 24828 47424 24840
rect 47624 25216 47682 25228
rect 47624 24840 47636 25216
rect 47670 24840 47682 25216
rect 47624 24828 47682 24840
rect 47882 25216 47940 25228
rect 47882 24840 47894 25216
rect 47928 24840 47940 25216
rect 47882 24828 47940 24840
rect 48140 25216 48198 25228
rect 48140 24840 48152 25216
rect 48186 24840 48198 25216
rect 48140 24828 48198 24840
rect 48398 25216 48456 25228
rect 48398 24840 48410 25216
rect 48444 24840 48456 25216
rect 48398 24828 48456 24840
rect 48656 25216 48714 25228
rect 48656 24840 48668 25216
rect 48702 24840 48714 25216
rect 48656 24828 48714 24840
rect 48914 25216 48972 25228
rect 48914 24840 48926 25216
rect 48960 24840 48972 25216
rect 48914 24828 48972 24840
rect 49222 24833 49274 24845
rect 49222 24799 49230 24833
rect 49264 24799 49274 24833
rect 49222 24765 49274 24799
rect 49222 24731 49230 24765
rect 49264 24731 49274 24765
rect 49222 24697 49274 24731
rect 49222 24663 49230 24697
rect 49264 24663 49274 24697
rect 49222 24645 49274 24663
rect 49304 24833 49356 24845
rect 49304 24799 49314 24833
rect 49348 24799 49356 24833
rect 49304 24765 49356 24799
rect 49304 24731 49314 24765
rect 49348 24731 49356 24765
rect 49304 24697 49356 24731
rect 49304 24663 49314 24697
rect 49348 24663 49356 24697
rect 49304 24645 49356 24663
rect 47366 23216 47424 23228
rect 47366 22840 47378 23216
rect 47412 22840 47424 23216
rect 47366 22828 47424 22840
rect 47624 23216 47682 23228
rect 47624 22840 47636 23216
rect 47670 22840 47682 23216
rect 47624 22828 47682 22840
rect 47882 23216 47940 23228
rect 47882 22840 47894 23216
rect 47928 22840 47940 23216
rect 47882 22828 47940 22840
rect 48140 23216 48198 23228
rect 48140 22840 48152 23216
rect 48186 22840 48198 23216
rect 48140 22828 48198 22840
rect 48398 23216 48456 23228
rect 48398 22840 48410 23216
rect 48444 22840 48456 23216
rect 48398 22828 48456 22840
rect 48656 23216 48714 23228
rect 48656 22840 48668 23216
rect 48702 22840 48714 23216
rect 48656 22828 48714 22840
rect 48914 23216 48972 23228
rect 48914 22840 48926 23216
rect 48960 22840 48972 23216
rect 48914 22828 48972 22840
rect 49222 22833 49274 22845
rect 49222 22799 49230 22833
rect 49264 22799 49274 22833
rect 49222 22765 49274 22799
rect 49222 22731 49230 22765
rect 49264 22731 49274 22765
rect 49222 22697 49274 22731
rect 49222 22663 49230 22697
rect 49264 22663 49274 22697
rect 49222 22645 49274 22663
rect 49304 22833 49356 22845
rect 49304 22799 49314 22833
rect 49348 22799 49356 22833
rect 49304 22765 49356 22799
rect 49304 22731 49314 22765
rect 49348 22731 49356 22765
rect 49304 22697 49356 22731
rect 49304 22663 49314 22697
rect 49348 22663 49356 22697
rect 49304 22645 49356 22663
rect 71426 26968 71484 26980
rect 71426 26392 71438 26968
rect 71472 26392 71484 26968
rect 71426 26380 71484 26392
rect 72444 26968 72502 26980
rect 72444 26392 72456 26968
rect 72490 26392 72502 26968
rect 72444 26380 72502 26392
rect 73462 26968 73520 26980
rect 73462 26392 73474 26968
rect 73508 26392 73520 26968
rect 73462 26380 73520 26392
rect 74480 26968 74538 26980
rect 74480 26392 74492 26968
rect 74526 26392 74538 26968
rect 74480 26380 74538 26392
rect 75498 26968 75556 26980
rect 75498 26392 75510 26968
rect 75544 26392 75556 26968
rect 75498 26380 75556 26392
rect 76516 26968 76574 26980
rect 76516 26392 76528 26968
rect 76562 26392 76574 26968
rect 76516 26380 76574 26392
rect 77534 26968 77592 26980
rect 77534 26392 77546 26968
rect 77580 26392 77592 26968
rect 77534 26380 77592 26392
rect 78552 26968 78610 26980
rect 78552 26392 78564 26968
rect 78598 26392 78610 26968
rect 78552 26380 78610 26392
rect 79570 26968 79628 26980
rect 79570 26392 79582 26968
rect 79616 26392 79628 26968
rect 79570 26380 79628 26392
rect 80588 26968 80646 26980
rect 80588 26392 80600 26968
rect 80634 26392 80646 26968
rect 80588 26380 80646 26392
rect 81606 26968 81664 26980
rect 81606 26392 81618 26968
rect 81652 26392 81664 26968
rect 81606 26380 81664 26392
rect 82624 26968 82682 26980
rect 82624 26392 82636 26968
rect 82670 26392 82682 26968
rect 82624 26380 82682 26392
rect 83642 26968 83700 26980
rect 83642 26392 83654 26968
rect 83688 26392 83700 26968
rect 83642 26380 83700 26392
rect 84660 26968 84718 26980
rect 84660 26392 84672 26968
rect 84706 26392 84718 26968
rect 84660 26380 84718 26392
rect 85678 26968 85736 26980
rect 85678 26392 85690 26968
rect 85724 26392 85736 26968
rect 85678 26380 85736 26392
rect 86696 26968 86754 26980
rect 86696 26392 86708 26968
rect 86742 26392 86754 26968
rect 86696 26380 86754 26392
rect 87714 26968 87772 26980
rect 87714 26392 87726 26968
rect 87760 26392 87772 26968
rect 87714 26380 87772 26392
rect 71426 25832 71484 25844
rect 71426 25256 71438 25832
rect 71472 25256 71484 25832
rect 71426 25244 71484 25256
rect 72444 25832 72502 25844
rect 72444 25256 72456 25832
rect 72490 25256 72502 25832
rect 72444 25244 72502 25256
rect 73462 25832 73520 25844
rect 73462 25256 73474 25832
rect 73508 25256 73520 25832
rect 73462 25244 73520 25256
rect 74480 25832 74538 25844
rect 74480 25256 74492 25832
rect 74526 25256 74538 25832
rect 74480 25244 74538 25256
rect 75498 25832 75556 25844
rect 75498 25256 75510 25832
rect 75544 25256 75556 25832
rect 75498 25244 75556 25256
rect 76516 25832 76574 25844
rect 76516 25256 76528 25832
rect 76562 25256 76574 25832
rect 76516 25244 76574 25256
rect 77534 25832 77592 25844
rect 77534 25256 77546 25832
rect 77580 25256 77592 25832
rect 77534 25244 77592 25256
rect 78552 25832 78610 25844
rect 78552 25256 78564 25832
rect 78598 25256 78610 25832
rect 78552 25244 78610 25256
rect 79570 25832 79628 25844
rect 79570 25256 79582 25832
rect 79616 25256 79628 25832
rect 79570 25244 79628 25256
rect 80588 25832 80646 25844
rect 80588 25256 80600 25832
rect 80634 25256 80646 25832
rect 80588 25244 80646 25256
rect 81606 25832 81664 25844
rect 81606 25256 81618 25832
rect 81652 25256 81664 25832
rect 81606 25244 81664 25256
rect 82624 25832 82682 25844
rect 82624 25256 82636 25832
rect 82670 25256 82682 25832
rect 82624 25244 82682 25256
rect 83642 25832 83700 25844
rect 83642 25256 83654 25832
rect 83688 25256 83700 25832
rect 83642 25244 83700 25256
rect 84660 25832 84718 25844
rect 84660 25256 84672 25832
rect 84706 25256 84718 25832
rect 84660 25244 84718 25256
rect 85678 25832 85736 25844
rect 85678 25256 85690 25832
rect 85724 25256 85736 25832
rect 85678 25244 85736 25256
rect 86696 25832 86754 25844
rect 86696 25256 86708 25832
rect 86742 25256 86754 25832
rect 86696 25244 86754 25256
rect 87714 25832 87772 25844
rect 87714 25256 87726 25832
rect 87760 25256 87772 25832
rect 87714 25244 87772 25256
rect 71426 24696 71484 24708
rect 71426 24120 71438 24696
rect 71472 24120 71484 24696
rect 71426 24108 71484 24120
rect 72444 24696 72502 24708
rect 72444 24120 72456 24696
rect 72490 24120 72502 24696
rect 72444 24108 72502 24120
rect 73462 24696 73520 24708
rect 73462 24120 73474 24696
rect 73508 24120 73520 24696
rect 73462 24108 73520 24120
rect 74480 24696 74538 24708
rect 74480 24120 74492 24696
rect 74526 24120 74538 24696
rect 74480 24108 74538 24120
rect 75498 24696 75556 24708
rect 75498 24120 75510 24696
rect 75544 24120 75556 24696
rect 75498 24108 75556 24120
rect 76516 24696 76574 24708
rect 76516 24120 76528 24696
rect 76562 24120 76574 24696
rect 76516 24108 76574 24120
rect 77534 24696 77592 24708
rect 77534 24120 77546 24696
rect 77580 24120 77592 24696
rect 77534 24108 77592 24120
rect 78552 24696 78610 24708
rect 78552 24120 78564 24696
rect 78598 24120 78610 24696
rect 78552 24108 78610 24120
rect 79570 24696 79628 24708
rect 79570 24120 79582 24696
rect 79616 24120 79628 24696
rect 79570 24108 79628 24120
rect 80588 24696 80646 24708
rect 80588 24120 80600 24696
rect 80634 24120 80646 24696
rect 80588 24108 80646 24120
rect 81606 24696 81664 24708
rect 81606 24120 81618 24696
rect 81652 24120 81664 24696
rect 81606 24108 81664 24120
rect 82624 24696 82682 24708
rect 82624 24120 82636 24696
rect 82670 24120 82682 24696
rect 82624 24108 82682 24120
rect 83642 24696 83700 24708
rect 83642 24120 83654 24696
rect 83688 24120 83700 24696
rect 83642 24108 83700 24120
rect 84660 24696 84718 24708
rect 84660 24120 84672 24696
rect 84706 24120 84718 24696
rect 84660 24108 84718 24120
rect 85678 24696 85736 24708
rect 85678 24120 85690 24696
rect 85724 24120 85736 24696
rect 85678 24108 85736 24120
rect 86696 24696 86754 24708
rect 86696 24120 86708 24696
rect 86742 24120 86754 24696
rect 86696 24108 86754 24120
rect 87714 24696 87772 24708
rect 87714 24120 87726 24696
rect 87760 24120 87772 24696
rect 87714 24108 87772 24120
rect 72412 22922 72470 22934
rect 72412 22346 72424 22922
rect 72458 22346 72470 22922
rect 72412 22334 72470 22346
rect 73430 22922 73488 22934
rect 73430 22346 73442 22922
rect 73476 22346 73488 22922
rect 73430 22334 73488 22346
rect 74448 22922 74506 22934
rect 74448 22346 74460 22922
rect 74494 22346 74506 22922
rect 74448 22334 74506 22346
rect 75466 22922 75524 22934
rect 75466 22346 75478 22922
rect 75512 22346 75524 22922
rect 75466 22334 75524 22346
rect 76484 22922 76542 22934
rect 76484 22346 76496 22922
rect 76530 22346 76542 22922
rect 76484 22334 76542 22346
rect 77502 22922 77560 22934
rect 77502 22346 77514 22922
rect 77548 22346 77560 22922
rect 77502 22334 77560 22346
rect 78520 22922 78578 22934
rect 78520 22346 78532 22922
rect 78566 22346 78578 22922
rect 78520 22334 78578 22346
rect 79538 22922 79596 22934
rect 79538 22346 79550 22922
rect 79584 22346 79596 22922
rect 79538 22334 79596 22346
rect 80556 22922 80614 22934
rect 80556 22346 80568 22922
rect 80602 22346 80614 22922
rect 80556 22334 80614 22346
rect 81574 22922 81632 22934
rect 81574 22346 81586 22922
rect 81620 22346 81632 22922
rect 81574 22334 81632 22346
rect 82592 22922 82650 22934
rect 82592 22346 82604 22922
rect 82638 22346 82650 22922
rect 82592 22334 82650 22346
rect 83610 22922 83668 22934
rect 83610 22346 83622 22922
rect 83656 22346 83668 22922
rect 83610 22334 83668 22346
rect 84628 22922 84686 22934
rect 84628 22346 84640 22922
rect 84674 22346 84686 22922
rect 84628 22334 84686 22346
rect 85646 22922 85704 22934
rect 85646 22346 85658 22922
rect 85692 22346 85704 22922
rect 85646 22334 85704 22346
rect 86664 22922 86722 22934
rect 86664 22346 86676 22922
rect 86710 22346 86722 22922
rect 86664 22334 86722 22346
rect 87682 22922 87740 22934
rect 87682 22346 87694 22922
rect 87728 22346 87740 22922
rect 87682 22334 87740 22346
rect 68564 21838 68622 21850
rect 68564 21462 68576 21838
rect 68610 21462 68622 21838
rect 68564 21450 68622 21462
rect 68782 21838 68840 21850
rect 68782 21462 68794 21838
rect 68828 21462 68840 21838
rect 68782 21450 68840 21462
rect 69000 21838 69058 21850
rect 69000 21462 69012 21838
rect 69046 21462 69058 21838
rect 69000 21450 69058 21462
rect 69218 21838 69276 21850
rect 69218 21462 69230 21838
rect 69264 21462 69276 21838
rect 69218 21450 69276 21462
rect 69436 21838 69494 21850
rect 69436 21462 69448 21838
rect 69482 21462 69494 21838
rect 69436 21450 69494 21462
rect 69654 21838 69712 21850
rect 69654 21462 69666 21838
rect 69700 21462 69712 21838
rect 69654 21450 69712 21462
rect 69872 21838 69930 21850
rect 69872 21462 69884 21838
rect 69918 21462 69930 21838
rect 69872 21450 69930 21462
rect 70090 21838 70148 21850
rect 70090 21462 70102 21838
rect 70136 21462 70148 21838
rect 70090 21450 70148 21462
rect 70308 21838 70366 21850
rect 70308 21462 70320 21838
rect 70354 21462 70366 21838
rect 70308 21450 70366 21462
rect 70526 21838 70584 21850
rect 70526 21462 70538 21838
rect 70572 21462 70584 21838
rect 70526 21450 70584 21462
rect 70744 21838 70802 21850
rect 70744 21462 70756 21838
rect 70790 21462 70802 21838
rect 70744 21450 70802 21462
rect 72412 21666 72470 21678
rect 72412 21090 72424 21666
rect 72458 21090 72470 21666
rect 72412 21078 72470 21090
rect 73430 21666 73488 21678
rect 73430 21090 73442 21666
rect 73476 21090 73488 21666
rect 73430 21078 73488 21090
rect 74448 21666 74506 21678
rect 74448 21090 74460 21666
rect 74494 21090 74506 21666
rect 74448 21078 74506 21090
rect 75466 21666 75524 21678
rect 75466 21090 75478 21666
rect 75512 21090 75524 21666
rect 75466 21078 75524 21090
rect 76484 21666 76542 21678
rect 76484 21090 76496 21666
rect 76530 21090 76542 21666
rect 76484 21078 76542 21090
rect 77502 21666 77560 21678
rect 77502 21090 77514 21666
rect 77548 21090 77560 21666
rect 77502 21078 77560 21090
rect 78520 21666 78578 21678
rect 78520 21090 78532 21666
rect 78566 21090 78578 21666
rect 78520 21078 78578 21090
rect 79538 21666 79596 21678
rect 79538 21090 79550 21666
rect 79584 21090 79596 21666
rect 79538 21078 79596 21090
rect 80556 21666 80614 21678
rect 80556 21090 80568 21666
rect 80602 21090 80614 21666
rect 80556 21078 80614 21090
rect 81574 21666 81632 21678
rect 81574 21090 81586 21666
rect 81620 21090 81632 21666
rect 81574 21078 81632 21090
rect 82592 21666 82650 21678
rect 82592 21090 82604 21666
rect 82638 21090 82650 21666
rect 82592 21078 82650 21090
rect 83610 21666 83668 21678
rect 83610 21090 83622 21666
rect 83656 21090 83668 21666
rect 83610 21078 83668 21090
rect 84628 21666 84686 21678
rect 84628 21090 84640 21666
rect 84674 21090 84686 21666
rect 84628 21078 84686 21090
rect 85646 21666 85704 21678
rect 85646 21090 85658 21666
rect 85692 21090 85704 21666
rect 85646 21078 85704 21090
rect 86664 21666 86722 21678
rect 86664 21090 86676 21666
rect 86710 21090 86722 21666
rect 86664 21078 86722 21090
rect 87682 21666 87740 21678
rect 87682 21090 87694 21666
rect 87728 21090 87740 21666
rect 87682 21078 87740 21090
rect 68564 20900 68622 20912
rect 68564 20524 68576 20900
rect 68610 20524 68622 20900
rect 68564 20512 68622 20524
rect 68782 20900 68840 20912
rect 68782 20524 68794 20900
rect 68828 20524 68840 20900
rect 68782 20512 68840 20524
rect 69000 20900 69058 20912
rect 69000 20524 69012 20900
rect 69046 20524 69058 20900
rect 69000 20512 69058 20524
rect 69218 20900 69276 20912
rect 69218 20524 69230 20900
rect 69264 20524 69276 20900
rect 69218 20512 69276 20524
rect 69436 20900 69494 20912
rect 69436 20524 69448 20900
rect 69482 20524 69494 20900
rect 69436 20512 69494 20524
rect 69654 20900 69712 20912
rect 69654 20524 69666 20900
rect 69700 20524 69712 20900
rect 69654 20512 69712 20524
rect 69872 20900 69930 20912
rect 69872 20524 69884 20900
rect 69918 20524 69930 20900
rect 69872 20512 69930 20524
rect 70090 20900 70148 20912
rect 70090 20524 70102 20900
rect 70136 20524 70148 20900
rect 70090 20512 70148 20524
rect 70308 20900 70366 20912
rect 70308 20524 70320 20900
rect 70354 20524 70366 20900
rect 70308 20512 70366 20524
rect 70526 20900 70584 20912
rect 70526 20524 70538 20900
rect 70572 20524 70584 20900
rect 70526 20512 70584 20524
rect 70744 20900 70802 20912
rect 70744 20524 70756 20900
rect 70790 20524 70802 20900
rect 70744 20512 70802 20524
rect 72412 20410 72470 20422
rect 68564 19962 68622 19974
rect 68564 19586 68576 19962
rect 68610 19586 68622 19962
rect 68564 19574 68622 19586
rect 68782 19962 68840 19974
rect 68782 19586 68794 19962
rect 68828 19586 68840 19962
rect 68782 19574 68840 19586
rect 69000 19962 69058 19974
rect 69000 19586 69012 19962
rect 69046 19586 69058 19962
rect 69000 19574 69058 19586
rect 69218 19962 69276 19974
rect 69218 19586 69230 19962
rect 69264 19586 69276 19962
rect 69218 19574 69276 19586
rect 69436 19962 69494 19974
rect 69436 19586 69448 19962
rect 69482 19586 69494 19962
rect 69436 19574 69494 19586
rect 69654 19962 69712 19974
rect 69654 19586 69666 19962
rect 69700 19586 69712 19962
rect 69654 19574 69712 19586
rect 69872 19962 69930 19974
rect 69872 19586 69884 19962
rect 69918 19586 69930 19962
rect 69872 19574 69930 19586
rect 70090 19962 70148 19974
rect 70090 19586 70102 19962
rect 70136 19586 70148 19962
rect 70090 19574 70148 19586
rect 70308 19962 70366 19974
rect 70308 19586 70320 19962
rect 70354 19586 70366 19962
rect 70308 19574 70366 19586
rect 70526 19962 70584 19974
rect 70526 19586 70538 19962
rect 70572 19586 70584 19962
rect 70526 19574 70584 19586
rect 70744 19962 70802 19974
rect 70744 19586 70756 19962
rect 70790 19586 70802 19962
rect 72412 19834 72424 20410
rect 72458 19834 72470 20410
rect 72412 19822 72470 19834
rect 73430 20410 73488 20422
rect 73430 19834 73442 20410
rect 73476 19834 73488 20410
rect 73430 19822 73488 19834
rect 74448 20410 74506 20422
rect 74448 19834 74460 20410
rect 74494 19834 74506 20410
rect 74448 19822 74506 19834
rect 75466 20410 75524 20422
rect 75466 19834 75478 20410
rect 75512 19834 75524 20410
rect 75466 19822 75524 19834
rect 76484 20410 76542 20422
rect 76484 19834 76496 20410
rect 76530 19834 76542 20410
rect 76484 19822 76542 19834
rect 77502 20410 77560 20422
rect 77502 19834 77514 20410
rect 77548 19834 77560 20410
rect 77502 19822 77560 19834
rect 78520 20410 78578 20422
rect 78520 19834 78532 20410
rect 78566 19834 78578 20410
rect 78520 19822 78578 19834
rect 79538 20410 79596 20422
rect 79538 19834 79550 20410
rect 79584 19834 79596 20410
rect 79538 19822 79596 19834
rect 80556 20410 80614 20422
rect 80556 19834 80568 20410
rect 80602 19834 80614 20410
rect 80556 19822 80614 19834
rect 81574 20410 81632 20422
rect 81574 19834 81586 20410
rect 81620 19834 81632 20410
rect 81574 19822 81632 19834
rect 82592 20410 82650 20422
rect 82592 19834 82604 20410
rect 82638 19834 82650 20410
rect 82592 19822 82650 19834
rect 83610 20410 83668 20422
rect 83610 19834 83622 20410
rect 83656 19834 83668 20410
rect 83610 19822 83668 19834
rect 84628 20410 84686 20422
rect 84628 19834 84640 20410
rect 84674 19834 84686 20410
rect 84628 19822 84686 19834
rect 85646 20410 85704 20422
rect 85646 19834 85658 20410
rect 85692 19834 85704 20410
rect 85646 19822 85704 19834
rect 86664 20410 86722 20422
rect 86664 19834 86676 20410
rect 86710 19834 86722 20410
rect 86664 19822 86722 19834
rect 87682 20410 87740 20422
rect 87682 19834 87694 20410
rect 87728 19834 87740 20410
rect 87682 19822 87740 19834
rect 70744 19574 70802 19586
rect 72412 19154 72470 19166
rect 68564 19024 68622 19036
rect 68564 18648 68576 19024
rect 68610 18648 68622 19024
rect 68564 18636 68622 18648
rect 68782 19024 68840 19036
rect 68782 18648 68794 19024
rect 68828 18648 68840 19024
rect 68782 18636 68840 18648
rect 69000 19024 69058 19036
rect 69000 18648 69012 19024
rect 69046 18648 69058 19024
rect 69000 18636 69058 18648
rect 69218 19024 69276 19036
rect 69218 18648 69230 19024
rect 69264 18648 69276 19024
rect 69218 18636 69276 18648
rect 69436 19024 69494 19036
rect 69436 18648 69448 19024
rect 69482 18648 69494 19024
rect 69436 18636 69494 18648
rect 69654 19024 69712 19036
rect 69654 18648 69666 19024
rect 69700 18648 69712 19024
rect 69654 18636 69712 18648
rect 69872 19024 69930 19036
rect 69872 18648 69884 19024
rect 69918 18648 69930 19024
rect 69872 18636 69930 18648
rect 70090 19024 70148 19036
rect 70090 18648 70102 19024
rect 70136 18648 70148 19024
rect 70090 18636 70148 18648
rect 70308 19024 70366 19036
rect 70308 18648 70320 19024
rect 70354 18648 70366 19024
rect 70308 18636 70366 18648
rect 70526 19024 70584 19036
rect 70526 18648 70538 19024
rect 70572 18648 70584 19024
rect 70526 18636 70584 18648
rect 70744 19024 70802 19036
rect 70744 18648 70756 19024
rect 70790 18648 70802 19024
rect 70744 18636 70802 18648
rect 72412 18578 72424 19154
rect 72458 18578 72470 19154
rect 72412 18566 72470 18578
rect 73430 19154 73488 19166
rect 73430 18578 73442 19154
rect 73476 18578 73488 19154
rect 73430 18566 73488 18578
rect 74448 19154 74506 19166
rect 74448 18578 74460 19154
rect 74494 18578 74506 19154
rect 74448 18566 74506 18578
rect 75466 19154 75524 19166
rect 75466 18578 75478 19154
rect 75512 18578 75524 19154
rect 75466 18566 75524 18578
rect 76484 19154 76542 19166
rect 76484 18578 76496 19154
rect 76530 18578 76542 19154
rect 76484 18566 76542 18578
rect 77502 19154 77560 19166
rect 77502 18578 77514 19154
rect 77548 18578 77560 19154
rect 77502 18566 77560 18578
rect 78520 19154 78578 19166
rect 78520 18578 78532 19154
rect 78566 18578 78578 19154
rect 78520 18566 78578 18578
rect 79538 19154 79596 19166
rect 79538 18578 79550 19154
rect 79584 18578 79596 19154
rect 79538 18566 79596 18578
rect 80556 19154 80614 19166
rect 80556 18578 80568 19154
rect 80602 18578 80614 19154
rect 80556 18566 80614 18578
rect 81574 19154 81632 19166
rect 81574 18578 81586 19154
rect 81620 18578 81632 19154
rect 81574 18566 81632 18578
rect 82592 19154 82650 19166
rect 82592 18578 82604 19154
rect 82638 18578 82650 19154
rect 82592 18566 82650 18578
rect 83610 19154 83668 19166
rect 83610 18578 83622 19154
rect 83656 18578 83668 19154
rect 83610 18566 83668 18578
rect 84628 19154 84686 19166
rect 84628 18578 84640 19154
rect 84674 18578 84686 19154
rect 84628 18566 84686 18578
rect 85646 19154 85704 19166
rect 85646 18578 85658 19154
rect 85692 18578 85704 19154
rect 85646 18566 85704 18578
rect 86664 19154 86722 19166
rect 86664 18578 86676 19154
rect 86710 18578 86722 19154
rect 86664 18566 86722 18578
rect 87682 19154 87740 19166
rect 87682 18578 87694 19154
rect 87728 18578 87740 19154
rect 87682 18566 87740 18578
rect -12992 16086 -12934 16098
rect -12992 15710 -12980 16086
rect -12946 15710 -12934 16086
rect -12992 15698 -12934 15710
rect -12734 16086 -12676 16098
rect -12734 15710 -12722 16086
rect -12688 15710 -12676 16086
rect -12734 15698 -12676 15710
rect -12476 16086 -12418 16098
rect -12476 15710 -12464 16086
rect -12430 15710 -12418 16086
rect -12476 15698 -12418 15710
rect -12218 16086 -12160 16098
rect -12218 15710 -12206 16086
rect -12172 15710 -12160 16086
rect -12218 15698 -12160 15710
rect -11960 16086 -11902 16098
rect -11960 15710 -11948 16086
rect -11914 15710 -11902 16086
rect -11960 15698 -11902 15710
rect -11702 16086 -11644 16098
rect -11702 15710 -11690 16086
rect -11656 15710 -11644 16086
rect -11702 15698 -11644 15710
rect -11444 16086 -11386 16098
rect -11444 15710 -11432 16086
rect -11398 15710 -11386 16086
rect -11444 15698 -11386 15710
rect -11136 15703 -11084 15715
rect -11136 15669 -11128 15703
rect -11094 15669 -11084 15703
rect -11136 15635 -11084 15669
rect -11136 15601 -11128 15635
rect -11094 15601 -11084 15635
rect -11136 15567 -11084 15601
rect -11136 15533 -11128 15567
rect -11094 15533 -11084 15567
rect -11136 15515 -11084 15533
rect -11054 15703 -11002 15715
rect -11054 15669 -11044 15703
rect -11010 15669 -11002 15703
rect -11054 15635 -11002 15669
rect -11054 15601 -11044 15635
rect -11010 15601 -11002 15635
rect -11054 15567 -11002 15601
rect -11054 15533 -11044 15567
rect -11010 15533 -11002 15567
rect -11054 15515 -11002 15533
rect -10392 16086 -10334 16098
rect -10392 15710 -10380 16086
rect -10346 15710 -10334 16086
rect -10392 15698 -10334 15710
rect -10134 16086 -10076 16098
rect -10134 15710 -10122 16086
rect -10088 15710 -10076 16086
rect -10134 15698 -10076 15710
rect -9876 16086 -9818 16098
rect -9876 15710 -9864 16086
rect -9830 15710 -9818 16086
rect -9876 15698 -9818 15710
rect -9618 16086 -9560 16098
rect -9618 15710 -9606 16086
rect -9572 15710 -9560 16086
rect -9618 15698 -9560 15710
rect -9360 16086 -9302 16098
rect -9360 15710 -9348 16086
rect -9314 15710 -9302 16086
rect -9360 15698 -9302 15710
rect -9102 16086 -9044 16098
rect -9102 15710 -9090 16086
rect -9056 15710 -9044 16086
rect -9102 15698 -9044 15710
rect -8844 16086 -8786 16098
rect -8844 15710 -8832 16086
rect -8798 15710 -8786 16086
rect -8844 15698 -8786 15710
rect -8536 15703 -8484 15715
rect -8536 15669 -8528 15703
rect -8494 15669 -8484 15703
rect -8536 15635 -8484 15669
rect -8536 15601 -8528 15635
rect -8494 15601 -8484 15635
rect -8536 15567 -8484 15601
rect -8536 15533 -8528 15567
rect -8494 15533 -8484 15567
rect -8536 15515 -8484 15533
rect -8454 15703 -8402 15715
rect -8454 15669 -8444 15703
rect -8410 15669 -8402 15703
rect -8454 15635 -8402 15669
rect -8454 15601 -8444 15635
rect -8410 15601 -8402 15635
rect -8454 15567 -8402 15601
rect -8454 15533 -8444 15567
rect -8410 15533 -8402 15567
rect -8454 15515 -8402 15533
rect -8036 15703 -7984 15715
rect -8036 15669 -8028 15703
rect -7994 15669 -7984 15703
rect -8036 15635 -7984 15669
rect -8036 15601 -8028 15635
rect -7994 15601 -7984 15635
rect -8036 15567 -7984 15601
rect -8036 15533 -8028 15567
rect -7994 15533 -7984 15567
rect -8036 15515 -7984 15533
rect -7954 15703 -7902 15715
rect -7954 15669 -7944 15703
rect -7910 15669 -7902 15703
rect -7954 15635 -7902 15669
rect -7954 15601 -7944 15635
rect -7910 15601 -7902 15635
rect -7954 15567 -7902 15601
rect -7954 15533 -7944 15567
rect -7910 15533 -7902 15567
rect -7954 15515 -7902 15533
rect 48792 8252 48850 8264
rect 48792 7876 48804 8252
rect 48838 7876 48850 8252
rect 48792 7864 48850 7876
rect 49050 8252 49108 8264
rect 49050 7876 49062 8252
rect 49096 7876 49108 8252
rect 49050 7864 49108 7876
rect 49308 8252 49366 8264
rect 49308 7876 49320 8252
rect 49354 7876 49366 8252
rect 49308 7864 49366 7876
rect 49566 8252 49624 8264
rect 49566 7876 49578 8252
rect 49612 7876 49624 8252
rect 49566 7864 49624 7876
rect 49824 8252 49882 8264
rect 49824 7876 49836 8252
rect 49870 7876 49882 8252
rect 49824 7864 49882 7876
rect 50082 8252 50140 8264
rect 50082 7876 50094 8252
rect 50128 7876 50140 8252
rect 50082 7864 50140 7876
rect 50340 8252 50398 8264
rect 50340 7876 50352 8252
rect 50386 7876 50398 8252
rect 50340 7864 50398 7876
rect 50648 7869 50700 7881
rect 50648 7835 50656 7869
rect 50690 7835 50700 7869
rect 50648 7801 50700 7835
rect 50648 7767 50656 7801
rect 50690 7767 50700 7801
rect 50648 7733 50700 7767
rect 50648 7699 50656 7733
rect 50690 7699 50700 7733
rect 50648 7681 50700 7699
rect 50730 7869 50782 7881
rect 50730 7835 50740 7869
rect 50774 7835 50782 7869
rect 50730 7801 50782 7835
rect 50730 7767 50740 7801
rect 50774 7767 50782 7801
rect 50730 7733 50782 7767
rect 50730 7699 50740 7733
rect 50774 7699 50782 7733
rect 50730 7681 50782 7699
rect 48792 6288 48850 6300
rect 48792 5912 48804 6288
rect 48838 5912 48850 6288
rect 48792 5900 48850 5912
rect 49050 6288 49108 6300
rect 49050 5912 49062 6288
rect 49096 5912 49108 6288
rect 49050 5900 49108 5912
rect 49308 6288 49366 6300
rect 49308 5912 49320 6288
rect 49354 5912 49366 6288
rect 49308 5900 49366 5912
rect 49566 6288 49624 6300
rect 49566 5912 49578 6288
rect 49612 5912 49624 6288
rect 49566 5900 49624 5912
rect 49824 6288 49882 6300
rect 49824 5912 49836 6288
rect 49870 5912 49882 6288
rect 49824 5900 49882 5912
rect 50082 6288 50140 6300
rect 50082 5912 50094 6288
rect 50128 5912 50140 6288
rect 50082 5900 50140 5912
rect 50340 6288 50398 6300
rect 50340 5912 50352 6288
rect 50386 5912 50398 6288
rect 50340 5900 50398 5912
rect 50648 5905 50700 5917
rect 50648 5871 50656 5905
rect 50690 5871 50700 5905
rect 50648 5837 50700 5871
rect 50648 5803 50656 5837
rect 50690 5803 50700 5837
rect 50648 5769 50700 5803
rect 50648 5735 50656 5769
rect 50690 5735 50700 5769
rect 50648 5717 50700 5735
rect 50730 5905 50782 5917
rect 50730 5871 50740 5905
rect 50774 5871 50782 5905
rect 50730 5837 50782 5871
rect 50730 5803 50740 5837
rect 50774 5803 50782 5837
rect 50730 5769 50782 5803
rect 50730 5735 50740 5769
rect 50774 5735 50782 5769
rect 50730 5717 50782 5735
rect 48792 4288 48850 4300
rect 48792 3912 48804 4288
rect 48838 3912 48850 4288
rect 48792 3900 48850 3912
rect 49050 4288 49108 4300
rect 49050 3912 49062 4288
rect 49096 3912 49108 4288
rect 49050 3900 49108 3912
rect 49308 4288 49366 4300
rect 49308 3912 49320 4288
rect 49354 3912 49366 4288
rect 49308 3900 49366 3912
rect 49566 4288 49624 4300
rect 49566 3912 49578 4288
rect 49612 3912 49624 4288
rect 49566 3900 49624 3912
rect 49824 4288 49882 4300
rect 49824 3912 49836 4288
rect 49870 3912 49882 4288
rect 49824 3900 49882 3912
rect 50082 4288 50140 4300
rect 50082 3912 50094 4288
rect 50128 3912 50140 4288
rect 50082 3900 50140 3912
rect 50340 4288 50398 4300
rect 50340 3912 50352 4288
rect 50386 3912 50398 4288
rect 50340 3900 50398 3912
rect 50648 3905 50700 3917
rect 50648 3871 50656 3905
rect 50690 3871 50700 3905
rect 50648 3837 50700 3871
rect 50648 3803 50656 3837
rect 50690 3803 50700 3837
rect 50648 3769 50700 3803
rect 50648 3735 50656 3769
rect 50690 3735 50700 3769
rect 50648 3717 50700 3735
rect 50730 3905 50782 3917
rect 50730 3871 50740 3905
rect 50774 3871 50782 3905
rect 50730 3837 50782 3871
rect 50730 3803 50740 3837
rect 50774 3803 50782 3837
rect 50730 3769 50782 3803
rect 50730 3735 50740 3769
rect 50774 3735 50782 3769
rect 50730 3717 50782 3735
rect 48792 2198 48850 2210
rect 48792 1822 48804 2198
rect 48838 1822 48850 2198
rect 48792 1810 48850 1822
rect 49050 2198 49108 2210
rect 49050 1822 49062 2198
rect 49096 1822 49108 2198
rect 49050 1810 49108 1822
rect 49308 2198 49366 2210
rect 49308 1822 49320 2198
rect 49354 1822 49366 2198
rect 49308 1810 49366 1822
rect 49566 2198 49624 2210
rect 49566 1822 49578 2198
rect 49612 1822 49624 2198
rect 49566 1810 49624 1822
rect 49824 2198 49882 2210
rect 49824 1822 49836 2198
rect 49870 1822 49882 2198
rect 49824 1810 49882 1822
rect 50082 2198 50140 2210
rect 50082 1822 50094 2198
rect 50128 1822 50140 2198
rect 50082 1810 50140 1822
rect 50340 2198 50398 2210
rect 50340 1822 50352 2198
rect 50386 1822 50398 2198
rect 50340 1810 50398 1822
rect 50648 1815 50700 1827
rect 50648 1781 50656 1815
rect 50690 1781 50700 1815
rect 50648 1747 50700 1781
rect 50648 1713 50656 1747
rect 50690 1713 50700 1747
rect 50648 1679 50700 1713
rect 50648 1645 50656 1679
rect 50690 1645 50700 1679
rect 50648 1627 50700 1645
rect 50730 1815 50782 1827
rect 50730 1781 50740 1815
rect 50774 1781 50782 1815
rect 50730 1747 50782 1781
rect 50730 1713 50740 1747
rect 50774 1713 50782 1747
rect 50730 1679 50782 1713
rect 50730 1645 50740 1679
rect 50774 1645 50782 1679
rect 50730 1627 50782 1645
<< ndiffc >>
rect 49230 24479 49264 24513
rect 49230 24411 49264 24445
rect 49314 24479 49348 24513
rect 49314 24411 49348 24445
rect 47378 24116 47412 24292
rect 47636 24116 47670 24292
rect 47894 24116 47928 24292
rect 48152 24116 48186 24292
rect 48410 24116 48444 24292
rect 48668 24116 48702 24292
rect 48926 24116 48960 24292
rect 49230 22479 49264 22513
rect 49230 22411 49264 22445
rect 49314 22479 49348 22513
rect 49314 22411 49348 22445
rect 47378 22116 47412 22292
rect 47636 22116 47670 22292
rect 47894 22116 47928 22292
rect 48152 22116 48186 22292
rect 48410 22116 48444 22292
rect 48668 22116 48702 22292
rect 48926 22116 48960 22292
rect -11128 15349 -11094 15383
rect -11128 15281 -11094 15315
rect -11044 15349 -11010 15383
rect -8528 15349 -8494 15383
rect -11044 15281 -11010 15315
rect -12980 14986 -12946 15162
rect -12722 14986 -12688 15162
rect -12464 14986 -12430 15162
rect -12206 14986 -12172 15162
rect -11948 14986 -11914 15162
rect -11690 14986 -11656 15162
rect -11432 14986 -11398 15162
rect -8528 15281 -8494 15315
rect -8444 15349 -8410 15383
rect -8444 15281 -8410 15315
rect -8028 15349 -7994 15383
rect -8028 15281 -7994 15315
rect -7944 15349 -7910 15383
rect -7944 15281 -7910 15315
rect -10380 14986 -10346 15162
rect -10122 14986 -10088 15162
rect -9864 14986 -9830 15162
rect -9606 14986 -9572 15162
rect -9348 14986 -9314 15162
rect -9090 14986 -9056 15162
rect -8832 14986 -8798 15162
rect 13532 14234 13566 14810
rect 14550 14234 14584 14810
rect 15568 14234 15602 14810
rect 16586 14234 16620 14810
rect 17604 14234 17638 14810
rect 18622 14234 18656 14810
rect 19640 14234 19674 14810
rect 20658 14234 20692 14810
rect 21676 14234 21710 14810
rect 22694 14234 22728 14810
rect 23712 14234 23746 14810
rect 24730 14234 24764 14810
rect 25748 14234 25782 14810
rect 26766 14234 26800 14810
rect 27784 14234 27818 14810
rect 28802 14234 28836 14810
rect 29820 14234 29854 14810
rect 30838 14234 30872 14810
rect 31856 14234 31890 14810
rect 32874 14234 32908 14810
rect 33892 14234 33926 14810
rect 1766 13440 1800 14016
rect 2784 13440 2818 14016
rect 3802 13440 3836 14016
rect 4820 13440 4854 14016
rect 5838 13440 5872 14016
rect 6856 13440 6890 14016
rect 7874 13440 7908 14016
rect 8892 13440 8926 14016
rect 9910 13440 9944 14016
rect 10928 13440 10962 14016
rect 1766 12622 1800 13198
rect 2784 12622 2818 13198
rect 3802 12622 3836 13198
rect 4820 12622 4854 13198
rect 5838 12622 5872 13198
rect 6856 12622 6890 13198
rect 7874 12622 7908 13198
rect 8892 12622 8926 13198
rect 9910 12622 9944 13198
rect 10928 12622 10962 13198
rect 13532 13000 13566 13576
rect 14550 13000 14584 13576
rect 15568 13000 15602 13576
rect 16586 13000 16620 13576
rect 17604 13000 17638 13576
rect 18622 13000 18656 13576
rect 19640 13000 19674 13576
rect 20658 13000 20692 13576
rect 21676 13000 21710 13576
rect 22694 13000 22728 13576
rect 23712 13000 23746 13576
rect 24730 13000 24764 13576
rect 25748 13000 25782 13576
rect 26766 13000 26800 13576
rect 27784 13000 27818 13576
rect 28802 13000 28836 13576
rect 29820 13000 29854 13576
rect 30838 13000 30872 13576
rect 31856 13000 31890 13576
rect 32874 13000 32908 13576
rect 33892 13000 33926 13576
rect 1766 11804 1800 12380
rect 2784 11804 2818 12380
rect 3802 11804 3836 12380
rect 4820 11804 4854 12380
rect 5838 11804 5872 12380
rect 6856 11804 6890 12380
rect 7874 11804 7908 12380
rect 8892 11804 8926 12380
rect 9910 11804 9944 12380
rect 10928 11804 10962 12380
rect 13532 11768 13566 12344
rect 14550 11768 14584 12344
rect 15568 11768 15602 12344
rect 16586 11768 16620 12344
rect 17604 11768 17638 12344
rect 18622 11768 18656 12344
rect 19640 11768 19674 12344
rect 20658 11768 20692 12344
rect 21676 11768 21710 12344
rect 22694 11768 22728 12344
rect 23712 11768 23746 12344
rect 24730 11768 24764 12344
rect 25748 11768 25782 12344
rect 26766 11768 26800 12344
rect 27784 11768 27818 12344
rect 28802 11768 28836 12344
rect 29820 11768 29854 12344
rect 30838 11768 30872 12344
rect 31856 11768 31890 12344
rect 32874 11768 32908 12344
rect 33892 11768 33926 12344
rect 1766 10986 1800 11562
rect 2784 10986 2818 11562
rect 3802 10986 3836 11562
rect 4820 10986 4854 11562
rect 5838 10986 5872 11562
rect 6856 10986 6890 11562
rect 7874 10986 7908 11562
rect 8892 10986 8926 11562
rect 9910 10986 9944 11562
rect 10928 10986 10962 11562
rect 1766 10168 1800 10744
rect 2784 10168 2818 10744
rect 3802 10168 3836 10744
rect 4820 10168 4854 10744
rect 5838 10168 5872 10744
rect 6856 10168 6890 10744
rect 7874 10168 7908 10744
rect 8892 10168 8926 10744
rect 9910 10168 9944 10744
rect 10928 10168 10962 10744
rect 13530 10534 13564 11110
rect 14548 10534 14582 11110
rect 15566 10534 15600 11110
rect 16584 10534 16618 11110
rect 17602 10534 17636 11110
rect 18620 10534 18654 11110
rect 19638 10534 19672 11110
rect 20656 10534 20690 11110
rect 21674 10534 21708 11110
rect 22692 10534 22726 11110
rect 23710 10534 23744 11110
rect 24728 10534 24762 11110
rect 25746 10534 25780 11110
rect 26764 10534 26798 11110
rect 27782 10534 27816 11110
rect 28800 10534 28834 11110
rect 29818 10534 29852 11110
rect 30836 10534 30870 11110
rect 31854 10534 31888 11110
rect 32872 10534 32906 11110
rect 33890 10534 33924 11110
rect 1766 9350 1800 9926
rect 2784 9350 2818 9926
rect 3802 9350 3836 9926
rect 4820 9350 4854 9926
rect 5838 9350 5872 9926
rect 6856 9350 6890 9926
rect 7874 9350 7908 9926
rect 8892 9350 8926 9926
rect 9910 9350 9944 9926
rect 10928 9350 10962 9926
rect 13530 9300 13564 9876
rect 14548 9300 14582 9876
rect 15566 9300 15600 9876
rect 16584 9300 16618 9876
rect 17602 9300 17636 9876
rect 18620 9300 18654 9876
rect 19638 9300 19672 9876
rect 20656 9300 20690 9876
rect 21674 9300 21708 9876
rect 22692 9300 22726 9876
rect 23710 9300 23744 9876
rect 24728 9300 24762 9876
rect 25746 9300 25780 9876
rect 26764 9300 26798 9876
rect 27782 9300 27816 9876
rect 28800 9300 28834 9876
rect 29818 9300 29852 9876
rect 30836 9300 30870 9876
rect 31854 9300 31888 9876
rect 32872 9300 32906 9876
rect 33890 9300 33924 9876
rect 1766 8532 1800 9108
rect 2784 8532 2818 9108
rect 3802 8532 3836 9108
rect 4820 8532 4854 9108
rect 5838 8532 5872 9108
rect 6856 8532 6890 9108
rect 7874 8532 7908 9108
rect 8892 8532 8926 9108
rect 9910 8532 9944 9108
rect 10928 8532 10962 9108
rect 1766 7714 1800 8290
rect 2784 7714 2818 8290
rect 3802 7714 3836 8290
rect 4820 7714 4854 8290
rect 5838 7714 5872 8290
rect 6856 7714 6890 8290
rect 7874 7714 7908 8290
rect 8892 7714 8926 8290
rect 9910 7714 9944 8290
rect 10928 7714 10962 8290
rect 13530 8068 13564 8644
rect 14548 8068 14582 8644
rect 15566 8068 15600 8644
rect 16584 8068 16618 8644
rect 17602 8068 17636 8644
rect 18620 8068 18654 8644
rect 19638 8068 19672 8644
rect 20656 8068 20690 8644
rect 21674 8068 21708 8644
rect 22692 8068 22726 8644
rect 23710 8068 23744 8644
rect 24728 8068 24762 8644
rect 25746 8068 25780 8644
rect 26764 8068 26798 8644
rect 27782 8068 27816 8644
rect 28800 8068 28834 8644
rect 29818 8068 29852 8644
rect 30836 8068 30870 8644
rect 31854 8068 31888 8644
rect 32872 8068 32906 8644
rect 33890 8068 33924 8644
rect 8626 6730 8660 6906
rect 8844 6730 8878 6906
rect 9062 6730 9096 6906
rect 9280 6730 9314 6906
rect 9498 6730 9532 6906
rect 9716 6730 9750 6906
rect 9934 6730 9968 6906
rect 10152 6730 10186 6906
rect 10370 6730 10404 6906
rect 10588 6730 10622 6906
rect 10806 6730 10840 6906
rect 13530 6834 13564 7410
rect 14548 6834 14582 7410
rect 15566 6834 15600 7410
rect 16584 6834 16618 7410
rect 17602 6834 17636 7410
rect 18620 6834 18654 7410
rect 19638 6834 19672 7410
rect 20656 6834 20690 7410
rect 21674 6834 21708 7410
rect 22692 6834 22726 7410
rect 23710 6834 23744 7410
rect 24728 6834 24762 7410
rect 25746 6834 25780 7410
rect 26764 6834 26798 7410
rect 27782 6834 27816 7410
rect 28800 6834 28834 7410
rect 29818 6834 29852 7410
rect 30836 6834 30870 7410
rect 31854 6834 31888 7410
rect 32872 6834 32906 7410
rect 33890 6834 33924 7410
rect 8626 5898 8660 6074
rect 8844 5898 8878 6074
rect 9062 5898 9096 6074
rect 9280 5898 9314 6074
rect 9498 5898 9532 6074
rect 9716 5898 9750 6074
rect 9934 5898 9968 6074
rect 10152 5898 10186 6074
rect 10370 5898 10404 6074
rect 10588 5898 10622 6074
rect 10806 5898 10840 6074
rect 13530 5600 13564 6176
rect 14548 5600 14582 6176
rect 15566 5600 15600 6176
rect 16584 5600 16618 6176
rect 17602 5600 17636 6176
rect 18620 5600 18654 6176
rect 19638 5600 19672 6176
rect 20656 5600 20690 6176
rect 21674 5600 21708 6176
rect 22692 5600 22726 6176
rect 23710 5600 23744 6176
rect 24728 5600 24762 6176
rect 25746 5600 25780 6176
rect 26764 5600 26798 6176
rect 27782 5600 27816 6176
rect 28800 5600 28834 6176
rect 29818 5600 29852 6176
rect 30836 5600 30870 6176
rect 31854 5600 31888 6176
rect 32872 5600 32906 6176
rect 33890 5600 33924 6176
rect 1545 4171 1579 4747
rect 2563 4171 2597 4747
rect 3581 4171 3615 4747
rect 4599 4171 4633 4747
rect 5617 4171 5651 4747
rect 6635 4171 6669 4747
rect 7653 4171 7687 4747
rect 8540 4172 8574 4748
rect 8838 4172 8872 4748
rect 9136 4172 9170 4748
rect 9434 4172 9468 4748
rect 9732 4172 9766 4748
rect 10030 4172 10064 4748
rect 10328 4172 10362 4748
rect 10626 4172 10660 4748
rect 10924 4172 10958 4748
rect 11222 4172 11256 4748
rect 11520 4172 11554 4748
rect 11818 4172 11852 4748
rect 13530 4368 13564 4944
rect 14548 4368 14582 4944
rect 15566 4368 15600 4944
rect 16584 4368 16618 4944
rect 17602 4368 17636 4944
rect 18620 4368 18654 4944
rect 19638 4368 19672 4944
rect 20656 4368 20690 4944
rect 21674 4368 21708 4944
rect 22692 4368 22726 4944
rect 23710 4368 23744 4944
rect 24728 4368 24762 4944
rect 25746 4368 25780 4944
rect 26764 4368 26798 4944
rect 27782 4368 27816 4944
rect 28800 4368 28834 4944
rect 29818 4368 29852 4944
rect 30836 4368 30870 4944
rect 31854 4368 31888 4944
rect 32872 4368 32906 4944
rect 33890 4368 33924 4944
rect 1544 3058 1578 3634
rect 2562 3058 2596 3634
rect 3580 3058 3614 3634
rect 4598 3058 4632 3634
rect 5616 3058 5650 3634
rect 6634 3058 6668 3634
rect 7652 3058 7686 3634
rect 8540 3060 8574 3636
rect 8838 3060 8872 3636
rect 9136 3060 9170 3636
rect 9434 3060 9468 3636
rect 9732 3060 9766 3636
rect 10030 3060 10064 3636
rect 10328 3060 10362 3636
rect 10626 3060 10660 3636
rect 10924 3060 10958 3636
rect 11222 3060 11256 3636
rect 11520 3060 11554 3636
rect 11818 3060 11852 3636
rect 13530 3134 13564 3710
rect 14548 3134 14582 3710
rect 15566 3134 15600 3710
rect 16584 3134 16618 3710
rect 17602 3134 17636 3710
rect 18620 3134 18654 3710
rect 19638 3134 19672 3710
rect 20656 3134 20690 3710
rect 21674 3134 21708 3710
rect 22692 3134 22726 3710
rect 23710 3134 23744 3710
rect 24728 3134 24762 3710
rect 25746 3134 25780 3710
rect 26764 3134 26798 3710
rect 27782 3134 27816 3710
rect 28800 3134 28834 3710
rect 29818 3134 29852 3710
rect 30836 3134 30870 3710
rect 31854 3134 31888 3710
rect 32872 3134 32906 3710
rect 33890 3134 33924 3710
rect 1545 1947 1579 2523
rect 2563 1947 2597 2523
rect 3581 1947 3615 2523
rect 4599 1947 4633 2523
rect 5617 1947 5651 2523
rect 6635 1947 6669 2523
rect 7653 1947 7687 2523
rect 8538 1948 8572 2524
rect 8836 1948 8870 2524
rect 9134 1948 9168 2524
rect 9432 1948 9466 2524
rect 9730 1948 9764 2524
rect 10028 1948 10062 2524
rect 10326 1948 10360 2524
rect 10624 1948 10658 2524
rect 10922 1948 10956 2524
rect 11220 1948 11254 2524
rect 11518 1948 11552 2524
rect 11816 1948 11850 2524
rect 13530 1900 13564 2476
rect 14548 1900 14582 2476
rect 15566 1900 15600 2476
rect 16584 1900 16618 2476
rect 17602 1900 17636 2476
rect 18620 1900 18654 2476
rect 19638 1900 19672 2476
rect 20656 1900 20690 2476
rect 21674 1900 21708 2476
rect 22692 1900 22726 2476
rect 23710 1900 23744 2476
rect 24728 1900 24762 2476
rect 25746 1900 25780 2476
rect 26764 1900 26798 2476
rect 27782 1900 27816 2476
rect 28800 1900 28834 2476
rect 29818 1900 29852 2476
rect 30836 1900 30870 2476
rect 31854 1900 31888 2476
rect 32872 1900 32906 2476
rect 33890 1900 33924 2476
rect 1544 834 1578 1410
rect 2562 834 2596 1410
rect 3580 834 3614 1410
rect 4598 834 4632 1410
rect 5616 834 5650 1410
rect 6634 834 6668 1410
rect 7652 834 7686 1410
rect 8538 838 8572 1414
rect 8836 838 8870 1414
rect 9134 838 9168 1414
rect 9432 838 9466 1414
rect 9730 838 9764 1414
rect 10028 838 10062 1414
rect 10326 838 10360 1414
rect 10624 838 10658 1414
rect 10922 838 10956 1414
rect 11220 838 11254 1414
rect 11518 838 11552 1414
rect 11816 838 11850 1414
rect 13530 668 13564 1244
rect 14548 668 14582 1244
rect 15566 668 15600 1244
rect 16584 668 16618 1244
rect 17602 668 17636 1244
rect 18620 668 18654 1244
rect 19638 668 19672 1244
rect 20656 668 20690 1244
rect 21674 668 21708 1244
rect 22692 668 22726 1244
rect 23710 668 23744 1244
rect 24728 668 24762 1244
rect 25746 668 25780 1244
rect 26764 668 26798 1244
rect 27782 668 27816 1244
rect 28800 668 28834 1244
rect 29818 668 29852 1244
rect 30836 668 30870 1244
rect 31854 668 31888 1244
rect 32872 668 32906 1244
rect 33890 668 33924 1244
rect 50656 7515 50690 7549
rect 50656 7447 50690 7481
rect 50740 7515 50774 7549
rect 50740 7447 50774 7481
rect 48804 7152 48838 7328
rect 49062 7152 49096 7328
rect 49320 7152 49354 7328
rect 49578 7152 49612 7328
rect 49836 7152 49870 7328
rect 50094 7152 50128 7328
rect 50352 7152 50386 7328
rect 50656 5551 50690 5585
rect 50656 5483 50690 5517
rect 50740 5551 50774 5585
rect 50740 5483 50774 5517
rect 48804 5188 48838 5364
rect 49062 5188 49096 5364
rect 49320 5188 49354 5364
rect 49578 5188 49612 5364
rect 49836 5188 49870 5364
rect 50094 5188 50128 5364
rect 50352 5188 50386 5364
rect 50656 3551 50690 3585
rect 50656 3483 50690 3517
rect 50740 3551 50774 3585
rect 50740 3483 50774 3517
rect 48804 3188 48838 3364
rect 49062 3188 49096 3364
rect 49320 3188 49354 3364
rect 49578 3188 49612 3364
rect 49836 3188 49870 3364
rect 50094 3188 50128 3364
rect 50352 3188 50386 3364
rect 50656 1461 50690 1495
rect 50656 1393 50690 1427
rect 50740 1461 50774 1495
rect 50740 1393 50774 1427
rect 48804 1098 48838 1274
rect 49062 1098 49096 1274
rect 49320 1098 49354 1274
rect 49578 1098 49612 1274
rect 49836 1098 49870 1274
rect 50094 1098 50128 1274
rect 50352 1098 50386 1274
rect 67532 14234 67566 14810
rect 68550 14234 68584 14810
rect 69568 14234 69602 14810
rect 70586 14234 70620 14810
rect 71604 14234 71638 14810
rect 72622 14234 72656 14810
rect 73640 14234 73674 14810
rect 74658 14234 74692 14810
rect 75676 14234 75710 14810
rect 76694 14234 76728 14810
rect 77712 14234 77746 14810
rect 78730 14234 78764 14810
rect 79748 14234 79782 14810
rect 80766 14234 80800 14810
rect 81784 14234 81818 14810
rect 82802 14234 82836 14810
rect 83820 14234 83854 14810
rect 84838 14234 84872 14810
rect 85856 14234 85890 14810
rect 86874 14234 86908 14810
rect 87892 14234 87926 14810
rect 55766 13440 55800 14016
rect 56784 13440 56818 14016
rect 57802 13440 57836 14016
rect 58820 13440 58854 14016
rect 59838 13440 59872 14016
rect 60856 13440 60890 14016
rect 61874 13440 61908 14016
rect 62892 13440 62926 14016
rect 63910 13440 63944 14016
rect 64928 13440 64962 14016
rect 55766 12622 55800 13198
rect 56784 12622 56818 13198
rect 57802 12622 57836 13198
rect 58820 12622 58854 13198
rect 59838 12622 59872 13198
rect 60856 12622 60890 13198
rect 61874 12622 61908 13198
rect 62892 12622 62926 13198
rect 63910 12622 63944 13198
rect 64928 12622 64962 13198
rect 67532 13000 67566 13576
rect 68550 13000 68584 13576
rect 69568 13000 69602 13576
rect 70586 13000 70620 13576
rect 71604 13000 71638 13576
rect 72622 13000 72656 13576
rect 73640 13000 73674 13576
rect 74658 13000 74692 13576
rect 75676 13000 75710 13576
rect 76694 13000 76728 13576
rect 77712 13000 77746 13576
rect 78730 13000 78764 13576
rect 79748 13000 79782 13576
rect 80766 13000 80800 13576
rect 81784 13000 81818 13576
rect 82802 13000 82836 13576
rect 83820 13000 83854 13576
rect 84838 13000 84872 13576
rect 85856 13000 85890 13576
rect 86874 13000 86908 13576
rect 87892 13000 87926 13576
rect 55766 11804 55800 12380
rect 56784 11804 56818 12380
rect 57802 11804 57836 12380
rect 58820 11804 58854 12380
rect 59838 11804 59872 12380
rect 60856 11804 60890 12380
rect 61874 11804 61908 12380
rect 62892 11804 62926 12380
rect 63910 11804 63944 12380
rect 64928 11804 64962 12380
rect 67532 11768 67566 12344
rect 68550 11768 68584 12344
rect 69568 11768 69602 12344
rect 70586 11768 70620 12344
rect 71604 11768 71638 12344
rect 72622 11768 72656 12344
rect 73640 11768 73674 12344
rect 74658 11768 74692 12344
rect 75676 11768 75710 12344
rect 76694 11768 76728 12344
rect 77712 11768 77746 12344
rect 78730 11768 78764 12344
rect 79748 11768 79782 12344
rect 80766 11768 80800 12344
rect 81784 11768 81818 12344
rect 82802 11768 82836 12344
rect 83820 11768 83854 12344
rect 84838 11768 84872 12344
rect 85856 11768 85890 12344
rect 86874 11768 86908 12344
rect 87892 11768 87926 12344
rect 55766 10986 55800 11562
rect 56784 10986 56818 11562
rect 57802 10986 57836 11562
rect 58820 10986 58854 11562
rect 59838 10986 59872 11562
rect 60856 10986 60890 11562
rect 61874 10986 61908 11562
rect 62892 10986 62926 11562
rect 63910 10986 63944 11562
rect 64928 10986 64962 11562
rect 55766 10168 55800 10744
rect 56784 10168 56818 10744
rect 57802 10168 57836 10744
rect 58820 10168 58854 10744
rect 59838 10168 59872 10744
rect 60856 10168 60890 10744
rect 61874 10168 61908 10744
rect 62892 10168 62926 10744
rect 63910 10168 63944 10744
rect 64928 10168 64962 10744
rect 67530 10534 67564 11110
rect 68548 10534 68582 11110
rect 69566 10534 69600 11110
rect 70584 10534 70618 11110
rect 71602 10534 71636 11110
rect 72620 10534 72654 11110
rect 73638 10534 73672 11110
rect 74656 10534 74690 11110
rect 75674 10534 75708 11110
rect 76692 10534 76726 11110
rect 77710 10534 77744 11110
rect 78728 10534 78762 11110
rect 79746 10534 79780 11110
rect 80764 10534 80798 11110
rect 81782 10534 81816 11110
rect 82800 10534 82834 11110
rect 83818 10534 83852 11110
rect 84836 10534 84870 11110
rect 85854 10534 85888 11110
rect 86872 10534 86906 11110
rect 87890 10534 87924 11110
rect 55766 9350 55800 9926
rect 56784 9350 56818 9926
rect 57802 9350 57836 9926
rect 58820 9350 58854 9926
rect 59838 9350 59872 9926
rect 60856 9350 60890 9926
rect 61874 9350 61908 9926
rect 62892 9350 62926 9926
rect 63910 9350 63944 9926
rect 64928 9350 64962 9926
rect 67530 9300 67564 9876
rect 68548 9300 68582 9876
rect 69566 9300 69600 9876
rect 70584 9300 70618 9876
rect 71602 9300 71636 9876
rect 72620 9300 72654 9876
rect 73638 9300 73672 9876
rect 74656 9300 74690 9876
rect 75674 9300 75708 9876
rect 76692 9300 76726 9876
rect 77710 9300 77744 9876
rect 78728 9300 78762 9876
rect 79746 9300 79780 9876
rect 80764 9300 80798 9876
rect 81782 9300 81816 9876
rect 82800 9300 82834 9876
rect 83818 9300 83852 9876
rect 84836 9300 84870 9876
rect 85854 9300 85888 9876
rect 86872 9300 86906 9876
rect 87890 9300 87924 9876
rect 55766 8532 55800 9108
rect 56784 8532 56818 9108
rect 57802 8532 57836 9108
rect 58820 8532 58854 9108
rect 59838 8532 59872 9108
rect 60856 8532 60890 9108
rect 61874 8532 61908 9108
rect 62892 8532 62926 9108
rect 63910 8532 63944 9108
rect 64928 8532 64962 9108
rect 55766 7714 55800 8290
rect 56784 7714 56818 8290
rect 57802 7714 57836 8290
rect 58820 7714 58854 8290
rect 59838 7714 59872 8290
rect 60856 7714 60890 8290
rect 61874 7714 61908 8290
rect 62892 7714 62926 8290
rect 63910 7714 63944 8290
rect 64928 7714 64962 8290
rect 67530 8068 67564 8644
rect 68548 8068 68582 8644
rect 69566 8068 69600 8644
rect 70584 8068 70618 8644
rect 71602 8068 71636 8644
rect 72620 8068 72654 8644
rect 73638 8068 73672 8644
rect 74656 8068 74690 8644
rect 75674 8068 75708 8644
rect 76692 8068 76726 8644
rect 77710 8068 77744 8644
rect 78728 8068 78762 8644
rect 79746 8068 79780 8644
rect 80764 8068 80798 8644
rect 81782 8068 81816 8644
rect 82800 8068 82834 8644
rect 83818 8068 83852 8644
rect 84836 8068 84870 8644
rect 85854 8068 85888 8644
rect 86872 8068 86906 8644
rect 87890 8068 87924 8644
rect 62626 6730 62660 6906
rect 62844 6730 62878 6906
rect 63062 6730 63096 6906
rect 63280 6730 63314 6906
rect 63498 6730 63532 6906
rect 63716 6730 63750 6906
rect 63934 6730 63968 6906
rect 64152 6730 64186 6906
rect 64370 6730 64404 6906
rect 64588 6730 64622 6906
rect 64806 6730 64840 6906
rect 67530 6834 67564 7410
rect 68548 6834 68582 7410
rect 69566 6834 69600 7410
rect 70584 6834 70618 7410
rect 71602 6834 71636 7410
rect 72620 6834 72654 7410
rect 73638 6834 73672 7410
rect 74656 6834 74690 7410
rect 75674 6834 75708 7410
rect 76692 6834 76726 7410
rect 77710 6834 77744 7410
rect 78728 6834 78762 7410
rect 79746 6834 79780 7410
rect 80764 6834 80798 7410
rect 81782 6834 81816 7410
rect 82800 6834 82834 7410
rect 83818 6834 83852 7410
rect 84836 6834 84870 7410
rect 85854 6834 85888 7410
rect 86872 6834 86906 7410
rect 87890 6834 87924 7410
rect 62626 5898 62660 6074
rect 62844 5898 62878 6074
rect 63062 5898 63096 6074
rect 63280 5898 63314 6074
rect 63498 5898 63532 6074
rect 63716 5898 63750 6074
rect 63934 5898 63968 6074
rect 64152 5898 64186 6074
rect 64370 5898 64404 6074
rect 64588 5898 64622 6074
rect 64806 5898 64840 6074
rect 67530 5600 67564 6176
rect 68548 5600 68582 6176
rect 69566 5600 69600 6176
rect 70584 5600 70618 6176
rect 71602 5600 71636 6176
rect 72620 5600 72654 6176
rect 73638 5600 73672 6176
rect 74656 5600 74690 6176
rect 75674 5600 75708 6176
rect 76692 5600 76726 6176
rect 77710 5600 77744 6176
rect 78728 5600 78762 6176
rect 79746 5600 79780 6176
rect 80764 5600 80798 6176
rect 81782 5600 81816 6176
rect 82800 5600 82834 6176
rect 83818 5600 83852 6176
rect 84836 5600 84870 6176
rect 85854 5600 85888 6176
rect 86872 5600 86906 6176
rect 87890 5600 87924 6176
rect 55545 4171 55579 4747
rect 56563 4171 56597 4747
rect 57581 4171 57615 4747
rect 58599 4171 58633 4747
rect 59617 4171 59651 4747
rect 60635 4171 60669 4747
rect 61653 4171 61687 4747
rect 62540 4172 62574 4748
rect 62838 4172 62872 4748
rect 63136 4172 63170 4748
rect 63434 4172 63468 4748
rect 63732 4172 63766 4748
rect 64030 4172 64064 4748
rect 64328 4172 64362 4748
rect 64626 4172 64660 4748
rect 64924 4172 64958 4748
rect 65222 4172 65256 4748
rect 65520 4172 65554 4748
rect 65818 4172 65852 4748
rect 67530 4368 67564 4944
rect 68548 4368 68582 4944
rect 69566 4368 69600 4944
rect 70584 4368 70618 4944
rect 71602 4368 71636 4944
rect 72620 4368 72654 4944
rect 73638 4368 73672 4944
rect 74656 4368 74690 4944
rect 75674 4368 75708 4944
rect 76692 4368 76726 4944
rect 77710 4368 77744 4944
rect 78728 4368 78762 4944
rect 79746 4368 79780 4944
rect 80764 4368 80798 4944
rect 81782 4368 81816 4944
rect 82800 4368 82834 4944
rect 83818 4368 83852 4944
rect 84836 4368 84870 4944
rect 85854 4368 85888 4944
rect 86872 4368 86906 4944
rect 87890 4368 87924 4944
rect 55544 3058 55578 3634
rect 56562 3058 56596 3634
rect 57580 3058 57614 3634
rect 58598 3058 58632 3634
rect 59616 3058 59650 3634
rect 60634 3058 60668 3634
rect 61652 3058 61686 3634
rect 62540 3060 62574 3636
rect 62838 3060 62872 3636
rect 63136 3060 63170 3636
rect 63434 3060 63468 3636
rect 63732 3060 63766 3636
rect 64030 3060 64064 3636
rect 64328 3060 64362 3636
rect 64626 3060 64660 3636
rect 64924 3060 64958 3636
rect 65222 3060 65256 3636
rect 65520 3060 65554 3636
rect 65818 3060 65852 3636
rect 67530 3134 67564 3710
rect 68548 3134 68582 3710
rect 69566 3134 69600 3710
rect 70584 3134 70618 3710
rect 71602 3134 71636 3710
rect 72620 3134 72654 3710
rect 73638 3134 73672 3710
rect 74656 3134 74690 3710
rect 75674 3134 75708 3710
rect 76692 3134 76726 3710
rect 77710 3134 77744 3710
rect 78728 3134 78762 3710
rect 79746 3134 79780 3710
rect 80764 3134 80798 3710
rect 81782 3134 81816 3710
rect 82800 3134 82834 3710
rect 83818 3134 83852 3710
rect 84836 3134 84870 3710
rect 85854 3134 85888 3710
rect 86872 3134 86906 3710
rect 87890 3134 87924 3710
rect 55545 1947 55579 2523
rect 56563 1947 56597 2523
rect 57581 1947 57615 2523
rect 58599 1947 58633 2523
rect 59617 1947 59651 2523
rect 60635 1947 60669 2523
rect 61653 1947 61687 2523
rect 62538 1948 62572 2524
rect 62836 1948 62870 2524
rect 63134 1948 63168 2524
rect 63432 1948 63466 2524
rect 63730 1948 63764 2524
rect 64028 1948 64062 2524
rect 64326 1948 64360 2524
rect 64624 1948 64658 2524
rect 64922 1948 64956 2524
rect 65220 1948 65254 2524
rect 65518 1948 65552 2524
rect 65816 1948 65850 2524
rect 67530 1900 67564 2476
rect 68548 1900 68582 2476
rect 69566 1900 69600 2476
rect 70584 1900 70618 2476
rect 71602 1900 71636 2476
rect 72620 1900 72654 2476
rect 73638 1900 73672 2476
rect 74656 1900 74690 2476
rect 75674 1900 75708 2476
rect 76692 1900 76726 2476
rect 77710 1900 77744 2476
rect 78728 1900 78762 2476
rect 79746 1900 79780 2476
rect 80764 1900 80798 2476
rect 81782 1900 81816 2476
rect 82800 1900 82834 2476
rect 83818 1900 83852 2476
rect 84836 1900 84870 2476
rect 85854 1900 85888 2476
rect 86872 1900 86906 2476
rect 87890 1900 87924 2476
rect 55544 834 55578 1410
rect 56562 834 56596 1410
rect 57580 834 57614 1410
rect 58598 834 58632 1410
rect 59616 834 59650 1410
rect 60634 834 60668 1410
rect 61652 834 61686 1410
rect 62538 838 62572 1414
rect 62836 838 62870 1414
rect 63134 838 63168 1414
rect 63432 838 63466 1414
rect 63730 838 63764 1414
rect 64028 838 64062 1414
rect 64326 838 64360 1414
rect 64624 838 64658 1414
rect 64922 838 64956 1414
rect 65220 838 65254 1414
rect 65518 838 65552 1414
rect 65816 838 65850 1414
rect 67530 668 67564 1244
rect 68548 668 68582 1244
rect 69566 668 69600 1244
rect 70584 668 70618 1244
rect 71602 668 71636 1244
rect 72620 668 72654 1244
rect 73638 668 73672 1244
rect 74656 668 74690 1244
rect 75674 668 75708 1244
rect 76692 668 76726 1244
rect 77710 668 77744 1244
rect 78728 668 78762 1244
rect 79746 668 79780 1244
rect 80764 668 80798 1244
rect 81782 668 81816 1244
rect 82800 668 82834 1244
rect 83818 668 83852 1244
rect 84836 668 84870 1244
rect 85854 668 85888 1244
rect 86872 668 86906 1244
rect 87890 668 87924 1244
<< pdiffc >>
rect 17438 26392 17472 26968
rect 18456 26392 18490 26968
rect 19474 26392 19508 26968
rect 20492 26392 20526 26968
rect 21510 26392 21544 26968
rect 22528 26392 22562 26968
rect 23546 26392 23580 26968
rect 24564 26392 24598 26968
rect 25582 26392 25616 26968
rect 26600 26392 26634 26968
rect 27618 26392 27652 26968
rect 28636 26392 28670 26968
rect 29654 26392 29688 26968
rect 30672 26392 30706 26968
rect 31690 26392 31724 26968
rect 32708 26392 32742 26968
rect 33726 26392 33760 26968
rect 17438 25256 17472 25832
rect 18456 25256 18490 25832
rect 19474 25256 19508 25832
rect 20492 25256 20526 25832
rect 21510 25256 21544 25832
rect 22528 25256 22562 25832
rect 23546 25256 23580 25832
rect 24564 25256 24598 25832
rect 25582 25256 25616 25832
rect 26600 25256 26634 25832
rect 27618 25256 27652 25832
rect 28636 25256 28670 25832
rect 29654 25256 29688 25832
rect 30672 25256 30706 25832
rect 31690 25256 31724 25832
rect 32708 25256 32742 25832
rect 33726 25256 33760 25832
rect 17438 24120 17472 24696
rect 18456 24120 18490 24696
rect 19474 24120 19508 24696
rect 20492 24120 20526 24696
rect 21510 24120 21544 24696
rect 22528 24120 22562 24696
rect 23546 24120 23580 24696
rect 24564 24120 24598 24696
rect 25582 24120 25616 24696
rect 26600 24120 26634 24696
rect 27618 24120 27652 24696
rect 28636 24120 28670 24696
rect 29654 24120 29688 24696
rect 30672 24120 30706 24696
rect 31690 24120 31724 24696
rect 32708 24120 32742 24696
rect 33726 24120 33760 24696
rect 18424 22346 18458 22922
rect 19442 22346 19476 22922
rect 20460 22346 20494 22922
rect 21478 22346 21512 22922
rect 22496 22346 22530 22922
rect 23514 22346 23548 22922
rect 24532 22346 24566 22922
rect 25550 22346 25584 22922
rect 26568 22346 26602 22922
rect 27586 22346 27620 22922
rect 28604 22346 28638 22922
rect 29622 22346 29656 22922
rect 30640 22346 30674 22922
rect 31658 22346 31692 22922
rect 32676 22346 32710 22922
rect 33694 22346 33728 22922
rect 14576 21462 14610 21838
rect 14794 21462 14828 21838
rect 15012 21462 15046 21838
rect 15230 21462 15264 21838
rect 15448 21462 15482 21838
rect 15666 21462 15700 21838
rect 15884 21462 15918 21838
rect 16102 21462 16136 21838
rect 16320 21462 16354 21838
rect 16538 21462 16572 21838
rect 16756 21462 16790 21838
rect 18424 21090 18458 21666
rect 19442 21090 19476 21666
rect 20460 21090 20494 21666
rect 21478 21090 21512 21666
rect 22496 21090 22530 21666
rect 23514 21090 23548 21666
rect 24532 21090 24566 21666
rect 25550 21090 25584 21666
rect 26568 21090 26602 21666
rect 27586 21090 27620 21666
rect 28604 21090 28638 21666
rect 29622 21090 29656 21666
rect 30640 21090 30674 21666
rect 31658 21090 31692 21666
rect 32676 21090 32710 21666
rect 33694 21090 33728 21666
rect 14576 20524 14610 20900
rect 14794 20524 14828 20900
rect 15012 20524 15046 20900
rect 15230 20524 15264 20900
rect 15448 20524 15482 20900
rect 15666 20524 15700 20900
rect 15884 20524 15918 20900
rect 16102 20524 16136 20900
rect 16320 20524 16354 20900
rect 16538 20524 16572 20900
rect 16756 20524 16790 20900
rect 14576 19586 14610 19962
rect 14794 19586 14828 19962
rect 15012 19586 15046 19962
rect 15230 19586 15264 19962
rect 15448 19586 15482 19962
rect 15666 19586 15700 19962
rect 15884 19586 15918 19962
rect 16102 19586 16136 19962
rect 16320 19586 16354 19962
rect 16538 19586 16572 19962
rect 16756 19586 16790 19962
rect 18424 19834 18458 20410
rect 19442 19834 19476 20410
rect 20460 19834 20494 20410
rect 21478 19834 21512 20410
rect 22496 19834 22530 20410
rect 23514 19834 23548 20410
rect 24532 19834 24566 20410
rect 25550 19834 25584 20410
rect 26568 19834 26602 20410
rect 27586 19834 27620 20410
rect 28604 19834 28638 20410
rect 29622 19834 29656 20410
rect 30640 19834 30674 20410
rect 31658 19834 31692 20410
rect 32676 19834 32710 20410
rect 33694 19834 33728 20410
rect 14576 18648 14610 19024
rect 14794 18648 14828 19024
rect 15012 18648 15046 19024
rect 15230 18648 15264 19024
rect 15448 18648 15482 19024
rect 15666 18648 15700 19024
rect 15884 18648 15918 19024
rect 16102 18648 16136 19024
rect 16320 18648 16354 19024
rect 16538 18648 16572 19024
rect 16756 18648 16790 19024
rect 18424 18578 18458 19154
rect 19442 18578 19476 19154
rect 20460 18578 20494 19154
rect 21478 18578 21512 19154
rect 22496 18578 22530 19154
rect 23514 18578 23548 19154
rect 24532 18578 24566 19154
rect 25550 18578 25584 19154
rect 26568 18578 26602 19154
rect 27586 18578 27620 19154
rect 28604 18578 28638 19154
rect 29622 18578 29656 19154
rect 30640 18578 30674 19154
rect 31658 18578 31692 19154
rect 32676 18578 32710 19154
rect 33694 18578 33728 19154
rect 47378 24840 47412 25216
rect 47636 24840 47670 25216
rect 47894 24840 47928 25216
rect 48152 24840 48186 25216
rect 48410 24840 48444 25216
rect 48668 24840 48702 25216
rect 48926 24840 48960 25216
rect 49230 24799 49264 24833
rect 49230 24731 49264 24765
rect 49230 24663 49264 24697
rect 49314 24799 49348 24833
rect 49314 24731 49348 24765
rect 49314 24663 49348 24697
rect 47378 22840 47412 23216
rect 47636 22840 47670 23216
rect 47894 22840 47928 23216
rect 48152 22840 48186 23216
rect 48410 22840 48444 23216
rect 48668 22840 48702 23216
rect 48926 22840 48960 23216
rect 49230 22799 49264 22833
rect 49230 22731 49264 22765
rect 49230 22663 49264 22697
rect 49314 22799 49348 22833
rect 49314 22731 49348 22765
rect 49314 22663 49348 22697
rect 71438 26392 71472 26968
rect 72456 26392 72490 26968
rect 73474 26392 73508 26968
rect 74492 26392 74526 26968
rect 75510 26392 75544 26968
rect 76528 26392 76562 26968
rect 77546 26392 77580 26968
rect 78564 26392 78598 26968
rect 79582 26392 79616 26968
rect 80600 26392 80634 26968
rect 81618 26392 81652 26968
rect 82636 26392 82670 26968
rect 83654 26392 83688 26968
rect 84672 26392 84706 26968
rect 85690 26392 85724 26968
rect 86708 26392 86742 26968
rect 87726 26392 87760 26968
rect 71438 25256 71472 25832
rect 72456 25256 72490 25832
rect 73474 25256 73508 25832
rect 74492 25256 74526 25832
rect 75510 25256 75544 25832
rect 76528 25256 76562 25832
rect 77546 25256 77580 25832
rect 78564 25256 78598 25832
rect 79582 25256 79616 25832
rect 80600 25256 80634 25832
rect 81618 25256 81652 25832
rect 82636 25256 82670 25832
rect 83654 25256 83688 25832
rect 84672 25256 84706 25832
rect 85690 25256 85724 25832
rect 86708 25256 86742 25832
rect 87726 25256 87760 25832
rect 71438 24120 71472 24696
rect 72456 24120 72490 24696
rect 73474 24120 73508 24696
rect 74492 24120 74526 24696
rect 75510 24120 75544 24696
rect 76528 24120 76562 24696
rect 77546 24120 77580 24696
rect 78564 24120 78598 24696
rect 79582 24120 79616 24696
rect 80600 24120 80634 24696
rect 81618 24120 81652 24696
rect 82636 24120 82670 24696
rect 83654 24120 83688 24696
rect 84672 24120 84706 24696
rect 85690 24120 85724 24696
rect 86708 24120 86742 24696
rect 87726 24120 87760 24696
rect 72424 22346 72458 22922
rect 73442 22346 73476 22922
rect 74460 22346 74494 22922
rect 75478 22346 75512 22922
rect 76496 22346 76530 22922
rect 77514 22346 77548 22922
rect 78532 22346 78566 22922
rect 79550 22346 79584 22922
rect 80568 22346 80602 22922
rect 81586 22346 81620 22922
rect 82604 22346 82638 22922
rect 83622 22346 83656 22922
rect 84640 22346 84674 22922
rect 85658 22346 85692 22922
rect 86676 22346 86710 22922
rect 87694 22346 87728 22922
rect 68576 21462 68610 21838
rect 68794 21462 68828 21838
rect 69012 21462 69046 21838
rect 69230 21462 69264 21838
rect 69448 21462 69482 21838
rect 69666 21462 69700 21838
rect 69884 21462 69918 21838
rect 70102 21462 70136 21838
rect 70320 21462 70354 21838
rect 70538 21462 70572 21838
rect 70756 21462 70790 21838
rect 72424 21090 72458 21666
rect 73442 21090 73476 21666
rect 74460 21090 74494 21666
rect 75478 21090 75512 21666
rect 76496 21090 76530 21666
rect 77514 21090 77548 21666
rect 78532 21090 78566 21666
rect 79550 21090 79584 21666
rect 80568 21090 80602 21666
rect 81586 21090 81620 21666
rect 82604 21090 82638 21666
rect 83622 21090 83656 21666
rect 84640 21090 84674 21666
rect 85658 21090 85692 21666
rect 86676 21090 86710 21666
rect 87694 21090 87728 21666
rect 68576 20524 68610 20900
rect 68794 20524 68828 20900
rect 69012 20524 69046 20900
rect 69230 20524 69264 20900
rect 69448 20524 69482 20900
rect 69666 20524 69700 20900
rect 69884 20524 69918 20900
rect 70102 20524 70136 20900
rect 70320 20524 70354 20900
rect 70538 20524 70572 20900
rect 70756 20524 70790 20900
rect 68576 19586 68610 19962
rect 68794 19586 68828 19962
rect 69012 19586 69046 19962
rect 69230 19586 69264 19962
rect 69448 19586 69482 19962
rect 69666 19586 69700 19962
rect 69884 19586 69918 19962
rect 70102 19586 70136 19962
rect 70320 19586 70354 19962
rect 70538 19586 70572 19962
rect 70756 19586 70790 19962
rect 72424 19834 72458 20410
rect 73442 19834 73476 20410
rect 74460 19834 74494 20410
rect 75478 19834 75512 20410
rect 76496 19834 76530 20410
rect 77514 19834 77548 20410
rect 78532 19834 78566 20410
rect 79550 19834 79584 20410
rect 80568 19834 80602 20410
rect 81586 19834 81620 20410
rect 82604 19834 82638 20410
rect 83622 19834 83656 20410
rect 84640 19834 84674 20410
rect 85658 19834 85692 20410
rect 86676 19834 86710 20410
rect 87694 19834 87728 20410
rect 68576 18648 68610 19024
rect 68794 18648 68828 19024
rect 69012 18648 69046 19024
rect 69230 18648 69264 19024
rect 69448 18648 69482 19024
rect 69666 18648 69700 19024
rect 69884 18648 69918 19024
rect 70102 18648 70136 19024
rect 70320 18648 70354 19024
rect 70538 18648 70572 19024
rect 70756 18648 70790 19024
rect 72424 18578 72458 19154
rect 73442 18578 73476 19154
rect 74460 18578 74494 19154
rect 75478 18578 75512 19154
rect 76496 18578 76530 19154
rect 77514 18578 77548 19154
rect 78532 18578 78566 19154
rect 79550 18578 79584 19154
rect 80568 18578 80602 19154
rect 81586 18578 81620 19154
rect 82604 18578 82638 19154
rect 83622 18578 83656 19154
rect 84640 18578 84674 19154
rect 85658 18578 85692 19154
rect 86676 18578 86710 19154
rect 87694 18578 87728 19154
rect -12980 15710 -12946 16086
rect -12722 15710 -12688 16086
rect -12464 15710 -12430 16086
rect -12206 15710 -12172 16086
rect -11948 15710 -11914 16086
rect -11690 15710 -11656 16086
rect -11432 15710 -11398 16086
rect -11128 15669 -11094 15703
rect -11128 15601 -11094 15635
rect -11128 15533 -11094 15567
rect -11044 15669 -11010 15703
rect -11044 15601 -11010 15635
rect -11044 15533 -11010 15567
rect -10380 15710 -10346 16086
rect -10122 15710 -10088 16086
rect -9864 15710 -9830 16086
rect -9606 15710 -9572 16086
rect -9348 15710 -9314 16086
rect -9090 15710 -9056 16086
rect -8832 15710 -8798 16086
rect -8528 15669 -8494 15703
rect -8528 15601 -8494 15635
rect -8528 15533 -8494 15567
rect -8444 15669 -8410 15703
rect -8444 15601 -8410 15635
rect -8444 15533 -8410 15567
rect -8028 15669 -7994 15703
rect -8028 15601 -7994 15635
rect -8028 15533 -7994 15567
rect -7944 15669 -7910 15703
rect -7944 15601 -7910 15635
rect -7944 15533 -7910 15567
rect 48804 7876 48838 8252
rect 49062 7876 49096 8252
rect 49320 7876 49354 8252
rect 49578 7876 49612 8252
rect 49836 7876 49870 8252
rect 50094 7876 50128 8252
rect 50352 7876 50386 8252
rect 50656 7835 50690 7869
rect 50656 7767 50690 7801
rect 50656 7699 50690 7733
rect 50740 7835 50774 7869
rect 50740 7767 50774 7801
rect 50740 7699 50774 7733
rect 48804 5912 48838 6288
rect 49062 5912 49096 6288
rect 49320 5912 49354 6288
rect 49578 5912 49612 6288
rect 49836 5912 49870 6288
rect 50094 5912 50128 6288
rect 50352 5912 50386 6288
rect 50656 5871 50690 5905
rect 50656 5803 50690 5837
rect 50656 5735 50690 5769
rect 50740 5871 50774 5905
rect 50740 5803 50774 5837
rect 50740 5735 50774 5769
rect 48804 3912 48838 4288
rect 49062 3912 49096 4288
rect 49320 3912 49354 4288
rect 49578 3912 49612 4288
rect 49836 3912 49870 4288
rect 50094 3912 50128 4288
rect 50352 3912 50386 4288
rect 50656 3871 50690 3905
rect 50656 3803 50690 3837
rect 50656 3735 50690 3769
rect 50740 3871 50774 3905
rect 50740 3803 50774 3837
rect 50740 3735 50774 3769
rect 48804 1822 48838 2198
rect 49062 1822 49096 2198
rect 49320 1822 49354 2198
rect 49578 1822 49612 2198
rect 49836 1822 49870 2198
rect 50094 1822 50128 2198
rect 50352 1822 50386 2198
rect 50656 1781 50690 1815
rect 50656 1713 50690 1747
rect 50656 1645 50690 1679
rect 50740 1781 50774 1815
rect 50740 1713 50774 1747
rect 50740 1645 50774 1679
<< psubdiff >>
rect 47264 24444 47360 24478
rect 48978 24444 49074 24478
rect 47264 24382 47298 24444
rect 49040 24382 49074 24444
rect 47264 23964 47298 24026
rect 49040 23964 49074 24026
rect 47264 23930 47360 23964
rect 48978 23930 49074 23964
rect 47264 22444 47360 22478
rect 48978 22444 49074 22478
rect 47264 22382 47298 22444
rect 49040 22382 49074 22444
rect 47264 21964 47298 22026
rect 49040 21964 49074 22026
rect 47264 21930 47360 21964
rect 48978 21930 49074 21964
rect -13094 15314 -12998 15348
rect -11380 15314 -11284 15348
rect -13094 15252 -13060 15314
rect -11318 15252 -11284 15314
rect -10494 15314 -10398 15348
rect -8780 15314 -8684 15348
rect -13094 14834 -13060 14896
rect -10494 15252 -10460 15314
rect -11318 14834 -11284 14896
rect -13094 14800 -12998 14834
rect -11380 14800 -11284 14834
rect -8718 15252 -8684 15314
rect -10494 14834 -10460 14896
rect -1372 15262 -1210 15362
rect 35710 15262 35872 15362
rect -8718 14834 -8684 14896
rect -10494 14800 -10398 14834
rect -8780 14800 -8684 14834
rect -1372 15200 -1272 15262
rect 35772 15200 35872 15262
rect 2282 14318 2364 14342
rect 2282 14284 2306 14318
rect 2340 14284 2364 14318
rect 2282 14260 2364 14284
rect 3300 14318 3382 14342
rect 3300 14284 3324 14318
rect 3358 14284 3382 14318
rect 3300 14260 3382 14284
rect 4318 14318 4400 14342
rect 4318 14284 4342 14318
rect 4376 14284 4400 14318
rect 4318 14260 4400 14284
rect 5336 14318 5418 14342
rect 5336 14284 5360 14318
rect 5394 14284 5418 14318
rect 5336 14260 5418 14284
rect 6354 14318 6436 14342
rect 6354 14284 6378 14318
rect 6412 14284 6436 14318
rect 6354 14260 6436 14284
rect 7372 14318 7454 14342
rect 7372 14284 7396 14318
rect 7430 14284 7454 14318
rect 7372 14260 7454 14284
rect 8390 14318 8472 14342
rect 8390 14284 8414 14318
rect 8448 14284 8472 14318
rect 8390 14260 8472 14284
rect 9408 14318 9490 14342
rect 9408 14284 9432 14318
rect 9466 14284 9490 14318
rect 9408 14260 9490 14284
rect 10426 14318 10508 14342
rect 10426 14284 10450 14318
rect 10484 14284 10508 14318
rect 10426 14260 10508 14284
rect 14016 13926 14098 13950
rect 14016 13892 14040 13926
rect 14074 13892 14098 13926
rect 14016 13868 14098 13892
rect 15034 13926 15116 13950
rect 15034 13892 15058 13926
rect 15092 13892 15116 13926
rect 15034 13868 15116 13892
rect 16052 13926 16134 13950
rect 16052 13892 16076 13926
rect 16110 13892 16134 13926
rect 16052 13868 16134 13892
rect 17070 13926 17152 13950
rect 17070 13892 17094 13926
rect 17128 13892 17152 13926
rect 17070 13868 17152 13892
rect 18088 13926 18170 13950
rect 18088 13892 18112 13926
rect 18146 13892 18170 13926
rect 18088 13868 18170 13892
rect 19106 13926 19188 13950
rect 19106 13892 19130 13926
rect 19164 13892 19188 13926
rect 19106 13868 19188 13892
rect 20124 13926 20206 13950
rect 20124 13892 20148 13926
rect 20182 13892 20206 13926
rect 20124 13868 20206 13892
rect 21142 13926 21224 13950
rect 21142 13892 21166 13926
rect 21200 13892 21224 13926
rect 21142 13868 21224 13892
rect 22160 13926 22242 13950
rect 22160 13892 22184 13926
rect 22218 13892 22242 13926
rect 22160 13868 22242 13892
rect 23178 13926 23260 13950
rect 23178 13892 23202 13926
rect 23236 13892 23260 13926
rect 23178 13868 23260 13892
rect 24196 13926 24278 13950
rect 24196 13892 24220 13926
rect 24254 13892 24278 13926
rect 24196 13868 24278 13892
rect 25214 13926 25296 13950
rect 25214 13892 25238 13926
rect 25272 13892 25296 13926
rect 25214 13868 25296 13892
rect 26232 13926 26314 13950
rect 26232 13892 26256 13926
rect 26290 13892 26314 13926
rect 26232 13868 26314 13892
rect 27250 13926 27332 13950
rect 27250 13892 27274 13926
rect 27308 13892 27332 13926
rect 27250 13868 27332 13892
rect 28268 13926 28350 13950
rect 28268 13892 28292 13926
rect 28326 13892 28350 13926
rect 28268 13868 28350 13892
rect 29286 13926 29368 13950
rect 29286 13892 29310 13926
rect 29344 13892 29368 13926
rect 29286 13868 29368 13892
rect 30304 13926 30386 13950
rect 30304 13892 30328 13926
rect 30362 13892 30386 13926
rect 30304 13868 30386 13892
rect 31322 13926 31404 13950
rect 31322 13892 31346 13926
rect 31380 13892 31404 13926
rect 31322 13868 31404 13892
rect 32340 13926 32422 13950
rect 32340 13892 32364 13926
rect 32398 13892 32422 13926
rect 32340 13868 32422 13892
rect 33358 13926 33440 13950
rect 33358 13892 33382 13926
rect 33416 13892 33440 13926
rect 33358 13868 33440 13892
rect 1744 13336 1826 13360
rect 1744 13302 1768 13336
rect 1802 13302 1826 13336
rect 1744 13278 1826 13302
rect 2762 13336 2844 13360
rect 2762 13302 2786 13336
rect 2820 13302 2844 13336
rect 2762 13278 2844 13302
rect 3780 13336 3862 13360
rect 3780 13302 3804 13336
rect 3838 13302 3862 13336
rect 3780 13278 3862 13302
rect 4798 13336 4880 13360
rect 4798 13302 4822 13336
rect 4856 13302 4880 13336
rect 4798 13278 4880 13302
rect 5816 13336 5898 13360
rect 5816 13302 5840 13336
rect 5874 13302 5898 13336
rect 5816 13278 5898 13302
rect 6834 13336 6916 13360
rect 6834 13302 6858 13336
rect 6892 13302 6916 13336
rect 6834 13278 6916 13302
rect 7852 13336 7934 13360
rect 7852 13302 7876 13336
rect 7910 13302 7934 13336
rect 7852 13278 7934 13302
rect 8870 13336 8952 13360
rect 8870 13302 8894 13336
rect 8928 13302 8952 13336
rect 8870 13278 8952 13302
rect 9888 13336 9970 13360
rect 9888 13302 9912 13336
rect 9946 13302 9970 13336
rect 9888 13278 9970 13302
rect 10906 13336 10988 13360
rect 10906 13302 10930 13336
rect 10964 13302 10988 13336
rect 10906 13278 10988 13302
rect 14004 12690 14086 12714
rect 14004 12656 14028 12690
rect 14062 12656 14086 12690
rect 14004 12632 14086 12656
rect 15022 12690 15104 12714
rect 15022 12656 15046 12690
rect 15080 12656 15104 12690
rect 15022 12632 15104 12656
rect 16040 12690 16122 12714
rect 16040 12656 16064 12690
rect 16098 12656 16122 12690
rect 16040 12632 16122 12656
rect 17058 12690 17140 12714
rect 17058 12656 17082 12690
rect 17116 12656 17140 12690
rect 17058 12632 17140 12656
rect 18076 12690 18158 12714
rect 18076 12656 18100 12690
rect 18134 12656 18158 12690
rect 18076 12632 18158 12656
rect 19094 12690 19176 12714
rect 19094 12656 19118 12690
rect 19152 12656 19176 12690
rect 19094 12632 19176 12656
rect 20112 12690 20194 12714
rect 20112 12656 20136 12690
rect 20170 12656 20194 12690
rect 20112 12632 20194 12656
rect 21130 12690 21212 12714
rect 21130 12656 21154 12690
rect 21188 12656 21212 12690
rect 21130 12632 21212 12656
rect 22148 12690 22230 12714
rect 22148 12656 22172 12690
rect 22206 12656 22230 12690
rect 22148 12632 22230 12656
rect 23166 12690 23248 12714
rect 23166 12656 23190 12690
rect 23224 12656 23248 12690
rect 23166 12632 23248 12656
rect 24184 12690 24266 12714
rect 24184 12656 24208 12690
rect 24242 12656 24266 12690
rect 24184 12632 24266 12656
rect 25202 12690 25284 12714
rect 25202 12656 25226 12690
rect 25260 12656 25284 12690
rect 25202 12632 25284 12656
rect 26220 12690 26302 12714
rect 26220 12656 26244 12690
rect 26278 12656 26302 12690
rect 26220 12632 26302 12656
rect 27238 12690 27320 12714
rect 27238 12656 27262 12690
rect 27296 12656 27320 12690
rect 27238 12632 27320 12656
rect 28256 12690 28338 12714
rect 28256 12656 28280 12690
rect 28314 12656 28338 12690
rect 28256 12632 28338 12656
rect 29274 12690 29356 12714
rect 29274 12656 29298 12690
rect 29332 12656 29356 12690
rect 29274 12632 29356 12656
rect 30292 12690 30374 12714
rect 30292 12656 30316 12690
rect 30350 12656 30374 12690
rect 30292 12632 30374 12656
rect 31310 12690 31392 12714
rect 31310 12656 31334 12690
rect 31368 12656 31392 12690
rect 31310 12632 31392 12656
rect 32328 12690 32410 12714
rect 32328 12656 32352 12690
rect 32386 12656 32410 12690
rect 32328 12632 32410 12656
rect 33346 12690 33428 12714
rect 33346 12656 33370 12690
rect 33404 12656 33428 12690
rect 33346 12632 33428 12656
rect 1744 12518 1826 12542
rect 1744 12484 1768 12518
rect 1802 12484 1826 12518
rect 1744 12460 1826 12484
rect 2762 12518 2844 12542
rect 2762 12484 2786 12518
rect 2820 12484 2844 12518
rect 2762 12460 2844 12484
rect 3780 12518 3862 12542
rect 3780 12484 3804 12518
rect 3838 12484 3862 12518
rect 3780 12460 3862 12484
rect 4798 12518 4880 12542
rect 4798 12484 4822 12518
rect 4856 12484 4880 12518
rect 4798 12460 4880 12484
rect 5816 12518 5898 12542
rect 5816 12484 5840 12518
rect 5874 12484 5898 12518
rect 5816 12460 5898 12484
rect 6834 12518 6916 12542
rect 6834 12484 6858 12518
rect 6892 12484 6916 12518
rect 6834 12460 6916 12484
rect 7852 12518 7934 12542
rect 7852 12484 7876 12518
rect 7910 12484 7934 12518
rect 7852 12460 7934 12484
rect 8870 12518 8952 12542
rect 8870 12484 8894 12518
rect 8928 12484 8952 12518
rect 8870 12460 8952 12484
rect 9888 12518 9970 12542
rect 9888 12484 9912 12518
rect 9946 12484 9970 12518
rect 9888 12460 9970 12484
rect 10906 12518 10988 12542
rect 10906 12484 10930 12518
rect 10964 12484 10988 12518
rect 10906 12460 10988 12484
rect 1744 11700 1826 11724
rect 1744 11666 1768 11700
rect 1802 11666 1826 11700
rect 1744 11642 1826 11666
rect 2762 11700 2844 11724
rect 2762 11666 2786 11700
rect 2820 11666 2844 11700
rect 2762 11642 2844 11666
rect 3780 11700 3862 11724
rect 3780 11666 3804 11700
rect 3838 11666 3862 11700
rect 3780 11642 3862 11666
rect 4798 11700 4880 11724
rect 4798 11666 4822 11700
rect 4856 11666 4880 11700
rect 4798 11642 4880 11666
rect 5816 11700 5898 11724
rect 5816 11666 5840 11700
rect 5874 11666 5898 11700
rect 5816 11642 5898 11666
rect 6834 11700 6916 11724
rect 6834 11666 6858 11700
rect 6892 11666 6916 11700
rect 6834 11642 6916 11666
rect 7852 11700 7934 11724
rect 7852 11666 7876 11700
rect 7910 11666 7934 11700
rect 7852 11642 7934 11666
rect 8870 11700 8952 11724
rect 8870 11666 8894 11700
rect 8928 11666 8952 11700
rect 8870 11642 8952 11666
rect 9888 11700 9970 11724
rect 9888 11666 9912 11700
rect 9946 11666 9970 11700
rect 9888 11642 9970 11666
rect 10906 11700 10988 11724
rect 10906 11666 10930 11700
rect 10964 11666 10988 11700
rect 10906 11642 10988 11666
rect 14016 11456 14098 11480
rect 14016 11422 14040 11456
rect 14074 11422 14098 11456
rect 14016 11398 14098 11422
rect 15034 11456 15116 11480
rect 15034 11422 15058 11456
rect 15092 11422 15116 11456
rect 15034 11398 15116 11422
rect 16052 11456 16134 11480
rect 16052 11422 16076 11456
rect 16110 11422 16134 11456
rect 16052 11398 16134 11422
rect 17070 11456 17152 11480
rect 17070 11422 17094 11456
rect 17128 11422 17152 11456
rect 17070 11398 17152 11422
rect 18088 11456 18170 11480
rect 18088 11422 18112 11456
rect 18146 11422 18170 11456
rect 18088 11398 18170 11422
rect 19106 11456 19188 11480
rect 19106 11422 19130 11456
rect 19164 11422 19188 11456
rect 19106 11398 19188 11422
rect 20124 11456 20206 11480
rect 20124 11422 20148 11456
rect 20182 11422 20206 11456
rect 20124 11398 20206 11422
rect 21142 11456 21224 11480
rect 21142 11422 21166 11456
rect 21200 11422 21224 11456
rect 21142 11398 21224 11422
rect 22160 11456 22242 11480
rect 22160 11422 22184 11456
rect 22218 11422 22242 11456
rect 22160 11398 22242 11422
rect 23178 11456 23260 11480
rect 23178 11422 23202 11456
rect 23236 11422 23260 11456
rect 23178 11398 23260 11422
rect 24196 11456 24278 11480
rect 24196 11422 24220 11456
rect 24254 11422 24278 11456
rect 24196 11398 24278 11422
rect 25214 11456 25296 11480
rect 25214 11422 25238 11456
rect 25272 11422 25296 11456
rect 25214 11398 25296 11422
rect 26232 11456 26314 11480
rect 26232 11422 26256 11456
rect 26290 11422 26314 11456
rect 26232 11398 26314 11422
rect 27250 11456 27332 11480
rect 27250 11422 27274 11456
rect 27308 11422 27332 11456
rect 27250 11398 27332 11422
rect 28268 11456 28350 11480
rect 28268 11422 28292 11456
rect 28326 11422 28350 11456
rect 28268 11398 28350 11422
rect 29286 11456 29368 11480
rect 29286 11422 29310 11456
rect 29344 11422 29368 11456
rect 29286 11398 29368 11422
rect 30304 11456 30386 11480
rect 30304 11422 30328 11456
rect 30362 11422 30386 11456
rect 30304 11398 30386 11422
rect 31322 11456 31404 11480
rect 31322 11422 31346 11456
rect 31380 11422 31404 11456
rect 31322 11398 31404 11422
rect 32340 11456 32422 11480
rect 32340 11422 32364 11456
rect 32398 11422 32422 11456
rect 32340 11398 32422 11422
rect 33358 11456 33440 11480
rect 33358 11422 33382 11456
rect 33416 11422 33440 11456
rect 33358 11398 33440 11422
rect 1744 10882 1826 10906
rect 1744 10848 1768 10882
rect 1802 10848 1826 10882
rect 1744 10824 1826 10848
rect 2762 10882 2844 10906
rect 2762 10848 2786 10882
rect 2820 10848 2844 10882
rect 2762 10824 2844 10848
rect 3780 10882 3862 10906
rect 3780 10848 3804 10882
rect 3838 10848 3862 10882
rect 3780 10824 3862 10848
rect 4798 10882 4880 10906
rect 4798 10848 4822 10882
rect 4856 10848 4880 10882
rect 4798 10824 4880 10848
rect 5816 10882 5898 10906
rect 5816 10848 5840 10882
rect 5874 10848 5898 10882
rect 5816 10824 5898 10848
rect 6834 10882 6916 10906
rect 6834 10848 6858 10882
rect 6892 10848 6916 10882
rect 6834 10824 6916 10848
rect 7852 10882 7934 10906
rect 7852 10848 7876 10882
rect 7910 10848 7934 10882
rect 7852 10824 7934 10848
rect 8870 10882 8952 10906
rect 8870 10848 8894 10882
rect 8928 10848 8952 10882
rect 8870 10824 8952 10848
rect 9888 10882 9970 10906
rect 9888 10848 9912 10882
rect 9946 10848 9970 10882
rect 9888 10824 9970 10848
rect 10906 10882 10988 10906
rect 10906 10848 10930 10882
rect 10964 10848 10988 10882
rect 10906 10824 10988 10848
rect 14016 10236 14098 10260
rect 14016 10202 14040 10236
rect 14074 10202 14098 10236
rect 14016 10178 14098 10202
rect 15034 10236 15116 10260
rect 15034 10202 15058 10236
rect 15092 10202 15116 10236
rect 15034 10178 15116 10202
rect 16052 10236 16134 10260
rect 16052 10202 16076 10236
rect 16110 10202 16134 10236
rect 16052 10178 16134 10202
rect 17070 10236 17152 10260
rect 17070 10202 17094 10236
rect 17128 10202 17152 10236
rect 17070 10178 17152 10202
rect 18088 10236 18170 10260
rect 18088 10202 18112 10236
rect 18146 10202 18170 10236
rect 18088 10178 18170 10202
rect 19106 10236 19188 10260
rect 19106 10202 19130 10236
rect 19164 10202 19188 10236
rect 19106 10178 19188 10202
rect 20124 10236 20206 10260
rect 20124 10202 20148 10236
rect 20182 10202 20206 10236
rect 20124 10178 20206 10202
rect 21142 10236 21224 10260
rect 21142 10202 21166 10236
rect 21200 10202 21224 10236
rect 21142 10178 21224 10202
rect 22160 10236 22242 10260
rect 22160 10202 22184 10236
rect 22218 10202 22242 10236
rect 22160 10178 22242 10202
rect 23178 10236 23260 10260
rect 23178 10202 23202 10236
rect 23236 10202 23260 10236
rect 23178 10178 23260 10202
rect 24196 10236 24278 10260
rect 24196 10202 24220 10236
rect 24254 10202 24278 10236
rect 24196 10178 24278 10202
rect 25214 10236 25296 10260
rect 25214 10202 25238 10236
rect 25272 10202 25296 10236
rect 25214 10178 25296 10202
rect 26232 10236 26314 10260
rect 26232 10202 26256 10236
rect 26290 10202 26314 10236
rect 26232 10178 26314 10202
rect 27250 10236 27332 10260
rect 27250 10202 27274 10236
rect 27308 10202 27332 10236
rect 27250 10178 27332 10202
rect 28268 10236 28350 10260
rect 28268 10202 28292 10236
rect 28326 10202 28350 10236
rect 28268 10178 28350 10202
rect 29286 10236 29368 10260
rect 29286 10202 29310 10236
rect 29344 10202 29368 10236
rect 29286 10178 29368 10202
rect 30304 10236 30386 10260
rect 30304 10202 30328 10236
rect 30362 10202 30386 10236
rect 30304 10178 30386 10202
rect 31322 10236 31404 10260
rect 31322 10202 31346 10236
rect 31380 10202 31404 10236
rect 31322 10178 31404 10202
rect 32340 10236 32422 10260
rect 32340 10202 32364 10236
rect 32398 10202 32422 10236
rect 32340 10178 32422 10202
rect 33358 10236 33440 10260
rect 33358 10202 33382 10236
rect 33416 10202 33440 10236
rect 33358 10178 33440 10202
rect 1744 10064 1826 10088
rect 1744 10030 1768 10064
rect 1802 10030 1826 10064
rect 1744 10006 1826 10030
rect 2762 10064 2844 10088
rect 2762 10030 2786 10064
rect 2820 10030 2844 10064
rect 2762 10006 2844 10030
rect 3780 10064 3862 10088
rect 3780 10030 3804 10064
rect 3838 10030 3862 10064
rect 3780 10006 3862 10030
rect 4798 10064 4880 10088
rect 4798 10030 4822 10064
rect 4856 10030 4880 10064
rect 4798 10006 4880 10030
rect 5816 10064 5898 10088
rect 5816 10030 5840 10064
rect 5874 10030 5898 10064
rect 5816 10006 5898 10030
rect 6834 10064 6916 10088
rect 6834 10030 6858 10064
rect 6892 10030 6916 10064
rect 6834 10006 6916 10030
rect 7852 10064 7934 10088
rect 7852 10030 7876 10064
rect 7910 10030 7934 10064
rect 7852 10006 7934 10030
rect 8870 10064 8952 10088
rect 8870 10030 8894 10064
rect 8928 10030 8952 10064
rect 8870 10006 8952 10030
rect 9888 10064 9970 10088
rect 9888 10030 9912 10064
rect 9946 10030 9970 10064
rect 9888 10006 9970 10030
rect 10906 10064 10988 10088
rect 10906 10030 10930 10064
rect 10964 10030 10988 10064
rect 10906 10006 10988 10030
rect 1744 9246 1826 9270
rect 1744 9212 1768 9246
rect 1802 9212 1826 9246
rect 1744 9188 1826 9212
rect 2762 9246 2844 9270
rect 2762 9212 2786 9246
rect 2820 9212 2844 9246
rect 2762 9188 2844 9212
rect 3780 9246 3862 9270
rect 3780 9212 3804 9246
rect 3838 9212 3862 9246
rect 3780 9188 3862 9212
rect 4798 9246 4880 9270
rect 4798 9212 4822 9246
rect 4856 9212 4880 9246
rect 4798 9188 4880 9212
rect 5816 9246 5898 9270
rect 5816 9212 5840 9246
rect 5874 9212 5898 9246
rect 5816 9188 5898 9212
rect 6834 9246 6916 9270
rect 6834 9212 6858 9246
rect 6892 9212 6916 9246
rect 6834 9188 6916 9212
rect 7852 9246 7934 9270
rect 7852 9212 7876 9246
rect 7910 9212 7934 9246
rect 7852 9188 7934 9212
rect 8870 9246 8952 9270
rect 8870 9212 8894 9246
rect 8928 9212 8952 9246
rect 8870 9188 8952 9212
rect 9888 9246 9970 9270
rect 9888 9212 9912 9246
rect 9946 9212 9970 9246
rect 9888 9188 9970 9212
rect 10906 9246 10988 9270
rect 10906 9212 10930 9246
rect 10964 9212 10988 9246
rect 10906 9188 10988 9212
rect 14030 8988 14112 9012
rect 14030 8954 14054 8988
rect 14088 8954 14112 8988
rect 14030 8930 14112 8954
rect 15048 8988 15130 9012
rect 15048 8954 15072 8988
rect 15106 8954 15130 8988
rect 15048 8930 15130 8954
rect 16066 8988 16148 9012
rect 16066 8954 16090 8988
rect 16124 8954 16148 8988
rect 16066 8930 16148 8954
rect 17084 8988 17166 9012
rect 17084 8954 17108 8988
rect 17142 8954 17166 8988
rect 17084 8930 17166 8954
rect 18102 8988 18184 9012
rect 18102 8954 18126 8988
rect 18160 8954 18184 8988
rect 18102 8930 18184 8954
rect 19120 8988 19202 9012
rect 19120 8954 19144 8988
rect 19178 8954 19202 8988
rect 19120 8930 19202 8954
rect 20138 8988 20220 9012
rect 20138 8954 20162 8988
rect 20196 8954 20220 8988
rect 20138 8930 20220 8954
rect 21156 8988 21238 9012
rect 21156 8954 21180 8988
rect 21214 8954 21238 8988
rect 21156 8930 21238 8954
rect 22174 8988 22256 9012
rect 22174 8954 22198 8988
rect 22232 8954 22256 8988
rect 22174 8930 22256 8954
rect 23192 8988 23274 9012
rect 23192 8954 23216 8988
rect 23250 8954 23274 8988
rect 23192 8930 23274 8954
rect 24210 8988 24292 9012
rect 24210 8954 24234 8988
rect 24268 8954 24292 8988
rect 24210 8930 24292 8954
rect 25228 8988 25310 9012
rect 25228 8954 25252 8988
rect 25286 8954 25310 8988
rect 25228 8930 25310 8954
rect 26246 8988 26328 9012
rect 26246 8954 26270 8988
rect 26304 8954 26328 8988
rect 26246 8930 26328 8954
rect 27264 8988 27346 9012
rect 27264 8954 27288 8988
rect 27322 8954 27346 8988
rect 27264 8930 27346 8954
rect 28282 8988 28364 9012
rect 28282 8954 28306 8988
rect 28340 8954 28364 8988
rect 28282 8930 28364 8954
rect 29300 8988 29382 9012
rect 29300 8954 29324 8988
rect 29358 8954 29382 8988
rect 29300 8930 29382 8954
rect 30318 8988 30400 9012
rect 30318 8954 30342 8988
rect 30376 8954 30400 8988
rect 30318 8930 30400 8954
rect 31336 8988 31418 9012
rect 31336 8954 31360 8988
rect 31394 8954 31418 8988
rect 31336 8930 31418 8954
rect 32354 8988 32436 9012
rect 32354 8954 32378 8988
rect 32412 8954 32436 8988
rect 32354 8930 32436 8954
rect 33372 8988 33454 9012
rect 33372 8954 33396 8988
rect 33430 8954 33454 8988
rect 33372 8930 33454 8954
rect 1744 8428 1826 8452
rect 1744 8394 1768 8428
rect 1802 8394 1826 8428
rect 1744 8370 1826 8394
rect 2762 8428 2844 8452
rect 2762 8394 2786 8428
rect 2820 8394 2844 8428
rect 2762 8370 2844 8394
rect 3780 8428 3862 8452
rect 3780 8394 3804 8428
rect 3838 8394 3862 8428
rect 3780 8370 3862 8394
rect 4798 8428 4880 8452
rect 4798 8394 4822 8428
rect 4856 8394 4880 8428
rect 4798 8370 4880 8394
rect 5816 8428 5898 8452
rect 5816 8394 5840 8428
rect 5874 8394 5898 8428
rect 5816 8370 5898 8394
rect 6834 8428 6916 8452
rect 6834 8394 6858 8428
rect 6892 8394 6916 8428
rect 6834 8370 6916 8394
rect 7852 8428 7934 8452
rect 7852 8394 7876 8428
rect 7910 8394 7934 8428
rect 7852 8370 7934 8394
rect 8870 8428 8952 8452
rect 8870 8394 8894 8428
rect 8928 8394 8952 8428
rect 8870 8370 8952 8394
rect 9888 8428 9970 8452
rect 9888 8394 9912 8428
rect 9946 8394 9970 8428
rect 9888 8370 9970 8394
rect 10906 8428 10988 8452
rect 10906 8394 10930 8428
rect 10964 8394 10988 8428
rect 10906 8370 10988 8394
rect 14016 7766 14098 7790
rect 14016 7732 14040 7766
rect 14074 7732 14098 7766
rect 14016 7708 14098 7732
rect 15034 7766 15116 7790
rect 15034 7732 15058 7766
rect 15092 7732 15116 7766
rect 15034 7708 15116 7732
rect 16052 7766 16134 7790
rect 16052 7732 16076 7766
rect 16110 7732 16134 7766
rect 16052 7708 16134 7732
rect 17070 7766 17152 7790
rect 17070 7732 17094 7766
rect 17128 7732 17152 7766
rect 17070 7708 17152 7732
rect 18088 7766 18170 7790
rect 18088 7732 18112 7766
rect 18146 7732 18170 7766
rect 18088 7708 18170 7732
rect 19106 7766 19188 7790
rect 19106 7732 19130 7766
rect 19164 7732 19188 7766
rect 19106 7708 19188 7732
rect 20124 7766 20206 7790
rect 20124 7732 20148 7766
rect 20182 7732 20206 7766
rect 20124 7708 20206 7732
rect 21142 7766 21224 7790
rect 21142 7732 21166 7766
rect 21200 7732 21224 7766
rect 21142 7708 21224 7732
rect 22160 7766 22242 7790
rect 22160 7732 22184 7766
rect 22218 7732 22242 7766
rect 22160 7708 22242 7732
rect 23178 7766 23260 7790
rect 23178 7732 23202 7766
rect 23236 7732 23260 7766
rect 23178 7708 23260 7732
rect 24196 7766 24278 7790
rect 24196 7732 24220 7766
rect 24254 7732 24278 7766
rect 24196 7708 24278 7732
rect 25214 7766 25296 7790
rect 25214 7732 25238 7766
rect 25272 7732 25296 7766
rect 25214 7708 25296 7732
rect 26232 7766 26314 7790
rect 26232 7732 26256 7766
rect 26290 7732 26314 7766
rect 26232 7708 26314 7732
rect 27250 7766 27332 7790
rect 27250 7732 27274 7766
rect 27308 7732 27332 7766
rect 27250 7708 27332 7732
rect 28268 7766 28350 7790
rect 28268 7732 28292 7766
rect 28326 7732 28350 7766
rect 28268 7708 28350 7732
rect 29286 7766 29368 7790
rect 29286 7732 29310 7766
rect 29344 7732 29368 7766
rect 29286 7708 29368 7732
rect 30304 7766 30386 7790
rect 30304 7732 30328 7766
rect 30362 7732 30386 7766
rect 30304 7708 30386 7732
rect 31322 7766 31404 7790
rect 31322 7732 31346 7766
rect 31380 7732 31404 7766
rect 31322 7708 31404 7732
rect 32340 7766 32422 7790
rect 32340 7732 32364 7766
rect 32398 7732 32422 7766
rect 32340 7708 32422 7732
rect 33358 7766 33440 7790
rect 33358 7732 33382 7766
rect 33416 7732 33440 7766
rect 33358 7708 33440 7732
rect 2254 7386 2336 7410
rect 2254 7352 2278 7386
rect 2312 7352 2336 7386
rect 2254 7328 2336 7352
rect 3272 7386 3354 7410
rect 3272 7352 3296 7386
rect 3330 7352 3354 7386
rect 3272 7328 3354 7352
rect 4290 7386 4372 7410
rect 4290 7352 4314 7386
rect 4348 7352 4372 7386
rect 4290 7328 4372 7352
rect 5308 7386 5390 7410
rect 5308 7352 5332 7386
rect 5366 7352 5390 7386
rect 5308 7328 5390 7352
rect 6326 7386 6408 7410
rect 6326 7352 6350 7386
rect 6384 7352 6408 7386
rect 6326 7328 6408 7352
rect 7344 7386 7426 7410
rect 7344 7352 7368 7386
rect 7402 7352 7426 7386
rect 7344 7328 7426 7352
rect 8362 7386 8444 7410
rect 8362 7352 8386 7386
rect 8420 7352 8444 7386
rect 8362 7328 8444 7352
rect 9380 7386 9462 7410
rect 9380 7352 9404 7386
rect 9438 7352 9462 7386
rect 9380 7328 9462 7352
rect 10398 7386 10480 7410
rect 10398 7352 10422 7386
rect 10456 7352 10480 7386
rect 10398 7328 10480 7352
rect 14016 6518 14098 6542
rect 14016 6484 14040 6518
rect 14074 6484 14098 6518
rect 14016 6460 14098 6484
rect 15034 6518 15116 6542
rect 15034 6484 15058 6518
rect 15092 6484 15116 6518
rect 15034 6460 15116 6484
rect 16052 6518 16134 6542
rect 16052 6484 16076 6518
rect 16110 6484 16134 6518
rect 16052 6460 16134 6484
rect 17070 6518 17152 6542
rect 17070 6484 17094 6518
rect 17128 6484 17152 6518
rect 17070 6460 17152 6484
rect 18088 6518 18170 6542
rect 18088 6484 18112 6518
rect 18146 6484 18170 6518
rect 18088 6460 18170 6484
rect 19106 6518 19188 6542
rect 19106 6484 19130 6518
rect 19164 6484 19188 6518
rect 19106 6460 19188 6484
rect 20124 6518 20206 6542
rect 20124 6484 20148 6518
rect 20182 6484 20206 6518
rect 20124 6460 20206 6484
rect 21142 6518 21224 6542
rect 21142 6484 21166 6518
rect 21200 6484 21224 6518
rect 21142 6460 21224 6484
rect 22160 6518 22242 6542
rect 22160 6484 22184 6518
rect 22218 6484 22242 6518
rect 22160 6460 22242 6484
rect 23178 6518 23260 6542
rect 23178 6484 23202 6518
rect 23236 6484 23260 6518
rect 23178 6460 23260 6484
rect 24196 6518 24278 6542
rect 24196 6484 24220 6518
rect 24254 6484 24278 6518
rect 24196 6460 24278 6484
rect 25214 6518 25296 6542
rect 25214 6484 25238 6518
rect 25272 6484 25296 6518
rect 25214 6460 25296 6484
rect 26232 6518 26314 6542
rect 26232 6484 26256 6518
rect 26290 6484 26314 6518
rect 26232 6460 26314 6484
rect 27250 6518 27332 6542
rect 27250 6484 27274 6518
rect 27308 6484 27332 6518
rect 27250 6460 27332 6484
rect 28268 6518 28350 6542
rect 28268 6484 28292 6518
rect 28326 6484 28350 6518
rect 28268 6460 28350 6484
rect 29286 6518 29368 6542
rect 29286 6484 29310 6518
rect 29344 6484 29368 6518
rect 29286 6460 29368 6484
rect 30304 6518 30386 6542
rect 30304 6484 30328 6518
rect 30362 6484 30386 6518
rect 30304 6460 30386 6484
rect 31322 6518 31404 6542
rect 31322 6484 31346 6518
rect 31380 6484 31404 6518
rect 31322 6460 31404 6484
rect 32340 6518 32422 6542
rect 32340 6484 32364 6518
rect 32398 6484 32422 6518
rect 32340 6460 32422 6484
rect 33358 6518 33440 6542
rect 33358 6484 33382 6518
rect 33416 6484 33440 6518
rect 33358 6460 33440 6484
rect 8332 6410 8414 6434
rect 8332 6376 8356 6410
rect 8390 6376 8414 6410
rect 8332 6352 8414 6376
rect 9350 6410 9432 6434
rect 9350 6376 9374 6410
rect 9408 6376 9432 6410
rect 9350 6352 9432 6376
rect 10368 6410 10450 6434
rect 10368 6376 10392 6410
rect 10426 6376 10450 6410
rect 10368 6352 10450 6376
rect 11386 6410 11468 6434
rect 11386 6376 11410 6410
rect 11444 6376 11468 6410
rect 11386 6352 11468 6376
rect 14030 5298 14112 5322
rect 14030 5264 14054 5298
rect 14088 5264 14112 5298
rect 14030 5240 14112 5264
rect 15048 5298 15130 5322
rect 15048 5264 15072 5298
rect 15106 5264 15130 5298
rect 15048 5240 15130 5264
rect 16066 5298 16148 5322
rect 16066 5264 16090 5298
rect 16124 5264 16148 5298
rect 16066 5240 16148 5264
rect 17084 5298 17166 5322
rect 17084 5264 17108 5298
rect 17142 5264 17166 5298
rect 17084 5240 17166 5264
rect 18102 5298 18184 5322
rect 18102 5264 18126 5298
rect 18160 5264 18184 5298
rect 18102 5240 18184 5264
rect 19120 5298 19202 5322
rect 19120 5264 19144 5298
rect 19178 5264 19202 5298
rect 19120 5240 19202 5264
rect 20138 5298 20220 5322
rect 20138 5264 20162 5298
rect 20196 5264 20220 5298
rect 20138 5240 20220 5264
rect 21156 5298 21238 5322
rect 21156 5264 21180 5298
rect 21214 5264 21238 5298
rect 21156 5240 21238 5264
rect 22174 5298 22256 5322
rect 22174 5264 22198 5298
rect 22232 5264 22256 5298
rect 22174 5240 22256 5264
rect 23192 5298 23274 5322
rect 23192 5264 23216 5298
rect 23250 5264 23274 5298
rect 23192 5240 23274 5264
rect 24210 5298 24292 5322
rect 24210 5264 24234 5298
rect 24268 5264 24292 5298
rect 24210 5240 24292 5264
rect 25228 5298 25310 5322
rect 25228 5264 25252 5298
rect 25286 5264 25310 5298
rect 25228 5240 25310 5264
rect 26246 5298 26328 5322
rect 26246 5264 26270 5298
rect 26304 5264 26328 5298
rect 26246 5240 26328 5264
rect 27264 5298 27346 5322
rect 27264 5264 27288 5298
rect 27322 5264 27346 5298
rect 27264 5240 27346 5264
rect 28282 5298 28364 5322
rect 28282 5264 28306 5298
rect 28340 5264 28364 5298
rect 28282 5240 28364 5264
rect 29300 5298 29382 5322
rect 29300 5264 29324 5298
rect 29358 5264 29382 5298
rect 29300 5240 29382 5264
rect 30318 5298 30400 5322
rect 30318 5264 30342 5298
rect 30376 5264 30400 5298
rect 30318 5240 30400 5264
rect 31336 5298 31418 5322
rect 31336 5264 31360 5298
rect 31394 5264 31418 5298
rect 31336 5240 31418 5264
rect 32354 5298 32436 5322
rect 32354 5264 32378 5298
rect 32412 5264 32436 5298
rect 32354 5240 32436 5264
rect 33372 5298 33454 5322
rect 33372 5264 33396 5298
rect 33430 5264 33454 5298
rect 33372 5240 33454 5264
rect 8630 5122 8712 5146
rect 2038 5066 2120 5090
rect 2038 5032 2062 5066
rect 2096 5032 2120 5066
rect 2038 5008 2120 5032
rect 3056 5066 3138 5090
rect 3056 5032 3080 5066
rect 3114 5032 3138 5066
rect 3056 5008 3138 5032
rect 4074 5066 4156 5090
rect 4074 5032 4098 5066
rect 4132 5032 4156 5066
rect 4074 5008 4156 5032
rect 5092 5066 5174 5090
rect 5092 5032 5116 5066
rect 5150 5032 5174 5066
rect 5092 5008 5174 5032
rect 6110 5066 6192 5090
rect 6110 5032 6134 5066
rect 6168 5032 6192 5066
rect 6110 5008 6192 5032
rect 7128 5066 7210 5090
rect 7128 5032 7152 5066
rect 7186 5032 7210 5066
rect 8630 5088 8654 5122
rect 8688 5088 8712 5122
rect 8630 5064 8712 5088
rect 9648 5122 9730 5146
rect 9648 5088 9672 5122
rect 9706 5088 9730 5122
rect 9648 5064 9730 5088
rect 10666 5122 10748 5146
rect 10666 5088 10690 5122
rect 10724 5088 10748 5122
rect 10666 5064 10748 5088
rect 11684 5122 11766 5146
rect 11684 5088 11708 5122
rect 11742 5088 11766 5122
rect 11684 5064 11766 5088
rect 7128 5008 7210 5032
rect 14030 4050 14112 4074
rect 14030 4016 14054 4050
rect 14088 4016 14112 4050
rect 14030 3992 14112 4016
rect 15048 4050 15130 4074
rect 15048 4016 15072 4050
rect 15106 4016 15130 4050
rect 15048 3992 15130 4016
rect 16066 4050 16148 4074
rect 16066 4016 16090 4050
rect 16124 4016 16148 4050
rect 16066 3992 16148 4016
rect 17084 4050 17166 4074
rect 17084 4016 17108 4050
rect 17142 4016 17166 4050
rect 17084 3992 17166 4016
rect 18102 4050 18184 4074
rect 18102 4016 18126 4050
rect 18160 4016 18184 4050
rect 18102 3992 18184 4016
rect 19120 4050 19202 4074
rect 19120 4016 19144 4050
rect 19178 4016 19202 4050
rect 19120 3992 19202 4016
rect 20138 4050 20220 4074
rect 20138 4016 20162 4050
rect 20196 4016 20220 4050
rect 20138 3992 20220 4016
rect 21156 4050 21238 4074
rect 21156 4016 21180 4050
rect 21214 4016 21238 4050
rect 21156 3992 21238 4016
rect 22174 4050 22256 4074
rect 22174 4016 22198 4050
rect 22232 4016 22256 4050
rect 22174 3992 22256 4016
rect 23192 4050 23274 4074
rect 23192 4016 23216 4050
rect 23250 4016 23274 4050
rect 23192 3992 23274 4016
rect 24210 4050 24292 4074
rect 24210 4016 24234 4050
rect 24268 4016 24292 4050
rect 24210 3992 24292 4016
rect 25228 4050 25310 4074
rect 25228 4016 25252 4050
rect 25286 4016 25310 4050
rect 25228 3992 25310 4016
rect 26246 4050 26328 4074
rect 26246 4016 26270 4050
rect 26304 4016 26328 4050
rect 26246 3992 26328 4016
rect 27264 4050 27346 4074
rect 27264 4016 27288 4050
rect 27322 4016 27346 4050
rect 27264 3992 27346 4016
rect 28282 4050 28364 4074
rect 28282 4016 28306 4050
rect 28340 4016 28364 4050
rect 28282 3992 28364 4016
rect 29300 4050 29382 4074
rect 29300 4016 29324 4050
rect 29358 4016 29382 4050
rect 29300 3992 29382 4016
rect 30318 4050 30400 4074
rect 30318 4016 30342 4050
rect 30376 4016 30400 4050
rect 30318 3992 30400 4016
rect 31336 4050 31418 4074
rect 31336 4016 31360 4050
rect 31394 4016 31418 4050
rect 31336 3992 31418 4016
rect 32354 4050 32436 4074
rect 32354 4016 32378 4050
rect 32412 4016 32436 4050
rect 32354 3992 32436 4016
rect 33372 4050 33454 4074
rect 33372 4016 33396 4050
rect 33430 4016 33454 4050
rect 33372 3992 33454 4016
rect 2052 3940 2134 3964
rect 2052 3906 2076 3940
rect 2110 3906 2134 3940
rect 2052 3882 2134 3906
rect 3070 3940 3152 3964
rect 3070 3906 3094 3940
rect 3128 3906 3152 3940
rect 3070 3882 3152 3906
rect 4088 3940 4170 3964
rect 4088 3906 4112 3940
rect 4146 3906 4170 3940
rect 4088 3882 4170 3906
rect 5106 3940 5188 3964
rect 5106 3906 5130 3940
rect 5164 3906 5188 3940
rect 5106 3882 5188 3906
rect 6124 3940 6206 3964
rect 6124 3906 6148 3940
rect 6182 3906 6206 3940
rect 6124 3882 6206 3906
rect 7142 3940 7224 3964
rect 7142 3906 7166 3940
rect 7200 3906 7224 3940
rect 7142 3882 7224 3906
rect 8590 3928 8672 3952
rect 8590 3894 8614 3928
rect 8648 3894 8672 3928
rect 8590 3870 8672 3894
rect 9608 3928 9690 3952
rect 9608 3894 9632 3928
rect 9666 3894 9690 3928
rect 9608 3870 9690 3894
rect 10626 3928 10708 3952
rect 10626 3894 10650 3928
rect 10684 3894 10708 3928
rect 10626 3870 10708 3894
rect 11644 3928 11726 3952
rect 11644 3894 11668 3928
rect 11702 3894 11726 3928
rect 11644 3870 11726 3894
rect 2026 2814 2108 2838
rect 2026 2780 2050 2814
rect 2084 2780 2108 2814
rect 2026 2756 2108 2780
rect 3044 2814 3126 2838
rect 3044 2780 3068 2814
rect 3102 2780 3126 2814
rect 3044 2756 3126 2780
rect 4062 2814 4144 2838
rect 4062 2780 4086 2814
rect 4120 2780 4144 2814
rect 4062 2756 4144 2780
rect 5080 2814 5162 2838
rect 5080 2780 5104 2814
rect 5138 2780 5162 2814
rect 5080 2756 5162 2780
rect 6098 2814 6180 2838
rect 6098 2780 6122 2814
rect 6156 2780 6180 2814
rect 6098 2756 6180 2780
rect 7116 2814 7198 2838
rect 7116 2780 7140 2814
rect 7174 2780 7198 2814
rect 7116 2756 7198 2780
rect 8590 2814 8672 2838
rect 8590 2780 8614 2814
rect 8648 2780 8672 2814
rect 8590 2756 8672 2780
rect 9608 2814 9690 2838
rect 9608 2780 9632 2814
rect 9666 2780 9690 2814
rect 9608 2756 9690 2780
rect 10626 2814 10708 2838
rect 10626 2780 10650 2814
rect 10684 2780 10708 2814
rect 10626 2756 10708 2780
rect 11644 2814 11726 2838
rect 11644 2780 11668 2814
rect 11702 2780 11726 2814
rect 11644 2756 11726 2780
rect 14016 2828 14098 2852
rect 14016 2794 14040 2828
rect 14074 2794 14098 2828
rect 14016 2770 14098 2794
rect 15034 2828 15116 2852
rect 15034 2794 15058 2828
rect 15092 2794 15116 2828
rect 15034 2770 15116 2794
rect 16052 2828 16134 2852
rect 16052 2794 16076 2828
rect 16110 2794 16134 2828
rect 16052 2770 16134 2794
rect 17070 2828 17152 2852
rect 17070 2794 17094 2828
rect 17128 2794 17152 2828
rect 17070 2770 17152 2794
rect 18088 2828 18170 2852
rect 18088 2794 18112 2828
rect 18146 2794 18170 2828
rect 18088 2770 18170 2794
rect 19106 2828 19188 2852
rect 19106 2794 19130 2828
rect 19164 2794 19188 2828
rect 19106 2770 19188 2794
rect 20124 2828 20206 2852
rect 20124 2794 20148 2828
rect 20182 2794 20206 2828
rect 20124 2770 20206 2794
rect 21142 2828 21224 2852
rect 21142 2794 21166 2828
rect 21200 2794 21224 2828
rect 21142 2770 21224 2794
rect 22160 2828 22242 2852
rect 22160 2794 22184 2828
rect 22218 2794 22242 2828
rect 22160 2770 22242 2794
rect 23178 2828 23260 2852
rect 23178 2794 23202 2828
rect 23236 2794 23260 2828
rect 23178 2770 23260 2794
rect 24196 2828 24278 2852
rect 24196 2794 24220 2828
rect 24254 2794 24278 2828
rect 24196 2770 24278 2794
rect 25214 2828 25296 2852
rect 25214 2794 25238 2828
rect 25272 2794 25296 2828
rect 25214 2770 25296 2794
rect 26232 2828 26314 2852
rect 26232 2794 26256 2828
rect 26290 2794 26314 2828
rect 26232 2770 26314 2794
rect 27250 2828 27332 2852
rect 27250 2794 27274 2828
rect 27308 2794 27332 2828
rect 27250 2770 27332 2794
rect 28268 2828 28350 2852
rect 28268 2794 28292 2828
rect 28326 2794 28350 2828
rect 28268 2770 28350 2794
rect 29286 2828 29368 2852
rect 29286 2794 29310 2828
rect 29344 2794 29368 2828
rect 29286 2770 29368 2794
rect 30304 2828 30386 2852
rect 30304 2794 30328 2828
rect 30362 2794 30386 2828
rect 30304 2770 30386 2794
rect 31322 2828 31404 2852
rect 31322 2794 31346 2828
rect 31380 2794 31404 2828
rect 31322 2770 31404 2794
rect 32340 2828 32422 2852
rect 32340 2794 32364 2828
rect 32398 2794 32422 2828
rect 32340 2770 32422 2794
rect 33358 2828 33440 2852
rect 33358 2794 33382 2828
rect 33416 2794 33440 2828
rect 33358 2770 33440 2794
rect 2052 1716 2134 1740
rect 2052 1682 2076 1716
rect 2110 1682 2134 1716
rect 2052 1658 2134 1682
rect 3070 1716 3152 1740
rect 3070 1682 3094 1716
rect 3128 1682 3152 1716
rect 3070 1658 3152 1682
rect 4088 1716 4170 1740
rect 4088 1682 4112 1716
rect 4146 1682 4170 1716
rect 4088 1658 4170 1682
rect 5106 1716 5188 1740
rect 5106 1682 5130 1716
rect 5164 1682 5188 1716
rect 5106 1658 5188 1682
rect 6124 1716 6206 1740
rect 6124 1682 6148 1716
rect 6182 1682 6206 1716
rect 6124 1658 6206 1682
rect 7142 1716 7224 1740
rect 7142 1682 7166 1716
rect 7200 1682 7224 1716
rect 7142 1658 7224 1682
rect 8644 1702 8726 1726
rect 8644 1668 8668 1702
rect 8702 1668 8726 1702
rect 8644 1644 8726 1668
rect 9662 1702 9744 1726
rect 9662 1668 9686 1702
rect 9720 1668 9744 1702
rect 9662 1644 9744 1668
rect 10680 1702 10762 1726
rect 10680 1668 10704 1702
rect 10738 1668 10762 1702
rect 10680 1644 10762 1668
rect 11698 1702 11780 1726
rect 11698 1668 11722 1702
rect 11756 1668 11780 1702
rect 11698 1644 11780 1668
rect 14016 1608 14098 1632
rect 14016 1574 14040 1608
rect 14074 1574 14098 1608
rect 14016 1550 14098 1574
rect 15034 1608 15116 1632
rect 15034 1574 15058 1608
rect 15092 1574 15116 1608
rect 15034 1550 15116 1574
rect 16052 1608 16134 1632
rect 16052 1574 16076 1608
rect 16110 1574 16134 1608
rect 16052 1550 16134 1574
rect 17070 1608 17152 1632
rect 17070 1574 17094 1608
rect 17128 1574 17152 1608
rect 17070 1550 17152 1574
rect 18088 1608 18170 1632
rect 18088 1574 18112 1608
rect 18146 1574 18170 1608
rect 18088 1550 18170 1574
rect 19106 1608 19188 1632
rect 19106 1574 19130 1608
rect 19164 1574 19188 1608
rect 19106 1550 19188 1574
rect 20124 1608 20206 1632
rect 20124 1574 20148 1608
rect 20182 1574 20206 1608
rect 20124 1550 20206 1574
rect 21142 1608 21224 1632
rect 21142 1574 21166 1608
rect 21200 1574 21224 1608
rect 21142 1550 21224 1574
rect 22160 1608 22242 1632
rect 22160 1574 22184 1608
rect 22218 1574 22242 1608
rect 22160 1550 22242 1574
rect 23178 1608 23260 1632
rect 23178 1574 23202 1608
rect 23236 1574 23260 1608
rect 23178 1550 23260 1574
rect 24196 1608 24278 1632
rect 24196 1574 24220 1608
rect 24254 1574 24278 1608
rect 24196 1550 24278 1574
rect 25214 1608 25296 1632
rect 25214 1574 25238 1608
rect 25272 1574 25296 1608
rect 25214 1550 25296 1574
rect 26232 1608 26314 1632
rect 26232 1574 26256 1608
rect 26290 1574 26314 1608
rect 26232 1550 26314 1574
rect 27250 1608 27332 1632
rect 27250 1574 27274 1608
rect 27308 1574 27332 1608
rect 27250 1550 27332 1574
rect 28268 1608 28350 1632
rect 28268 1574 28292 1608
rect 28326 1574 28350 1608
rect 28268 1550 28350 1574
rect 29286 1608 29368 1632
rect 29286 1574 29310 1608
rect 29344 1574 29368 1608
rect 29286 1550 29368 1574
rect 30304 1608 30386 1632
rect 30304 1574 30328 1608
rect 30362 1574 30386 1608
rect 30304 1550 30386 1574
rect 31322 1608 31404 1632
rect 31322 1574 31346 1608
rect 31380 1574 31404 1608
rect 31322 1550 31404 1574
rect 32340 1608 32422 1632
rect 32340 1574 32364 1608
rect 32398 1574 32422 1608
rect 32340 1550 32422 1574
rect 33358 1608 33440 1632
rect 33358 1574 33382 1608
rect 33416 1574 33440 1608
rect 33358 1550 33440 1574
rect 2026 522 2108 546
rect 2026 488 2050 522
rect 2084 488 2108 522
rect 2026 464 2108 488
rect 3044 522 3126 546
rect 3044 488 3068 522
rect 3102 488 3126 522
rect 3044 464 3126 488
rect 4062 522 4144 546
rect 4062 488 4086 522
rect 4120 488 4144 522
rect 4062 464 4144 488
rect 5080 522 5162 546
rect 5080 488 5104 522
rect 5138 488 5162 522
rect 5080 464 5162 488
rect 6098 522 6180 546
rect 6098 488 6122 522
rect 6156 488 6180 522
rect 6098 464 6180 488
rect 7116 522 7198 546
rect 7116 488 7140 522
rect 7174 488 7198 522
rect 7116 464 7198 488
rect 8618 468 8700 492
rect 8618 434 8642 468
rect 8676 434 8700 468
rect 8618 410 8700 434
rect 9636 468 9718 492
rect 9636 434 9660 468
rect 9694 434 9718 468
rect 9636 410 9718 434
rect 10654 468 10736 492
rect 10654 434 10678 468
rect 10712 434 10736 468
rect 10654 410 10736 434
rect 11672 468 11754 492
rect 11672 434 11696 468
rect 11730 434 11754 468
rect 11672 410 11754 434
rect -1372 -582 -1272 -520
rect 52628 15262 52790 15362
rect 89710 15262 89872 15362
rect 52628 15200 52728 15262
rect 48690 7480 48786 7514
rect 50404 7480 50500 7514
rect 48690 7418 48724 7480
rect 50466 7418 50500 7480
rect 48690 7000 48724 7062
rect 50466 7000 50500 7062
rect 48690 6966 48786 7000
rect 50404 6966 50500 7000
rect 48690 5516 48786 5550
rect 50404 5516 50500 5550
rect 48690 5454 48724 5516
rect 50466 5454 50500 5516
rect 48690 5036 48724 5098
rect 50466 5036 50500 5098
rect 48690 5002 48786 5036
rect 50404 5002 50500 5036
rect 48690 3516 48786 3550
rect 50404 3516 50500 3550
rect 48690 3454 48724 3516
rect 50466 3454 50500 3516
rect 48690 3036 48724 3098
rect 50466 3036 50500 3098
rect 48690 3002 48786 3036
rect 50404 3002 50500 3036
rect 48690 1426 48786 1460
rect 50404 1426 50500 1460
rect 48690 1364 48724 1426
rect 50466 1364 50500 1426
rect 48690 946 48724 1008
rect 50466 946 50500 1008
rect 48690 912 48786 946
rect 50404 912 50500 946
rect 35772 -582 35872 -520
rect -1372 -682 -1210 -582
rect 35710 -682 35872 -582
rect 89772 15200 89872 15262
rect 56282 14318 56364 14342
rect 56282 14284 56306 14318
rect 56340 14284 56364 14318
rect 56282 14260 56364 14284
rect 57300 14318 57382 14342
rect 57300 14284 57324 14318
rect 57358 14284 57382 14318
rect 57300 14260 57382 14284
rect 58318 14318 58400 14342
rect 58318 14284 58342 14318
rect 58376 14284 58400 14318
rect 58318 14260 58400 14284
rect 59336 14318 59418 14342
rect 59336 14284 59360 14318
rect 59394 14284 59418 14318
rect 59336 14260 59418 14284
rect 60354 14318 60436 14342
rect 60354 14284 60378 14318
rect 60412 14284 60436 14318
rect 60354 14260 60436 14284
rect 61372 14318 61454 14342
rect 61372 14284 61396 14318
rect 61430 14284 61454 14318
rect 61372 14260 61454 14284
rect 62390 14318 62472 14342
rect 62390 14284 62414 14318
rect 62448 14284 62472 14318
rect 62390 14260 62472 14284
rect 63408 14318 63490 14342
rect 63408 14284 63432 14318
rect 63466 14284 63490 14318
rect 63408 14260 63490 14284
rect 64426 14318 64508 14342
rect 64426 14284 64450 14318
rect 64484 14284 64508 14318
rect 64426 14260 64508 14284
rect 68016 13926 68098 13950
rect 68016 13892 68040 13926
rect 68074 13892 68098 13926
rect 68016 13868 68098 13892
rect 69034 13926 69116 13950
rect 69034 13892 69058 13926
rect 69092 13892 69116 13926
rect 69034 13868 69116 13892
rect 70052 13926 70134 13950
rect 70052 13892 70076 13926
rect 70110 13892 70134 13926
rect 70052 13868 70134 13892
rect 71070 13926 71152 13950
rect 71070 13892 71094 13926
rect 71128 13892 71152 13926
rect 71070 13868 71152 13892
rect 72088 13926 72170 13950
rect 72088 13892 72112 13926
rect 72146 13892 72170 13926
rect 72088 13868 72170 13892
rect 73106 13926 73188 13950
rect 73106 13892 73130 13926
rect 73164 13892 73188 13926
rect 73106 13868 73188 13892
rect 74124 13926 74206 13950
rect 74124 13892 74148 13926
rect 74182 13892 74206 13926
rect 74124 13868 74206 13892
rect 75142 13926 75224 13950
rect 75142 13892 75166 13926
rect 75200 13892 75224 13926
rect 75142 13868 75224 13892
rect 76160 13926 76242 13950
rect 76160 13892 76184 13926
rect 76218 13892 76242 13926
rect 76160 13868 76242 13892
rect 77178 13926 77260 13950
rect 77178 13892 77202 13926
rect 77236 13892 77260 13926
rect 77178 13868 77260 13892
rect 78196 13926 78278 13950
rect 78196 13892 78220 13926
rect 78254 13892 78278 13926
rect 78196 13868 78278 13892
rect 79214 13926 79296 13950
rect 79214 13892 79238 13926
rect 79272 13892 79296 13926
rect 79214 13868 79296 13892
rect 80232 13926 80314 13950
rect 80232 13892 80256 13926
rect 80290 13892 80314 13926
rect 80232 13868 80314 13892
rect 81250 13926 81332 13950
rect 81250 13892 81274 13926
rect 81308 13892 81332 13926
rect 81250 13868 81332 13892
rect 82268 13926 82350 13950
rect 82268 13892 82292 13926
rect 82326 13892 82350 13926
rect 82268 13868 82350 13892
rect 83286 13926 83368 13950
rect 83286 13892 83310 13926
rect 83344 13892 83368 13926
rect 83286 13868 83368 13892
rect 84304 13926 84386 13950
rect 84304 13892 84328 13926
rect 84362 13892 84386 13926
rect 84304 13868 84386 13892
rect 85322 13926 85404 13950
rect 85322 13892 85346 13926
rect 85380 13892 85404 13926
rect 85322 13868 85404 13892
rect 86340 13926 86422 13950
rect 86340 13892 86364 13926
rect 86398 13892 86422 13926
rect 86340 13868 86422 13892
rect 87358 13926 87440 13950
rect 87358 13892 87382 13926
rect 87416 13892 87440 13926
rect 87358 13868 87440 13892
rect 55744 13336 55826 13360
rect 55744 13302 55768 13336
rect 55802 13302 55826 13336
rect 55744 13278 55826 13302
rect 56762 13336 56844 13360
rect 56762 13302 56786 13336
rect 56820 13302 56844 13336
rect 56762 13278 56844 13302
rect 57780 13336 57862 13360
rect 57780 13302 57804 13336
rect 57838 13302 57862 13336
rect 57780 13278 57862 13302
rect 58798 13336 58880 13360
rect 58798 13302 58822 13336
rect 58856 13302 58880 13336
rect 58798 13278 58880 13302
rect 59816 13336 59898 13360
rect 59816 13302 59840 13336
rect 59874 13302 59898 13336
rect 59816 13278 59898 13302
rect 60834 13336 60916 13360
rect 60834 13302 60858 13336
rect 60892 13302 60916 13336
rect 60834 13278 60916 13302
rect 61852 13336 61934 13360
rect 61852 13302 61876 13336
rect 61910 13302 61934 13336
rect 61852 13278 61934 13302
rect 62870 13336 62952 13360
rect 62870 13302 62894 13336
rect 62928 13302 62952 13336
rect 62870 13278 62952 13302
rect 63888 13336 63970 13360
rect 63888 13302 63912 13336
rect 63946 13302 63970 13336
rect 63888 13278 63970 13302
rect 64906 13336 64988 13360
rect 64906 13302 64930 13336
rect 64964 13302 64988 13336
rect 64906 13278 64988 13302
rect 68004 12690 68086 12714
rect 68004 12656 68028 12690
rect 68062 12656 68086 12690
rect 68004 12632 68086 12656
rect 69022 12690 69104 12714
rect 69022 12656 69046 12690
rect 69080 12656 69104 12690
rect 69022 12632 69104 12656
rect 70040 12690 70122 12714
rect 70040 12656 70064 12690
rect 70098 12656 70122 12690
rect 70040 12632 70122 12656
rect 71058 12690 71140 12714
rect 71058 12656 71082 12690
rect 71116 12656 71140 12690
rect 71058 12632 71140 12656
rect 72076 12690 72158 12714
rect 72076 12656 72100 12690
rect 72134 12656 72158 12690
rect 72076 12632 72158 12656
rect 73094 12690 73176 12714
rect 73094 12656 73118 12690
rect 73152 12656 73176 12690
rect 73094 12632 73176 12656
rect 74112 12690 74194 12714
rect 74112 12656 74136 12690
rect 74170 12656 74194 12690
rect 74112 12632 74194 12656
rect 75130 12690 75212 12714
rect 75130 12656 75154 12690
rect 75188 12656 75212 12690
rect 75130 12632 75212 12656
rect 76148 12690 76230 12714
rect 76148 12656 76172 12690
rect 76206 12656 76230 12690
rect 76148 12632 76230 12656
rect 77166 12690 77248 12714
rect 77166 12656 77190 12690
rect 77224 12656 77248 12690
rect 77166 12632 77248 12656
rect 78184 12690 78266 12714
rect 78184 12656 78208 12690
rect 78242 12656 78266 12690
rect 78184 12632 78266 12656
rect 79202 12690 79284 12714
rect 79202 12656 79226 12690
rect 79260 12656 79284 12690
rect 79202 12632 79284 12656
rect 80220 12690 80302 12714
rect 80220 12656 80244 12690
rect 80278 12656 80302 12690
rect 80220 12632 80302 12656
rect 81238 12690 81320 12714
rect 81238 12656 81262 12690
rect 81296 12656 81320 12690
rect 81238 12632 81320 12656
rect 82256 12690 82338 12714
rect 82256 12656 82280 12690
rect 82314 12656 82338 12690
rect 82256 12632 82338 12656
rect 83274 12690 83356 12714
rect 83274 12656 83298 12690
rect 83332 12656 83356 12690
rect 83274 12632 83356 12656
rect 84292 12690 84374 12714
rect 84292 12656 84316 12690
rect 84350 12656 84374 12690
rect 84292 12632 84374 12656
rect 85310 12690 85392 12714
rect 85310 12656 85334 12690
rect 85368 12656 85392 12690
rect 85310 12632 85392 12656
rect 86328 12690 86410 12714
rect 86328 12656 86352 12690
rect 86386 12656 86410 12690
rect 86328 12632 86410 12656
rect 87346 12690 87428 12714
rect 87346 12656 87370 12690
rect 87404 12656 87428 12690
rect 87346 12632 87428 12656
rect 55744 12518 55826 12542
rect 55744 12484 55768 12518
rect 55802 12484 55826 12518
rect 55744 12460 55826 12484
rect 56762 12518 56844 12542
rect 56762 12484 56786 12518
rect 56820 12484 56844 12518
rect 56762 12460 56844 12484
rect 57780 12518 57862 12542
rect 57780 12484 57804 12518
rect 57838 12484 57862 12518
rect 57780 12460 57862 12484
rect 58798 12518 58880 12542
rect 58798 12484 58822 12518
rect 58856 12484 58880 12518
rect 58798 12460 58880 12484
rect 59816 12518 59898 12542
rect 59816 12484 59840 12518
rect 59874 12484 59898 12518
rect 59816 12460 59898 12484
rect 60834 12518 60916 12542
rect 60834 12484 60858 12518
rect 60892 12484 60916 12518
rect 60834 12460 60916 12484
rect 61852 12518 61934 12542
rect 61852 12484 61876 12518
rect 61910 12484 61934 12518
rect 61852 12460 61934 12484
rect 62870 12518 62952 12542
rect 62870 12484 62894 12518
rect 62928 12484 62952 12518
rect 62870 12460 62952 12484
rect 63888 12518 63970 12542
rect 63888 12484 63912 12518
rect 63946 12484 63970 12518
rect 63888 12460 63970 12484
rect 64906 12518 64988 12542
rect 64906 12484 64930 12518
rect 64964 12484 64988 12518
rect 64906 12460 64988 12484
rect 55744 11700 55826 11724
rect 55744 11666 55768 11700
rect 55802 11666 55826 11700
rect 55744 11642 55826 11666
rect 56762 11700 56844 11724
rect 56762 11666 56786 11700
rect 56820 11666 56844 11700
rect 56762 11642 56844 11666
rect 57780 11700 57862 11724
rect 57780 11666 57804 11700
rect 57838 11666 57862 11700
rect 57780 11642 57862 11666
rect 58798 11700 58880 11724
rect 58798 11666 58822 11700
rect 58856 11666 58880 11700
rect 58798 11642 58880 11666
rect 59816 11700 59898 11724
rect 59816 11666 59840 11700
rect 59874 11666 59898 11700
rect 59816 11642 59898 11666
rect 60834 11700 60916 11724
rect 60834 11666 60858 11700
rect 60892 11666 60916 11700
rect 60834 11642 60916 11666
rect 61852 11700 61934 11724
rect 61852 11666 61876 11700
rect 61910 11666 61934 11700
rect 61852 11642 61934 11666
rect 62870 11700 62952 11724
rect 62870 11666 62894 11700
rect 62928 11666 62952 11700
rect 62870 11642 62952 11666
rect 63888 11700 63970 11724
rect 63888 11666 63912 11700
rect 63946 11666 63970 11700
rect 63888 11642 63970 11666
rect 64906 11700 64988 11724
rect 64906 11666 64930 11700
rect 64964 11666 64988 11700
rect 64906 11642 64988 11666
rect 68016 11456 68098 11480
rect 68016 11422 68040 11456
rect 68074 11422 68098 11456
rect 68016 11398 68098 11422
rect 69034 11456 69116 11480
rect 69034 11422 69058 11456
rect 69092 11422 69116 11456
rect 69034 11398 69116 11422
rect 70052 11456 70134 11480
rect 70052 11422 70076 11456
rect 70110 11422 70134 11456
rect 70052 11398 70134 11422
rect 71070 11456 71152 11480
rect 71070 11422 71094 11456
rect 71128 11422 71152 11456
rect 71070 11398 71152 11422
rect 72088 11456 72170 11480
rect 72088 11422 72112 11456
rect 72146 11422 72170 11456
rect 72088 11398 72170 11422
rect 73106 11456 73188 11480
rect 73106 11422 73130 11456
rect 73164 11422 73188 11456
rect 73106 11398 73188 11422
rect 74124 11456 74206 11480
rect 74124 11422 74148 11456
rect 74182 11422 74206 11456
rect 74124 11398 74206 11422
rect 75142 11456 75224 11480
rect 75142 11422 75166 11456
rect 75200 11422 75224 11456
rect 75142 11398 75224 11422
rect 76160 11456 76242 11480
rect 76160 11422 76184 11456
rect 76218 11422 76242 11456
rect 76160 11398 76242 11422
rect 77178 11456 77260 11480
rect 77178 11422 77202 11456
rect 77236 11422 77260 11456
rect 77178 11398 77260 11422
rect 78196 11456 78278 11480
rect 78196 11422 78220 11456
rect 78254 11422 78278 11456
rect 78196 11398 78278 11422
rect 79214 11456 79296 11480
rect 79214 11422 79238 11456
rect 79272 11422 79296 11456
rect 79214 11398 79296 11422
rect 80232 11456 80314 11480
rect 80232 11422 80256 11456
rect 80290 11422 80314 11456
rect 80232 11398 80314 11422
rect 81250 11456 81332 11480
rect 81250 11422 81274 11456
rect 81308 11422 81332 11456
rect 81250 11398 81332 11422
rect 82268 11456 82350 11480
rect 82268 11422 82292 11456
rect 82326 11422 82350 11456
rect 82268 11398 82350 11422
rect 83286 11456 83368 11480
rect 83286 11422 83310 11456
rect 83344 11422 83368 11456
rect 83286 11398 83368 11422
rect 84304 11456 84386 11480
rect 84304 11422 84328 11456
rect 84362 11422 84386 11456
rect 84304 11398 84386 11422
rect 85322 11456 85404 11480
rect 85322 11422 85346 11456
rect 85380 11422 85404 11456
rect 85322 11398 85404 11422
rect 86340 11456 86422 11480
rect 86340 11422 86364 11456
rect 86398 11422 86422 11456
rect 86340 11398 86422 11422
rect 87358 11456 87440 11480
rect 87358 11422 87382 11456
rect 87416 11422 87440 11456
rect 87358 11398 87440 11422
rect 55744 10882 55826 10906
rect 55744 10848 55768 10882
rect 55802 10848 55826 10882
rect 55744 10824 55826 10848
rect 56762 10882 56844 10906
rect 56762 10848 56786 10882
rect 56820 10848 56844 10882
rect 56762 10824 56844 10848
rect 57780 10882 57862 10906
rect 57780 10848 57804 10882
rect 57838 10848 57862 10882
rect 57780 10824 57862 10848
rect 58798 10882 58880 10906
rect 58798 10848 58822 10882
rect 58856 10848 58880 10882
rect 58798 10824 58880 10848
rect 59816 10882 59898 10906
rect 59816 10848 59840 10882
rect 59874 10848 59898 10882
rect 59816 10824 59898 10848
rect 60834 10882 60916 10906
rect 60834 10848 60858 10882
rect 60892 10848 60916 10882
rect 60834 10824 60916 10848
rect 61852 10882 61934 10906
rect 61852 10848 61876 10882
rect 61910 10848 61934 10882
rect 61852 10824 61934 10848
rect 62870 10882 62952 10906
rect 62870 10848 62894 10882
rect 62928 10848 62952 10882
rect 62870 10824 62952 10848
rect 63888 10882 63970 10906
rect 63888 10848 63912 10882
rect 63946 10848 63970 10882
rect 63888 10824 63970 10848
rect 64906 10882 64988 10906
rect 64906 10848 64930 10882
rect 64964 10848 64988 10882
rect 64906 10824 64988 10848
rect 68016 10236 68098 10260
rect 68016 10202 68040 10236
rect 68074 10202 68098 10236
rect 68016 10178 68098 10202
rect 69034 10236 69116 10260
rect 69034 10202 69058 10236
rect 69092 10202 69116 10236
rect 69034 10178 69116 10202
rect 70052 10236 70134 10260
rect 70052 10202 70076 10236
rect 70110 10202 70134 10236
rect 70052 10178 70134 10202
rect 71070 10236 71152 10260
rect 71070 10202 71094 10236
rect 71128 10202 71152 10236
rect 71070 10178 71152 10202
rect 72088 10236 72170 10260
rect 72088 10202 72112 10236
rect 72146 10202 72170 10236
rect 72088 10178 72170 10202
rect 73106 10236 73188 10260
rect 73106 10202 73130 10236
rect 73164 10202 73188 10236
rect 73106 10178 73188 10202
rect 74124 10236 74206 10260
rect 74124 10202 74148 10236
rect 74182 10202 74206 10236
rect 74124 10178 74206 10202
rect 75142 10236 75224 10260
rect 75142 10202 75166 10236
rect 75200 10202 75224 10236
rect 75142 10178 75224 10202
rect 76160 10236 76242 10260
rect 76160 10202 76184 10236
rect 76218 10202 76242 10236
rect 76160 10178 76242 10202
rect 77178 10236 77260 10260
rect 77178 10202 77202 10236
rect 77236 10202 77260 10236
rect 77178 10178 77260 10202
rect 78196 10236 78278 10260
rect 78196 10202 78220 10236
rect 78254 10202 78278 10236
rect 78196 10178 78278 10202
rect 79214 10236 79296 10260
rect 79214 10202 79238 10236
rect 79272 10202 79296 10236
rect 79214 10178 79296 10202
rect 80232 10236 80314 10260
rect 80232 10202 80256 10236
rect 80290 10202 80314 10236
rect 80232 10178 80314 10202
rect 81250 10236 81332 10260
rect 81250 10202 81274 10236
rect 81308 10202 81332 10236
rect 81250 10178 81332 10202
rect 82268 10236 82350 10260
rect 82268 10202 82292 10236
rect 82326 10202 82350 10236
rect 82268 10178 82350 10202
rect 83286 10236 83368 10260
rect 83286 10202 83310 10236
rect 83344 10202 83368 10236
rect 83286 10178 83368 10202
rect 84304 10236 84386 10260
rect 84304 10202 84328 10236
rect 84362 10202 84386 10236
rect 84304 10178 84386 10202
rect 85322 10236 85404 10260
rect 85322 10202 85346 10236
rect 85380 10202 85404 10236
rect 85322 10178 85404 10202
rect 86340 10236 86422 10260
rect 86340 10202 86364 10236
rect 86398 10202 86422 10236
rect 86340 10178 86422 10202
rect 87358 10236 87440 10260
rect 87358 10202 87382 10236
rect 87416 10202 87440 10236
rect 87358 10178 87440 10202
rect 55744 10064 55826 10088
rect 55744 10030 55768 10064
rect 55802 10030 55826 10064
rect 55744 10006 55826 10030
rect 56762 10064 56844 10088
rect 56762 10030 56786 10064
rect 56820 10030 56844 10064
rect 56762 10006 56844 10030
rect 57780 10064 57862 10088
rect 57780 10030 57804 10064
rect 57838 10030 57862 10064
rect 57780 10006 57862 10030
rect 58798 10064 58880 10088
rect 58798 10030 58822 10064
rect 58856 10030 58880 10064
rect 58798 10006 58880 10030
rect 59816 10064 59898 10088
rect 59816 10030 59840 10064
rect 59874 10030 59898 10064
rect 59816 10006 59898 10030
rect 60834 10064 60916 10088
rect 60834 10030 60858 10064
rect 60892 10030 60916 10064
rect 60834 10006 60916 10030
rect 61852 10064 61934 10088
rect 61852 10030 61876 10064
rect 61910 10030 61934 10064
rect 61852 10006 61934 10030
rect 62870 10064 62952 10088
rect 62870 10030 62894 10064
rect 62928 10030 62952 10064
rect 62870 10006 62952 10030
rect 63888 10064 63970 10088
rect 63888 10030 63912 10064
rect 63946 10030 63970 10064
rect 63888 10006 63970 10030
rect 64906 10064 64988 10088
rect 64906 10030 64930 10064
rect 64964 10030 64988 10064
rect 64906 10006 64988 10030
rect 55744 9246 55826 9270
rect 55744 9212 55768 9246
rect 55802 9212 55826 9246
rect 55744 9188 55826 9212
rect 56762 9246 56844 9270
rect 56762 9212 56786 9246
rect 56820 9212 56844 9246
rect 56762 9188 56844 9212
rect 57780 9246 57862 9270
rect 57780 9212 57804 9246
rect 57838 9212 57862 9246
rect 57780 9188 57862 9212
rect 58798 9246 58880 9270
rect 58798 9212 58822 9246
rect 58856 9212 58880 9246
rect 58798 9188 58880 9212
rect 59816 9246 59898 9270
rect 59816 9212 59840 9246
rect 59874 9212 59898 9246
rect 59816 9188 59898 9212
rect 60834 9246 60916 9270
rect 60834 9212 60858 9246
rect 60892 9212 60916 9246
rect 60834 9188 60916 9212
rect 61852 9246 61934 9270
rect 61852 9212 61876 9246
rect 61910 9212 61934 9246
rect 61852 9188 61934 9212
rect 62870 9246 62952 9270
rect 62870 9212 62894 9246
rect 62928 9212 62952 9246
rect 62870 9188 62952 9212
rect 63888 9246 63970 9270
rect 63888 9212 63912 9246
rect 63946 9212 63970 9246
rect 63888 9188 63970 9212
rect 64906 9246 64988 9270
rect 64906 9212 64930 9246
rect 64964 9212 64988 9246
rect 64906 9188 64988 9212
rect 68030 8988 68112 9012
rect 68030 8954 68054 8988
rect 68088 8954 68112 8988
rect 68030 8930 68112 8954
rect 69048 8988 69130 9012
rect 69048 8954 69072 8988
rect 69106 8954 69130 8988
rect 69048 8930 69130 8954
rect 70066 8988 70148 9012
rect 70066 8954 70090 8988
rect 70124 8954 70148 8988
rect 70066 8930 70148 8954
rect 71084 8988 71166 9012
rect 71084 8954 71108 8988
rect 71142 8954 71166 8988
rect 71084 8930 71166 8954
rect 72102 8988 72184 9012
rect 72102 8954 72126 8988
rect 72160 8954 72184 8988
rect 72102 8930 72184 8954
rect 73120 8988 73202 9012
rect 73120 8954 73144 8988
rect 73178 8954 73202 8988
rect 73120 8930 73202 8954
rect 74138 8988 74220 9012
rect 74138 8954 74162 8988
rect 74196 8954 74220 8988
rect 74138 8930 74220 8954
rect 75156 8988 75238 9012
rect 75156 8954 75180 8988
rect 75214 8954 75238 8988
rect 75156 8930 75238 8954
rect 76174 8988 76256 9012
rect 76174 8954 76198 8988
rect 76232 8954 76256 8988
rect 76174 8930 76256 8954
rect 77192 8988 77274 9012
rect 77192 8954 77216 8988
rect 77250 8954 77274 8988
rect 77192 8930 77274 8954
rect 78210 8988 78292 9012
rect 78210 8954 78234 8988
rect 78268 8954 78292 8988
rect 78210 8930 78292 8954
rect 79228 8988 79310 9012
rect 79228 8954 79252 8988
rect 79286 8954 79310 8988
rect 79228 8930 79310 8954
rect 80246 8988 80328 9012
rect 80246 8954 80270 8988
rect 80304 8954 80328 8988
rect 80246 8930 80328 8954
rect 81264 8988 81346 9012
rect 81264 8954 81288 8988
rect 81322 8954 81346 8988
rect 81264 8930 81346 8954
rect 82282 8988 82364 9012
rect 82282 8954 82306 8988
rect 82340 8954 82364 8988
rect 82282 8930 82364 8954
rect 83300 8988 83382 9012
rect 83300 8954 83324 8988
rect 83358 8954 83382 8988
rect 83300 8930 83382 8954
rect 84318 8988 84400 9012
rect 84318 8954 84342 8988
rect 84376 8954 84400 8988
rect 84318 8930 84400 8954
rect 85336 8988 85418 9012
rect 85336 8954 85360 8988
rect 85394 8954 85418 8988
rect 85336 8930 85418 8954
rect 86354 8988 86436 9012
rect 86354 8954 86378 8988
rect 86412 8954 86436 8988
rect 86354 8930 86436 8954
rect 87372 8988 87454 9012
rect 87372 8954 87396 8988
rect 87430 8954 87454 8988
rect 87372 8930 87454 8954
rect 55744 8428 55826 8452
rect 55744 8394 55768 8428
rect 55802 8394 55826 8428
rect 55744 8370 55826 8394
rect 56762 8428 56844 8452
rect 56762 8394 56786 8428
rect 56820 8394 56844 8428
rect 56762 8370 56844 8394
rect 57780 8428 57862 8452
rect 57780 8394 57804 8428
rect 57838 8394 57862 8428
rect 57780 8370 57862 8394
rect 58798 8428 58880 8452
rect 58798 8394 58822 8428
rect 58856 8394 58880 8428
rect 58798 8370 58880 8394
rect 59816 8428 59898 8452
rect 59816 8394 59840 8428
rect 59874 8394 59898 8428
rect 59816 8370 59898 8394
rect 60834 8428 60916 8452
rect 60834 8394 60858 8428
rect 60892 8394 60916 8428
rect 60834 8370 60916 8394
rect 61852 8428 61934 8452
rect 61852 8394 61876 8428
rect 61910 8394 61934 8428
rect 61852 8370 61934 8394
rect 62870 8428 62952 8452
rect 62870 8394 62894 8428
rect 62928 8394 62952 8428
rect 62870 8370 62952 8394
rect 63888 8428 63970 8452
rect 63888 8394 63912 8428
rect 63946 8394 63970 8428
rect 63888 8370 63970 8394
rect 64906 8428 64988 8452
rect 64906 8394 64930 8428
rect 64964 8394 64988 8428
rect 64906 8370 64988 8394
rect 68016 7766 68098 7790
rect 68016 7732 68040 7766
rect 68074 7732 68098 7766
rect 68016 7708 68098 7732
rect 69034 7766 69116 7790
rect 69034 7732 69058 7766
rect 69092 7732 69116 7766
rect 69034 7708 69116 7732
rect 70052 7766 70134 7790
rect 70052 7732 70076 7766
rect 70110 7732 70134 7766
rect 70052 7708 70134 7732
rect 71070 7766 71152 7790
rect 71070 7732 71094 7766
rect 71128 7732 71152 7766
rect 71070 7708 71152 7732
rect 72088 7766 72170 7790
rect 72088 7732 72112 7766
rect 72146 7732 72170 7766
rect 72088 7708 72170 7732
rect 73106 7766 73188 7790
rect 73106 7732 73130 7766
rect 73164 7732 73188 7766
rect 73106 7708 73188 7732
rect 74124 7766 74206 7790
rect 74124 7732 74148 7766
rect 74182 7732 74206 7766
rect 74124 7708 74206 7732
rect 75142 7766 75224 7790
rect 75142 7732 75166 7766
rect 75200 7732 75224 7766
rect 75142 7708 75224 7732
rect 76160 7766 76242 7790
rect 76160 7732 76184 7766
rect 76218 7732 76242 7766
rect 76160 7708 76242 7732
rect 77178 7766 77260 7790
rect 77178 7732 77202 7766
rect 77236 7732 77260 7766
rect 77178 7708 77260 7732
rect 78196 7766 78278 7790
rect 78196 7732 78220 7766
rect 78254 7732 78278 7766
rect 78196 7708 78278 7732
rect 79214 7766 79296 7790
rect 79214 7732 79238 7766
rect 79272 7732 79296 7766
rect 79214 7708 79296 7732
rect 80232 7766 80314 7790
rect 80232 7732 80256 7766
rect 80290 7732 80314 7766
rect 80232 7708 80314 7732
rect 81250 7766 81332 7790
rect 81250 7732 81274 7766
rect 81308 7732 81332 7766
rect 81250 7708 81332 7732
rect 82268 7766 82350 7790
rect 82268 7732 82292 7766
rect 82326 7732 82350 7766
rect 82268 7708 82350 7732
rect 83286 7766 83368 7790
rect 83286 7732 83310 7766
rect 83344 7732 83368 7766
rect 83286 7708 83368 7732
rect 84304 7766 84386 7790
rect 84304 7732 84328 7766
rect 84362 7732 84386 7766
rect 84304 7708 84386 7732
rect 85322 7766 85404 7790
rect 85322 7732 85346 7766
rect 85380 7732 85404 7766
rect 85322 7708 85404 7732
rect 86340 7766 86422 7790
rect 86340 7732 86364 7766
rect 86398 7732 86422 7766
rect 86340 7708 86422 7732
rect 87358 7766 87440 7790
rect 87358 7732 87382 7766
rect 87416 7732 87440 7766
rect 87358 7708 87440 7732
rect 56254 7386 56336 7410
rect 56254 7352 56278 7386
rect 56312 7352 56336 7386
rect 56254 7328 56336 7352
rect 57272 7386 57354 7410
rect 57272 7352 57296 7386
rect 57330 7352 57354 7386
rect 57272 7328 57354 7352
rect 58290 7386 58372 7410
rect 58290 7352 58314 7386
rect 58348 7352 58372 7386
rect 58290 7328 58372 7352
rect 59308 7386 59390 7410
rect 59308 7352 59332 7386
rect 59366 7352 59390 7386
rect 59308 7328 59390 7352
rect 60326 7386 60408 7410
rect 60326 7352 60350 7386
rect 60384 7352 60408 7386
rect 60326 7328 60408 7352
rect 61344 7386 61426 7410
rect 61344 7352 61368 7386
rect 61402 7352 61426 7386
rect 61344 7328 61426 7352
rect 62362 7386 62444 7410
rect 62362 7352 62386 7386
rect 62420 7352 62444 7386
rect 62362 7328 62444 7352
rect 63380 7386 63462 7410
rect 63380 7352 63404 7386
rect 63438 7352 63462 7386
rect 63380 7328 63462 7352
rect 64398 7386 64480 7410
rect 64398 7352 64422 7386
rect 64456 7352 64480 7386
rect 64398 7328 64480 7352
rect 68016 6518 68098 6542
rect 68016 6484 68040 6518
rect 68074 6484 68098 6518
rect 68016 6460 68098 6484
rect 69034 6518 69116 6542
rect 69034 6484 69058 6518
rect 69092 6484 69116 6518
rect 69034 6460 69116 6484
rect 70052 6518 70134 6542
rect 70052 6484 70076 6518
rect 70110 6484 70134 6518
rect 70052 6460 70134 6484
rect 71070 6518 71152 6542
rect 71070 6484 71094 6518
rect 71128 6484 71152 6518
rect 71070 6460 71152 6484
rect 72088 6518 72170 6542
rect 72088 6484 72112 6518
rect 72146 6484 72170 6518
rect 72088 6460 72170 6484
rect 73106 6518 73188 6542
rect 73106 6484 73130 6518
rect 73164 6484 73188 6518
rect 73106 6460 73188 6484
rect 74124 6518 74206 6542
rect 74124 6484 74148 6518
rect 74182 6484 74206 6518
rect 74124 6460 74206 6484
rect 75142 6518 75224 6542
rect 75142 6484 75166 6518
rect 75200 6484 75224 6518
rect 75142 6460 75224 6484
rect 76160 6518 76242 6542
rect 76160 6484 76184 6518
rect 76218 6484 76242 6518
rect 76160 6460 76242 6484
rect 77178 6518 77260 6542
rect 77178 6484 77202 6518
rect 77236 6484 77260 6518
rect 77178 6460 77260 6484
rect 78196 6518 78278 6542
rect 78196 6484 78220 6518
rect 78254 6484 78278 6518
rect 78196 6460 78278 6484
rect 79214 6518 79296 6542
rect 79214 6484 79238 6518
rect 79272 6484 79296 6518
rect 79214 6460 79296 6484
rect 80232 6518 80314 6542
rect 80232 6484 80256 6518
rect 80290 6484 80314 6518
rect 80232 6460 80314 6484
rect 81250 6518 81332 6542
rect 81250 6484 81274 6518
rect 81308 6484 81332 6518
rect 81250 6460 81332 6484
rect 82268 6518 82350 6542
rect 82268 6484 82292 6518
rect 82326 6484 82350 6518
rect 82268 6460 82350 6484
rect 83286 6518 83368 6542
rect 83286 6484 83310 6518
rect 83344 6484 83368 6518
rect 83286 6460 83368 6484
rect 84304 6518 84386 6542
rect 84304 6484 84328 6518
rect 84362 6484 84386 6518
rect 84304 6460 84386 6484
rect 85322 6518 85404 6542
rect 85322 6484 85346 6518
rect 85380 6484 85404 6518
rect 85322 6460 85404 6484
rect 86340 6518 86422 6542
rect 86340 6484 86364 6518
rect 86398 6484 86422 6518
rect 86340 6460 86422 6484
rect 87358 6518 87440 6542
rect 87358 6484 87382 6518
rect 87416 6484 87440 6518
rect 87358 6460 87440 6484
rect 62332 6410 62414 6434
rect 62332 6376 62356 6410
rect 62390 6376 62414 6410
rect 62332 6352 62414 6376
rect 63350 6410 63432 6434
rect 63350 6376 63374 6410
rect 63408 6376 63432 6410
rect 63350 6352 63432 6376
rect 64368 6410 64450 6434
rect 64368 6376 64392 6410
rect 64426 6376 64450 6410
rect 64368 6352 64450 6376
rect 65386 6410 65468 6434
rect 65386 6376 65410 6410
rect 65444 6376 65468 6410
rect 65386 6352 65468 6376
rect 68030 5298 68112 5322
rect 68030 5264 68054 5298
rect 68088 5264 68112 5298
rect 68030 5240 68112 5264
rect 69048 5298 69130 5322
rect 69048 5264 69072 5298
rect 69106 5264 69130 5298
rect 69048 5240 69130 5264
rect 70066 5298 70148 5322
rect 70066 5264 70090 5298
rect 70124 5264 70148 5298
rect 70066 5240 70148 5264
rect 71084 5298 71166 5322
rect 71084 5264 71108 5298
rect 71142 5264 71166 5298
rect 71084 5240 71166 5264
rect 72102 5298 72184 5322
rect 72102 5264 72126 5298
rect 72160 5264 72184 5298
rect 72102 5240 72184 5264
rect 73120 5298 73202 5322
rect 73120 5264 73144 5298
rect 73178 5264 73202 5298
rect 73120 5240 73202 5264
rect 74138 5298 74220 5322
rect 74138 5264 74162 5298
rect 74196 5264 74220 5298
rect 74138 5240 74220 5264
rect 75156 5298 75238 5322
rect 75156 5264 75180 5298
rect 75214 5264 75238 5298
rect 75156 5240 75238 5264
rect 76174 5298 76256 5322
rect 76174 5264 76198 5298
rect 76232 5264 76256 5298
rect 76174 5240 76256 5264
rect 77192 5298 77274 5322
rect 77192 5264 77216 5298
rect 77250 5264 77274 5298
rect 77192 5240 77274 5264
rect 78210 5298 78292 5322
rect 78210 5264 78234 5298
rect 78268 5264 78292 5298
rect 78210 5240 78292 5264
rect 79228 5298 79310 5322
rect 79228 5264 79252 5298
rect 79286 5264 79310 5298
rect 79228 5240 79310 5264
rect 80246 5298 80328 5322
rect 80246 5264 80270 5298
rect 80304 5264 80328 5298
rect 80246 5240 80328 5264
rect 81264 5298 81346 5322
rect 81264 5264 81288 5298
rect 81322 5264 81346 5298
rect 81264 5240 81346 5264
rect 82282 5298 82364 5322
rect 82282 5264 82306 5298
rect 82340 5264 82364 5298
rect 82282 5240 82364 5264
rect 83300 5298 83382 5322
rect 83300 5264 83324 5298
rect 83358 5264 83382 5298
rect 83300 5240 83382 5264
rect 84318 5298 84400 5322
rect 84318 5264 84342 5298
rect 84376 5264 84400 5298
rect 84318 5240 84400 5264
rect 85336 5298 85418 5322
rect 85336 5264 85360 5298
rect 85394 5264 85418 5298
rect 85336 5240 85418 5264
rect 86354 5298 86436 5322
rect 86354 5264 86378 5298
rect 86412 5264 86436 5298
rect 86354 5240 86436 5264
rect 87372 5298 87454 5322
rect 87372 5264 87396 5298
rect 87430 5264 87454 5298
rect 87372 5240 87454 5264
rect 62630 5122 62712 5146
rect 56038 5066 56120 5090
rect 56038 5032 56062 5066
rect 56096 5032 56120 5066
rect 56038 5008 56120 5032
rect 57056 5066 57138 5090
rect 57056 5032 57080 5066
rect 57114 5032 57138 5066
rect 57056 5008 57138 5032
rect 58074 5066 58156 5090
rect 58074 5032 58098 5066
rect 58132 5032 58156 5066
rect 58074 5008 58156 5032
rect 59092 5066 59174 5090
rect 59092 5032 59116 5066
rect 59150 5032 59174 5066
rect 59092 5008 59174 5032
rect 60110 5066 60192 5090
rect 60110 5032 60134 5066
rect 60168 5032 60192 5066
rect 60110 5008 60192 5032
rect 61128 5066 61210 5090
rect 61128 5032 61152 5066
rect 61186 5032 61210 5066
rect 62630 5088 62654 5122
rect 62688 5088 62712 5122
rect 62630 5064 62712 5088
rect 63648 5122 63730 5146
rect 63648 5088 63672 5122
rect 63706 5088 63730 5122
rect 63648 5064 63730 5088
rect 64666 5122 64748 5146
rect 64666 5088 64690 5122
rect 64724 5088 64748 5122
rect 64666 5064 64748 5088
rect 65684 5122 65766 5146
rect 65684 5088 65708 5122
rect 65742 5088 65766 5122
rect 65684 5064 65766 5088
rect 61128 5008 61210 5032
rect 68030 4050 68112 4074
rect 68030 4016 68054 4050
rect 68088 4016 68112 4050
rect 68030 3992 68112 4016
rect 69048 4050 69130 4074
rect 69048 4016 69072 4050
rect 69106 4016 69130 4050
rect 69048 3992 69130 4016
rect 70066 4050 70148 4074
rect 70066 4016 70090 4050
rect 70124 4016 70148 4050
rect 70066 3992 70148 4016
rect 71084 4050 71166 4074
rect 71084 4016 71108 4050
rect 71142 4016 71166 4050
rect 71084 3992 71166 4016
rect 72102 4050 72184 4074
rect 72102 4016 72126 4050
rect 72160 4016 72184 4050
rect 72102 3992 72184 4016
rect 73120 4050 73202 4074
rect 73120 4016 73144 4050
rect 73178 4016 73202 4050
rect 73120 3992 73202 4016
rect 74138 4050 74220 4074
rect 74138 4016 74162 4050
rect 74196 4016 74220 4050
rect 74138 3992 74220 4016
rect 75156 4050 75238 4074
rect 75156 4016 75180 4050
rect 75214 4016 75238 4050
rect 75156 3992 75238 4016
rect 76174 4050 76256 4074
rect 76174 4016 76198 4050
rect 76232 4016 76256 4050
rect 76174 3992 76256 4016
rect 77192 4050 77274 4074
rect 77192 4016 77216 4050
rect 77250 4016 77274 4050
rect 77192 3992 77274 4016
rect 78210 4050 78292 4074
rect 78210 4016 78234 4050
rect 78268 4016 78292 4050
rect 78210 3992 78292 4016
rect 79228 4050 79310 4074
rect 79228 4016 79252 4050
rect 79286 4016 79310 4050
rect 79228 3992 79310 4016
rect 80246 4050 80328 4074
rect 80246 4016 80270 4050
rect 80304 4016 80328 4050
rect 80246 3992 80328 4016
rect 81264 4050 81346 4074
rect 81264 4016 81288 4050
rect 81322 4016 81346 4050
rect 81264 3992 81346 4016
rect 82282 4050 82364 4074
rect 82282 4016 82306 4050
rect 82340 4016 82364 4050
rect 82282 3992 82364 4016
rect 83300 4050 83382 4074
rect 83300 4016 83324 4050
rect 83358 4016 83382 4050
rect 83300 3992 83382 4016
rect 84318 4050 84400 4074
rect 84318 4016 84342 4050
rect 84376 4016 84400 4050
rect 84318 3992 84400 4016
rect 85336 4050 85418 4074
rect 85336 4016 85360 4050
rect 85394 4016 85418 4050
rect 85336 3992 85418 4016
rect 86354 4050 86436 4074
rect 86354 4016 86378 4050
rect 86412 4016 86436 4050
rect 86354 3992 86436 4016
rect 87372 4050 87454 4074
rect 87372 4016 87396 4050
rect 87430 4016 87454 4050
rect 87372 3992 87454 4016
rect 56052 3940 56134 3964
rect 56052 3906 56076 3940
rect 56110 3906 56134 3940
rect 56052 3882 56134 3906
rect 57070 3940 57152 3964
rect 57070 3906 57094 3940
rect 57128 3906 57152 3940
rect 57070 3882 57152 3906
rect 58088 3940 58170 3964
rect 58088 3906 58112 3940
rect 58146 3906 58170 3940
rect 58088 3882 58170 3906
rect 59106 3940 59188 3964
rect 59106 3906 59130 3940
rect 59164 3906 59188 3940
rect 59106 3882 59188 3906
rect 60124 3940 60206 3964
rect 60124 3906 60148 3940
rect 60182 3906 60206 3940
rect 60124 3882 60206 3906
rect 61142 3940 61224 3964
rect 61142 3906 61166 3940
rect 61200 3906 61224 3940
rect 61142 3882 61224 3906
rect 62590 3928 62672 3952
rect 62590 3894 62614 3928
rect 62648 3894 62672 3928
rect 62590 3870 62672 3894
rect 63608 3928 63690 3952
rect 63608 3894 63632 3928
rect 63666 3894 63690 3928
rect 63608 3870 63690 3894
rect 64626 3928 64708 3952
rect 64626 3894 64650 3928
rect 64684 3894 64708 3928
rect 64626 3870 64708 3894
rect 65644 3928 65726 3952
rect 65644 3894 65668 3928
rect 65702 3894 65726 3928
rect 65644 3870 65726 3894
rect 56026 2814 56108 2838
rect 56026 2780 56050 2814
rect 56084 2780 56108 2814
rect 56026 2756 56108 2780
rect 57044 2814 57126 2838
rect 57044 2780 57068 2814
rect 57102 2780 57126 2814
rect 57044 2756 57126 2780
rect 58062 2814 58144 2838
rect 58062 2780 58086 2814
rect 58120 2780 58144 2814
rect 58062 2756 58144 2780
rect 59080 2814 59162 2838
rect 59080 2780 59104 2814
rect 59138 2780 59162 2814
rect 59080 2756 59162 2780
rect 60098 2814 60180 2838
rect 60098 2780 60122 2814
rect 60156 2780 60180 2814
rect 60098 2756 60180 2780
rect 61116 2814 61198 2838
rect 61116 2780 61140 2814
rect 61174 2780 61198 2814
rect 61116 2756 61198 2780
rect 62590 2814 62672 2838
rect 62590 2780 62614 2814
rect 62648 2780 62672 2814
rect 62590 2756 62672 2780
rect 63608 2814 63690 2838
rect 63608 2780 63632 2814
rect 63666 2780 63690 2814
rect 63608 2756 63690 2780
rect 64626 2814 64708 2838
rect 64626 2780 64650 2814
rect 64684 2780 64708 2814
rect 64626 2756 64708 2780
rect 65644 2814 65726 2838
rect 65644 2780 65668 2814
rect 65702 2780 65726 2814
rect 65644 2756 65726 2780
rect 68016 2828 68098 2852
rect 68016 2794 68040 2828
rect 68074 2794 68098 2828
rect 68016 2770 68098 2794
rect 69034 2828 69116 2852
rect 69034 2794 69058 2828
rect 69092 2794 69116 2828
rect 69034 2770 69116 2794
rect 70052 2828 70134 2852
rect 70052 2794 70076 2828
rect 70110 2794 70134 2828
rect 70052 2770 70134 2794
rect 71070 2828 71152 2852
rect 71070 2794 71094 2828
rect 71128 2794 71152 2828
rect 71070 2770 71152 2794
rect 72088 2828 72170 2852
rect 72088 2794 72112 2828
rect 72146 2794 72170 2828
rect 72088 2770 72170 2794
rect 73106 2828 73188 2852
rect 73106 2794 73130 2828
rect 73164 2794 73188 2828
rect 73106 2770 73188 2794
rect 74124 2828 74206 2852
rect 74124 2794 74148 2828
rect 74182 2794 74206 2828
rect 74124 2770 74206 2794
rect 75142 2828 75224 2852
rect 75142 2794 75166 2828
rect 75200 2794 75224 2828
rect 75142 2770 75224 2794
rect 76160 2828 76242 2852
rect 76160 2794 76184 2828
rect 76218 2794 76242 2828
rect 76160 2770 76242 2794
rect 77178 2828 77260 2852
rect 77178 2794 77202 2828
rect 77236 2794 77260 2828
rect 77178 2770 77260 2794
rect 78196 2828 78278 2852
rect 78196 2794 78220 2828
rect 78254 2794 78278 2828
rect 78196 2770 78278 2794
rect 79214 2828 79296 2852
rect 79214 2794 79238 2828
rect 79272 2794 79296 2828
rect 79214 2770 79296 2794
rect 80232 2828 80314 2852
rect 80232 2794 80256 2828
rect 80290 2794 80314 2828
rect 80232 2770 80314 2794
rect 81250 2828 81332 2852
rect 81250 2794 81274 2828
rect 81308 2794 81332 2828
rect 81250 2770 81332 2794
rect 82268 2828 82350 2852
rect 82268 2794 82292 2828
rect 82326 2794 82350 2828
rect 82268 2770 82350 2794
rect 83286 2828 83368 2852
rect 83286 2794 83310 2828
rect 83344 2794 83368 2828
rect 83286 2770 83368 2794
rect 84304 2828 84386 2852
rect 84304 2794 84328 2828
rect 84362 2794 84386 2828
rect 84304 2770 84386 2794
rect 85322 2828 85404 2852
rect 85322 2794 85346 2828
rect 85380 2794 85404 2828
rect 85322 2770 85404 2794
rect 86340 2828 86422 2852
rect 86340 2794 86364 2828
rect 86398 2794 86422 2828
rect 86340 2770 86422 2794
rect 87358 2828 87440 2852
rect 87358 2794 87382 2828
rect 87416 2794 87440 2828
rect 87358 2770 87440 2794
rect 56052 1716 56134 1740
rect 56052 1682 56076 1716
rect 56110 1682 56134 1716
rect 56052 1658 56134 1682
rect 57070 1716 57152 1740
rect 57070 1682 57094 1716
rect 57128 1682 57152 1716
rect 57070 1658 57152 1682
rect 58088 1716 58170 1740
rect 58088 1682 58112 1716
rect 58146 1682 58170 1716
rect 58088 1658 58170 1682
rect 59106 1716 59188 1740
rect 59106 1682 59130 1716
rect 59164 1682 59188 1716
rect 59106 1658 59188 1682
rect 60124 1716 60206 1740
rect 60124 1682 60148 1716
rect 60182 1682 60206 1716
rect 60124 1658 60206 1682
rect 61142 1716 61224 1740
rect 61142 1682 61166 1716
rect 61200 1682 61224 1716
rect 61142 1658 61224 1682
rect 62644 1702 62726 1726
rect 62644 1668 62668 1702
rect 62702 1668 62726 1702
rect 62644 1644 62726 1668
rect 63662 1702 63744 1726
rect 63662 1668 63686 1702
rect 63720 1668 63744 1702
rect 63662 1644 63744 1668
rect 64680 1702 64762 1726
rect 64680 1668 64704 1702
rect 64738 1668 64762 1702
rect 64680 1644 64762 1668
rect 65698 1702 65780 1726
rect 65698 1668 65722 1702
rect 65756 1668 65780 1702
rect 65698 1644 65780 1668
rect 68016 1608 68098 1632
rect 68016 1574 68040 1608
rect 68074 1574 68098 1608
rect 68016 1550 68098 1574
rect 69034 1608 69116 1632
rect 69034 1574 69058 1608
rect 69092 1574 69116 1608
rect 69034 1550 69116 1574
rect 70052 1608 70134 1632
rect 70052 1574 70076 1608
rect 70110 1574 70134 1608
rect 70052 1550 70134 1574
rect 71070 1608 71152 1632
rect 71070 1574 71094 1608
rect 71128 1574 71152 1608
rect 71070 1550 71152 1574
rect 72088 1608 72170 1632
rect 72088 1574 72112 1608
rect 72146 1574 72170 1608
rect 72088 1550 72170 1574
rect 73106 1608 73188 1632
rect 73106 1574 73130 1608
rect 73164 1574 73188 1608
rect 73106 1550 73188 1574
rect 74124 1608 74206 1632
rect 74124 1574 74148 1608
rect 74182 1574 74206 1608
rect 74124 1550 74206 1574
rect 75142 1608 75224 1632
rect 75142 1574 75166 1608
rect 75200 1574 75224 1608
rect 75142 1550 75224 1574
rect 76160 1608 76242 1632
rect 76160 1574 76184 1608
rect 76218 1574 76242 1608
rect 76160 1550 76242 1574
rect 77178 1608 77260 1632
rect 77178 1574 77202 1608
rect 77236 1574 77260 1608
rect 77178 1550 77260 1574
rect 78196 1608 78278 1632
rect 78196 1574 78220 1608
rect 78254 1574 78278 1608
rect 78196 1550 78278 1574
rect 79214 1608 79296 1632
rect 79214 1574 79238 1608
rect 79272 1574 79296 1608
rect 79214 1550 79296 1574
rect 80232 1608 80314 1632
rect 80232 1574 80256 1608
rect 80290 1574 80314 1608
rect 80232 1550 80314 1574
rect 81250 1608 81332 1632
rect 81250 1574 81274 1608
rect 81308 1574 81332 1608
rect 81250 1550 81332 1574
rect 82268 1608 82350 1632
rect 82268 1574 82292 1608
rect 82326 1574 82350 1608
rect 82268 1550 82350 1574
rect 83286 1608 83368 1632
rect 83286 1574 83310 1608
rect 83344 1574 83368 1608
rect 83286 1550 83368 1574
rect 84304 1608 84386 1632
rect 84304 1574 84328 1608
rect 84362 1574 84386 1608
rect 84304 1550 84386 1574
rect 85322 1608 85404 1632
rect 85322 1574 85346 1608
rect 85380 1574 85404 1608
rect 85322 1550 85404 1574
rect 86340 1608 86422 1632
rect 86340 1574 86364 1608
rect 86398 1574 86422 1608
rect 86340 1550 86422 1574
rect 87358 1608 87440 1632
rect 87358 1574 87382 1608
rect 87416 1574 87440 1608
rect 87358 1550 87440 1574
rect 56026 522 56108 546
rect 56026 488 56050 522
rect 56084 488 56108 522
rect 56026 464 56108 488
rect 57044 522 57126 546
rect 57044 488 57068 522
rect 57102 488 57126 522
rect 57044 464 57126 488
rect 58062 522 58144 546
rect 58062 488 58086 522
rect 58120 488 58144 522
rect 58062 464 58144 488
rect 59080 522 59162 546
rect 59080 488 59104 522
rect 59138 488 59162 522
rect 59080 464 59162 488
rect 60098 522 60180 546
rect 60098 488 60122 522
rect 60156 488 60180 522
rect 60098 464 60180 488
rect 61116 522 61198 546
rect 61116 488 61140 522
rect 61174 488 61198 522
rect 61116 464 61198 488
rect 62618 468 62700 492
rect 62618 434 62642 468
rect 62676 434 62700 468
rect 62618 410 62700 434
rect 63636 468 63718 492
rect 63636 434 63660 468
rect 63694 434 63718 468
rect 63636 410 63718 434
rect 64654 468 64736 492
rect 64654 434 64678 468
rect 64712 434 64736 468
rect 64654 410 64736 434
rect 65672 468 65754 492
rect 65672 434 65696 468
rect 65730 434 65754 468
rect 65672 410 65754 434
rect 52628 -582 52728 -520
rect 89772 -582 89872 -520
rect 52628 -682 52790 -582
rect 89710 -682 89872 -582
<< nsubdiff >>
rect 11328 28162 11490 28262
rect 35610 28162 35772 28262
rect 11328 28100 11428 28162
rect 35672 28100 35772 28162
rect 18940 26142 19022 26168
rect 18940 26108 18964 26142
rect 18998 26108 19022 26142
rect 18940 26084 19022 26108
rect 19958 26142 20040 26168
rect 19958 26108 19982 26142
rect 20016 26108 20040 26142
rect 19958 26084 20040 26108
rect 20976 26142 21058 26168
rect 20976 26108 21000 26142
rect 21034 26108 21058 26142
rect 20976 26084 21058 26108
rect 21994 26142 22076 26168
rect 21994 26108 22018 26142
rect 22052 26108 22076 26142
rect 21994 26084 22076 26108
rect 23012 26142 23094 26168
rect 23012 26108 23036 26142
rect 23070 26108 23094 26142
rect 23012 26084 23094 26108
rect 24030 26142 24112 26168
rect 24030 26108 24054 26142
rect 24088 26108 24112 26142
rect 24030 26084 24112 26108
rect 25048 26142 25130 26168
rect 25048 26108 25072 26142
rect 25106 26108 25130 26142
rect 25048 26084 25130 26108
rect 26066 26142 26148 26168
rect 26066 26108 26090 26142
rect 26124 26108 26148 26142
rect 26066 26084 26148 26108
rect 27084 26142 27166 26168
rect 27084 26108 27108 26142
rect 27142 26108 27166 26142
rect 27084 26084 27166 26108
rect 28102 26142 28184 26168
rect 28102 26108 28126 26142
rect 28160 26108 28184 26142
rect 28102 26084 28184 26108
rect 29120 26142 29202 26168
rect 29120 26108 29144 26142
rect 29178 26108 29202 26142
rect 29120 26084 29202 26108
rect 30138 26142 30220 26168
rect 30138 26108 30162 26142
rect 30196 26108 30220 26142
rect 30138 26084 30220 26108
rect 31156 26142 31238 26168
rect 31156 26108 31180 26142
rect 31214 26108 31238 26142
rect 31156 26084 31238 26108
rect 32174 26142 32256 26168
rect 32174 26108 32198 26142
rect 32232 26108 32256 26142
rect 32174 26084 32256 26108
rect 33192 26142 33274 26168
rect 33192 26108 33216 26142
rect 33250 26108 33274 26142
rect 33192 26084 33274 26108
rect 17922 24990 18004 25016
rect 17922 24956 17946 24990
rect 17980 24956 18004 24990
rect 17922 24932 18004 24956
rect 18940 24990 19022 25016
rect 18940 24956 18964 24990
rect 18998 24956 19022 24990
rect 18940 24932 19022 24956
rect 19958 24990 20040 25016
rect 19958 24956 19982 24990
rect 20016 24956 20040 24990
rect 19958 24932 20040 24956
rect 20976 24990 21058 25016
rect 20976 24956 21000 24990
rect 21034 24956 21058 24990
rect 20976 24932 21058 24956
rect 21994 24990 22076 25016
rect 21994 24956 22018 24990
rect 22052 24956 22076 24990
rect 21994 24932 22076 24956
rect 23012 24990 23094 25016
rect 23012 24956 23036 24990
rect 23070 24956 23094 24990
rect 23012 24932 23094 24956
rect 24030 24990 24112 25016
rect 24030 24956 24054 24990
rect 24088 24956 24112 24990
rect 24030 24932 24112 24956
rect 25048 24990 25130 25016
rect 25048 24956 25072 24990
rect 25106 24956 25130 24990
rect 25048 24932 25130 24956
rect 26066 24990 26148 25016
rect 26066 24956 26090 24990
rect 26124 24956 26148 24990
rect 26066 24932 26148 24956
rect 27084 24990 27166 25016
rect 27084 24956 27108 24990
rect 27142 24956 27166 24990
rect 27084 24932 27166 24956
rect 28102 24990 28184 25016
rect 28102 24956 28126 24990
rect 28160 24956 28184 24990
rect 28102 24932 28184 24956
rect 29120 24990 29202 25016
rect 29120 24956 29144 24990
rect 29178 24956 29202 24990
rect 29120 24932 29202 24956
rect 30138 24990 30220 25016
rect 30138 24956 30162 24990
rect 30196 24956 30220 24990
rect 30138 24932 30220 24956
rect 31156 24990 31238 25016
rect 31156 24956 31180 24990
rect 31214 24956 31238 24990
rect 31156 24932 31238 24956
rect 32174 24990 32256 25016
rect 32174 24956 32198 24990
rect 32232 24956 32256 24990
rect 32174 24932 32256 24956
rect 33192 24990 33274 25016
rect 33192 24956 33216 24990
rect 33250 24956 33274 24990
rect 33192 24932 33274 24956
rect 18940 23546 19022 23572
rect 18940 23512 18964 23546
rect 18998 23512 19022 23546
rect 18940 23488 19022 23512
rect 19958 23546 20040 23572
rect 19958 23512 19982 23546
rect 20016 23512 20040 23546
rect 19958 23488 20040 23512
rect 20976 23546 21058 23572
rect 20976 23512 21000 23546
rect 21034 23512 21058 23546
rect 20976 23488 21058 23512
rect 21994 23546 22076 23572
rect 21994 23512 22018 23546
rect 22052 23512 22076 23546
rect 21994 23488 22076 23512
rect 23012 23546 23094 23572
rect 23012 23512 23036 23546
rect 23070 23512 23094 23546
rect 23012 23488 23094 23512
rect 24030 23546 24112 23572
rect 24030 23512 24054 23546
rect 24088 23512 24112 23546
rect 24030 23488 24112 23512
rect 25048 23546 25130 23572
rect 25048 23512 25072 23546
rect 25106 23512 25130 23546
rect 25048 23488 25130 23512
rect 26066 23546 26148 23572
rect 26066 23512 26090 23546
rect 26124 23512 26148 23546
rect 26066 23488 26148 23512
rect 27084 23546 27166 23572
rect 27084 23512 27108 23546
rect 27142 23512 27166 23546
rect 27084 23488 27166 23512
rect 28102 23546 28184 23572
rect 28102 23512 28126 23546
rect 28160 23512 28184 23546
rect 28102 23488 28184 23512
rect 29120 23546 29202 23572
rect 29120 23512 29144 23546
rect 29178 23512 29202 23546
rect 29120 23488 29202 23512
rect 30138 23546 30220 23572
rect 30138 23512 30162 23546
rect 30196 23512 30220 23546
rect 30138 23488 30220 23512
rect 31156 23546 31238 23572
rect 31156 23512 31180 23546
rect 31214 23512 31238 23546
rect 31156 23488 31238 23512
rect 32174 23546 32256 23572
rect 32174 23512 32198 23546
rect 32232 23512 32256 23546
rect 32174 23488 32256 23512
rect 33192 23546 33274 23572
rect 33192 23512 33216 23546
rect 33250 23512 33274 23546
rect 33192 23488 33274 23512
rect 14666 22274 14748 22300
rect 14666 22240 14690 22274
rect 14724 22240 14748 22274
rect 14666 22216 14748 22240
rect 15684 22274 15766 22300
rect 15684 22240 15708 22274
rect 15742 22240 15766 22274
rect 15684 22216 15766 22240
rect 16702 22274 16784 22300
rect 16702 22240 16726 22274
rect 16760 22240 16784 22274
rect 16702 22216 16784 22240
rect 18940 22034 19022 22060
rect 18940 22000 18964 22034
rect 18998 22000 19022 22034
rect 18940 21976 19022 22000
rect 19958 22034 20040 22060
rect 19958 22000 19982 22034
rect 20016 22000 20040 22034
rect 19958 21976 20040 22000
rect 20976 22034 21058 22060
rect 20976 22000 21000 22034
rect 21034 22000 21058 22034
rect 20976 21976 21058 22000
rect 21994 22034 22076 22060
rect 21994 22000 22018 22034
rect 22052 22000 22076 22034
rect 21994 21976 22076 22000
rect 23012 22034 23094 22060
rect 23012 22000 23036 22034
rect 23070 22000 23094 22034
rect 23012 21976 23094 22000
rect 24030 22034 24112 22060
rect 24030 22000 24054 22034
rect 24088 22000 24112 22034
rect 24030 21976 24112 22000
rect 25048 22034 25130 22060
rect 25048 22000 25072 22034
rect 25106 22000 25130 22034
rect 25048 21976 25130 22000
rect 26066 22034 26148 22060
rect 26066 22000 26090 22034
rect 26124 22000 26148 22034
rect 26066 21976 26148 22000
rect 27084 22034 27166 22060
rect 27084 22000 27108 22034
rect 27142 22000 27166 22034
rect 27084 21976 27166 22000
rect 28102 22034 28184 22060
rect 28102 22000 28126 22034
rect 28160 22000 28184 22034
rect 28102 21976 28184 22000
rect 29120 22034 29202 22060
rect 29120 22000 29144 22034
rect 29178 22000 29202 22034
rect 29120 21976 29202 22000
rect 30138 22034 30220 22060
rect 30138 22000 30162 22034
rect 30196 22000 30220 22034
rect 30138 21976 30220 22000
rect 31156 22034 31238 22060
rect 31156 22000 31180 22034
rect 31214 22000 31238 22034
rect 31156 21976 31238 22000
rect 32174 22034 32256 22060
rect 32174 22000 32198 22034
rect 32232 22000 32256 22034
rect 32174 21976 32256 22000
rect 33192 22034 33274 22060
rect 33192 22000 33216 22034
rect 33250 22000 33274 22034
rect 33192 21976 33274 22000
rect 14624 21190 14706 21216
rect 14624 21156 14648 21190
rect 14682 21156 14706 21190
rect 14624 21132 14706 21156
rect 15642 21190 15724 21216
rect 15642 21156 15666 21190
rect 15700 21156 15724 21190
rect 15642 21132 15724 21156
rect 16660 21190 16742 21216
rect 16660 21156 16684 21190
rect 16718 21156 16742 21190
rect 16660 21132 16742 21156
rect 18898 20766 18980 20792
rect 18898 20732 18922 20766
rect 18956 20732 18980 20766
rect 18898 20708 18980 20732
rect 19916 20766 19998 20792
rect 19916 20732 19940 20766
rect 19974 20732 19998 20766
rect 19916 20708 19998 20732
rect 20934 20766 21016 20792
rect 20934 20732 20958 20766
rect 20992 20732 21016 20766
rect 20934 20708 21016 20732
rect 21952 20766 22034 20792
rect 21952 20732 21976 20766
rect 22010 20732 22034 20766
rect 21952 20708 22034 20732
rect 22970 20766 23052 20792
rect 22970 20732 22994 20766
rect 23028 20732 23052 20766
rect 22970 20708 23052 20732
rect 23988 20766 24070 20792
rect 23988 20732 24012 20766
rect 24046 20732 24070 20766
rect 23988 20708 24070 20732
rect 25006 20766 25088 20792
rect 25006 20732 25030 20766
rect 25064 20732 25088 20766
rect 25006 20708 25088 20732
rect 26024 20766 26106 20792
rect 26024 20732 26048 20766
rect 26082 20732 26106 20766
rect 26024 20708 26106 20732
rect 27042 20766 27124 20792
rect 27042 20732 27066 20766
rect 27100 20732 27124 20766
rect 27042 20708 27124 20732
rect 28060 20766 28142 20792
rect 28060 20732 28084 20766
rect 28118 20732 28142 20766
rect 28060 20708 28142 20732
rect 29078 20766 29160 20792
rect 29078 20732 29102 20766
rect 29136 20732 29160 20766
rect 29078 20708 29160 20732
rect 30096 20766 30178 20792
rect 30096 20732 30120 20766
rect 30154 20732 30178 20766
rect 30096 20708 30178 20732
rect 31114 20766 31196 20792
rect 31114 20732 31138 20766
rect 31172 20732 31196 20766
rect 31114 20708 31196 20732
rect 32132 20766 32214 20792
rect 32132 20732 32156 20766
rect 32190 20732 32214 20766
rect 32132 20708 32214 20732
rect 33150 20766 33232 20792
rect 33150 20732 33174 20766
rect 33208 20732 33232 20766
rect 33150 20708 33232 20732
rect 14596 20248 14678 20274
rect 14596 20214 14620 20248
rect 14654 20214 14678 20248
rect 14596 20190 14678 20214
rect 15614 20248 15696 20274
rect 15614 20214 15638 20248
rect 15672 20214 15696 20248
rect 15614 20190 15696 20214
rect 16632 20248 16714 20274
rect 16632 20214 16656 20248
rect 16690 20214 16714 20248
rect 16632 20190 16714 20214
rect 18898 19528 18980 19554
rect 18898 19494 18922 19528
rect 18956 19494 18980 19528
rect 18898 19470 18980 19494
rect 19916 19528 19998 19554
rect 19916 19494 19940 19528
rect 19974 19494 19998 19528
rect 19916 19470 19998 19494
rect 20934 19528 21016 19554
rect 20934 19494 20958 19528
rect 20992 19494 21016 19528
rect 20934 19470 21016 19494
rect 21952 19528 22034 19554
rect 21952 19494 21976 19528
rect 22010 19494 22034 19528
rect 21952 19470 22034 19494
rect 22970 19528 23052 19554
rect 22970 19494 22994 19528
rect 23028 19494 23052 19528
rect 22970 19470 23052 19494
rect 23988 19528 24070 19554
rect 23988 19494 24012 19528
rect 24046 19494 24070 19528
rect 23988 19470 24070 19494
rect 25006 19528 25088 19554
rect 25006 19494 25030 19528
rect 25064 19494 25088 19528
rect 25006 19470 25088 19494
rect 26024 19528 26106 19554
rect 26024 19494 26048 19528
rect 26082 19494 26106 19528
rect 26024 19470 26106 19494
rect 27042 19528 27124 19554
rect 27042 19494 27066 19528
rect 27100 19494 27124 19528
rect 27042 19470 27124 19494
rect 28060 19528 28142 19554
rect 28060 19494 28084 19528
rect 28118 19494 28142 19528
rect 28060 19470 28142 19494
rect 29078 19528 29160 19554
rect 29078 19494 29102 19528
rect 29136 19494 29160 19528
rect 29078 19470 29160 19494
rect 30096 19528 30178 19554
rect 30096 19494 30120 19528
rect 30154 19494 30178 19528
rect 30096 19470 30178 19494
rect 31114 19528 31196 19554
rect 31114 19494 31138 19528
rect 31172 19494 31196 19528
rect 31114 19470 31196 19494
rect 32132 19528 32214 19554
rect 32132 19494 32156 19528
rect 32190 19494 32214 19528
rect 32132 19470 32214 19494
rect 33150 19528 33232 19554
rect 33150 19494 33174 19528
rect 33208 19494 33232 19528
rect 33150 19470 33232 19494
rect 14596 19334 14678 19360
rect 14596 19300 14620 19334
rect 14654 19300 14678 19334
rect 14596 19276 14678 19300
rect 15614 19334 15696 19360
rect 15614 19300 15638 19334
rect 15672 19300 15696 19334
rect 15614 19276 15696 19300
rect 16632 19334 16714 19360
rect 16632 19300 16656 19334
rect 16690 19300 16714 19334
rect 16632 19276 16714 19300
rect 11328 17758 11428 17820
rect 65328 28162 65490 28262
rect 89610 28162 89772 28262
rect 65328 28100 65428 28162
rect 47264 25377 47360 25411
rect 48978 25377 49074 25411
rect 47264 25315 47298 25377
rect 49040 25315 49074 25377
rect 47264 24679 47298 24741
rect 49040 24679 49074 24741
rect 47264 24645 47360 24679
rect 48978 24645 49074 24679
rect 47264 23377 47360 23411
rect 48978 23377 49074 23411
rect 47264 23315 47298 23377
rect 49040 23315 49074 23377
rect 47264 22679 47298 22741
rect 49040 22679 49074 22741
rect 47264 22645 47360 22679
rect 48978 22645 49074 22679
rect 35672 17758 35772 17820
rect 11328 17658 11490 17758
rect 35610 17658 35772 17758
rect 89672 28100 89772 28162
rect 72940 26142 73022 26168
rect 72940 26108 72964 26142
rect 72998 26108 73022 26142
rect 72940 26084 73022 26108
rect 73958 26142 74040 26168
rect 73958 26108 73982 26142
rect 74016 26108 74040 26142
rect 73958 26084 74040 26108
rect 74976 26142 75058 26168
rect 74976 26108 75000 26142
rect 75034 26108 75058 26142
rect 74976 26084 75058 26108
rect 75994 26142 76076 26168
rect 75994 26108 76018 26142
rect 76052 26108 76076 26142
rect 75994 26084 76076 26108
rect 77012 26142 77094 26168
rect 77012 26108 77036 26142
rect 77070 26108 77094 26142
rect 77012 26084 77094 26108
rect 78030 26142 78112 26168
rect 78030 26108 78054 26142
rect 78088 26108 78112 26142
rect 78030 26084 78112 26108
rect 79048 26142 79130 26168
rect 79048 26108 79072 26142
rect 79106 26108 79130 26142
rect 79048 26084 79130 26108
rect 80066 26142 80148 26168
rect 80066 26108 80090 26142
rect 80124 26108 80148 26142
rect 80066 26084 80148 26108
rect 81084 26142 81166 26168
rect 81084 26108 81108 26142
rect 81142 26108 81166 26142
rect 81084 26084 81166 26108
rect 82102 26142 82184 26168
rect 82102 26108 82126 26142
rect 82160 26108 82184 26142
rect 82102 26084 82184 26108
rect 83120 26142 83202 26168
rect 83120 26108 83144 26142
rect 83178 26108 83202 26142
rect 83120 26084 83202 26108
rect 84138 26142 84220 26168
rect 84138 26108 84162 26142
rect 84196 26108 84220 26142
rect 84138 26084 84220 26108
rect 85156 26142 85238 26168
rect 85156 26108 85180 26142
rect 85214 26108 85238 26142
rect 85156 26084 85238 26108
rect 86174 26142 86256 26168
rect 86174 26108 86198 26142
rect 86232 26108 86256 26142
rect 86174 26084 86256 26108
rect 87192 26142 87274 26168
rect 87192 26108 87216 26142
rect 87250 26108 87274 26142
rect 87192 26084 87274 26108
rect 71922 24990 72004 25016
rect 71922 24956 71946 24990
rect 71980 24956 72004 24990
rect 71922 24932 72004 24956
rect 72940 24990 73022 25016
rect 72940 24956 72964 24990
rect 72998 24956 73022 24990
rect 72940 24932 73022 24956
rect 73958 24990 74040 25016
rect 73958 24956 73982 24990
rect 74016 24956 74040 24990
rect 73958 24932 74040 24956
rect 74976 24990 75058 25016
rect 74976 24956 75000 24990
rect 75034 24956 75058 24990
rect 74976 24932 75058 24956
rect 75994 24990 76076 25016
rect 75994 24956 76018 24990
rect 76052 24956 76076 24990
rect 75994 24932 76076 24956
rect 77012 24990 77094 25016
rect 77012 24956 77036 24990
rect 77070 24956 77094 24990
rect 77012 24932 77094 24956
rect 78030 24990 78112 25016
rect 78030 24956 78054 24990
rect 78088 24956 78112 24990
rect 78030 24932 78112 24956
rect 79048 24990 79130 25016
rect 79048 24956 79072 24990
rect 79106 24956 79130 24990
rect 79048 24932 79130 24956
rect 80066 24990 80148 25016
rect 80066 24956 80090 24990
rect 80124 24956 80148 24990
rect 80066 24932 80148 24956
rect 81084 24990 81166 25016
rect 81084 24956 81108 24990
rect 81142 24956 81166 24990
rect 81084 24932 81166 24956
rect 82102 24990 82184 25016
rect 82102 24956 82126 24990
rect 82160 24956 82184 24990
rect 82102 24932 82184 24956
rect 83120 24990 83202 25016
rect 83120 24956 83144 24990
rect 83178 24956 83202 24990
rect 83120 24932 83202 24956
rect 84138 24990 84220 25016
rect 84138 24956 84162 24990
rect 84196 24956 84220 24990
rect 84138 24932 84220 24956
rect 85156 24990 85238 25016
rect 85156 24956 85180 24990
rect 85214 24956 85238 24990
rect 85156 24932 85238 24956
rect 86174 24990 86256 25016
rect 86174 24956 86198 24990
rect 86232 24956 86256 24990
rect 86174 24932 86256 24956
rect 87192 24990 87274 25016
rect 87192 24956 87216 24990
rect 87250 24956 87274 24990
rect 87192 24932 87274 24956
rect 72940 23546 73022 23572
rect 72940 23512 72964 23546
rect 72998 23512 73022 23546
rect 72940 23488 73022 23512
rect 73958 23546 74040 23572
rect 73958 23512 73982 23546
rect 74016 23512 74040 23546
rect 73958 23488 74040 23512
rect 74976 23546 75058 23572
rect 74976 23512 75000 23546
rect 75034 23512 75058 23546
rect 74976 23488 75058 23512
rect 75994 23546 76076 23572
rect 75994 23512 76018 23546
rect 76052 23512 76076 23546
rect 75994 23488 76076 23512
rect 77012 23546 77094 23572
rect 77012 23512 77036 23546
rect 77070 23512 77094 23546
rect 77012 23488 77094 23512
rect 78030 23546 78112 23572
rect 78030 23512 78054 23546
rect 78088 23512 78112 23546
rect 78030 23488 78112 23512
rect 79048 23546 79130 23572
rect 79048 23512 79072 23546
rect 79106 23512 79130 23546
rect 79048 23488 79130 23512
rect 80066 23546 80148 23572
rect 80066 23512 80090 23546
rect 80124 23512 80148 23546
rect 80066 23488 80148 23512
rect 81084 23546 81166 23572
rect 81084 23512 81108 23546
rect 81142 23512 81166 23546
rect 81084 23488 81166 23512
rect 82102 23546 82184 23572
rect 82102 23512 82126 23546
rect 82160 23512 82184 23546
rect 82102 23488 82184 23512
rect 83120 23546 83202 23572
rect 83120 23512 83144 23546
rect 83178 23512 83202 23546
rect 83120 23488 83202 23512
rect 84138 23546 84220 23572
rect 84138 23512 84162 23546
rect 84196 23512 84220 23546
rect 84138 23488 84220 23512
rect 85156 23546 85238 23572
rect 85156 23512 85180 23546
rect 85214 23512 85238 23546
rect 85156 23488 85238 23512
rect 86174 23546 86256 23572
rect 86174 23512 86198 23546
rect 86232 23512 86256 23546
rect 86174 23488 86256 23512
rect 87192 23546 87274 23572
rect 87192 23512 87216 23546
rect 87250 23512 87274 23546
rect 87192 23488 87274 23512
rect 68666 22274 68748 22300
rect 68666 22240 68690 22274
rect 68724 22240 68748 22274
rect 68666 22216 68748 22240
rect 69684 22274 69766 22300
rect 69684 22240 69708 22274
rect 69742 22240 69766 22274
rect 69684 22216 69766 22240
rect 70702 22274 70784 22300
rect 70702 22240 70726 22274
rect 70760 22240 70784 22274
rect 70702 22216 70784 22240
rect 72940 22034 73022 22060
rect 72940 22000 72964 22034
rect 72998 22000 73022 22034
rect 72940 21976 73022 22000
rect 73958 22034 74040 22060
rect 73958 22000 73982 22034
rect 74016 22000 74040 22034
rect 73958 21976 74040 22000
rect 74976 22034 75058 22060
rect 74976 22000 75000 22034
rect 75034 22000 75058 22034
rect 74976 21976 75058 22000
rect 75994 22034 76076 22060
rect 75994 22000 76018 22034
rect 76052 22000 76076 22034
rect 75994 21976 76076 22000
rect 77012 22034 77094 22060
rect 77012 22000 77036 22034
rect 77070 22000 77094 22034
rect 77012 21976 77094 22000
rect 78030 22034 78112 22060
rect 78030 22000 78054 22034
rect 78088 22000 78112 22034
rect 78030 21976 78112 22000
rect 79048 22034 79130 22060
rect 79048 22000 79072 22034
rect 79106 22000 79130 22034
rect 79048 21976 79130 22000
rect 80066 22034 80148 22060
rect 80066 22000 80090 22034
rect 80124 22000 80148 22034
rect 80066 21976 80148 22000
rect 81084 22034 81166 22060
rect 81084 22000 81108 22034
rect 81142 22000 81166 22034
rect 81084 21976 81166 22000
rect 82102 22034 82184 22060
rect 82102 22000 82126 22034
rect 82160 22000 82184 22034
rect 82102 21976 82184 22000
rect 83120 22034 83202 22060
rect 83120 22000 83144 22034
rect 83178 22000 83202 22034
rect 83120 21976 83202 22000
rect 84138 22034 84220 22060
rect 84138 22000 84162 22034
rect 84196 22000 84220 22034
rect 84138 21976 84220 22000
rect 85156 22034 85238 22060
rect 85156 22000 85180 22034
rect 85214 22000 85238 22034
rect 85156 21976 85238 22000
rect 86174 22034 86256 22060
rect 86174 22000 86198 22034
rect 86232 22000 86256 22034
rect 86174 21976 86256 22000
rect 87192 22034 87274 22060
rect 87192 22000 87216 22034
rect 87250 22000 87274 22034
rect 87192 21976 87274 22000
rect 68624 21190 68706 21216
rect 68624 21156 68648 21190
rect 68682 21156 68706 21190
rect 68624 21132 68706 21156
rect 69642 21190 69724 21216
rect 69642 21156 69666 21190
rect 69700 21156 69724 21190
rect 69642 21132 69724 21156
rect 70660 21190 70742 21216
rect 70660 21156 70684 21190
rect 70718 21156 70742 21190
rect 70660 21132 70742 21156
rect 72898 20766 72980 20792
rect 72898 20732 72922 20766
rect 72956 20732 72980 20766
rect 72898 20708 72980 20732
rect 73916 20766 73998 20792
rect 73916 20732 73940 20766
rect 73974 20732 73998 20766
rect 73916 20708 73998 20732
rect 74934 20766 75016 20792
rect 74934 20732 74958 20766
rect 74992 20732 75016 20766
rect 74934 20708 75016 20732
rect 75952 20766 76034 20792
rect 75952 20732 75976 20766
rect 76010 20732 76034 20766
rect 75952 20708 76034 20732
rect 76970 20766 77052 20792
rect 76970 20732 76994 20766
rect 77028 20732 77052 20766
rect 76970 20708 77052 20732
rect 77988 20766 78070 20792
rect 77988 20732 78012 20766
rect 78046 20732 78070 20766
rect 77988 20708 78070 20732
rect 79006 20766 79088 20792
rect 79006 20732 79030 20766
rect 79064 20732 79088 20766
rect 79006 20708 79088 20732
rect 80024 20766 80106 20792
rect 80024 20732 80048 20766
rect 80082 20732 80106 20766
rect 80024 20708 80106 20732
rect 81042 20766 81124 20792
rect 81042 20732 81066 20766
rect 81100 20732 81124 20766
rect 81042 20708 81124 20732
rect 82060 20766 82142 20792
rect 82060 20732 82084 20766
rect 82118 20732 82142 20766
rect 82060 20708 82142 20732
rect 83078 20766 83160 20792
rect 83078 20732 83102 20766
rect 83136 20732 83160 20766
rect 83078 20708 83160 20732
rect 84096 20766 84178 20792
rect 84096 20732 84120 20766
rect 84154 20732 84178 20766
rect 84096 20708 84178 20732
rect 85114 20766 85196 20792
rect 85114 20732 85138 20766
rect 85172 20732 85196 20766
rect 85114 20708 85196 20732
rect 86132 20766 86214 20792
rect 86132 20732 86156 20766
rect 86190 20732 86214 20766
rect 86132 20708 86214 20732
rect 87150 20766 87232 20792
rect 87150 20732 87174 20766
rect 87208 20732 87232 20766
rect 87150 20708 87232 20732
rect 68596 20248 68678 20274
rect 68596 20214 68620 20248
rect 68654 20214 68678 20248
rect 68596 20190 68678 20214
rect 69614 20248 69696 20274
rect 69614 20214 69638 20248
rect 69672 20214 69696 20248
rect 69614 20190 69696 20214
rect 70632 20248 70714 20274
rect 70632 20214 70656 20248
rect 70690 20214 70714 20248
rect 70632 20190 70714 20214
rect 72898 19528 72980 19554
rect 72898 19494 72922 19528
rect 72956 19494 72980 19528
rect 72898 19470 72980 19494
rect 73916 19528 73998 19554
rect 73916 19494 73940 19528
rect 73974 19494 73998 19528
rect 73916 19470 73998 19494
rect 74934 19528 75016 19554
rect 74934 19494 74958 19528
rect 74992 19494 75016 19528
rect 74934 19470 75016 19494
rect 75952 19528 76034 19554
rect 75952 19494 75976 19528
rect 76010 19494 76034 19528
rect 75952 19470 76034 19494
rect 76970 19528 77052 19554
rect 76970 19494 76994 19528
rect 77028 19494 77052 19528
rect 76970 19470 77052 19494
rect 77988 19528 78070 19554
rect 77988 19494 78012 19528
rect 78046 19494 78070 19528
rect 77988 19470 78070 19494
rect 79006 19528 79088 19554
rect 79006 19494 79030 19528
rect 79064 19494 79088 19528
rect 79006 19470 79088 19494
rect 80024 19528 80106 19554
rect 80024 19494 80048 19528
rect 80082 19494 80106 19528
rect 80024 19470 80106 19494
rect 81042 19528 81124 19554
rect 81042 19494 81066 19528
rect 81100 19494 81124 19528
rect 81042 19470 81124 19494
rect 82060 19528 82142 19554
rect 82060 19494 82084 19528
rect 82118 19494 82142 19528
rect 82060 19470 82142 19494
rect 83078 19528 83160 19554
rect 83078 19494 83102 19528
rect 83136 19494 83160 19528
rect 83078 19470 83160 19494
rect 84096 19528 84178 19554
rect 84096 19494 84120 19528
rect 84154 19494 84178 19528
rect 84096 19470 84178 19494
rect 85114 19528 85196 19554
rect 85114 19494 85138 19528
rect 85172 19494 85196 19528
rect 85114 19470 85196 19494
rect 86132 19528 86214 19554
rect 86132 19494 86156 19528
rect 86190 19494 86214 19528
rect 86132 19470 86214 19494
rect 87150 19528 87232 19554
rect 87150 19494 87174 19528
rect 87208 19494 87232 19528
rect 87150 19470 87232 19494
rect 68596 19334 68678 19360
rect 68596 19300 68620 19334
rect 68654 19300 68678 19334
rect 68596 19276 68678 19300
rect 69614 19334 69696 19360
rect 69614 19300 69638 19334
rect 69672 19300 69696 19334
rect 69614 19276 69696 19300
rect 70632 19334 70714 19360
rect 70632 19300 70656 19334
rect 70690 19300 70714 19334
rect 70632 19276 70714 19300
rect 65328 17758 65428 17820
rect 89672 17758 89772 17820
rect 65328 17658 65490 17758
rect 89610 17658 89772 17758
rect -13094 16247 -12998 16281
rect -11380 16247 -11284 16281
rect -13094 16185 -13060 16247
rect -11318 16185 -11284 16247
rect -13094 15549 -13060 15611
rect -10494 16247 -10398 16281
rect -8780 16247 -8684 16281
rect -10494 16185 -10460 16247
rect -11318 15549 -11284 15611
rect -13094 15515 -12998 15549
rect -11380 15515 -11284 15549
rect -8718 16185 -8684 16247
rect -10494 15549 -10460 15611
rect -8718 15549 -8684 15611
rect -10494 15515 -10398 15549
rect -8780 15515 -8684 15549
rect 48690 8413 48786 8447
rect 50404 8413 50500 8447
rect 48690 8351 48724 8413
rect 50466 8351 50500 8413
rect 48690 7715 48724 7777
rect 50466 7715 50500 7777
rect 48690 7681 48786 7715
rect 50404 7681 50500 7715
rect 48690 6449 48786 6483
rect 50404 6449 50500 6483
rect 48690 6387 48724 6449
rect 50466 6387 50500 6449
rect 48690 5751 48724 5813
rect 50466 5751 50500 5813
rect 48690 5717 48786 5751
rect 50404 5717 50500 5751
rect 48690 4449 48786 4483
rect 50404 4449 50500 4483
rect 48690 4387 48724 4449
rect 50466 4387 50500 4449
rect 48690 3751 48724 3813
rect 50466 3751 50500 3813
rect 48690 3717 48786 3751
rect 50404 3717 50500 3751
rect 48690 2359 48786 2393
rect 50404 2359 50500 2393
rect 48690 2297 48724 2359
rect 50466 2297 50500 2359
rect 48690 1661 48724 1723
rect 50466 1661 50500 1723
rect 48690 1627 48786 1661
rect 50404 1627 50500 1661
<< psubdiffcont >>
rect 47360 24444 48978 24478
rect 47264 24026 47298 24382
rect 49040 24026 49074 24382
rect 47360 23930 48978 23964
rect 47360 22444 48978 22478
rect 47264 22026 47298 22382
rect 49040 22026 49074 22382
rect 47360 21930 48978 21964
rect -12998 15314 -11380 15348
rect -13094 14896 -13060 15252
rect -10398 15314 -8780 15348
rect -11318 14896 -11284 15252
rect -12998 14800 -11380 14834
rect -10494 14896 -10460 15252
rect -8718 14896 -8684 15252
rect -1210 15262 35710 15362
rect -10398 14800 -8780 14834
rect -1372 -520 -1272 15200
rect 2306 14284 2340 14318
rect 3324 14284 3358 14318
rect 4342 14284 4376 14318
rect 5360 14284 5394 14318
rect 6378 14284 6412 14318
rect 7396 14284 7430 14318
rect 8414 14284 8448 14318
rect 9432 14284 9466 14318
rect 10450 14284 10484 14318
rect 14040 13892 14074 13926
rect 15058 13892 15092 13926
rect 16076 13892 16110 13926
rect 17094 13892 17128 13926
rect 18112 13892 18146 13926
rect 19130 13892 19164 13926
rect 20148 13892 20182 13926
rect 21166 13892 21200 13926
rect 22184 13892 22218 13926
rect 23202 13892 23236 13926
rect 24220 13892 24254 13926
rect 25238 13892 25272 13926
rect 26256 13892 26290 13926
rect 27274 13892 27308 13926
rect 28292 13892 28326 13926
rect 29310 13892 29344 13926
rect 30328 13892 30362 13926
rect 31346 13892 31380 13926
rect 32364 13892 32398 13926
rect 33382 13892 33416 13926
rect 1768 13302 1802 13336
rect 2786 13302 2820 13336
rect 3804 13302 3838 13336
rect 4822 13302 4856 13336
rect 5840 13302 5874 13336
rect 6858 13302 6892 13336
rect 7876 13302 7910 13336
rect 8894 13302 8928 13336
rect 9912 13302 9946 13336
rect 10930 13302 10964 13336
rect 14028 12656 14062 12690
rect 15046 12656 15080 12690
rect 16064 12656 16098 12690
rect 17082 12656 17116 12690
rect 18100 12656 18134 12690
rect 19118 12656 19152 12690
rect 20136 12656 20170 12690
rect 21154 12656 21188 12690
rect 22172 12656 22206 12690
rect 23190 12656 23224 12690
rect 24208 12656 24242 12690
rect 25226 12656 25260 12690
rect 26244 12656 26278 12690
rect 27262 12656 27296 12690
rect 28280 12656 28314 12690
rect 29298 12656 29332 12690
rect 30316 12656 30350 12690
rect 31334 12656 31368 12690
rect 32352 12656 32386 12690
rect 33370 12656 33404 12690
rect 1768 12484 1802 12518
rect 2786 12484 2820 12518
rect 3804 12484 3838 12518
rect 4822 12484 4856 12518
rect 5840 12484 5874 12518
rect 6858 12484 6892 12518
rect 7876 12484 7910 12518
rect 8894 12484 8928 12518
rect 9912 12484 9946 12518
rect 10930 12484 10964 12518
rect 1768 11666 1802 11700
rect 2786 11666 2820 11700
rect 3804 11666 3838 11700
rect 4822 11666 4856 11700
rect 5840 11666 5874 11700
rect 6858 11666 6892 11700
rect 7876 11666 7910 11700
rect 8894 11666 8928 11700
rect 9912 11666 9946 11700
rect 10930 11666 10964 11700
rect 14040 11422 14074 11456
rect 15058 11422 15092 11456
rect 16076 11422 16110 11456
rect 17094 11422 17128 11456
rect 18112 11422 18146 11456
rect 19130 11422 19164 11456
rect 20148 11422 20182 11456
rect 21166 11422 21200 11456
rect 22184 11422 22218 11456
rect 23202 11422 23236 11456
rect 24220 11422 24254 11456
rect 25238 11422 25272 11456
rect 26256 11422 26290 11456
rect 27274 11422 27308 11456
rect 28292 11422 28326 11456
rect 29310 11422 29344 11456
rect 30328 11422 30362 11456
rect 31346 11422 31380 11456
rect 32364 11422 32398 11456
rect 33382 11422 33416 11456
rect 1768 10848 1802 10882
rect 2786 10848 2820 10882
rect 3804 10848 3838 10882
rect 4822 10848 4856 10882
rect 5840 10848 5874 10882
rect 6858 10848 6892 10882
rect 7876 10848 7910 10882
rect 8894 10848 8928 10882
rect 9912 10848 9946 10882
rect 10930 10848 10964 10882
rect 14040 10202 14074 10236
rect 15058 10202 15092 10236
rect 16076 10202 16110 10236
rect 17094 10202 17128 10236
rect 18112 10202 18146 10236
rect 19130 10202 19164 10236
rect 20148 10202 20182 10236
rect 21166 10202 21200 10236
rect 22184 10202 22218 10236
rect 23202 10202 23236 10236
rect 24220 10202 24254 10236
rect 25238 10202 25272 10236
rect 26256 10202 26290 10236
rect 27274 10202 27308 10236
rect 28292 10202 28326 10236
rect 29310 10202 29344 10236
rect 30328 10202 30362 10236
rect 31346 10202 31380 10236
rect 32364 10202 32398 10236
rect 33382 10202 33416 10236
rect 1768 10030 1802 10064
rect 2786 10030 2820 10064
rect 3804 10030 3838 10064
rect 4822 10030 4856 10064
rect 5840 10030 5874 10064
rect 6858 10030 6892 10064
rect 7876 10030 7910 10064
rect 8894 10030 8928 10064
rect 9912 10030 9946 10064
rect 10930 10030 10964 10064
rect 1768 9212 1802 9246
rect 2786 9212 2820 9246
rect 3804 9212 3838 9246
rect 4822 9212 4856 9246
rect 5840 9212 5874 9246
rect 6858 9212 6892 9246
rect 7876 9212 7910 9246
rect 8894 9212 8928 9246
rect 9912 9212 9946 9246
rect 10930 9212 10964 9246
rect 14054 8954 14088 8988
rect 15072 8954 15106 8988
rect 16090 8954 16124 8988
rect 17108 8954 17142 8988
rect 18126 8954 18160 8988
rect 19144 8954 19178 8988
rect 20162 8954 20196 8988
rect 21180 8954 21214 8988
rect 22198 8954 22232 8988
rect 23216 8954 23250 8988
rect 24234 8954 24268 8988
rect 25252 8954 25286 8988
rect 26270 8954 26304 8988
rect 27288 8954 27322 8988
rect 28306 8954 28340 8988
rect 29324 8954 29358 8988
rect 30342 8954 30376 8988
rect 31360 8954 31394 8988
rect 32378 8954 32412 8988
rect 33396 8954 33430 8988
rect 1768 8394 1802 8428
rect 2786 8394 2820 8428
rect 3804 8394 3838 8428
rect 4822 8394 4856 8428
rect 5840 8394 5874 8428
rect 6858 8394 6892 8428
rect 7876 8394 7910 8428
rect 8894 8394 8928 8428
rect 9912 8394 9946 8428
rect 10930 8394 10964 8428
rect 14040 7732 14074 7766
rect 15058 7732 15092 7766
rect 16076 7732 16110 7766
rect 17094 7732 17128 7766
rect 18112 7732 18146 7766
rect 19130 7732 19164 7766
rect 20148 7732 20182 7766
rect 21166 7732 21200 7766
rect 22184 7732 22218 7766
rect 23202 7732 23236 7766
rect 24220 7732 24254 7766
rect 25238 7732 25272 7766
rect 26256 7732 26290 7766
rect 27274 7732 27308 7766
rect 28292 7732 28326 7766
rect 29310 7732 29344 7766
rect 30328 7732 30362 7766
rect 31346 7732 31380 7766
rect 32364 7732 32398 7766
rect 33382 7732 33416 7766
rect 2278 7352 2312 7386
rect 3296 7352 3330 7386
rect 4314 7352 4348 7386
rect 5332 7352 5366 7386
rect 6350 7352 6384 7386
rect 7368 7352 7402 7386
rect 8386 7352 8420 7386
rect 9404 7352 9438 7386
rect 10422 7352 10456 7386
rect 14040 6484 14074 6518
rect 15058 6484 15092 6518
rect 16076 6484 16110 6518
rect 17094 6484 17128 6518
rect 18112 6484 18146 6518
rect 19130 6484 19164 6518
rect 20148 6484 20182 6518
rect 21166 6484 21200 6518
rect 22184 6484 22218 6518
rect 23202 6484 23236 6518
rect 24220 6484 24254 6518
rect 25238 6484 25272 6518
rect 26256 6484 26290 6518
rect 27274 6484 27308 6518
rect 28292 6484 28326 6518
rect 29310 6484 29344 6518
rect 30328 6484 30362 6518
rect 31346 6484 31380 6518
rect 32364 6484 32398 6518
rect 33382 6484 33416 6518
rect 8356 6376 8390 6410
rect 9374 6376 9408 6410
rect 10392 6376 10426 6410
rect 11410 6376 11444 6410
rect 14054 5264 14088 5298
rect 15072 5264 15106 5298
rect 16090 5264 16124 5298
rect 17108 5264 17142 5298
rect 18126 5264 18160 5298
rect 19144 5264 19178 5298
rect 20162 5264 20196 5298
rect 21180 5264 21214 5298
rect 22198 5264 22232 5298
rect 23216 5264 23250 5298
rect 24234 5264 24268 5298
rect 25252 5264 25286 5298
rect 26270 5264 26304 5298
rect 27288 5264 27322 5298
rect 28306 5264 28340 5298
rect 29324 5264 29358 5298
rect 30342 5264 30376 5298
rect 31360 5264 31394 5298
rect 32378 5264 32412 5298
rect 33396 5264 33430 5298
rect 2062 5032 2096 5066
rect 3080 5032 3114 5066
rect 4098 5032 4132 5066
rect 5116 5032 5150 5066
rect 6134 5032 6168 5066
rect 7152 5032 7186 5066
rect 8654 5088 8688 5122
rect 9672 5088 9706 5122
rect 10690 5088 10724 5122
rect 11708 5088 11742 5122
rect 14054 4016 14088 4050
rect 15072 4016 15106 4050
rect 16090 4016 16124 4050
rect 17108 4016 17142 4050
rect 18126 4016 18160 4050
rect 19144 4016 19178 4050
rect 20162 4016 20196 4050
rect 21180 4016 21214 4050
rect 22198 4016 22232 4050
rect 23216 4016 23250 4050
rect 24234 4016 24268 4050
rect 25252 4016 25286 4050
rect 26270 4016 26304 4050
rect 27288 4016 27322 4050
rect 28306 4016 28340 4050
rect 29324 4016 29358 4050
rect 30342 4016 30376 4050
rect 31360 4016 31394 4050
rect 32378 4016 32412 4050
rect 33396 4016 33430 4050
rect 2076 3906 2110 3940
rect 3094 3906 3128 3940
rect 4112 3906 4146 3940
rect 5130 3906 5164 3940
rect 6148 3906 6182 3940
rect 7166 3906 7200 3940
rect 8614 3894 8648 3928
rect 9632 3894 9666 3928
rect 10650 3894 10684 3928
rect 11668 3894 11702 3928
rect 2050 2780 2084 2814
rect 3068 2780 3102 2814
rect 4086 2780 4120 2814
rect 5104 2780 5138 2814
rect 6122 2780 6156 2814
rect 7140 2780 7174 2814
rect 8614 2780 8648 2814
rect 9632 2780 9666 2814
rect 10650 2780 10684 2814
rect 11668 2780 11702 2814
rect 14040 2794 14074 2828
rect 15058 2794 15092 2828
rect 16076 2794 16110 2828
rect 17094 2794 17128 2828
rect 18112 2794 18146 2828
rect 19130 2794 19164 2828
rect 20148 2794 20182 2828
rect 21166 2794 21200 2828
rect 22184 2794 22218 2828
rect 23202 2794 23236 2828
rect 24220 2794 24254 2828
rect 25238 2794 25272 2828
rect 26256 2794 26290 2828
rect 27274 2794 27308 2828
rect 28292 2794 28326 2828
rect 29310 2794 29344 2828
rect 30328 2794 30362 2828
rect 31346 2794 31380 2828
rect 32364 2794 32398 2828
rect 33382 2794 33416 2828
rect 2076 1682 2110 1716
rect 3094 1682 3128 1716
rect 4112 1682 4146 1716
rect 5130 1682 5164 1716
rect 6148 1682 6182 1716
rect 7166 1682 7200 1716
rect 8668 1668 8702 1702
rect 9686 1668 9720 1702
rect 10704 1668 10738 1702
rect 11722 1668 11756 1702
rect 14040 1574 14074 1608
rect 15058 1574 15092 1608
rect 16076 1574 16110 1608
rect 17094 1574 17128 1608
rect 18112 1574 18146 1608
rect 19130 1574 19164 1608
rect 20148 1574 20182 1608
rect 21166 1574 21200 1608
rect 22184 1574 22218 1608
rect 23202 1574 23236 1608
rect 24220 1574 24254 1608
rect 25238 1574 25272 1608
rect 26256 1574 26290 1608
rect 27274 1574 27308 1608
rect 28292 1574 28326 1608
rect 29310 1574 29344 1608
rect 30328 1574 30362 1608
rect 31346 1574 31380 1608
rect 32364 1574 32398 1608
rect 33382 1574 33416 1608
rect 2050 488 2084 522
rect 3068 488 3102 522
rect 4086 488 4120 522
rect 5104 488 5138 522
rect 6122 488 6156 522
rect 7140 488 7174 522
rect 8642 434 8676 468
rect 9660 434 9694 468
rect 10678 434 10712 468
rect 11696 434 11730 468
rect 35772 -520 35872 15200
rect 52790 15262 89710 15362
rect 48786 7480 50404 7514
rect 48690 7062 48724 7418
rect 50466 7062 50500 7418
rect 48786 6966 50404 7000
rect 48786 5516 50404 5550
rect 48690 5098 48724 5454
rect 50466 5098 50500 5454
rect 48786 5002 50404 5036
rect 48786 3516 50404 3550
rect 48690 3098 48724 3454
rect 50466 3098 50500 3454
rect 48786 3002 50404 3036
rect 48786 1426 50404 1460
rect 48690 1008 48724 1364
rect 50466 1008 50500 1364
rect 48786 912 50404 946
rect -1210 -682 35710 -582
rect 52628 -520 52728 15200
rect 56306 14284 56340 14318
rect 57324 14284 57358 14318
rect 58342 14284 58376 14318
rect 59360 14284 59394 14318
rect 60378 14284 60412 14318
rect 61396 14284 61430 14318
rect 62414 14284 62448 14318
rect 63432 14284 63466 14318
rect 64450 14284 64484 14318
rect 68040 13892 68074 13926
rect 69058 13892 69092 13926
rect 70076 13892 70110 13926
rect 71094 13892 71128 13926
rect 72112 13892 72146 13926
rect 73130 13892 73164 13926
rect 74148 13892 74182 13926
rect 75166 13892 75200 13926
rect 76184 13892 76218 13926
rect 77202 13892 77236 13926
rect 78220 13892 78254 13926
rect 79238 13892 79272 13926
rect 80256 13892 80290 13926
rect 81274 13892 81308 13926
rect 82292 13892 82326 13926
rect 83310 13892 83344 13926
rect 84328 13892 84362 13926
rect 85346 13892 85380 13926
rect 86364 13892 86398 13926
rect 87382 13892 87416 13926
rect 55768 13302 55802 13336
rect 56786 13302 56820 13336
rect 57804 13302 57838 13336
rect 58822 13302 58856 13336
rect 59840 13302 59874 13336
rect 60858 13302 60892 13336
rect 61876 13302 61910 13336
rect 62894 13302 62928 13336
rect 63912 13302 63946 13336
rect 64930 13302 64964 13336
rect 68028 12656 68062 12690
rect 69046 12656 69080 12690
rect 70064 12656 70098 12690
rect 71082 12656 71116 12690
rect 72100 12656 72134 12690
rect 73118 12656 73152 12690
rect 74136 12656 74170 12690
rect 75154 12656 75188 12690
rect 76172 12656 76206 12690
rect 77190 12656 77224 12690
rect 78208 12656 78242 12690
rect 79226 12656 79260 12690
rect 80244 12656 80278 12690
rect 81262 12656 81296 12690
rect 82280 12656 82314 12690
rect 83298 12656 83332 12690
rect 84316 12656 84350 12690
rect 85334 12656 85368 12690
rect 86352 12656 86386 12690
rect 87370 12656 87404 12690
rect 55768 12484 55802 12518
rect 56786 12484 56820 12518
rect 57804 12484 57838 12518
rect 58822 12484 58856 12518
rect 59840 12484 59874 12518
rect 60858 12484 60892 12518
rect 61876 12484 61910 12518
rect 62894 12484 62928 12518
rect 63912 12484 63946 12518
rect 64930 12484 64964 12518
rect 55768 11666 55802 11700
rect 56786 11666 56820 11700
rect 57804 11666 57838 11700
rect 58822 11666 58856 11700
rect 59840 11666 59874 11700
rect 60858 11666 60892 11700
rect 61876 11666 61910 11700
rect 62894 11666 62928 11700
rect 63912 11666 63946 11700
rect 64930 11666 64964 11700
rect 68040 11422 68074 11456
rect 69058 11422 69092 11456
rect 70076 11422 70110 11456
rect 71094 11422 71128 11456
rect 72112 11422 72146 11456
rect 73130 11422 73164 11456
rect 74148 11422 74182 11456
rect 75166 11422 75200 11456
rect 76184 11422 76218 11456
rect 77202 11422 77236 11456
rect 78220 11422 78254 11456
rect 79238 11422 79272 11456
rect 80256 11422 80290 11456
rect 81274 11422 81308 11456
rect 82292 11422 82326 11456
rect 83310 11422 83344 11456
rect 84328 11422 84362 11456
rect 85346 11422 85380 11456
rect 86364 11422 86398 11456
rect 87382 11422 87416 11456
rect 55768 10848 55802 10882
rect 56786 10848 56820 10882
rect 57804 10848 57838 10882
rect 58822 10848 58856 10882
rect 59840 10848 59874 10882
rect 60858 10848 60892 10882
rect 61876 10848 61910 10882
rect 62894 10848 62928 10882
rect 63912 10848 63946 10882
rect 64930 10848 64964 10882
rect 68040 10202 68074 10236
rect 69058 10202 69092 10236
rect 70076 10202 70110 10236
rect 71094 10202 71128 10236
rect 72112 10202 72146 10236
rect 73130 10202 73164 10236
rect 74148 10202 74182 10236
rect 75166 10202 75200 10236
rect 76184 10202 76218 10236
rect 77202 10202 77236 10236
rect 78220 10202 78254 10236
rect 79238 10202 79272 10236
rect 80256 10202 80290 10236
rect 81274 10202 81308 10236
rect 82292 10202 82326 10236
rect 83310 10202 83344 10236
rect 84328 10202 84362 10236
rect 85346 10202 85380 10236
rect 86364 10202 86398 10236
rect 87382 10202 87416 10236
rect 55768 10030 55802 10064
rect 56786 10030 56820 10064
rect 57804 10030 57838 10064
rect 58822 10030 58856 10064
rect 59840 10030 59874 10064
rect 60858 10030 60892 10064
rect 61876 10030 61910 10064
rect 62894 10030 62928 10064
rect 63912 10030 63946 10064
rect 64930 10030 64964 10064
rect 55768 9212 55802 9246
rect 56786 9212 56820 9246
rect 57804 9212 57838 9246
rect 58822 9212 58856 9246
rect 59840 9212 59874 9246
rect 60858 9212 60892 9246
rect 61876 9212 61910 9246
rect 62894 9212 62928 9246
rect 63912 9212 63946 9246
rect 64930 9212 64964 9246
rect 68054 8954 68088 8988
rect 69072 8954 69106 8988
rect 70090 8954 70124 8988
rect 71108 8954 71142 8988
rect 72126 8954 72160 8988
rect 73144 8954 73178 8988
rect 74162 8954 74196 8988
rect 75180 8954 75214 8988
rect 76198 8954 76232 8988
rect 77216 8954 77250 8988
rect 78234 8954 78268 8988
rect 79252 8954 79286 8988
rect 80270 8954 80304 8988
rect 81288 8954 81322 8988
rect 82306 8954 82340 8988
rect 83324 8954 83358 8988
rect 84342 8954 84376 8988
rect 85360 8954 85394 8988
rect 86378 8954 86412 8988
rect 87396 8954 87430 8988
rect 55768 8394 55802 8428
rect 56786 8394 56820 8428
rect 57804 8394 57838 8428
rect 58822 8394 58856 8428
rect 59840 8394 59874 8428
rect 60858 8394 60892 8428
rect 61876 8394 61910 8428
rect 62894 8394 62928 8428
rect 63912 8394 63946 8428
rect 64930 8394 64964 8428
rect 68040 7732 68074 7766
rect 69058 7732 69092 7766
rect 70076 7732 70110 7766
rect 71094 7732 71128 7766
rect 72112 7732 72146 7766
rect 73130 7732 73164 7766
rect 74148 7732 74182 7766
rect 75166 7732 75200 7766
rect 76184 7732 76218 7766
rect 77202 7732 77236 7766
rect 78220 7732 78254 7766
rect 79238 7732 79272 7766
rect 80256 7732 80290 7766
rect 81274 7732 81308 7766
rect 82292 7732 82326 7766
rect 83310 7732 83344 7766
rect 84328 7732 84362 7766
rect 85346 7732 85380 7766
rect 86364 7732 86398 7766
rect 87382 7732 87416 7766
rect 56278 7352 56312 7386
rect 57296 7352 57330 7386
rect 58314 7352 58348 7386
rect 59332 7352 59366 7386
rect 60350 7352 60384 7386
rect 61368 7352 61402 7386
rect 62386 7352 62420 7386
rect 63404 7352 63438 7386
rect 64422 7352 64456 7386
rect 68040 6484 68074 6518
rect 69058 6484 69092 6518
rect 70076 6484 70110 6518
rect 71094 6484 71128 6518
rect 72112 6484 72146 6518
rect 73130 6484 73164 6518
rect 74148 6484 74182 6518
rect 75166 6484 75200 6518
rect 76184 6484 76218 6518
rect 77202 6484 77236 6518
rect 78220 6484 78254 6518
rect 79238 6484 79272 6518
rect 80256 6484 80290 6518
rect 81274 6484 81308 6518
rect 82292 6484 82326 6518
rect 83310 6484 83344 6518
rect 84328 6484 84362 6518
rect 85346 6484 85380 6518
rect 86364 6484 86398 6518
rect 87382 6484 87416 6518
rect 62356 6376 62390 6410
rect 63374 6376 63408 6410
rect 64392 6376 64426 6410
rect 65410 6376 65444 6410
rect 68054 5264 68088 5298
rect 69072 5264 69106 5298
rect 70090 5264 70124 5298
rect 71108 5264 71142 5298
rect 72126 5264 72160 5298
rect 73144 5264 73178 5298
rect 74162 5264 74196 5298
rect 75180 5264 75214 5298
rect 76198 5264 76232 5298
rect 77216 5264 77250 5298
rect 78234 5264 78268 5298
rect 79252 5264 79286 5298
rect 80270 5264 80304 5298
rect 81288 5264 81322 5298
rect 82306 5264 82340 5298
rect 83324 5264 83358 5298
rect 84342 5264 84376 5298
rect 85360 5264 85394 5298
rect 86378 5264 86412 5298
rect 87396 5264 87430 5298
rect 56062 5032 56096 5066
rect 57080 5032 57114 5066
rect 58098 5032 58132 5066
rect 59116 5032 59150 5066
rect 60134 5032 60168 5066
rect 61152 5032 61186 5066
rect 62654 5088 62688 5122
rect 63672 5088 63706 5122
rect 64690 5088 64724 5122
rect 65708 5088 65742 5122
rect 68054 4016 68088 4050
rect 69072 4016 69106 4050
rect 70090 4016 70124 4050
rect 71108 4016 71142 4050
rect 72126 4016 72160 4050
rect 73144 4016 73178 4050
rect 74162 4016 74196 4050
rect 75180 4016 75214 4050
rect 76198 4016 76232 4050
rect 77216 4016 77250 4050
rect 78234 4016 78268 4050
rect 79252 4016 79286 4050
rect 80270 4016 80304 4050
rect 81288 4016 81322 4050
rect 82306 4016 82340 4050
rect 83324 4016 83358 4050
rect 84342 4016 84376 4050
rect 85360 4016 85394 4050
rect 86378 4016 86412 4050
rect 87396 4016 87430 4050
rect 56076 3906 56110 3940
rect 57094 3906 57128 3940
rect 58112 3906 58146 3940
rect 59130 3906 59164 3940
rect 60148 3906 60182 3940
rect 61166 3906 61200 3940
rect 62614 3894 62648 3928
rect 63632 3894 63666 3928
rect 64650 3894 64684 3928
rect 65668 3894 65702 3928
rect 56050 2780 56084 2814
rect 57068 2780 57102 2814
rect 58086 2780 58120 2814
rect 59104 2780 59138 2814
rect 60122 2780 60156 2814
rect 61140 2780 61174 2814
rect 62614 2780 62648 2814
rect 63632 2780 63666 2814
rect 64650 2780 64684 2814
rect 65668 2780 65702 2814
rect 68040 2794 68074 2828
rect 69058 2794 69092 2828
rect 70076 2794 70110 2828
rect 71094 2794 71128 2828
rect 72112 2794 72146 2828
rect 73130 2794 73164 2828
rect 74148 2794 74182 2828
rect 75166 2794 75200 2828
rect 76184 2794 76218 2828
rect 77202 2794 77236 2828
rect 78220 2794 78254 2828
rect 79238 2794 79272 2828
rect 80256 2794 80290 2828
rect 81274 2794 81308 2828
rect 82292 2794 82326 2828
rect 83310 2794 83344 2828
rect 84328 2794 84362 2828
rect 85346 2794 85380 2828
rect 86364 2794 86398 2828
rect 87382 2794 87416 2828
rect 56076 1682 56110 1716
rect 57094 1682 57128 1716
rect 58112 1682 58146 1716
rect 59130 1682 59164 1716
rect 60148 1682 60182 1716
rect 61166 1682 61200 1716
rect 62668 1668 62702 1702
rect 63686 1668 63720 1702
rect 64704 1668 64738 1702
rect 65722 1668 65756 1702
rect 68040 1574 68074 1608
rect 69058 1574 69092 1608
rect 70076 1574 70110 1608
rect 71094 1574 71128 1608
rect 72112 1574 72146 1608
rect 73130 1574 73164 1608
rect 74148 1574 74182 1608
rect 75166 1574 75200 1608
rect 76184 1574 76218 1608
rect 77202 1574 77236 1608
rect 78220 1574 78254 1608
rect 79238 1574 79272 1608
rect 80256 1574 80290 1608
rect 81274 1574 81308 1608
rect 82292 1574 82326 1608
rect 83310 1574 83344 1608
rect 84328 1574 84362 1608
rect 85346 1574 85380 1608
rect 86364 1574 86398 1608
rect 87382 1574 87416 1608
rect 56050 488 56084 522
rect 57068 488 57102 522
rect 58086 488 58120 522
rect 59104 488 59138 522
rect 60122 488 60156 522
rect 61140 488 61174 522
rect 62642 434 62676 468
rect 63660 434 63694 468
rect 64678 434 64712 468
rect 65696 434 65730 468
rect 89772 -520 89872 15200
rect 52790 -682 89710 -582
<< nsubdiffcont >>
rect 11490 28162 35610 28262
rect 11328 17820 11428 28100
rect 18964 26108 18998 26142
rect 19982 26108 20016 26142
rect 21000 26108 21034 26142
rect 22018 26108 22052 26142
rect 23036 26108 23070 26142
rect 24054 26108 24088 26142
rect 25072 26108 25106 26142
rect 26090 26108 26124 26142
rect 27108 26108 27142 26142
rect 28126 26108 28160 26142
rect 29144 26108 29178 26142
rect 30162 26108 30196 26142
rect 31180 26108 31214 26142
rect 32198 26108 32232 26142
rect 33216 26108 33250 26142
rect 17946 24956 17980 24990
rect 18964 24956 18998 24990
rect 19982 24956 20016 24990
rect 21000 24956 21034 24990
rect 22018 24956 22052 24990
rect 23036 24956 23070 24990
rect 24054 24956 24088 24990
rect 25072 24956 25106 24990
rect 26090 24956 26124 24990
rect 27108 24956 27142 24990
rect 28126 24956 28160 24990
rect 29144 24956 29178 24990
rect 30162 24956 30196 24990
rect 31180 24956 31214 24990
rect 32198 24956 32232 24990
rect 33216 24956 33250 24990
rect 18964 23512 18998 23546
rect 19982 23512 20016 23546
rect 21000 23512 21034 23546
rect 22018 23512 22052 23546
rect 23036 23512 23070 23546
rect 24054 23512 24088 23546
rect 25072 23512 25106 23546
rect 26090 23512 26124 23546
rect 27108 23512 27142 23546
rect 28126 23512 28160 23546
rect 29144 23512 29178 23546
rect 30162 23512 30196 23546
rect 31180 23512 31214 23546
rect 32198 23512 32232 23546
rect 33216 23512 33250 23546
rect 14690 22240 14724 22274
rect 15708 22240 15742 22274
rect 16726 22240 16760 22274
rect 18964 22000 18998 22034
rect 19982 22000 20016 22034
rect 21000 22000 21034 22034
rect 22018 22000 22052 22034
rect 23036 22000 23070 22034
rect 24054 22000 24088 22034
rect 25072 22000 25106 22034
rect 26090 22000 26124 22034
rect 27108 22000 27142 22034
rect 28126 22000 28160 22034
rect 29144 22000 29178 22034
rect 30162 22000 30196 22034
rect 31180 22000 31214 22034
rect 32198 22000 32232 22034
rect 33216 22000 33250 22034
rect 14648 21156 14682 21190
rect 15666 21156 15700 21190
rect 16684 21156 16718 21190
rect 18922 20732 18956 20766
rect 19940 20732 19974 20766
rect 20958 20732 20992 20766
rect 21976 20732 22010 20766
rect 22994 20732 23028 20766
rect 24012 20732 24046 20766
rect 25030 20732 25064 20766
rect 26048 20732 26082 20766
rect 27066 20732 27100 20766
rect 28084 20732 28118 20766
rect 29102 20732 29136 20766
rect 30120 20732 30154 20766
rect 31138 20732 31172 20766
rect 32156 20732 32190 20766
rect 33174 20732 33208 20766
rect 14620 20214 14654 20248
rect 15638 20214 15672 20248
rect 16656 20214 16690 20248
rect 18922 19494 18956 19528
rect 19940 19494 19974 19528
rect 20958 19494 20992 19528
rect 21976 19494 22010 19528
rect 22994 19494 23028 19528
rect 24012 19494 24046 19528
rect 25030 19494 25064 19528
rect 26048 19494 26082 19528
rect 27066 19494 27100 19528
rect 28084 19494 28118 19528
rect 29102 19494 29136 19528
rect 30120 19494 30154 19528
rect 31138 19494 31172 19528
rect 32156 19494 32190 19528
rect 33174 19494 33208 19528
rect 14620 19300 14654 19334
rect 15638 19300 15672 19334
rect 16656 19300 16690 19334
rect 35672 17820 35772 28100
rect 65490 28162 89610 28262
rect 47360 25377 48978 25411
rect 47264 24741 47298 25315
rect 49040 24741 49074 25315
rect 47360 24645 48978 24679
rect 47360 23377 48978 23411
rect 47264 22741 47298 23315
rect 49040 22741 49074 23315
rect 47360 22645 48978 22679
rect 11490 17658 35610 17758
rect 65328 17820 65428 28100
rect 72964 26108 72998 26142
rect 73982 26108 74016 26142
rect 75000 26108 75034 26142
rect 76018 26108 76052 26142
rect 77036 26108 77070 26142
rect 78054 26108 78088 26142
rect 79072 26108 79106 26142
rect 80090 26108 80124 26142
rect 81108 26108 81142 26142
rect 82126 26108 82160 26142
rect 83144 26108 83178 26142
rect 84162 26108 84196 26142
rect 85180 26108 85214 26142
rect 86198 26108 86232 26142
rect 87216 26108 87250 26142
rect 71946 24956 71980 24990
rect 72964 24956 72998 24990
rect 73982 24956 74016 24990
rect 75000 24956 75034 24990
rect 76018 24956 76052 24990
rect 77036 24956 77070 24990
rect 78054 24956 78088 24990
rect 79072 24956 79106 24990
rect 80090 24956 80124 24990
rect 81108 24956 81142 24990
rect 82126 24956 82160 24990
rect 83144 24956 83178 24990
rect 84162 24956 84196 24990
rect 85180 24956 85214 24990
rect 86198 24956 86232 24990
rect 87216 24956 87250 24990
rect 72964 23512 72998 23546
rect 73982 23512 74016 23546
rect 75000 23512 75034 23546
rect 76018 23512 76052 23546
rect 77036 23512 77070 23546
rect 78054 23512 78088 23546
rect 79072 23512 79106 23546
rect 80090 23512 80124 23546
rect 81108 23512 81142 23546
rect 82126 23512 82160 23546
rect 83144 23512 83178 23546
rect 84162 23512 84196 23546
rect 85180 23512 85214 23546
rect 86198 23512 86232 23546
rect 87216 23512 87250 23546
rect 68690 22240 68724 22274
rect 69708 22240 69742 22274
rect 70726 22240 70760 22274
rect 72964 22000 72998 22034
rect 73982 22000 74016 22034
rect 75000 22000 75034 22034
rect 76018 22000 76052 22034
rect 77036 22000 77070 22034
rect 78054 22000 78088 22034
rect 79072 22000 79106 22034
rect 80090 22000 80124 22034
rect 81108 22000 81142 22034
rect 82126 22000 82160 22034
rect 83144 22000 83178 22034
rect 84162 22000 84196 22034
rect 85180 22000 85214 22034
rect 86198 22000 86232 22034
rect 87216 22000 87250 22034
rect 68648 21156 68682 21190
rect 69666 21156 69700 21190
rect 70684 21156 70718 21190
rect 72922 20732 72956 20766
rect 73940 20732 73974 20766
rect 74958 20732 74992 20766
rect 75976 20732 76010 20766
rect 76994 20732 77028 20766
rect 78012 20732 78046 20766
rect 79030 20732 79064 20766
rect 80048 20732 80082 20766
rect 81066 20732 81100 20766
rect 82084 20732 82118 20766
rect 83102 20732 83136 20766
rect 84120 20732 84154 20766
rect 85138 20732 85172 20766
rect 86156 20732 86190 20766
rect 87174 20732 87208 20766
rect 68620 20214 68654 20248
rect 69638 20214 69672 20248
rect 70656 20214 70690 20248
rect 72922 19494 72956 19528
rect 73940 19494 73974 19528
rect 74958 19494 74992 19528
rect 75976 19494 76010 19528
rect 76994 19494 77028 19528
rect 78012 19494 78046 19528
rect 79030 19494 79064 19528
rect 80048 19494 80082 19528
rect 81066 19494 81100 19528
rect 82084 19494 82118 19528
rect 83102 19494 83136 19528
rect 84120 19494 84154 19528
rect 85138 19494 85172 19528
rect 86156 19494 86190 19528
rect 87174 19494 87208 19528
rect 68620 19300 68654 19334
rect 69638 19300 69672 19334
rect 70656 19300 70690 19334
rect 89672 17820 89772 28100
rect 65490 17658 89610 17758
rect -12998 16247 -11380 16281
rect -13094 15611 -13060 16185
rect -11318 15611 -11284 16185
rect -10398 16247 -8780 16281
rect -12998 15515 -11380 15549
rect -10494 15611 -10460 16185
rect -8718 15611 -8684 16185
rect -10398 15515 -8780 15549
rect 48786 8413 50404 8447
rect 48690 7777 48724 8351
rect 50466 7777 50500 8351
rect 48786 7681 50404 7715
rect 48786 6449 50404 6483
rect 48690 5813 48724 6387
rect 50466 5813 50500 6387
rect 48786 5717 50404 5751
rect 48786 4449 50404 4483
rect 48690 3813 48724 4387
rect 50466 3813 50500 4387
rect 48786 3717 50404 3751
rect 48786 2359 50404 2393
rect 48690 1723 48724 2297
rect 50466 1723 50500 2297
rect 48786 1627 50404 1661
<< poly >>
rect 17670 27061 18258 27077
rect 17670 27044 17686 27061
rect 17484 27027 17686 27044
rect 18242 27044 18258 27061
rect 18688 27061 19276 27077
rect 18688 27044 18704 27061
rect 18242 27027 18444 27044
rect 17484 26980 18444 27027
rect 18502 27027 18704 27044
rect 19260 27044 19276 27061
rect 19706 27061 20294 27077
rect 19706 27044 19722 27061
rect 19260 27027 19462 27044
rect 18502 26980 19462 27027
rect 19520 27027 19722 27044
rect 20278 27044 20294 27061
rect 20724 27061 21312 27077
rect 20724 27044 20740 27061
rect 20278 27027 20480 27044
rect 19520 26980 20480 27027
rect 20538 27027 20740 27044
rect 21296 27044 21312 27061
rect 21742 27061 22330 27077
rect 21742 27044 21758 27061
rect 21296 27027 21498 27044
rect 20538 26980 21498 27027
rect 21556 27027 21758 27044
rect 22314 27044 22330 27061
rect 22760 27061 23348 27077
rect 22760 27044 22776 27061
rect 22314 27027 22516 27044
rect 21556 26980 22516 27027
rect 22574 27027 22776 27044
rect 23332 27044 23348 27061
rect 23778 27061 24366 27077
rect 23778 27044 23794 27061
rect 23332 27027 23534 27044
rect 22574 26980 23534 27027
rect 23592 27027 23794 27044
rect 24350 27044 24366 27061
rect 24796 27061 25384 27077
rect 24796 27044 24812 27061
rect 24350 27027 24552 27044
rect 23592 26980 24552 27027
rect 24610 27027 24812 27044
rect 25368 27044 25384 27061
rect 25814 27061 26402 27077
rect 25814 27044 25830 27061
rect 25368 27027 25570 27044
rect 24610 26980 25570 27027
rect 25628 27027 25830 27044
rect 26386 27044 26402 27061
rect 26832 27061 27420 27077
rect 26832 27044 26848 27061
rect 26386 27027 26588 27044
rect 25628 26980 26588 27027
rect 26646 27027 26848 27044
rect 27404 27044 27420 27061
rect 27850 27061 28438 27077
rect 27850 27044 27866 27061
rect 27404 27027 27606 27044
rect 26646 26980 27606 27027
rect 27664 27027 27866 27044
rect 28422 27044 28438 27061
rect 28868 27061 29456 27077
rect 28868 27044 28884 27061
rect 28422 27027 28624 27044
rect 27664 26980 28624 27027
rect 28682 27027 28884 27044
rect 29440 27044 29456 27061
rect 29886 27061 30474 27077
rect 29886 27044 29902 27061
rect 29440 27027 29642 27044
rect 28682 26980 29642 27027
rect 29700 27027 29902 27044
rect 30458 27044 30474 27061
rect 30904 27061 31492 27077
rect 30904 27044 30920 27061
rect 30458 27027 30660 27044
rect 29700 26980 30660 27027
rect 30718 27027 30920 27044
rect 31476 27044 31492 27061
rect 31922 27061 32510 27077
rect 31922 27044 31938 27061
rect 31476 27027 31678 27044
rect 30718 26980 31678 27027
rect 31736 27027 31938 27044
rect 32494 27044 32510 27061
rect 32940 27061 33528 27077
rect 32940 27044 32956 27061
rect 32494 27027 32696 27044
rect 31736 26980 32696 27027
rect 32754 27027 32956 27044
rect 33512 27044 33528 27061
rect 33512 27027 33714 27044
rect 32754 26980 33714 27027
rect 17484 26333 18444 26380
rect 17484 26316 17686 26333
rect 17670 26299 17686 26316
rect 18242 26316 18444 26333
rect 18502 26333 19462 26380
rect 18502 26316 18704 26333
rect 18242 26299 18258 26316
rect 17670 26283 18258 26299
rect 18688 26299 18704 26316
rect 19260 26316 19462 26333
rect 19520 26333 20480 26380
rect 19520 26316 19722 26333
rect 19260 26299 19276 26316
rect 18688 26283 19276 26299
rect 19706 26299 19722 26316
rect 20278 26316 20480 26333
rect 20538 26333 21498 26380
rect 20538 26316 20740 26333
rect 20278 26299 20294 26316
rect 19706 26283 20294 26299
rect 20724 26299 20740 26316
rect 21296 26316 21498 26333
rect 21556 26333 22516 26380
rect 21556 26316 21758 26333
rect 21296 26299 21312 26316
rect 20724 26283 21312 26299
rect 21742 26299 21758 26316
rect 22314 26316 22516 26333
rect 22574 26333 23534 26380
rect 22574 26316 22776 26333
rect 22314 26299 22330 26316
rect 21742 26283 22330 26299
rect 22760 26299 22776 26316
rect 23332 26316 23534 26333
rect 23592 26333 24552 26380
rect 23592 26316 23794 26333
rect 23332 26299 23348 26316
rect 22760 26283 23348 26299
rect 23778 26299 23794 26316
rect 24350 26316 24552 26333
rect 24610 26333 25570 26380
rect 24610 26316 24812 26333
rect 24350 26299 24366 26316
rect 23778 26283 24366 26299
rect 24796 26299 24812 26316
rect 25368 26316 25570 26333
rect 25628 26333 26588 26380
rect 25628 26316 25830 26333
rect 25368 26299 25384 26316
rect 24796 26283 25384 26299
rect 25814 26299 25830 26316
rect 26386 26316 26588 26333
rect 26646 26333 27606 26380
rect 26646 26316 26848 26333
rect 26386 26299 26402 26316
rect 25814 26283 26402 26299
rect 26832 26299 26848 26316
rect 27404 26316 27606 26333
rect 27664 26333 28624 26380
rect 27664 26316 27866 26333
rect 27404 26299 27420 26316
rect 26832 26283 27420 26299
rect 27850 26299 27866 26316
rect 28422 26316 28624 26333
rect 28682 26333 29642 26380
rect 28682 26316 28884 26333
rect 28422 26299 28438 26316
rect 27850 26283 28438 26299
rect 28868 26299 28884 26316
rect 29440 26316 29642 26333
rect 29700 26333 30660 26380
rect 29700 26316 29902 26333
rect 29440 26299 29456 26316
rect 28868 26283 29456 26299
rect 29886 26299 29902 26316
rect 30458 26316 30660 26333
rect 30718 26333 31678 26380
rect 30718 26316 30920 26333
rect 30458 26299 30474 26316
rect 29886 26283 30474 26299
rect 30904 26299 30920 26316
rect 31476 26316 31678 26333
rect 31736 26333 32696 26380
rect 31736 26316 31938 26333
rect 31476 26299 31492 26316
rect 30904 26283 31492 26299
rect 31922 26299 31938 26316
rect 32494 26316 32696 26333
rect 32754 26333 33714 26380
rect 32754 26316 32956 26333
rect 32494 26299 32510 26316
rect 31922 26283 32510 26299
rect 32940 26299 32956 26316
rect 33512 26316 33714 26333
rect 33512 26299 33528 26316
rect 32940 26283 33528 26299
rect 17670 25925 18258 25941
rect 17670 25908 17686 25925
rect 17484 25891 17686 25908
rect 18242 25908 18258 25925
rect 18688 25925 19276 25941
rect 18688 25908 18704 25925
rect 18242 25891 18444 25908
rect 17484 25844 18444 25891
rect 18502 25891 18704 25908
rect 19260 25908 19276 25925
rect 19706 25925 20294 25941
rect 19706 25908 19722 25925
rect 19260 25891 19462 25908
rect 18502 25844 19462 25891
rect 19520 25891 19722 25908
rect 20278 25908 20294 25925
rect 20724 25925 21312 25941
rect 20724 25908 20740 25925
rect 20278 25891 20480 25908
rect 19520 25844 20480 25891
rect 20538 25891 20740 25908
rect 21296 25908 21312 25925
rect 21742 25925 22330 25941
rect 21742 25908 21758 25925
rect 21296 25891 21498 25908
rect 20538 25844 21498 25891
rect 21556 25891 21758 25908
rect 22314 25908 22330 25925
rect 22760 25925 23348 25941
rect 22760 25908 22776 25925
rect 22314 25891 22516 25908
rect 21556 25844 22516 25891
rect 22574 25891 22776 25908
rect 23332 25908 23348 25925
rect 23778 25925 24366 25941
rect 23778 25908 23794 25925
rect 23332 25891 23534 25908
rect 22574 25844 23534 25891
rect 23592 25891 23794 25908
rect 24350 25908 24366 25925
rect 24796 25925 25384 25941
rect 24796 25908 24812 25925
rect 24350 25891 24552 25908
rect 23592 25844 24552 25891
rect 24610 25891 24812 25908
rect 25368 25908 25384 25925
rect 25814 25925 26402 25941
rect 25814 25908 25830 25925
rect 25368 25891 25570 25908
rect 24610 25844 25570 25891
rect 25628 25891 25830 25908
rect 26386 25908 26402 25925
rect 26832 25925 27420 25941
rect 26832 25908 26848 25925
rect 26386 25891 26588 25908
rect 25628 25844 26588 25891
rect 26646 25891 26848 25908
rect 27404 25908 27420 25925
rect 27850 25925 28438 25941
rect 27850 25908 27866 25925
rect 27404 25891 27606 25908
rect 26646 25844 27606 25891
rect 27664 25891 27866 25908
rect 28422 25908 28438 25925
rect 28868 25925 29456 25941
rect 28868 25908 28884 25925
rect 28422 25891 28624 25908
rect 27664 25844 28624 25891
rect 28682 25891 28884 25908
rect 29440 25908 29456 25925
rect 29886 25925 30474 25941
rect 29886 25908 29902 25925
rect 29440 25891 29642 25908
rect 28682 25844 29642 25891
rect 29700 25891 29902 25908
rect 30458 25908 30474 25925
rect 30904 25925 31492 25941
rect 30904 25908 30920 25925
rect 30458 25891 30660 25908
rect 29700 25844 30660 25891
rect 30718 25891 30920 25908
rect 31476 25908 31492 25925
rect 31922 25925 32510 25941
rect 31922 25908 31938 25925
rect 31476 25891 31678 25908
rect 30718 25844 31678 25891
rect 31736 25891 31938 25908
rect 32494 25908 32510 25925
rect 32940 25925 33528 25941
rect 32940 25908 32956 25925
rect 32494 25891 32696 25908
rect 31736 25844 32696 25891
rect 32754 25891 32956 25908
rect 33512 25908 33528 25925
rect 33512 25891 33714 25908
rect 32754 25844 33714 25891
rect 17484 25197 18444 25244
rect 17484 25180 17686 25197
rect 17670 25163 17686 25180
rect 18242 25180 18444 25197
rect 18502 25197 19462 25244
rect 18502 25180 18704 25197
rect 18242 25163 18258 25180
rect 17670 25147 18258 25163
rect 18688 25163 18704 25180
rect 19260 25180 19462 25197
rect 19520 25197 20480 25244
rect 19520 25180 19722 25197
rect 19260 25163 19276 25180
rect 18688 25147 19276 25163
rect 19706 25163 19722 25180
rect 20278 25180 20480 25197
rect 20538 25197 21498 25244
rect 20538 25180 20740 25197
rect 20278 25163 20294 25180
rect 19706 25147 20294 25163
rect 20724 25163 20740 25180
rect 21296 25180 21498 25197
rect 21556 25197 22516 25244
rect 21556 25180 21758 25197
rect 21296 25163 21312 25180
rect 20724 25147 21312 25163
rect 21742 25163 21758 25180
rect 22314 25180 22516 25197
rect 22574 25197 23534 25244
rect 22574 25180 22776 25197
rect 22314 25163 22330 25180
rect 21742 25147 22330 25163
rect 22760 25163 22776 25180
rect 23332 25180 23534 25197
rect 23592 25197 24552 25244
rect 23592 25180 23794 25197
rect 23332 25163 23348 25180
rect 22760 25147 23348 25163
rect 23778 25163 23794 25180
rect 24350 25180 24552 25197
rect 24610 25197 25570 25244
rect 24610 25180 24812 25197
rect 24350 25163 24366 25180
rect 23778 25147 24366 25163
rect 24796 25163 24812 25180
rect 25368 25180 25570 25197
rect 25628 25197 26588 25244
rect 25628 25180 25830 25197
rect 25368 25163 25384 25180
rect 24796 25147 25384 25163
rect 25814 25163 25830 25180
rect 26386 25180 26588 25197
rect 26646 25197 27606 25244
rect 26646 25180 26848 25197
rect 26386 25163 26402 25180
rect 25814 25147 26402 25163
rect 26832 25163 26848 25180
rect 27404 25180 27606 25197
rect 27664 25197 28624 25244
rect 27664 25180 27866 25197
rect 27404 25163 27420 25180
rect 26832 25147 27420 25163
rect 27850 25163 27866 25180
rect 28422 25180 28624 25197
rect 28682 25197 29642 25244
rect 28682 25180 28884 25197
rect 28422 25163 28438 25180
rect 27850 25147 28438 25163
rect 28868 25163 28884 25180
rect 29440 25180 29642 25197
rect 29700 25197 30660 25244
rect 29700 25180 29902 25197
rect 29440 25163 29456 25180
rect 28868 25147 29456 25163
rect 29886 25163 29902 25180
rect 30458 25180 30660 25197
rect 30718 25197 31678 25244
rect 30718 25180 30920 25197
rect 30458 25163 30474 25180
rect 29886 25147 30474 25163
rect 30904 25163 30920 25180
rect 31476 25180 31678 25197
rect 31736 25197 32696 25244
rect 31736 25180 31938 25197
rect 31476 25163 31492 25180
rect 30904 25147 31492 25163
rect 31922 25163 31938 25180
rect 32494 25180 32696 25197
rect 32754 25197 33714 25244
rect 32754 25180 32956 25197
rect 32494 25163 32510 25180
rect 31922 25147 32510 25163
rect 32940 25163 32956 25180
rect 33512 25180 33714 25197
rect 33512 25163 33528 25180
rect 32940 25147 33528 25163
rect 17670 24789 18258 24805
rect 17670 24772 17686 24789
rect 17484 24755 17686 24772
rect 18242 24772 18258 24789
rect 18688 24789 19276 24805
rect 18688 24772 18704 24789
rect 18242 24755 18444 24772
rect 17484 24708 18444 24755
rect 18502 24755 18704 24772
rect 19260 24772 19276 24789
rect 19706 24789 20294 24805
rect 19706 24772 19722 24789
rect 19260 24755 19462 24772
rect 18502 24708 19462 24755
rect 19520 24755 19722 24772
rect 20278 24772 20294 24789
rect 20724 24789 21312 24805
rect 20724 24772 20740 24789
rect 20278 24755 20480 24772
rect 19520 24708 20480 24755
rect 20538 24755 20740 24772
rect 21296 24772 21312 24789
rect 21742 24789 22330 24805
rect 21742 24772 21758 24789
rect 21296 24755 21498 24772
rect 20538 24708 21498 24755
rect 21556 24755 21758 24772
rect 22314 24772 22330 24789
rect 22760 24789 23348 24805
rect 22760 24772 22776 24789
rect 22314 24755 22516 24772
rect 21556 24708 22516 24755
rect 22574 24755 22776 24772
rect 23332 24772 23348 24789
rect 23778 24789 24366 24805
rect 23778 24772 23794 24789
rect 23332 24755 23534 24772
rect 22574 24708 23534 24755
rect 23592 24755 23794 24772
rect 24350 24772 24366 24789
rect 24796 24789 25384 24805
rect 24796 24772 24812 24789
rect 24350 24755 24552 24772
rect 23592 24708 24552 24755
rect 24610 24755 24812 24772
rect 25368 24772 25384 24789
rect 25814 24789 26402 24805
rect 25814 24772 25830 24789
rect 25368 24755 25570 24772
rect 24610 24708 25570 24755
rect 25628 24755 25830 24772
rect 26386 24772 26402 24789
rect 26832 24789 27420 24805
rect 26832 24772 26848 24789
rect 26386 24755 26588 24772
rect 25628 24708 26588 24755
rect 26646 24755 26848 24772
rect 27404 24772 27420 24789
rect 27850 24789 28438 24805
rect 27850 24772 27866 24789
rect 27404 24755 27606 24772
rect 26646 24708 27606 24755
rect 27664 24755 27866 24772
rect 28422 24772 28438 24789
rect 28868 24789 29456 24805
rect 28868 24772 28884 24789
rect 28422 24755 28624 24772
rect 27664 24708 28624 24755
rect 28682 24755 28884 24772
rect 29440 24772 29456 24789
rect 29886 24789 30474 24805
rect 29886 24772 29902 24789
rect 29440 24755 29642 24772
rect 28682 24708 29642 24755
rect 29700 24755 29902 24772
rect 30458 24772 30474 24789
rect 30904 24789 31492 24805
rect 30904 24772 30920 24789
rect 30458 24755 30660 24772
rect 29700 24708 30660 24755
rect 30718 24755 30920 24772
rect 31476 24772 31492 24789
rect 31922 24789 32510 24805
rect 31922 24772 31938 24789
rect 31476 24755 31678 24772
rect 30718 24708 31678 24755
rect 31736 24755 31938 24772
rect 32494 24772 32510 24789
rect 32940 24789 33528 24805
rect 32940 24772 32956 24789
rect 32494 24755 32696 24772
rect 31736 24708 32696 24755
rect 32754 24755 32956 24772
rect 33512 24772 33528 24789
rect 33512 24755 33714 24772
rect 32754 24708 33714 24755
rect 17484 24061 18444 24108
rect 17484 24044 17686 24061
rect 17670 24027 17686 24044
rect 18242 24044 18444 24061
rect 18502 24061 19462 24108
rect 18502 24044 18704 24061
rect 18242 24027 18258 24044
rect 17670 24011 18258 24027
rect 18688 24027 18704 24044
rect 19260 24044 19462 24061
rect 19520 24061 20480 24108
rect 19520 24044 19722 24061
rect 19260 24027 19276 24044
rect 18688 24011 19276 24027
rect 19706 24027 19722 24044
rect 20278 24044 20480 24061
rect 20538 24061 21498 24108
rect 20538 24044 20740 24061
rect 20278 24027 20294 24044
rect 19706 24011 20294 24027
rect 20724 24027 20740 24044
rect 21296 24044 21498 24061
rect 21556 24061 22516 24108
rect 21556 24044 21758 24061
rect 21296 24027 21312 24044
rect 20724 24011 21312 24027
rect 21742 24027 21758 24044
rect 22314 24044 22516 24061
rect 22574 24061 23534 24108
rect 22574 24044 22776 24061
rect 22314 24027 22330 24044
rect 21742 24011 22330 24027
rect 22760 24027 22776 24044
rect 23332 24044 23534 24061
rect 23592 24061 24552 24108
rect 23592 24044 23794 24061
rect 23332 24027 23348 24044
rect 22760 24011 23348 24027
rect 23778 24027 23794 24044
rect 24350 24044 24552 24061
rect 24610 24061 25570 24108
rect 24610 24044 24812 24061
rect 24350 24027 24366 24044
rect 23778 24011 24366 24027
rect 24796 24027 24812 24044
rect 25368 24044 25570 24061
rect 25628 24061 26588 24108
rect 25628 24044 25830 24061
rect 25368 24027 25384 24044
rect 24796 24011 25384 24027
rect 25814 24027 25830 24044
rect 26386 24044 26588 24061
rect 26646 24061 27606 24108
rect 26646 24044 26848 24061
rect 26386 24027 26402 24044
rect 25814 24011 26402 24027
rect 26832 24027 26848 24044
rect 27404 24044 27606 24061
rect 27664 24061 28624 24108
rect 27664 24044 27866 24061
rect 27404 24027 27420 24044
rect 26832 24011 27420 24027
rect 27850 24027 27866 24044
rect 28422 24044 28624 24061
rect 28682 24061 29642 24108
rect 28682 24044 28884 24061
rect 28422 24027 28438 24044
rect 27850 24011 28438 24027
rect 28868 24027 28884 24044
rect 29440 24044 29642 24061
rect 29700 24061 30660 24108
rect 29700 24044 29902 24061
rect 29440 24027 29456 24044
rect 28868 24011 29456 24027
rect 29886 24027 29902 24044
rect 30458 24044 30660 24061
rect 30718 24061 31678 24108
rect 30718 24044 30920 24061
rect 30458 24027 30474 24044
rect 29886 24011 30474 24027
rect 30904 24027 30920 24044
rect 31476 24044 31678 24061
rect 31736 24061 32696 24108
rect 31736 24044 31938 24061
rect 31476 24027 31492 24044
rect 30904 24011 31492 24027
rect 31922 24027 31938 24044
rect 32494 24044 32696 24061
rect 32754 24061 33714 24108
rect 32754 24044 32956 24061
rect 32494 24027 32510 24044
rect 31922 24011 32510 24027
rect 32940 24027 32956 24044
rect 33512 24044 33714 24061
rect 33512 24027 33528 24044
rect 32940 24011 33528 24027
rect 18656 23015 19244 23031
rect 18656 22998 18672 23015
rect 18470 22981 18672 22998
rect 19228 22998 19244 23015
rect 19674 23015 20262 23031
rect 19674 22998 19690 23015
rect 19228 22981 19430 22998
rect 18470 22934 19430 22981
rect 19488 22981 19690 22998
rect 20246 22998 20262 23015
rect 20692 23015 21280 23031
rect 20692 22998 20708 23015
rect 20246 22981 20448 22998
rect 19488 22934 20448 22981
rect 20506 22981 20708 22998
rect 21264 22998 21280 23015
rect 21710 23015 22298 23031
rect 21710 22998 21726 23015
rect 21264 22981 21466 22998
rect 20506 22934 21466 22981
rect 21524 22981 21726 22998
rect 22282 22998 22298 23015
rect 22728 23015 23316 23031
rect 22728 22998 22744 23015
rect 22282 22981 22484 22998
rect 21524 22934 22484 22981
rect 22542 22981 22744 22998
rect 23300 22998 23316 23015
rect 23746 23015 24334 23031
rect 23746 22998 23762 23015
rect 23300 22981 23502 22998
rect 22542 22934 23502 22981
rect 23560 22981 23762 22998
rect 24318 22998 24334 23015
rect 24764 23015 25352 23031
rect 24764 22998 24780 23015
rect 24318 22981 24520 22998
rect 23560 22934 24520 22981
rect 24578 22981 24780 22998
rect 25336 22998 25352 23015
rect 25782 23015 26370 23031
rect 25782 22998 25798 23015
rect 25336 22981 25538 22998
rect 24578 22934 25538 22981
rect 25596 22981 25798 22998
rect 26354 22998 26370 23015
rect 26800 23015 27388 23031
rect 26800 22998 26816 23015
rect 26354 22981 26556 22998
rect 25596 22934 26556 22981
rect 26614 22981 26816 22998
rect 27372 22998 27388 23015
rect 27818 23015 28406 23031
rect 27818 22998 27834 23015
rect 27372 22981 27574 22998
rect 26614 22934 27574 22981
rect 27632 22981 27834 22998
rect 28390 22998 28406 23015
rect 28836 23015 29424 23031
rect 28836 22998 28852 23015
rect 28390 22981 28592 22998
rect 27632 22934 28592 22981
rect 28650 22981 28852 22998
rect 29408 22998 29424 23015
rect 29854 23015 30442 23031
rect 29854 22998 29870 23015
rect 29408 22981 29610 22998
rect 28650 22934 29610 22981
rect 29668 22981 29870 22998
rect 30426 22998 30442 23015
rect 30872 23015 31460 23031
rect 30872 22998 30888 23015
rect 30426 22981 30628 22998
rect 29668 22934 30628 22981
rect 30686 22981 30888 22998
rect 31444 22998 31460 23015
rect 31890 23015 32478 23031
rect 31890 22998 31906 23015
rect 31444 22981 31646 22998
rect 30686 22934 31646 22981
rect 31704 22981 31906 22998
rect 32462 22998 32478 23015
rect 32908 23015 33496 23031
rect 32908 22998 32924 23015
rect 32462 22981 32664 22998
rect 31704 22934 32664 22981
rect 32722 22981 32924 22998
rect 33480 22998 33496 23015
rect 33480 22981 33682 22998
rect 32722 22934 33682 22981
rect 18470 22287 19430 22334
rect 18470 22270 18672 22287
rect 18656 22253 18672 22270
rect 19228 22270 19430 22287
rect 19488 22287 20448 22334
rect 19488 22270 19690 22287
rect 19228 22253 19244 22270
rect 18656 22237 19244 22253
rect 19674 22253 19690 22270
rect 20246 22270 20448 22287
rect 20506 22287 21466 22334
rect 20506 22270 20708 22287
rect 20246 22253 20262 22270
rect 19674 22237 20262 22253
rect 20692 22253 20708 22270
rect 21264 22270 21466 22287
rect 21524 22287 22484 22334
rect 21524 22270 21726 22287
rect 21264 22253 21280 22270
rect 20692 22237 21280 22253
rect 21710 22253 21726 22270
rect 22282 22270 22484 22287
rect 22542 22287 23502 22334
rect 22542 22270 22744 22287
rect 22282 22253 22298 22270
rect 21710 22237 22298 22253
rect 22728 22253 22744 22270
rect 23300 22270 23502 22287
rect 23560 22287 24520 22334
rect 23560 22270 23762 22287
rect 23300 22253 23316 22270
rect 22728 22237 23316 22253
rect 23746 22253 23762 22270
rect 24318 22270 24520 22287
rect 24578 22287 25538 22334
rect 24578 22270 24780 22287
rect 24318 22253 24334 22270
rect 23746 22237 24334 22253
rect 24764 22253 24780 22270
rect 25336 22270 25538 22287
rect 25596 22287 26556 22334
rect 25596 22270 25798 22287
rect 25336 22253 25352 22270
rect 24764 22237 25352 22253
rect 25782 22253 25798 22270
rect 26354 22270 26556 22287
rect 26614 22287 27574 22334
rect 26614 22270 26816 22287
rect 26354 22253 26370 22270
rect 25782 22237 26370 22253
rect 26800 22253 26816 22270
rect 27372 22270 27574 22287
rect 27632 22287 28592 22334
rect 27632 22270 27834 22287
rect 27372 22253 27388 22270
rect 26800 22237 27388 22253
rect 27818 22253 27834 22270
rect 28390 22270 28592 22287
rect 28650 22287 29610 22334
rect 28650 22270 28852 22287
rect 28390 22253 28406 22270
rect 27818 22237 28406 22253
rect 28836 22253 28852 22270
rect 29408 22270 29610 22287
rect 29668 22287 30628 22334
rect 29668 22270 29870 22287
rect 29408 22253 29424 22270
rect 28836 22237 29424 22253
rect 29854 22253 29870 22270
rect 30426 22270 30628 22287
rect 30686 22287 31646 22334
rect 30686 22270 30888 22287
rect 30426 22253 30442 22270
rect 29854 22237 30442 22253
rect 30872 22253 30888 22270
rect 31444 22270 31646 22287
rect 31704 22287 32664 22334
rect 31704 22270 31906 22287
rect 31444 22253 31460 22270
rect 30872 22237 31460 22253
rect 31890 22253 31906 22270
rect 32462 22270 32664 22287
rect 32722 22287 33682 22334
rect 32722 22270 32924 22287
rect 32462 22253 32478 22270
rect 31890 22237 32478 22253
rect 32908 22253 32924 22270
rect 33480 22270 33682 22287
rect 33480 22253 33496 22270
rect 32908 22237 33496 22253
rect 14648 21931 14756 21947
rect 14648 21914 14664 21931
rect 14622 21897 14664 21914
rect 14740 21914 14756 21931
rect 14866 21931 14974 21947
rect 14866 21914 14882 21931
rect 14740 21897 14782 21914
rect 14622 21850 14782 21897
rect 14840 21897 14882 21914
rect 14958 21914 14974 21931
rect 15084 21931 15192 21947
rect 15084 21914 15100 21931
rect 14958 21897 15000 21914
rect 14840 21850 15000 21897
rect 15058 21897 15100 21914
rect 15176 21914 15192 21931
rect 15302 21931 15410 21947
rect 15302 21914 15318 21931
rect 15176 21897 15218 21914
rect 15058 21850 15218 21897
rect 15276 21897 15318 21914
rect 15394 21914 15410 21931
rect 15520 21931 15628 21947
rect 15520 21914 15536 21931
rect 15394 21897 15436 21914
rect 15276 21850 15436 21897
rect 15494 21897 15536 21914
rect 15612 21914 15628 21931
rect 15738 21931 15846 21947
rect 15738 21914 15754 21931
rect 15612 21897 15654 21914
rect 15494 21850 15654 21897
rect 15712 21897 15754 21914
rect 15830 21914 15846 21931
rect 15956 21931 16064 21947
rect 15956 21914 15972 21931
rect 15830 21897 15872 21914
rect 15712 21850 15872 21897
rect 15930 21897 15972 21914
rect 16048 21914 16064 21931
rect 16174 21931 16282 21947
rect 16174 21914 16190 21931
rect 16048 21897 16090 21914
rect 15930 21850 16090 21897
rect 16148 21897 16190 21914
rect 16266 21914 16282 21931
rect 16392 21931 16500 21947
rect 16392 21914 16408 21931
rect 16266 21897 16308 21914
rect 16148 21850 16308 21897
rect 16366 21897 16408 21914
rect 16484 21914 16500 21931
rect 16610 21931 16718 21947
rect 16610 21914 16626 21931
rect 16484 21897 16526 21914
rect 16366 21850 16526 21897
rect 16584 21897 16626 21914
rect 16702 21914 16718 21931
rect 16702 21897 16744 21914
rect 16584 21850 16744 21897
rect 18656 21759 19244 21775
rect 18656 21742 18672 21759
rect 18470 21725 18672 21742
rect 19228 21742 19244 21759
rect 19674 21759 20262 21775
rect 19674 21742 19690 21759
rect 19228 21725 19430 21742
rect 18470 21678 19430 21725
rect 19488 21725 19690 21742
rect 20246 21742 20262 21759
rect 20692 21759 21280 21775
rect 20692 21742 20708 21759
rect 20246 21725 20448 21742
rect 19488 21678 20448 21725
rect 20506 21725 20708 21742
rect 21264 21742 21280 21759
rect 21710 21759 22298 21775
rect 21710 21742 21726 21759
rect 21264 21725 21466 21742
rect 20506 21678 21466 21725
rect 21524 21725 21726 21742
rect 22282 21742 22298 21759
rect 22728 21759 23316 21775
rect 22728 21742 22744 21759
rect 22282 21725 22484 21742
rect 21524 21678 22484 21725
rect 22542 21725 22744 21742
rect 23300 21742 23316 21759
rect 23746 21759 24334 21775
rect 23746 21742 23762 21759
rect 23300 21725 23502 21742
rect 22542 21678 23502 21725
rect 23560 21725 23762 21742
rect 24318 21742 24334 21759
rect 24764 21759 25352 21775
rect 24764 21742 24780 21759
rect 24318 21725 24520 21742
rect 23560 21678 24520 21725
rect 24578 21725 24780 21742
rect 25336 21742 25352 21759
rect 25782 21759 26370 21775
rect 25782 21742 25798 21759
rect 25336 21725 25538 21742
rect 24578 21678 25538 21725
rect 25596 21725 25798 21742
rect 26354 21742 26370 21759
rect 26800 21759 27388 21775
rect 26800 21742 26816 21759
rect 26354 21725 26556 21742
rect 25596 21678 26556 21725
rect 26614 21725 26816 21742
rect 27372 21742 27388 21759
rect 27818 21759 28406 21775
rect 27818 21742 27834 21759
rect 27372 21725 27574 21742
rect 26614 21678 27574 21725
rect 27632 21725 27834 21742
rect 28390 21742 28406 21759
rect 28836 21759 29424 21775
rect 28836 21742 28852 21759
rect 28390 21725 28592 21742
rect 27632 21678 28592 21725
rect 28650 21725 28852 21742
rect 29408 21742 29424 21759
rect 29854 21759 30442 21775
rect 29854 21742 29870 21759
rect 29408 21725 29610 21742
rect 28650 21678 29610 21725
rect 29668 21725 29870 21742
rect 30426 21742 30442 21759
rect 30872 21759 31460 21775
rect 30872 21742 30888 21759
rect 30426 21725 30628 21742
rect 29668 21678 30628 21725
rect 30686 21725 30888 21742
rect 31444 21742 31460 21759
rect 31890 21759 32478 21775
rect 31890 21742 31906 21759
rect 31444 21725 31646 21742
rect 30686 21678 31646 21725
rect 31704 21725 31906 21742
rect 32462 21742 32478 21759
rect 32908 21759 33496 21775
rect 32908 21742 32924 21759
rect 32462 21725 32664 21742
rect 31704 21678 32664 21725
rect 32722 21725 32924 21742
rect 33480 21742 33496 21759
rect 33480 21725 33682 21742
rect 32722 21678 33682 21725
rect 14622 21403 14782 21450
rect 14622 21386 14664 21403
rect 14648 21369 14664 21386
rect 14740 21386 14782 21403
rect 14840 21403 15000 21450
rect 14840 21386 14882 21403
rect 14740 21369 14756 21386
rect 14648 21353 14756 21369
rect 14866 21369 14882 21386
rect 14958 21386 15000 21403
rect 15058 21403 15218 21450
rect 15058 21386 15100 21403
rect 14958 21369 14974 21386
rect 14866 21353 14974 21369
rect 15084 21369 15100 21386
rect 15176 21386 15218 21403
rect 15276 21403 15436 21450
rect 15276 21386 15318 21403
rect 15176 21369 15192 21386
rect 15084 21353 15192 21369
rect 15302 21369 15318 21386
rect 15394 21386 15436 21403
rect 15494 21403 15654 21450
rect 15494 21386 15536 21403
rect 15394 21369 15410 21386
rect 15302 21353 15410 21369
rect 15520 21369 15536 21386
rect 15612 21386 15654 21403
rect 15712 21403 15872 21450
rect 15712 21386 15754 21403
rect 15612 21369 15628 21386
rect 15520 21353 15628 21369
rect 15738 21369 15754 21386
rect 15830 21386 15872 21403
rect 15930 21403 16090 21450
rect 15930 21386 15972 21403
rect 15830 21369 15846 21386
rect 15738 21353 15846 21369
rect 15956 21369 15972 21386
rect 16048 21386 16090 21403
rect 16148 21403 16308 21450
rect 16148 21386 16190 21403
rect 16048 21369 16064 21386
rect 15956 21353 16064 21369
rect 16174 21369 16190 21386
rect 16266 21386 16308 21403
rect 16366 21403 16526 21450
rect 16366 21386 16408 21403
rect 16266 21369 16282 21386
rect 16174 21353 16282 21369
rect 16392 21369 16408 21386
rect 16484 21386 16526 21403
rect 16584 21403 16744 21450
rect 16584 21386 16626 21403
rect 16484 21369 16500 21386
rect 16392 21353 16500 21369
rect 16610 21369 16626 21386
rect 16702 21386 16744 21403
rect 16702 21369 16718 21386
rect 16610 21353 16718 21369
rect 18470 21031 19430 21078
rect 18470 21014 18672 21031
rect 14648 20993 14756 21009
rect 14648 20976 14664 20993
rect 14622 20959 14664 20976
rect 14740 20976 14756 20993
rect 14866 20993 14974 21009
rect 14866 20976 14882 20993
rect 14740 20959 14782 20976
rect 14622 20912 14782 20959
rect 14840 20959 14882 20976
rect 14958 20976 14974 20993
rect 15084 20993 15192 21009
rect 15084 20976 15100 20993
rect 14958 20959 15000 20976
rect 14840 20912 15000 20959
rect 15058 20959 15100 20976
rect 15176 20976 15192 20993
rect 15302 20993 15410 21009
rect 15302 20976 15318 20993
rect 15176 20959 15218 20976
rect 15058 20912 15218 20959
rect 15276 20959 15318 20976
rect 15394 20976 15410 20993
rect 15520 20993 15628 21009
rect 15520 20976 15536 20993
rect 15394 20959 15436 20976
rect 15276 20912 15436 20959
rect 15494 20959 15536 20976
rect 15612 20976 15628 20993
rect 15738 20993 15846 21009
rect 15738 20976 15754 20993
rect 15612 20959 15654 20976
rect 15494 20912 15654 20959
rect 15712 20959 15754 20976
rect 15830 20976 15846 20993
rect 15956 20993 16064 21009
rect 15956 20976 15972 20993
rect 15830 20959 15872 20976
rect 15712 20912 15872 20959
rect 15930 20959 15972 20976
rect 16048 20976 16064 20993
rect 16174 20993 16282 21009
rect 16174 20976 16190 20993
rect 16048 20959 16090 20976
rect 15930 20912 16090 20959
rect 16148 20959 16190 20976
rect 16266 20976 16282 20993
rect 16392 20993 16500 21009
rect 16392 20976 16408 20993
rect 16266 20959 16308 20976
rect 16148 20912 16308 20959
rect 16366 20959 16408 20976
rect 16484 20976 16500 20993
rect 16610 20993 16718 21009
rect 16610 20976 16626 20993
rect 16484 20959 16526 20976
rect 16366 20912 16526 20959
rect 16584 20959 16626 20976
rect 16702 20976 16718 20993
rect 18656 20997 18672 21014
rect 19228 21014 19430 21031
rect 19488 21031 20448 21078
rect 19488 21014 19690 21031
rect 19228 20997 19244 21014
rect 18656 20981 19244 20997
rect 19674 20997 19690 21014
rect 20246 21014 20448 21031
rect 20506 21031 21466 21078
rect 20506 21014 20708 21031
rect 20246 20997 20262 21014
rect 19674 20981 20262 20997
rect 20692 20997 20708 21014
rect 21264 21014 21466 21031
rect 21524 21031 22484 21078
rect 21524 21014 21726 21031
rect 21264 20997 21280 21014
rect 20692 20981 21280 20997
rect 21710 20997 21726 21014
rect 22282 21014 22484 21031
rect 22542 21031 23502 21078
rect 22542 21014 22744 21031
rect 22282 20997 22298 21014
rect 21710 20981 22298 20997
rect 22728 20997 22744 21014
rect 23300 21014 23502 21031
rect 23560 21031 24520 21078
rect 23560 21014 23762 21031
rect 23300 20997 23316 21014
rect 22728 20981 23316 20997
rect 23746 20997 23762 21014
rect 24318 21014 24520 21031
rect 24578 21031 25538 21078
rect 24578 21014 24780 21031
rect 24318 20997 24334 21014
rect 23746 20981 24334 20997
rect 24764 20997 24780 21014
rect 25336 21014 25538 21031
rect 25596 21031 26556 21078
rect 25596 21014 25798 21031
rect 25336 20997 25352 21014
rect 24764 20981 25352 20997
rect 25782 20997 25798 21014
rect 26354 21014 26556 21031
rect 26614 21031 27574 21078
rect 26614 21014 26816 21031
rect 26354 20997 26370 21014
rect 25782 20981 26370 20997
rect 26800 20997 26816 21014
rect 27372 21014 27574 21031
rect 27632 21031 28592 21078
rect 27632 21014 27834 21031
rect 27372 20997 27388 21014
rect 26800 20981 27388 20997
rect 27818 20997 27834 21014
rect 28390 21014 28592 21031
rect 28650 21031 29610 21078
rect 28650 21014 28852 21031
rect 28390 20997 28406 21014
rect 27818 20981 28406 20997
rect 28836 20997 28852 21014
rect 29408 21014 29610 21031
rect 29668 21031 30628 21078
rect 29668 21014 29870 21031
rect 29408 20997 29424 21014
rect 28836 20981 29424 20997
rect 29854 20997 29870 21014
rect 30426 21014 30628 21031
rect 30686 21031 31646 21078
rect 30686 21014 30888 21031
rect 30426 20997 30442 21014
rect 29854 20981 30442 20997
rect 30872 20997 30888 21014
rect 31444 21014 31646 21031
rect 31704 21031 32664 21078
rect 31704 21014 31906 21031
rect 31444 20997 31460 21014
rect 30872 20981 31460 20997
rect 31890 20997 31906 21014
rect 32462 21014 32664 21031
rect 32722 21031 33682 21078
rect 32722 21014 32924 21031
rect 32462 20997 32478 21014
rect 31890 20981 32478 20997
rect 32908 20997 32924 21014
rect 33480 21014 33682 21031
rect 33480 20997 33496 21014
rect 32908 20981 33496 20997
rect 16702 20959 16744 20976
rect 16584 20912 16744 20959
rect 14622 20465 14782 20512
rect 14622 20448 14664 20465
rect 14648 20431 14664 20448
rect 14740 20448 14782 20465
rect 14840 20465 15000 20512
rect 14840 20448 14882 20465
rect 14740 20431 14756 20448
rect 14648 20415 14756 20431
rect 14866 20431 14882 20448
rect 14958 20448 15000 20465
rect 15058 20465 15218 20512
rect 15058 20448 15100 20465
rect 14958 20431 14974 20448
rect 14866 20415 14974 20431
rect 15084 20431 15100 20448
rect 15176 20448 15218 20465
rect 15276 20465 15436 20512
rect 15276 20448 15318 20465
rect 15176 20431 15192 20448
rect 15084 20415 15192 20431
rect 15302 20431 15318 20448
rect 15394 20448 15436 20465
rect 15494 20465 15654 20512
rect 15494 20448 15536 20465
rect 15394 20431 15410 20448
rect 15302 20415 15410 20431
rect 15520 20431 15536 20448
rect 15612 20448 15654 20465
rect 15712 20465 15872 20512
rect 15712 20448 15754 20465
rect 15612 20431 15628 20448
rect 15520 20415 15628 20431
rect 15738 20431 15754 20448
rect 15830 20448 15872 20465
rect 15930 20465 16090 20512
rect 15930 20448 15972 20465
rect 15830 20431 15846 20448
rect 15738 20415 15846 20431
rect 15956 20431 15972 20448
rect 16048 20448 16090 20465
rect 16148 20465 16308 20512
rect 16148 20448 16190 20465
rect 16048 20431 16064 20448
rect 15956 20415 16064 20431
rect 16174 20431 16190 20448
rect 16266 20448 16308 20465
rect 16366 20465 16526 20512
rect 16366 20448 16408 20465
rect 16266 20431 16282 20448
rect 16174 20415 16282 20431
rect 16392 20431 16408 20448
rect 16484 20448 16526 20465
rect 16584 20465 16744 20512
rect 18656 20503 19244 20519
rect 18656 20486 18672 20503
rect 16584 20448 16626 20465
rect 16484 20431 16500 20448
rect 16392 20415 16500 20431
rect 16610 20431 16626 20448
rect 16702 20448 16744 20465
rect 18470 20469 18672 20486
rect 19228 20486 19244 20503
rect 19674 20503 20262 20519
rect 19674 20486 19690 20503
rect 19228 20469 19430 20486
rect 16702 20431 16718 20448
rect 16610 20415 16718 20431
rect 18470 20422 19430 20469
rect 19488 20469 19690 20486
rect 20246 20486 20262 20503
rect 20692 20503 21280 20519
rect 20692 20486 20708 20503
rect 20246 20469 20448 20486
rect 19488 20422 20448 20469
rect 20506 20469 20708 20486
rect 21264 20486 21280 20503
rect 21710 20503 22298 20519
rect 21710 20486 21726 20503
rect 21264 20469 21466 20486
rect 20506 20422 21466 20469
rect 21524 20469 21726 20486
rect 22282 20486 22298 20503
rect 22728 20503 23316 20519
rect 22728 20486 22744 20503
rect 22282 20469 22484 20486
rect 21524 20422 22484 20469
rect 22542 20469 22744 20486
rect 23300 20486 23316 20503
rect 23746 20503 24334 20519
rect 23746 20486 23762 20503
rect 23300 20469 23502 20486
rect 22542 20422 23502 20469
rect 23560 20469 23762 20486
rect 24318 20486 24334 20503
rect 24764 20503 25352 20519
rect 24764 20486 24780 20503
rect 24318 20469 24520 20486
rect 23560 20422 24520 20469
rect 24578 20469 24780 20486
rect 25336 20486 25352 20503
rect 25782 20503 26370 20519
rect 25782 20486 25798 20503
rect 25336 20469 25538 20486
rect 24578 20422 25538 20469
rect 25596 20469 25798 20486
rect 26354 20486 26370 20503
rect 26800 20503 27388 20519
rect 26800 20486 26816 20503
rect 26354 20469 26556 20486
rect 25596 20422 26556 20469
rect 26614 20469 26816 20486
rect 27372 20486 27388 20503
rect 27818 20503 28406 20519
rect 27818 20486 27834 20503
rect 27372 20469 27574 20486
rect 26614 20422 27574 20469
rect 27632 20469 27834 20486
rect 28390 20486 28406 20503
rect 28836 20503 29424 20519
rect 28836 20486 28852 20503
rect 28390 20469 28592 20486
rect 27632 20422 28592 20469
rect 28650 20469 28852 20486
rect 29408 20486 29424 20503
rect 29854 20503 30442 20519
rect 29854 20486 29870 20503
rect 29408 20469 29610 20486
rect 28650 20422 29610 20469
rect 29668 20469 29870 20486
rect 30426 20486 30442 20503
rect 30872 20503 31460 20519
rect 30872 20486 30888 20503
rect 30426 20469 30628 20486
rect 29668 20422 30628 20469
rect 30686 20469 30888 20486
rect 31444 20486 31460 20503
rect 31890 20503 32478 20519
rect 31890 20486 31906 20503
rect 31444 20469 31646 20486
rect 30686 20422 31646 20469
rect 31704 20469 31906 20486
rect 32462 20486 32478 20503
rect 32908 20503 33496 20519
rect 32908 20486 32924 20503
rect 32462 20469 32664 20486
rect 31704 20422 32664 20469
rect 32722 20469 32924 20486
rect 33480 20486 33496 20503
rect 33480 20469 33682 20486
rect 32722 20422 33682 20469
rect 14648 20055 14756 20071
rect 14648 20038 14664 20055
rect 14622 20021 14664 20038
rect 14740 20038 14756 20055
rect 14866 20055 14974 20071
rect 14866 20038 14882 20055
rect 14740 20021 14782 20038
rect 14622 19974 14782 20021
rect 14840 20021 14882 20038
rect 14958 20038 14974 20055
rect 15084 20055 15192 20071
rect 15084 20038 15100 20055
rect 14958 20021 15000 20038
rect 14840 19974 15000 20021
rect 15058 20021 15100 20038
rect 15176 20038 15192 20055
rect 15302 20055 15410 20071
rect 15302 20038 15318 20055
rect 15176 20021 15218 20038
rect 15058 19974 15218 20021
rect 15276 20021 15318 20038
rect 15394 20038 15410 20055
rect 15520 20055 15628 20071
rect 15520 20038 15536 20055
rect 15394 20021 15436 20038
rect 15276 19974 15436 20021
rect 15494 20021 15536 20038
rect 15612 20038 15628 20055
rect 15738 20055 15846 20071
rect 15738 20038 15754 20055
rect 15612 20021 15654 20038
rect 15494 19974 15654 20021
rect 15712 20021 15754 20038
rect 15830 20038 15846 20055
rect 15956 20055 16064 20071
rect 15956 20038 15972 20055
rect 15830 20021 15872 20038
rect 15712 19974 15872 20021
rect 15930 20021 15972 20038
rect 16048 20038 16064 20055
rect 16174 20055 16282 20071
rect 16174 20038 16190 20055
rect 16048 20021 16090 20038
rect 15930 19974 16090 20021
rect 16148 20021 16190 20038
rect 16266 20038 16282 20055
rect 16392 20055 16500 20071
rect 16392 20038 16408 20055
rect 16266 20021 16308 20038
rect 16148 19974 16308 20021
rect 16366 20021 16408 20038
rect 16484 20038 16500 20055
rect 16610 20055 16718 20071
rect 16610 20038 16626 20055
rect 16484 20021 16526 20038
rect 16366 19974 16526 20021
rect 16584 20021 16626 20038
rect 16702 20038 16718 20055
rect 16702 20021 16744 20038
rect 16584 19974 16744 20021
rect 18470 19775 19430 19822
rect 18470 19758 18672 19775
rect 18656 19741 18672 19758
rect 19228 19758 19430 19775
rect 19488 19775 20448 19822
rect 19488 19758 19690 19775
rect 19228 19741 19244 19758
rect 18656 19725 19244 19741
rect 19674 19741 19690 19758
rect 20246 19758 20448 19775
rect 20506 19775 21466 19822
rect 20506 19758 20708 19775
rect 20246 19741 20262 19758
rect 19674 19725 20262 19741
rect 20692 19741 20708 19758
rect 21264 19758 21466 19775
rect 21524 19775 22484 19822
rect 21524 19758 21726 19775
rect 21264 19741 21280 19758
rect 20692 19725 21280 19741
rect 21710 19741 21726 19758
rect 22282 19758 22484 19775
rect 22542 19775 23502 19822
rect 22542 19758 22744 19775
rect 22282 19741 22298 19758
rect 21710 19725 22298 19741
rect 22728 19741 22744 19758
rect 23300 19758 23502 19775
rect 23560 19775 24520 19822
rect 23560 19758 23762 19775
rect 23300 19741 23316 19758
rect 22728 19725 23316 19741
rect 23746 19741 23762 19758
rect 24318 19758 24520 19775
rect 24578 19775 25538 19822
rect 24578 19758 24780 19775
rect 24318 19741 24334 19758
rect 23746 19725 24334 19741
rect 24764 19741 24780 19758
rect 25336 19758 25538 19775
rect 25596 19775 26556 19822
rect 25596 19758 25798 19775
rect 25336 19741 25352 19758
rect 24764 19725 25352 19741
rect 25782 19741 25798 19758
rect 26354 19758 26556 19775
rect 26614 19775 27574 19822
rect 26614 19758 26816 19775
rect 26354 19741 26370 19758
rect 25782 19725 26370 19741
rect 26800 19741 26816 19758
rect 27372 19758 27574 19775
rect 27632 19775 28592 19822
rect 27632 19758 27834 19775
rect 27372 19741 27388 19758
rect 26800 19725 27388 19741
rect 27818 19741 27834 19758
rect 28390 19758 28592 19775
rect 28650 19775 29610 19822
rect 28650 19758 28852 19775
rect 28390 19741 28406 19758
rect 27818 19725 28406 19741
rect 28836 19741 28852 19758
rect 29408 19758 29610 19775
rect 29668 19775 30628 19822
rect 29668 19758 29870 19775
rect 29408 19741 29424 19758
rect 28836 19725 29424 19741
rect 29854 19741 29870 19758
rect 30426 19758 30628 19775
rect 30686 19775 31646 19822
rect 30686 19758 30888 19775
rect 30426 19741 30442 19758
rect 29854 19725 30442 19741
rect 30872 19741 30888 19758
rect 31444 19758 31646 19775
rect 31704 19775 32664 19822
rect 31704 19758 31906 19775
rect 31444 19741 31460 19758
rect 30872 19725 31460 19741
rect 31890 19741 31906 19758
rect 32462 19758 32664 19775
rect 32722 19775 33682 19822
rect 32722 19758 32924 19775
rect 32462 19741 32478 19758
rect 31890 19725 32478 19741
rect 32908 19741 32924 19758
rect 33480 19758 33682 19775
rect 33480 19741 33496 19758
rect 32908 19725 33496 19741
rect 14622 19527 14782 19574
rect 14622 19510 14664 19527
rect 14648 19493 14664 19510
rect 14740 19510 14782 19527
rect 14840 19527 15000 19574
rect 14840 19510 14882 19527
rect 14740 19493 14756 19510
rect 14648 19477 14756 19493
rect 14866 19493 14882 19510
rect 14958 19510 15000 19527
rect 15058 19527 15218 19574
rect 15058 19510 15100 19527
rect 14958 19493 14974 19510
rect 14866 19477 14974 19493
rect 15084 19493 15100 19510
rect 15176 19510 15218 19527
rect 15276 19527 15436 19574
rect 15276 19510 15318 19527
rect 15176 19493 15192 19510
rect 15084 19477 15192 19493
rect 15302 19493 15318 19510
rect 15394 19510 15436 19527
rect 15494 19527 15654 19574
rect 15494 19510 15536 19527
rect 15394 19493 15410 19510
rect 15302 19477 15410 19493
rect 15520 19493 15536 19510
rect 15612 19510 15654 19527
rect 15712 19527 15872 19574
rect 15712 19510 15754 19527
rect 15612 19493 15628 19510
rect 15520 19477 15628 19493
rect 15738 19493 15754 19510
rect 15830 19510 15872 19527
rect 15930 19527 16090 19574
rect 15930 19510 15972 19527
rect 15830 19493 15846 19510
rect 15738 19477 15846 19493
rect 15956 19493 15972 19510
rect 16048 19510 16090 19527
rect 16148 19527 16308 19574
rect 16148 19510 16190 19527
rect 16048 19493 16064 19510
rect 15956 19477 16064 19493
rect 16174 19493 16190 19510
rect 16266 19510 16308 19527
rect 16366 19527 16526 19574
rect 16366 19510 16408 19527
rect 16266 19493 16282 19510
rect 16174 19477 16282 19493
rect 16392 19493 16408 19510
rect 16484 19510 16526 19527
rect 16584 19527 16744 19574
rect 16584 19510 16626 19527
rect 16484 19493 16500 19510
rect 16392 19477 16500 19493
rect 16610 19493 16626 19510
rect 16702 19510 16744 19527
rect 16702 19493 16718 19510
rect 16610 19477 16718 19493
rect 18656 19247 19244 19263
rect 18656 19230 18672 19247
rect 18470 19213 18672 19230
rect 19228 19230 19244 19247
rect 19674 19247 20262 19263
rect 19674 19230 19690 19247
rect 19228 19213 19430 19230
rect 18470 19166 19430 19213
rect 19488 19213 19690 19230
rect 20246 19230 20262 19247
rect 20692 19247 21280 19263
rect 20692 19230 20708 19247
rect 20246 19213 20448 19230
rect 19488 19166 20448 19213
rect 20506 19213 20708 19230
rect 21264 19230 21280 19247
rect 21710 19247 22298 19263
rect 21710 19230 21726 19247
rect 21264 19213 21466 19230
rect 20506 19166 21466 19213
rect 21524 19213 21726 19230
rect 22282 19230 22298 19247
rect 22728 19247 23316 19263
rect 22728 19230 22744 19247
rect 22282 19213 22484 19230
rect 21524 19166 22484 19213
rect 22542 19213 22744 19230
rect 23300 19230 23316 19247
rect 23746 19247 24334 19263
rect 23746 19230 23762 19247
rect 23300 19213 23502 19230
rect 22542 19166 23502 19213
rect 23560 19213 23762 19230
rect 24318 19230 24334 19247
rect 24764 19247 25352 19263
rect 24764 19230 24780 19247
rect 24318 19213 24520 19230
rect 23560 19166 24520 19213
rect 24578 19213 24780 19230
rect 25336 19230 25352 19247
rect 25782 19247 26370 19263
rect 25782 19230 25798 19247
rect 25336 19213 25538 19230
rect 24578 19166 25538 19213
rect 25596 19213 25798 19230
rect 26354 19230 26370 19247
rect 26800 19247 27388 19263
rect 26800 19230 26816 19247
rect 26354 19213 26556 19230
rect 25596 19166 26556 19213
rect 26614 19213 26816 19230
rect 27372 19230 27388 19247
rect 27818 19247 28406 19263
rect 27818 19230 27834 19247
rect 27372 19213 27574 19230
rect 26614 19166 27574 19213
rect 27632 19213 27834 19230
rect 28390 19230 28406 19247
rect 28836 19247 29424 19263
rect 28836 19230 28852 19247
rect 28390 19213 28592 19230
rect 27632 19166 28592 19213
rect 28650 19213 28852 19230
rect 29408 19230 29424 19247
rect 29854 19247 30442 19263
rect 29854 19230 29870 19247
rect 29408 19213 29610 19230
rect 28650 19166 29610 19213
rect 29668 19213 29870 19230
rect 30426 19230 30442 19247
rect 30872 19247 31460 19263
rect 30872 19230 30888 19247
rect 30426 19213 30628 19230
rect 29668 19166 30628 19213
rect 30686 19213 30888 19230
rect 31444 19230 31460 19247
rect 31890 19247 32478 19263
rect 31890 19230 31906 19247
rect 31444 19213 31646 19230
rect 30686 19166 31646 19213
rect 31704 19213 31906 19230
rect 32462 19230 32478 19247
rect 32908 19247 33496 19263
rect 32908 19230 32924 19247
rect 32462 19213 32664 19230
rect 31704 19166 32664 19213
rect 32722 19213 32924 19230
rect 33480 19230 33496 19247
rect 33480 19213 33682 19230
rect 32722 19166 33682 19213
rect 14648 19117 14756 19133
rect 14648 19100 14664 19117
rect 14622 19083 14664 19100
rect 14740 19100 14756 19117
rect 14866 19117 14974 19133
rect 14866 19100 14882 19117
rect 14740 19083 14782 19100
rect 14622 19036 14782 19083
rect 14840 19083 14882 19100
rect 14958 19100 14974 19117
rect 15084 19117 15192 19133
rect 15084 19100 15100 19117
rect 14958 19083 15000 19100
rect 14840 19036 15000 19083
rect 15058 19083 15100 19100
rect 15176 19100 15192 19117
rect 15302 19117 15410 19133
rect 15302 19100 15318 19117
rect 15176 19083 15218 19100
rect 15058 19036 15218 19083
rect 15276 19083 15318 19100
rect 15394 19100 15410 19117
rect 15520 19117 15628 19133
rect 15520 19100 15536 19117
rect 15394 19083 15436 19100
rect 15276 19036 15436 19083
rect 15494 19083 15536 19100
rect 15612 19100 15628 19117
rect 15738 19117 15846 19133
rect 15738 19100 15754 19117
rect 15612 19083 15654 19100
rect 15494 19036 15654 19083
rect 15712 19083 15754 19100
rect 15830 19100 15846 19117
rect 15956 19117 16064 19133
rect 15956 19100 15972 19117
rect 15830 19083 15872 19100
rect 15712 19036 15872 19083
rect 15930 19083 15972 19100
rect 16048 19100 16064 19117
rect 16174 19117 16282 19133
rect 16174 19100 16190 19117
rect 16048 19083 16090 19100
rect 15930 19036 16090 19083
rect 16148 19083 16190 19100
rect 16266 19100 16282 19117
rect 16392 19117 16500 19133
rect 16392 19100 16408 19117
rect 16266 19083 16308 19100
rect 16148 19036 16308 19083
rect 16366 19083 16408 19100
rect 16484 19100 16500 19117
rect 16610 19117 16718 19133
rect 16610 19100 16626 19117
rect 16484 19083 16526 19100
rect 16366 19036 16526 19083
rect 16584 19083 16626 19100
rect 16702 19100 16718 19117
rect 16702 19083 16744 19100
rect 16584 19036 16744 19083
rect 14622 18589 14782 18636
rect 14622 18572 14664 18589
rect 14648 18555 14664 18572
rect 14740 18572 14782 18589
rect 14840 18589 15000 18636
rect 14840 18572 14882 18589
rect 14740 18555 14756 18572
rect 14648 18539 14756 18555
rect 14866 18555 14882 18572
rect 14958 18572 15000 18589
rect 15058 18589 15218 18636
rect 15058 18572 15100 18589
rect 14958 18555 14974 18572
rect 14866 18539 14974 18555
rect 15084 18555 15100 18572
rect 15176 18572 15218 18589
rect 15276 18589 15436 18636
rect 15276 18572 15318 18589
rect 15176 18555 15192 18572
rect 15084 18539 15192 18555
rect 15302 18555 15318 18572
rect 15394 18572 15436 18589
rect 15494 18589 15654 18636
rect 15494 18572 15536 18589
rect 15394 18555 15410 18572
rect 15302 18539 15410 18555
rect 15520 18555 15536 18572
rect 15612 18572 15654 18589
rect 15712 18589 15872 18636
rect 15712 18572 15754 18589
rect 15612 18555 15628 18572
rect 15520 18539 15628 18555
rect 15738 18555 15754 18572
rect 15830 18572 15872 18589
rect 15930 18589 16090 18636
rect 15930 18572 15972 18589
rect 15830 18555 15846 18572
rect 15738 18539 15846 18555
rect 15956 18555 15972 18572
rect 16048 18572 16090 18589
rect 16148 18589 16308 18636
rect 16148 18572 16190 18589
rect 16048 18555 16064 18572
rect 15956 18539 16064 18555
rect 16174 18555 16190 18572
rect 16266 18572 16308 18589
rect 16366 18589 16526 18636
rect 16366 18572 16408 18589
rect 16266 18555 16282 18572
rect 16174 18539 16282 18555
rect 16392 18555 16408 18572
rect 16484 18572 16526 18589
rect 16584 18589 16744 18636
rect 16584 18572 16626 18589
rect 16484 18555 16500 18572
rect 16392 18539 16500 18555
rect 16610 18555 16626 18572
rect 16702 18572 16744 18589
rect 16702 18555 16718 18572
rect 16610 18539 16718 18555
rect 18470 18519 19430 18566
rect 18470 18502 18672 18519
rect 18656 18485 18672 18502
rect 19228 18502 19430 18519
rect 19488 18519 20448 18566
rect 19488 18502 19690 18519
rect 19228 18485 19244 18502
rect 18656 18469 19244 18485
rect 19674 18485 19690 18502
rect 20246 18502 20448 18519
rect 20506 18519 21466 18566
rect 20506 18502 20708 18519
rect 20246 18485 20262 18502
rect 19674 18469 20262 18485
rect 20692 18485 20708 18502
rect 21264 18502 21466 18519
rect 21524 18519 22484 18566
rect 21524 18502 21726 18519
rect 21264 18485 21280 18502
rect 20692 18469 21280 18485
rect 21710 18485 21726 18502
rect 22282 18502 22484 18519
rect 22542 18519 23502 18566
rect 22542 18502 22744 18519
rect 22282 18485 22298 18502
rect 21710 18469 22298 18485
rect 22728 18485 22744 18502
rect 23300 18502 23502 18519
rect 23560 18519 24520 18566
rect 23560 18502 23762 18519
rect 23300 18485 23316 18502
rect 22728 18469 23316 18485
rect 23746 18485 23762 18502
rect 24318 18502 24520 18519
rect 24578 18519 25538 18566
rect 24578 18502 24780 18519
rect 24318 18485 24334 18502
rect 23746 18469 24334 18485
rect 24764 18485 24780 18502
rect 25336 18502 25538 18519
rect 25596 18519 26556 18566
rect 25596 18502 25798 18519
rect 25336 18485 25352 18502
rect 24764 18469 25352 18485
rect 25782 18485 25798 18502
rect 26354 18502 26556 18519
rect 26614 18519 27574 18566
rect 26614 18502 26816 18519
rect 26354 18485 26370 18502
rect 25782 18469 26370 18485
rect 26800 18485 26816 18502
rect 27372 18502 27574 18519
rect 27632 18519 28592 18566
rect 27632 18502 27834 18519
rect 27372 18485 27388 18502
rect 26800 18469 27388 18485
rect 27818 18485 27834 18502
rect 28390 18502 28592 18519
rect 28650 18519 29610 18566
rect 28650 18502 28852 18519
rect 28390 18485 28406 18502
rect 27818 18469 28406 18485
rect 28836 18485 28852 18502
rect 29408 18502 29610 18519
rect 29668 18519 30628 18566
rect 29668 18502 29870 18519
rect 29408 18485 29424 18502
rect 28836 18469 29424 18485
rect 29854 18485 29870 18502
rect 30426 18502 30628 18519
rect 30686 18519 31646 18566
rect 30686 18502 30888 18519
rect 30426 18485 30442 18502
rect 29854 18469 30442 18485
rect 30872 18485 30888 18502
rect 31444 18502 31646 18519
rect 31704 18519 32664 18566
rect 31704 18502 31906 18519
rect 31444 18485 31460 18502
rect 30872 18469 31460 18485
rect 31890 18485 31906 18502
rect 32462 18502 32664 18519
rect 32722 18519 33682 18566
rect 32722 18502 32924 18519
rect 32462 18485 32478 18502
rect 31890 18469 32478 18485
rect 32908 18485 32924 18502
rect 33480 18502 33682 18519
rect 33480 18485 33496 18502
rect 32908 18469 33496 18485
rect 47458 25309 47590 25325
rect 47458 25292 47474 25309
rect 47424 25275 47474 25292
rect 47574 25292 47590 25309
rect 47716 25309 47848 25325
rect 47716 25292 47732 25309
rect 47574 25275 47624 25292
rect 47424 25228 47624 25275
rect 47682 25275 47732 25292
rect 47832 25292 47848 25309
rect 47974 25309 48106 25325
rect 47974 25292 47990 25309
rect 47832 25275 47882 25292
rect 47682 25228 47882 25275
rect 47940 25275 47990 25292
rect 48090 25292 48106 25309
rect 48232 25309 48364 25325
rect 48232 25292 48248 25309
rect 48090 25275 48140 25292
rect 47940 25228 48140 25275
rect 48198 25275 48248 25292
rect 48348 25292 48364 25309
rect 48490 25309 48622 25325
rect 48490 25292 48506 25309
rect 48348 25275 48398 25292
rect 48198 25228 48398 25275
rect 48456 25275 48506 25292
rect 48606 25292 48622 25309
rect 48748 25309 48880 25325
rect 48748 25292 48764 25309
rect 48606 25275 48656 25292
rect 48456 25228 48656 25275
rect 48714 25275 48764 25292
rect 48864 25292 48880 25309
rect 48864 25275 48914 25292
rect 48714 25228 48914 25275
rect 47424 24781 47624 24828
rect 47424 24764 47474 24781
rect 47458 24747 47474 24764
rect 47574 24764 47624 24781
rect 47682 24781 47882 24828
rect 47682 24764 47732 24781
rect 47574 24747 47590 24764
rect 47458 24731 47590 24747
rect 47716 24747 47732 24764
rect 47832 24764 47882 24781
rect 47940 24781 48140 24828
rect 47940 24764 47990 24781
rect 47832 24747 47848 24764
rect 47716 24731 47848 24747
rect 47974 24747 47990 24764
rect 48090 24764 48140 24781
rect 48198 24781 48398 24828
rect 48198 24764 48248 24781
rect 48090 24747 48106 24764
rect 47974 24731 48106 24747
rect 48232 24747 48248 24764
rect 48348 24764 48398 24781
rect 48456 24781 48656 24828
rect 48456 24764 48506 24781
rect 48348 24747 48364 24764
rect 48232 24731 48364 24747
rect 48490 24747 48506 24764
rect 48606 24764 48656 24781
rect 48714 24781 48914 24828
rect 48714 24764 48764 24781
rect 48606 24747 48622 24764
rect 48490 24731 48622 24747
rect 48748 24747 48764 24764
rect 48864 24764 48914 24781
rect 48864 24747 48880 24764
rect 48748 24731 48880 24747
rect 49274 24845 49304 24871
rect 49274 24613 49304 24645
rect 49274 24597 49360 24613
rect 49274 24563 49310 24597
rect 49344 24563 49360 24597
rect 49274 24547 49360 24563
rect 49274 24525 49304 24547
rect 47458 24376 47590 24392
rect 47458 24359 47474 24376
rect 47424 24342 47474 24359
rect 47574 24359 47590 24376
rect 47716 24376 47848 24392
rect 47716 24359 47732 24376
rect 47574 24342 47624 24359
rect 47424 24304 47624 24342
rect 47682 24342 47732 24359
rect 47832 24359 47848 24376
rect 47974 24376 48106 24392
rect 47974 24359 47990 24376
rect 47832 24342 47882 24359
rect 47682 24304 47882 24342
rect 47940 24342 47990 24359
rect 48090 24359 48106 24376
rect 48232 24376 48364 24392
rect 48232 24359 48248 24376
rect 48090 24342 48140 24359
rect 47940 24304 48140 24342
rect 48198 24342 48248 24359
rect 48348 24359 48364 24376
rect 48490 24376 48622 24392
rect 48490 24359 48506 24376
rect 48348 24342 48398 24359
rect 48198 24304 48398 24342
rect 48456 24342 48506 24359
rect 48606 24359 48622 24376
rect 48748 24376 48880 24392
rect 48748 24359 48764 24376
rect 48606 24342 48656 24359
rect 48456 24304 48656 24342
rect 48714 24342 48764 24359
rect 48864 24359 48880 24376
rect 48864 24342 48914 24359
rect 48714 24304 48914 24342
rect 47424 24066 47624 24104
rect 47424 24049 47474 24066
rect 47458 24032 47474 24049
rect 47574 24049 47624 24066
rect 47682 24066 47882 24104
rect 47682 24049 47732 24066
rect 47574 24032 47590 24049
rect 47458 24016 47590 24032
rect 47716 24032 47732 24049
rect 47832 24049 47882 24066
rect 47940 24066 48140 24104
rect 47940 24049 47990 24066
rect 47832 24032 47848 24049
rect 47716 24016 47848 24032
rect 47974 24032 47990 24049
rect 48090 24049 48140 24066
rect 48198 24066 48398 24104
rect 48198 24049 48248 24066
rect 48090 24032 48106 24049
rect 47974 24016 48106 24032
rect 48232 24032 48248 24049
rect 48348 24049 48398 24066
rect 48456 24066 48656 24104
rect 48456 24049 48506 24066
rect 48348 24032 48364 24049
rect 48232 24016 48364 24032
rect 48490 24032 48506 24049
rect 48606 24049 48656 24066
rect 48714 24066 48914 24104
rect 48714 24049 48764 24066
rect 48606 24032 48622 24049
rect 48490 24016 48622 24032
rect 48748 24032 48764 24049
rect 48864 24049 48914 24066
rect 48864 24032 48880 24049
rect 48748 24016 48880 24032
rect 49274 24369 49304 24395
rect 47458 23309 47590 23325
rect 47458 23292 47474 23309
rect 47424 23275 47474 23292
rect 47574 23292 47590 23309
rect 47716 23309 47848 23325
rect 47716 23292 47732 23309
rect 47574 23275 47624 23292
rect 47424 23228 47624 23275
rect 47682 23275 47732 23292
rect 47832 23292 47848 23309
rect 47974 23309 48106 23325
rect 47974 23292 47990 23309
rect 47832 23275 47882 23292
rect 47682 23228 47882 23275
rect 47940 23275 47990 23292
rect 48090 23292 48106 23309
rect 48232 23309 48364 23325
rect 48232 23292 48248 23309
rect 48090 23275 48140 23292
rect 47940 23228 48140 23275
rect 48198 23275 48248 23292
rect 48348 23292 48364 23309
rect 48490 23309 48622 23325
rect 48490 23292 48506 23309
rect 48348 23275 48398 23292
rect 48198 23228 48398 23275
rect 48456 23275 48506 23292
rect 48606 23292 48622 23309
rect 48748 23309 48880 23325
rect 48748 23292 48764 23309
rect 48606 23275 48656 23292
rect 48456 23228 48656 23275
rect 48714 23275 48764 23292
rect 48864 23292 48880 23309
rect 48864 23275 48914 23292
rect 48714 23228 48914 23275
rect 47424 22781 47624 22828
rect 47424 22764 47474 22781
rect 47458 22747 47474 22764
rect 47574 22764 47624 22781
rect 47682 22781 47882 22828
rect 47682 22764 47732 22781
rect 47574 22747 47590 22764
rect 47458 22731 47590 22747
rect 47716 22747 47732 22764
rect 47832 22764 47882 22781
rect 47940 22781 48140 22828
rect 47940 22764 47990 22781
rect 47832 22747 47848 22764
rect 47716 22731 47848 22747
rect 47974 22747 47990 22764
rect 48090 22764 48140 22781
rect 48198 22781 48398 22828
rect 48198 22764 48248 22781
rect 48090 22747 48106 22764
rect 47974 22731 48106 22747
rect 48232 22747 48248 22764
rect 48348 22764 48398 22781
rect 48456 22781 48656 22828
rect 48456 22764 48506 22781
rect 48348 22747 48364 22764
rect 48232 22731 48364 22747
rect 48490 22747 48506 22764
rect 48606 22764 48656 22781
rect 48714 22781 48914 22828
rect 48714 22764 48764 22781
rect 48606 22747 48622 22764
rect 48490 22731 48622 22747
rect 48748 22747 48764 22764
rect 48864 22764 48914 22781
rect 48864 22747 48880 22764
rect 48748 22731 48880 22747
rect 49274 22845 49304 22871
rect 49274 22613 49304 22645
rect 49274 22597 49360 22613
rect 49274 22563 49310 22597
rect 49344 22563 49360 22597
rect 49274 22547 49360 22563
rect 49274 22525 49304 22547
rect 47458 22376 47590 22392
rect 47458 22359 47474 22376
rect 47424 22342 47474 22359
rect 47574 22359 47590 22376
rect 47716 22376 47848 22392
rect 47716 22359 47732 22376
rect 47574 22342 47624 22359
rect 47424 22304 47624 22342
rect 47682 22342 47732 22359
rect 47832 22359 47848 22376
rect 47974 22376 48106 22392
rect 47974 22359 47990 22376
rect 47832 22342 47882 22359
rect 47682 22304 47882 22342
rect 47940 22342 47990 22359
rect 48090 22359 48106 22376
rect 48232 22376 48364 22392
rect 48232 22359 48248 22376
rect 48090 22342 48140 22359
rect 47940 22304 48140 22342
rect 48198 22342 48248 22359
rect 48348 22359 48364 22376
rect 48490 22376 48622 22392
rect 48490 22359 48506 22376
rect 48348 22342 48398 22359
rect 48198 22304 48398 22342
rect 48456 22342 48506 22359
rect 48606 22359 48622 22376
rect 48748 22376 48880 22392
rect 48748 22359 48764 22376
rect 48606 22342 48656 22359
rect 48456 22304 48656 22342
rect 48714 22342 48764 22359
rect 48864 22359 48880 22376
rect 48864 22342 48914 22359
rect 48714 22304 48914 22342
rect 47424 22066 47624 22104
rect 47424 22049 47474 22066
rect 47458 22032 47474 22049
rect 47574 22049 47624 22066
rect 47682 22066 47882 22104
rect 47682 22049 47732 22066
rect 47574 22032 47590 22049
rect 47458 22016 47590 22032
rect 47716 22032 47732 22049
rect 47832 22049 47882 22066
rect 47940 22066 48140 22104
rect 47940 22049 47990 22066
rect 47832 22032 47848 22049
rect 47716 22016 47848 22032
rect 47974 22032 47990 22049
rect 48090 22049 48140 22066
rect 48198 22066 48398 22104
rect 48198 22049 48248 22066
rect 48090 22032 48106 22049
rect 47974 22016 48106 22032
rect 48232 22032 48248 22049
rect 48348 22049 48398 22066
rect 48456 22066 48656 22104
rect 48456 22049 48506 22066
rect 48348 22032 48364 22049
rect 48232 22016 48364 22032
rect 48490 22032 48506 22049
rect 48606 22049 48656 22066
rect 48714 22066 48914 22104
rect 48714 22049 48764 22066
rect 48606 22032 48622 22049
rect 48490 22016 48622 22032
rect 48748 22032 48764 22049
rect 48864 22049 48914 22066
rect 48864 22032 48880 22049
rect 48748 22016 48880 22032
rect 49274 22369 49304 22395
rect 71670 27061 72258 27077
rect 71670 27044 71686 27061
rect 71484 27027 71686 27044
rect 72242 27044 72258 27061
rect 72688 27061 73276 27077
rect 72688 27044 72704 27061
rect 72242 27027 72444 27044
rect 71484 26980 72444 27027
rect 72502 27027 72704 27044
rect 73260 27044 73276 27061
rect 73706 27061 74294 27077
rect 73706 27044 73722 27061
rect 73260 27027 73462 27044
rect 72502 26980 73462 27027
rect 73520 27027 73722 27044
rect 74278 27044 74294 27061
rect 74724 27061 75312 27077
rect 74724 27044 74740 27061
rect 74278 27027 74480 27044
rect 73520 26980 74480 27027
rect 74538 27027 74740 27044
rect 75296 27044 75312 27061
rect 75742 27061 76330 27077
rect 75742 27044 75758 27061
rect 75296 27027 75498 27044
rect 74538 26980 75498 27027
rect 75556 27027 75758 27044
rect 76314 27044 76330 27061
rect 76760 27061 77348 27077
rect 76760 27044 76776 27061
rect 76314 27027 76516 27044
rect 75556 26980 76516 27027
rect 76574 27027 76776 27044
rect 77332 27044 77348 27061
rect 77778 27061 78366 27077
rect 77778 27044 77794 27061
rect 77332 27027 77534 27044
rect 76574 26980 77534 27027
rect 77592 27027 77794 27044
rect 78350 27044 78366 27061
rect 78796 27061 79384 27077
rect 78796 27044 78812 27061
rect 78350 27027 78552 27044
rect 77592 26980 78552 27027
rect 78610 27027 78812 27044
rect 79368 27044 79384 27061
rect 79814 27061 80402 27077
rect 79814 27044 79830 27061
rect 79368 27027 79570 27044
rect 78610 26980 79570 27027
rect 79628 27027 79830 27044
rect 80386 27044 80402 27061
rect 80832 27061 81420 27077
rect 80832 27044 80848 27061
rect 80386 27027 80588 27044
rect 79628 26980 80588 27027
rect 80646 27027 80848 27044
rect 81404 27044 81420 27061
rect 81850 27061 82438 27077
rect 81850 27044 81866 27061
rect 81404 27027 81606 27044
rect 80646 26980 81606 27027
rect 81664 27027 81866 27044
rect 82422 27044 82438 27061
rect 82868 27061 83456 27077
rect 82868 27044 82884 27061
rect 82422 27027 82624 27044
rect 81664 26980 82624 27027
rect 82682 27027 82884 27044
rect 83440 27044 83456 27061
rect 83886 27061 84474 27077
rect 83886 27044 83902 27061
rect 83440 27027 83642 27044
rect 82682 26980 83642 27027
rect 83700 27027 83902 27044
rect 84458 27044 84474 27061
rect 84904 27061 85492 27077
rect 84904 27044 84920 27061
rect 84458 27027 84660 27044
rect 83700 26980 84660 27027
rect 84718 27027 84920 27044
rect 85476 27044 85492 27061
rect 85922 27061 86510 27077
rect 85922 27044 85938 27061
rect 85476 27027 85678 27044
rect 84718 26980 85678 27027
rect 85736 27027 85938 27044
rect 86494 27044 86510 27061
rect 86940 27061 87528 27077
rect 86940 27044 86956 27061
rect 86494 27027 86696 27044
rect 85736 26980 86696 27027
rect 86754 27027 86956 27044
rect 87512 27044 87528 27061
rect 87512 27027 87714 27044
rect 86754 26980 87714 27027
rect 71484 26333 72444 26380
rect 71484 26316 71686 26333
rect 71670 26299 71686 26316
rect 72242 26316 72444 26333
rect 72502 26333 73462 26380
rect 72502 26316 72704 26333
rect 72242 26299 72258 26316
rect 71670 26283 72258 26299
rect 72688 26299 72704 26316
rect 73260 26316 73462 26333
rect 73520 26333 74480 26380
rect 73520 26316 73722 26333
rect 73260 26299 73276 26316
rect 72688 26283 73276 26299
rect 73706 26299 73722 26316
rect 74278 26316 74480 26333
rect 74538 26333 75498 26380
rect 74538 26316 74740 26333
rect 74278 26299 74294 26316
rect 73706 26283 74294 26299
rect 74724 26299 74740 26316
rect 75296 26316 75498 26333
rect 75556 26333 76516 26380
rect 75556 26316 75758 26333
rect 75296 26299 75312 26316
rect 74724 26283 75312 26299
rect 75742 26299 75758 26316
rect 76314 26316 76516 26333
rect 76574 26333 77534 26380
rect 76574 26316 76776 26333
rect 76314 26299 76330 26316
rect 75742 26283 76330 26299
rect 76760 26299 76776 26316
rect 77332 26316 77534 26333
rect 77592 26333 78552 26380
rect 77592 26316 77794 26333
rect 77332 26299 77348 26316
rect 76760 26283 77348 26299
rect 77778 26299 77794 26316
rect 78350 26316 78552 26333
rect 78610 26333 79570 26380
rect 78610 26316 78812 26333
rect 78350 26299 78366 26316
rect 77778 26283 78366 26299
rect 78796 26299 78812 26316
rect 79368 26316 79570 26333
rect 79628 26333 80588 26380
rect 79628 26316 79830 26333
rect 79368 26299 79384 26316
rect 78796 26283 79384 26299
rect 79814 26299 79830 26316
rect 80386 26316 80588 26333
rect 80646 26333 81606 26380
rect 80646 26316 80848 26333
rect 80386 26299 80402 26316
rect 79814 26283 80402 26299
rect 80832 26299 80848 26316
rect 81404 26316 81606 26333
rect 81664 26333 82624 26380
rect 81664 26316 81866 26333
rect 81404 26299 81420 26316
rect 80832 26283 81420 26299
rect 81850 26299 81866 26316
rect 82422 26316 82624 26333
rect 82682 26333 83642 26380
rect 82682 26316 82884 26333
rect 82422 26299 82438 26316
rect 81850 26283 82438 26299
rect 82868 26299 82884 26316
rect 83440 26316 83642 26333
rect 83700 26333 84660 26380
rect 83700 26316 83902 26333
rect 83440 26299 83456 26316
rect 82868 26283 83456 26299
rect 83886 26299 83902 26316
rect 84458 26316 84660 26333
rect 84718 26333 85678 26380
rect 84718 26316 84920 26333
rect 84458 26299 84474 26316
rect 83886 26283 84474 26299
rect 84904 26299 84920 26316
rect 85476 26316 85678 26333
rect 85736 26333 86696 26380
rect 85736 26316 85938 26333
rect 85476 26299 85492 26316
rect 84904 26283 85492 26299
rect 85922 26299 85938 26316
rect 86494 26316 86696 26333
rect 86754 26333 87714 26380
rect 86754 26316 86956 26333
rect 86494 26299 86510 26316
rect 85922 26283 86510 26299
rect 86940 26299 86956 26316
rect 87512 26316 87714 26333
rect 87512 26299 87528 26316
rect 86940 26283 87528 26299
rect 71670 25925 72258 25941
rect 71670 25908 71686 25925
rect 71484 25891 71686 25908
rect 72242 25908 72258 25925
rect 72688 25925 73276 25941
rect 72688 25908 72704 25925
rect 72242 25891 72444 25908
rect 71484 25844 72444 25891
rect 72502 25891 72704 25908
rect 73260 25908 73276 25925
rect 73706 25925 74294 25941
rect 73706 25908 73722 25925
rect 73260 25891 73462 25908
rect 72502 25844 73462 25891
rect 73520 25891 73722 25908
rect 74278 25908 74294 25925
rect 74724 25925 75312 25941
rect 74724 25908 74740 25925
rect 74278 25891 74480 25908
rect 73520 25844 74480 25891
rect 74538 25891 74740 25908
rect 75296 25908 75312 25925
rect 75742 25925 76330 25941
rect 75742 25908 75758 25925
rect 75296 25891 75498 25908
rect 74538 25844 75498 25891
rect 75556 25891 75758 25908
rect 76314 25908 76330 25925
rect 76760 25925 77348 25941
rect 76760 25908 76776 25925
rect 76314 25891 76516 25908
rect 75556 25844 76516 25891
rect 76574 25891 76776 25908
rect 77332 25908 77348 25925
rect 77778 25925 78366 25941
rect 77778 25908 77794 25925
rect 77332 25891 77534 25908
rect 76574 25844 77534 25891
rect 77592 25891 77794 25908
rect 78350 25908 78366 25925
rect 78796 25925 79384 25941
rect 78796 25908 78812 25925
rect 78350 25891 78552 25908
rect 77592 25844 78552 25891
rect 78610 25891 78812 25908
rect 79368 25908 79384 25925
rect 79814 25925 80402 25941
rect 79814 25908 79830 25925
rect 79368 25891 79570 25908
rect 78610 25844 79570 25891
rect 79628 25891 79830 25908
rect 80386 25908 80402 25925
rect 80832 25925 81420 25941
rect 80832 25908 80848 25925
rect 80386 25891 80588 25908
rect 79628 25844 80588 25891
rect 80646 25891 80848 25908
rect 81404 25908 81420 25925
rect 81850 25925 82438 25941
rect 81850 25908 81866 25925
rect 81404 25891 81606 25908
rect 80646 25844 81606 25891
rect 81664 25891 81866 25908
rect 82422 25908 82438 25925
rect 82868 25925 83456 25941
rect 82868 25908 82884 25925
rect 82422 25891 82624 25908
rect 81664 25844 82624 25891
rect 82682 25891 82884 25908
rect 83440 25908 83456 25925
rect 83886 25925 84474 25941
rect 83886 25908 83902 25925
rect 83440 25891 83642 25908
rect 82682 25844 83642 25891
rect 83700 25891 83902 25908
rect 84458 25908 84474 25925
rect 84904 25925 85492 25941
rect 84904 25908 84920 25925
rect 84458 25891 84660 25908
rect 83700 25844 84660 25891
rect 84718 25891 84920 25908
rect 85476 25908 85492 25925
rect 85922 25925 86510 25941
rect 85922 25908 85938 25925
rect 85476 25891 85678 25908
rect 84718 25844 85678 25891
rect 85736 25891 85938 25908
rect 86494 25908 86510 25925
rect 86940 25925 87528 25941
rect 86940 25908 86956 25925
rect 86494 25891 86696 25908
rect 85736 25844 86696 25891
rect 86754 25891 86956 25908
rect 87512 25908 87528 25925
rect 87512 25891 87714 25908
rect 86754 25844 87714 25891
rect 71484 25197 72444 25244
rect 71484 25180 71686 25197
rect 71670 25163 71686 25180
rect 72242 25180 72444 25197
rect 72502 25197 73462 25244
rect 72502 25180 72704 25197
rect 72242 25163 72258 25180
rect 71670 25147 72258 25163
rect 72688 25163 72704 25180
rect 73260 25180 73462 25197
rect 73520 25197 74480 25244
rect 73520 25180 73722 25197
rect 73260 25163 73276 25180
rect 72688 25147 73276 25163
rect 73706 25163 73722 25180
rect 74278 25180 74480 25197
rect 74538 25197 75498 25244
rect 74538 25180 74740 25197
rect 74278 25163 74294 25180
rect 73706 25147 74294 25163
rect 74724 25163 74740 25180
rect 75296 25180 75498 25197
rect 75556 25197 76516 25244
rect 75556 25180 75758 25197
rect 75296 25163 75312 25180
rect 74724 25147 75312 25163
rect 75742 25163 75758 25180
rect 76314 25180 76516 25197
rect 76574 25197 77534 25244
rect 76574 25180 76776 25197
rect 76314 25163 76330 25180
rect 75742 25147 76330 25163
rect 76760 25163 76776 25180
rect 77332 25180 77534 25197
rect 77592 25197 78552 25244
rect 77592 25180 77794 25197
rect 77332 25163 77348 25180
rect 76760 25147 77348 25163
rect 77778 25163 77794 25180
rect 78350 25180 78552 25197
rect 78610 25197 79570 25244
rect 78610 25180 78812 25197
rect 78350 25163 78366 25180
rect 77778 25147 78366 25163
rect 78796 25163 78812 25180
rect 79368 25180 79570 25197
rect 79628 25197 80588 25244
rect 79628 25180 79830 25197
rect 79368 25163 79384 25180
rect 78796 25147 79384 25163
rect 79814 25163 79830 25180
rect 80386 25180 80588 25197
rect 80646 25197 81606 25244
rect 80646 25180 80848 25197
rect 80386 25163 80402 25180
rect 79814 25147 80402 25163
rect 80832 25163 80848 25180
rect 81404 25180 81606 25197
rect 81664 25197 82624 25244
rect 81664 25180 81866 25197
rect 81404 25163 81420 25180
rect 80832 25147 81420 25163
rect 81850 25163 81866 25180
rect 82422 25180 82624 25197
rect 82682 25197 83642 25244
rect 82682 25180 82884 25197
rect 82422 25163 82438 25180
rect 81850 25147 82438 25163
rect 82868 25163 82884 25180
rect 83440 25180 83642 25197
rect 83700 25197 84660 25244
rect 83700 25180 83902 25197
rect 83440 25163 83456 25180
rect 82868 25147 83456 25163
rect 83886 25163 83902 25180
rect 84458 25180 84660 25197
rect 84718 25197 85678 25244
rect 84718 25180 84920 25197
rect 84458 25163 84474 25180
rect 83886 25147 84474 25163
rect 84904 25163 84920 25180
rect 85476 25180 85678 25197
rect 85736 25197 86696 25244
rect 85736 25180 85938 25197
rect 85476 25163 85492 25180
rect 84904 25147 85492 25163
rect 85922 25163 85938 25180
rect 86494 25180 86696 25197
rect 86754 25197 87714 25244
rect 86754 25180 86956 25197
rect 86494 25163 86510 25180
rect 85922 25147 86510 25163
rect 86940 25163 86956 25180
rect 87512 25180 87714 25197
rect 87512 25163 87528 25180
rect 86940 25147 87528 25163
rect 71670 24789 72258 24805
rect 71670 24772 71686 24789
rect 71484 24755 71686 24772
rect 72242 24772 72258 24789
rect 72688 24789 73276 24805
rect 72688 24772 72704 24789
rect 72242 24755 72444 24772
rect 71484 24708 72444 24755
rect 72502 24755 72704 24772
rect 73260 24772 73276 24789
rect 73706 24789 74294 24805
rect 73706 24772 73722 24789
rect 73260 24755 73462 24772
rect 72502 24708 73462 24755
rect 73520 24755 73722 24772
rect 74278 24772 74294 24789
rect 74724 24789 75312 24805
rect 74724 24772 74740 24789
rect 74278 24755 74480 24772
rect 73520 24708 74480 24755
rect 74538 24755 74740 24772
rect 75296 24772 75312 24789
rect 75742 24789 76330 24805
rect 75742 24772 75758 24789
rect 75296 24755 75498 24772
rect 74538 24708 75498 24755
rect 75556 24755 75758 24772
rect 76314 24772 76330 24789
rect 76760 24789 77348 24805
rect 76760 24772 76776 24789
rect 76314 24755 76516 24772
rect 75556 24708 76516 24755
rect 76574 24755 76776 24772
rect 77332 24772 77348 24789
rect 77778 24789 78366 24805
rect 77778 24772 77794 24789
rect 77332 24755 77534 24772
rect 76574 24708 77534 24755
rect 77592 24755 77794 24772
rect 78350 24772 78366 24789
rect 78796 24789 79384 24805
rect 78796 24772 78812 24789
rect 78350 24755 78552 24772
rect 77592 24708 78552 24755
rect 78610 24755 78812 24772
rect 79368 24772 79384 24789
rect 79814 24789 80402 24805
rect 79814 24772 79830 24789
rect 79368 24755 79570 24772
rect 78610 24708 79570 24755
rect 79628 24755 79830 24772
rect 80386 24772 80402 24789
rect 80832 24789 81420 24805
rect 80832 24772 80848 24789
rect 80386 24755 80588 24772
rect 79628 24708 80588 24755
rect 80646 24755 80848 24772
rect 81404 24772 81420 24789
rect 81850 24789 82438 24805
rect 81850 24772 81866 24789
rect 81404 24755 81606 24772
rect 80646 24708 81606 24755
rect 81664 24755 81866 24772
rect 82422 24772 82438 24789
rect 82868 24789 83456 24805
rect 82868 24772 82884 24789
rect 82422 24755 82624 24772
rect 81664 24708 82624 24755
rect 82682 24755 82884 24772
rect 83440 24772 83456 24789
rect 83886 24789 84474 24805
rect 83886 24772 83902 24789
rect 83440 24755 83642 24772
rect 82682 24708 83642 24755
rect 83700 24755 83902 24772
rect 84458 24772 84474 24789
rect 84904 24789 85492 24805
rect 84904 24772 84920 24789
rect 84458 24755 84660 24772
rect 83700 24708 84660 24755
rect 84718 24755 84920 24772
rect 85476 24772 85492 24789
rect 85922 24789 86510 24805
rect 85922 24772 85938 24789
rect 85476 24755 85678 24772
rect 84718 24708 85678 24755
rect 85736 24755 85938 24772
rect 86494 24772 86510 24789
rect 86940 24789 87528 24805
rect 86940 24772 86956 24789
rect 86494 24755 86696 24772
rect 85736 24708 86696 24755
rect 86754 24755 86956 24772
rect 87512 24772 87528 24789
rect 87512 24755 87714 24772
rect 86754 24708 87714 24755
rect 71484 24061 72444 24108
rect 71484 24044 71686 24061
rect 71670 24027 71686 24044
rect 72242 24044 72444 24061
rect 72502 24061 73462 24108
rect 72502 24044 72704 24061
rect 72242 24027 72258 24044
rect 71670 24011 72258 24027
rect 72688 24027 72704 24044
rect 73260 24044 73462 24061
rect 73520 24061 74480 24108
rect 73520 24044 73722 24061
rect 73260 24027 73276 24044
rect 72688 24011 73276 24027
rect 73706 24027 73722 24044
rect 74278 24044 74480 24061
rect 74538 24061 75498 24108
rect 74538 24044 74740 24061
rect 74278 24027 74294 24044
rect 73706 24011 74294 24027
rect 74724 24027 74740 24044
rect 75296 24044 75498 24061
rect 75556 24061 76516 24108
rect 75556 24044 75758 24061
rect 75296 24027 75312 24044
rect 74724 24011 75312 24027
rect 75742 24027 75758 24044
rect 76314 24044 76516 24061
rect 76574 24061 77534 24108
rect 76574 24044 76776 24061
rect 76314 24027 76330 24044
rect 75742 24011 76330 24027
rect 76760 24027 76776 24044
rect 77332 24044 77534 24061
rect 77592 24061 78552 24108
rect 77592 24044 77794 24061
rect 77332 24027 77348 24044
rect 76760 24011 77348 24027
rect 77778 24027 77794 24044
rect 78350 24044 78552 24061
rect 78610 24061 79570 24108
rect 78610 24044 78812 24061
rect 78350 24027 78366 24044
rect 77778 24011 78366 24027
rect 78796 24027 78812 24044
rect 79368 24044 79570 24061
rect 79628 24061 80588 24108
rect 79628 24044 79830 24061
rect 79368 24027 79384 24044
rect 78796 24011 79384 24027
rect 79814 24027 79830 24044
rect 80386 24044 80588 24061
rect 80646 24061 81606 24108
rect 80646 24044 80848 24061
rect 80386 24027 80402 24044
rect 79814 24011 80402 24027
rect 80832 24027 80848 24044
rect 81404 24044 81606 24061
rect 81664 24061 82624 24108
rect 81664 24044 81866 24061
rect 81404 24027 81420 24044
rect 80832 24011 81420 24027
rect 81850 24027 81866 24044
rect 82422 24044 82624 24061
rect 82682 24061 83642 24108
rect 82682 24044 82884 24061
rect 82422 24027 82438 24044
rect 81850 24011 82438 24027
rect 82868 24027 82884 24044
rect 83440 24044 83642 24061
rect 83700 24061 84660 24108
rect 83700 24044 83902 24061
rect 83440 24027 83456 24044
rect 82868 24011 83456 24027
rect 83886 24027 83902 24044
rect 84458 24044 84660 24061
rect 84718 24061 85678 24108
rect 84718 24044 84920 24061
rect 84458 24027 84474 24044
rect 83886 24011 84474 24027
rect 84904 24027 84920 24044
rect 85476 24044 85678 24061
rect 85736 24061 86696 24108
rect 85736 24044 85938 24061
rect 85476 24027 85492 24044
rect 84904 24011 85492 24027
rect 85922 24027 85938 24044
rect 86494 24044 86696 24061
rect 86754 24061 87714 24108
rect 86754 24044 86956 24061
rect 86494 24027 86510 24044
rect 85922 24011 86510 24027
rect 86940 24027 86956 24044
rect 87512 24044 87714 24061
rect 87512 24027 87528 24044
rect 86940 24011 87528 24027
rect 72656 23015 73244 23031
rect 72656 22998 72672 23015
rect 72470 22981 72672 22998
rect 73228 22998 73244 23015
rect 73674 23015 74262 23031
rect 73674 22998 73690 23015
rect 73228 22981 73430 22998
rect 72470 22934 73430 22981
rect 73488 22981 73690 22998
rect 74246 22998 74262 23015
rect 74692 23015 75280 23031
rect 74692 22998 74708 23015
rect 74246 22981 74448 22998
rect 73488 22934 74448 22981
rect 74506 22981 74708 22998
rect 75264 22998 75280 23015
rect 75710 23015 76298 23031
rect 75710 22998 75726 23015
rect 75264 22981 75466 22998
rect 74506 22934 75466 22981
rect 75524 22981 75726 22998
rect 76282 22998 76298 23015
rect 76728 23015 77316 23031
rect 76728 22998 76744 23015
rect 76282 22981 76484 22998
rect 75524 22934 76484 22981
rect 76542 22981 76744 22998
rect 77300 22998 77316 23015
rect 77746 23015 78334 23031
rect 77746 22998 77762 23015
rect 77300 22981 77502 22998
rect 76542 22934 77502 22981
rect 77560 22981 77762 22998
rect 78318 22998 78334 23015
rect 78764 23015 79352 23031
rect 78764 22998 78780 23015
rect 78318 22981 78520 22998
rect 77560 22934 78520 22981
rect 78578 22981 78780 22998
rect 79336 22998 79352 23015
rect 79782 23015 80370 23031
rect 79782 22998 79798 23015
rect 79336 22981 79538 22998
rect 78578 22934 79538 22981
rect 79596 22981 79798 22998
rect 80354 22998 80370 23015
rect 80800 23015 81388 23031
rect 80800 22998 80816 23015
rect 80354 22981 80556 22998
rect 79596 22934 80556 22981
rect 80614 22981 80816 22998
rect 81372 22998 81388 23015
rect 81818 23015 82406 23031
rect 81818 22998 81834 23015
rect 81372 22981 81574 22998
rect 80614 22934 81574 22981
rect 81632 22981 81834 22998
rect 82390 22998 82406 23015
rect 82836 23015 83424 23031
rect 82836 22998 82852 23015
rect 82390 22981 82592 22998
rect 81632 22934 82592 22981
rect 82650 22981 82852 22998
rect 83408 22998 83424 23015
rect 83854 23015 84442 23031
rect 83854 22998 83870 23015
rect 83408 22981 83610 22998
rect 82650 22934 83610 22981
rect 83668 22981 83870 22998
rect 84426 22998 84442 23015
rect 84872 23015 85460 23031
rect 84872 22998 84888 23015
rect 84426 22981 84628 22998
rect 83668 22934 84628 22981
rect 84686 22981 84888 22998
rect 85444 22998 85460 23015
rect 85890 23015 86478 23031
rect 85890 22998 85906 23015
rect 85444 22981 85646 22998
rect 84686 22934 85646 22981
rect 85704 22981 85906 22998
rect 86462 22998 86478 23015
rect 86908 23015 87496 23031
rect 86908 22998 86924 23015
rect 86462 22981 86664 22998
rect 85704 22934 86664 22981
rect 86722 22981 86924 22998
rect 87480 22998 87496 23015
rect 87480 22981 87682 22998
rect 86722 22934 87682 22981
rect 72470 22287 73430 22334
rect 72470 22270 72672 22287
rect 72656 22253 72672 22270
rect 73228 22270 73430 22287
rect 73488 22287 74448 22334
rect 73488 22270 73690 22287
rect 73228 22253 73244 22270
rect 72656 22237 73244 22253
rect 73674 22253 73690 22270
rect 74246 22270 74448 22287
rect 74506 22287 75466 22334
rect 74506 22270 74708 22287
rect 74246 22253 74262 22270
rect 73674 22237 74262 22253
rect 74692 22253 74708 22270
rect 75264 22270 75466 22287
rect 75524 22287 76484 22334
rect 75524 22270 75726 22287
rect 75264 22253 75280 22270
rect 74692 22237 75280 22253
rect 75710 22253 75726 22270
rect 76282 22270 76484 22287
rect 76542 22287 77502 22334
rect 76542 22270 76744 22287
rect 76282 22253 76298 22270
rect 75710 22237 76298 22253
rect 76728 22253 76744 22270
rect 77300 22270 77502 22287
rect 77560 22287 78520 22334
rect 77560 22270 77762 22287
rect 77300 22253 77316 22270
rect 76728 22237 77316 22253
rect 77746 22253 77762 22270
rect 78318 22270 78520 22287
rect 78578 22287 79538 22334
rect 78578 22270 78780 22287
rect 78318 22253 78334 22270
rect 77746 22237 78334 22253
rect 78764 22253 78780 22270
rect 79336 22270 79538 22287
rect 79596 22287 80556 22334
rect 79596 22270 79798 22287
rect 79336 22253 79352 22270
rect 78764 22237 79352 22253
rect 79782 22253 79798 22270
rect 80354 22270 80556 22287
rect 80614 22287 81574 22334
rect 80614 22270 80816 22287
rect 80354 22253 80370 22270
rect 79782 22237 80370 22253
rect 80800 22253 80816 22270
rect 81372 22270 81574 22287
rect 81632 22287 82592 22334
rect 81632 22270 81834 22287
rect 81372 22253 81388 22270
rect 80800 22237 81388 22253
rect 81818 22253 81834 22270
rect 82390 22270 82592 22287
rect 82650 22287 83610 22334
rect 82650 22270 82852 22287
rect 82390 22253 82406 22270
rect 81818 22237 82406 22253
rect 82836 22253 82852 22270
rect 83408 22270 83610 22287
rect 83668 22287 84628 22334
rect 83668 22270 83870 22287
rect 83408 22253 83424 22270
rect 82836 22237 83424 22253
rect 83854 22253 83870 22270
rect 84426 22270 84628 22287
rect 84686 22287 85646 22334
rect 84686 22270 84888 22287
rect 84426 22253 84442 22270
rect 83854 22237 84442 22253
rect 84872 22253 84888 22270
rect 85444 22270 85646 22287
rect 85704 22287 86664 22334
rect 85704 22270 85906 22287
rect 85444 22253 85460 22270
rect 84872 22237 85460 22253
rect 85890 22253 85906 22270
rect 86462 22270 86664 22287
rect 86722 22287 87682 22334
rect 86722 22270 86924 22287
rect 86462 22253 86478 22270
rect 85890 22237 86478 22253
rect 86908 22253 86924 22270
rect 87480 22270 87682 22287
rect 87480 22253 87496 22270
rect 86908 22237 87496 22253
rect 68648 21931 68756 21947
rect 68648 21914 68664 21931
rect 68622 21897 68664 21914
rect 68740 21914 68756 21931
rect 68866 21931 68974 21947
rect 68866 21914 68882 21931
rect 68740 21897 68782 21914
rect 68622 21850 68782 21897
rect 68840 21897 68882 21914
rect 68958 21914 68974 21931
rect 69084 21931 69192 21947
rect 69084 21914 69100 21931
rect 68958 21897 69000 21914
rect 68840 21850 69000 21897
rect 69058 21897 69100 21914
rect 69176 21914 69192 21931
rect 69302 21931 69410 21947
rect 69302 21914 69318 21931
rect 69176 21897 69218 21914
rect 69058 21850 69218 21897
rect 69276 21897 69318 21914
rect 69394 21914 69410 21931
rect 69520 21931 69628 21947
rect 69520 21914 69536 21931
rect 69394 21897 69436 21914
rect 69276 21850 69436 21897
rect 69494 21897 69536 21914
rect 69612 21914 69628 21931
rect 69738 21931 69846 21947
rect 69738 21914 69754 21931
rect 69612 21897 69654 21914
rect 69494 21850 69654 21897
rect 69712 21897 69754 21914
rect 69830 21914 69846 21931
rect 69956 21931 70064 21947
rect 69956 21914 69972 21931
rect 69830 21897 69872 21914
rect 69712 21850 69872 21897
rect 69930 21897 69972 21914
rect 70048 21914 70064 21931
rect 70174 21931 70282 21947
rect 70174 21914 70190 21931
rect 70048 21897 70090 21914
rect 69930 21850 70090 21897
rect 70148 21897 70190 21914
rect 70266 21914 70282 21931
rect 70392 21931 70500 21947
rect 70392 21914 70408 21931
rect 70266 21897 70308 21914
rect 70148 21850 70308 21897
rect 70366 21897 70408 21914
rect 70484 21914 70500 21931
rect 70610 21931 70718 21947
rect 70610 21914 70626 21931
rect 70484 21897 70526 21914
rect 70366 21850 70526 21897
rect 70584 21897 70626 21914
rect 70702 21914 70718 21931
rect 70702 21897 70744 21914
rect 70584 21850 70744 21897
rect 72656 21759 73244 21775
rect 72656 21742 72672 21759
rect 72470 21725 72672 21742
rect 73228 21742 73244 21759
rect 73674 21759 74262 21775
rect 73674 21742 73690 21759
rect 73228 21725 73430 21742
rect 72470 21678 73430 21725
rect 73488 21725 73690 21742
rect 74246 21742 74262 21759
rect 74692 21759 75280 21775
rect 74692 21742 74708 21759
rect 74246 21725 74448 21742
rect 73488 21678 74448 21725
rect 74506 21725 74708 21742
rect 75264 21742 75280 21759
rect 75710 21759 76298 21775
rect 75710 21742 75726 21759
rect 75264 21725 75466 21742
rect 74506 21678 75466 21725
rect 75524 21725 75726 21742
rect 76282 21742 76298 21759
rect 76728 21759 77316 21775
rect 76728 21742 76744 21759
rect 76282 21725 76484 21742
rect 75524 21678 76484 21725
rect 76542 21725 76744 21742
rect 77300 21742 77316 21759
rect 77746 21759 78334 21775
rect 77746 21742 77762 21759
rect 77300 21725 77502 21742
rect 76542 21678 77502 21725
rect 77560 21725 77762 21742
rect 78318 21742 78334 21759
rect 78764 21759 79352 21775
rect 78764 21742 78780 21759
rect 78318 21725 78520 21742
rect 77560 21678 78520 21725
rect 78578 21725 78780 21742
rect 79336 21742 79352 21759
rect 79782 21759 80370 21775
rect 79782 21742 79798 21759
rect 79336 21725 79538 21742
rect 78578 21678 79538 21725
rect 79596 21725 79798 21742
rect 80354 21742 80370 21759
rect 80800 21759 81388 21775
rect 80800 21742 80816 21759
rect 80354 21725 80556 21742
rect 79596 21678 80556 21725
rect 80614 21725 80816 21742
rect 81372 21742 81388 21759
rect 81818 21759 82406 21775
rect 81818 21742 81834 21759
rect 81372 21725 81574 21742
rect 80614 21678 81574 21725
rect 81632 21725 81834 21742
rect 82390 21742 82406 21759
rect 82836 21759 83424 21775
rect 82836 21742 82852 21759
rect 82390 21725 82592 21742
rect 81632 21678 82592 21725
rect 82650 21725 82852 21742
rect 83408 21742 83424 21759
rect 83854 21759 84442 21775
rect 83854 21742 83870 21759
rect 83408 21725 83610 21742
rect 82650 21678 83610 21725
rect 83668 21725 83870 21742
rect 84426 21742 84442 21759
rect 84872 21759 85460 21775
rect 84872 21742 84888 21759
rect 84426 21725 84628 21742
rect 83668 21678 84628 21725
rect 84686 21725 84888 21742
rect 85444 21742 85460 21759
rect 85890 21759 86478 21775
rect 85890 21742 85906 21759
rect 85444 21725 85646 21742
rect 84686 21678 85646 21725
rect 85704 21725 85906 21742
rect 86462 21742 86478 21759
rect 86908 21759 87496 21775
rect 86908 21742 86924 21759
rect 86462 21725 86664 21742
rect 85704 21678 86664 21725
rect 86722 21725 86924 21742
rect 87480 21742 87496 21759
rect 87480 21725 87682 21742
rect 86722 21678 87682 21725
rect 68622 21403 68782 21450
rect 68622 21386 68664 21403
rect 68648 21369 68664 21386
rect 68740 21386 68782 21403
rect 68840 21403 69000 21450
rect 68840 21386 68882 21403
rect 68740 21369 68756 21386
rect 68648 21353 68756 21369
rect 68866 21369 68882 21386
rect 68958 21386 69000 21403
rect 69058 21403 69218 21450
rect 69058 21386 69100 21403
rect 68958 21369 68974 21386
rect 68866 21353 68974 21369
rect 69084 21369 69100 21386
rect 69176 21386 69218 21403
rect 69276 21403 69436 21450
rect 69276 21386 69318 21403
rect 69176 21369 69192 21386
rect 69084 21353 69192 21369
rect 69302 21369 69318 21386
rect 69394 21386 69436 21403
rect 69494 21403 69654 21450
rect 69494 21386 69536 21403
rect 69394 21369 69410 21386
rect 69302 21353 69410 21369
rect 69520 21369 69536 21386
rect 69612 21386 69654 21403
rect 69712 21403 69872 21450
rect 69712 21386 69754 21403
rect 69612 21369 69628 21386
rect 69520 21353 69628 21369
rect 69738 21369 69754 21386
rect 69830 21386 69872 21403
rect 69930 21403 70090 21450
rect 69930 21386 69972 21403
rect 69830 21369 69846 21386
rect 69738 21353 69846 21369
rect 69956 21369 69972 21386
rect 70048 21386 70090 21403
rect 70148 21403 70308 21450
rect 70148 21386 70190 21403
rect 70048 21369 70064 21386
rect 69956 21353 70064 21369
rect 70174 21369 70190 21386
rect 70266 21386 70308 21403
rect 70366 21403 70526 21450
rect 70366 21386 70408 21403
rect 70266 21369 70282 21386
rect 70174 21353 70282 21369
rect 70392 21369 70408 21386
rect 70484 21386 70526 21403
rect 70584 21403 70744 21450
rect 70584 21386 70626 21403
rect 70484 21369 70500 21386
rect 70392 21353 70500 21369
rect 70610 21369 70626 21386
rect 70702 21386 70744 21403
rect 70702 21369 70718 21386
rect 70610 21353 70718 21369
rect 72470 21031 73430 21078
rect 72470 21014 72672 21031
rect 68648 20993 68756 21009
rect 68648 20976 68664 20993
rect 68622 20959 68664 20976
rect 68740 20976 68756 20993
rect 68866 20993 68974 21009
rect 68866 20976 68882 20993
rect 68740 20959 68782 20976
rect 68622 20912 68782 20959
rect 68840 20959 68882 20976
rect 68958 20976 68974 20993
rect 69084 20993 69192 21009
rect 69084 20976 69100 20993
rect 68958 20959 69000 20976
rect 68840 20912 69000 20959
rect 69058 20959 69100 20976
rect 69176 20976 69192 20993
rect 69302 20993 69410 21009
rect 69302 20976 69318 20993
rect 69176 20959 69218 20976
rect 69058 20912 69218 20959
rect 69276 20959 69318 20976
rect 69394 20976 69410 20993
rect 69520 20993 69628 21009
rect 69520 20976 69536 20993
rect 69394 20959 69436 20976
rect 69276 20912 69436 20959
rect 69494 20959 69536 20976
rect 69612 20976 69628 20993
rect 69738 20993 69846 21009
rect 69738 20976 69754 20993
rect 69612 20959 69654 20976
rect 69494 20912 69654 20959
rect 69712 20959 69754 20976
rect 69830 20976 69846 20993
rect 69956 20993 70064 21009
rect 69956 20976 69972 20993
rect 69830 20959 69872 20976
rect 69712 20912 69872 20959
rect 69930 20959 69972 20976
rect 70048 20976 70064 20993
rect 70174 20993 70282 21009
rect 70174 20976 70190 20993
rect 70048 20959 70090 20976
rect 69930 20912 70090 20959
rect 70148 20959 70190 20976
rect 70266 20976 70282 20993
rect 70392 20993 70500 21009
rect 70392 20976 70408 20993
rect 70266 20959 70308 20976
rect 70148 20912 70308 20959
rect 70366 20959 70408 20976
rect 70484 20976 70500 20993
rect 70610 20993 70718 21009
rect 70610 20976 70626 20993
rect 70484 20959 70526 20976
rect 70366 20912 70526 20959
rect 70584 20959 70626 20976
rect 70702 20976 70718 20993
rect 72656 20997 72672 21014
rect 73228 21014 73430 21031
rect 73488 21031 74448 21078
rect 73488 21014 73690 21031
rect 73228 20997 73244 21014
rect 72656 20981 73244 20997
rect 73674 20997 73690 21014
rect 74246 21014 74448 21031
rect 74506 21031 75466 21078
rect 74506 21014 74708 21031
rect 74246 20997 74262 21014
rect 73674 20981 74262 20997
rect 74692 20997 74708 21014
rect 75264 21014 75466 21031
rect 75524 21031 76484 21078
rect 75524 21014 75726 21031
rect 75264 20997 75280 21014
rect 74692 20981 75280 20997
rect 75710 20997 75726 21014
rect 76282 21014 76484 21031
rect 76542 21031 77502 21078
rect 76542 21014 76744 21031
rect 76282 20997 76298 21014
rect 75710 20981 76298 20997
rect 76728 20997 76744 21014
rect 77300 21014 77502 21031
rect 77560 21031 78520 21078
rect 77560 21014 77762 21031
rect 77300 20997 77316 21014
rect 76728 20981 77316 20997
rect 77746 20997 77762 21014
rect 78318 21014 78520 21031
rect 78578 21031 79538 21078
rect 78578 21014 78780 21031
rect 78318 20997 78334 21014
rect 77746 20981 78334 20997
rect 78764 20997 78780 21014
rect 79336 21014 79538 21031
rect 79596 21031 80556 21078
rect 79596 21014 79798 21031
rect 79336 20997 79352 21014
rect 78764 20981 79352 20997
rect 79782 20997 79798 21014
rect 80354 21014 80556 21031
rect 80614 21031 81574 21078
rect 80614 21014 80816 21031
rect 80354 20997 80370 21014
rect 79782 20981 80370 20997
rect 80800 20997 80816 21014
rect 81372 21014 81574 21031
rect 81632 21031 82592 21078
rect 81632 21014 81834 21031
rect 81372 20997 81388 21014
rect 80800 20981 81388 20997
rect 81818 20997 81834 21014
rect 82390 21014 82592 21031
rect 82650 21031 83610 21078
rect 82650 21014 82852 21031
rect 82390 20997 82406 21014
rect 81818 20981 82406 20997
rect 82836 20997 82852 21014
rect 83408 21014 83610 21031
rect 83668 21031 84628 21078
rect 83668 21014 83870 21031
rect 83408 20997 83424 21014
rect 82836 20981 83424 20997
rect 83854 20997 83870 21014
rect 84426 21014 84628 21031
rect 84686 21031 85646 21078
rect 84686 21014 84888 21031
rect 84426 20997 84442 21014
rect 83854 20981 84442 20997
rect 84872 20997 84888 21014
rect 85444 21014 85646 21031
rect 85704 21031 86664 21078
rect 85704 21014 85906 21031
rect 85444 20997 85460 21014
rect 84872 20981 85460 20997
rect 85890 20997 85906 21014
rect 86462 21014 86664 21031
rect 86722 21031 87682 21078
rect 86722 21014 86924 21031
rect 86462 20997 86478 21014
rect 85890 20981 86478 20997
rect 86908 20997 86924 21014
rect 87480 21014 87682 21031
rect 87480 20997 87496 21014
rect 86908 20981 87496 20997
rect 70702 20959 70744 20976
rect 70584 20912 70744 20959
rect 68622 20465 68782 20512
rect 68622 20448 68664 20465
rect 68648 20431 68664 20448
rect 68740 20448 68782 20465
rect 68840 20465 69000 20512
rect 68840 20448 68882 20465
rect 68740 20431 68756 20448
rect 68648 20415 68756 20431
rect 68866 20431 68882 20448
rect 68958 20448 69000 20465
rect 69058 20465 69218 20512
rect 69058 20448 69100 20465
rect 68958 20431 68974 20448
rect 68866 20415 68974 20431
rect 69084 20431 69100 20448
rect 69176 20448 69218 20465
rect 69276 20465 69436 20512
rect 69276 20448 69318 20465
rect 69176 20431 69192 20448
rect 69084 20415 69192 20431
rect 69302 20431 69318 20448
rect 69394 20448 69436 20465
rect 69494 20465 69654 20512
rect 69494 20448 69536 20465
rect 69394 20431 69410 20448
rect 69302 20415 69410 20431
rect 69520 20431 69536 20448
rect 69612 20448 69654 20465
rect 69712 20465 69872 20512
rect 69712 20448 69754 20465
rect 69612 20431 69628 20448
rect 69520 20415 69628 20431
rect 69738 20431 69754 20448
rect 69830 20448 69872 20465
rect 69930 20465 70090 20512
rect 69930 20448 69972 20465
rect 69830 20431 69846 20448
rect 69738 20415 69846 20431
rect 69956 20431 69972 20448
rect 70048 20448 70090 20465
rect 70148 20465 70308 20512
rect 70148 20448 70190 20465
rect 70048 20431 70064 20448
rect 69956 20415 70064 20431
rect 70174 20431 70190 20448
rect 70266 20448 70308 20465
rect 70366 20465 70526 20512
rect 70366 20448 70408 20465
rect 70266 20431 70282 20448
rect 70174 20415 70282 20431
rect 70392 20431 70408 20448
rect 70484 20448 70526 20465
rect 70584 20465 70744 20512
rect 72656 20503 73244 20519
rect 72656 20486 72672 20503
rect 70584 20448 70626 20465
rect 70484 20431 70500 20448
rect 70392 20415 70500 20431
rect 70610 20431 70626 20448
rect 70702 20448 70744 20465
rect 72470 20469 72672 20486
rect 73228 20486 73244 20503
rect 73674 20503 74262 20519
rect 73674 20486 73690 20503
rect 73228 20469 73430 20486
rect 70702 20431 70718 20448
rect 70610 20415 70718 20431
rect 72470 20422 73430 20469
rect 73488 20469 73690 20486
rect 74246 20486 74262 20503
rect 74692 20503 75280 20519
rect 74692 20486 74708 20503
rect 74246 20469 74448 20486
rect 73488 20422 74448 20469
rect 74506 20469 74708 20486
rect 75264 20486 75280 20503
rect 75710 20503 76298 20519
rect 75710 20486 75726 20503
rect 75264 20469 75466 20486
rect 74506 20422 75466 20469
rect 75524 20469 75726 20486
rect 76282 20486 76298 20503
rect 76728 20503 77316 20519
rect 76728 20486 76744 20503
rect 76282 20469 76484 20486
rect 75524 20422 76484 20469
rect 76542 20469 76744 20486
rect 77300 20486 77316 20503
rect 77746 20503 78334 20519
rect 77746 20486 77762 20503
rect 77300 20469 77502 20486
rect 76542 20422 77502 20469
rect 77560 20469 77762 20486
rect 78318 20486 78334 20503
rect 78764 20503 79352 20519
rect 78764 20486 78780 20503
rect 78318 20469 78520 20486
rect 77560 20422 78520 20469
rect 78578 20469 78780 20486
rect 79336 20486 79352 20503
rect 79782 20503 80370 20519
rect 79782 20486 79798 20503
rect 79336 20469 79538 20486
rect 78578 20422 79538 20469
rect 79596 20469 79798 20486
rect 80354 20486 80370 20503
rect 80800 20503 81388 20519
rect 80800 20486 80816 20503
rect 80354 20469 80556 20486
rect 79596 20422 80556 20469
rect 80614 20469 80816 20486
rect 81372 20486 81388 20503
rect 81818 20503 82406 20519
rect 81818 20486 81834 20503
rect 81372 20469 81574 20486
rect 80614 20422 81574 20469
rect 81632 20469 81834 20486
rect 82390 20486 82406 20503
rect 82836 20503 83424 20519
rect 82836 20486 82852 20503
rect 82390 20469 82592 20486
rect 81632 20422 82592 20469
rect 82650 20469 82852 20486
rect 83408 20486 83424 20503
rect 83854 20503 84442 20519
rect 83854 20486 83870 20503
rect 83408 20469 83610 20486
rect 82650 20422 83610 20469
rect 83668 20469 83870 20486
rect 84426 20486 84442 20503
rect 84872 20503 85460 20519
rect 84872 20486 84888 20503
rect 84426 20469 84628 20486
rect 83668 20422 84628 20469
rect 84686 20469 84888 20486
rect 85444 20486 85460 20503
rect 85890 20503 86478 20519
rect 85890 20486 85906 20503
rect 85444 20469 85646 20486
rect 84686 20422 85646 20469
rect 85704 20469 85906 20486
rect 86462 20486 86478 20503
rect 86908 20503 87496 20519
rect 86908 20486 86924 20503
rect 86462 20469 86664 20486
rect 85704 20422 86664 20469
rect 86722 20469 86924 20486
rect 87480 20486 87496 20503
rect 87480 20469 87682 20486
rect 86722 20422 87682 20469
rect 68648 20055 68756 20071
rect 68648 20038 68664 20055
rect 68622 20021 68664 20038
rect 68740 20038 68756 20055
rect 68866 20055 68974 20071
rect 68866 20038 68882 20055
rect 68740 20021 68782 20038
rect 68622 19974 68782 20021
rect 68840 20021 68882 20038
rect 68958 20038 68974 20055
rect 69084 20055 69192 20071
rect 69084 20038 69100 20055
rect 68958 20021 69000 20038
rect 68840 19974 69000 20021
rect 69058 20021 69100 20038
rect 69176 20038 69192 20055
rect 69302 20055 69410 20071
rect 69302 20038 69318 20055
rect 69176 20021 69218 20038
rect 69058 19974 69218 20021
rect 69276 20021 69318 20038
rect 69394 20038 69410 20055
rect 69520 20055 69628 20071
rect 69520 20038 69536 20055
rect 69394 20021 69436 20038
rect 69276 19974 69436 20021
rect 69494 20021 69536 20038
rect 69612 20038 69628 20055
rect 69738 20055 69846 20071
rect 69738 20038 69754 20055
rect 69612 20021 69654 20038
rect 69494 19974 69654 20021
rect 69712 20021 69754 20038
rect 69830 20038 69846 20055
rect 69956 20055 70064 20071
rect 69956 20038 69972 20055
rect 69830 20021 69872 20038
rect 69712 19974 69872 20021
rect 69930 20021 69972 20038
rect 70048 20038 70064 20055
rect 70174 20055 70282 20071
rect 70174 20038 70190 20055
rect 70048 20021 70090 20038
rect 69930 19974 70090 20021
rect 70148 20021 70190 20038
rect 70266 20038 70282 20055
rect 70392 20055 70500 20071
rect 70392 20038 70408 20055
rect 70266 20021 70308 20038
rect 70148 19974 70308 20021
rect 70366 20021 70408 20038
rect 70484 20038 70500 20055
rect 70610 20055 70718 20071
rect 70610 20038 70626 20055
rect 70484 20021 70526 20038
rect 70366 19974 70526 20021
rect 70584 20021 70626 20038
rect 70702 20038 70718 20055
rect 70702 20021 70744 20038
rect 70584 19974 70744 20021
rect 72470 19775 73430 19822
rect 72470 19758 72672 19775
rect 72656 19741 72672 19758
rect 73228 19758 73430 19775
rect 73488 19775 74448 19822
rect 73488 19758 73690 19775
rect 73228 19741 73244 19758
rect 72656 19725 73244 19741
rect 73674 19741 73690 19758
rect 74246 19758 74448 19775
rect 74506 19775 75466 19822
rect 74506 19758 74708 19775
rect 74246 19741 74262 19758
rect 73674 19725 74262 19741
rect 74692 19741 74708 19758
rect 75264 19758 75466 19775
rect 75524 19775 76484 19822
rect 75524 19758 75726 19775
rect 75264 19741 75280 19758
rect 74692 19725 75280 19741
rect 75710 19741 75726 19758
rect 76282 19758 76484 19775
rect 76542 19775 77502 19822
rect 76542 19758 76744 19775
rect 76282 19741 76298 19758
rect 75710 19725 76298 19741
rect 76728 19741 76744 19758
rect 77300 19758 77502 19775
rect 77560 19775 78520 19822
rect 77560 19758 77762 19775
rect 77300 19741 77316 19758
rect 76728 19725 77316 19741
rect 77746 19741 77762 19758
rect 78318 19758 78520 19775
rect 78578 19775 79538 19822
rect 78578 19758 78780 19775
rect 78318 19741 78334 19758
rect 77746 19725 78334 19741
rect 78764 19741 78780 19758
rect 79336 19758 79538 19775
rect 79596 19775 80556 19822
rect 79596 19758 79798 19775
rect 79336 19741 79352 19758
rect 78764 19725 79352 19741
rect 79782 19741 79798 19758
rect 80354 19758 80556 19775
rect 80614 19775 81574 19822
rect 80614 19758 80816 19775
rect 80354 19741 80370 19758
rect 79782 19725 80370 19741
rect 80800 19741 80816 19758
rect 81372 19758 81574 19775
rect 81632 19775 82592 19822
rect 81632 19758 81834 19775
rect 81372 19741 81388 19758
rect 80800 19725 81388 19741
rect 81818 19741 81834 19758
rect 82390 19758 82592 19775
rect 82650 19775 83610 19822
rect 82650 19758 82852 19775
rect 82390 19741 82406 19758
rect 81818 19725 82406 19741
rect 82836 19741 82852 19758
rect 83408 19758 83610 19775
rect 83668 19775 84628 19822
rect 83668 19758 83870 19775
rect 83408 19741 83424 19758
rect 82836 19725 83424 19741
rect 83854 19741 83870 19758
rect 84426 19758 84628 19775
rect 84686 19775 85646 19822
rect 84686 19758 84888 19775
rect 84426 19741 84442 19758
rect 83854 19725 84442 19741
rect 84872 19741 84888 19758
rect 85444 19758 85646 19775
rect 85704 19775 86664 19822
rect 85704 19758 85906 19775
rect 85444 19741 85460 19758
rect 84872 19725 85460 19741
rect 85890 19741 85906 19758
rect 86462 19758 86664 19775
rect 86722 19775 87682 19822
rect 86722 19758 86924 19775
rect 86462 19741 86478 19758
rect 85890 19725 86478 19741
rect 86908 19741 86924 19758
rect 87480 19758 87682 19775
rect 87480 19741 87496 19758
rect 86908 19725 87496 19741
rect 68622 19527 68782 19574
rect 68622 19510 68664 19527
rect 68648 19493 68664 19510
rect 68740 19510 68782 19527
rect 68840 19527 69000 19574
rect 68840 19510 68882 19527
rect 68740 19493 68756 19510
rect 68648 19477 68756 19493
rect 68866 19493 68882 19510
rect 68958 19510 69000 19527
rect 69058 19527 69218 19574
rect 69058 19510 69100 19527
rect 68958 19493 68974 19510
rect 68866 19477 68974 19493
rect 69084 19493 69100 19510
rect 69176 19510 69218 19527
rect 69276 19527 69436 19574
rect 69276 19510 69318 19527
rect 69176 19493 69192 19510
rect 69084 19477 69192 19493
rect 69302 19493 69318 19510
rect 69394 19510 69436 19527
rect 69494 19527 69654 19574
rect 69494 19510 69536 19527
rect 69394 19493 69410 19510
rect 69302 19477 69410 19493
rect 69520 19493 69536 19510
rect 69612 19510 69654 19527
rect 69712 19527 69872 19574
rect 69712 19510 69754 19527
rect 69612 19493 69628 19510
rect 69520 19477 69628 19493
rect 69738 19493 69754 19510
rect 69830 19510 69872 19527
rect 69930 19527 70090 19574
rect 69930 19510 69972 19527
rect 69830 19493 69846 19510
rect 69738 19477 69846 19493
rect 69956 19493 69972 19510
rect 70048 19510 70090 19527
rect 70148 19527 70308 19574
rect 70148 19510 70190 19527
rect 70048 19493 70064 19510
rect 69956 19477 70064 19493
rect 70174 19493 70190 19510
rect 70266 19510 70308 19527
rect 70366 19527 70526 19574
rect 70366 19510 70408 19527
rect 70266 19493 70282 19510
rect 70174 19477 70282 19493
rect 70392 19493 70408 19510
rect 70484 19510 70526 19527
rect 70584 19527 70744 19574
rect 70584 19510 70626 19527
rect 70484 19493 70500 19510
rect 70392 19477 70500 19493
rect 70610 19493 70626 19510
rect 70702 19510 70744 19527
rect 70702 19493 70718 19510
rect 70610 19477 70718 19493
rect 72656 19247 73244 19263
rect 72656 19230 72672 19247
rect 72470 19213 72672 19230
rect 73228 19230 73244 19247
rect 73674 19247 74262 19263
rect 73674 19230 73690 19247
rect 73228 19213 73430 19230
rect 72470 19166 73430 19213
rect 73488 19213 73690 19230
rect 74246 19230 74262 19247
rect 74692 19247 75280 19263
rect 74692 19230 74708 19247
rect 74246 19213 74448 19230
rect 73488 19166 74448 19213
rect 74506 19213 74708 19230
rect 75264 19230 75280 19247
rect 75710 19247 76298 19263
rect 75710 19230 75726 19247
rect 75264 19213 75466 19230
rect 74506 19166 75466 19213
rect 75524 19213 75726 19230
rect 76282 19230 76298 19247
rect 76728 19247 77316 19263
rect 76728 19230 76744 19247
rect 76282 19213 76484 19230
rect 75524 19166 76484 19213
rect 76542 19213 76744 19230
rect 77300 19230 77316 19247
rect 77746 19247 78334 19263
rect 77746 19230 77762 19247
rect 77300 19213 77502 19230
rect 76542 19166 77502 19213
rect 77560 19213 77762 19230
rect 78318 19230 78334 19247
rect 78764 19247 79352 19263
rect 78764 19230 78780 19247
rect 78318 19213 78520 19230
rect 77560 19166 78520 19213
rect 78578 19213 78780 19230
rect 79336 19230 79352 19247
rect 79782 19247 80370 19263
rect 79782 19230 79798 19247
rect 79336 19213 79538 19230
rect 78578 19166 79538 19213
rect 79596 19213 79798 19230
rect 80354 19230 80370 19247
rect 80800 19247 81388 19263
rect 80800 19230 80816 19247
rect 80354 19213 80556 19230
rect 79596 19166 80556 19213
rect 80614 19213 80816 19230
rect 81372 19230 81388 19247
rect 81818 19247 82406 19263
rect 81818 19230 81834 19247
rect 81372 19213 81574 19230
rect 80614 19166 81574 19213
rect 81632 19213 81834 19230
rect 82390 19230 82406 19247
rect 82836 19247 83424 19263
rect 82836 19230 82852 19247
rect 82390 19213 82592 19230
rect 81632 19166 82592 19213
rect 82650 19213 82852 19230
rect 83408 19230 83424 19247
rect 83854 19247 84442 19263
rect 83854 19230 83870 19247
rect 83408 19213 83610 19230
rect 82650 19166 83610 19213
rect 83668 19213 83870 19230
rect 84426 19230 84442 19247
rect 84872 19247 85460 19263
rect 84872 19230 84888 19247
rect 84426 19213 84628 19230
rect 83668 19166 84628 19213
rect 84686 19213 84888 19230
rect 85444 19230 85460 19247
rect 85890 19247 86478 19263
rect 85890 19230 85906 19247
rect 85444 19213 85646 19230
rect 84686 19166 85646 19213
rect 85704 19213 85906 19230
rect 86462 19230 86478 19247
rect 86908 19247 87496 19263
rect 86908 19230 86924 19247
rect 86462 19213 86664 19230
rect 85704 19166 86664 19213
rect 86722 19213 86924 19230
rect 87480 19230 87496 19247
rect 87480 19213 87682 19230
rect 86722 19166 87682 19213
rect 68648 19117 68756 19133
rect 68648 19100 68664 19117
rect 68622 19083 68664 19100
rect 68740 19100 68756 19117
rect 68866 19117 68974 19133
rect 68866 19100 68882 19117
rect 68740 19083 68782 19100
rect 68622 19036 68782 19083
rect 68840 19083 68882 19100
rect 68958 19100 68974 19117
rect 69084 19117 69192 19133
rect 69084 19100 69100 19117
rect 68958 19083 69000 19100
rect 68840 19036 69000 19083
rect 69058 19083 69100 19100
rect 69176 19100 69192 19117
rect 69302 19117 69410 19133
rect 69302 19100 69318 19117
rect 69176 19083 69218 19100
rect 69058 19036 69218 19083
rect 69276 19083 69318 19100
rect 69394 19100 69410 19117
rect 69520 19117 69628 19133
rect 69520 19100 69536 19117
rect 69394 19083 69436 19100
rect 69276 19036 69436 19083
rect 69494 19083 69536 19100
rect 69612 19100 69628 19117
rect 69738 19117 69846 19133
rect 69738 19100 69754 19117
rect 69612 19083 69654 19100
rect 69494 19036 69654 19083
rect 69712 19083 69754 19100
rect 69830 19100 69846 19117
rect 69956 19117 70064 19133
rect 69956 19100 69972 19117
rect 69830 19083 69872 19100
rect 69712 19036 69872 19083
rect 69930 19083 69972 19100
rect 70048 19100 70064 19117
rect 70174 19117 70282 19133
rect 70174 19100 70190 19117
rect 70048 19083 70090 19100
rect 69930 19036 70090 19083
rect 70148 19083 70190 19100
rect 70266 19100 70282 19117
rect 70392 19117 70500 19133
rect 70392 19100 70408 19117
rect 70266 19083 70308 19100
rect 70148 19036 70308 19083
rect 70366 19083 70408 19100
rect 70484 19100 70500 19117
rect 70610 19117 70718 19133
rect 70610 19100 70626 19117
rect 70484 19083 70526 19100
rect 70366 19036 70526 19083
rect 70584 19083 70626 19100
rect 70702 19100 70718 19117
rect 70702 19083 70744 19100
rect 70584 19036 70744 19083
rect 68622 18589 68782 18636
rect 68622 18572 68664 18589
rect 68648 18555 68664 18572
rect 68740 18572 68782 18589
rect 68840 18589 69000 18636
rect 68840 18572 68882 18589
rect 68740 18555 68756 18572
rect 68648 18539 68756 18555
rect 68866 18555 68882 18572
rect 68958 18572 69000 18589
rect 69058 18589 69218 18636
rect 69058 18572 69100 18589
rect 68958 18555 68974 18572
rect 68866 18539 68974 18555
rect 69084 18555 69100 18572
rect 69176 18572 69218 18589
rect 69276 18589 69436 18636
rect 69276 18572 69318 18589
rect 69176 18555 69192 18572
rect 69084 18539 69192 18555
rect 69302 18555 69318 18572
rect 69394 18572 69436 18589
rect 69494 18589 69654 18636
rect 69494 18572 69536 18589
rect 69394 18555 69410 18572
rect 69302 18539 69410 18555
rect 69520 18555 69536 18572
rect 69612 18572 69654 18589
rect 69712 18589 69872 18636
rect 69712 18572 69754 18589
rect 69612 18555 69628 18572
rect 69520 18539 69628 18555
rect 69738 18555 69754 18572
rect 69830 18572 69872 18589
rect 69930 18589 70090 18636
rect 69930 18572 69972 18589
rect 69830 18555 69846 18572
rect 69738 18539 69846 18555
rect 69956 18555 69972 18572
rect 70048 18572 70090 18589
rect 70148 18589 70308 18636
rect 70148 18572 70190 18589
rect 70048 18555 70064 18572
rect 69956 18539 70064 18555
rect 70174 18555 70190 18572
rect 70266 18572 70308 18589
rect 70366 18589 70526 18636
rect 70366 18572 70408 18589
rect 70266 18555 70282 18572
rect 70174 18539 70282 18555
rect 70392 18555 70408 18572
rect 70484 18572 70526 18589
rect 70584 18589 70744 18636
rect 70584 18572 70626 18589
rect 70484 18555 70500 18572
rect 70392 18539 70500 18555
rect 70610 18555 70626 18572
rect 70702 18572 70744 18589
rect 70702 18555 70718 18572
rect 70610 18539 70718 18555
rect 72470 18519 73430 18566
rect 72470 18502 72672 18519
rect 72656 18485 72672 18502
rect 73228 18502 73430 18519
rect 73488 18519 74448 18566
rect 73488 18502 73690 18519
rect 73228 18485 73244 18502
rect 72656 18469 73244 18485
rect 73674 18485 73690 18502
rect 74246 18502 74448 18519
rect 74506 18519 75466 18566
rect 74506 18502 74708 18519
rect 74246 18485 74262 18502
rect 73674 18469 74262 18485
rect 74692 18485 74708 18502
rect 75264 18502 75466 18519
rect 75524 18519 76484 18566
rect 75524 18502 75726 18519
rect 75264 18485 75280 18502
rect 74692 18469 75280 18485
rect 75710 18485 75726 18502
rect 76282 18502 76484 18519
rect 76542 18519 77502 18566
rect 76542 18502 76744 18519
rect 76282 18485 76298 18502
rect 75710 18469 76298 18485
rect 76728 18485 76744 18502
rect 77300 18502 77502 18519
rect 77560 18519 78520 18566
rect 77560 18502 77762 18519
rect 77300 18485 77316 18502
rect 76728 18469 77316 18485
rect 77746 18485 77762 18502
rect 78318 18502 78520 18519
rect 78578 18519 79538 18566
rect 78578 18502 78780 18519
rect 78318 18485 78334 18502
rect 77746 18469 78334 18485
rect 78764 18485 78780 18502
rect 79336 18502 79538 18519
rect 79596 18519 80556 18566
rect 79596 18502 79798 18519
rect 79336 18485 79352 18502
rect 78764 18469 79352 18485
rect 79782 18485 79798 18502
rect 80354 18502 80556 18519
rect 80614 18519 81574 18566
rect 80614 18502 80816 18519
rect 80354 18485 80370 18502
rect 79782 18469 80370 18485
rect 80800 18485 80816 18502
rect 81372 18502 81574 18519
rect 81632 18519 82592 18566
rect 81632 18502 81834 18519
rect 81372 18485 81388 18502
rect 80800 18469 81388 18485
rect 81818 18485 81834 18502
rect 82390 18502 82592 18519
rect 82650 18519 83610 18566
rect 82650 18502 82852 18519
rect 82390 18485 82406 18502
rect 81818 18469 82406 18485
rect 82836 18485 82852 18502
rect 83408 18502 83610 18519
rect 83668 18519 84628 18566
rect 83668 18502 83870 18519
rect 83408 18485 83424 18502
rect 82836 18469 83424 18485
rect 83854 18485 83870 18502
rect 84426 18502 84628 18519
rect 84686 18519 85646 18566
rect 84686 18502 84888 18519
rect 84426 18485 84442 18502
rect 83854 18469 84442 18485
rect 84872 18485 84888 18502
rect 85444 18502 85646 18519
rect 85704 18519 86664 18566
rect 85704 18502 85906 18519
rect 85444 18485 85460 18502
rect 84872 18469 85460 18485
rect 85890 18485 85906 18502
rect 86462 18502 86664 18519
rect 86722 18519 87682 18566
rect 86722 18502 86924 18519
rect 86462 18485 86478 18502
rect 85890 18469 86478 18485
rect 86908 18485 86924 18502
rect 87480 18502 87682 18519
rect 87480 18485 87496 18502
rect 86908 18469 87496 18485
rect -12900 16179 -12768 16195
rect -12900 16162 -12884 16179
rect -12934 16145 -12884 16162
rect -12784 16162 -12768 16179
rect -12642 16179 -12510 16195
rect -12642 16162 -12626 16179
rect -12784 16145 -12734 16162
rect -12934 16098 -12734 16145
rect -12676 16145 -12626 16162
rect -12526 16162 -12510 16179
rect -12384 16179 -12252 16195
rect -12384 16162 -12368 16179
rect -12526 16145 -12476 16162
rect -12676 16098 -12476 16145
rect -12418 16145 -12368 16162
rect -12268 16162 -12252 16179
rect -12126 16179 -11994 16195
rect -12126 16162 -12110 16179
rect -12268 16145 -12218 16162
rect -12418 16098 -12218 16145
rect -12160 16145 -12110 16162
rect -12010 16162 -11994 16179
rect -11868 16179 -11736 16195
rect -11868 16162 -11852 16179
rect -12010 16145 -11960 16162
rect -12160 16098 -11960 16145
rect -11902 16145 -11852 16162
rect -11752 16162 -11736 16179
rect -11610 16179 -11478 16195
rect -11610 16162 -11594 16179
rect -11752 16145 -11702 16162
rect -11902 16098 -11702 16145
rect -11644 16145 -11594 16162
rect -11494 16162 -11478 16179
rect -11494 16145 -11444 16162
rect -11644 16098 -11444 16145
rect -12934 15651 -12734 15698
rect -12934 15634 -12884 15651
rect -12900 15617 -12884 15634
rect -12784 15634 -12734 15651
rect -12676 15651 -12476 15698
rect -12676 15634 -12626 15651
rect -12784 15617 -12768 15634
rect -12900 15601 -12768 15617
rect -12642 15617 -12626 15634
rect -12526 15634 -12476 15651
rect -12418 15651 -12218 15698
rect -12418 15634 -12368 15651
rect -12526 15617 -12510 15634
rect -12642 15601 -12510 15617
rect -12384 15617 -12368 15634
rect -12268 15634 -12218 15651
rect -12160 15651 -11960 15698
rect -12160 15634 -12110 15651
rect -12268 15617 -12252 15634
rect -12384 15601 -12252 15617
rect -12126 15617 -12110 15634
rect -12010 15634 -11960 15651
rect -11902 15651 -11702 15698
rect -11902 15634 -11852 15651
rect -12010 15617 -11994 15634
rect -12126 15601 -11994 15617
rect -11868 15617 -11852 15634
rect -11752 15634 -11702 15651
rect -11644 15651 -11444 15698
rect -11644 15634 -11594 15651
rect -11752 15617 -11736 15634
rect -11868 15601 -11736 15617
rect -11610 15617 -11594 15634
rect -11494 15634 -11444 15651
rect -11494 15617 -11478 15634
rect -11610 15601 -11478 15617
rect -11084 15715 -11054 15741
rect -10300 16179 -10168 16195
rect -10300 16162 -10284 16179
rect -10334 16145 -10284 16162
rect -10184 16162 -10168 16179
rect -10042 16179 -9910 16195
rect -10042 16162 -10026 16179
rect -10184 16145 -10134 16162
rect -10334 16098 -10134 16145
rect -10076 16145 -10026 16162
rect -9926 16162 -9910 16179
rect -9784 16179 -9652 16195
rect -9784 16162 -9768 16179
rect -9926 16145 -9876 16162
rect -10076 16098 -9876 16145
rect -9818 16145 -9768 16162
rect -9668 16162 -9652 16179
rect -9526 16179 -9394 16195
rect -9526 16162 -9510 16179
rect -9668 16145 -9618 16162
rect -9818 16098 -9618 16145
rect -9560 16145 -9510 16162
rect -9410 16162 -9394 16179
rect -9268 16179 -9136 16195
rect -9268 16162 -9252 16179
rect -9410 16145 -9360 16162
rect -9560 16098 -9360 16145
rect -9302 16145 -9252 16162
rect -9152 16162 -9136 16179
rect -9010 16179 -8878 16195
rect -9010 16162 -8994 16179
rect -9152 16145 -9102 16162
rect -9302 16098 -9102 16145
rect -9044 16145 -8994 16162
rect -8894 16162 -8878 16179
rect -8894 16145 -8844 16162
rect -9044 16098 -8844 16145
rect -10334 15651 -10134 15698
rect -10334 15634 -10284 15651
rect -10300 15617 -10284 15634
rect -10184 15634 -10134 15651
rect -10076 15651 -9876 15698
rect -10076 15634 -10026 15651
rect -10184 15617 -10168 15634
rect -10300 15601 -10168 15617
rect -10042 15617 -10026 15634
rect -9926 15634 -9876 15651
rect -9818 15651 -9618 15698
rect -9818 15634 -9768 15651
rect -9926 15617 -9910 15634
rect -10042 15601 -9910 15617
rect -9784 15617 -9768 15634
rect -9668 15634 -9618 15651
rect -9560 15651 -9360 15698
rect -9560 15634 -9510 15651
rect -9668 15617 -9652 15634
rect -9784 15601 -9652 15617
rect -9526 15617 -9510 15634
rect -9410 15634 -9360 15651
rect -9302 15651 -9102 15698
rect -9302 15634 -9252 15651
rect -9410 15617 -9394 15634
rect -9526 15601 -9394 15617
rect -9268 15617 -9252 15634
rect -9152 15634 -9102 15651
rect -9044 15651 -8844 15698
rect -9044 15634 -8994 15651
rect -9152 15617 -9136 15634
rect -9268 15601 -9136 15617
rect -9010 15617 -8994 15634
rect -8894 15634 -8844 15651
rect -8894 15617 -8878 15634
rect -9010 15601 -8878 15617
rect -8484 15715 -8454 15741
rect -7984 15715 -7954 15741
rect -11084 15483 -11054 15515
rect -8484 15483 -8454 15515
rect -7984 15483 -7954 15515
rect -11084 15467 -10998 15483
rect -11084 15433 -11048 15467
rect -11014 15433 -10998 15467
rect -11084 15417 -10998 15433
rect -8484 15467 -8398 15483
rect -8484 15433 -8448 15467
rect -8414 15433 -8398 15467
rect -8484 15417 -8398 15433
rect -7984 15467 -7898 15483
rect -7984 15433 -7948 15467
rect -7914 15433 -7898 15467
rect -7984 15417 -7898 15433
rect -11084 15395 -11054 15417
rect -8484 15395 -8454 15417
rect -7984 15395 -7954 15417
rect -12900 15246 -12768 15262
rect -12900 15229 -12884 15246
rect -12934 15212 -12884 15229
rect -12784 15229 -12768 15246
rect -12642 15246 -12510 15262
rect -12642 15229 -12626 15246
rect -12784 15212 -12734 15229
rect -12934 15174 -12734 15212
rect -12676 15212 -12626 15229
rect -12526 15229 -12510 15246
rect -12384 15246 -12252 15262
rect -12384 15229 -12368 15246
rect -12526 15212 -12476 15229
rect -12676 15174 -12476 15212
rect -12418 15212 -12368 15229
rect -12268 15229 -12252 15246
rect -12126 15246 -11994 15262
rect -12126 15229 -12110 15246
rect -12268 15212 -12218 15229
rect -12418 15174 -12218 15212
rect -12160 15212 -12110 15229
rect -12010 15229 -11994 15246
rect -11868 15246 -11736 15262
rect -11868 15229 -11852 15246
rect -12010 15212 -11960 15229
rect -12160 15174 -11960 15212
rect -11902 15212 -11852 15229
rect -11752 15229 -11736 15246
rect -11610 15246 -11478 15262
rect -11610 15229 -11594 15246
rect -11752 15212 -11702 15229
rect -11902 15174 -11702 15212
rect -11644 15212 -11594 15229
rect -11494 15229 -11478 15246
rect -11494 15212 -11444 15229
rect -11644 15174 -11444 15212
rect -12934 14936 -12734 14974
rect -12934 14919 -12884 14936
rect -12900 14902 -12884 14919
rect -12784 14919 -12734 14936
rect -12676 14936 -12476 14974
rect -12676 14919 -12626 14936
rect -12784 14902 -12768 14919
rect -12900 14886 -12768 14902
rect -12642 14902 -12626 14919
rect -12526 14919 -12476 14936
rect -12418 14936 -12218 14974
rect -12418 14919 -12368 14936
rect -12526 14902 -12510 14919
rect -12642 14886 -12510 14902
rect -12384 14902 -12368 14919
rect -12268 14919 -12218 14936
rect -12160 14936 -11960 14974
rect -12160 14919 -12110 14936
rect -12268 14902 -12252 14919
rect -12384 14886 -12252 14902
rect -12126 14902 -12110 14919
rect -12010 14919 -11960 14936
rect -11902 14936 -11702 14974
rect -11902 14919 -11852 14936
rect -12010 14902 -11994 14919
rect -12126 14886 -11994 14902
rect -11868 14902 -11852 14919
rect -11752 14919 -11702 14936
rect -11644 14936 -11444 14974
rect -11644 14919 -11594 14936
rect -11752 14902 -11736 14919
rect -11868 14886 -11736 14902
rect -11610 14902 -11594 14919
rect -11494 14919 -11444 14936
rect -11494 14902 -11478 14919
rect -11610 14886 -11478 14902
rect -11084 15239 -11054 15265
rect -10300 15246 -10168 15262
rect -10300 15229 -10284 15246
rect -10334 15212 -10284 15229
rect -10184 15229 -10168 15246
rect -10042 15246 -9910 15262
rect -10042 15229 -10026 15246
rect -10184 15212 -10134 15229
rect -10334 15174 -10134 15212
rect -10076 15212 -10026 15229
rect -9926 15229 -9910 15246
rect -9784 15246 -9652 15262
rect -9784 15229 -9768 15246
rect -9926 15212 -9876 15229
rect -10076 15174 -9876 15212
rect -9818 15212 -9768 15229
rect -9668 15229 -9652 15246
rect -9526 15246 -9394 15262
rect -9526 15229 -9510 15246
rect -9668 15212 -9618 15229
rect -9818 15174 -9618 15212
rect -9560 15212 -9510 15229
rect -9410 15229 -9394 15246
rect -9268 15246 -9136 15262
rect -9268 15229 -9252 15246
rect -9410 15212 -9360 15229
rect -9560 15174 -9360 15212
rect -9302 15212 -9252 15229
rect -9152 15229 -9136 15246
rect -9010 15246 -8878 15262
rect -9010 15229 -8994 15246
rect -9152 15212 -9102 15229
rect -9302 15174 -9102 15212
rect -9044 15212 -8994 15229
rect -8894 15229 -8878 15246
rect -8894 15212 -8844 15229
rect -9044 15174 -8844 15212
rect -10334 14936 -10134 14974
rect -10334 14919 -10284 14936
rect -10300 14902 -10284 14919
rect -10184 14919 -10134 14936
rect -10076 14936 -9876 14974
rect -10076 14919 -10026 14936
rect -10184 14902 -10168 14919
rect -10300 14886 -10168 14902
rect -10042 14902 -10026 14919
rect -9926 14919 -9876 14936
rect -9818 14936 -9618 14974
rect -9818 14919 -9768 14936
rect -9926 14902 -9910 14919
rect -10042 14886 -9910 14902
rect -9784 14902 -9768 14919
rect -9668 14919 -9618 14936
rect -9560 14936 -9360 14974
rect -9560 14919 -9510 14936
rect -9668 14902 -9652 14919
rect -9784 14886 -9652 14902
rect -9526 14902 -9510 14919
rect -9410 14919 -9360 14936
rect -9302 14936 -9102 14974
rect -9302 14919 -9252 14936
rect -9410 14902 -9394 14919
rect -9526 14886 -9394 14902
rect -9268 14902 -9252 14919
rect -9152 14919 -9102 14936
rect -9044 14936 -8844 14974
rect -9044 14919 -8994 14936
rect -9152 14902 -9136 14919
rect -9268 14886 -9136 14902
rect -9010 14902 -8994 14919
rect -8894 14919 -8844 14936
rect -8894 14902 -8878 14919
rect -9010 14886 -8878 14902
rect -8484 15239 -8454 15265
rect -7984 15239 -7954 15265
rect 13764 14894 14352 14910
rect 13764 14877 13780 14894
rect 13578 14860 13780 14877
rect 14336 14877 14352 14894
rect 14782 14894 15370 14910
rect 14782 14877 14798 14894
rect 14336 14860 14538 14877
rect 13578 14822 14538 14860
rect 14596 14860 14798 14877
rect 15354 14877 15370 14894
rect 15800 14894 16388 14910
rect 15800 14877 15816 14894
rect 15354 14860 15556 14877
rect 14596 14822 15556 14860
rect 15614 14860 15816 14877
rect 16372 14877 16388 14894
rect 16818 14894 17406 14910
rect 16818 14877 16834 14894
rect 16372 14860 16574 14877
rect 15614 14822 16574 14860
rect 16632 14860 16834 14877
rect 17390 14877 17406 14894
rect 17836 14894 18424 14910
rect 17836 14877 17852 14894
rect 17390 14860 17592 14877
rect 16632 14822 17592 14860
rect 17650 14860 17852 14877
rect 18408 14877 18424 14894
rect 18854 14894 19442 14910
rect 18854 14877 18870 14894
rect 18408 14860 18610 14877
rect 17650 14822 18610 14860
rect 18668 14860 18870 14877
rect 19426 14877 19442 14894
rect 19872 14894 20460 14910
rect 19872 14877 19888 14894
rect 19426 14860 19628 14877
rect 18668 14822 19628 14860
rect 19686 14860 19888 14877
rect 20444 14877 20460 14894
rect 20890 14894 21478 14910
rect 20890 14877 20906 14894
rect 20444 14860 20646 14877
rect 19686 14822 20646 14860
rect 20704 14860 20906 14877
rect 21462 14877 21478 14894
rect 21908 14894 22496 14910
rect 21908 14877 21924 14894
rect 21462 14860 21664 14877
rect 20704 14822 21664 14860
rect 21722 14860 21924 14877
rect 22480 14877 22496 14894
rect 22926 14894 23514 14910
rect 22926 14877 22942 14894
rect 22480 14860 22682 14877
rect 21722 14822 22682 14860
rect 22740 14860 22942 14877
rect 23498 14877 23514 14894
rect 23944 14894 24532 14910
rect 23944 14877 23960 14894
rect 23498 14860 23700 14877
rect 22740 14822 23700 14860
rect 23758 14860 23960 14877
rect 24516 14877 24532 14894
rect 24962 14894 25550 14910
rect 24962 14877 24978 14894
rect 24516 14860 24718 14877
rect 23758 14822 24718 14860
rect 24776 14860 24978 14877
rect 25534 14877 25550 14894
rect 25980 14894 26568 14910
rect 25980 14877 25996 14894
rect 25534 14860 25736 14877
rect 24776 14822 25736 14860
rect 25794 14860 25996 14877
rect 26552 14877 26568 14894
rect 26998 14894 27586 14910
rect 26998 14877 27014 14894
rect 26552 14860 26754 14877
rect 25794 14822 26754 14860
rect 26812 14860 27014 14877
rect 27570 14877 27586 14894
rect 28016 14894 28604 14910
rect 28016 14877 28032 14894
rect 27570 14860 27772 14877
rect 26812 14822 27772 14860
rect 27830 14860 28032 14877
rect 28588 14877 28604 14894
rect 29034 14894 29622 14910
rect 29034 14877 29050 14894
rect 28588 14860 28790 14877
rect 27830 14822 28790 14860
rect 28848 14860 29050 14877
rect 29606 14877 29622 14894
rect 30052 14894 30640 14910
rect 30052 14877 30068 14894
rect 29606 14860 29808 14877
rect 28848 14822 29808 14860
rect 29866 14860 30068 14877
rect 30624 14877 30640 14894
rect 31070 14894 31658 14910
rect 31070 14877 31086 14894
rect 30624 14860 30826 14877
rect 29866 14822 30826 14860
rect 30884 14860 31086 14877
rect 31642 14877 31658 14894
rect 32088 14894 32676 14910
rect 32088 14877 32104 14894
rect 31642 14860 31844 14877
rect 30884 14822 31844 14860
rect 31902 14860 32104 14877
rect 32660 14877 32676 14894
rect 33106 14894 33694 14910
rect 33106 14877 33122 14894
rect 32660 14860 32862 14877
rect 31902 14822 32862 14860
rect 32920 14860 33122 14877
rect 33678 14877 33694 14894
rect 33678 14860 33880 14877
rect 32920 14822 33880 14860
rect 13578 14184 14538 14222
rect 13578 14167 13780 14184
rect 13764 14150 13780 14167
rect 14336 14167 14538 14184
rect 14596 14184 15556 14222
rect 14596 14167 14798 14184
rect 14336 14150 14352 14167
rect 13764 14134 14352 14150
rect 14782 14150 14798 14167
rect 15354 14167 15556 14184
rect 15614 14184 16574 14222
rect 15614 14167 15816 14184
rect 15354 14150 15370 14167
rect 14782 14134 15370 14150
rect 15800 14150 15816 14167
rect 16372 14167 16574 14184
rect 16632 14184 17592 14222
rect 16632 14167 16834 14184
rect 16372 14150 16388 14167
rect 15800 14134 16388 14150
rect 16818 14150 16834 14167
rect 17390 14167 17592 14184
rect 17650 14184 18610 14222
rect 17650 14167 17852 14184
rect 17390 14150 17406 14167
rect 16818 14134 17406 14150
rect 17836 14150 17852 14167
rect 18408 14167 18610 14184
rect 18668 14184 19628 14222
rect 18668 14167 18870 14184
rect 18408 14150 18424 14167
rect 17836 14134 18424 14150
rect 18854 14150 18870 14167
rect 19426 14167 19628 14184
rect 19686 14184 20646 14222
rect 19686 14167 19888 14184
rect 19426 14150 19442 14167
rect 18854 14134 19442 14150
rect 19872 14150 19888 14167
rect 20444 14167 20646 14184
rect 20704 14184 21664 14222
rect 20704 14167 20906 14184
rect 20444 14150 20460 14167
rect 19872 14134 20460 14150
rect 20890 14150 20906 14167
rect 21462 14167 21664 14184
rect 21722 14184 22682 14222
rect 21722 14167 21924 14184
rect 21462 14150 21478 14167
rect 20890 14134 21478 14150
rect 21908 14150 21924 14167
rect 22480 14167 22682 14184
rect 22740 14184 23700 14222
rect 22740 14167 22942 14184
rect 22480 14150 22496 14167
rect 21908 14134 22496 14150
rect 22926 14150 22942 14167
rect 23498 14167 23700 14184
rect 23758 14184 24718 14222
rect 23758 14167 23960 14184
rect 23498 14150 23514 14167
rect 22926 14134 23514 14150
rect 23944 14150 23960 14167
rect 24516 14167 24718 14184
rect 24776 14184 25736 14222
rect 24776 14167 24978 14184
rect 24516 14150 24532 14167
rect 23944 14134 24532 14150
rect 24962 14150 24978 14167
rect 25534 14167 25736 14184
rect 25794 14184 26754 14222
rect 25794 14167 25996 14184
rect 25534 14150 25550 14167
rect 24962 14134 25550 14150
rect 25980 14150 25996 14167
rect 26552 14167 26754 14184
rect 26812 14184 27772 14222
rect 26812 14167 27014 14184
rect 26552 14150 26568 14167
rect 25980 14134 26568 14150
rect 26998 14150 27014 14167
rect 27570 14167 27772 14184
rect 27830 14184 28790 14222
rect 27830 14167 28032 14184
rect 27570 14150 27586 14167
rect 26998 14134 27586 14150
rect 28016 14150 28032 14167
rect 28588 14167 28790 14184
rect 28848 14184 29808 14222
rect 28848 14167 29050 14184
rect 28588 14150 28604 14167
rect 28016 14134 28604 14150
rect 29034 14150 29050 14167
rect 29606 14167 29808 14184
rect 29866 14184 30826 14222
rect 29866 14167 30068 14184
rect 29606 14150 29622 14167
rect 29034 14134 29622 14150
rect 30052 14150 30068 14167
rect 30624 14167 30826 14184
rect 30884 14184 31844 14222
rect 30884 14167 31086 14184
rect 30624 14150 30640 14167
rect 30052 14134 30640 14150
rect 31070 14150 31086 14167
rect 31642 14167 31844 14184
rect 31902 14184 32862 14222
rect 31902 14167 32104 14184
rect 31642 14150 31658 14167
rect 31070 14134 31658 14150
rect 32088 14150 32104 14167
rect 32660 14167 32862 14184
rect 32920 14184 33880 14222
rect 32920 14167 33122 14184
rect 32660 14150 32676 14167
rect 32088 14134 32676 14150
rect 33106 14150 33122 14167
rect 33678 14167 33880 14184
rect 33678 14150 33694 14167
rect 33106 14134 33694 14150
rect 1998 14100 2586 14116
rect 1998 14083 2014 14100
rect 1812 14066 2014 14083
rect 2570 14083 2586 14100
rect 3016 14100 3604 14116
rect 3016 14083 3032 14100
rect 2570 14066 2772 14083
rect 1812 14028 2772 14066
rect 2830 14066 3032 14083
rect 3588 14083 3604 14100
rect 4034 14100 4622 14116
rect 4034 14083 4050 14100
rect 3588 14066 3790 14083
rect 2830 14028 3790 14066
rect 3848 14066 4050 14083
rect 4606 14083 4622 14100
rect 5052 14100 5640 14116
rect 5052 14083 5068 14100
rect 4606 14066 4808 14083
rect 3848 14028 4808 14066
rect 4866 14066 5068 14083
rect 5624 14083 5640 14100
rect 6070 14100 6658 14116
rect 6070 14083 6086 14100
rect 5624 14066 5826 14083
rect 4866 14028 5826 14066
rect 5884 14066 6086 14083
rect 6642 14083 6658 14100
rect 7088 14100 7676 14116
rect 7088 14083 7104 14100
rect 6642 14066 6844 14083
rect 5884 14028 6844 14066
rect 6902 14066 7104 14083
rect 7660 14083 7676 14100
rect 8106 14100 8694 14116
rect 8106 14083 8122 14100
rect 7660 14066 7862 14083
rect 6902 14028 7862 14066
rect 7920 14066 8122 14083
rect 8678 14083 8694 14100
rect 9124 14100 9712 14116
rect 9124 14083 9140 14100
rect 8678 14066 8880 14083
rect 7920 14028 8880 14066
rect 8938 14066 9140 14083
rect 9696 14083 9712 14100
rect 10142 14100 10730 14116
rect 10142 14083 10158 14100
rect 9696 14066 9898 14083
rect 8938 14028 9898 14066
rect 9956 14066 10158 14083
rect 10714 14083 10730 14100
rect 10714 14066 10916 14083
rect 9956 14028 10916 14066
rect 13764 13660 14352 13676
rect 13764 13643 13780 13660
rect 13578 13626 13780 13643
rect 14336 13643 14352 13660
rect 14782 13660 15370 13676
rect 14782 13643 14798 13660
rect 14336 13626 14538 13643
rect 13578 13588 14538 13626
rect 14596 13626 14798 13643
rect 15354 13643 15370 13660
rect 15800 13660 16388 13676
rect 15800 13643 15816 13660
rect 15354 13626 15556 13643
rect 14596 13588 15556 13626
rect 15614 13626 15816 13643
rect 16372 13643 16388 13660
rect 16818 13660 17406 13676
rect 16818 13643 16834 13660
rect 16372 13626 16574 13643
rect 15614 13588 16574 13626
rect 16632 13626 16834 13643
rect 17390 13643 17406 13660
rect 17836 13660 18424 13676
rect 17836 13643 17852 13660
rect 17390 13626 17592 13643
rect 16632 13588 17592 13626
rect 17650 13626 17852 13643
rect 18408 13643 18424 13660
rect 18854 13660 19442 13676
rect 18854 13643 18870 13660
rect 18408 13626 18610 13643
rect 17650 13588 18610 13626
rect 18668 13626 18870 13643
rect 19426 13643 19442 13660
rect 19872 13660 20460 13676
rect 19872 13643 19888 13660
rect 19426 13626 19628 13643
rect 18668 13588 19628 13626
rect 19686 13626 19888 13643
rect 20444 13643 20460 13660
rect 20890 13660 21478 13676
rect 20890 13643 20906 13660
rect 20444 13626 20646 13643
rect 19686 13588 20646 13626
rect 20704 13626 20906 13643
rect 21462 13643 21478 13660
rect 21908 13660 22496 13676
rect 21908 13643 21924 13660
rect 21462 13626 21664 13643
rect 20704 13588 21664 13626
rect 21722 13626 21924 13643
rect 22480 13643 22496 13660
rect 22926 13660 23514 13676
rect 22926 13643 22942 13660
rect 22480 13626 22682 13643
rect 21722 13588 22682 13626
rect 22740 13626 22942 13643
rect 23498 13643 23514 13660
rect 23944 13660 24532 13676
rect 23944 13643 23960 13660
rect 23498 13626 23700 13643
rect 22740 13588 23700 13626
rect 23758 13626 23960 13643
rect 24516 13643 24532 13660
rect 24962 13660 25550 13676
rect 24962 13643 24978 13660
rect 24516 13626 24718 13643
rect 23758 13588 24718 13626
rect 24776 13626 24978 13643
rect 25534 13643 25550 13660
rect 25980 13660 26568 13676
rect 25980 13643 25996 13660
rect 25534 13626 25736 13643
rect 24776 13588 25736 13626
rect 25794 13626 25996 13643
rect 26552 13643 26568 13660
rect 26998 13660 27586 13676
rect 26998 13643 27014 13660
rect 26552 13626 26754 13643
rect 25794 13588 26754 13626
rect 26812 13626 27014 13643
rect 27570 13643 27586 13660
rect 28016 13660 28604 13676
rect 28016 13643 28032 13660
rect 27570 13626 27772 13643
rect 26812 13588 27772 13626
rect 27830 13626 28032 13643
rect 28588 13643 28604 13660
rect 29034 13660 29622 13676
rect 29034 13643 29050 13660
rect 28588 13626 28790 13643
rect 27830 13588 28790 13626
rect 28848 13626 29050 13643
rect 29606 13643 29622 13660
rect 30052 13660 30640 13676
rect 30052 13643 30068 13660
rect 29606 13626 29808 13643
rect 28848 13588 29808 13626
rect 29866 13626 30068 13643
rect 30624 13643 30640 13660
rect 31070 13660 31658 13676
rect 31070 13643 31086 13660
rect 30624 13626 30826 13643
rect 29866 13588 30826 13626
rect 30884 13626 31086 13643
rect 31642 13643 31658 13660
rect 32088 13660 32676 13676
rect 32088 13643 32104 13660
rect 31642 13626 31844 13643
rect 30884 13588 31844 13626
rect 31902 13626 32104 13643
rect 32660 13643 32676 13660
rect 33106 13660 33694 13676
rect 33106 13643 33122 13660
rect 32660 13626 32862 13643
rect 31902 13588 32862 13626
rect 32920 13626 33122 13643
rect 33678 13643 33694 13660
rect 33678 13626 33880 13643
rect 32920 13588 33880 13626
rect 1812 13390 2772 13428
rect 1812 13373 2014 13390
rect 1998 13356 2014 13373
rect 2570 13373 2772 13390
rect 2830 13390 3790 13428
rect 2830 13373 3032 13390
rect 2570 13356 2586 13373
rect 1998 13340 2586 13356
rect 3016 13356 3032 13373
rect 3588 13373 3790 13390
rect 3848 13390 4808 13428
rect 3848 13373 4050 13390
rect 3588 13356 3604 13373
rect 3016 13340 3604 13356
rect 1998 13282 2586 13298
rect 1998 13265 2014 13282
rect 1812 13248 2014 13265
rect 2570 13265 2586 13282
rect 4034 13356 4050 13373
rect 4606 13373 4808 13390
rect 4866 13390 5826 13428
rect 4866 13373 5068 13390
rect 4606 13356 4622 13373
rect 4034 13340 4622 13356
rect 3016 13282 3604 13298
rect 3016 13265 3032 13282
rect 2570 13248 2772 13265
rect 1812 13210 2772 13248
rect 2830 13248 3032 13265
rect 3588 13265 3604 13282
rect 5052 13356 5068 13373
rect 5624 13373 5826 13390
rect 5884 13390 6844 13428
rect 5884 13373 6086 13390
rect 5624 13356 5640 13373
rect 5052 13340 5640 13356
rect 4034 13282 4622 13298
rect 4034 13265 4050 13282
rect 3588 13248 3790 13265
rect 2830 13210 3790 13248
rect 3848 13248 4050 13265
rect 4606 13265 4622 13282
rect 6070 13356 6086 13373
rect 6642 13373 6844 13390
rect 6902 13390 7862 13428
rect 6902 13373 7104 13390
rect 6642 13356 6658 13373
rect 6070 13340 6658 13356
rect 5052 13282 5640 13298
rect 5052 13265 5068 13282
rect 4606 13248 4808 13265
rect 3848 13210 4808 13248
rect 4866 13248 5068 13265
rect 5624 13265 5640 13282
rect 7088 13356 7104 13373
rect 7660 13373 7862 13390
rect 7920 13390 8880 13428
rect 7920 13373 8122 13390
rect 7660 13356 7676 13373
rect 7088 13340 7676 13356
rect 6070 13282 6658 13298
rect 6070 13265 6086 13282
rect 5624 13248 5826 13265
rect 4866 13210 5826 13248
rect 5884 13248 6086 13265
rect 6642 13265 6658 13282
rect 8106 13356 8122 13373
rect 8678 13373 8880 13390
rect 8938 13390 9898 13428
rect 8938 13373 9140 13390
rect 8678 13356 8694 13373
rect 8106 13340 8694 13356
rect 7088 13282 7676 13298
rect 7088 13265 7104 13282
rect 6642 13248 6844 13265
rect 5884 13210 6844 13248
rect 6902 13248 7104 13265
rect 7660 13265 7676 13282
rect 9124 13356 9140 13373
rect 9696 13373 9898 13390
rect 9956 13390 10916 13428
rect 9956 13373 10158 13390
rect 9696 13356 9712 13373
rect 9124 13340 9712 13356
rect 8106 13282 8694 13298
rect 8106 13265 8122 13282
rect 7660 13248 7862 13265
rect 6902 13210 7862 13248
rect 7920 13248 8122 13265
rect 8678 13265 8694 13282
rect 10142 13356 10158 13373
rect 10714 13373 10916 13390
rect 10714 13356 10730 13373
rect 10142 13340 10730 13356
rect 9124 13282 9712 13298
rect 9124 13265 9140 13282
rect 8678 13248 8880 13265
rect 7920 13210 8880 13248
rect 8938 13248 9140 13265
rect 9696 13265 9712 13282
rect 10142 13282 10730 13298
rect 10142 13265 10158 13282
rect 9696 13248 9898 13265
rect 8938 13210 9898 13248
rect 9956 13248 10158 13265
rect 10714 13265 10730 13282
rect 10714 13248 10916 13265
rect 9956 13210 10916 13248
rect 13578 12950 14538 12988
rect 13578 12933 13780 12950
rect 13764 12916 13780 12933
rect 14336 12933 14538 12950
rect 14596 12950 15556 12988
rect 14596 12933 14798 12950
rect 14336 12916 14352 12933
rect 13764 12900 14352 12916
rect 14782 12916 14798 12933
rect 15354 12933 15556 12950
rect 15614 12950 16574 12988
rect 15614 12933 15816 12950
rect 15354 12916 15370 12933
rect 14782 12900 15370 12916
rect 15800 12916 15816 12933
rect 16372 12933 16574 12950
rect 16632 12950 17592 12988
rect 16632 12933 16834 12950
rect 16372 12916 16388 12933
rect 15800 12900 16388 12916
rect 16818 12916 16834 12933
rect 17390 12933 17592 12950
rect 17650 12950 18610 12988
rect 17650 12933 17852 12950
rect 17390 12916 17406 12933
rect 16818 12900 17406 12916
rect 17836 12916 17852 12933
rect 18408 12933 18610 12950
rect 18668 12950 19628 12988
rect 18668 12933 18870 12950
rect 18408 12916 18424 12933
rect 17836 12900 18424 12916
rect 18854 12916 18870 12933
rect 19426 12933 19628 12950
rect 19686 12950 20646 12988
rect 19686 12933 19888 12950
rect 19426 12916 19442 12933
rect 18854 12900 19442 12916
rect 19872 12916 19888 12933
rect 20444 12933 20646 12950
rect 20704 12950 21664 12988
rect 20704 12933 20906 12950
rect 20444 12916 20460 12933
rect 19872 12900 20460 12916
rect 20890 12916 20906 12933
rect 21462 12933 21664 12950
rect 21722 12950 22682 12988
rect 21722 12933 21924 12950
rect 21462 12916 21478 12933
rect 20890 12900 21478 12916
rect 21908 12916 21924 12933
rect 22480 12933 22682 12950
rect 22740 12950 23700 12988
rect 22740 12933 22942 12950
rect 22480 12916 22496 12933
rect 21908 12900 22496 12916
rect 22926 12916 22942 12933
rect 23498 12933 23700 12950
rect 23758 12950 24718 12988
rect 23758 12933 23960 12950
rect 23498 12916 23514 12933
rect 22926 12900 23514 12916
rect 23944 12916 23960 12933
rect 24516 12933 24718 12950
rect 24776 12950 25736 12988
rect 24776 12933 24978 12950
rect 24516 12916 24532 12933
rect 23944 12900 24532 12916
rect 24962 12916 24978 12933
rect 25534 12933 25736 12950
rect 25794 12950 26754 12988
rect 25794 12933 25996 12950
rect 25534 12916 25550 12933
rect 24962 12900 25550 12916
rect 25980 12916 25996 12933
rect 26552 12933 26754 12950
rect 26812 12950 27772 12988
rect 26812 12933 27014 12950
rect 26552 12916 26568 12933
rect 25980 12900 26568 12916
rect 26998 12916 27014 12933
rect 27570 12933 27772 12950
rect 27830 12950 28790 12988
rect 27830 12933 28032 12950
rect 27570 12916 27586 12933
rect 26998 12900 27586 12916
rect 28016 12916 28032 12933
rect 28588 12933 28790 12950
rect 28848 12950 29808 12988
rect 28848 12933 29050 12950
rect 28588 12916 28604 12933
rect 28016 12900 28604 12916
rect 29034 12916 29050 12933
rect 29606 12933 29808 12950
rect 29866 12950 30826 12988
rect 29866 12933 30068 12950
rect 29606 12916 29622 12933
rect 29034 12900 29622 12916
rect 30052 12916 30068 12933
rect 30624 12933 30826 12950
rect 30884 12950 31844 12988
rect 30884 12933 31086 12950
rect 30624 12916 30640 12933
rect 30052 12900 30640 12916
rect 31070 12916 31086 12933
rect 31642 12933 31844 12950
rect 31902 12950 32862 12988
rect 31902 12933 32104 12950
rect 31642 12916 31658 12933
rect 31070 12900 31658 12916
rect 32088 12916 32104 12933
rect 32660 12933 32862 12950
rect 32920 12950 33880 12988
rect 32920 12933 33122 12950
rect 32660 12916 32676 12933
rect 32088 12900 32676 12916
rect 33106 12916 33122 12933
rect 33678 12933 33880 12950
rect 33678 12916 33694 12933
rect 33106 12900 33694 12916
rect 1812 12572 2772 12610
rect 1812 12555 2014 12572
rect 1998 12538 2014 12555
rect 2570 12555 2772 12572
rect 2830 12572 3790 12610
rect 2830 12555 3032 12572
rect 2570 12538 2586 12555
rect 1998 12522 2586 12538
rect 3016 12538 3032 12555
rect 3588 12555 3790 12572
rect 3848 12572 4808 12610
rect 3848 12555 4050 12572
rect 3588 12538 3604 12555
rect 3016 12522 3604 12538
rect 1998 12464 2586 12480
rect 1998 12447 2014 12464
rect 1812 12430 2014 12447
rect 2570 12447 2586 12464
rect 4034 12538 4050 12555
rect 4606 12555 4808 12572
rect 4866 12572 5826 12610
rect 4866 12555 5068 12572
rect 4606 12538 4622 12555
rect 4034 12522 4622 12538
rect 3016 12464 3604 12480
rect 3016 12447 3032 12464
rect 2570 12430 2772 12447
rect 1812 12392 2772 12430
rect 2830 12430 3032 12447
rect 3588 12447 3604 12464
rect 5052 12538 5068 12555
rect 5624 12555 5826 12572
rect 5884 12572 6844 12610
rect 5884 12555 6086 12572
rect 5624 12538 5640 12555
rect 5052 12522 5640 12538
rect 4034 12464 4622 12480
rect 4034 12447 4050 12464
rect 3588 12430 3790 12447
rect 2830 12392 3790 12430
rect 3848 12430 4050 12447
rect 4606 12447 4622 12464
rect 6070 12538 6086 12555
rect 6642 12555 6844 12572
rect 6902 12572 7862 12610
rect 6902 12555 7104 12572
rect 6642 12538 6658 12555
rect 6070 12522 6658 12538
rect 5052 12464 5640 12480
rect 5052 12447 5068 12464
rect 4606 12430 4808 12447
rect 3848 12392 4808 12430
rect 4866 12430 5068 12447
rect 5624 12447 5640 12464
rect 7088 12538 7104 12555
rect 7660 12555 7862 12572
rect 7920 12572 8880 12610
rect 7920 12555 8122 12572
rect 7660 12538 7676 12555
rect 7088 12522 7676 12538
rect 6070 12464 6658 12480
rect 6070 12447 6086 12464
rect 5624 12430 5826 12447
rect 4866 12392 5826 12430
rect 5884 12430 6086 12447
rect 6642 12447 6658 12464
rect 8106 12538 8122 12555
rect 8678 12555 8880 12572
rect 8938 12572 9898 12610
rect 8938 12555 9140 12572
rect 8678 12538 8694 12555
rect 8106 12522 8694 12538
rect 7088 12464 7676 12480
rect 7088 12447 7104 12464
rect 6642 12430 6844 12447
rect 5884 12392 6844 12430
rect 6902 12430 7104 12447
rect 7660 12447 7676 12464
rect 9124 12538 9140 12555
rect 9696 12555 9898 12572
rect 9956 12572 10916 12610
rect 9956 12555 10158 12572
rect 9696 12538 9712 12555
rect 9124 12522 9712 12538
rect 8106 12464 8694 12480
rect 8106 12447 8122 12464
rect 7660 12430 7862 12447
rect 6902 12392 7862 12430
rect 7920 12430 8122 12447
rect 8678 12447 8694 12464
rect 10142 12538 10158 12555
rect 10714 12555 10916 12572
rect 10714 12538 10730 12555
rect 10142 12522 10730 12538
rect 9124 12464 9712 12480
rect 9124 12447 9140 12464
rect 8678 12430 8880 12447
rect 7920 12392 8880 12430
rect 8938 12430 9140 12447
rect 9696 12447 9712 12464
rect 10142 12464 10730 12480
rect 10142 12447 10158 12464
rect 9696 12430 9898 12447
rect 8938 12392 9898 12430
rect 9956 12430 10158 12447
rect 10714 12447 10730 12464
rect 10714 12430 10916 12447
rect 9956 12392 10916 12430
rect 13764 12428 14352 12444
rect 13764 12411 13780 12428
rect 13578 12394 13780 12411
rect 14336 12411 14352 12428
rect 14782 12428 15370 12444
rect 14782 12411 14798 12428
rect 14336 12394 14538 12411
rect 13578 12356 14538 12394
rect 14596 12394 14798 12411
rect 15354 12411 15370 12428
rect 15800 12428 16388 12444
rect 15800 12411 15816 12428
rect 15354 12394 15556 12411
rect 14596 12356 15556 12394
rect 15614 12394 15816 12411
rect 16372 12411 16388 12428
rect 16818 12428 17406 12444
rect 16818 12411 16834 12428
rect 16372 12394 16574 12411
rect 15614 12356 16574 12394
rect 16632 12394 16834 12411
rect 17390 12411 17406 12428
rect 17836 12428 18424 12444
rect 17836 12411 17852 12428
rect 17390 12394 17592 12411
rect 16632 12356 17592 12394
rect 17650 12394 17852 12411
rect 18408 12411 18424 12428
rect 18854 12428 19442 12444
rect 18854 12411 18870 12428
rect 18408 12394 18610 12411
rect 17650 12356 18610 12394
rect 18668 12394 18870 12411
rect 19426 12411 19442 12428
rect 19872 12428 20460 12444
rect 19872 12411 19888 12428
rect 19426 12394 19628 12411
rect 18668 12356 19628 12394
rect 19686 12394 19888 12411
rect 20444 12411 20460 12428
rect 20890 12428 21478 12444
rect 20890 12411 20906 12428
rect 20444 12394 20646 12411
rect 19686 12356 20646 12394
rect 20704 12394 20906 12411
rect 21462 12411 21478 12428
rect 21908 12428 22496 12444
rect 21908 12411 21924 12428
rect 21462 12394 21664 12411
rect 20704 12356 21664 12394
rect 21722 12394 21924 12411
rect 22480 12411 22496 12428
rect 22926 12428 23514 12444
rect 22926 12411 22942 12428
rect 22480 12394 22682 12411
rect 21722 12356 22682 12394
rect 22740 12394 22942 12411
rect 23498 12411 23514 12428
rect 23944 12428 24532 12444
rect 23944 12411 23960 12428
rect 23498 12394 23700 12411
rect 22740 12356 23700 12394
rect 23758 12394 23960 12411
rect 24516 12411 24532 12428
rect 24962 12428 25550 12444
rect 24962 12411 24978 12428
rect 24516 12394 24718 12411
rect 23758 12356 24718 12394
rect 24776 12394 24978 12411
rect 25534 12411 25550 12428
rect 25980 12428 26568 12444
rect 25980 12411 25996 12428
rect 25534 12394 25736 12411
rect 24776 12356 25736 12394
rect 25794 12394 25996 12411
rect 26552 12411 26568 12428
rect 26998 12428 27586 12444
rect 26998 12411 27014 12428
rect 26552 12394 26754 12411
rect 25794 12356 26754 12394
rect 26812 12394 27014 12411
rect 27570 12411 27586 12428
rect 28016 12428 28604 12444
rect 28016 12411 28032 12428
rect 27570 12394 27772 12411
rect 26812 12356 27772 12394
rect 27830 12394 28032 12411
rect 28588 12411 28604 12428
rect 29034 12428 29622 12444
rect 29034 12411 29050 12428
rect 28588 12394 28790 12411
rect 27830 12356 28790 12394
rect 28848 12394 29050 12411
rect 29606 12411 29622 12428
rect 30052 12428 30640 12444
rect 30052 12411 30068 12428
rect 29606 12394 29808 12411
rect 28848 12356 29808 12394
rect 29866 12394 30068 12411
rect 30624 12411 30640 12428
rect 31070 12428 31658 12444
rect 31070 12411 31086 12428
rect 30624 12394 30826 12411
rect 29866 12356 30826 12394
rect 30884 12394 31086 12411
rect 31642 12411 31658 12428
rect 32088 12428 32676 12444
rect 32088 12411 32104 12428
rect 31642 12394 31844 12411
rect 30884 12356 31844 12394
rect 31902 12394 32104 12411
rect 32660 12411 32676 12428
rect 33106 12428 33694 12444
rect 33106 12411 33122 12428
rect 32660 12394 32862 12411
rect 31902 12356 32862 12394
rect 32920 12394 33122 12411
rect 33678 12411 33694 12428
rect 33678 12394 33880 12411
rect 32920 12356 33880 12394
rect 1812 11754 2772 11792
rect 1812 11737 2014 11754
rect 1998 11720 2014 11737
rect 2570 11737 2772 11754
rect 2830 11754 3790 11792
rect 2830 11737 3032 11754
rect 2570 11720 2586 11737
rect 1998 11704 2586 11720
rect 3016 11720 3032 11737
rect 3588 11737 3790 11754
rect 3848 11754 4808 11792
rect 3848 11737 4050 11754
rect 3588 11720 3604 11737
rect 3016 11704 3604 11720
rect 1998 11646 2586 11662
rect 1998 11629 2014 11646
rect 1812 11612 2014 11629
rect 2570 11629 2586 11646
rect 4034 11720 4050 11737
rect 4606 11737 4808 11754
rect 4866 11754 5826 11792
rect 4866 11737 5068 11754
rect 4606 11720 4622 11737
rect 4034 11704 4622 11720
rect 3016 11646 3604 11662
rect 3016 11629 3032 11646
rect 2570 11612 2772 11629
rect 1812 11574 2772 11612
rect 2830 11612 3032 11629
rect 3588 11629 3604 11646
rect 5052 11720 5068 11737
rect 5624 11737 5826 11754
rect 5884 11754 6844 11792
rect 5884 11737 6086 11754
rect 5624 11720 5640 11737
rect 5052 11704 5640 11720
rect 4034 11646 4622 11662
rect 4034 11629 4050 11646
rect 3588 11612 3790 11629
rect 2830 11574 3790 11612
rect 3848 11612 4050 11629
rect 4606 11629 4622 11646
rect 6070 11720 6086 11737
rect 6642 11737 6844 11754
rect 6902 11754 7862 11792
rect 6902 11737 7104 11754
rect 6642 11720 6658 11737
rect 6070 11704 6658 11720
rect 5052 11646 5640 11662
rect 5052 11629 5068 11646
rect 4606 11612 4808 11629
rect 3848 11574 4808 11612
rect 4866 11612 5068 11629
rect 5624 11629 5640 11646
rect 7088 11720 7104 11737
rect 7660 11737 7862 11754
rect 7920 11754 8880 11792
rect 7920 11737 8122 11754
rect 7660 11720 7676 11737
rect 7088 11704 7676 11720
rect 6070 11646 6658 11662
rect 6070 11629 6086 11646
rect 5624 11612 5826 11629
rect 4866 11574 5826 11612
rect 5884 11612 6086 11629
rect 6642 11629 6658 11646
rect 8106 11720 8122 11737
rect 8678 11737 8880 11754
rect 8938 11754 9898 11792
rect 8938 11737 9140 11754
rect 8678 11720 8694 11737
rect 8106 11704 8694 11720
rect 7088 11646 7676 11662
rect 7088 11629 7104 11646
rect 6642 11612 6844 11629
rect 5884 11574 6844 11612
rect 6902 11612 7104 11629
rect 7660 11629 7676 11646
rect 9124 11720 9140 11737
rect 9696 11737 9898 11754
rect 9956 11754 10916 11792
rect 9956 11737 10158 11754
rect 9696 11720 9712 11737
rect 9124 11704 9712 11720
rect 8106 11646 8694 11662
rect 8106 11629 8122 11646
rect 7660 11612 7862 11629
rect 6902 11574 7862 11612
rect 7920 11612 8122 11629
rect 8678 11629 8694 11646
rect 10142 11720 10158 11737
rect 10714 11737 10916 11754
rect 10714 11720 10730 11737
rect 10142 11704 10730 11720
rect 9124 11646 9712 11662
rect 9124 11629 9140 11646
rect 8678 11612 8880 11629
rect 7920 11574 8880 11612
rect 8938 11612 9140 11629
rect 9696 11629 9712 11646
rect 13578 11718 14538 11756
rect 13578 11701 13780 11718
rect 13764 11684 13780 11701
rect 14336 11701 14538 11718
rect 14596 11718 15556 11756
rect 14596 11701 14798 11718
rect 14336 11684 14352 11701
rect 13764 11668 14352 11684
rect 14782 11684 14798 11701
rect 15354 11701 15556 11718
rect 15614 11718 16574 11756
rect 15614 11701 15816 11718
rect 15354 11684 15370 11701
rect 14782 11668 15370 11684
rect 15800 11684 15816 11701
rect 16372 11701 16574 11718
rect 16632 11718 17592 11756
rect 16632 11701 16834 11718
rect 16372 11684 16388 11701
rect 15800 11668 16388 11684
rect 16818 11684 16834 11701
rect 17390 11701 17592 11718
rect 17650 11718 18610 11756
rect 17650 11701 17852 11718
rect 17390 11684 17406 11701
rect 16818 11668 17406 11684
rect 17836 11684 17852 11701
rect 18408 11701 18610 11718
rect 18668 11718 19628 11756
rect 18668 11701 18870 11718
rect 18408 11684 18424 11701
rect 17836 11668 18424 11684
rect 18854 11684 18870 11701
rect 19426 11701 19628 11718
rect 19686 11718 20646 11756
rect 19686 11701 19888 11718
rect 19426 11684 19442 11701
rect 18854 11668 19442 11684
rect 19872 11684 19888 11701
rect 20444 11701 20646 11718
rect 20704 11718 21664 11756
rect 20704 11701 20906 11718
rect 20444 11684 20460 11701
rect 19872 11668 20460 11684
rect 20890 11684 20906 11701
rect 21462 11701 21664 11718
rect 21722 11718 22682 11756
rect 21722 11701 21924 11718
rect 21462 11684 21478 11701
rect 20890 11668 21478 11684
rect 21908 11684 21924 11701
rect 22480 11701 22682 11718
rect 22740 11718 23700 11756
rect 22740 11701 22942 11718
rect 22480 11684 22496 11701
rect 21908 11668 22496 11684
rect 22926 11684 22942 11701
rect 23498 11701 23700 11718
rect 23758 11718 24718 11756
rect 23758 11701 23960 11718
rect 23498 11684 23514 11701
rect 22926 11668 23514 11684
rect 23944 11684 23960 11701
rect 24516 11701 24718 11718
rect 24776 11718 25736 11756
rect 24776 11701 24978 11718
rect 24516 11684 24532 11701
rect 23944 11668 24532 11684
rect 24962 11684 24978 11701
rect 25534 11701 25736 11718
rect 25794 11718 26754 11756
rect 25794 11701 25996 11718
rect 25534 11684 25550 11701
rect 24962 11668 25550 11684
rect 25980 11684 25996 11701
rect 26552 11701 26754 11718
rect 26812 11718 27772 11756
rect 26812 11701 27014 11718
rect 26552 11684 26568 11701
rect 25980 11668 26568 11684
rect 26998 11684 27014 11701
rect 27570 11701 27772 11718
rect 27830 11718 28790 11756
rect 27830 11701 28032 11718
rect 27570 11684 27586 11701
rect 26998 11668 27586 11684
rect 28016 11684 28032 11701
rect 28588 11701 28790 11718
rect 28848 11718 29808 11756
rect 28848 11701 29050 11718
rect 28588 11684 28604 11701
rect 28016 11668 28604 11684
rect 29034 11684 29050 11701
rect 29606 11701 29808 11718
rect 29866 11718 30826 11756
rect 29866 11701 30068 11718
rect 29606 11684 29622 11701
rect 29034 11668 29622 11684
rect 30052 11684 30068 11701
rect 30624 11701 30826 11718
rect 30884 11718 31844 11756
rect 30884 11701 31086 11718
rect 30624 11684 30640 11701
rect 30052 11668 30640 11684
rect 31070 11684 31086 11701
rect 31642 11701 31844 11718
rect 31902 11718 32862 11756
rect 31902 11701 32104 11718
rect 31642 11684 31658 11701
rect 31070 11668 31658 11684
rect 32088 11684 32104 11701
rect 32660 11701 32862 11718
rect 32920 11718 33880 11756
rect 32920 11701 33122 11718
rect 32660 11684 32676 11701
rect 32088 11668 32676 11684
rect 33106 11684 33122 11701
rect 33678 11701 33880 11718
rect 33678 11684 33694 11701
rect 33106 11668 33694 11684
rect 10142 11646 10730 11662
rect 10142 11629 10158 11646
rect 9696 11612 9898 11629
rect 8938 11574 9898 11612
rect 9956 11612 10158 11629
rect 10714 11629 10730 11646
rect 10714 11612 10916 11629
rect 9956 11574 10916 11612
rect 13762 11194 14350 11210
rect 13762 11177 13778 11194
rect 13576 11160 13778 11177
rect 14334 11177 14350 11194
rect 14780 11194 15368 11210
rect 14780 11177 14796 11194
rect 14334 11160 14536 11177
rect 13576 11122 14536 11160
rect 14594 11160 14796 11177
rect 15352 11177 15368 11194
rect 15798 11194 16386 11210
rect 15798 11177 15814 11194
rect 15352 11160 15554 11177
rect 14594 11122 15554 11160
rect 15612 11160 15814 11177
rect 16370 11177 16386 11194
rect 16816 11194 17404 11210
rect 16816 11177 16832 11194
rect 16370 11160 16572 11177
rect 15612 11122 16572 11160
rect 16630 11160 16832 11177
rect 17388 11177 17404 11194
rect 17834 11194 18422 11210
rect 17834 11177 17850 11194
rect 17388 11160 17590 11177
rect 16630 11122 17590 11160
rect 17648 11160 17850 11177
rect 18406 11177 18422 11194
rect 18852 11194 19440 11210
rect 18852 11177 18868 11194
rect 18406 11160 18608 11177
rect 17648 11122 18608 11160
rect 18666 11160 18868 11177
rect 19424 11177 19440 11194
rect 19870 11194 20458 11210
rect 19870 11177 19886 11194
rect 19424 11160 19626 11177
rect 18666 11122 19626 11160
rect 19684 11160 19886 11177
rect 20442 11177 20458 11194
rect 20888 11194 21476 11210
rect 20888 11177 20904 11194
rect 20442 11160 20644 11177
rect 19684 11122 20644 11160
rect 20702 11160 20904 11177
rect 21460 11177 21476 11194
rect 21906 11194 22494 11210
rect 21906 11177 21922 11194
rect 21460 11160 21662 11177
rect 20702 11122 21662 11160
rect 21720 11160 21922 11177
rect 22478 11177 22494 11194
rect 22924 11194 23512 11210
rect 22924 11177 22940 11194
rect 22478 11160 22680 11177
rect 21720 11122 22680 11160
rect 22738 11160 22940 11177
rect 23496 11177 23512 11194
rect 23942 11194 24530 11210
rect 23942 11177 23958 11194
rect 23496 11160 23698 11177
rect 22738 11122 23698 11160
rect 23756 11160 23958 11177
rect 24514 11177 24530 11194
rect 24960 11194 25548 11210
rect 24960 11177 24976 11194
rect 24514 11160 24716 11177
rect 23756 11122 24716 11160
rect 24774 11160 24976 11177
rect 25532 11177 25548 11194
rect 25978 11194 26566 11210
rect 25978 11177 25994 11194
rect 25532 11160 25734 11177
rect 24774 11122 25734 11160
rect 25792 11160 25994 11177
rect 26550 11177 26566 11194
rect 26996 11194 27584 11210
rect 26996 11177 27012 11194
rect 26550 11160 26752 11177
rect 25792 11122 26752 11160
rect 26810 11160 27012 11177
rect 27568 11177 27584 11194
rect 28014 11194 28602 11210
rect 28014 11177 28030 11194
rect 27568 11160 27770 11177
rect 26810 11122 27770 11160
rect 27828 11160 28030 11177
rect 28586 11177 28602 11194
rect 29032 11194 29620 11210
rect 29032 11177 29048 11194
rect 28586 11160 28788 11177
rect 27828 11122 28788 11160
rect 28846 11160 29048 11177
rect 29604 11177 29620 11194
rect 30050 11194 30638 11210
rect 30050 11177 30066 11194
rect 29604 11160 29806 11177
rect 28846 11122 29806 11160
rect 29864 11160 30066 11177
rect 30622 11177 30638 11194
rect 31068 11194 31656 11210
rect 31068 11177 31084 11194
rect 30622 11160 30824 11177
rect 29864 11122 30824 11160
rect 30882 11160 31084 11177
rect 31640 11177 31656 11194
rect 32086 11194 32674 11210
rect 32086 11177 32102 11194
rect 31640 11160 31842 11177
rect 30882 11122 31842 11160
rect 31900 11160 32102 11177
rect 32658 11177 32674 11194
rect 33104 11194 33692 11210
rect 33104 11177 33120 11194
rect 32658 11160 32860 11177
rect 31900 11122 32860 11160
rect 32918 11160 33120 11177
rect 33676 11177 33692 11194
rect 33676 11160 33878 11177
rect 32918 11122 33878 11160
rect 1812 10936 2772 10974
rect 1812 10919 2014 10936
rect 1998 10902 2014 10919
rect 2570 10919 2772 10936
rect 2830 10936 3790 10974
rect 2830 10919 3032 10936
rect 2570 10902 2586 10919
rect 1998 10886 2586 10902
rect 3016 10902 3032 10919
rect 3588 10919 3790 10936
rect 3848 10936 4808 10974
rect 3848 10919 4050 10936
rect 3588 10902 3604 10919
rect 3016 10886 3604 10902
rect 1998 10828 2586 10844
rect 1998 10811 2014 10828
rect 1812 10794 2014 10811
rect 2570 10811 2586 10828
rect 4034 10902 4050 10919
rect 4606 10919 4808 10936
rect 4866 10936 5826 10974
rect 4866 10919 5068 10936
rect 4606 10902 4622 10919
rect 4034 10886 4622 10902
rect 3016 10828 3604 10844
rect 3016 10811 3032 10828
rect 2570 10794 2772 10811
rect 1812 10756 2772 10794
rect 2830 10794 3032 10811
rect 3588 10811 3604 10828
rect 5052 10902 5068 10919
rect 5624 10919 5826 10936
rect 5884 10936 6844 10974
rect 5884 10919 6086 10936
rect 5624 10902 5640 10919
rect 5052 10886 5640 10902
rect 4034 10828 4622 10844
rect 4034 10811 4050 10828
rect 3588 10794 3790 10811
rect 2830 10756 3790 10794
rect 3848 10794 4050 10811
rect 4606 10811 4622 10828
rect 6070 10902 6086 10919
rect 6642 10919 6844 10936
rect 6902 10936 7862 10974
rect 6902 10919 7104 10936
rect 6642 10902 6658 10919
rect 6070 10886 6658 10902
rect 5052 10828 5640 10844
rect 5052 10811 5068 10828
rect 4606 10794 4808 10811
rect 3848 10756 4808 10794
rect 4866 10794 5068 10811
rect 5624 10811 5640 10828
rect 7088 10902 7104 10919
rect 7660 10919 7862 10936
rect 7920 10936 8880 10974
rect 7920 10919 8122 10936
rect 7660 10902 7676 10919
rect 7088 10886 7676 10902
rect 6070 10828 6658 10844
rect 6070 10811 6086 10828
rect 5624 10794 5826 10811
rect 4866 10756 5826 10794
rect 5884 10794 6086 10811
rect 6642 10811 6658 10828
rect 8106 10902 8122 10919
rect 8678 10919 8880 10936
rect 8938 10936 9898 10974
rect 8938 10919 9140 10936
rect 8678 10902 8694 10919
rect 8106 10886 8694 10902
rect 7088 10828 7676 10844
rect 7088 10811 7104 10828
rect 6642 10794 6844 10811
rect 5884 10756 6844 10794
rect 6902 10794 7104 10811
rect 7660 10811 7676 10828
rect 9124 10902 9140 10919
rect 9696 10919 9898 10936
rect 9956 10936 10916 10974
rect 9956 10919 10158 10936
rect 9696 10902 9712 10919
rect 9124 10886 9712 10902
rect 8106 10828 8694 10844
rect 8106 10811 8122 10828
rect 7660 10794 7862 10811
rect 6902 10756 7862 10794
rect 7920 10794 8122 10811
rect 8678 10811 8694 10828
rect 10142 10902 10158 10919
rect 10714 10919 10916 10936
rect 10714 10902 10730 10919
rect 10142 10886 10730 10902
rect 9124 10828 9712 10844
rect 9124 10811 9140 10828
rect 8678 10794 8880 10811
rect 7920 10756 8880 10794
rect 8938 10794 9140 10811
rect 9696 10811 9712 10828
rect 10142 10828 10730 10844
rect 10142 10811 10158 10828
rect 9696 10794 9898 10811
rect 8938 10756 9898 10794
rect 9956 10794 10158 10811
rect 10714 10811 10730 10828
rect 10714 10794 10916 10811
rect 9956 10756 10916 10794
rect 13576 10484 14536 10522
rect 13576 10467 13778 10484
rect 13762 10450 13778 10467
rect 14334 10467 14536 10484
rect 14594 10484 15554 10522
rect 14594 10467 14796 10484
rect 14334 10450 14350 10467
rect 13762 10434 14350 10450
rect 14780 10450 14796 10467
rect 15352 10467 15554 10484
rect 15612 10484 16572 10522
rect 15612 10467 15814 10484
rect 15352 10450 15368 10467
rect 14780 10434 15368 10450
rect 15798 10450 15814 10467
rect 16370 10467 16572 10484
rect 16630 10484 17590 10522
rect 16630 10467 16832 10484
rect 16370 10450 16386 10467
rect 15798 10434 16386 10450
rect 16816 10450 16832 10467
rect 17388 10467 17590 10484
rect 17648 10484 18608 10522
rect 17648 10467 17850 10484
rect 17388 10450 17404 10467
rect 16816 10434 17404 10450
rect 17834 10450 17850 10467
rect 18406 10467 18608 10484
rect 18666 10484 19626 10522
rect 18666 10467 18868 10484
rect 18406 10450 18422 10467
rect 17834 10434 18422 10450
rect 18852 10450 18868 10467
rect 19424 10467 19626 10484
rect 19684 10484 20644 10522
rect 19684 10467 19886 10484
rect 19424 10450 19440 10467
rect 18852 10434 19440 10450
rect 19870 10450 19886 10467
rect 20442 10467 20644 10484
rect 20702 10484 21662 10522
rect 20702 10467 20904 10484
rect 20442 10450 20458 10467
rect 19870 10434 20458 10450
rect 20888 10450 20904 10467
rect 21460 10467 21662 10484
rect 21720 10484 22680 10522
rect 21720 10467 21922 10484
rect 21460 10450 21476 10467
rect 20888 10434 21476 10450
rect 21906 10450 21922 10467
rect 22478 10467 22680 10484
rect 22738 10484 23698 10522
rect 22738 10467 22940 10484
rect 22478 10450 22494 10467
rect 21906 10434 22494 10450
rect 22924 10450 22940 10467
rect 23496 10467 23698 10484
rect 23756 10484 24716 10522
rect 23756 10467 23958 10484
rect 23496 10450 23512 10467
rect 22924 10434 23512 10450
rect 23942 10450 23958 10467
rect 24514 10467 24716 10484
rect 24774 10484 25734 10522
rect 24774 10467 24976 10484
rect 24514 10450 24530 10467
rect 23942 10434 24530 10450
rect 24960 10450 24976 10467
rect 25532 10467 25734 10484
rect 25792 10484 26752 10522
rect 25792 10467 25994 10484
rect 25532 10450 25548 10467
rect 24960 10434 25548 10450
rect 25978 10450 25994 10467
rect 26550 10467 26752 10484
rect 26810 10484 27770 10522
rect 26810 10467 27012 10484
rect 26550 10450 26566 10467
rect 25978 10434 26566 10450
rect 26996 10450 27012 10467
rect 27568 10467 27770 10484
rect 27828 10484 28788 10522
rect 27828 10467 28030 10484
rect 27568 10450 27584 10467
rect 26996 10434 27584 10450
rect 28014 10450 28030 10467
rect 28586 10467 28788 10484
rect 28846 10484 29806 10522
rect 28846 10467 29048 10484
rect 28586 10450 28602 10467
rect 28014 10434 28602 10450
rect 29032 10450 29048 10467
rect 29604 10467 29806 10484
rect 29864 10484 30824 10522
rect 29864 10467 30066 10484
rect 29604 10450 29620 10467
rect 29032 10434 29620 10450
rect 30050 10450 30066 10467
rect 30622 10467 30824 10484
rect 30882 10484 31842 10522
rect 30882 10467 31084 10484
rect 30622 10450 30638 10467
rect 30050 10434 30638 10450
rect 31068 10450 31084 10467
rect 31640 10467 31842 10484
rect 31900 10484 32860 10522
rect 31900 10467 32102 10484
rect 31640 10450 31656 10467
rect 31068 10434 31656 10450
rect 32086 10450 32102 10467
rect 32658 10467 32860 10484
rect 32918 10484 33878 10522
rect 32918 10467 33120 10484
rect 32658 10450 32674 10467
rect 32086 10434 32674 10450
rect 33104 10450 33120 10467
rect 33676 10467 33878 10484
rect 33676 10450 33692 10467
rect 33104 10434 33692 10450
rect 1812 10118 2772 10156
rect 1812 10101 2014 10118
rect 1998 10084 2014 10101
rect 2570 10101 2772 10118
rect 2830 10118 3790 10156
rect 2830 10101 3032 10118
rect 2570 10084 2586 10101
rect 1998 10068 2586 10084
rect 3016 10084 3032 10101
rect 3588 10101 3790 10118
rect 3848 10118 4808 10156
rect 3848 10101 4050 10118
rect 3588 10084 3604 10101
rect 3016 10068 3604 10084
rect 1998 10010 2586 10026
rect 1998 9993 2014 10010
rect 1812 9976 2014 9993
rect 2570 9993 2586 10010
rect 4034 10084 4050 10101
rect 4606 10101 4808 10118
rect 4866 10118 5826 10156
rect 4866 10101 5068 10118
rect 4606 10084 4622 10101
rect 4034 10068 4622 10084
rect 3016 10010 3604 10026
rect 3016 9993 3032 10010
rect 2570 9976 2772 9993
rect 1812 9938 2772 9976
rect 2830 9976 3032 9993
rect 3588 9993 3604 10010
rect 5052 10084 5068 10101
rect 5624 10101 5826 10118
rect 5884 10118 6844 10156
rect 5884 10101 6086 10118
rect 5624 10084 5640 10101
rect 5052 10068 5640 10084
rect 4034 10010 4622 10026
rect 4034 9993 4050 10010
rect 3588 9976 3790 9993
rect 2830 9938 3790 9976
rect 3848 9976 4050 9993
rect 4606 9993 4622 10010
rect 6070 10084 6086 10101
rect 6642 10101 6844 10118
rect 6902 10118 7862 10156
rect 6902 10101 7104 10118
rect 6642 10084 6658 10101
rect 6070 10068 6658 10084
rect 5052 10010 5640 10026
rect 5052 9993 5068 10010
rect 4606 9976 4808 9993
rect 3848 9938 4808 9976
rect 4866 9976 5068 9993
rect 5624 9993 5640 10010
rect 7088 10084 7104 10101
rect 7660 10101 7862 10118
rect 7920 10118 8880 10156
rect 7920 10101 8122 10118
rect 7660 10084 7676 10101
rect 7088 10068 7676 10084
rect 6070 10010 6658 10026
rect 6070 9993 6086 10010
rect 5624 9976 5826 9993
rect 4866 9938 5826 9976
rect 5884 9976 6086 9993
rect 6642 9993 6658 10010
rect 8106 10084 8122 10101
rect 8678 10101 8880 10118
rect 8938 10118 9898 10156
rect 8938 10101 9140 10118
rect 8678 10084 8694 10101
rect 8106 10068 8694 10084
rect 7088 10010 7676 10026
rect 7088 9993 7104 10010
rect 6642 9976 6844 9993
rect 5884 9938 6844 9976
rect 6902 9976 7104 9993
rect 7660 9993 7676 10010
rect 9124 10084 9140 10101
rect 9696 10101 9898 10118
rect 9956 10118 10916 10156
rect 9956 10101 10158 10118
rect 9696 10084 9712 10101
rect 9124 10068 9712 10084
rect 8106 10010 8694 10026
rect 8106 9993 8122 10010
rect 7660 9976 7862 9993
rect 6902 9938 7862 9976
rect 7920 9976 8122 9993
rect 8678 9993 8694 10010
rect 10142 10084 10158 10101
rect 10714 10101 10916 10118
rect 10714 10084 10730 10101
rect 10142 10068 10730 10084
rect 9124 10010 9712 10026
rect 9124 9993 9140 10010
rect 8678 9976 8880 9993
rect 7920 9938 8880 9976
rect 8938 9976 9140 9993
rect 9696 9993 9712 10010
rect 10142 10010 10730 10026
rect 10142 9993 10158 10010
rect 9696 9976 9898 9993
rect 8938 9938 9898 9976
rect 9956 9976 10158 9993
rect 10714 9993 10730 10010
rect 10714 9976 10916 9993
rect 9956 9938 10916 9976
rect 13762 9960 14350 9976
rect 13762 9943 13778 9960
rect 13576 9926 13778 9943
rect 14334 9943 14350 9960
rect 14780 9960 15368 9976
rect 14780 9943 14796 9960
rect 14334 9926 14536 9943
rect 13576 9888 14536 9926
rect 14594 9926 14796 9943
rect 15352 9943 15368 9960
rect 15798 9960 16386 9976
rect 15798 9943 15814 9960
rect 15352 9926 15554 9943
rect 14594 9888 15554 9926
rect 15612 9926 15814 9943
rect 16370 9943 16386 9960
rect 16816 9960 17404 9976
rect 16816 9943 16832 9960
rect 16370 9926 16572 9943
rect 15612 9888 16572 9926
rect 16630 9926 16832 9943
rect 17388 9943 17404 9960
rect 17834 9960 18422 9976
rect 17834 9943 17850 9960
rect 17388 9926 17590 9943
rect 16630 9888 17590 9926
rect 17648 9926 17850 9943
rect 18406 9943 18422 9960
rect 18852 9960 19440 9976
rect 18852 9943 18868 9960
rect 18406 9926 18608 9943
rect 17648 9888 18608 9926
rect 18666 9926 18868 9943
rect 19424 9943 19440 9960
rect 19870 9960 20458 9976
rect 19870 9943 19886 9960
rect 19424 9926 19626 9943
rect 18666 9888 19626 9926
rect 19684 9926 19886 9943
rect 20442 9943 20458 9960
rect 20888 9960 21476 9976
rect 20888 9943 20904 9960
rect 20442 9926 20644 9943
rect 19684 9888 20644 9926
rect 20702 9926 20904 9943
rect 21460 9943 21476 9960
rect 21906 9960 22494 9976
rect 21906 9943 21922 9960
rect 21460 9926 21662 9943
rect 20702 9888 21662 9926
rect 21720 9926 21922 9943
rect 22478 9943 22494 9960
rect 22924 9960 23512 9976
rect 22924 9943 22940 9960
rect 22478 9926 22680 9943
rect 21720 9888 22680 9926
rect 22738 9926 22940 9943
rect 23496 9943 23512 9960
rect 23942 9960 24530 9976
rect 23942 9943 23958 9960
rect 23496 9926 23698 9943
rect 22738 9888 23698 9926
rect 23756 9926 23958 9943
rect 24514 9943 24530 9960
rect 24960 9960 25548 9976
rect 24960 9943 24976 9960
rect 24514 9926 24716 9943
rect 23756 9888 24716 9926
rect 24774 9926 24976 9943
rect 25532 9943 25548 9960
rect 25978 9960 26566 9976
rect 25978 9943 25994 9960
rect 25532 9926 25734 9943
rect 24774 9888 25734 9926
rect 25792 9926 25994 9943
rect 26550 9943 26566 9960
rect 26996 9960 27584 9976
rect 26996 9943 27012 9960
rect 26550 9926 26752 9943
rect 25792 9888 26752 9926
rect 26810 9926 27012 9943
rect 27568 9943 27584 9960
rect 28014 9960 28602 9976
rect 28014 9943 28030 9960
rect 27568 9926 27770 9943
rect 26810 9888 27770 9926
rect 27828 9926 28030 9943
rect 28586 9943 28602 9960
rect 29032 9960 29620 9976
rect 29032 9943 29048 9960
rect 28586 9926 28788 9943
rect 27828 9888 28788 9926
rect 28846 9926 29048 9943
rect 29604 9943 29620 9960
rect 30050 9960 30638 9976
rect 30050 9943 30066 9960
rect 29604 9926 29806 9943
rect 28846 9888 29806 9926
rect 29864 9926 30066 9943
rect 30622 9943 30638 9960
rect 31068 9960 31656 9976
rect 31068 9943 31084 9960
rect 30622 9926 30824 9943
rect 29864 9888 30824 9926
rect 30882 9926 31084 9943
rect 31640 9943 31656 9960
rect 32086 9960 32674 9976
rect 32086 9943 32102 9960
rect 31640 9926 31842 9943
rect 30882 9888 31842 9926
rect 31900 9926 32102 9943
rect 32658 9943 32674 9960
rect 33104 9960 33692 9976
rect 33104 9943 33120 9960
rect 32658 9926 32860 9943
rect 31900 9888 32860 9926
rect 32918 9926 33120 9943
rect 33676 9943 33692 9960
rect 33676 9926 33878 9943
rect 32918 9888 33878 9926
rect 1812 9300 2772 9338
rect 1812 9283 2014 9300
rect 1998 9266 2014 9283
rect 2570 9283 2772 9300
rect 2830 9300 3790 9338
rect 2830 9283 3032 9300
rect 2570 9266 2586 9283
rect 1998 9250 2586 9266
rect 3016 9266 3032 9283
rect 3588 9283 3790 9300
rect 3848 9300 4808 9338
rect 3848 9283 4050 9300
rect 3588 9266 3604 9283
rect 3016 9250 3604 9266
rect 1998 9192 2586 9208
rect 1998 9175 2014 9192
rect 1812 9158 2014 9175
rect 2570 9175 2586 9192
rect 4034 9266 4050 9283
rect 4606 9283 4808 9300
rect 4866 9300 5826 9338
rect 4866 9283 5068 9300
rect 4606 9266 4622 9283
rect 4034 9250 4622 9266
rect 3016 9192 3604 9208
rect 3016 9175 3032 9192
rect 2570 9158 2772 9175
rect 1812 9120 2772 9158
rect 2830 9158 3032 9175
rect 3588 9175 3604 9192
rect 5052 9266 5068 9283
rect 5624 9283 5826 9300
rect 5884 9300 6844 9338
rect 5884 9283 6086 9300
rect 5624 9266 5640 9283
rect 5052 9250 5640 9266
rect 4034 9192 4622 9208
rect 4034 9175 4050 9192
rect 3588 9158 3790 9175
rect 2830 9120 3790 9158
rect 3848 9158 4050 9175
rect 4606 9175 4622 9192
rect 6070 9266 6086 9283
rect 6642 9283 6844 9300
rect 6902 9300 7862 9338
rect 6902 9283 7104 9300
rect 6642 9266 6658 9283
rect 6070 9250 6658 9266
rect 5052 9192 5640 9208
rect 5052 9175 5068 9192
rect 4606 9158 4808 9175
rect 3848 9120 4808 9158
rect 4866 9158 5068 9175
rect 5624 9175 5640 9192
rect 7088 9266 7104 9283
rect 7660 9283 7862 9300
rect 7920 9300 8880 9338
rect 7920 9283 8122 9300
rect 7660 9266 7676 9283
rect 7088 9250 7676 9266
rect 6070 9192 6658 9208
rect 6070 9175 6086 9192
rect 5624 9158 5826 9175
rect 4866 9120 5826 9158
rect 5884 9158 6086 9175
rect 6642 9175 6658 9192
rect 8106 9266 8122 9283
rect 8678 9283 8880 9300
rect 8938 9300 9898 9338
rect 8938 9283 9140 9300
rect 8678 9266 8694 9283
rect 8106 9250 8694 9266
rect 7088 9192 7676 9208
rect 7088 9175 7104 9192
rect 6642 9158 6844 9175
rect 5884 9120 6844 9158
rect 6902 9158 7104 9175
rect 7660 9175 7676 9192
rect 9124 9266 9140 9283
rect 9696 9283 9898 9300
rect 9956 9300 10916 9338
rect 9956 9283 10158 9300
rect 9696 9266 9712 9283
rect 9124 9250 9712 9266
rect 8106 9192 8694 9208
rect 8106 9175 8122 9192
rect 7660 9158 7862 9175
rect 6902 9120 7862 9158
rect 7920 9158 8122 9175
rect 8678 9175 8694 9192
rect 10142 9266 10158 9283
rect 10714 9283 10916 9300
rect 10714 9266 10730 9283
rect 10142 9250 10730 9266
rect 9124 9192 9712 9208
rect 9124 9175 9140 9192
rect 8678 9158 8880 9175
rect 7920 9120 8880 9158
rect 8938 9158 9140 9175
rect 9696 9175 9712 9192
rect 13576 9250 14536 9288
rect 13576 9233 13778 9250
rect 10142 9192 10730 9208
rect 10142 9175 10158 9192
rect 9696 9158 9898 9175
rect 8938 9120 9898 9158
rect 9956 9158 10158 9175
rect 10714 9175 10730 9192
rect 13762 9216 13778 9233
rect 14334 9233 14536 9250
rect 14594 9250 15554 9288
rect 14594 9233 14796 9250
rect 14334 9216 14350 9233
rect 13762 9200 14350 9216
rect 14780 9216 14796 9233
rect 15352 9233 15554 9250
rect 15612 9250 16572 9288
rect 15612 9233 15814 9250
rect 15352 9216 15368 9233
rect 14780 9200 15368 9216
rect 15798 9216 15814 9233
rect 16370 9233 16572 9250
rect 16630 9250 17590 9288
rect 16630 9233 16832 9250
rect 16370 9216 16386 9233
rect 15798 9200 16386 9216
rect 16816 9216 16832 9233
rect 17388 9233 17590 9250
rect 17648 9250 18608 9288
rect 17648 9233 17850 9250
rect 17388 9216 17404 9233
rect 16816 9200 17404 9216
rect 17834 9216 17850 9233
rect 18406 9233 18608 9250
rect 18666 9250 19626 9288
rect 18666 9233 18868 9250
rect 18406 9216 18422 9233
rect 17834 9200 18422 9216
rect 18852 9216 18868 9233
rect 19424 9233 19626 9250
rect 19684 9250 20644 9288
rect 19684 9233 19886 9250
rect 19424 9216 19440 9233
rect 18852 9200 19440 9216
rect 19870 9216 19886 9233
rect 20442 9233 20644 9250
rect 20702 9250 21662 9288
rect 20702 9233 20904 9250
rect 20442 9216 20458 9233
rect 19870 9200 20458 9216
rect 20888 9216 20904 9233
rect 21460 9233 21662 9250
rect 21720 9250 22680 9288
rect 21720 9233 21922 9250
rect 21460 9216 21476 9233
rect 20888 9200 21476 9216
rect 21906 9216 21922 9233
rect 22478 9233 22680 9250
rect 22738 9250 23698 9288
rect 22738 9233 22940 9250
rect 22478 9216 22494 9233
rect 21906 9200 22494 9216
rect 22924 9216 22940 9233
rect 23496 9233 23698 9250
rect 23756 9250 24716 9288
rect 23756 9233 23958 9250
rect 23496 9216 23512 9233
rect 22924 9200 23512 9216
rect 23942 9216 23958 9233
rect 24514 9233 24716 9250
rect 24774 9250 25734 9288
rect 24774 9233 24976 9250
rect 24514 9216 24530 9233
rect 23942 9200 24530 9216
rect 24960 9216 24976 9233
rect 25532 9233 25734 9250
rect 25792 9250 26752 9288
rect 25792 9233 25994 9250
rect 25532 9216 25548 9233
rect 24960 9200 25548 9216
rect 25978 9216 25994 9233
rect 26550 9233 26752 9250
rect 26810 9250 27770 9288
rect 26810 9233 27012 9250
rect 26550 9216 26566 9233
rect 25978 9200 26566 9216
rect 26996 9216 27012 9233
rect 27568 9233 27770 9250
rect 27828 9250 28788 9288
rect 27828 9233 28030 9250
rect 27568 9216 27584 9233
rect 26996 9200 27584 9216
rect 28014 9216 28030 9233
rect 28586 9233 28788 9250
rect 28846 9250 29806 9288
rect 28846 9233 29048 9250
rect 28586 9216 28602 9233
rect 28014 9200 28602 9216
rect 29032 9216 29048 9233
rect 29604 9233 29806 9250
rect 29864 9250 30824 9288
rect 29864 9233 30066 9250
rect 29604 9216 29620 9233
rect 29032 9200 29620 9216
rect 30050 9216 30066 9233
rect 30622 9233 30824 9250
rect 30882 9250 31842 9288
rect 30882 9233 31084 9250
rect 30622 9216 30638 9233
rect 30050 9200 30638 9216
rect 31068 9216 31084 9233
rect 31640 9233 31842 9250
rect 31900 9250 32860 9288
rect 31900 9233 32102 9250
rect 31640 9216 31656 9233
rect 31068 9200 31656 9216
rect 32086 9216 32102 9233
rect 32658 9233 32860 9250
rect 32918 9250 33878 9288
rect 32918 9233 33120 9250
rect 32658 9216 32674 9233
rect 32086 9200 32674 9216
rect 33104 9216 33120 9233
rect 33676 9233 33878 9250
rect 33676 9216 33692 9233
rect 33104 9200 33692 9216
rect 10714 9158 10916 9175
rect 9956 9120 10916 9158
rect 13762 8728 14350 8744
rect 13762 8711 13778 8728
rect 13576 8694 13778 8711
rect 14334 8711 14350 8728
rect 14780 8728 15368 8744
rect 14780 8711 14796 8728
rect 14334 8694 14536 8711
rect 13576 8656 14536 8694
rect 14594 8694 14796 8711
rect 15352 8711 15368 8728
rect 15798 8728 16386 8744
rect 15798 8711 15814 8728
rect 15352 8694 15554 8711
rect 14594 8656 15554 8694
rect 15612 8694 15814 8711
rect 16370 8711 16386 8728
rect 16816 8728 17404 8744
rect 16816 8711 16832 8728
rect 16370 8694 16572 8711
rect 15612 8656 16572 8694
rect 16630 8694 16832 8711
rect 17388 8711 17404 8728
rect 17834 8728 18422 8744
rect 17834 8711 17850 8728
rect 17388 8694 17590 8711
rect 16630 8656 17590 8694
rect 17648 8694 17850 8711
rect 18406 8711 18422 8728
rect 18852 8728 19440 8744
rect 18852 8711 18868 8728
rect 18406 8694 18608 8711
rect 17648 8656 18608 8694
rect 18666 8694 18868 8711
rect 19424 8711 19440 8728
rect 19870 8728 20458 8744
rect 19870 8711 19886 8728
rect 19424 8694 19626 8711
rect 18666 8656 19626 8694
rect 19684 8694 19886 8711
rect 20442 8711 20458 8728
rect 20888 8728 21476 8744
rect 20888 8711 20904 8728
rect 20442 8694 20644 8711
rect 19684 8656 20644 8694
rect 20702 8694 20904 8711
rect 21460 8711 21476 8728
rect 21906 8728 22494 8744
rect 21906 8711 21922 8728
rect 21460 8694 21662 8711
rect 20702 8656 21662 8694
rect 21720 8694 21922 8711
rect 22478 8711 22494 8728
rect 22924 8728 23512 8744
rect 22924 8711 22940 8728
rect 22478 8694 22680 8711
rect 21720 8656 22680 8694
rect 22738 8694 22940 8711
rect 23496 8711 23512 8728
rect 23942 8728 24530 8744
rect 23942 8711 23958 8728
rect 23496 8694 23698 8711
rect 22738 8656 23698 8694
rect 23756 8694 23958 8711
rect 24514 8711 24530 8728
rect 24960 8728 25548 8744
rect 24960 8711 24976 8728
rect 24514 8694 24716 8711
rect 23756 8656 24716 8694
rect 24774 8694 24976 8711
rect 25532 8711 25548 8728
rect 25978 8728 26566 8744
rect 25978 8711 25994 8728
rect 25532 8694 25734 8711
rect 24774 8656 25734 8694
rect 25792 8694 25994 8711
rect 26550 8711 26566 8728
rect 26996 8728 27584 8744
rect 26996 8711 27012 8728
rect 26550 8694 26752 8711
rect 25792 8656 26752 8694
rect 26810 8694 27012 8711
rect 27568 8711 27584 8728
rect 28014 8728 28602 8744
rect 28014 8711 28030 8728
rect 27568 8694 27770 8711
rect 26810 8656 27770 8694
rect 27828 8694 28030 8711
rect 28586 8711 28602 8728
rect 29032 8728 29620 8744
rect 29032 8711 29048 8728
rect 28586 8694 28788 8711
rect 27828 8656 28788 8694
rect 28846 8694 29048 8711
rect 29604 8711 29620 8728
rect 30050 8728 30638 8744
rect 30050 8711 30066 8728
rect 29604 8694 29806 8711
rect 28846 8656 29806 8694
rect 29864 8694 30066 8711
rect 30622 8711 30638 8728
rect 31068 8728 31656 8744
rect 31068 8711 31084 8728
rect 30622 8694 30824 8711
rect 29864 8656 30824 8694
rect 30882 8694 31084 8711
rect 31640 8711 31656 8728
rect 32086 8728 32674 8744
rect 32086 8711 32102 8728
rect 31640 8694 31842 8711
rect 30882 8656 31842 8694
rect 31900 8694 32102 8711
rect 32658 8711 32674 8728
rect 33104 8728 33692 8744
rect 33104 8711 33120 8728
rect 32658 8694 32860 8711
rect 31900 8656 32860 8694
rect 32918 8694 33120 8711
rect 33676 8711 33692 8728
rect 33676 8694 33878 8711
rect 32918 8656 33878 8694
rect 1812 8482 2772 8520
rect 1812 8465 2014 8482
rect 1998 8448 2014 8465
rect 2570 8465 2772 8482
rect 2830 8482 3790 8520
rect 2830 8465 3032 8482
rect 2570 8448 2586 8465
rect 1998 8432 2586 8448
rect 3016 8448 3032 8465
rect 3588 8465 3790 8482
rect 3848 8482 4808 8520
rect 3848 8465 4050 8482
rect 3588 8448 3604 8465
rect 3016 8432 3604 8448
rect 1998 8374 2586 8390
rect 1998 8357 2014 8374
rect 1812 8340 2014 8357
rect 2570 8357 2586 8374
rect 4034 8448 4050 8465
rect 4606 8465 4808 8482
rect 4866 8482 5826 8520
rect 4866 8465 5068 8482
rect 4606 8448 4622 8465
rect 4034 8432 4622 8448
rect 3016 8374 3604 8390
rect 3016 8357 3032 8374
rect 2570 8340 2772 8357
rect 1812 8302 2772 8340
rect 2830 8340 3032 8357
rect 3588 8357 3604 8374
rect 5052 8448 5068 8465
rect 5624 8465 5826 8482
rect 5884 8482 6844 8520
rect 5884 8465 6086 8482
rect 5624 8448 5640 8465
rect 5052 8432 5640 8448
rect 4034 8374 4622 8390
rect 4034 8357 4050 8374
rect 3588 8340 3790 8357
rect 2830 8302 3790 8340
rect 3848 8340 4050 8357
rect 4606 8357 4622 8374
rect 6070 8448 6086 8465
rect 6642 8465 6844 8482
rect 6902 8482 7862 8520
rect 6902 8465 7104 8482
rect 6642 8448 6658 8465
rect 6070 8432 6658 8448
rect 5052 8374 5640 8390
rect 5052 8357 5068 8374
rect 4606 8340 4808 8357
rect 3848 8302 4808 8340
rect 4866 8340 5068 8357
rect 5624 8357 5640 8374
rect 7088 8448 7104 8465
rect 7660 8465 7862 8482
rect 7920 8482 8880 8520
rect 7920 8465 8122 8482
rect 7660 8448 7676 8465
rect 7088 8432 7676 8448
rect 6070 8374 6658 8390
rect 6070 8357 6086 8374
rect 5624 8340 5826 8357
rect 4866 8302 5826 8340
rect 5884 8340 6086 8357
rect 6642 8357 6658 8374
rect 8106 8448 8122 8465
rect 8678 8465 8880 8482
rect 8938 8482 9898 8520
rect 8938 8465 9140 8482
rect 8678 8448 8694 8465
rect 8106 8432 8694 8448
rect 7088 8374 7676 8390
rect 7088 8357 7104 8374
rect 6642 8340 6844 8357
rect 5884 8302 6844 8340
rect 6902 8340 7104 8357
rect 7660 8357 7676 8374
rect 9124 8448 9140 8465
rect 9696 8465 9898 8482
rect 9956 8482 10916 8520
rect 9956 8465 10158 8482
rect 9696 8448 9712 8465
rect 9124 8432 9712 8448
rect 8106 8374 8694 8390
rect 8106 8357 8122 8374
rect 7660 8340 7862 8357
rect 6902 8302 7862 8340
rect 7920 8340 8122 8357
rect 8678 8357 8694 8374
rect 10142 8448 10158 8465
rect 10714 8465 10916 8482
rect 10714 8448 10730 8465
rect 10142 8432 10730 8448
rect 9124 8374 9712 8390
rect 9124 8357 9140 8374
rect 8678 8340 8880 8357
rect 7920 8302 8880 8340
rect 8938 8340 9140 8357
rect 9696 8357 9712 8374
rect 10142 8374 10730 8390
rect 10142 8357 10158 8374
rect 9696 8340 9898 8357
rect 8938 8302 9898 8340
rect 9956 8340 10158 8357
rect 10714 8357 10730 8374
rect 10714 8340 10916 8357
rect 9956 8302 10916 8340
rect 13576 8018 14536 8056
rect 13576 8001 13778 8018
rect 13762 7984 13778 8001
rect 14334 8001 14536 8018
rect 14594 8018 15554 8056
rect 14594 8001 14796 8018
rect 14334 7984 14350 8001
rect 13762 7968 14350 7984
rect 14780 7984 14796 8001
rect 15352 8001 15554 8018
rect 15612 8018 16572 8056
rect 15612 8001 15814 8018
rect 15352 7984 15368 8001
rect 14780 7968 15368 7984
rect 15798 7984 15814 8001
rect 16370 8001 16572 8018
rect 16630 8018 17590 8056
rect 16630 8001 16832 8018
rect 16370 7984 16386 8001
rect 15798 7968 16386 7984
rect 16816 7984 16832 8001
rect 17388 8001 17590 8018
rect 17648 8018 18608 8056
rect 17648 8001 17850 8018
rect 17388 7984 17404 8001
rect 16816 7968 17404 7984
rect 17834 7984 17850 8001
rect 18406 8001 18608 8018
rect 18666 8018 19626 8056
rect 18666 8001 18868 8018
rect 18406 7984 18422 8001
rect 17834 7968 18422 7984
rect 18852 7984 18868 8001
rect 19424 8001 19626 8018
rect 19684 8018 20644 8056
rect 19684 8001 19886 8018
rect 19424 7984 19440 8001
rect 18852 7968 19440 7984
rect 19870 7984 19886 8001
rect 20442 8001 20644 8018
rect 20702 8018 21662 8056
rect 20702 8001 20904 8018
rect 20442 7984 20458 8001
rect 19870 7968 20458 7984
rect 20888 7984 20904 8001
rect 21460 8001 21662 8018
rect 21720 8018 22680 8056
rect 21720 8001 21922 8018
rect 21460 7984 21476 8001
rect 20888 7968 21476 7984
rect 21906 7984 21922 8001
rect 22478 8001 22680 8018
rect 22738 8018 23698 8056
rect 22738 8001 22940 8018
rect 22478 7984 22494 8001
rect 21906 7968 22494 7984
rect 22924 7984 22940 8001
rect 23496 8001 23698 8018
rect 23756 8018 24716 8056
rect 23756 8001 23958 8018
rect 23496 7984 23512 8001
rect 22924 7968 23512 7984
rect 23942 7984 23958 8001
rect 24514 8001 24716 8018
rect 24774 8018 25734 8056
rect 24774 8001 24976 8018
rect 24514 7984 24530 8001
rect 23942 7968 24530 7984
rect 24960 7984 24976 8001
rect 25532 8001 25734 8018
rect 25792 8018 26752 8056
rect 25792 8001 25994 8018
rect 25532 7984 25548 8001
rect 24960 7968 25548 7984
rect 25978 7984 25994 8001
rect 26550 8001 26752 8018
rect 26810 8018 27770 8056
rect 26810 8001 27012 8018
rect 26550 7984 26566 8001
rect 25978 7968 26566 7984
rect 26996 7984 27012 8001
rect 27568 8001 27770 8018
rect 27828 8018 28788 8056
rect 27828 8001 28030 8018
rect 27568 7984 27584 8001
rect 26996 7968 27584 7984
rect 28014 7984 28030 8001
rect 28586 8001 28788 8018
rect 28846 8018 29806 8056
rect 28846 8001 29048 8018
rect 28586 7984 28602 8001
rect 28014 7968 28602 7984
rect 29032 7984 29048 8001
rect 29604 8001 29806 8018
rect 29864 8018 30824 8056
rect 29864 8001 30066 8018
rect 29604 7984 29620 8001
rect 29032 7968 29620 7984
rect 30050 7984 30066 8001
rect 30622 8001 30824 8018
rect 30882 8018 31842 8056
rect 30882 8001 31084 8018
rect 30622 7984 30638 8001
rect 30050 7968 30638 7984
rect 31068 7984 31084 8001
rect 31640 8001 31842 8018
rect 31900 8018 32860 8056
rect 31900 8001 32102 8018
rect 31640 7984 31656 8001
rect 31068 7968 31656 7984
rect 32086 7984 32102 8001
rect 32658 8001 32860 8018
rect 32918 8018 33878 8056
rect 32918 8001 33120 8018
rect 32658 7984 32674 8001
rect 32086 7968 32674 7984
rect 33104 7984 33120 8001
rect 33676 8001 33878 8018
rect 33676 7984 33692 8001
rect 33104 7968 33692 7984
rect 1812 7664 2772 7702
rect 1812 7647 2014 7664
rect 1998 7630 2014 7647
rect 2570 7647 2772 7664
rect 2830 7664 3790 7702
rect 2830 7647 3032 7664
rect 2570 7630 2586 7647
rect 1998 7614 2586 7630
rect 3016 7630 3032 7647
rect 3588 7647 3790 7664
rect 3848 7664 4808 7702
rect 3848 7647 4050 7664
rect 3588 7630 3604 7647
rect 3016 7614 3604 7630
rect 4034 7630 4050 7647
rect 4606 7647 4808 7664
rect 4866 7664 5826 7702
rect 4866 7647 5068 7664
rect 4606 7630 4622 7647
rect 4034 7614 4622 7630
rect 5052 7630 5068 7647
rect 5624 7647 5826 7664
rect 5884 7664 6844 7702
rect 5884 7647 6086 7664
rect 5624 7630 5640 7647
rect 5052 7614 5640 7630
rect 6070 7630 6086 7647
rect 6642 7647 6844 7664
rect 6902 7664 7862 7702
rect 6902 7647 7104 7664
rect 6642 7630 6658 7647
rect 6070 7614 6658 7630
rect 7088 7630 7104 7647
rect 7660 7647 7862 7664
rect 7920 7664 8880 7702
rect 7920 7647 8122 7664
rect 7660 7630 7676 7647
rect 7088 7614 7676 7630
rect 8106 7630 8122 7647
rect 8678 7647 8880 7664
rect 8938 7664 9898 7702
rect 8938 7647 9140 7664
rect 8678 7630 8694 7647
rect 8106 7614 8694 7630
rect 9124 7630 9140 7647
rect 9696 7647 9898 7664
rect 9956 7664 10916 7702
rect 9956 7647 10158 7664
rect 9696 7630 9712 7647
rect 9124 7614 9712 7630
rect 10142 7630 10158 7647
rect 10714 7647 10916 7664
rect 10714 7630 10730 7647
rect 10142 7614 10730 7630
rect 13762 7494 14350 7510
rect 13762 7477 13778 7494
rect 13576 7460 13778 7477
rect 14334 7477 14350 7494
rect 14780 7494 15368 7510
rect 14780 7477 14796 7494
rect 14334 7460 14536 7477
rect 13576 7422 14536 7460
rect 14594 7460 14796 7477
rect 15352 7477 15368 7494
rect 15798 7494 16386 7510
rect 15798 7477 15814 7494
rect 15352 7460 15554 7477
rect 14594 7422 15554 7460
rect 15612 7460 15814 7477
rect 16370 7477 16386 7494
rect 16816 7494 17404 7510
rect 16816 7477 16832 7494
rect 16370 7460 16572 7477
rect 15612 7422 16572 7460
rect 16630 7460 16832 7477
rect 17388 7477 17404 7494
rect 17834 7494 18422 7510
rect 17834 7477 17850 7494
rect 17388 7460 17590 7477
rect 16630 7422 17590 7460
rect 17648 7460 17850 7477
rect 18406 7477 18422 7494
rect 18852 7494 19440 7510
rect 18852 7477 18868 7494
rect 18406 7460 18608 7477
rect 17648 7422 18608 7460
rect 18666 7460 18868 7477
rect 19424 7477 19440 7494
rect 19870 7494 20458 7510
rect 19870 7477 19886 7494
rect 19424 7460 19626 7477
rect 18666 7422 19626 7460
rect 19684 7460 19886 7477
rect 20442 7477 20458 7494
rect 20888 7494 21476 7510
rect 20888 7477 20904 7494
rect 20442 7460 20644 7477
rect 19684 7422 20644 7460
rect 20702 7460 20904 7477
rect 21460 7477 21476 7494
rect 21906 7494 22494 7510
rect 21906 7477 21922 7494
rect 21460 7460 21662 7477
rect 20702 7422 21662 7460
rect 21720 7460 21922 7477
rect 22478 7477 22494 7494
rect 22924 7494 23512 7510
rect 22924 7477 22940 7494
rect 22478 7460 22680 7477
rect 21720 7422 22680 7460
rect 22738 7460 22940 7477
rect 23496 7477 23512 7494
rect 23942 7494 24530 7510
rect 23942 7477 23958 7494
rect 23496 7460 23698 7477
rect 22738 7422 23698 7460
rect 23756 7460 23958 7477
rect 24514 7477 24530 7494
rect 24960 7494 25548 7510
rect 24960 7477 24976 7494
rect 24514 7460 24716 7477
rect 23756 7422 24716 7460
rect 24774 7460 24976 7477
rect 25532 7477 25548 7494
rect 25978 7494 26566 7510
rect 25978 7477 25994 7494
rect 25532 7460 25734 7477
rect 24774 7422 25734 7460
rect 25792 7460 25994 7477
rect 26550 7477 26566 7494
rect 26996 7494 27584 7510
rect 26996 7477 27012 7494
rect 26550 7460 26752 7477
rect 25792 7422 26752 7460
rect 26810 7460 27012 7477
rect 27568 7477 27584 7494
rect 28014 7494 28602 7510
rect 28014 7477 28030 7494
rect 27568 7460 27770 7477
rect 26810 7422 27770 7460
rect 27828 7460 28030 7477
rect 28586 7477 28602 7494
rect 29032 7494 29620 7510
rect 29032 7477 29048 7494
rect 28586 7460 28788 7477
rect 27828 7422 28788 7460
rect 28846 7460 29048 7477
rect 29604 7477 29620 7494
rect 30050 7494 30638 7510
rect 30050 7477 30066 7494
rect 29604 7460 29806 7477
rect 28846 7422 29806 7460
rect 29864 7460 30066 7477
rect 30622 7477 30638 7494
rect 31068 7494 31656 7510
rect 31068 7477 31084 7494
rect 30622 7460 30824 7477
rect 29864 7422 30824 7460
rect 30882 7460 31084 7477
rect 31640 7477 31656 7494
rect 32086 7494 32674 7510
rect 32086 7477 32102 7494
rect 31640 7460 31842 7477
rect 30882 7422 31842 7460
rect 31900 7460 32102 7477
rect 32658 7477 32674 7494
rect 33104 7494 33692 7510
rect 33104 7477 33120 7494
rect 32658 7460 32860 7477
rect 31900 7422 32860 7460
rect 32918 7460 33120 7477
rect 33676 7477 33692 7494
rect 33676 7460 33878 7477
rect 32918 7422 33878 7460
rect 8698 6990 8806 7006
rect 8698 6973 8714 6990
rect 8672 6956 8714 6973
rect 8790 6973 8806 6990
rect 8916 6990 9024 7006
rect 8916 6973 8932 6990
rect 8790 6956 8832 6973
rect 8672 6918 8832 6956
rect 8890 6956 8932 6973
rect 9008 6973 9024 6990
rect 9134 6990 9242 7006
rect 9134 6973 9150 6990
rect 9008 6956 9050 6973
rect 8890 6918 9050 6956
rect 9108 6956 9150 6973
rect 9226 6973 9242 6990
rect 9352 6990 9460 7006
rect 9352 6973 9368 6990
rect 9226 6956 9268 6973
rect 9108 6918 9268 6956
rect 9326 6956 9368 6973
rect 9444 6973 9460 6990
rect 9570 6990 9678 7006
rect 9570 6973 9586 6990
rect 9444 6956 9486 6973
rect 9326 6918 9486 6956
rect 9544 6956 9586 6973
rect 9662 6973 9678 6990
rect 9788 6990 9896 7006
rect 9788 6973 9804 6990
rect 9662 6956 9704 6973
rect 9544 6918 9704 6956
rect 9762 6956 9804 6973
rect 9880 6973 9896 6990
rect 10006 6990 10114 7006
rect 10006 6973 10022 6990
rect 9880 6956 9922 6973
rect 9762 6918 9922 6956
rect 9980 6956 10022 6973
rect 10098 6973 10114 6990
rect 10224 6990 10332 7006
rect 10224 6973 10240 6990
rect 10098 6956 10140 6973
rect 9980 6918 10140 6956
rect 10198 6956 10240 6973
rect 10316 6973 10332 6990
rect 10442 6990 10550 7006
rect 10442 6973 10458 6990
rect 10316 6956 10358 6973
rect 10198 6918 10358 6956
rect 10416 6956 10458 6973
rect 10534 6973 10550 6990
rect 10660 6990 10768 7006
rect 10660 6973 10676 6990
rect 10534 6956 10576 6973
rect 10416 6918 10576 6956
rect 10634 6956 10676 6973
rect 10752 6973 10768 6990
rect 10752 6956 10794 6973
rect 10634 6918 10794 6956
rect 13576 6784 14536 6822
rect 13576 6767 13778 6784
rect 13762 6750 13778 6767
rect 14334 6767 14536 6784
rect 14594 6784 15554 6822
rect 14594 6767 14796 6784
rect 14334 6750 14350 6767
rect 13762 6734 14350 6750
rect 14780 6750 14796 6767
rect 15352 6767 15554 6784
rect 15612 6784 16572 6822
rect 15612 6767 15814 6784
rect 15352 6750 15368 6767
rect 14780 6734 15368 6750
rect 15798 6750 15814 6767
rect 16370 6767 16572 6784
rect 16630 6784 17590 6822
rect 16630 6767 16832 6784
rect 16370 6750 16386 6767
rect 15798 6734 16386 6750
rect 16816 6750 16832 6767
rect 17388 6767 17590 6784
rect 17648 6784 18608 6822
rect 17648 6767 17850 6784
rect 17388 6750 17404 6767
rect 16816 6734 17404 6750
rect 17834 6750 17850 6767
rect 18406 6767 18608 6784
rect 18666 6784 19626 6822
rect 18666 6767 18868 6784
rect 18406 6750 18422 6767
rect 17834 6734 18422 6750
rect 18852 6750 18868 6767
rect 19424 6767 19626 6784
rect 19684 6784 20644 6822
rect 19684 6767 19886 6784
rect 19424 6750 19440 6767
rect 18852 6734 19440 6750
rect 19870 6750 19886 6767
rect 20442 6767 20644 6784
rect 20702 6784 21662 6822
rect 20702 6767 20904 6784
rect 20442 6750 20458 6767
rect 19870 6734 20458 6750
rect 20888 6750 20904 6767
rect 21460 6767 21662 6784
rect 21720 6784 22680 6822
rect 21720 6767 21922 6784
rect 21460 6750 21476 6767
rect 20888 6734 21476 6750
rect 21906 6750 21922 6767
rect 22478 6767 22680 6784
rect 22738 6784 23698 6822
rect 22738 6767 22940 6784
rect 22478 6750 22494 6767
rect 21906 6734 22494 6750
rect 22924 6750 22940 6767
rect 23496 6767 23698 6784
rect 23756 6784 24716 6822
rect 23756 6767 23958 6784
rect 23496 6750 23512 6767
rect 22924 6734 23512 6750
rect 23942 6750 23958 6767
rect 24514 6767 24716 6784
rect 24774 6784 25734 6822
rect 24774 6767 24976 6784
rect 24514 6750 24530 6767
rect 23942 6734 24530 6750
rect 24960 6750 24976 6767
rect 25532 6767 25734 6784
rect 25792 6784 26752 6822
rect 25792 6767 25994 6784
rect 25532 6750 25548 6767
rect 24960 6734 25548 6750
rect 25978 6750 25994 6767
rect 26550 6767 26752 6784
rect 26810 6784 27770 6822
rect 26810 6767 27012 6784
rect 26550 6750 26566 6767
rect 25978 6734 26566 6750
rect 26996 6750 27012 6767
rect 27568 6767 27770 6784
rect 27828 6784 28788 6822
rect 27828 6767 28030 6784
rect 27568 6750 27584 6767
rect 26996 6734 27584 6750
rect 28014 6750 28030 6767
rect 28586 6767 28788 6784
rect 28846 6784 29806 6822
rect 28846 6767 29048 6784
rect 28586 6750 28602 6767
rect 28014 6734 28602 6750
rect 29032 6750 29048 6767
rect 29604 6767 29806 6784
rect 29864 6784 30824 6822
rect 29864 6767 30066 6784
rect 29604 6750 29620 6767
rect 29032 6734 29620 6750
rect 30050 6750 30066 6767
rect 30622 6767 30824 6784
rect 30882 6784 31842 6822
rect 30882 6767 31084 6784
rect 30622 6750 30638 6767
rect 30050 6734 30638 6750
rect 31068 6750 31084 6767
rect 31640 6767 31842 6784
rect 31900 6784 32860 6822
rect 31900 6767 32102 6784
rect 31640 6750 31656 6767
rect 31068 6734 31656 6750
rect 32086 6750 32102 6767
rect 32658 6767 32860 6784
rect 32918 6784 33878 6822
rect 32918 6767 33120 6784
rect 32658 6750 32674 6767
rect 32086 6734 32674 6750
rect 33104 6750 33120 6767
rect 33676 6767 33878 6784
rect 33676 6750 33692 6767
rect 33104 6734 33692 6750
rect 8672 6680 8832 6718
rect 8672 6663 8714 6680
rect 8698 6646 8714 6663
rect 8790 6663 8832 6680
rect 8890 6680 9050 6718
rect 8890 6663 8932 6680
rect 8790 6646 8806 6663
rect 8698 6630 8806 6646
rect 8916 6646 8932 6663
rect 9008 6663 9050 6680
rect 9108 6680 9268 6718
rect 9108 6663 9150 6680
rect 9008 6646 9024 6663
rect 8916 6630 9024 6646
rect 9134 6646 9150 6663
rect 9226 6663 9268 6680
rect 9326 6680 9486 6718
rect 9326 6663 9368 6680
rect 9226 6646 9242 6663
rect 9134 6630 9242 6646
rect 9352 6646 9368 6663
rect 9444 6663 9486 6680
rect 9544 6680 9704 6718
rect 9544 6663 9586 6680
rect 9444 6646 9460 6663
rect 9352 6630 9460 6646
rect 9570 6646 9586 6663
rect 9662 6663 9704 6680
rect 9762 6680 9922 6718
rect 9762 6663 9804 6680
rect 9662 6646 9678 6663
rect 9570 6630 9678 6646
rect 9788 6646 9804 6663
rect 9880 6663 9922 6680
rect 9980 6680 10140 6718
rect 9980 6663 10022 6680
rect 9880 6646 9896 6663
rect 9788 6630 9896 6646
rect 10006 6646 10022 6663
rect 10098 6663 10140 6680
rect 10198 6680 10358 6718
rect 10198 6663 10240 6680
rect 10098 6646 10114 6663
rect 10006 6630 10114 6646
rect 10224 6646 10240 6663
rect 10316 6663 10358 6680
rect 10416 6680 10576 6718
rect 10416 6663 10458 6680
rect 10316 6646 10332 6663
rect 10224 6630 10332 6646
rect 10442 6646 10458 6663
rect 10534 6663 10576 6680
rect 10634 6680 10794 6718
rect 10634 6663 10676 6680
rect 10534 6646 10550 6663
rect 10442 6630 10550 6646
rect 10660 6646 10676 6663
rect 10752 6663 10794 6680
rect 10752 6646 10768 6663
rect 10660 6630 10768 6646
rect 13762 6260 14350 6276
rect 13762 6243 13778 6260
rect 13576 6226 13778 6243
rect 14334 6243 14350 6260
rect 14780 6260 15368 6276
rect 14780 6243 14796 6260
rect 14334 6226 14536 6243
rect 13576 6188 14536 6226
rect 14594 6226 14796 6243
rect 15352 6243 15368 6260
rect 15798 6260 16386 6276
rect 15798 6243 15814 6260
rect 15352 6226 15554 6243
rect 14594 6188 15554 6226
rect 15612 6226 15814 6243
rect 16370 6243 16386 6260
rect 16816 6260 17404 6276
rect 16816 6243 16832 6260
rect 16370 6226 16572 6243
rect 15612 6188 16572 6226
rect 16630 6226 16832 6243
rect 17388 6243 17404 6260
rect 17834 6260 18422 6276
rect 17834 6243 17850 6260
rect 17388 6226 17590 6243
rect 16630 6188 17590 6226
rect 17648 6226 17850 6243
rect 18406 6243 18422 6260
rect 18852 6260 19440 6276
rect 18852 6243 18868 6260
rect 18406 6226 18608 6243
rect 17648 6188 18608 6226
rect 18666 6226 18868 6243
rect 19424 6243 19440 6260
rect 19870 6260 20458 6276
rect 19870 6243 19886 6260
rect 19424 6226 19626 6243
rect 18666 6188 19626 6226
rect 19684 6226 19886 6243
rect 20442 6243 20458 6260
rect 20888 6260 21476 6276
rect 20888 6243 20904 6260
rect 20442 6226 20644 6243
rect 19684 6188 20644 6226
rect 20702 6226 20904 6243
rect 21460 6243 21476 6260
rect 21906 6260 22494 6276
rect 21906 6243 21922 6260
rect 21460 6226 21662 6243
rect 20702 6188 21662 6226
rect 21720 6226 21922 6243
rect 22478 6243 22494 6260
rect 22924 6260 23512 6276
rect 22924 6243 22940 6260
rect 22478 6226 22680 6243
rect 21720 6188 22680 6226
rect 22738 6226 22940 6243
rect 23496 6243 23512 6260
rect 23942 6260 24530 6276
rect 23942 6243 23958 6260
rect 23496 6226 23698 6243
rect 22738 6188 23698 6226
rect 23756 6226 23958 6243
rect 24514 6243 24530 6260
rect 24960 6260 25548 6276
rect 24960 6243 24976 6260
rect 24514 6226 24716 6243
rect 23756 6188 24716 6226
rect 24774 6226 24976 6243
rect 25532 6243 25548 6260
rect 25978 6260 26566 6276
rect 25978 6243 25994 6260
rect 25532 6226 25734 6243
rect 24774 6188 25734 6226
rect 25792 6226 25994 6243
rect 26550 6243 26566 6260
rect 26996 6260 27584 6276
rect 26996 6243 27012 6260
rect 26550 6226 26752 6243
rect 25792 6188 26752 6226
rect 26810 6226 27012 6243
rect 27568 6243 27584 6260
rect 28014 6260 28602 6276
rect 28014 6243 28030 6260
rect 27568 6226 27770 6243
rect 26810 6188 27770 6226
rect 27828 6226 28030 6243
rect 28586 6243 28602 6260
rect 29032 6260 29620 6276
rect 29032 6243 29048 6260
rect 28586 6226 28788 6243
rect 27828 6188 28788 6226
rect 28846 6226 29048 6243
rect 29604 6243 29620 6260
rect 30050 6260 30638 6276
rect 30050 6243 30066 6260
rect 29604 6226 29806 6243
rect 28846 6188 29806 6226
rect 29864 6226 30066 6243
rect 30622 6243 30638 6260
rect 31068 6260 31656 6276
rect 31068 6243 31084 6260
rect 30622 6226 30824 6243
rect 29864 6188 30824 6226
rect 30882 6226 31084 6243
rect 31640 6243 31656 6260
rect 32086 6260 32674 6276
rect 32086 6243 32102 6260
rect 31640 6226 31842 6243
rect 30882 6188 31842 6226
rect 31900 6226 32102 6243
rect 32658 6243 32674 6260
rect 33104 6260 33692 6276
rect 33104 6243 33120 6260
rect 32658 6226 32860 6243
rect 31900 6188 32860 6226
rect 32918 6226 33120 6243
rect 33676 6243 33692 6260
rect 33676 6226 33878 6243
rect 32918 6188 33878 6226
rect 8698 6158 8806 6174
rect 8698 6141 8714 6158
rect 8672 6124 8714 6141
rect 8790 6141 8806 6158
rect 8916 6158 9024 6174
rect 8916 6141 8932 6158
rect 8790 6124 8832 6141
rect 8672 6086 8832 6124
rect 8890 6124 8932 6141
rect 9008 6141 9024 6158
rect 9134 6158 9242 6174
rect 9134 6141 9150 6158
rect 9008 6124 9050 6141
rect 8890 6086 9050 6124
rect 9108 6124 9150 6141
rect 9226 6141 9242 6158
rect 9352 6158 9460 6174
rect 9352 6141 9368 6158
rect 9226 6124 9268 6141
rect 9108 6086 9268 6124
rect 9326 6124 9368 6141
rect 9444 6141 9460 6158
rect 9570 6158 9678 6174
rect 9570 6141 9586 6158
rect 9444 6124 9486 6141
rect 9326 6086 9486 6124
rect 9544 6124 9586 6141
rect 9662 6141 9678 6158
rect 9788 6158 9896 6174
rect 9788 6141 9804 6158
rect 9662 6124 9704 6141
rect 9544 6086 9704 6124
rect 9762 6124 9804 6141
rect 9880 6141 9896 6158
rect 10006 6158 10114 6174
rect 10006 6141 10022 6158
rect 9880 6124 9922 6141
rect 9762 6086 9922 6124
rect 9980 6124 10022 6141
rect 10098 6141 10114 6158
rect 10224 6158 10332 6174
rect 10224 6141 10240 6158
rect 10098 6124 10140 6141
rect 9980 6086 10140 6124
rect 10198 6124 10240 6141
rect 10316 6141 10332 6158
rect 10442 6158 10550 6174
rect 10442 6141 10458 6158
rect 10316 6124 10358 6141
rect 10198 6086 10358 6124
rect 10416 6124 10458 6141
rect 10534 6141 10550 6158
rect 10660 6158 10768 6174
rect 10660 6141 10676 6158
rect 10534 6124 10576 6141
rect 10416 6086 10576 6124
rect 10634 6124 10676 6141
rect 10752 6141 10768 6158
rect 10752 6124 10794 6141
rect 10634 6086 10794 6124
rect 8672 5848 8832 5886
rect 8672 5831 8714 5848
rect 8698 5814 8714 5831
rect 8790 5831 8832 5848
rect 8890 5848 9050 5886
rect 8890 5831 8932 5848
rect 8790 5814 8806 5831
rect 8698 5798 8806 5814
rect 8916 5814 8932 5831
rect 9008 5831 9050 5848
rect 9108 5848 9268 5886
rect 9108 5831 9150 5848
rect 9008 5814 9024 5831
rect 8916 5798 9024 5814
rect 9134 5814 9150 5831
rect 9226 5831 9268 5848
rect 9326 5848 9486 5886
rect 9326 5831 9368 5848
rect 9226 5814 9242 5831
rect 9134 5798 9242 5814
rect 9352 5814 9368 5831
rect 9444 5831 9486 5848
rect 9544 5848 9704 5886
rect 9544 5831 9586 5848
rect 9444 5814 9460 5831
rect 9352 5798 9460 5814
rect 9570 5814 9586 5831
rect 9662 5831 9704 5848
rect 9762 5848 9922 5886
rect 9762 5831 9804 5848
rect 9662 5814 9678 5831
rect 9570 5798 9678 5814
rect 9788 5814 9804 5831
rect 9880 5831 9922 5848
rect 9980 5848 10140 5886
rect 9980 5831 10022 5848
rect 9880 5814 9896 5831
rect 9788 5798 9896 5814
rect 10006 5814 10022 5831
rect 10098 5831 10140 5848
rect 10198 5848 10358 5886
rect 10198 5831 10240 5848
rect 10098 5814 10114 5831
rect 10006 5798 10114 5814
rect 10224 5814 10240 5831
rect 10316 5831 10358 5848
rect 10416 5848 10576 5886
rect 10416 5831 10458 5848
rect 10316 5814 10332 5831
rect 10224 5798 10332 5814
rect 10442 5814 10458 5831
rect 10534 5831 10576 5848
rect 10634 5848 10794 5886
rect 10634 5831 10676 5848
rect 10534 5814 10550 5831
rect 10442 5798 10550 5814
rect 10660 5814 10676 5831
rect 10752 5831 10794 5848
rect 10752 5814 10768 5831
rect 10660 5798 10768 5814
rect 13576 5550 14536 5588
rect 13576 5533 13778 5550
rect 13762 5516 13778 5533
rect 14334 5533 14536 5550
rect 14594 5550 15554 5588
rect 14594 5533 14796 5550
rect 14334 5516 14350 5533
rect 13762 5500 14350 5516
rect 14780 5516 14796 5533
rect 15352 5533 15554 5550
rect 15612 5550 16572 5588
rect 15612 5533 15814 5550
rect 15352 5516 15368 5533
rect 14780 5500 15368 5516
rect 15798 5516 15814 5533
rect 16370 5533 16572 5550
rect 16630 5550 17590 5588
rect 16630 5533 16832 5550
rect 16370 5516 16386 5533
rect 15798 5500 16386 5516
rect 16816 5516 16832 5533
rect 17388 5533 17590 5550
rect 17648 5550 18608 5588
rect 17648 5533 17850 5550
rect 17388 5516 17404 5533
rect 16816 5500 17404 5516
rect 17834 5516 17850 5533
rect 18406 5533 18608 5550
rect 18666 5550 19626 5588
rect 18666 5533 18868 5550
rect 18406 5516 18422 5533
rect 17834 5500 18422 5516
rect 18852 5516 18868 5533
rect 19424 5533 19626 5550
rect 19684 5550 20644 5588
rect 19684 5533 19886 5550
rect 19424 5516 19440 5533
rect 18852 5500 19440 5516
rect 19870 5516 19886 5533
rect 20442 5533 20644 5550
rect 20702 5550 21662 5588
rect 20702 5533 20904 5550
rect 20442 5516 20458 5533
rect 19870 5500 20458 5516
rect 20888 5516 20904 5533
rect 21460 5533 21662 5550
rect 21720 5550 22680 5588
rect 21720 5533 21922 5550
rect 21460 5516 21476 5533
rect 20888 5500 21476 5516
rect 21906 5516 21922 5533
rect 22478 5533 22680 5550
rect 22738 5550 23698 5588
rect 22738 5533 22940 5550
rect 22478 5516 22494 5533
rect 21906 5500 22494 5516
rect 22924 5516 22940 5533
rect 23496 5533 23698 5550
rect 23756 5550 24716 5588
rect 23756 5533 23958 5550
rect 23496 5516 23512 5533
rect 22924 5500 23512 5516
rect 23942 5516 23958 5533
rect 24514 5533 24716 5550
rect 24774 5550 25734 5588
rect 24774 5533 24976 5550
rect 24514 5516 24530 5533
rect 23942 5500 24530 5516
rect 24960 5516 24976 5533
rect 25532 5533 25734 5550
rect 25792 5550 26752 5588
rect 25792 5533 25994 5550
rect 25532 5516 25548 5533
rect 24960 5500 25548 5516
rect 25978 5516 25994 5533
rect 26550 5533 26752 5550
rect 26810 5550 27770 5588
rect 26810 5533 27012 5550
rect 26550 5516 26566 5533
rect 25978 5500 26566 5516
rect 26996 5516 27012 5533
rect 27568 5533 27770 5550
rect 27828 5550 28788 5588
rect 27828 5533 28030 5550
rect 27568 5516 27584 5533
rect 26996 5500 27584 5516
rect 28014 5516 28030 5533
rect 28586 5533 28788 5550
rect 28846 5550 29806 5588
rect 28846 5533 29048 5550
rect 28586 5516 28602 5533
rect 28014 5500 28602 5516
rect 29032 5516 29048 5533
rect 29604 5533 29806 5550
rect 29864 5550 30824 5588
rect 29864 5533 30066 5550
rect 29604 5516 29620 5533
rect 29032 5500 29620 5516
rect 30050 5516 30066 5533
rect 30622 5533 30824 5550
rect 30882 5550 31842 5588
rect 30882 5533 31084 5550
rect 30622 5516 30638 5533
rect 30050 5500 30638 5516
rect 31068 5516 31084 5533
rect 31640 5533 31842 5550
rect 31900 5550 32860 5588
rect 31900 5533 32102 5550
rect 31640 5516 31656 5533
rect 31068 5500 31656 5516
rect 32086 5516 32102 5533
rect 32658 5533 32860 5550
rect 32918 5550 33878 5588
rect 32918 5533 33120 5550
rect 32658 5516 32674 5533
rect 32086 5500 32674 5516
rect 33104 5516 33120 5533
rect 33676 5533 33878 5550
rect 33676 5516 33692 5533
rect 33104 5500 33692 5516
rect 13762 5028 14350 5044
rect 13762 5011 13778 5028
rect 13576 4994 13778 5011
rect 14334 5011 14350 5028
rect 14780 5028 15368 5044
rect 14780 5011 14796 5028
rect 14334 4994 14536 5011
rect 13576 4956 14536 4994
rect 14594 4994 14796 5011
rect 15352 5011 15368 5028
rect 15798 5028 16386 5044
rect 15798 5011 15814 5028
rect 15352 4994 15554 5011
rect 14594 4956 15554 4994
rect 15612 4994 15814 5011
rect 16370 5011 16386 5028
rect 16816 5028 17404 5044
rect 16816 5011 16832 5028
rect 16370 4994 16572 5011
rect 15612 4956 16572 4994
rect 16630 4994 16832 5011
rect 17388 5011 17404 5028
rect 17834 5028 18422 5044
rect 17834 5011 17850 5028
rect 17388 4994 17590 5011
rect 16630 4956 17590 4994
rect 17648 4994 17850 5011
rect 18406 5011 18422 5028
rect 18852 5028 19440 5044
rect 18852 5011 18868 5028
rect 18406 4994 18608 5011
rect 17648 4956 18608 4994
rect 18666 4994 18868 5011
rect 19424 5011 19440 5028
rect 19870 5028 20458 5044
rect 19870 5011 19886 5028
rect 19424 4994 19626 5011
rect 18666 4956 19626 4994
rect 19684 4994 19886 5011
rect 20442 5011 20458 5028
rect 20888 5028 21476 5044
rect 20888 5011 20904 5028
rect 20442 4994 20644 5011
rect 19684 4956 20644 4994
rect 20702 4994 20904 5011
rect 21460 5011 21476 5028
rect 21906 5028 22494 5044
rect 21906 5011 21922 5028
rect 21460 4994 21662 5011
rect 20702 4956 21662 4994
rect 21720 4994 21922 5011
rect 22478 5011 22494 5028
rect 22924 5028 23512 5044
rect 22924 5011 22940 5028
rect 22478 4994 22680 5011
rect 21720 4956 22680 4994
rect 22738 4994 22940 5011
rect 23496 5011 23512 5028
rect 23942 5028 24530 5044
rect 23942 5011 23958 5028
rect 23496 4994 23698 5011
rect 22738 4956 23698 4994
rect 23756 4994 23958 5011
rect 24514 5011 24530 5028
rect 24960 5028 25548 5044
rect 24960 5011 24976 5028
rect 24514 4994 24716 5011
rect 23756 4956 24716 4994
rect 24774 4994 24976 5011
rect 25532 5011 25548 5028
rect 25978 5028 26566 5044
rect 25978 5011 25994 5028
rect 25532 4994 25734 5011
rect 24774 4956 25734 4994
rect 25792 4994 25994 5011
rect 26550 5011 26566 5028
rect 26996 5028 27584 5044
rect 26996 5011 27012 5028
rect 26550 4994 26752 5011
rect 25792 4956 26752 4994
rect 26810 4994 27012 5011
rect 27568 5011 27584 5028
rect 28014 5028 28602 5044
rect 28014 5011 28030 5028
rect 27568 4994 27770 5011
rect 26810 4956 27770 4994
rect 27828 4994 28030 5011
rect 28586 5011 28602 5028
rect 29032 5028 29620 5044
rect 29032 5011 29048 5028
rect 28586 4994 28788 5011
rect 27828 4956 28788 4994
rect 28846 4994 29048 5011
rect 29604 5011 29620 5028
rect 30050 5028 30638 5044
rect 30050 5011 30066 5028
rect 29604 4994 29806 5011
rect 28846 4956 29806 4994
rect 29864 4994 30066 5011
rect 30622 5011 30638 5028
rect 31068 5028 31656 5044
rect 31068 5011 31084 5028
rect 30622 4994 30824 5011
rect 29864 4956 30824 4994
rect 30882 4994 31084 5011
rect 31640 5011 31656 5028
rect 32086 5028 32674 5044
rect 32086 5011 32102 5028
rect 31640 4994 31842 5011
rect 30882 4956 31842 4994
rect 31900 4994 32102 5011
rect 32658 5011 32674 5028
rect 33104 5028 33692 5044
rect 33104 5011 33120 5028
rect 32658 4994 32860 5011
rect 31900 4956 32860 4994
rect 32918 4994 33120 5011
rect 33676 5011 33692 5028
rect 33676 4994 33878 5011
rect 32918 4956 33878 4994
rect 1777 4831 2365 4847
rect 1777 4814 1793 4831
rect 1591 4797 1793 4814
rect 2349 4814 2365 4831
rect 2795 4831 3383 4847
rect 2795 4814 2811 4831
rect 2349 4797 2551 4814
rect 1591 4759 2551 4797
rect 2609 4797 2811 4814
rect 3367 4814 3383 4831
rect 3813 4831 4401 4847
rect 3813 4814 3829 4831
rect 3367 4797 3569 4814
rect 2609 4759 3569 4797
rect 3627 4797 3829 4814
rect 4385 4814 4401 4831
rect 4831 4831 5419 4847
rect 4831 4814 4847 4831
rect 4385 4797 4587 4814
rect 3627 4759 4587 4797
rect 4645 4797 4847 4814
rect 5403 4814 5419 4831
rect 5849 4831 6437 4847
rect 5849 4814 5865 4831
rect 5403 4797 5605 4814
rect 4645 4759 5605 4797
rect 5663 4797 5865 4814
rect 6421 4814 6437 4831
rect 6867 4831 7455 4847
rect 6867 4814 6883 4831
rect 6421 4797 6623 4814
rect 5663 4759 6623 4797
rect 6681 4797 6883 4814
rect 7439 4814 7455 4831
rect 8628 4832 8784 4848
rect 8628 4815 8644 4832
rect 7439 4797 7641 4814
rect 6681 4759 7641 4797
rect 8586 4798 8644 4815
rect 8768 4815 8784 4832
rect 8926 4832 9082 4848
rect 8926 4815 8942 4832
rect 8768 4798 8826 4815
rect 8586 4760 8826 4798
rect 8884 4798 8942 4815
rect 9066 4815 9082 4832
rect 9224 4832 9380 4848
rect 9224 4815 9240 4832
rect 9066 4798 9124 4815
rect 8884 4760 9124 4798
rect 9182 4798 9240 4815
rect 9364 4815 9380 4832
rect 9522 4832 9678 4848
rect 9522 4815 9538 4832
rect 9364 4798 9422 4815
rect 9182 4760 9422 4798
rect 9480 4798 9538 4815
rect 9662 4815 9678 4832
rect 9820 4832 9976 4848
rect 9820 4815 9836 4832
rect 9662 4798 9720 4815
rect 9480 4760 9720 4798
rect 9778 4798 9836 4815
rect 9960 4815 9976 4832
rect 10118 4832 10274 4848
rect 10118 4815 10134 4832
rect 9960 4798 10018 4815
rect 9778 4760 10018 4798
rect 10076 4798 10134 4815
rect 10258 4815 10274 4832
rect 10416 4832 10572 4848
rect 10416 4815 10432 4832
rect 10258 4798 10316 4815
rect 10076 4760 10316 4798
rect 10374 4798 10432 4815
rect 10556 4815 10572 4832
rect 10714 4832 10870 4848
rect 10714 4815 10730 4832
rect 10556 4798 10614 4815
rect 10374 4760 10614 4798
rect 10672 4798 10730 4815
rect 10854 4815 10870 4832
rect 11012 4832 11168 4848
rect 11012 4815 11028 4832
rect 10854 4798 10912 4815
rect 10672 4760 10912 4798
rect 10970 4798 11028 4815
rect 11152 4815 11168 4832
rect 11310 4832 11466 4848
rect 11310 4815 11326 4832
rect 11152 4798 11210 4815
rect 10970 4760 11210 4798
rect 11268 4798 11326 4815
rect 11450 4815 11466 4832
rect 11608 4832 11764 4848
rect 11608 4815 11624 4832
rect 11450 4798 11508 4815
rect 11268 4760 11508 4798
rect 11566 4798 11624 4815
rect 11748 4815 11764 4832
rect 11748 4798 11806 4815
rect 11566 4760 11806 4798
rect 13576 4318 14536 4356
rect 13576 4301 13778 4318
rect 13762 4284 13778 4301
rect 14334 4301 14536 4318
rect 14594 4318 15554 4356
rect 14594 4301 14796 4318
rect 14334 4284 14350 4301
rect 13762 4268 14350 4284
rect 14780 4284 14796 4301
rect 15352 4301 15554 4318
rect 15612 4318 16572 4356
rect 15612 4301 15814 4318
rect 15352 4284 15368 4301
rect 14780 4268 15368 4284
rect 15798 4284 15814 4301
rect 16370 4301 16572 4318
rect 16630 4318 17590 4356
rect 16630 4301 16832 4318
rect 16370 4284 16386 4301
rect 15798 4268 16386 4284
rect 16816 4284 16832 4301
rect 17388 4301 17590 4318
rect 17648 4318 18608 4356
rect 17648 4301 17850 4318
rect 17388 4284 17404 4301
rect 16816 4268 17404 4284
rect 17834 4284 17850 4301
rect 18406 4301 18608 4318
rect 18666 4318 19626 4356
rect 18666 4301 18868 4318
rect 18406 4284 18422 4301
rect 17834 4268 18422 4284
rect 18852 4284 18868 4301
rect 19424 4301 19626 4318
rect 19684 4318 20644 4356
rect 19684 4301 19886 4318
rect 19424 4284 19440 4301
rect 18852 4268 19440 4284
rect 19870 4284 19886 4301
rect 20442 4301 20644 4318
rect 20702 4318 21662 4356
rect 20702 4301 20904 4318
rect 20442 4284 20458 4301
rect 19870 4268 20458 4284
rect 20888 4284 20904 4301
rect 21460 4301 21662 4318
rect 21720 4318 22680 4356
rect 21720 4301 21922 4318
rect 21460 4284 21476 4301
rect 20888 4268 21476 4284
rect 21906 4284 21922 4301
rect 22478 4301 22680 4318
rect 22738 4318 23698 4356
rect 22738 4301 22940 4318
rect 22478 4284 22494 4301
rect 21906 4268 22494 4284
rect 22924 4284 22940 4301
rect 23496 4301 23698 4318
rect 23756 4318 24716 4356
rect 23756 4301 23958 4318
rect 23496 4284 23512 4301
rect 22924 4268 23512 4284
rect 23942 4284 23958 4301
rect 24514 4301 24716 4318
rect 24774 4318 25734 4356
rect 24774 4301 24976 4318
rect 24514 4284 24530 4301
rect 23942 4268 24530 4284
rect 24960 4284 24976 4301
rect 25532 4301 25734 4318
rect 25792 4318 26752 4356
rect 25792 4301 25994 4318
rect 25532 4284 25548 4301
rect 24960 4268 25548 4284
rect 25978 4284 25994 4301
rect 26550 4301 26752 4318
rect 26810 4318 27770 4356
rect 26810 4301 27012 4318
rect 26550 4284 26566 4301
rect 25978 4268 26566 4284
rect 26996 4284 27012 4301
rect 27568 4301 27770 4318
rect 27828 4318 28788 4356
rect 27828 4301 28030 4318
rect 27568 4284 27584 4301
rect 26996 4268 27584 4284
rect 28014 4284 28030 4301
rect 28586 4301 28788 4318
rect 28846 4318 29806 4356
rect 28846 4301 29048 4318
rect 28586 4284 28602 4301
rect 28014 4268 28602 4284
rect 29032 4284 29048 4301
rect 29604 4301 29806 4318
rect 29864 4318 30824 4356
rect 29864 4301 30066 4318
rect 29604 4284 29620 4301
rect 29032 4268 29620 4284
rect 30050 4284 30066 4301
rect 30622 4301 30824 4318
rect 30882 4318 31842 4356
rect 30882 4301 31084 4318
rect 30622 4284 30638 4301
rect 30050 4268 30638 4284
rect 31068 4284 31084 4301
rect 31640 4301 31842 4318
rect 31900 4318 32860 4356
rect 31900 4301 32102 4318
rect 31640 4284 31656 4301
rect 31068 4268 31656 4284
rect 32086 4284 32102 4301
rect 32658 4301 32860 4318
rect 32918 4318 33878 4356
rect 32918 4301 33120 4318
rect 32658 4284 32674 4301
rect 32086 4268 32674 4284
rect 33104 4284 33120 4301
rect 33676 4301 33878 4318
rect 33676 4284 33692 4301
rect 33104 4268 33692 4284
rect 1591 4121 2551 4159
rect 1591 4104 1793 4121
rect 1777 4087 1793 4104
rect 2349 4104 2551 4121
rect 2609 4121 3569 4159
rect 2609 4104 2811 4121
rect 2349 4087 2365 4104
rect 1777 4071 2365 4087
rect 2795 4087 2811 4104
rect 3367 4104 3569 4121
rect 3627 4121 4587 4159
rect 3627 4104 3829 4121
rect 3367 4087 3383 4104
rect 2795 4071 3383 4087
rect 3813 4087 3829 4104
rect 4385 4104 4587 4121
rect 4645 4121 5605 4159
rect 4645 4104 4847 4121
rect 4385 4087 4401 4104
rect 3813 4071 4401 4087
rect 4831 4087 4847 4104
rect 5403 4104 5605 4121
rect 5663 4121 6623 4159
rect 5663 4104 5865 4121
rect 5403 4087 5419 4104
rect 4831 4071 5419 4087
rect 5849 4087 5865 4104
rect 6421 4104 6623 4121
rect 6681 4121 7641 4159
rect 6681 4104 6883 4121
rect 6421 4087 6437 4104
rect 5849 4071 6437 4087
rect 6867 4087 6883 4104
rect 7439 4104 7641 4121
rect 8586 4122 8826 4160
rect 8586 4105 8644 4122
rect 7439 4087 7455 4104
rect 6867 4071 7455 4087
rect 8628 4088 8644 4105
rect 8768 4105 8826 4122
rect 8884 4122 9124 4160
rect 8884 4105 8942 4122
rect 8768 4088 8784 4105
rect 8628 4072 8784 4088
rect 8926 4088 8942 4105
rect 9066 4105 9124 4122
rect 9182 4122 9422 4160
rect 9182 4105 9240 4122
rect 9066 4088 9082 4105
rect 8926 4072 9082 4088
rect 9224 4088 9240 4105
rect 9364 4105 9422 4122
rect 9480 4122 9720 4160
rect 9480 4105 9538 4122
rect 9364 4088 9380 4105
rect 9224 4072 9380 4088
rect 9522 4088 9538 4105
rect 9662 4105 9720 4122
rect 9778 4122 10018 4160
rect 9778 4105 9836 4122
rect 9662 4088 9678 4105
rect 9522 4072 9678 4088
rect 9820 4088 9836 4105
rect 9960 4105 10018 4122
rect 10076 4122 10316 4160
rect 10076 4105 10134 4122
rect 9960 4088 9976 4105
rect 9820 4072 9976 4088
rect 10118 4088 10134 4105
rect 10258 4105 10316 4122
rect 10374 4122 10614 4160
rect 10374 4105 10432 4122
rect 10258 4088 10274 4105
rect 10118 4072 10274 4088
rect 10416 4088 10432 4105
rect 10556 4105 10614 4122
rect 10672 4122 10912 4160
rect 10672 4105 10730 4122
rect 10556 4088 10572 4105
rect 10416 4072 10572 4088
rect 10714 4088 10730 4105
rect 10854 4105 10912 4122
rect 10970 4122 11210 4160
rect 10970 4105 11028 4122
rect 10854 4088 10870 4105
rect 10714 4072 10870 4088
rect 11012 4088 11028 4105
rect 11152 4105 11210 4122
rect 11268 4122 11508 4160
rect 11268 4105 11326 4122
rect 11152 4088 11168 4105
rect 11012 4072 11168 4088
rect 11310 4088 11326 4105
rect 11450 4105 11508 4122
rect 11566 4122 11806 4160
rect 11566 4105 11624 4122
rect 11450 4088 11466 4105
rect 11310 4072 11466 4088
rect 11608 4088 11624 4105
rect 11748 4105 11806 4122
rect 11748 4088 11764 4105
rect 11608 4072 11764 4088
rect 13762 3794 14350 3810
rect 13762 3777 13778 3794
rect 13576 3760 13778 3777
rect 14334 3777 14350 3794
rect 14780 3794 15368 3810
rect 14780 3777 14796 3794
rect 14334 3760 14536 3777
rect 1776 3718 2364 3734
rect 1776 3701 1792 3718
rect 1590 3684 1792 3701
rect 2348 3701 2364 3718
rect 2794 3718 3382 3734
rect 2794 3701 2810 3718
rect 2348 3684 2550 3701
rect 1590 3646 2550 3684
rect 2608 3684 2810 3701
rect 3366 3701 3382 3718
rect 3812 3718 4400 3734
rect 3812 3701 3828 3718
rect 3366 3684 3568 3701
rect 2608 3646 3568 3684
rect 3626 3684 3828 3701
rect 4384 3701 4400 3718
rect 4830 3718 5418 3734
rect 4830 3701 4846 3718
rect 4384 3684 4586 3701
rect 3626 3646 4586 3684
rect 4644 3684 4846 3701
rect 5402 3701 5418 3718
rect 5848 3718 6436 3734
rect 5848 3701 5864 3718
rect 5402 3684 5604 3701
rect 4644 3646 5604 3684
rect 5662 3684 5864 3701
rect 6420 3701 6436 3718
rect 6866 3718 7454 3734
rect 6866 3701 6882 3718
rect 6420 3684 6622 3701
rect 5662 3646 6622 3684
rect 6680 3684 6882 3701
rect 7438 3701 7454 3718
rect 8628 3720 8784 3736
rect 8628 3703 8644 3720
rect 7438 3684 7640 3701
rect 6680 3646 7640 3684
rect 8586 3686 8644 3703
rect 8768 3703 8784 3720
rect 8926 3720 9082 3736
rect 8926 3703 8942 3720
rect 8768 3686 8826 3703
rect 8586 3648 8826 3686
rect 8884 3686 8942 3703
rect 9066 3703 9082 3720
rect 9224 3720 9380 3736
rect 9224 3703 9240 3720
rect 9066 3686 9124 3703
rect 8884 3648 9124 3686
rect 9182 3686 9240 3703
rect 9364 3703 9380 3720
rect 9522 3720 9678 3736
rect 9522 3703 9538 3720
rect 9364 3686 9422 3703
rect 9182 3648 9422 3686
rect 9480 3686 9538 3703
rect 9662 3703 9678 3720
rect 9820 3720 9976 3736
rect 9820 3703 9836 3720
rect 9662 3686 9720 3703
rect 9480 3648 9720 3686
rect 9778 3686 9836 3703
rect 9960 3703 9976 3720
rect 10118 3720 10274 3736
rect 10118 3703 10134 3720
rect 9960 3686 10018 3703
rect 9778 3648 10018 3686
rect 10076 3686 10134 3703
rect 10258 3703 10274 3720
rect 10416 3720 10572 3736
rect 10416 3703 10432 3720
rect 10258 3686 10316 3703
rect 10076 3648 10316 3686
rect 10374 3686 10432 3703
rect 10556 3703 10572 3720
rect 10714 3720 10870 3736
rect 10714 3703 10730 3720
rect 10556 3686 10614 3703
rect 10374 3648 10614 3686
rect 10672 3686 10730 3703
rect 10854 3703 10870 3720
rect 11012 3720 11168 3736
rect 11012 3703 11028 3720
rect 10854 3686 10912 3703
rect 10672 3648 10912 3686
rect 10970 3686 11028 3703
rect 11152 3703 11168 3720
rect 11310 3720 11466 3736
rect 11310 3703 11326 3720
rect 11152 3686 11210 3703
rect 10970 3648 11210 3686
rect 11268 3686 11326 3703
rect 11450 3703 11466 3720
rect 11608 3720 11764 3736
rect 13576 3722 14536 3760
rect 14594 3760 14796 3777
rect 15352 3777 15368 3794
rect 15798 3794 16386 3810
rect 15798 3777 15814 3794
rect 15352 3760 15554 3777
rect 14594 3722 15554 3760
rect 15612 3760 15814 3777
rect 16370 3777 16386 3794
rect 16816 3794 17404 3810
rect 16816 3777 16832 3794
rect 16370 3760 16572 3777
rect 15612 3722 16572 3760
rect 16630 3760 16832 3777
rect 17388 3777 17404 3794
rect 17834 3794 18422 3810
rect 17834 3777 17850 3794
rect 17388 3760 17590 3777
rect 16630 3722 17590 3760
rect 17648 3760 17850 3777
rect 18406 3777 18422 3794
rect 18852 3794 19440 3810
rect 18852 3777 18868 3794
rect 18406 3760 18608 3777
rect 17648 3722 18608 3760
rect 18666 3760 18868 3777
rect 19424 3777 19440 3794
rect 19870 3794 20458 3810
rect 19870 3777 19886 3794
rect 19424 3760 19626 3777
rect 18666 3722 19626 3760
rect 19684 3760 19886 3777
rect 20442 3777 20458 3794
rect 20888 3794 21476 3810
rect 20888 3777 20904 3794
rect 20442 3760 20644 3777
rect 19684 3722 20644 3760
rect 20702 3760 20904 3777
rect 21460 3777 21476 3794
rect 21906 3794 22494 3810
rect 21906 3777 21922 3794
rect 21460 3760 21662 3777
rect 20702 3722 21662 3760
rect 21720 3760 21922 3777
rect 22478 3777 22494 3794
rect 22924 3794 23512 3810
rect 22924 3777 22940 3794
rect 22478 3760 22680 3777
rect 21720 3722 22680 3760
rect 22738 3760 22940 3777
rect 23496 3777 23512 3794
rect 23942 3794 24530 3810
rect 23942 3777 23958 3794
rect 23496 3760 23698 3777
rect 22738 3722 23698 3760
rect 23756 3760 23958 3777
rect 24514 3777 24530 3794
rect 24960 3794 25548 3810
rect 24960 3777 24976 3794
rect 24514 3760 24716 3777
rect 23756 3722 24716 3760
rect 24774 3760 24976 3777
rect 25532 3777 25548 3794
rect 25978 3794 26566 3810
rect 25978 3777 25994 3794
rect 25532 3760 25734 3777
rect 24774 3722 25734 3760
rect 25792 3760 25994 3777
rect 26550 3777 26566 3794
rect 26996 3794 27584 3810
rect 26996 3777 27012 3794
rect 26550 3760 26752 3777
rect 25792 3722 26752 3760
rect 26810 3760 27012 3777
rect 27568 3777 27584 3794
rect 28014 3794 28602 3810
rect 28014 3777 28030 3794
rect 27568 3760 27770 3777
rect 26810 3722 27770 3760
rect 27828 3760 28030 3777
rect 28586 3777 28602 3794
rect 29032 3794 29620 3810
rect 29032 3777 29048 3794
rect 28586 3760 28788 3777
rect 27828 3722 28788 3760
rect 28846 3760 29048 3777
rect 29604 3777 29620 3794
rect 30050 3794 30638 3810
rect 30050 3777 30066 3794
rect 29604 3760 29806 3777
rect 28846 3722 29806 3760
rect 29864 3760 30066 3777
rect 30622 3777 30638 3794
rect 31068 3794 31656 3810
rect 31068 3777 31084 3794
rect 30622 3760 30824 3777
rect 29864 3722 30824 3760
rect 30882 3760 31084 3777
rect 31640 3777 31656 3794
rect 32086 3794 32674 3810
rect 32086 3777 32102 3794
rect 31640 3760 31842 3777
rect 30882 3722 31842 3760
rect 31900 3760 32102 3777
rect 32658 3777 32674 3794
rect 33104 3794 33692 3810
rect 33104 3777 33120 3794
rect 32658 3760 32860 3777
rect 31900 3722 32860 3760
rect 32918 3760 33120 3777
rect 33676 3777 33692 3794
rect 33676 3760 33878 3777
rect 32918 3722 33878 3760
rect 11608 3703 11624 3720
rect 11450 3686 11508 3703
rect 11268 3648 11508 3686
rect 11566 3686 11624 3703
rect 11748 3703 11764 3720
rect 11748 3686 11806 3703
rect 11566 3648 11806 3686
rect 13576 3084 14536 3122
rect 13576 3067 13778 3084
rect 13762 3050 13778 3067
rect 14334 3067 14536 3084
rect 14594 3084 15554 3122
rect 14594 3067 14796 3084
rect 14334 3050 14350 3067
rect 1590 3008 2550 3046
rect 1590 2991 1792 3008
rect 1776 2974 1792 2991
rect 2348 2991 2550 3008
rect 2608 3008 3568 3046
rect 2608 2991 2810 3008
rect 2348 2974 2364 2991
rect 1776 2958 2364 2974
rect 2794 2974 2810 2991
rect 3366 2991 3568 3008
rect 3626 3008 4586 3046
rect 3626 2991 3828 3008
rect 3366 2974 3382 2991
rect 2794 2958 3382 2974
rect 3812 2974 3828 2991
rect 4384 2991 4586 3008
rect 4644 3008 5604 3046
rect 4644 2991 4846 3008
rect 4384 2974 4400 2991
rect 3812 2958 4400 2974
rect 4830 2974 4846 2991
rect 5402 2991 5604 3008
rect 5662 3008 6622 3046
rect 5662 2991 5864 3008
rect 5402 2974 5418 2991
rect 4830 2958 5418 2974
rect 5848 2974 5864 2991
rect 6420 2991 6622 3008
rect 6680 3008 7640 3046
rect 6680 2991 6882 3008
rect 6420 2974 6436 2991
rect 5848 2958 6436 2974
rect 6866 2974 6882 2991
rect 7438 2991 7640 3008
rect 8586 3010 8826 3048
rect 8586 2993 8644 3010
rect 7438 2974 7454 2991
rect 6866 2958 7454 2974
rect 8628 2976 8644 2993
rect 8768 2993 8826 3010
rect 8884 3010 9124 3048
rect 8884 2993 8942 3010
rect 8768 2976 8784 2993
rect 8628 2960 8784 2976
rect 8926 2976 8942 2993
rect 9066 2993 9124 3010
rect 9182 3010 9422 3048
rect 9182 2993 9240 3010
rect 9066 2976 9082 2993
rect 8926 2960 9082 2976
rect 9224 2976 9240 2993
rect 9364 2993 9422 3010
rect 9480 3010 9720 3048
rect 9480 2993 9538 3010
rect 9364 2976 9380 2993
rect 9224 2960 9380 2976
rect 9522 2976 9538 2993
rect 9662 2993 9720 3010
rect 9778 3010 10018 3048
rect 9778 2993 9836 3010
rect 9662 2976 9678 2993
rect 9522 2960 9678 2976
rect 9820 2976 9836 2993
rect 9960 2993 10018 3010
rect 10076 3010 10316 3048
rect 10076 2993 10134 3010
rect 9960 2976 9976 2993
rect 9820 2960 9976 2976
rect 10118 2976 10134 2993
rect 10258 2993 10316 3010
rect 10374 3010 10614 3048
rect 10374 2993 10432 3010
rect 10258 2976 10274 2993
rect 10118 2960 10274 2976
rect 10416 2976 10432 2993
rect 10556 2993 10614 3010
rect 10672 3010 10912 3048
rect 10672 2993 10730 3010
rect 10556 2976 10572 2993
rect 10416 2960 10572 2976
rect 10714 2976 10730 2993
rect 10854 2993 10912 3010
rect 10970 3010 11210 3048
rect 10970 2993 11028 3010
rect 10854 2976 10870 2993
rect 10714 2960 10870 2976
rect 11012 2976 11028 2993
rect 11152 2993 11210 3010
rect 11268 3010 11508 3048
rect 11268 2993 11326 3010
rect 11152 2976 11168 2993
rect 11012 2960 11168 2976
rect 11310 2976 11326 2993
rect 11450 2993 11508 3010
rect 11566 3010 11806 3048
rect 13762 3034 14350 3050
rect 14780 3050 14796 3067
rect 15352 3067 15554 3084
rect 15612 3084 16572 3122
rect 15612 3067 15814 3084
rect 15352 3050 15368 3067
rect 14780 3034 15368 3050
rect 15798 3050 15814 3067
rect 16370 3067 16572 3084
rect 16630 3084 17590 3122
rect 16630 3067 16832 3084
rect 16370 3050 16386 3067
rect 15798 3034 16386 3050
rect 16816 3050 16832 3067
rect 17388 3067 17590 3084
rect 17648 3084 18608 3122
rect 17648 3067 17850 3084
rect 17388 3050 17404 3067
rect 16816 3034 17404 3050
rect 17834 3050 17850 3067
rect 18406 3067 18608 3084
rect 18666 3084 19626 3122
rect 18666 3067 18868 3084
rect 18406 3050 18422 3067
rect 17834 3034 18422 3050
rect 18852 3050 18868 3067
rect 19424 3067 19626 3084
rect 19684 3084 20644 3122
rect 19684 3067 19886 3084
rect 19424 3050 19440 3067
rect 18852 3034 19440 3050
rect 19870 3050 19886 3067
rect 20442 3067 20644 3084
rect 20702 3084 21662 3122
rect 20702 3067 20904 3084
rect 20442 3050 20458 3067
rect 19870 3034 20458 3050
rect 20888 3050 20904 3067
rect 21460 3067 21662 3084
rect 21720 3084 22680 3122
rect 21720 3067 21922 3084
rect 21460 3050 21476 3067
rect 20888 3034 21476 3050
rect 21906 3050 21922 3067
rect 22478 3067 22680 3084
rect 22738 3084 23698 3122
rect 22738 3067 22940 3084
rect 22478 3050 22494 3067
rect 21906 3034 22494 3050
rect 22924 3050 22940 3067
rect 23496 3067 23698 3084
rect 23756 3084 24716 3122
rect 23756 3067 23958 3084
rect 23496 3050 23512 3067
rect 22924 3034 23512 3050
rect 23942 3050 23958 3067
rect 24514 3067 24716 3084
rect 24774 3084 25734 3122
rect 24774 3067 24976 3084
rect 24514 3050 24530 3067
rect 23942 3034 24530 3050
rect 24960 3050 24976 3067
rect 25532 3067 25734 3084
rect 25792 3084 26752 3122
rect 25792 3067 25994 3084
rect 25532 3050 25548 3067
rect 24960 3034 25548 3050
rect 25978 3050 25994 3067
rect 26550 3067 26752 3084
rect 26810 3084 27770 3122
rect 26810 3067 27012 3084
rect 26550 3050 26566 3067
rect 25978 3034 26566 3050
rect 26996 3050 27012 3067
rect 27568 3067 27770 3084
rect 27828 3084 28788 3122
rect 27828 3067 28030 3084
rect 27568 3050 27584 3067
rect 26996 3034 27584 3050
rect 28014 3050 28030 3067
rect 28586 3067 28788 3084
rect 28846 3084 29806 3122
rect 28846 3067 29048 3084
rect 28586 3050 28602 3067
rect 28014 3034 28602 3050
rect 29032 3050 29048 3067
rect 29604 3067 29806 3084
rect 29864 3084 30824 3122
rect 29864 3067 30066 3084
rect 29604 3050 29620 3067
rect 29032 3034 29620 3050
rect 30050 3050 30066 3067
rect 30622 3067 30824 3084
rect 30882 3084 31842 3122
rect 30882 3067 31084 3084
rect 30622 3050 30638 3067
rect 30050 3034 30638 3050
rect 31068 3050 31084 3067
rect 31640 3067 31842 3084
rect 31900 3084 32860 3122
rect 31900 3067 32102 3084
rect 31640 3050 31656 3067
rect 31068 3034 31656 3050
rect 32086 3050 32102 3067
rect 32658 3067 32860 3084
rect 32918 3084 33878 3122
rect 32918 3067 33120 3084
rect 32658 3050 32674 3067
rect 32086 3034 32674 3050
rect 33104 3050 33120 3067
rect 33676 3067 33878 3084
rect 33676 3050 33692 3067
rect 33104 3034 33692 3050
rect 11566 2993 11624 3010
rect 11450 2976 11466 2993
rect 11310 2960 11466 2976
rect 11608 2976 11624 2993
rect 11748 2993 11806 3010
rect 11748 2976 11764 2993
rect 11608 2960 11764 2976
rect 1777 2607 2365 2623
rect 1777 2590 1793 2607
rect 1591 2573 1793 2590
rect 2349 2590 2365 2607
rect 2795 2607 3383 2623
rect 2795 2590 2811 2607
rect 2349 2573 2551 2590
rect 1591 2535 2551 2573
rect 2609 2573 2811 2590
rect 3367 2590 3383 2607
rect 3813 2607 4401 2623
rect 3813 2590 3829 2607
rect 3367 2573 3569 2590
rect 2609 2535 3569 2573
rect 3627 2573 3829 2590
rect 4385 2590 4401 2607
rect 4831 2607 5419 2623
rect 4831 2590 4847 2607
rect 4385 2573 4587 2590
rect 3627 2535 4587 2573
rect 4645 2573 4847 2590
rect 5403 2590 5419 2607
rect 5849 2607 6437 2623
rect 5849 2590 5865 2607
rect 5403 2573 5605 2590
rect 4645 2535 5605 2573
rect 5663 2573 5865 2590
rect 6421 2590 6437 2607
rect 6867 2607 7455 2623
rect 6867 2590 6883 2607
rect 6421 2573 6623 2590
rect 5663 2535 6623 2573
rect 6681 2573 6883 2590
rect 7439 2590 7455 2607
rect 8626 2608 8782 2624
rect 8626 2591 8642 2608
rect 7439 2573 7641 2590
rect 6681 2535 7641 2573
rect 8584 2574 8642 2591
rect 8766 2591 8782 2608
rect 8924 2608 9080 2624
rect 8924 2591 8940 2608
rect 8766 2574 8824 2591
rect 8584 2536 8824 2574
rect 8882 2574 8940 2591
rect 9064 2591 9080 2608
rect 9222 2608 9378 2624
rect 9222 2591 9238 2608
rect 9064 2574 9122 2591
rect 8882 2536 9122 2574
rect 9180 2574 9238 2591
rect 9362 2591 9378 2608
rect 9520 2608 9676 2624
rect 9520 2591 9536 2608
rect 9362 2574 9420 2591
rect 9180 2536 9420 2574
rect 9478 2574 9536 2591
rect 9660 2591 9676 2608
rect 9818 2608 9974 2624
rect 9818 2591 9834 2608
rect 9660 2574 9718 2591
rect 9478 2536 9718 2574
rect 9776 2574 9834 2591
rect 9958 2591 9974 2608
rect 10116 2608 10272 2624
rect 10116 2591 10132 2608
rect 9958 2574 10016 2591
rect 9776 2536 10016 2574
rect 10074 2574 10132 2591
rect 10256 2591 10272 2608
rect 10414 2608 10570 2624
rect 10414 2591 10430 2608
rect 10256 2574 10314 2591
rect 10074 2536 10314 2574
rect 10372 2574 10430 2591
rect 10554 2591 10570 2608
rect 10712 2608 10868 2624
rect 10712 2591 10728 2608
rect 10554 2574 10612 2591
rect 10372 2536 10612 2574
rect 10670 2574 10728 2591
rect 10852 2591 10868 2608
rect 11010 2608 11166 2624
rect 11010 2591 11026 2608
rect 10852 2574 10910 2591
rect 10670 2536 10910 2574
rect 10968 2574 11026 2591
rect 11150 2591 11166 2608
rect 11308 2608 11464 2624
rect 11308 2591 11324 2608
rect 11150 2574 11208 2591
rect 10968 2536 11208 2574
rect 11266 2574 11324 2591
rect 11448 2591 11464 2608
rect 11606 2608 11762 2624
rect 11606 2591 11622 2608
rect 11448 2574 11506 2591
rect 11266 2536 11506 2574
rect 11564 2574 11622 2591
rect 11746 2591 11762 2608
rect 11746 2574 11804 2591
rect 11564 2536 11804 2574
rect 13762 2560 14350 2576
rect 13762 2543 13778 2560
rect 13576 2526 13778 2543
rect 14334 2543 14350 2560
rect 14780 2560 15368 2576
rect 14780 2543 14796 2560
rect 14334 2526 14536 2543
rect 13576 2488 14536 2526
rect 14594 2526 14796 2543
rect 15352 2543 15368 2560
rect 15798 2560 16386 2576
rect 15798 2543 15814 2560
rect 15352 2526 15554 2543
rect 14594 2488 15554 2526
rect 15612 2526 15814 2543
rect 16370 2543 16386 2560
rect 16816 2560 17404 2576
rect 16816 2543 16832 2560
rect 16370 2526 16572 2543
rect 15612 2488 16572 2526
rect 16630 2526 16832 2543
rect 17388 2543 17404 2560
rect 17834 2560 18422 2576
rect 17834 2543 17850 2560
rect 17388 2526 17590 2543
rect 16630 2488 17590 2526
rect 17648 2526 17850 2543
rect 18406 2543 18422 2560
rect 18852 2560 19440 2576
rect 18852 2543 18868 2560
rect 18406 2526 18608 2543
rect 17648 2488 18608 2526
rect 18666 2526 18868 2543
rect 19424 2543 19440 2560
rect 19870 2560 20458 2576
rect 19870 2543 19886 2560
rect 19424 2526 19626 2543
rect 18666 2488 19626 2526
rect 19684 2526 19886 2543
rect 20442 2543 20458 2560
rect 20888 2560 21476 2576
rect 20888 2543 20904 2560
rect 20442 2526 20644 2543
rect 19684 2488 20644 2526
rect 20702 2526 20904 2543
rect 21460 2543 21476 2560
rect 21906 2560 22494 2576
rect 21906 2543 21922 2560
rect 21460 2526 21662 2543
rect 20702 2488 21662 2526
rect 21720 2526 21922 2543
rect 22478 2543 22494 2560
rect 22924 2560 23512 2576
rect 22924 2543 22940 2560
rect 22478 2526 22680 2543
rect 21720 2488 22680 2526
rect 22738 2526 22940 2543
rect 23496 2543 23512 2560
rect 23942 2560 24530 2576
rect 23942 2543 23958 2560
rect 23496 2526 23698 2543
rect 22738 2488 23698 2526
rect 23756 2526 23958 2543
rect 24514 2543 24530 2560
rect 24960 2560 25548 2576
rect 24960 2543 24976 2560
rect 24514 2526 24716 2543
rect 23756 2488 24716 2526
rect 24774 2526 24976 2543
rect 25532 2543 25548 2560
rect 25978 2560 26566 2576
rect 25978 2543 25994 2560
rect 25532 2526 25734 2543
rect 24774 2488 25734 2526
rect 25792 2526 25994 2543
rect 26550 2543 26566 2560
rect 26996 2560 27584 2576
rect 26996 2543 27012 2560
rect 26550 2526 26752 2543
rect 25792 2488 26752 2526
rect 26810 2526 27012 2543
rect 27568 2543 27584 2560
rect 28014 2560 28602 2576
rect 28014 2543 28030 2560
rect 27568 2526 27770 2543
rect 26810 2488 27770 2526
rect 27828 2526 28030 2543
rect 28586 2543 28602 2560
rect 29032 2560 29620 2576
rect 29032 2543 29048 2560
rect 28586 2526 28788 2543
rect 27828 2488 28788 2526
rect 28846 2526 29048 2543
rect 29604 2543 29620 2560
rect 30050 2560 30638 2576
rect 30050 2543 30066 2560
rect 29604 2526 29806 2543
rect 28846 2488 29806 2526
rect 29864 2526 30066 2543
rect 30622 2543 30638 2560
rect 31068 2560 31656 2576
rect 31068 2543 31084 2560
rect 30622 2526 30824 2543
rect 29864 2488 30824 2526
rect 30882 2526 31084 2543
rect 31640 2543 31656 2560
rect 32086 2560 32674 2576
rect 32086 2543 32102 2560
rect 31640 2526 31842 2543
rect 30882 2488 31842 2526
rect 31900 2526 32102 2543
rect 32658 2543 32674 2560
rect 33104 2560 33692 2576
rect 33104 2543 33120 2560
rect 32658 2526 32860 2543
rect 31900 2488 32860 2526
rect 32918 2526 33120 2543
rect 33676 2543 33692 2560
rect 33676 2526 33878 2543
rect 32918 2488 33878 2526
rect 1591 1897 2551 1935
rect 1591 1880 1793 1897
rect 1777 1863 1793 1880
rect 2349 1880 2551 1897
rect 2609 1897 3569 1935
rect 2609 1880 2811 1897
rect 2349 1863 2365 1880
rect 1777 1847 2365 1863
rect 2795 1863 2811 1880
rect 3367 1880 3569 1897
rect 3627 1897 4587 1935
rect 3627 1880 3829 1897
rect 3367 1863 3383 1880
rect 2795 1847 3383 1863
rect 3813 1863 3829 1880
rect 4385 1880 4587 1897
rect 4645 1897 5605 1935
rect 4645 1880 4847 1897
rect 4385 1863 4401 1880
rect 3813 1847 4401 1863
rect 4831 1863 4847 1880
rect 5403 1880 5605 1897
rect 5663 1897 6623 1935
rect 5663 1880 5865 1897
rect 5403 1863 5419 1880
rect 4831 1847 5419 1863
rect 5849 1863 5865 1880
rect 6421 1880 6623 1897
rect 6681 1897 7641 1935
rect 6681 1880 6883 1897
rect 6421 1863 6437 1880
rect 5849 1847 6437 1863
rect 6867 1863 6883 1880
rect 7439 1880 7641 1897
rect 8584 1898 8824 1936
rect 8584 1881 8642 1898
rect 7439 1863 7455 1880
rect 6867 1847 7455 1863
rect 8626 1864 8642 1881
rect 8766 1881 8824 1898
rect 8882 1898 9122 1936
rect 8882 1881 8940 1898
rect 8766 1864 8782 1881
rect 8626 1848 8782 1864
rect 8924 1864 8940 1881
rect 9064 1881 9122 1898
rect 9180 1898 9420 1936
rect 9180 1881 9238 1898
rect 9064 1864 9080 1881
rect 8924 1848 9080 1864
rect 9222 1864 9238 1881
rect 9362 1881 9420 1898
rect 9478 1898 9718 1936
rect 9478 1881 9536 1898
rect 9362 1864 9378 1881
rect 9222 1848 9378 1864
rect 9520 1864 9536 1881
rect 9660 1881 9718 1898
rect 9776 1898 10016 1936
rect 9776 1881 9834 1898
rect 9660 1864 9676 1881
rect 9520 1848 9676 1864
rect 9818 1864 9834 1881
rect 9958 1881 10016 1898
rect 10074 1898 10314 1936
rect 10074 1881 10132 1898
rect 9958 1864 9974 1881
rect 9818 1848 9974 1864
rect 10116 1864 10132 1881
rect 10256 1881 10314 1898
rect 10372 1898 10612 1936
rect 10372 1881 10430 1898
rect 10256 1864 10272 1881
rect 10116 1848 10272 1864
rect 10414 1864 10430 1881
rect 10554 1881 10612 1898
rect 10670 1898 10910 1936
rect 10670 1881 10728 1898
rect 10554 1864 10570 1881
rect 10414 1848 10570 1864
rect 10712 1864 10728 1881
rect 10852 1881 10910 1898
rect 10968 1898 11208 1936
rect 10968 1881 11026 1898
rect 10852 1864 10868 1881
rect 10712 1848 10868 1864
rect 11010 1864 11026 1881
rect 11150 1881 11208 1898
rect 11266 1898 11506 1936
rect 11266 1881 11324 1898
rect 11150 1864 11166 1881
rect 11010 1848 11166 1864
rect 11308 1864 11324 1881
rect 11448 1881 11506 1898
rect 11564 1898 11804 1936
rect 11564 1881 11622 1898
rect 11448 1864 11464 1881
rect 11308 1848 11464 1864
rect 11606 1864 11622 1881
rect 11746 1881 11804 1898
rect 11746 1864 11762 1881
rect 11606 1848 11762 1864
rect 13576 1850 14536 1888
rect 13576 1833 13778 1850
rect 13762 1816 13778 1833
rect 14334 1833 14536 1850
rect 14594 1850 15554 1888
rect 14594 1833 14796 1850
rect 14334 1816 14350 1833
rect 13762 1800 14350 1816
rect 14780 1816 14796 1833
rect 15352 1833 15554 1850
rect 15612 1850 16572 1888
rect 15612 1833 15814 1850
rect 15352 1816 15368 1833
rect 14780 1800 15368 1816
rect 15798 1816 15814 1833
rect 16370 1833 16572 1850
rect 16630 1850 17590 1888
rect 16630 1833 16832 1850
rect 16370 1816 16386 1833
rect 15798 1800 16386 1816
rect 16816 1816 16832 1833
rect 17388 1833 17590 1850
rect 17648 1850 18608 1888
rect 17648 1833 17850 1850
rect 17388 1816 17404 1833
rect 16816 1800 17404 1816
rect 17834 1816 17850 1833
rect 18406 1833 18608 1850
rect 18666 1850 19626 1888
rect 18666 1833 18868 1850
rect 18406 1816 18422 1833
rect 17834 1800 18422 1816
rect 18852 1816 18868 1833
rect 19424 1833 19626 1850
rect 19684 1850 20644 1888
rect 19684 1833 19886 1850
rect 19424 1816 19440 1833
rect 18852 1800 19440 1816
rect 19870 1816 19886 1833
rect 20442 1833 20644 1850
rect 20702 1850 21662 1888
rect 20702 1833 20904 1850
rect 20442 1816 20458 1833
rect 19870 1800 20458 1816
rect 20888 1816 20904 1833
rect 21460 1833 21662 1850
rect 21720 1850 22680 1888
rect 21720 1833 21922 1850
rect 21460 1816 21476 1833
rect 20888 1800 21476 1816
rect 21906 1816 21922 1833
rect 22478 1833 22680 1850
rect 22738 1850 23698 1888
rect 22738 1833 22940 1850
rect 22478 1816 22494 1833
rect 21906 1800 22494 1816
rect 22924 1816 22940 1833
rect 23496 1833 23698 1850
rect 23756 1850 24716 1888
rect 23756 1833 23958 1850
rect 23496 1816 23512 1833
rect 22924 1800 23512 1816
rect 23942 1816 23958 1833
rect 24514 1833 24716 1850
rect 24774 1850 25734 1888
rect 24774 1833 24976 1850
rect 24514 1816 24530 1833
rect 23942 1800 24530 1816
rect 24960 1816 24976 1833
rect 25532 1833 25734 1850
rect 25792 1850 26752 1888
rect 25792 1833 25994 1850
rect 25532 1816 25548 1833
rect 24960 1800 25548 1816
rect 25978 1816 25994 1833
rect 26550 1833 26752 1850
rect 26810 1850 27770 1888
rect 26810 1833 27012 1850
rect 26550 1816 26566 1833
rect 25978 1800 26566 1816
rect 26996 1816 27012 1833
rect 27568 1833 27770 1850
rect 27828 1850 28788 1888
rect 27828 1833 28030 1850
rect 27568 1816 27584 1833
rect 26996 1800 27584 1816
rect 28014 1816 28030 1833
rect 28586 1833 28788 1850
rect 28846 1850 29806 1888
rect 28846 1833 29048 1850
rect 28586 1816 28602 1833
rect 28014 1800 28602 1816
rect 29032 1816 29048 1833
rect 29604 1833 29806 1850
rect 29864 1850 30824 1888
rect 29864 1833 30066 1850
rect 29604 1816 29620 1833
rect 29032 1800 29620 1816
rect 30050 1816 30066 1833
rect 30622 1833 30824 1850
rect 30882 1850 31842 1888
rect 30882 1833 31084 1850
rect 30622 1816 30638 1833
rect 30050 1800 30638 1816
rect 31068 1816 31084 1833
rect 31640 1833 31842 1850
rect 31900 1850 32860 1888
rect 31900 1833 32102 1850
rect 31640 1816 31656 1833
rect 31068 1800 31656 1816
rect 32086 1816 32102 1833
rect 32658 1833 32860 1850
rect 32918 1850 33878 1888
rect 32918 1833 33120 1850
rect 32658 1816 32674 1833
rect 32086 1800 32674 1816
rect 33104 1816 33120 1833
rect 33676 1833 33878 1850
rect 33676 1816 33692 1833
rect 33104 1800 33692 1816
rect 1776 1494 2364 1510
rect 1776 1477 1792 1494
rect 1590 1460 1792 1477
rect 2348 1477 2364 1494
rect 2794 1494 3382 1510
rect 2794 1477 2810 1494
rect 2348 1460 2550 1477
rect 1590 1422 2550 1460
rect 2608 1460 2810 1477
rect 3366 1477 3382 1494
rect 3812 1494 4400 1510
rect 3812 1477 3828 1494
rect 3366 1460 3568 1477
rect 2608 1422 3568 1460
rect 3626 1460 3828 1477
rect 4384 1477 4400 1494
rect 4830 1494 5418 1510
rect 4830 1477 4846 1494
rect 4384 1460 4586 1477
rect 3626 1422 4586 1460
rect 4644 1460 4846 1477
rect 5402 1477 5418 1494
rect 5848 1494 6436 1510
rect 5848 1477 5864 1494
rect 5402 1460 5604 1477
rect 4644 1422 5604 1460
rect 5662 1460 5864 1477
rect 6420 1477 6436 1494
rect 6866 1494 7454 1510
rect 6866 1477 6882 1494
rect 6420 1460 6622 1477
rect 5662 1422 6622 1460
rect 6680 1460 6882 1477
rect 7438 1477 7454 1494
rect 8626 1498 8782 1514
rect 8626 1481 8642 1498
rect 7438 1460 7640 1477
rect 6680 1422 7640 1460
rect 8584 1464 8642 1481
rect 8766 1481 8782 1498
rect 8924 1498 9080 1514
rect 8924 1481 8940 1498
rect 8766 1464 8824 1481
rect 8584 1426 8824 1464
rect 8882 1464 8940 1481
rect 9064 1481 9080 1498
rect 9222 1498 9378 1514
rect 9222 1481 9238 1498
rect 9064 1464 9122 1481
rect 8882 1426 9122 1464
rect 9180 1464 9238 1481
rect 9362 1481 9378 1498
rect 9520 1498 9676 1514
rect 9520 1481 9536 1498
rect 9362 1464 9420 1481
rect 9180 1426 9420 1464
rect 9478 1464 9536 1481
rect 9660 1481 9676 1498
rect 9818 1498 9974 1514
rect 9818 1481 9834 1498
rect 9660 1464 9718 1481
rect 9478 1426 9718 1464
rect 9776 1464 9834 1481
rect 9958 1481 9974 1498
rect 10116 1498 10272 1514
rect 10116 1481 10132 1498
rect 9958 1464 10016 1481
rect 9776 1426 10016 1464
rect 10074 1464 10132 1481
rect 10256 1481 10272 1498
rect 10414 1498 10570 1514
rect 10414 1481 10430 1498
rect 10256 1464 10314 1481
rect 10074 1426 10314 1464
rect 10372 1464 10430 1481
rect 10554 1481 10570 1498
rect 10712 1498 10868 1514
rect 10712 1481 10728 1498
rect 10554 1464 10612 1481
rect 10372 1426 10612 1464
rect 10670 1464 10728 1481
rect 10852 1481 10868 1498
rect 11010 1498 11166 1514
rect 11010 1481 11026 1498
rect 10852 1464 10910 1481
rect 10670 1426 10910 1464
rect 10968 1464 11026 1481
rect 11150 1481 11166 1498
rect 11308 1498 11464 1514
rect 11308 1481 11324 1498
rect 11150 1464 11208 1481
rect 10968 1426 11208 1464
rect 11266 1464 11324 1481
rect 11448 1481 11464 1498
rect 11606 1498 11762 1514
rect 11606 1481 11622 1498
rect 11448 1464 11506 1481
rect 11266 1426 11506 1464
rect 11564 1464 11622 1481
rect 11746 1481 11762 1498
rect 11746 1464 11804 1481
rect 11564 1426 11804 1464
rect 13762 1328 14350 1344
rect 13762 1311 13778 1328
rect 13576 1294 13778 1311
rect 14334 1311 14350 1328
rect 14780 1328 15368 1344
rect 14780 1311 14796 1328
rect 14334 1294 14536 1311
rect 13576 1256 14536 1294
rect 14594 1294 14796 1311
rect 15352 1311 15368 1328
rect 15798 1328 16386 1344
rect 15798 1311 15814 1328
rect 15352 1294 15554 1311
rect 14594 1256 15554 1294
rect 15612 1294 15814 1311
rect 16370 1311 16386 1328
rect 16816 1328 17404 1344
rect 16816 1311 16832 1328
rect 16370 1294 16572 1311
rect 15612 1256 16572 1294
rect 16630 1294 16832 1311
rect 17388 1311 17404 1328
rect 17834 1328 18422 1344
rect 17834 1311 17850 1328
rect 17388 1294 17590 1311
rect 16630 1256 17590 1294
rect 17648 1294 17850 1311
rect 18406 1311 18422 1328
rect 18852 1328 19440 1344
rect 18852 1311 18868 1328
rect 18406 1294 18608 1311
rect 17648 1256 18608 1294
rect 18666 1294 18868 1311
rect 19424 1311 19440 1328
rect 19870 1328 20458 1344
rect 19870 1311 19886 1328
rect 19424 1294 19626 1311
rect 18666 1256 19626 1294
rect 19684 1294 19886 1311
rect 20442 1311 20458 1328
rect 20888 1328 21476 1344
rect 20888 1311 20904 1328
rect 20442 1294 20644 1311
rect 19684 1256 20644 1294
rect 20702 1294 20904 1311
rect 21460 1311 21476 1328
rect 21906 1328 22494 1344
rect 21906 1311 21922 1328
rect 21460 1294 21662 1311
rect 20702 1256 21662 1294
rect 21720 1294 21922 1311
rect 22478 1311 22494 1328
rect 22924 1328 23512 1344
rect 22924 1311 22940 1328
rect 22478 1294 22680 1311
rect 21720 1256 22680 1294
rect 22738 1294 22940 1311
rect 23496 1311 23512 1328
rect 23942 1328 24530 1344
rect 23942 1311 23958 1328
rect 23496 1294 23698 1311
rect 22738 1256 23698 1294
rect 23756 1294 23958 1311
rect 24514 1311 24530 1328
rect 24960 1328 25548 1344
rect 24960 1311 24976 1328
rect 24514 1294 24716 1311
rect 23756 1256 24716 1294
rect 24774 1294 24976 1311
rect 25532 1311 25548 1328
rect 25978 1328 26566 1344
rect 25978 1311 25994 1328
rect 25532 1294 25734 1311
rect 24774 1256 25734 1294
rect 25792 1294 25994 1311
rect 26550 1311 26566 1328
rect 26996 1328 27584 1344
rect 26996 1311 27012 1328
rect 26550 1294 26752 1311
rect 25792 1256 26752 1294
rect 26810 1294 27012 1311
rect 27568 1311 27584 1328
rect 28014 1328 28602 1344
rect 28014 1311 28030 1328
rect 27568 1294 27770 1311
rect 26810 1256 27770 1294
rect 27828 1294 28030 1311
rect 28586 1311 28602 1328
rect 29032 1328 29620 1344
rect 29032 1311 29048 1328
rect 28586 1294 28788 1311
rect 27828 1256 28788 1294
rect 28846 1294 29048 1311
rect 29604 1311 29620 1328
rect 30050 1328 30638 1344
rect 30050 1311 30066 1328
rect 29604 1294 29806 1311
rect 28846 1256 29806 1294
rect 29864 1294 30066 1311
rect 30622 1311 30638 1328
rect 31068 1328 31656 1344
rect 31068 1311 31084 1328
rect 30622 1294 30824 1311
rect 29864 1256 30824 1294
rect 30882 1294 31084 1311
rect 31640 1311 31656 1328
rect 32086 1328 32674 1344
rect 32086 1311 32102 1328
rect 31640 1294 31842 1311
rect 30882 1256 31842 1294
rect 31900 1294 32102 1311
rect 32658 1311 32674 1328
rect 33104 1328 33692 1344
rect 33104 1311 33120 1328
rect 32658 1294 32860 1311
rect 31900 1256 32860 1294
rect 32918 1294 33120 1311
rect 33676 1311 33692 1328
rect 33676 1294 33878 1311
rect 32918 1256 33878 1294
rect 1590 784 2550 822
rect 1590 767 1792 784
rect 1776 750 1792 767
rect 2348 767 2550 784
rect 2608 784 3568 822
rect 2608 767 2810 784
rect 2348 750 2364 767
rect 1776 734 2364 750
rect 2794 750 2810 767
rect 3366 767 3568 784
rect 3626 784 4586 822
rect 3626 767 3828 784
rect 3366 750 3382 767
rect 2794 734 3382 750
rect 3812 750 3828 767
rect 4384 767 4586 784
rect 4644 784 5604 822
rect 4644 767 4846 784
rect 4384 750 4400 767
rect 3812 734 4400 750
rect 4830 750 4846 767
rect 5402 767 5604 784
rect 5662 784 6622 822
rect 5662 767 5864 784
rect 5402 750 5418 767
rect 4830 734 5418 750
rect 5848 750 5864 767
rect 6420 767 6622 784
rect 6680 784 7640 822
rect 6680 767 6882 784
rect 6420 750 6436 767
rect 5848 734 6436 750
rect 6866 750 6882 767
rect 7438 767 7640 784
rect 8584 788 8824 826
rect 8584 771 8642 788
rect 7438 750 7454 767
rect 6866 734 7454 750
rect 8626 754 8642 771
rect 8766 771 8824 788
rect 8882 788 9122 826
rect 8882 771 8940 788
rect 8766 754 8782 771
rect 8626 738 8782 754
rect 8924 754 8940 771
rect 9064 771 9122 788
rect 9180 788 9420 826
rect 9180 771 9238 788
rect 9064 754 9080 771
rect 8924 738 9080 754
rect 9222 754 9238 771
rect 9362 771 9420 788
rect 9478 788 9718 826
rect 9478 771 9536 788
rect 9362 754 9378 771
rect 9222 738 9378 754
rect 9520 754 9536 771
rect 9660 771 9718 788
rect 9776 788 10016 826
rect 9776 771 9834 788
rect 9660 754 9676 771
rect 9520 738 9676 754
rect 9818 754 9834 771
rect 9958 771 10016 788
rect 10074 788 10314 826
rect 10074 771 10132 788
rect 9958 754 9974 771
rect 9818 738 9974 754
rect 10116 754 10132 771
rect 10256 771 10314 788
rect 10372 788 10612 826
rect 10372 771 10430 788
rect 10256 754 10272 771
rect 10116 738 10272 754
rect 10414 754 10430 771
rect 10554 771 10612 788
rect 10670 788 10910 826
rect 10670 771 10728 788
rect 10554 754 10570 771
rect 10414 738 10570 754
rect 10712 754 10728 771
rect 10852 771 10910 788
rect 10968 788 11208 826
rect 10968 771 11026 788
rect 10852 754 10868 771
rect 10712 738 10868 754
rect 11010 754 11026 771
rect 11150 771 11208 788
rect 11266 788 11506 826
rect 11266 771 11324 788
rect 11150 754 11166 771
rect 11010 738 11166 754
rect 11308 754 11324 771
rect 11448 771 11506 788
rect 11564 788 11804 826
rect 11564 771 11622 788
rect 11448 754 11464 771
rect 11308 738 11464 754
rect 11606 754 11622 771
rect 11746 771 11804 788
rect 11746 754 11762 771
rect 11606 738 11762 754
rect 13576 618 14536 656
rect 13576 601 13778 618
rect 13762 584 13778 601
rect 14334 601 14536 618
rect 14594 618 15554 656
rect 14594 601 14796 618
rect 14334 584 14350 601
rect 13762 568 14350 584
rect 14780 584 14796 601
rect 15352 601 15554 618
rect 15612 618 16572 656
rect 15612 601 15814 618
rect 15352 584 15368 601
rect 14780 568 15368 584
rect 15798 584 15814 601
rect 16370 601 16572 618
rect 16630 618 17590 656
rect 16630 601 16832 618
rect 16370 584 16386 601
rect 15798 568 16386 584
rect 16816 584 16832 601
rect 17388 601 17590 618
rect 17648 618 18608 656
rect 17648 601 17850 618
rect 17388 584 17404 601
rect 16816 568 17404 584
rect 17834 584 17850 601
rect 18406 601 18608 618
rect 18666 618 19626 656
rect 18666 601 18868 618
rect 18406 584 18422 601
rect 17834 568 18422 584
rect 18852 584 18868 601
rect 19424 601 19626 618
rect 19684 618 20644 656
rect 19684 601 19886 618
rect 19424 584 19440 601
rect 18852 568 19440 584
rect 19870 584 19886 601
rect 20442 601 20644 618
rect 20702 618 21662 656
rect 20702 601 20904 618
rect 20442 584 20458 601
rect 19870 568 20458 584
rect 20888 584 20904 601
rect 21460 601 21662 618
rect 21720 618 22680 656
rect 21720 601 21922 618
rect 21460 584 21476 601
rect 20888 568 21476 584
rect 21906 584 21922 601
rect 22478 601 22680 618
rect 22738 618 23698 656
rect 22738 601 22940 618
rect 22478 584 22494 601
rect 21906 568 22494 584
rect 22924 584 22940 601
rect 23496 601 23698 618
rect 23756 618 24716 656
rect 23756 601 23958 618
rect 23496 584 23512 601
rect 22924 568 23512 584
rect 23942 584 23958 601
rect 24514 601 24716 618
rect 24774 618 25734 656
rect 24774 601 24976 618
rect 24514 584 24530 601
rect 23942 568 24530 584
rect 24960 584 24976 601
rect 25532 601 25734 618
rect 25792 618 26752 656
rect 25792 601 25994 618
rect 25532 584 25548 601
rect 24960 568 25548 584
rect 25978 584 25994 601
rect 26550 601 26752 618
rect 26810 618 27770 656
rect 26810 601 27012 618
rect 26550 584 26566 601
rect 25978 568 26566 584
rect 26996 584 27012 601
rect 27568 601 27770 618
rect 27828 618 28788 656
rect 27828 601 28030 618
rect 27568 584 27584 601
rect 26996 568 27584 584
rect 28014 584 28030 601
rect 28586 601 28788 618
rect 28846 618 29806 656
rect 28846 601 29048 618
rect 28586 584 28602 601
rect 28014 568 28602 584
rect 29032 584 29048 601
rect 29604 601 29806 618
rect 29864 618 30824 656
rect 29864 601 30066 618
rect 29604 584 29620 601
rect 29032 568 29620 584
rect 30050 584 30066 601
rect 30622 601 30824 618
rect 30882 618 31842 656
rect 30882 601 31084 618
rect 30622 584 30638 601
rect 30050 568 30638 584
rect 31068 584 31084 601
rect 31640 601 31842 618
rect 31900 618 32860 656
rect 31900 601 32102 618
rect 31640 584 31656 601
rect 31068 568 31656 584
rect 32086 584 32102 601
rect 32658 601 32860 618
rect 32918 618 33878 656
rect 32918 601 33120 618
rect 32658 584 32674 601
rect 32086 568 32674 584
rect 33104 584 33120 601
rect 33676 601 33878 618
rect 33676 584 33692 601
rect 33104 568 33692 584
rect 48884 8345 49016 8361
rect 48884 8328 48900 8345
rect 48850 8311 48900 8328
rect 49000 8328 49016 8345
rect 49142 8345 49274 8361
rect 49142 8328 49158 8345
rect 49000 8311 49050 8328
rect 48850 8264 49050 8311
rect 49108 8311 49158 8328
rect 49258 8328 49274 8345
rect 49400 8345 49532 8361
rect 49400 8328 49416 8345
rect 49258 8311 49308 8328
rect 49108 8264 49308 8311
rect 49366 8311 49416 8328
rect 49516 8328 49532 8345
rect 49658 8345 49790 8361
rect 49658 8328 49674 8345
rect 49516 8311 49566 8328
rect 49366 8264 49566 8311
rect 49624 8311 49674 8328
rect 49774 8328 49790 8345
rect 49916 8345 50048 8361
rect 49916 8328 49932 8345
rect 49774 8311 49824 8328
rect 49624 8264 49824 8311
rect 49882 8311 49932 8328
rect 50032 8328 50048 8345
rect 50174 8345 50306 8361
rect 50174 8328 50190 8345
rect 50032 8311 50082 8328
rect 49882 8264 50082 8311
rect 50140 8311 50190 8328
rect 50290 8328 50306 8345
rect 50290 8311 50340 8328
rect 50140 8264 50340 8311
rect 48850 7817 49050 7864
rect 48850 7800 48900 7817
rect 48884 7783 48900 7800
rect 49000 7800 49050 7817
rect 49108 7817 49308 7864
rect 49108 7800 49158 7817
rect 49000 7783 49016 7800
rect 48884 7767 49016 7783
rect 49142 7783 49158 7800
rect 49258 7800 49308 7817
rect 49366 7817 49566 7864
rect 49366 7800 49416 7817
rect 49258 7783 49274 7800
rect 49142 7767 49274 7783
rect 49400 7783 49416 7800
rect 49516 7800 49566 7817
rect 49624 7817 49824 7864
rect 49624 7800 49674 7817
rect 49516 7783 49532 7800
rect 49400 7767 49532 7783
rect 49658 7783 49674 7800
rect 49774 7800 49824 7817
rect 49882 7817 50082 7864
rect 49882 7800 49932 7817
rect 49774 7783 49790 7800
rect 49658 7767 49790 7783
rect 49916 7783 49932 7800
rect 50032 7800 50082 7817
rect 50140 7817 50340 7864
rect 50140 7800 50190 7817
rect 50032 7783 50048 7800
rect 49916 7767 50048 7783
rect 50174 7783 50190 7800
rect 50290 7800 50340 7817
rect 50290 7783 50306 7800
rect 50174 7767 50306 7783
rect 50700 7881 50730 7907
rect 50700 7649 50730 7681
rect 50700 7633 50786 7649
rect 50700 7599 50736 7633
rect 50770 7599 50786 7633
rect 50700 7583 50786 7599
rect 50700 7561 50730 7583
rect 48884 7412 49016 7428
rect 48884 7395 48900 7412
rect 48850 7378 48900 7395
rect 49000 7395 49016 7412
rect 49142 7412 49274 7428
rect 49142 7395 49158 7412
rect 49000 7378 49050 7395
rect 48850 7340 49050 7378
rect 49108 7378 49158 7395
rect 49258 7395 49274 7412
rect 49400 7412 49532 7428
rect 49400 7395 49416 7412
rect 49258 7378 49308 7395
rect 49108 7340 49308 7378
rect 49366 7378 49416 7395
rect 49516 7395 49532 7412
rect 49658 7412 49790 7428
rect 49658 7395 49674 7412
rect 49516 7378 49566 7395
rect 49366 7340 49566 7378
rect 49624 7378 49674 7395
rect 49774 7395 49790 7412
rect 49916 7412 50048 7428
rect 49916 7395 49932 7412
rect 49774 7378 49824 7395
rect 49624 7340 49824 7378
rect 49882 7378 49932 7395
rect 50032 7395 50048 7412
rect 50174 7412 50306 7428
rect 50174 7395 50190 7412
rect 50032 7378 50082 7395
rect 49882 7340 50082 7378
rect 50140 7378 50190 7395
rect 50290 7395 50306 7412
rect 50290 7378 50340 7395
rect 50140 7340 50340 7378
rect 48850 7102 49050 7140
rect 48850 7085 48900 7102
rect 48884 7068 48900 7085
rect 49000 7085 49050 7102
rect 49108 7102 49308 7140
rect 49108 7085 49158 7102
rect 49000 7068 49016 7085
rect 48884 7052 49016 7068
rect 49142 7068 49158 7085
rect 49258 7085 49308 7102
rect 49366 7102 49566 7140
rect 49366 7085 49416 7102
rect 49258 7068 49274 7085
rect 49142 7052 49274 7068
rect 49400 7068 49416 7085
rect 49516 7085 49566 7102
rect 49624 7102 49824 7140
rect 49624 7085 49674 7102
rect 49516 7068 49532 7085
rect 49400 7052 49532 7068
rect 49658 7068 49674 7085
rect 49774 7085 49824 7102
rect 49882 7102 50082 7140
rect 49882 7085 49932 7102
rect 49774 7068 49790 7085
rect 49658 7052 49790 7068
rect 49916 7068 49932 7085
rect 50032 7085 50082 7102
rect 50140 7102 50340 7140
rect 50140 7085 50190 7102
rect 50032 7068 50048 7085
rect 49916 7052 50048 7068
rect 50174 7068 50190 7085
rect 50290 7085 50340 7102
rect 50290 7068 50306 7085
rect 50174 7052 50306 7068
rect 50700 7405 50730 7431
rect 48884 6381 49016 6397
rect 48884 6364 48900 6381
rect 48850 6347 48900 6364
rect 49000 6364 49016 6381
rect 49142 6381 49274 6397
rect 49142 6364 49158 6381
rect 49000 6347 49050 6364
rect 48850 6300 49050 6347
rect 49108 6347 49158 6364
rect 49258 6364 49274 6381
rect 49400 6381 49532 6397
rect 49400 6364 49416 6381
rect 49258 6347 49308 6364
rect 49108 6300 49308 6347
rect 49366 6347 49416 6364
rect 49516 6364 49532 6381
rect 49658 6381 49790 6397
rect 49658 6364 49674 6381
rect 49516 6347 49566 6364
rect 49366 6300 49566 6347
rect 49624 6347 49674 6364
rect 49774 6364 49790 6381
rect 49916 6381 50048 6397
rect 49916 6364 49932 6381
rect 49774 6347 49824 6364
rect 49624 6300 49824 6347
rect 49882 6347 49932 6364
rect 50032 6364 50048 6381
rect 50174 6381 50306 6397
rect 50174 6364 50190 6381
rect 50032 6347 50082 6364
rect 49882 6300 50082 6347
rect 50140 6347 50190 6364
rect 50290 6364 50306 6381
rect 50290 6347 50340 6364
rect 50140 6300 50340 6347
rect 48850 5853 49050 5900
rect 48850 5836 48900 5853
rect 48884 5819 48900 5836
rect 49000 5836 49050 5853
rect 49108 5853 49308 5900
rect 49108 5836 49158 5853
rect 49000 5819 49016 5836
rect 48884 5803 49016 5819
rect 49142 5819 49158 5836
rect 49258 5836 49308 5853
rect 49366 5853 49566 5900
rect 49366 5836 49416 5853
rect 49258 5819 49274 5836
rect 49142 5803 49274 5819
rect 49400 5819 49416 5836
rect 49516 5836 49566 5853
rect 49624 5853 49824 5900
rect 49624 5836 49674 5853
rect 49516 5819 49532 5836
rect 49400 5803 49532 5819
rect 49658 5819 49674 5836
rect 49774 5836 49824 5853
rect 49882 5853 50082 5900
rect 49882 5836 49932 5853
rect 49774 5819 49790 5836
rect 49658 5803 49790 5819
rect 49916 5819 49932 5836
rect 50032 5836 50082 5853
rect 50140 5853 50340 5900
rect 50140 5836 50190 5853
rect 50032 5819 50048 5836
rect 49916 5803 50048 5819
rect 50174 5819 50190 5836
rect 50290 5836 50340 5853
rect 50290 5819 50306 5836
rect 50174 5803 50306 5819
rect 50700 5917 50730 5943
rect 50700 5685 50730 5717
rect 50700 5669 50786 5685
rect 50700 5635 50736 5669
rect 50770 5635 50786 5669
rect 50700 5619 50786 5635
rect 50700 5597 50730 5619
rect 48884 5448 49016 5464
rect 48884 5431 48900 5448
rect 48850 5414 48900 5431
rect 49000 5431 49016 5448
rect 49142 5448 49274 5464
rect 49142 5431 49158 5448
rect 49000 5414 49050 5431
rect 48850 5376 49050 5414
rect 49108 5414 49158 5431
rect 49258 5431 49274 5448
rect 49400 5448 49532 5464
rect 49400 5431 49416 5448
rect 49258 5414 49308 5431
rect 49108 5376 49308 5414
rect 49366 5414 49416 5431
rect 49516 5431 49532 5448
rect 49658 5448 49790 5464
rect 49658 5431 49674 5448
rect 49516 5414 49566 5431
rect 49366 5376 49566 5414
rect 49624 5414 49674 5431
rect 49774 5431 49790 5448
rect 49916 5448 50048 5464
rect 49916 5431 49932 5448
rect 49774 5414 49824 5431
rect 49624 5376 49824 5414
rect 49882 5414 49932 5431
rect 50032 5431 50048 5448
rect 50174 5448 50306 5464
rect 50174 5431 50190 5448
rect 50032 5414 50082 5431
rect 49882 5376 50082 5414
rect 50140 5414 50190 5431
rect 50290 5431 50306 5448
rect 50290 5414 50340 5431
rect 50140 5376 50340 5414
rect 48850 5138 49050 5176
rect 48850 5121 48900 5138
rect 48884 5104 48900 5121
rect 49000 5121 49050 5138
rect 49108 5138 49308 5176
rect 49108 5121 49158 5138
rect 49000 5104 49016 5121
rect 48884 5088 49016 5104
rect 49142 5104 49158 5121
rect 49258 5121 49308 5138
rect 49366 5138 49566 5176
rect 49366 5121 49416 5138
rect 49258 5104 49274 5121
rect 49142 5088 49274 5104
rect 49400 5104 49416 5121
rect 49516 5121 49566 5138
rect 49624 5138 49824 5176
rect 49624 5121 49674 5138
rect 49516 5104 49532 5121
rect 49400 5088 49532 5104
rect 49658 5104 49674 5121
rect 49774 5121 49824 5138
rect 49882 5138 50082 5176
rect 49882 5121 49932 5138
rect 49774 5104 49790 5121
rect 49658 5088 49790 5104
rect 49916 5104 49932 5121
rect 50032 5121 50082 5138
rect 50140 5138 50340 5176
rect 50140 5121 50190 5138
rect 50032 5104 50048 5121
rect 49916 5088 50048 5104
rect 50174 5104 50190 5121
rect 50290 5121 50340 5138
rect 50290 5104 50306 5121
rect 50174 5088 50306 5104
rect 50700 5441 50730 5467
rect 48884 4381 49016 4397
rect 48884 4364 48900 4381
rect 48850 4347 48900 4364
rect 49000 4364 49016 4381
rect 49142 4381 49274 4397
rect 49142 4364 49158 4381
rect 49000 4347 49050 4364
rect 48850 4300 49050 4347
rect 49108 4347 49158 4364
rect 49258 4364 49274 4381
rect 49400 4381 49532 4397
rect 49400 4364 49416 4381
rect 49258 4347 49308 4364
rect 49108 4300 49308 4347
rect 49366 4347 49416 4364
rect 49516 4364 49532 4381
rect 49658 4381 49790 4397
rect 49658 4364 49674 4381
rect 49516 4347 49566 4364
rect 49366 4300 49566 4347
rect 49624 4347 49674 4364
rect 49774 4364 49790 4381
rect 49916 4381 50048 4397
rect 49916 4364 49932 4381
rect 49774 4347 49824 4364
rect 49624 4300 49824 4347
rect 49882 4347 49932 4364
rect 50032 4364 50048 4381
rect 50174 4381 50306 4397
rect 50174 4364 50190 4381
rect 50032 4347 50082 4364
rect 49882 4300 50082 4347
rect 50140 4347 50190 4364
rect 50290 4364 50306 4381
rect 50290 4347 50340 4364
rect 50140 4300 50340 4347
rect 48850 3853 49050 3900
rect 48850 3836 48900 3853
rect 48884 3819 48900 3836
rect 49000 3836 49050 3853
rect 49108 3853 49308 3900
rect 49108 3836 49158 3853
rect 49000 3819 49016 3836
rect 48884 3803 49016 3819
rect 49142 3819 49158 3836
rect 49258 3836 49308 3853
rect 49366 3853 49566 3900
rect 49366 3836 49416 3853
rect 49258 3819 49274 3836
rect 49142 3803 49274 3819
rect 49400 3819 49416 3836
rect 49516 3836 49566 3853
rect 49624 3853 49824 3900
rect 49624 3836 49674 3853
rect 49516 3819 49532 3836
rect 49400 3803 49532 3819
rect 49658 3819 49674 3836
rect 49774 3836 49824 3853
rect 49882 3853 50082 3900
rect 49882 3836 49932 3853
rect 49774 3819 49790 3836
rect 49658 3803 49790 3819
rect 49916 3819 49932 3836
rect 50032 3836 50082 3853
rect 50140 3853 50340 3900
rect 50140 3836 50190 3853
rect 50032 3819 50048 3836
rect 49916 3803 50048 3819
rect 50174 3819 50190 3836
rect 50290 3836 50340 3853
rect 50290 3819 50306 3836
rect 50174 3803 50306 3819
rect 50700 3917 50730 3943
rect 50700 3685 50730 3717
rect 50700 3669 50786 3685
rect 50700 3635 50736 3669
rect 50770 3635 50786 3669
rect 50700 3619 50786 3635
rect 50700 3597 50730 3619
rect 48884 3448 49016 3464
rect 48884 3431 48900 3448
rect 48850 3414 48900 3431
rect 49000 3431 49016 3448
rect 49142 3448 49274 3464
rect 49142 3431 49158 3448
rect 49000 3414 49050 3431
rect 48850 3376 49050 3414
rect 49108 3414 49158 3431
rect 49258 3431 49274 3448
rect 49400 3448 49532 3464
rect 49400 3431 49416 3448
rect 49258 3414 49308 3431
rect 49108 3376 49308 3414
rect 49366 3414 49416 3431
rect 49516 3431 49532 3448
rect 49658 3448 49790 3464
rect 49658 3431 49674 3448
rect 49516 3414 49566 3431
rect 49366 3376 49566 3414
rect 49624 3414 49674 3431
rect 49774 3431 49790 3448
rect 49916 3448 50048 3464
rect 49916 3431 49932 3448
rect 49774 3414 49824 3431
rect 49624 3376 49824 3414
rect 49882 3414 49932 3431
rect 50032 3431 50048 3448
rect 50174 3448 50306 3464
rect 50174 3431 50190 3448
rect 50032 3414 50082 3431
rect 49882 3376 50082 3414
rect 50140 3414 50190 3431
rect 50290 3431 50306 3448
rect 50290 3414 50340 3431
rect 50140 3376 50340 3414
rect 48850 3138 49050 3176
rect 48850 3121 48900 3138
rect 48884 3104 48900 3121
rect 49000 3121 49050 3138
rect 49108 3138 49308 3176
rect 49108 3121 49158 3138
rect 49000 3104 49016 3121
rect 48884 3088 49016 3104
rect 49142 3104 49158 3121
rect 49258 3121 49308 3138
rect 49366 3138 49566 3176
rect 49366 3121 49416 3138
rect 49258 3104 49274 3121
rect 49142 3088 49274 3104
rect 49400 3104 49416 3121
rect 49516 3121 49566 3138
rect 49624 3138 49824 3176
rect 49624 3121 49674 3138
rect 49516 3104 49532 3121
rect 49400 3088 49532 3104
rect 49658 3104 49674 3121
rect 49774 3121 49824 3138
rect 49882 3138 50082 3176
rect 49882 3121 49932 3138
rect 49774 3104 49790 3121
rect 49658 3088 49790 3104
rect 49916 3104 49932 3121
rect 50032 3121 50082 3138
rect 50140 3138 50340 3176
rect 50140 3121 50190 3138
rect 50032 3104 50048 3121
rect 49916 3088 50048 3104
rect 50174 3104 50190 3121
rect 50290 3121 50340 3138
rect 50290 3104 50306 3121
rect 50174 3088 50306 3104
rect 50700 3441 50730 3467
rect 48884 2291 49016 2307
rect 48884 2274 48900 2291
rect 48850 2257 48900 2274
rect 49000 2274 49016 2291
rect 49142 2291 49274 2307
rect 49142 2274 49158 2291
rect 49000 2257 49050 2274
rect 48850 2210 49050 2257
rect 49108 2257 49158 2274
rect 49258 2274 49274 2291
rect 49400 2291 49532 2307
rect 49400 2274 49416 2291
rect 49258 2257 49308 2274
rect 49108 2210 49308 2257
rect 49366 2257 49416 2274
rect 49516 2274 49532 2291
rect 49658 2291 49790 2307
rect 49658 2274 49674 2291
rect 49516 2257 49566 2274
rect 49366 2210 49566 2257
rect 49624 2257 49674 2274
rect 49774 2274 49790 2291
rect 49916 2291 50048 2307
rect 49916 2274 49932 2291
rect 49774 2257 49824 2274
rect 49624 2210 49824 2257
rect 49882 2257 49932 2274
rect 50032 2274 50048 2291
rect 50174 2291 50306 2307
rect 50174 2274 50190 2291
rect 50032 2257 50082 2274
rect 49882 2210 50082 2257
rect 50140 2257 50190 2274
rect 50290 2274 50306 2291
rect 50290 2257 50340 2274
rect 50140 2210 50340 2257
rect 48850 1763 49050 1810
rect 48850 1746 48900 1763
rect 48884 1729 48900 1746
rect 49000 1746 49050 1763
rect 49108 1763 49308 1810
rect 49108 1746 49158 1763
rect 49000 1729 49016 1746
rect 48884 1713 49016 1729
rect 49142 1729 49158 1746
rect 49258 1746 49308 1763
rect 49366 1763 49566 1810
rect 49366 1746 49416 1763
rect 49258 1729 49274 1746
rect 49142 1713 49274 1729
rect 49400 1729 49416 1746
rect 49516 1746 49566 1763
rect 49624 1763 49824 1810
rect 49624 1746 49674 1763
rect 49516 1729 49532 1746
rect 49400 1713 49532 1729
rect 49658 1729 49674 1746
rect 49774 1746 49824 1763
rect 49882 1763 50082 1810
rect 49882 1746 49932 1763
rect 49774 1729 49790 1746
rect 49658 1713 49790 1729
rect 49916 1729 49932 1746
rect 50032 1746 50082 1763
rect 50140 1763 50340 1810
rect 50140 1746 50190 1763
rect 50032 1729 50048 1746
rect 49916 1713 50048 1729
rect 50174 1729 50190 1746
rect 50290 1746 50340 1763
rect 50290 1729 50306 1746
rect 50174 1713 50306 1729
rect 50700 1827 50730 1853
rect 50700 1595 50730 1627
rect 50700 1579 50786 1595
rect 50700 1545 50736 1579
rect 50770 1545 50786 1579
rect 50700 1529 50786 1545
rect 50700 1507 50730 1529
rect 48884 1358 49016 1374
rect 48884 1341 48900 1358
rect 48850 1324 48900 1341
rect 49000 1341 49016 1358
rect 49142 1358 49274 1374
rect 49142 1341 49158 1358
rect 49000 1324 49050 1341
rect 48850 1286 49050 1324
rect 49108 1324 49158 1341
rect 49258 1341 49274 1358
rect 49400 1358 49532 1374
rect 49400 1341 49416 1358
rect 49258 1324 49308 1341
rect 49108 1286 49308 1324
rect 49366 1324 49416 1341
rect 49516 1341 49532 1358
rect 49658 1358 49790 1374
rect 49658 1341 49674 1358
rect 49516 1324 49566 1341
rect 49366 1286 49566 1324
rect 49624 1324 49674 1341
rect 49774 1341 49790 1358
rect 49916 1358 50048 1374
rect 49916 1341 49932 1358
rect 49774 1324 49824 1341
rect 49624 1286 49824 1324
rect 49882 1324 49932 1341
rect 50032 1341 50048 1358
rect 50174 1358 50306 1374
rect 50174 1341 50190 1358
rect 50032 1324 50082 1341
rect 49882 1286 50082 1324
rect 50140 1324 50190 1341
rect 50290 1341 50306 1358
rect 50290 1324 50340 1341
rect 50140 1286 50340 1324
rect 48850 1048 49050 1086
rect 48850 1031 48900 1048
rect 48884 1014 48900 1031
rect 49000 1031 49050 1048
rect 49108 1048 49308 1086
rect 49108 1031 49158 1048
rect 49000 1014 49016 1031
rect 48884 998 49016 1014
rect 49142 1014 49158 1031
rect 49258 1031 49308 1048
rect 49366 1048 49566 1086
rect 49366 1031 49416 1048
rect 49258 1014 49274 1031
rect 49142 998 49274 1014
rect 49400 1014 49416 1031
rect 49516 1031 49566 1048
rect 49624 1048 49824 1086
rect 49624 1031 49674 1048
rect 49516 1014 49532 1031
rect 49400 998 49532 1014
rect 49658 1014 49674 1031
rect 49774 1031 49824 1048
rect 49882 1048 50082 1086
rect 49882 1031 49932 1048
rect 49774 1014 49790 1031
rect 49658 998 49790 1014
rect 49916 1014 49932 1031
rect 50032 1031 50082 1048
rect 50140 1048 50340 1086
rect 50140 1031 50190 1048
rect 50032 1014 50048 1031
rect 49916 998 50048 1014
rect 50174 1014 50190 1031
rect 50290 1031 50340 1048
rect 50290 1014 50306 1031
rect 50174 998 50306 1014
rect 50700 1351 50730 1377
rect 67764 14894 68352 14910
rect 67764 14877 67780 14894
rect 67578 14860 67780 14877
rect 68336 14877 68352 14894
rect 68782 14894 69370 14910
rect 68782 14877 68798 14894
rect 68336 14860 68538 14877
rect 67578 14822 68538 14860
rect 68596 14860 68798 14877
rect 69354 14877 69370 14894
rect 69800 14894 70388 14910
rect 69800 14877 69816 14894
rect 69354 14860 69556 14877
rect 68596 14822 69556 14860
rect 69614 14860 69816 14877
rect 70372 14877 70388 14894
rect 70818 14894 71406 14910
rect 70818 14877 70834 14894
rect 70372 14860 70574 14877
rect 69614 14822 70574 14860
rect 70632 14860 70834 14877
rect 71390 14877 71406 14894
rect 71836 14894 72424 14910
rect 71836 14877 71852 14894
rect 71390 14860 71592 14877
rect 70632 14822 71592 14860
rect 71650 14860 71852 14877
rect 72408 14877 72424 14894
rect 72854 14894 73442 14910
rect 72854 14877 72870 14894
rect 72408 14860 72610 14877
rect 71650 14822 72610 14860
rect 72668 14860 72870 14877
rect 73426 14877 73442 14894
rect 73872 14894 74460 14910
rect 73872 14877 73888 14894
rect 73426 14860 73628 14877
rect 72668 14822 73628 14860
rect 73686 14860 73888 14877
rect 74444 14877 74460 14894
rect 74890 14894 75478 14910
rect 74890 14877 74906 14894
rect 74444 14860 74646 14877
rect 73686 14822 74646 14860
rect 74704 14860 74906 14877
rect 75462 14877 75478 14894
rect 75908 14894 76496 14910
rect 75908 14877 75924 14894
rect 75462 14860 75664 14877
rect 74704 14822 75664 14860
rect 75722 14860 75924 14877
rect 76480 14877 76496 14894
rect 76926 14894 77514 14910
rect 76926 14877 76942 14894
rect 76480 14860 76682 14877
rect 75722 14822 76682 14860
rect 76740 14860 76942 14877
rect 77498 14877 77514 14894
rect 77944 14894 78532 14910
rect 77944 14877 77960 14894
rect 77498 14860 77700 14877
rect 76740 14822 77700 14860
rect 77758 14860 77960 14877
rect 78516 14877 78532 14894
rect 78962 14894 79550 14910
rect 78962 14877 78978 14894
rect 78516 14860 78718 14877
rect 77758 14822 78718 14860
rect 78776 14860 78978 14877
rect 79534 14877 79550 14894
rect 79980 14894 80568 14910
rect 79980 14877 79996 14894
rect 79534 14860 79736 14877
rect 78776 14822 79736 14860
rect 79794 14860 79996 14877
rect 80552 14877 80568 14894
rect 80998 14894 81586 14910
rect 80998 14877 81014 14894
rect 80552 14860 80754 14877
rect 79794 14822 80754 14860
rect 80812 14860 81014 14877
rect 81570 14877 81586 14894
rect 82016 14894 82604 14910
rect 82016 14877 82032 14894
rect 81570 14860 81772 14877
rect 80812 14822 81772 14860
rect 81830 14860 82032 14877
rect 82588 14877 82604 14894
rect 83034 14894 83622 14910
rect 83034 14877 83050 14894
rect 82588 14860 82790 14877
rect 81830 14822 82790 14860
rect 82848 14860 83050 14877
rect 83606 14877 83622 14894
rect 84052 14894 84640 14910
rect 84052 14877 84068 14894
rect 83606 14860 83808 14877
rect 82848 14822 83808 14860
rect 83866 14860 84068 14877
rect 84624 14877 84640 14894
rect 85070 14894 85658 14910
rect 85070 14877 85086 14894
rect 84624 14860 84826 14877
rect 83866 14822 84826 14860
rect 84884 14860 85086 14877
rect 85642 14877 85658 14894
rect 86088 14894 86676 14910
rect 86088 14877 86104 14894
rect 85642 14860 85844 14877
rect 84884 14822 85844 14860
rect 85902 14860 86104 14877
rect 86660 14877 86676 14894
rect 87106 14894 87694 14910
rect 87106 14877 87122 14894
rect 86660 14860 86862 14877
rect 85902 14822 86862 14860
rect 86920 14860 87122 14877
rect 87678 14877 87694 14894
rect 87678 14860 87880 14877
rect 86920 14822 87880 14860
rect 67578 14184 68538 14222
rect 67578 14167 67780 14184
rect 67764 14150 67780 14167
rect 68336 14167 68538 14184
rect 68596 14184 69556 14222
rect 68596 14167 68798 14184
rect 68336 14150 68352 14167
rect 67764 14134 68352 14150
rect 68782 14150 68798 14167
rect 69354 14167 69556 14184
rect 69614 14184 70574 14222
rect 69614 14167 69816 14184
rect 69354 14150 69370 14167
rect 68782 14134 69370 14150
rect 69800 14150 69816 14167
rect 70372 14167 70574 14184
rect 70632 14184 71592 14222
rect 70632 14167 70834 14184
rect 70372 14150 70388 14167
rect 69800 14134 70388 14150
rect 70818 14150 70834 14167
rect 71390 14167 71592 14184
rect 71650 14184 72610 14222
rect 71650 14167 71852 14184
rect 71390 14150 71406 14167
rect 70818 14134 71406 14150
rect 71836 14150 71852 14167
rect 72408 14167 72610 14184
rect 72668 14184 73628 14222
rect 72668 14167 72870 14184
rect 72408 14150 72424 14167
rect 71836 14134 72424 14150
rect 72854 14150 72870 14167
rect 73426 14167 73628 14184
rect 73686 14184 74646 14222
rect 73686 14167 73888 14184
rect 73426 14150 73442 14167
rect 72854 14134 73442 14150
rect 73872 14150 73888 14167
rect 74444 14167 74646 14184
rect 74704 14184 75664 14222
rect 74704 14167 74906 14184
rect 74444 14150 74460 14167
rect 73872 14134 74460 14150
rect 74890 14150 74906 14167
rect 75462 14167 75664 14184
rect 75722 14184 76682 14222
rect 75722 14167 75924 14184
rect 75462 14150 75478 14167
rect 74890 14134 75478 14150
rect 75908 14150 75924 14167
rect 76480 14167 76682 14184
rect 76740 14184 77700 14222
rect 76740 14167 76942 14184
rect 76480 14150 76496 14167
rect 75908 14134 76496 14150
rect 76926 14150 76942 14167
rect 77498 14167 77700 14184
rect 77758 14184 78718 14222
rect 77758 14167 77960 14184
rect 77498 14150 77514 14167
rect 76926 14134 77514 14150
rect 77944 14150 77960 14167
rect 78516 14167 78718 14184
rect 78776 14184 79736 14222
rect 78776 14167 78978 14184
rect 78516 14150 78532 14167
rect 77944 14134 78532 14150
rect 78962 14150 78978 14167
rect 79534 14167 79736 14184
rect 79794 14184 80754 14222
rect 79794 14167 79996 14184
rect 79534 14150 79550 14167
rect 78962 14134 79550 14150
rect 79980 14150 79996 14167
rect 80552 14167 80754 14184
rect 80812 14184 81772 14222
rect 80812 14167 81014 14184
rect 80552 14150 80568 14167
rect 79980 14134 80568 14150
rect 80998 14150 81014 14167
rect 81570 14167 81772 14184
rect 81830 14184 82790 14222
rect 81830 14167 82032 14184
rect 81570 14150 81586 14167
rect 80998 14134 81586 14150
rect 82016 14150 82032 14167
rect 82588 14167 82790 14184
rect 82848 14184 83808 14222
rect 82848 14167 83050 14184
rect 82588 14150 82604 14167
rect 82016 14134 82604 14150
rect 83034 14150 83050 14167
rect 83606 14167 83808 14184
rect 83866 14184 84826 14222
rect 83866 14167 84068 14184
rect 83606 14150 83622 14167
rect 83034 14134 83622 14150
rect 84052 14150 84068 14167
rect 84624 14167 84826 14184
rect 84884 14184 85844 14222
rect 84884 14167 85086 14184
rect 84624 14150 84640 14167
rect 84052 14134 84640 14150
rect 85070 14150 85086 14167
rect 85642 14167 85844 14184
rect 85902 14184 86862 14222
rect 85902 14167 86104 14184
rect 85642 14150 85658 14167
rect 85070 14134 85658 14150
rect 86088 14150 86104 14167
rect 86660 14167 86862 14184
rect 86920 14184 87880 14222
rect 86920 14167 87122 14184
rect 86660 14150 86676 14167
rect 86088 14134 86676 14150
rect 87106 14150 87122 14167
rect 87678 14167 87880 14184
rect 87678 14150 87694 14167
rect 87106 14134 87694 14150
rect 55998 14100 56586 14116
rect 55998 14083 56014 14100
rect 55812 14066 56014 14083
rect 56570 14083 56586 14100
rect 57016 14100 57604 14116
rect 57016 14083 57032 14100
rect 56570 14066 56772 14083
rect 55812 14028 56772 14066
rect 56830 14066 57032 14083
rect 57588 14083 57604 14100
rect 58034 14100 58622 14116
rect 58034 14083 58050 14100
rect 57588 14066 57790 14083
rect 56830 14028 57790 14066
rect 57848 14066 58050 14083
rect 58606 14083 58622 14100
rect 59052 14100 59640 14116
rect 59052 14083 59068 14100
rect 58606 14066 58808 14083
rect 57848 14028 58808 14066
rect 58866 14066 59068 14083
rect 59624 14083 59640 14100
rect 60070 14100 60658 14116
rect 60070 14083 60086 14100
rect 59624 14066 59826 14083
rect 58866 14028 59826 14066
rect 59884 14066 60086 14083
rect 60642 14083 60658 14100
rect 61088 14100 61676 14116
rect 61088 14083 61104 14100
rect 60642 14066 60844 14083
rect 59884 14028 60844 14066
rect 60902 14066 61104 14083
rect 61660 14083 61676 14100
rect 62106 14100 62694 14116
rect 62106 14083 62122 14100
rect 61660 14066 61862 14083
rect 60902 14028 61862 14066
rect 61920 14066 62122 14083
rect 62678 14083 62694 14100
rect 63124 14100 63712 14116
rect 63124 14083 63140 14100
rect 62678 14066 62880 14083
rect 61920 14028 62880 14066
rect 62938 14066 63140 14083
rect 63696 14083 63712 14100
rect 64142 14100 64730 14116
rect 64142 14083 64158 14100
rect 63696 14066 63898 14083
rect 62938 14028 63898 14066
rect 63956 14066 64158 14083
rect 64714 14083 64730 14100
rect 64714 14066 64916 14083
rect 63956 14028 64916 14066
rect 67764 13660 68352 13676
rect 67764 13643 67780 13660
rect 67578 13626 67780 13643
rect 68336 13643 68352 13660
rect 68782 13660 69370 13676
rect 68782 13643 68798 13660
rect 68336 13626 68538 13643
rect 67578 13588 68538 13626
rect 68596 13626 68798 13643
rect 69354 13643 69370 13660
rect 69800 13660 70388 13676
rect 69800 13643 69816 13660
rect 69354 13626 69556 13643
rect 68596 13588 69556 13626
rect 69614 13626 69816 13643
rect 70372 13643 70388 13660
rect 70818 13660 71406 13676
rect 70818 13643 70834 13660
rect 70372 13626 70574 13643
rect 69614 13588 70574 13626
rect 70632 13626 70834 13643
rect 71390 13643 71406 13660
rect 71836 13660 72424 13676
rect 71836 13643 71852 13660
rect 71390 13626 71592 13643
rect 70632 13588 71592 13626
rect 71650 13626 71852 13643
rect 72408 13643 72424 13660
rect 72854 13660 73442 13676
rect 72854 13643 72870 13660
rect 72408 13626 72610 13643
rect 71650 13588 72610 13626
rect 72668 13626 72870 13643
rect 73426 13643 73442 13660
rect 73872 13660 74460 13676
rect 73872 13643 73888 13660
rect 73426 13626 73628 13643
rect 72668 13588 73628 13626
rect 73686 13626 73888 13643
rect 74444 13643 74460 13660
rect 74890 13660 75478 13676
rect 74890 13643 74906 13660
rect 74444 13626 74646 13643
rect 73686 13588 74646 13626
rect 74704 13626 74906 13643
rect 75462 13643 75478 13660
rect 75908 13660 76496 13676
rect 75908 13643 75924 13660
rect 75462 13626 75664 13643
rect 74704 13588 75664 13626
rect 75722 13626 75924 13643
rect 76480 13643 76496 13660
rect 76926 13660 77514 13676
rect 76926 13643 76942 13660
rect 76480 13626 76682 13643
rect 75722 13588 76682 13626
rect 76740 13626 76942 13643
rect 77498 13643 77514 13660
rect 77944 13660 78532 13676
rect 77944 13643 77960 13660
rect 77498 13626 77700 13643
rect 76740 13588 77700 13626
rect 77758 13626 77960 13643
rect 78516 13643 78532 13660
rect 78962 13660 79550 13676
rect 78962 13643 78978 13660
rect 78516 13626 78718 13643
rect 77758 13588 78718 13626
rect 78776 13626 78978 13643
rect 79534 13643 79550 13660
rect 79980 13660 80568 13676
rect 79980 13643 79996 13660
rect 79534 13626 79736 13643
rect 78776 13588 79736 13626
rect 79794 13626 79996 13643
rect 80552 13643 80568 13660
rect 80998 13660 81586 13676
rect 80998 13643 81014 13660
rect 80552 13626 80754 13643
rect 79794 13588 80754 13626
rect 80812 13626 81014 13643
rect 81570 13643 81586 13660
rect 82016 13660 82604 13676
rect 82016 13643 82032 13660
rect 81570 13626 81772 13643
rect 80812 13588 81772 13626
rect 81830 13626 82032 13643
rect 82588 13643 82604 13660
rect 83034 13660 83622 13676
rect 83034 13643 83050 13660
rect 82588 13626 82790 13643
rect 81830 13588 82790 13626
rect 82848 13626 83050 13643
rect 83606 13643 83622 13660
rect 84052 13660 84640 13676
rect 84052 13643 84068 13660
rect 83606 13626 83808 13643
rect 82848 13588 83808 13626
rect 83866 13626 84068 13643
rect 84624 13643 84640 13660
rect 85070 13660 85658 13676
rect 85070 13643 85086 13660
rect 84624 13626 84826 13643
rect 83866 13588 84826 13626
rect 84884 13626 85086 13643
rect 85642 13643 85658 13660
rect 86088 13660 86676 13676
rect 86088 13643 86104 13660
rect 85642 13626 85844 13643
rect 84884 13588 85844 13626
rect 85902 13626 86104 13643
rect 86660 13643 86676 13660
rect 87106 13660 87694 13676
rect 87106 13643 87122 13660
rect 86660 13626 86862 13643
rect 85902 13588 86862 13626
rect 86920 13626 87122 13643
rect 87678 13643 87694 13660
rect 87678 13626 87880 13643
rect 86920 13588 87880 13626
rect 55812 13390 56772 13428
rect 55812 13373 56014 13390
rect 55998 13356 56014 13373
rect 56570 13373 56772 13390
rect 56830 13390 57790 13428
rect 56830 13373 57032 13390
rect 56570 13356 56586 13373
rect 55998 13340 56586 13356
rect 57016 13356 57032 13373
rect 57588 13373 57790 13390
rect 57848 13390 58808 13428
rect 57848 13373 58050 13390
rect 57588 13356 57604 13373
rect 57016 13340 57604 13356
rect 55998 13282 56586 13298
rect 55998 13265 56014 13282
rect 55812 13248 56014 13265
rect 56570 13265 56586 13282
rect 58034 13356 58050 13373
rect 58606 13373 58808 13390
rect 58866 13390 59826 13428
rect 58866 13373 59068 13390
rect 58606 13356 58622 13373
rect 58034 13340 58622 13356
rect 57016 13282 57604 13298
rect 57016 13265 57032 13282
rect 56570 13248 56772 13265
rect 55812 13210 56772 13248
rect 56830 13248 57032 13265
rect 57588 13265 57604 13282
rect 59052 13356 59068 13373
rect 59624 13373 59826 13390
rect 59884 13390 60844 13428
rect 59884 13373 60086 13390
rect 59624 13356 59640 13373
rect 59052 13340 59640 13356
rect 58034 13282 58622 13298
rect 58034 13265 58050 13282
rect 57588 13248 57790 13265
rect 56830 13210 57790 13248
rect 57848 13248 58050 13265
rect 58606 13265 58622 13282
rect 60070 13356 60086 13373
rect 60642 13373 60844 13390
rect 60902 13390 61862 13428
rect 60902 13373 61104 13390
rect 60642 13356 60658 13373
rect 60070 13340 60658 13356
rect 59052 13282 59640 13298
rect 59052 13265 59068 13282
rect 58606 13248 58808 13265
rect 57848 13210 58808 13248
rect 58866 13248 59068 13265
rect 59624 13265 59640 13282
rect 61088 13356 61104 13373
rect 61660 13373 61862 13390
rect 61920 13390 62880 13428
rect 61920 13373 62122 13390
rect 61660 13356 61676 13373
rect 61088 13340 61676 13356
rect 60070 13282 60658 13298
rect 60070 13265 60086 13282
rect 59624 13248 59826 13265
rect 58866 13210 59826 13248
rect 59884 13248 60086 13265
rect 60642 13265 60658 13282
rect 62106 13356 62122 13373
rect 62678 13373 62880 13390
rect 62938 13390 63898 13428
rect 62938 13373 63140 13390
rect 62678 13356 62694 13373
rect 62106 13340 62694 13356
rect 61088 13282 61676 13298
rect 61088 13265 61104 13282
rect 60642 13248 60844 13265
rect 59884 13210 60844 13248
rect 60902 13248 61104 13265
rect 61660 13265 61676 13282
rect 63124 13356 63140 13373
rect 63696 13373 63898 13390
rect 63956 13390 64916 13428
rect 63956 13373 64158 13390
rect 63696 13356 63712 13373
rect 63124 13340 63712 13356
rect 62106 13282 62694 13298
rect 62106 13265 62122 13282
rect 61660 13248 61862 13265
rect 60902 13210 61862 13248
rect 61920 13248 62122 13265
rect 62678 13265 62694 13282
rect 64142 13356 64158 13373
rect 64714 13373 64916 13390
rect 64714 13356 64730 13373
rect 64142 13340 64730 13356
rect 63124 13282 63712 13298
rect 63124 13265 63140 13282
rect 62678 13248 62880 13265
rect 61920 13210 62880 13248
rect 62938 13248 63140 13265
rect 63696 13265 63712 13282
rect 64142 13282 64730 13298
rect 64142 13265 64158 13282
rect 63696 13248 63898 13265
rect 62938 13210 63898 13248
rect 63956 13248 64158 13265
rect 64714 13265 64730 13282
rect 64714 13248 64916 13265
rect 63956 13210 64916 13248
rect 67578 12950 68538 12988
rect 67578 12933 67780 12950
rect 67764 12916 67780 12933
rect 68336 12933 68538 12950
rect 68596 12950 69556 12988
rect 68596 12933 68798 12950
rect 68336 12916 68352 12933
rect 67764 12900 68352 12916
rect 68782 12916 68798 12933
rect 69354 12933 69556 12950
rect 69614 12950 70574 12988
rect 69614 12933 69816 12950
rect 69354 12916 69370 12933
rect 68782 12900 69370 12916
rect 69800 12916 69816 12933
rect 70372 12933 70574 12950
rect 70632 12950 71592 12988
rect 70632 12933 70834 12950
rect 70372 12916 70388 12933
rect 69800 12900 70388 12916
rect 70818 12916 70834 12933
rect 71390 12933 71592 12950
rect 71650 12950 72610 12988
rect 71650 12933 71852 12950
rect 71390 12916 71406 12933
rect 70818 12900 71406 12916
rect 71836 12916 71852 12933
rect 72408 12933 72610 12950
rect 72668 12950 73628 12988
rect 72668 12933 72870 12950
rect 72408 12916 72424 12933
rect 71836 12900 72424 12916
rect 72854 12916 72870 12933
rect 73426 12933 73628 12950
rect 73686 12950 74646 12988
rect 73686 12933 73888 12950
rect 73426 12916 73442 12933
rect 72854 12900 73442 12916
rect 73872 12916 73888 12933
rect 74444 12933 74646 12950
rect 74704 12950 75664 12988
rect 74704 12933 74906 12950
rect 74444 12916 74460 12933
rect 73872 12900 74460 12916
rect 74890 12916 74906 12933
rect 75462 12933 75664 12950
rect 75722 12950 76682 12988
rect 75722 12933 75924 12950
rect 75462 12916 75478 12933
rect 74890 12900 75478 12916
rect 75908 12916 75924 12933
rect 76480 12933 76682 12950
rect 76740 12950 77700 12988
rect 76740 12933 76942 12950
rect 76480 12916 76496 12933
rect 75908 12900 76496 12916
rect 76926 12916 76942 12933
rect 77498 12933 77700 12950
rect 77758 12950 78718 12988
rect 77758 12933 77960 12950
rect 77498 12916 77514 12933
rect 76926 12900 77514 12916
rect 77944 12916 77960 12933
rect 78516 12933 78718 12950
rect 78776 12950 79736 12988
rect 78776 12933 78978 12950
rect 78516 12916 78532 12933
rect 77944 12900 78532 12916
rect 78962 12916 78978 12933
rect 79534 12933 79736 12950
rect 79794 12950 80754 12988
rect 79794 12933 79996 12950
rect 79534 12916 79550 12933
rect 78962 12900 79550 12916
rect 79980 12916 79996 12933
rect 80552 12933 80754 12950
rect 80812 12950 81772 12988
rect 80812 12933 81014 12950
rect 80552 12916 80568 12933
rect 79980 12900 80568 12916
rect 80998 12916 81014 12933
rect 81570 12933 81772 12950
rect 81830 12950 82790 12988
rect 81830 12933 82032 12950
rect 81570 12916 81586 12933
rect 80998 12900 81586 12916
rect 82016 12916 82032 12933
rect 82588 12933 82790 12950
rect 82848 12950 83808 12988
rect 82848 12933 83050 12950
rect 82588 12916 82604 12933
rect 82016 12900 82604 12916
rect 83034 12916 83050 12933
rect 83606 12933 83808 12950
rect 83866 12950 84826 12988
rect 83866 12933 84068 12950
rect 83606 12916 83622 12933
rect 83034 12900 83622 12916
rect 84052 12916 84068 12933
rect 84624 12933 84826 12950
rect 84884 12950 85844 12988
rect 84884 12933 85086 12950
rect 84624 12916 84640 12933
rect 84052 12900 84640 12916
rect 85070 12916 85086 12933
rect 85642 12933 85844 12950
rect 85902 12950 86862 12988
rect 85902 12933 86104 12950
rect 85642 12916 85658 12933
rect 85070 12900 85658 12916
rect 86088 12916 86104 12933
rect 86660 12933 86862 12950
rect 86920 12950 87880 12988
rect 86920 12933 87122 12950
rect 86660 12916 86676 12933
rect 86088 12900 86676 12916
rect 87106 12916 87122 12933
rect 87678 12933 87880 12950
rect 87678 12916 87694 12933
rect 87106 12900 87694 12916
rect 55812 12572 56772 12610
rect 55812 12555 56014 12572
rect 55998 12538 56014 12555
rect 56570 12555 56772 12572
rect 56830 12572 57790 12610
rect 56830 12555 57032 12572
rect 56570 12538 56586 12555
rect 55998 12522 56586 12538
rect 57016 12538 57032 12555
rect 57588 12555 57790 12572
rect 57848 12572 58808 12610
rect 57848 12555 58050 12572
rect 57588 12538 57604 12555
rect 57016 12522 57604 12538
rect 55998 12464 56586 12480
rect 55998 12447 56014 12464
rect 55812 12430 56014 12447
rect 56570 12447 56586 12464
rect 58034 12538 58050 12555
rect 58606 12555 58808 12572
rect 58866 12572 59826 12610
rect 58866 12555 59068 12572
rect 58606 12538 58622 12555
rect 58034 12522 58622 12538
rect 57016 12464 57604 12480
rect 57016 12447 57032 12464
rect 56570 12430 56772 12447
rect 55812 12392 56772 12430
rect 56830 12430 57032 12447
rect 57588 12447 57604 12464
rect 59052 12538 59068 12555
rect 59624 12555 59826 12572
rect 59884 12572 60844 12610
rect 59884 12555 60086 12572
rect 59624 12538 59640 12555
rect 59052 12522 59640 12538
rect 58034 12464 58622 12480
rect 58034 12447 58050 12464
rect 57588 12430 57790 12447
rect 56830 12392 57790 12430
rect 57848 12430 58050 12447
rect 58606 12447 58622 12464
rect 60070 12538 60086 12555
rect 60642 12555 60844 12572
rect 60902 12572 61862 12610
rect 60902 12555 61104 12572
rect 60642 12538 60658 12555
rect 60070 12522 60658 12538
rect 59052 12464 59640 12480
rect 59052 12447 59068 12464
rect 58606 12430 58808 12447
rect 57848 12392 58808 12430
rect 58866 12430 59068 12447
rect 59624 12447 59640 12464
rect 61088 12538 61104 12555
rect 61660 12555 61862 12572
rect 61920 12572 62880 12610
rect 61920 12555 62122 12572
rect 61660 12538 61676 12555
rect 61088 12522 61676 12538
rect 60070 12464 60658 12480
rect 60070 12447 60086 12464
rect 59624 12430 59826 12447
rect 58866 12392 59826 12430
rect 59884 12430 60086 12447
rect 60642 12447 60658 12464
rect 62106 12538 62122 12555
rect 62678 12555 62880 12572
rect 62938 12572 63898 12610
rect 62938 12555 63140 12572
rect 62678 12538 62694 12555
rect 62106 12522 62694 12538
rect 61088 12464 61676 12480
rect 61088 12447 61104 12464
rect 60642 12430 60844 12447
rect 59884 12392 60844 12430
rect 60902 12430 61104 12447
rect 61660 12447 61676 12464
rect 63124 12538 63140 12555
rect 63696 12555 63898 12572
rect 63956 12572 64916 12610
rect 63956 12555 64158 12572
rect 63696 12538 63712 12555
rect 63124 12522 63712 12538
rect 62106 12464 62694 12480
rect 62106 12447 62122 12464
rect 61660 12430 61862 12447
rect 60902 12392 61862 12430
rect 61920 12430 62122 12447
rect 62678 12447 62694 12464
rect 64142 12538 64158 12555
rect 64714 12555 64916 12572
rect 64714 12538 64730 12555
rect 64142 12522 64730 12538
rect 63124 12464 63712 12480
rect 63124 12447 63140 12464
rect 62678 12430 62880 12447
rect 61920 12392 62880 12430
rect 62938 12430 63140 12447
rect 63696 12447 63712 12464
rect 64142 12464 64730 12480
rect 64142 12447 64158 12464
rect 63696 12430 63898 12447
rect 62938 12392 63898 12430
rect 63956 12430 64158 12447
rect 64714 12447 64730 12464
rect 64714 12430 64916 12447
rect 63956 12392 64916 12430
rect 67764 12428 68352 12444
rect 67764 12411 67780 12428
rect 67578 12394 67780 12411
rect 68336 12411 68352 12428
rect 68782 12428 69370 12444
rect 68782 12411 68798 12428
rect 68336 12394 68538 12411
rect 67578 12356 68538 12394
rect 68596 12394 68798 12411
rect 69354 12411 69370 12428
rect 69800 12428 70388 12444
rect 69800 12411 69816 12428
rect 69354 12394 69556 12411
rect 68596 12356 69556 12394
rect 69614 12394 69816 12411
rect 70372 12411 70388 12428
rect 70818 12428 71406 12444
rect 70818 12411 70834 12428
rect 70372 12394 70574 12411
rect 69614 12356 70574 12394
rect 70632 12394 70834 12411
rect 71390 12411 71406 12428
rect 71836 12428 72424 12444
rect 71836 12411 71852 12428
rect 71390 12394 71592 12411
rect 70632 12356 71592 12394
rect 71650 12394 71852 12411
rect 72408 12411 72424 12428
rect 72854 12428 73442 12444
rect 72854 12411 72870 12428
rect 72408 12394 72610 12411
rect 71650 12356 72610 12394
rect 72668 12394 72870 12411
rect 73426 12411 73442 12428
rect 73872 12428 74460 12444
rect 73872 12411 73888 12428
rect 73426 12394 73628 12411
rect 72668 12356 73628 12394
rect 73686 12394 73888 12411
rect 74444 12411 74460 12428
rect 74890 12428 75478 12444
rect 74890 12411 74906 12428
rect 74444 12394 74646 12411
rect 73686 12356 74646 12394
rect 74704 12394 74906 12411
rect 75462 12411 75478 12428
rect 75908 12428 76496 12444
rect 75908 12411 75924 12428
rect 75462 12394 75664 12411
rect 74704 12356 75664 12394
rect 75722 12394 75924 12411
rect 76480 12411 76496 12428
rect 76926 12428 77514 12444
rect 76926 12411 76942 12428
rect 76480 12394 76682 12411
rect 75722 12356 76682 12394
rect 76740 12394 76942 12411
rect 77498 12411 77514 12428
rect 77944 12428 78532 12444
rect 77944 12411 77960 12428
rect 77498 12394 77700 12411
rect 76740 12356 77700 12394
rect 77758 12394 77960 12411
rect 78516 12411 78532 12428
rect 78962 12428 79550 12444
rect 78962 12411 78978 12428
rect 78516 12394 78718 12411
rect 77758 12356 78718 12394
rect 78776 12394 78978 12411
rect 79534 12411 79550 12428
rect 79980 12428 80568 12444
rect 79980 12411 79996 12428
rect 79534 12394 79736 12411
rect 78776 12356 79736 12394
rect 79794 12394 79996 12411
rect 80552 12411 80568 12428
rect 80998 12428 81586 12444
rect 80998 12411 81014 12428
rect 80552 12394 80754 12411
rect 79794 12356 80754 12394
rect 80812 12394 81014 12411
rect 81570 12411 81586 12428
rect 82016 12428 82604 12444
rect 82016 12411 82032 12428
rect 81570 12394 81772 12411
rect 80812 12356 81772 12394
rect 81830 12394 82032 12411
rect 82588 12411 82604 12428
rect 83034 12428 83622 12444
rect 83034 12411 83050 12428
rect 82588 12394 82790 12411
rect 81830 12356 82790 12394
rect 82848 12394 83050 12411
rect 83606 12411 83622 12428
rect 84052 12428 84640 12444
rect 84052 12411 84068 12428
rect 83606 12394 83808 12411
rect 82848 12356 83808 12394
rect 83866 12394 84068 12411
rect 84624 12411 84640 12428
rect 85070 12428 85658 12444
rect 85070 12411 85086 12428
rect 84624 12394 84826 12411
rect 83866 12356 84826 12394
rect 84884 12394 85086 12411
rect 85642 12411 85658 12428
rect 86088 12428 86676 12444
rect 86088 12411 86104 12428
rect 85642 12394 85844 12411
rect 84884 12356 85844 12394
rect 85902 12394 86104 12411
rect 86660 12411 86676 12428
rect 87106 12428 87694 12444
rect 87106 12411 87122 12428
rect 86660 12394 86862 12411
rect 85902 12356 86862 12394
rect 86920 12394 87122 12411
rect 87678 12411 87694 12428
rect 87678 12394 87880 12411
rect 86920 12356 87880 12394
rect 55812 11754 56772 11792
rect 55812 11737 56014 11754
rect 55998 11720 56014 11737
rect 56570 11737 56772 11754
rect 56830 11754 57790 11792
rect 56830 11737 57032 11754
rect 56570 11720 56586 11737
rect 55998 11704 56586 11720
rect 57016 11720 57032 11737
rect 57588 11737 57790 11754
rect 57848 11754 58808 11792
rect 57848 11737 58050 11754
rect 57588 11720 57604 11737
rect 57016 11704 57604 11720
rect 55998 11646 56586 11662
rect 55998 11629 56014 11646
rect 55812 11612 56014 11629
rect 56570 11629 56586 11646
rect 58034 11720 58050 11737
rect 58606 11737 58808 11754
rect 58866 11754 59826 11792
rect 58866 11737 59068 11754
rect 58606 11720 58622 11737
rect 58034 11704 58622 11720
rect 57016 11646 57604 11662
rect 57016 11629 57032 11646
rect 56570 11612 56772 11629
rect 55812 11574 56772 11612
rect 56830 11612 57032 11629
rect 57588 11629 57604 11646
rect 59052 11720 59068 11737
rect 59624 11737 59826 11754
rect 59884 11754 60844 11792
rect 59884 11737 60086 11754
rect 59624 11720 59640 11737
rect 59052 11704 59640 11720
rect 58034 11646 58622 11662
rect 58034 11629 58050 11646
rect 57588 11612 57790 11629
rect 56830 11574 57790 11612
rect 57848 11612 58050 11629
rect 58606 11629 58622 11646
rect 60070 11720 60086 11737
rect 60642 11737 60844 11754
rect 60902 11754 61862 11792
rect 60902 11737 61104 11754
rect 60642 11720 60658 11737
rect 60070 11704 60658 11720
rect 59052 11646 59640 11662
rect 59052 11629 59068 11646
rect 58606 11612 58808 11629
rect 57848 11574 58808 11612
rect 58866 11612 59068 11629
rect 59624 11629 59640 11646
rect 61088 11720 61104 11737
rect 61660 11737 61862 11754
rect 61920 11754 62880 11792
rect 61920 11737 62122 11754
rect 61660 11720 61676 11737
rect 61088 11704 61676 11720
rect 60070 11646 60658 11662
rect 60070 11629 60086 11646
rect 59624 11612 59826 11629
rect 58866 11574 59826 11612
rect 59884 11612 60086 11629
rect 60642 11629 60658 11646
rect 62106 11720 62122 11737
rect 62678 11737 62880 11754
rect 62938 11754 63898 11792
rect 62938 11737 63140 11754
rect 62678 11720 62694 11737
rect 62106 11704 62694 11720
rect 61088 11646 61676 11662
rect 61088 11629 61104 11646
rect 60642 11612 60844 11629
rect 59884 11574 60844 11612
rect 60902 11612 61104 11629
rect 61660 11629 61676 11646
rect 63124 11720 63140 11737
rect 63696 11737 63898 11754
rect 63956 11754 64916 11792
rect 63956 11737 64158 11754
rect 63696 11720 63712 11737
rect 63124 11704 63712 11720
rect 62106 11646 62694 11662
rect 62106 11629 62122 11646
rect 61660 11612 61862 11629
rect 60902 11574 61862 11612
rect 61920 11612 62122 11629
rect 62678 11629 62694 11646
rect 64142 11720 64158 11737
rect 64714 11737 64916 11754
rect 64714 11720 64730 11737
rect 64142 11704 64730 11720
rect 63124 11646 63712 11662
rect 63124 11629 63140 11646
rect 62678 11612 62880 11629
rect 61920 11574 62880 11612
rect 62938 11612 63140 11629
rect 63696 11629 63712 11646
rect 67578 11718 68538 11756
rect 67578 11701 67780 11718
rect 67764 11684 67780 11701
rect 68336 11701 68538 11718
rect 68596 11718 69556 11756
rect 68596 11701 68798 11718
rect 68336 11684 68352 11701
rect 67764 11668 68352 11684
rect 68782 11684 68798 11701
rect 69354 11701 69556 11718
rect 69614 11718 70574 11756
rect 69614 11701 69816 11718
rect 69354 11684 69370 11701
rect 68782 11668 69370 11684
rect 69800 11684 69816 11701
rect 70372 11701 70574 11718
rect 70632 11718 71592 11756
rect 70632 11701 70834 11718
rect 70372 11684 70388 11701
rect 69800 11668 70388 11684
rect 70818 11684 70834 11701
rect 71390 11701 71592 11718
rect 71650 11718 72610 11756
rect 71650 11701 71852 11718
rect 71390 11684 71406 11701
rect 70818 11668 71406 11684
rect 71836 11684 71852 11701
rect 72408 11701 72610 11718
rect 72668 11718 73628 11756
rect 72668 11701 72870 11718
rect 72408 11684 72424 11701
rect 71836 11668 72424 11684
rect 72854 11684 72870 11701
rect 73426 11701 73628 11718
rect 73686 11718 74646 11756
rect 73686 11701 73888 11718
rect 73426 11684 73442 11701
rect 72854 11668 73442 11684
rect 73872 11684 73888 11701
rect 74444 11701 74646 11718
rect 74704 11718 75664 11756
rect 74704 11701 74906 11718
rect 74444 11684 74460 11701
rect 73872 11668 74460 11684
rect 74890 11684 74906 11701
rect 75462 11701 75664 11718
rect 75722 11718 76682 11756
rect 75722 11701 75924 11718
rect 75462 11684 75478 11701
rect 74890 11668 75478 11684
rect 75908 11684 75924 11701
rect 76480 11701 76682 11718
rect 76740 11718 77700 11756
rect 76740 11701 76942 11718
rect 76480 11684 76496 11701
rect 75908 11668 76496 11684
rect 76926 11684 76942 11701
rect 77498 11701 77700 11718
rect 77758 11718 78718 11756
rect 77758 11701 77960 11718
rect 77498 11684 77514 11701
rect 76926 11668 77514 11684
rect 77944 11684 77960 11701
rect 78516 11701 78718 11718
rect 78776 11718 79736 11756
rect 78776 11701 78978 11718
rect 78516 11684 78532 11701
rect 77944 11668 78532 11684
rect 78962 11684 78978 11701
rect 79534 11701 79736 11718
rect 79794 11718 80754 11756
rect 79794 11701 79996 11718
rect 79534 11684 79550 11701
rect 78962 11668 79550 11684
rect 79980 11684 79996 11701
rect 80552 11701 80754 11718
rect 80812 11718 81772 11756
rect 80812 11701 81014 11718
rect 80552 11684 80568 11701
rect 79980 11668 80568 11684
rect 80998 11684 81014 11701
rect 81570 11701 81772 11718
rect 81830 11718 82790 11756
rect 81830 11701 82032 11718
rect 81570 11684 81586 11701
rect 80998 11668 81586 11684
rect 82016 11684 82032 11701
rect 82588 11701 82790 11718
rect 82848 11718 83808 11756
rect 82848 11701 83050 11718
rect 82588 11684 82604 11701
rect 82016 11668 82604 11684
rect 83034 11684 83050 11701
rect 83606 11701 83808 11718
rect 83866 11718 84826 11756
rect 83866 11701 84068 11718
rect 83606 11684 83622 11701
rect 83034 11668 83622 11684
rect 84052 11684 84068 11701
rect 84624 11701 84826 11718
rect 84884 11718 85844 11756
rect 84884 11701 85086 11718
rect 84624 11684 84640 11701
rect 84052 11668 84640 11684
rect 85070 11684 85086 11701
rect 85642 11701 85844 11718
rect 85902 11718 86862 11756
rect 85902 11701 86104 11718
rect 85642 11684 85658 11701
rect 85070 11668 85658 11684
rect 86088 11684 86104 11701
rect 86660 11701 86862 11718
rect 86920 11718 87880 11756
rect 86920 11701 87122 11718
rect 86660 11684 86676 11701
rect 86088 11668 86676 11684
rect 87106 11684 87122 11701
rect 87678 11701 87880 11718
rect 87678 11684 87694 11701
rect 87106 11668 87694 11684
rect 64142 11646 64730 11662
rect 64142 11629 64158 11646
rect 63696 11612 63898 11629
rect 62938 11574 63898 11612
rect 63956 11612 64158 11629
rect 64714 11629 64730 11646
rect 64714 11612 64916 11629
rect 63956 11574 64916 11612
rect 67762 11194 68350 11210
rect 67762 11177 67778 11194
rect 67576 11160 67778 11177
rect 68334 11177 68350 11194
rect 68780 11194 69368 11210
rect 68780 11177 68796 11194
rect 68334 11160 68536 11177
rect 67576 11122 68536 11160
rect 68594 11160 68796 11177
rect 69352 11177 69368 11194
rect 69798 11194 70386 11210
rect 69798 11177 69814 11194
rect 69352 11160 69554 11177
rect 68594 11122 69554 11160
rect 69612 11160 69814 11177
rect 70370 11177 70386 11194
rect 70816 11194 71404 11210
rect 70816 11177 70832 11194
rect 70370 11160 70572 11177
rect 69612 11122 70572 11160
rect 70630 11160 70832 11177
rect 71388 11177 71404 11194
rect 71834 11194 72422 11210
rect 71834 11177 71850 11194
rect 71388 11160 71590 11177
rect 70630 11122 71590 11160
rect 71648 11160 71850 11177
rect 72406 11177 72422 11194
rect 72852 11194 73440 11210
rect 72852 11177 72868 11194
rect 72406 11160 72608 11177
rect 71648 11122 72608 11160
rect 72666 11160 72868 11177
rect 73424 11177 73440 11194
rect 73870 11194 74458 11210
rect 73870 11177 73886 11194
rect 73424 11160 73626 11177
rect 72666 11122 73626 11160
rect 73684 11160 73886 11177
rect 74442 11177 74458 11194
rect 74888 11194 75476 11210
rect 74888 11177 74904 11194
rect 74442 11160 74644 11177
rect 73684 11122 74644 11160
rect 74702 11160 74904 11177
rect 75460 11177 75476 11194
rect 75906 11194 76494 11210
rect 75906 11177 75922 11194
rect 75460 11160 75662 11177
rect 74702 11122 75662 11160
rect 75720 11160 75922 11177
rect 76478 11177 76494 11194
rect 76924 11194 77512 11210
rect 76924 11177 76940 11194
rect 76478 11160 76680 11177
rect 75720 11122 76680 11160
rect 76738 11160 76940 11177
rect 77496 11177 77512 11194
rect 77942 11194 78530 11210
rect 77942 11177 77958 11194
rect 77496 11160 77698 11177
rect 76738 11122 77698 11160
rect 77756 11160 77958 11177
rect 78514 11177 78530 11194
rect 78960 11194 79548 11210
rect 78960 11177 78976 11194
rect 78514 11160 78716 11177
rect 77756 11122 78716 11160
rect 78774 11160 78976 11177
rect 79532 11177 79548 11194
rect 79978 11194 80566 11210
rect 79978 11177 79994 11194
rect 79532 11160 79734 11177
rect 78774 11122 79734 11160
rect 79792 11160 79994 11177
rect 80550 11177 80566 11194
rect 80996 11194 81584 11210
rect 80996 11177 81012 11194
rect 80550 11160 80752 11177
rect 79792 11122 80752 11160
rect 80810 11160 81012 11177
rect 81568 11177 81584 11194
rect 82014 11194 82602 11210
rect 82014 11177 82030 11194
rect 81568 11160 81770 11177
rect 80810 11122 81770 11160
rect 81828 11160 82030 11177
rect 82586 11177 82602 11194
rect 83032 11194 83620 11210
rect 83032 11177 83048 11194
rect 82586 11160 82788 11177
rect 81828 11122 82788 11160
rect 82846 11160 83048 11177
rect 83604 11177 83620 11194
rect 84050 11194 84638 11210
rect 84050 11177 84066 11194
rect 83604 11160 83806 11177
rect 82846 11122 83806 11160
rect 83864 11160 84066 11177
rect 84622 11177 84638 11194
rect 85068 11194 85656 11210
rect 85068 11177 85084 11194
rect 84622 11160 84824 11177
rect 83864 11122 84824 11160
rect 84882 11160 85084 11177
rect 85640 11177 85656 11194
rect 86086 11194 86674 11210
rect 86086 11177 86102 11194
rect 85640 11160 85842 11177
rect 84882 11122 85842 11160
rect 85900 11160 86102 11177
rect 86658 11177 86674 11194
rect 87104 11194 87692 11210
rect 87104 11177 87120 11194
rect 86658 11160 86860 11177
rect 85900 11122 86860 11160
rect 86918 11160 87120 11177
rect 87676 11177 87692 11194
rect 87676 11160 87878 11177
rect 86918 11122 87878 11160
rect 55812 10936 56772 10974
rect 55812 10919 56014 10936
rect 55998 10902 56014 10919
rect 56570 10919 56772 10936
rect 56830 10936 57790 10974
rect 56830 10919 57032 10936
rect 56570 10902 56586 10919
rect 55998 10886 56586 10902
rect 57016 10902 57032 10919
rect 57588 10919 57790 10936
rect 57848 10936 58808 10974
rect 57848 10919 58050 10936
rect 57588 10902 57604 10919
rect 57016 10886 57604 10902
rect 55998 10828 56586 10844
rect 55998 10811 56014 10828
rect 55812 10794 56014 10811
rect 56570 10811 56586 10828
rect 58034 10902 58050 10919
rect 58606 10919 58808 10936
rect 58866 10936 59826 10974
rect 58866 10919 59068 10936
rect 58606 10902 58622 10919
rect 58034 10886 58622 10902
rect 57016 10828 57604 10844
rect 57016 10811 57032 10828
rect 56570 10794 56772 10811
rect 55812 10756 56772 10794
rect 56830 10794 57032 10811
rect 57588 10811 57604 10828
rect 59052 10902 59068 10919
rect 59624 10919 59826 10936
rect 59884 10936 60844 10974
rect 59884 10919 60086 10936
rect 59624 10902 59640 10919
rect 59052 10886 59640 10902
rect 58034 10828 58622 10844
rect 58034 10811 58050 10828
rect 57588 10794 57790 10811
rect 56830 10756 57790 10794
rect 57848 10794 58050 10811
rect 58606 10811 58622 10828
rect 60070 10902 60086 10919
rect 60642 10919 60844 10936
rect 60902 10936 61862 10974
rect 60902 10919 61104 10936
rect 60642 10902 60658 10919
rect 60070 10886 60658 10902
rect 59052 10828 59640 10844
rect 59052 10811 59068 10828
rect 58606 10794 58808 10811
rect 57848 10756 58808 10794
rect 58866 10794 59068 10811
rect 59624 10811 59640 10828
rect 61088 10902 61104 10919
rect 61660 10919 61862 10936
rect 61920 10936 62880 10974
rect 61920 10919 62122 10936
rect 61660 10902 61676 10919
rect 61088 10886 61676 10902
rect 60070 10828 60658 10844
rect 60070 10811 60086 10828
rect 59624 10794 59826 10811
rect 58866 10756 59826 10794
rect 59884 10794 60086 10811
rect 60642 10811 60658 10828
rect 62106 10902 62122 10919
rect 62678 10919 62880 10936
rect 62938 10936 63898 10974
rect 62938 10919 63140 10936
rect 62678 10902 62694 10919
rect 62106 10886 62694 10902
rect 61088 10828 61676 10844
rect 61088 10811 61104 10828
rect 60642 10794 60844 10811
rect 59884 10756 60844 10794
rect 60902 10794 61104 10811
rect 61660 10811 61676 10828
rect 63124 10902 63140 10919
rect 63696 10919 63898 10936
rect 63956 10936 64916 10974
rect 63956 10919 64158 10936
rect 63696 10902 63712 10919
rect 63124 10886 63712 10902
rect 62106 10828 62694 10844
rect 62106 10811 62122 10828
rect 61660 10794 61862 10811
rect 60902 10756 61862 10794
rect 61920 10794 62122 10811
rect 62678 10811 62694 10828
rect 64142 10902 64158 10919
rect 64714 10919 64916 10936
rect 64714 10902 64730 10919
rect 64142 10886 64730 10902
rect 63124 10828 63712 10844
rect 63124 10811 63140 10828
rect 62678 10794 62880 10811
rect 61920 10756 62880 10794
rect 62938 10794 63140 10811
rect 63696 10811 63712 10828
rect 64142 10828 64730 10844
rect 64142 10811 64158 10828
rect 63696 10794 63898 10811
rect 62938 10756 63898 10794
rect 63956 10794 64158 10811
rect 64714 10811 64730 10828
rect 64714 10794 64916 10811
rect 63956 10756 64916 10794
rect 67576 10484 68536 10522
rect 67576 10467 67778 10484
rect 67762 10450 67778 10467
rect 68334 10467 68536 10484
rect 68594 10484 69554 10522
rect 68594 10467 68796 10484
rect 68334 10450 68350 10467
rect 67762 10434 68350 10450
rect 68780 10450 68796 10467
rect 69352 10467 69554 10484
rect 69612 10484 70572 10522
rect 69612 10467 69814 10484
rect 69352 10450 69368 10467
rect 68780 10434 69368 10450
rect 69798 10450 69814 10467
rect 70370 10467 70572 10484
rect 70630 10484 71590 10522
rect 70630 10467 70832 10484
rect 70370 10450 70386 10467
rect 69798 10434 70386 10450
rect 70816 10450 70832 10467
rect 71388 10467 71590 10484
rect 71648 10484 72608 10522
rect 71648 10467 71850 10484
rect 71388 10450 71404 10467
rect 70816 10434 71404 10450
rect 71834 10450 71850 10467
rect 72406 10467 72608 10484
rect 72666 10484 73626 10522
rect 72666 10467 72868 10484
rect 72406 10450 72422 10467
rect 71834 10434 72422 10450
rect 72852 10450 72868 10467
rect 73424 10467 73626 10484
rect 73684 10484 74644 10522
rect 73684 10467 73886 10484
rect 73424 10450 73440 10467
rect 72852 10434 73440 10450
rect 73870 10450 73886 10467
rect 74442 10467 74644 10484
rect 74702 10484 75662 10522
rect 74702 10467 74904 10484
rect 74442 10450 74458 10467
rect 73870 10434 74458 10450
rect 74888 10450 74904 10467
rect 75460 10467 75662 10484
rect 75720 10484 76680 10522
rect 75720 10467 75922 10484
rect 75460 10450 75476 10467
rect 74888 10434 75476 10450
rect 75906 10450 75922 10467
rect 76478 10467 76680 10484
rect 76738 10484 77698 10522
rect 76738 10467 76940 10484
rect 76478 10450 76494 10467
rect 75906 10434 76494 10450
rect 76924 10450 76940 10467
rect 77496 10467 77698 10484
rect 77756 10484 78716 10522
rect 77756 10467 77958 10484
rect 77496 10450 77512 10467
rect 76924 10434 77512 10450
rect 77942 10450 77958 10467
rect 78514 10467 78716 10484
rect 78774 10484 79734 10522
rect 78774 10467 78976 10484
rect 78514 10450 78530 10467
rect 77942 10434 78530 10450
rect 78960 10450 78976 10467
rect 79532 10467 79734 10484
rect 79792 10484 80752 10522
rect 79792 10467 79994 10484
rect 79532 10450 79548 10467
rect 78960 10434 79548 10450
rect 79978 10450 79994 10467
rect 80550 10467 80752 10484
rect 80810 10484 81770 10522
rect 80810 10467 81012 10484
rect 80550 10450 80566 10467
rect 79978 10434 80566 10450
rect 80996 10450 81012 10467
rect 81568 10467 81770 10484
rect 81828 10484 82788 10522
rect 81828 10467 82030 10484
rect 81568 10450 81584 10467
rect 80996 10434 81584 10450
rect 82014 10450 82030 10467
rect 82586 10467 82788 10484
rect 82846 10484 83806 10522
rect 82846 10467 83048 10484
rect 82586 10450 82602 10467
rect 82014 10434 82602 10450
rect 83032 10450 83048 10467
rect 83604 10467 83806 10484
rect 83864 10484 84824 10522
rect 83864 10467 84066 10484
rect 83604 10450 83620 10467
rect 83032 10434 83620 10450
rect 84050 10450 84066 10467
rect 84622 10467 84824 10484
rect 84882 10484 85842 10522
rect 84882 10467 85084 10484
rect 84622 10450 84638 10467
rect 84050 10434 84638 10450
rect 85068 10450 85084 10467
rect 85640 10467 85842 10484
rect 85900 10484 86860 10522
rect 85900 10467 86102 10484
rect 85640 10450 85656 10467
rect 85068 10434 85656 10450
rect 86086 10450 86102 10467
rect 86658 10467 86860 10484
rect 86918 10484 87878 10522
rect 86918 10467 87120 10484
rect 86658 10450 86674 10467
rect 86086 10434 86674 10450
rect 87104 10450 87120 10467
rect 87676 10467 87878 10484
rect 87676 10450 87692 10467
rect 87104 10434 87692 10450
rect 55812 10118 56772 10156
rect 55812 10101 56014 10118
rect 55998 10084 56014 10101
rect 56570 10101 56772 10118
rect 56830 10118 57790 10156
rect 56830 10101 57032 10118
rect 56570 10084 56586 10101
rect 55998 10068 56586 10084
rect 57016 10084 57032 10101
rect 57588 10101 57790 10118
rect 57848 10118 58808 10156
rect 57848 10101 58050 10118
rect 57588 10084 57604 10101
rect 57016 10068 57604 10084
rect 55998 10010 56586 10026
rect 55998 9993 56014 10010
rect 55812 9976 56014 9993
rect 56570 9993 56586 10010
rect 58034 10084 58050 10101
rect 58606 10101 58808 10118
rect 58866 10118 59826 10156
rect 58866 10101 59068 10118
rect 58606 10084 58622 10101
rect 58034 10068 58622 10084
rect 57016 10010 57604 10026
rect 57016 9993 57032 10010
rect 56570 9976 56772 9993
rect 55812 9938 56772 9976
rect 56830 9976 57032 9993
rect 57588 9993 57604 10010
rect 59052 10084 59068 10101
rect 59624 10101 59826 10118
rect 59884 10118 60844 10156
rect 59884 10101 60086 10118
rect 59624 10084 59640 10101
rect 59052 10068 59640 10084
rect 58034 10010 58622 10026
rect 58034 9993 58050 10010
rect 57588 9976 57790 9993
rect 56830 9938 57790 9976
rect 57848 9976 58050 9993
rect 58606 9993 58622 10010
rect 60070 10084 60086 10101
rect 60642 10101 60844 10118
rect 60902 10118 61862 10156
rect 60902 10101 61104 10118
rect 60642 10084 60658 10101
rect 60070 10068 60658 10084
rect 59052 10010 59640 10026
rect 59052 9993 59068 10010
rect 58606 9976 58808 9993
rect 57848 9938 58808 9976
rect 58866 9976 59068 9993
rect 59624 9993 59640 10010
rect 61088 10084 61104 10101
rect 61660 10101 61862 10118
rect 61920 10118 62880 10156
rect 61920 10101 62122 10118
rect 61660 10084 61676 10101
rect 61088 10068 61676 10084
rect 60070 10010 60658 10026
rect 60070 9993 60086 10010
rect 59624 9976 59826 9993
rect 58866 9938 59826 9976
rect 59884 9976 60086 9993
rect 60642 9993 60658 10010
rect 62106 10084 62122 10101
rect 62678 10101 62880 10118
rect 62938 10118 63898 10156
rect 62938 10101 63140 10118
rect 62678 10084 62694 10101
rect 62106 10068 62694 10084
rect 61088 10010 61676 10026
rect 61088 9993 61104 10010
rect 60642 9976 60844 9993
rect 59884 9938 60844 9976
rect 60902 9976 61104 9993
rect 61660 9993 61676 10010
rect 63124 10084 63140 10101
rect 63696 10101 63898 10118
rect 63956 10118 64916 10156
rect 63956 10101 64158 10118
rect 63696 10084 63712 10101
rect 63124 10068 63712 10084
rect 62106 10010 62694 10026
rect 62106 9993 62122 10010
rect 61660 9976 61862 9993
rect 60902 9938 61862 9976
rect 61920 9976 62122 9993
rect 62678 9993 62694 10010
rect 64142 10084 64158 10101
rect 64714 10101 64916 10118
rect 64714 10084 64730 10101
rect 64142 10068 64730 10084
rect 63124 10010 63712 10026
rect 63124 9993 63140 10010
rect 62678 9976 62880 9993
rect 61920 9938 62880 9976
rect 62938 9976 63140 9993
rect 63696 9993 63712 10010
rect 64142 10010 64730 10026
rect 64142 9993 64158 10010
rect 63696 9976 63898 9993
rect 62938 9938 63898 9976
rect 63956 9976 64158 9993
rect 64714 9993 64730 10010
rect 64714 9976 64916 9993
rect 63956 9938 64916 9976
rect 67762 9960 68350 9976
rect 67762 9943 67778 9960
rect 67576 9926 67778 9943
rect 68334 9943 68350 9960
rect 68780 9960 69368 9976
rect 68780 9943 68796 9960
rect 68334 9926 68536 9943
rect 67576 9888 68536 9926
rect 68594 9926 68796 9943
rect 69352 9943 69368 9960
rect 69798 9960 70386 9976
rect 69798 9943 69814 9960
rect 69352 9926 69554 9943
rect 68594 9888 69554 9926
rect 69612 9926 69814 9943
rect 70370 9943 70386 9960
rect 70816 9960 71404 9976
rect 70816 9943 70832 9960
rect 70370 9926 70572 9943
rect 69612 9888 70572 9926
rect 70630 9926 70832 9943
rect 71388 9943 71404 9960
rect 71834 9960 72422 9976
rect 71834 9943 71850 9960
rect 71388 9926 71590 9943
rect 70630 9888 71590 9926
rect 71648 9926 71850 9943
rect 72406 9943 72422 9960
rect 72852 9960 73440 9976
rect 72852 9943 72868 9960
rect 72406 9926 72608 9943
rect 71648 9888 72608 9926
rect 72666 9926 72868 9943
rect 73424 9943 73440 9960
rect 73870 9960 74458 9976
rect 73870 9943 73886 9960
rect 73424 9926 73626 9943
rect 72666 9888 73626 9926
rect 73684 9926 73886 9943
rect 74442 9943 74458 9960
rect 74888 9960 75476 9976
rect 74888 9943 74904 9960
rect 74442 9926 74644 9943
rect 73684 9888 74644 9926
rect 74702 9926 74904 9943
rect 75460 9943 75476 9960
rect 75906 9960 76494 9976
rect 75906 9943 75922 9960
rect 75460 9926 75662 9943
rect 74702 9888 75662 9926
rect 75720 9926 75922 9943
rect 76478 9943 76494 9960
rect 76924 9960 77512 9976
rect 76924 9943 76940 9960
rect 76478 9926 76680 9943
rect 75720 9888 76680 9926
rect 76738 9926 76940 9943
rect 77496 9943 77512 9960
rect 77942 9960 78530 9976
rect 77942 9943 77958 9960
rect 77496 9926 77698 9943
rect 76738 9888 77698 9926
rect 77756 9926 77958 9943
rect 78514 9943 78530 9960
rect 78960 9960 79548 9976
rect 78960 9943 78976 9960
rect 78514 9926 78716 9943
rect 77756 9888 78716 9926
rect 78774 9926 78976 9943
rect 79532 9943 79548 9960
rect 79978 9960 80566 9976
rect 79978 9943 79994 9960
rect 79532 9926 79734 9943
rect 78774 9888 79734 9926
rect 79792 9926 79994 9943
rect 80550 9943 80566 9960
rect 80996 9960 81584 9976
rect 80996 9943 81012 9960
rect 80550 9926 80752 9943
rect 79792 9888 80752 9926
rect 80810 9926 81012 9943
rect 81568 9943 81584 9960
rect 82014 9960 82602 9976
rect 82014 9943 82030 9960
rect 81568 9926 81770 9943
rect 80810 9888 81770 9926
rect 81828 9926 82030 9943
rect 82586 9943 82602 9960
rect 83032 9960 83620 9976
rect 83032 9943 83048 9960
rect 82586 9926 82788 9943
rect 81828 9888 82788 9926
rect 82846 9926 83048 9943
rect 83604 9943 83620 9960
rect 84050 9960 84638 9976
rect 84050 9943 84066 9960
rect 83604 9926 83806 9943
rect 82846 9888 83806 9926
rect 83864 9926 84066 9943
rect 84622 9943 84638 9960
rect 85068 9960 85656 9976
rect 85068 9943 85084 9960
rect 84622 9926 84824 9943
rect 83864 9888 84824 9926
rect 84882 9926 85084 9943
rect 85640 9943 85656 9960
rect 86086 9960 86674 9976
rect 86086 9943 86102 9960
rect 85640 9926 85842 9943
rect 84882 9888 85842 9926
rect 85900 9926 86102 9943
rect 86658 9943 86674 9960
rect 87104 9960 87692 9976
rect 87104 9943 87120 9960
rect 86658 9926 86860 9943
rect 85900 9888 86860 9926
rect 86918 9926 87120 9943
rect 87676 9943 87692 9960
rect 87676 9926 87878 9943
rect 86918 9888 87878 9926
rect 55812 9300 56772 9338
rect 55812 9283 56014 9300
rect 55998 9266 56014 9283
rect 56570 9283 56772 9300
rect 56830 9300 57790 9338
rect 56830 9283 57032 9300
rect 56570 9266 56586 9283
rect 55998 9250 56586 9266
rect 57016 9266 57032 9283
rect 57588 9283 57790 9300
rect 57848 9300 58808 9338
rect 57848 9283 58050 9300
rect 57588 9266 57604 9283
rect 57016 9250 57604 9266
rect 55998 9192 56586 9208
rect 55998 9175 56014 9192
rect 55812 9158 56014 9175
rect 56570 9175 56586 9192
rect 58034 9266 58050 9283
rect 58606 9283 58808 9300
rect 58866 9300 59826 9338
rect 58866 9283 59068 9300
rect 58606 9266 58622 9283
rect 58034 9250 58622 9266
rect 57016 9192 57604 9208
rect 57016 9175 57032 9192
rect 56570 9158 56772 9175
rect 55812 9120 56772 9158
rect 56830 9158 57032 9175
rect 57588 9175 57604 9192
rect 59052 9266 59068 9283
rect 59624 9283 59826 9300
rect 59884 9300 60844 9338
rect 59884 9283 60086 9300
rect 59624 9266 59640 9283
rect 59052 9250 59640 9266
rect 58034 9192 58622 9208
rect 58034 9175 58050 9192
rect 57588 9158 57790 9175
rect 56830 9120 57790 9158
rect 57848 9158 58050 9175
rect 58606 9175 58622 9192
rect 60070 9266 60086 9283
rect 60642 9283 60844 9300
rect 60902 9300 61862 9338
rect 60902 9283 61104 9300
rect 60642 9266 60658 9283
rect 60070 9250 60658 9266
rect 59052 9192 59640 9208
rect 59052 9175 59068 9192
rect 58606 9158 58808 9175
rect 57848 9120 58808 9158
rect 58866 9158 59068 9175
rect 59624 9175 59640 9192
rect 61088 9266 61104 9283
rect 61660 9283 61862 9300
rect 61920 9300 62880 9338
rect 61920 9283 62122 9300
rect 61660 9266 61676 9283
rect 61088 9250 61676 9266
rect 60070 9192 60658 9208
rect 60070 9175 60086 9192
rect 59624 9158 59826 9175
rect 58866 9120 59826 9158
rect 59884 9158 60086 9175
rect 60642 9175 60658 9192
rect 62106 9266 62122 9283
rect 62678 9283 62880 9300
rect 62938 9300 63898 9338
rect 62938 9283 63140 9300
rect 62678 9266 62694 9283
rect 62106 9250 62694 9266
rect 61088 9192 61676 9208
rect 61088 9175 61104 9192
rect 60642 9158 60844 9175
rect 59884 9120 60844 9158
rect 60902 9158 61104 9175
rect 61660 9175 61676 9192
rect 63124 9266 63140 9283
rect 63696 9283 63898 9300
rect 63956 9300 64916 9338
rect 63956 9283 64158 9300
rect 63696 9266 63712 9283
rect 63124 9250 63712 9266
rect 62106 9192 62694 9208
rect 62106 9175 62122 9192
rect 61660 9158 61862 9175
rect 60902 9120 61862 9158
rect 61920 9158 62122 9175
rect 62678 9175 62694 9192
rect 64142 9266 64158 9283
rect 64714 9283 64916 9300
rect 64714 9266 64730 9283
rect 64142 9250 64730 9266
rect 63124 9192 63712 9208
rect 63124 9175 63140 9192
rect 62678 9158 62880 9175
rect 61920 9120 62880 9158
rect 62938 9158 63140 9175
rect 63696 9175 63712 9192
rect 67576 9250 68536 9288
rect 67576 9233 67778 9250
rect 64142 9192 64730 9208
rect 64142 9175 64158 9192
rect 63696 9158 63898 9175
rect 62938 9120 63898 9158
rect 63956 9158 64158 9175
rect 64714 9175 64730 9192
rect 67762 9216 67778 9233
rect 68334 9233 68536 9250
rect 68594 9250 69554 9288
rect 68594 9233 68796 9250
rect 68334 9216 68350 9233
rect 67762 9200 68350 9216
rect 68780 9216 68796 9233
rect 69352 9233 69554 9250
rect 69612 9250 70572 9288
rect 69612 9233 69814 9250
rect 69352 9216 69368 9233
rect 68780 9200 69368 9216
rect 69798 9216 69814 9233
rect 70370 9233 70572 9250
rect 70630 9250 71590 9288
rect 70630 9233 70832 9250
rect 70370 9216 70386 9233
rect 69798 9200 70386 9216
rect 70816 9216 70832 9233
rect 71388 9233 71590 9250
rect 71648 9250 72608 9288
rect 71648 9233 71850 9250
rect 71388 9216 71404 9233
rect 70816 9200 71404 9216
rect 71834 9216 71850 9233
rect 72406 9233 72608 9250
rect 72666 9250 73626 9288
rect 72666 9233 72868 9250
rect 72406 9216 72422 9233
rect 71834 9200 72422 9216
rect 72852 9216 72868 9233
rect 73424 9233 73626 9250
rect 73684 9250 74644 9288
rect 73684 9233 73886 9250
rect 73424 9216 73440 9233
rect 72852 9200 73440 9216
rect 73870 9216 73886 9233
rect 74442 9233 74644 9250
rect 74702 9250 75662 9288
rect 74702 9233 74904 9250
rect 74442 9216 74458 9233
rect 73870 9200 74458 9216
rect 74888 9216 74904 9233
rect 75460 9233 75662 9250
rect 75720 9250 76680 9288
rect 75720 9233 75922 9250
rect 75460 9216 75476 9233
rect 74888 9200 75476 9216
rect 75906 9216 75922 9233
rect 76478 9233 76680 9250
rect 76738 9250 77698 9288
rect 76738 9233 76940 9250
rect 76478 9216 76494 9233
rect 75906 9200 76494 9216
rect 76924 9216 76940 9233
rect 77496 9233 77698 9250
rect 77756 9250 78716 9288
rect 77756 9233 77958 9250
rect 77496 9216 77512 9233
rect 76924 9200 77512 9216
rect 77942 9216 77958 9233
rect 78514 9233 78716 9250
rect 78774 9250 79734 9288
rect 78774 9233 78976 9250
rect 78514 9216 78530 9233
rect 77942 9200 78530 9216
rect 78960 9216 78976 9233
rect 79532 9233 79734 9250
rect 79792 9250 80752 9288
rect 79792 9233 79994 9250
rect 79532 9216 79548 9233
rect 78960 9200 79548 9216
rect 79978 9216 79994 9233
rect 80550 9233 80752 9250
rect 80810 9250 81770 9288
rect 80810 9233 81012 9250
rect 80550 9216 80566 9233
rect 79978 9200 80566 9216
rect 80996 9216 81012 9233
rect 81568 9233 81770 9250
rect 81828 9250 82788 9288
rect 81828 9233 82030 9250
rect 81568 9216 81584 9233
rect 80996 9200 81584 9216
rect 82014 9216 82030 9233
rect 82586 9233 82788 9250
rect 82846 9250 83806 9288
rect 82846 9233 83048 9250
rect 82586 9216 82602 9233
rect 82014 9200 82602 9216
rect 83032 9216 83048 9233
rect 83604 9233 83806 9250
rect 83864 9250 84824 9288
rect 83864 9233 84066 9250
rect 83604 9216 83620 9233
rect 83032 9200 83620 9216
rect 84050 9216 84066 9233
rect 84622 9233 84824 9250
rect 84882 9250 85842 9288
rect 84882 9233 85084 9250
rect 84622 9216 84638 9233
rect 84050 9200 84638 9216
rect 85068 9216 85084 9233
rect 85640 9233 85842 9250
rect 85900 9250 86860 9288
rect 85900 9233 86102 9250
rect 85640 9216 85656 9233
rect 85068 9200 85656 9216
rect 86086 9216 86102 9233
rect 86658 9233 86860 9250
rect 86918 9250 87878 9288
rect 86918 9233 87120 9250
rect 86658 9216 86674 9233
rect 86086 9200 86674 9216
rect 87104 9216 87120 9233
rect 87676 9233 87878 9250
rect 87676 9216 87692 9233
rect 87104 9200 87692 9216
rect 64714 9158 64916 9175
rect 63956 9120 64916 9158
rect 67762 8728 68350 8744
rect 67762 8711 67778 8728
rect 67576 8694 67778 8711
rect 68334 8711 68350 8728
rect 68780 8728 69368 8744
rect 68780 8711 68796 8728
rect 68334 8694 68536 8711
rect 67576 8656 68536 8694
rect 68594 8694 68796 8711
rect 69352 8711 69368 8728
rect 69798 8728 70386 8744
rect 69798 8711 69814 8728
rect 69352 8694 69554 8711
rect 68594 8656 69554 8694
rect 69612 8694 69814 8711
rect 70370 8711 70386 8728
rect 70816 8728 71404 8744
rect 70816 8711 70832 8728
rect 70370 8694 70572 8711
rect 69612 8656 70572 8694
rect 70630 8694 70832 8711
rect 71388 8711 71404 8728
rect 71834 8728 72422 8744
rect 71834 8711 71850 8728
rect 71388 8694 71590 8711
rect 70630 8656 71590 8694
rect 71648 8694 71850 8711
rect 72406 8711 72422 8728
rect 72852 8728 73440 8744
rect 72852 8711 72868 8728
rect 72406 8694 72608 8711
rect 71648 8656 72608 8694
rect 72666 8694 72868 8711
rect 73424 8711 73440 8728
rect 73870 8728 74458 8744
rect 73870 8711 73886 8728
rect 73424 8694 73626 8711
rect 72666 8656 73626 8694
rect 73684 8694 73886 8711
rect 74442 8711 74458 8728
rect 74888 8728 75476 8744
rect 74888 8711 74904 8728
rect 74442 8694 74644 8711
rect 73684 8656 74644 8694
rect 74702 8694 74904 8711
rect 75460 8711 75476 8728
rect 75906 8728 76494 8744
rect 75906 8711 75922 8728
rect 75460 8694 75662 8711
rect 74702 8656 75662 8694
rect 75720 8694 75922 8711
rect 76478 8711 76494 8728
rect 76924 8728 77512 8744
rect 76924 8711 76940 8728
rect 76478 8694 76680 8711
rect 75720 8656 76680 8694
rect 76738 8694 76940 8711
rect 77496 8711 77512 8728
rect 77942 8728 78530 8744
rect 77942 8711 77958 8728
rect 77496 8694 77698 8711
rect 76738 8656 77698 8694
rect 77756 8694 77958 8711
rect 78514 8711 78530 8728
rect 78960 8728 79548 8744
rect 78960 8711 78976 8728
rect 78514 8694 78716 8711
rect 77756 8656 78716 8694
rect 78774 8694 78976 8711
rect 79532 8711 79548 8728
rect 79978 8728 80566 8744
rect 79978 8711 79994 8728
rect 79532 8694 79734 8711
rect 78774 8656 79734 8694
rect 79792 8694 79994 8711
rect 80550 8711 80566 8728
rect 80996 8728 81584 8744
rect 80996 8711 81012 8728
rect 80550 8694 80752 8711
rect 79792 8656 80752 8694
rect 80810 8694 81012 8711
rect 81568 8711 81584 8728
rect 82014 8728 82602 8744
rect 82014 8711 82030 8728
rect 81568 8694 81770 8711
rect 80810 8656 81770 8694
rect 81828 8694 82030 8711
rect 82586 8711 82602 8728
rect 83032 8728 83620 8744
rect 83032 8711 83048 8728
rect 82586 8694 82788 8711
rect 81828 8656 82788 8694
rect 82846 8694 83048 8711
rect 83604 8711 83620 8728
rect 84050 8728 84638 8744
rect 84050 8711 84066 8728
rect 83604 8694 83806 8711
rect 82846 8656 83806 8694
rect 83864 8694 84066 8711
rect 84622 8711 84638 8728
rect 85068 8728 85656 8744
rect 85068 8711 85084 8728
rect 84622 8694 84824 8711
rect 83864 8656 84824 8694
rect 84882 8694 85084 8711
rect 85640 8711 85656 8728
rect 86086 8728 86674 8744
rect 86086 8711 86102 8728
rect 85640 8694 85842 8711
rect 84882 8656 85842 8694
rect 85900 8694 86102 8711
rect 86658 8711 86674 8728
rect 87104 8728 87692 8744
rect 87104 8711 87120 8728
rect 86658 8694 86860 8711
rect 85900 8656 86860 8694
rect 86918 8694 87120 8711
rect 87676 8711 87692 8728
rect 87676 8694 87878 8711
rect 86918 8656 87878 8694
rect 55812 8482 56772 8520
rect 55812 8465 56014 8482
rect 55998 8448 56014 8465
rect 56570 8465 56772 8482
rect 56830 8482 57790 8520
rect 56830 8465 57032 8482
rect 56570 8448 56586 8465
rect 55998 8432 56586 8448
rect 57016 8448 57032 8465
rect 57588 8465 57790 8482
rect 57848 8482 58808 8520
rect 57848 8465 58050 8482
rect 57588 8448 57604 8465
rect 57016 8432 57604 8448
rect 55998 8374 56586 8390
rect 55998 8357 56014 8374
rect 55812 8340 56014 8357
rect 56570 8357 56586 8374
rect 58034 8448 58050 8465
rect 58606 8465 58808 8482
rect 58866 8482 59826 8520
rect 58866 8465 59068 8482
rect 58606 8448 58622 8465
rect 58034 8432 58622 8448
rect 57016 8374 57604 8390
rect 57016 8357 57032 8374
rect 56570 8340 56772 8357
rect 55812 8302 56772 8340
rect 56830 8340 57032 8357
rect 57588 8357 57604 8374
rect 59052 8448 59068 8465
rect 59624 8465 59826 8482
rect 59884 8482 60844 8520
rect 59884 8465 60086 8482
rect 59624 8448 59640 8465
rect 59052 8432 59640 8448
rect 58034 8374 58622 8390
rect 58034 8357 58050 8374
rect 57588 8340 57790 8357
rect 56830 8302 57790 8340
rect 57848 8340 58050 8357
rect 58606 8357 58622 8374
rect 60070 8448 60086 8465
rect 60642 8465 60844 8482
rect 60902 8482 61862 8520
rect 60902 8465 61104 8482
rect 60642 8448 60658 8465
rect 60070 8432 60658 8448
rect 59052 8374 59640 8390
rect 59052 8357 59068 8374
rect 58606 8340 58808 8357
rect 57848 8302 58808 8340
rect 58866 8340 59068 8357
rect 59624 8357 59640 8374
rect 61088 8448 61104 8465
rect 61660 8465 61862 8482
rect 61920 8482 62880 8520
rect 61920 8465 62122 8482
rect 61660 8448 61676 8465
rect 61088 8432 61676 8448
rect 60070 8374 60658 8390
rect 60070 8357 60086 8374
rect 59624 8340 59826 8357
rect 58866 8302 59826 8340
rect 59884 8340 60086 8357
rect 60642 8357 60658 8374
rect 62106 8448 62122 8465
rect 62678 8465 62880 8482
rect 62938 8482 63898 8520
rect 62938 8465 63140 8482
rect 62678 8448 62694 8465
rect 62106 8432 62694 8448
rect 61088 8374 61676 8390
rect 61088 8357 61104 8374
rect 60642 8340 60844 8357
rect 59884 8302 60844 8340
rect 60902 8340 61104 8357
rect 61660 8357 61676 8374
rect 63124 8448 63140 8465
rect 63696 8465 63898 8482
rect 63956 8482 64916 8520
rect 63956 8465 64158 8482
rect 63696 8448 63712 8465
rect 63124 8432 63712 8448
rect 62106 8374 62694 8390
rect 62106 8357 62122 8374
rect 61660 8340 61862 8357
rect 60902 8302 61862 8340
rect 61920 8340 62122 8357
rect 62678 8357 62694 8374
rect 64142 8448 64158 8465
rect 64714 8465 64916 8482
rect 64714 8448 64730 8465
rect 64142 8432 64730 8448
rect 63124 8374 63712 8390
rect 63124 8357 63140 8374
rect 62678 8340 62880 8357
rect 61920 8302 62880 8340
rect 62938 8340 63140 8357
rect 63696 8357 63712 8374
rect 64142 8374 64730 8390
rect 64142 8357 64158 8374
rect 63696 8340 63898 8357
rect 62938 8302 63898 8340
rect 63956 8340 64158 8357
rect 64714 8357 64730 8374
rect 64714 8340 64916 8357
rect 63956 8302 64916 8340
rect 67576 8018 68536 8056
rect 67576 8001 67778 8018
rect 67762 7984 67778 8001
rect 68334 8001 68536 8018
rect 68594 8018 69554 8056
rect 68594 8001 68796 8018
rect 68334 7984 68350 8001
rect 67762 7968 68350 7984
rect 68780 7984 68796 8001
rect 69352 8001 69554 8018
rect 69612 8018 70572 8056
rect 69612 8001 69814 8018
rect 69352 7984 69368 8001
rect 68780 7968 69368 7984
rect 69798 7984 69814 8001
rect 70370 8001 70572 8018
rect 70630 8018 71590 8056
rect 70630 8001 70832 8018
rect 70370 7984 70386 8001
rect 69798 7968 70386 7984
rect 70816 7984 70832 8001
rect 71388 8001 71590 8018
rect 71648 8018 72608 8056
rect 71648 8001 71850 8018
rect 71388 7984 71404 8001
rect 70816 7968 71404 7984
rect 71834 7984 71850 8001
rect 72406 8001 72608 8018
rect 72666 8018 73626 8056
rect 72666 8001 72868 8018
rect 72406 7984 72422 8001
rect 71834 7968 72422 7984
rect 72852 7984 72868 8001
rect 73424 8001 73626 8018
rect 73684 8018 74644 8056
rect 73684 8001 73886 8018
rect 73424 7984 73440 8001
rect 72852 7968 73440 7984
rect 73870 7984 73886 8001
rect 74442 8001 74644 8018
rect 74702 8018 75662 8056
rect 74702 8001 74904 8018
rect 74442 7984 74458 8001
rect 73870 7968 74458 7984
rect 74888 7984 74904 8001
rect 75460 8001 75662 8018
rect 75720 8018 76680 8056
rect 75720 8001 75922 8018
rect 75460 7984 75476 8001
rect 74888 7968 75476 7984
rect 75906 7984 75922 8001
rect 76478 8001 76680 8018
rect 76738 8018 77698 8056
rect 76738 8001 76940 8018
rect 76478 7984 76494 8001
rect 75906 7968 76494 7984
rect 76924 7984 76940 8001
rect 77496 8001 77698 8018
rect 77756 8018 78716 8056
rect 77756 8001 77958 8018
rect 77496 7984 77512 8001
rect 76924 7968 77512 7984
rect 77942 7984 77958 8001
rect 78514 8001 78716 8018
rect 78774 8018 79734 8056
rect 78774 8001 78976 8018
rect 78514 7984 78530 8001
rect 77942 7968 78530 7984
rect 78960 7984 78976 8001
rect 79532 8001 79734 8018
rect 79792 8018 80752 8056
rect 79792 8001 79994 8018
rect 79532 7984 79548 8001
rect 78960 7968 79548 7984
rect 79978 7984 79994 8001
rect 80550 8001 80752 8018
rect 80810 8018 81770 8056
rect 80810 8001 81012 8018
rect 80550 7984 80566 8001
rect 79978 7968 80566 7984
rect 80996 7984 81012 8001
rect 81568 8001 81770 8018
rect 81828 8018 82788 8056
rect 81828 8001 82030 8018
rect 81568 7984 81584 8001
rect 80996 7968 81584 7984
rect 82014 7984 82030 8001
rect 82586 8001 82788 8018
rect 82846 8018 83806 8056
rect 82846 8001 83048 8018
rect 82586 7984 82602 8001
rect 82014 7968 82602 7984
rect 83032 7984 83048 8001
rect 83604 8001 83806 8018
rect 83864 8018 84824 8056
rect 83864 8001 84066 8018
rect 83604 7984 83620 8001
rect 83032 7968 83620 7984
rect 84050 7984 84066 8001
rect 84622 8001 84824 8018
rect 84882 8018 85842 8056
rect 84882 8001 85084 8018
rect 84622 7984 84638 8001
rect 84050 7968 84638 7984
rect 85068 7984 85084 8001
rect 85640 8001 85842 8018
rect 85900 8018 86860 8056
rect 85900 8001 86102 8018
rect 85640 7984 85656 8001
rect 85068 7968 85656 7984
rect 86086 7984 86102 8001
rect 86658 8001 86860 8018
rect 86918 8018 87878 8056
rect 86918 8001 87120 8018
rect 86658 7984 86674 8001
rect 86086 7968 86674 7984
rect 87104 7984 87120 8001
rect 87676 8001 87878 8018
rect 87676 7984 87692 8001
rect 87104 7968 87692 7984
rect 55812 7664 56772 7702
rect 55812 7647 56014 7664
rect 55998 7630 56014 7647
rect 56570 7647 56772 7664
rect 56830 7664 57790 7702
rect 56830 7647 57032 7664
rect 56570 7630 56586 7647
rect 55998 7614 56586 7630
rect 57016 7630 57032 7647
rect 57588 7647 57790 7664
rect 57848 7664 58808 7702
rect 57848 7647 58050 7664
rect 57588 7630 57604 7647
rect 57016 7614 57604 7630
rect 58034 7630 58050 7647
rect 58606 7647 58808 7664
rect 58866 7664 59826 7702
rect 58866 7647 59068 7664
rect 58606 7630 58622 7647
rect 58034 7614 58622 7630
rect 59052 7630 59068 7647
rect 59624 7647 59826 7664
rect 59884 7664 60844 7702
rect 59884 7647 60086 7664
rect 59624 7630 59640 7647
rect 59052 7614 59640 7630
rect 60070 7630 60086 7647
rect 60642 7647 60844 7664
rect 60902 7664 61862 7702
rect 60902 7647 61104 7664
rect 60642 7630 60658 7647
rect 60070 7614 60658 7630
rect 61088 7630 61104 7647
rect 61660 7647 61862 7664
rect 61920 7664 62880 7702
rect 61920 7647 62122 7664
rect 61660 7630 61676 7647
rect 61088 7614 61676 7630
rect 62106 7630 62122 7647
rect 62678 7647 62880 7664
rect 62938 7664 63898 7702
rect 62938 7647 63140 7664
rect 62678 7630 62694 7647
rect 62106 7614 62694 7630
rect 63124 7630 63140 7647
rect 63696 7647 63898 7664
rect 63956 7664 64916 7702
rect 63956 7647 64158 7664
rect 63696 7630 63712 7647
rect 63124 7614 63712 7630
rect 64142 7630 64158 7647
rect 64714 7647 64916 7664
rect 64714 7630 64730 7647
rect 64142 7614 64730 7630
rect 67762 7494 68350 7510
rect 67762 7477 67778 7494
rect 67576 7460 67778 7477
rect 68334 7477 68350 7494
rect 68780 7494 69368 7510
rect 68780 7477 68796 7494
rect 68334 7460 68536 7477
rect 67576 7422 68536 7460
rect 68594 7460 68796 7477
rect 69352 7477 69368 7494
rect 69798 7494 70386 7510
rect 69798 7477 69814 7494
rect 69352 7460 69554 7477
rect 68594 7422 69554 7460
rect 69612 7460 69814 7477
rect 70370 7477 70386 7494
rect 70816 7494 71404 7510
rect 70816 7477 70832 7494
rect 70370 7460 70572 7477
rect 69612 7422 70572 7460
rect 70630 7460 70832 7477
rect 71388 7477 71404 7494
rect 71834 7494 72422 7510
rect 71834 7477 71850 7494
rect 71388 7460 71590 7477
rect 70630 7422 71590 7460
rect 71648 7460 71850 7477
rect 72406 7477 72422 7494
rect 72852 7494 73440 7510
rect 72852 7477 72868 7494
rect 72406 7460 72608 7477
rect 71648 7422 72608 7460
rect 72666 7460 72868 7477
rect 73424 7477 73440 7494
rect 73870 7494 74458 7510
rect 73870 7477 73886 7494
rect 73424 7460 73626 7477
rect 72666 7422 73626 7460
rect 73684 7460 73886 7477
rect 74442 7477 74458 7494
rect 74888 7494 75476 7510
rect 74888 7477 74904 7494
rect 74442 7460 74644 7477
rect 73684 7422 74644 7460
rect 74702 7460 74904 7477
rect 75460 7477 75476 7494
rect 75906 7494 76494 7510
rect 75906 7477 75922 7494
rect 75460 7460 75662 7477
rect 74702 7422 75662 7460
rect 75720 7460 75922 7477
rect 76478 7477 76494 7494
rect 76924 7494 77512 7510
rect 76924 7477 76940 7494
rect 76478 7460 76680 7477
rect 75720 7422 76680 7460
rect 76738 7460 76940 7477
rect 77496 7477 77512 7494
rect 77942 7494 78530 7510
rect 77942 7477 77958 7494
rect 77496 7460 77698 7477
rect 76738 7422 77698 7460
rect 77756 7460 77958 7477
rect 78514 7477 78530 7494
rect 78960 7494 79548 7510
rect 78960 7477 78976 7494
rect 78514 7460 78716 7477
rect 77756 7422 78716 7460
rect 78774 7460 78976 7477
rect 79532 7477 79548 7494
rect 79978 7494 80566 7510
rect 79978 7477 79994 7494
rect 79532 7460 79734 7477
rect 78774 7422 79734 7460
rect 79792 7460 79994 7477
rect 80550 7477 80566 7494
rect 80996 7494 81584 7510
rect 80996 7477 81012 7494
rect 80550 7460 80752 7477
rect 79792 7422 80752 7460
rect 80810 7460 81012 7477
rect 81568 7477 81584 7494
rect 82014 7494 82602 7510
rect 82014 7477 82030 7494
rect 81568 7460 81770 7477
rect 80810 7422 81770 7460
rect 81828 7460 82030 7477
rect 82586 7477 82602 7494
rect 83032 7494 83620 7510
rect 83032 7477 83048 7494
rect 82586 7460 82788 7477
rect 81828 7422 82788 7460
rect 82846 7460 83048 7477
rect 83604 7477 83620 7494
rect 84050 7494 84638 7510
rect 84050 7477 84066 7494
rect 83604 7460 83806 7477
rect 82846 7422 83806 7460
rect 83864 7460 84066 7477
rect 84622 7477 84638 7494
rect 85068 7494 85656 7510
rect 85068 7477 85084 7494
rect 84622 7460 84824 7477
rect 83864 7422 84824 7460
rect 84882 7460 85084 7477
rect 85640 7477 85656 7494
rect 86086 7494 86674 7510
rect 86086 7477 86102 7494
rect 85640 7460 85842 7477
rect 84882 7422 85842 7460
rect 85900 7460 86102 7477
rect 86658 7477 86674 7494
rect 87104 7494 87692 7510
rect 87104 7477 87120 7494
rect 86658 7460 86860 7477
rect 85900 7422 86860 7460
rect 86918 7460 87120 7477
rect 87676 7477 87692 7494
rect 87676 7460 87878 7477
rect 86918 7422 87878 7460
rect 62698 6990 62806 7006
rect 62698 6973 62714 6990
rect 62672 6956 62714 6973
rect 62790 6973 62806 6990
rect 62916 6990 63024 7006
rect 62916 6973 62932 6990
rect 62790 6956 62832 6973
rect 62672 6918 62832 6956
rect 62890 6956 62932 6973
rect 63008 6973 63024 6990
rect 63134 6990 63242 7006
rect 63134 6973 63150 6990
rect 63008 6956 63050 6973
rect 62890 6918 63050 6956
rect 63108 6956 63150 6973
rect 63226 6973 63242 6990
rect 63352 6990 63460 7006
rect 63352 6973 63368 6990
rect 63226 6956 63268 6973
rect 63108 6918 63268 6956
rect 63326 6956 63368 6973
rect 63444 6973 63460 6990
rect 63570 6990 63678 7006
rect 63570 6973 63586 6990
rect 63444 6956 63486 6973
rect 63326 6918 63486 6956
rect 63544 6956 63586 6973
rect 63662 6973 63678 6990
rect 63788 6990 63896 7006
rect 63788 6973 63804 6990
rect 63662 6956 63704 6973
rect 63544 6918 63704 6956
rect 63762 6956 63804 6973
rect 63880 6973 63896 6990
rect 64006 6990 64114 7006
rect 64006 6973 64022 6990
rect 63880 6956 63922 6973
rect 63762 6918 63922 6956
rect 63980 6956 64022 6973
rect 64098 6973 64114 6990
rect 64224 6990 64332 7006
rect 64224 6973 64240 6990
rect 64098 6956 64140 6973
rect 63980 6918 64140 6956
rect 64198 6956 64240 6973
rect 64316 6973 64332 6990
rect 64442 6990 64550 7006
rect 64442 6973 64458 6990
rect 64316 6956 64358 6973
rect 64198 6918 64358 6956
rect 64416 6956 64458 6973
rect 64534 6973 64550 6990
rect 64660 6990 64768 7006
rect 64660 6973 64676 6990
rect 64534 6956 64576 6973
rect 64416 6918 64576 6956
rect 64634 6956 64676 6973
rect 64752 6973 64768 6990
rect 64752 6956 64794 6973
rect 64634 6918 64794 6956
rect 67576 6784 68536 6822
rect 67576 6767 67778 6784
rect 67762 6750 67778 6767
rect 68334 6767 68536 6784
rect 68594 6784 69554 6822
rect 68594 6767 68796 6784
rect 68334 6750 68350 6767
rect 67762 6734 68350 6750
rect 68780 6750 68796 6767
rect 69352 6767 69554 6784
rect 69612 6784 70572 6822
rect 69612 6767 69814 6784
rect 69352 6750 69368 6767
rect 68780 6734 69368 6750
rect 69798 6750 69814 6767
rect 70370 6767 70572 6784
rect 70630 6784 71590 6822
rect 70630 6767 70832 6784
rect 70370 6750 70386 6767
rect 69798 6734 70386 6750
rect 70816 6750 70832 6767
rect 71388 6767 71590 6784
rect 71648 6784 72608 6822
rect 71648 6767 71850 6784
rect 71388 6750 71404 6767
rect 70816 6734 71404 6750
rect 71834 6750 71850 6767
rect 72406 6767 72608 6784
rect 72666 6784 73626 6822
rect 72666 6767 72868 6784
rect 72406 6750 72422 6767
rect 71834 6734 72422 6750
rect 72852 6750 72868 6767
rect 73424 6767 73626 6784
rect 73684 6784 74644 6822
rect 73684 6767 73886 6784
rect 73424 6750 73440 6767
rect 72852 6734 73440 6750
rect 73870 6750 73886 6767
rect 74442 6767 74644 6784
rect 74702 6784 75662 6822
rect 74702 6767 74904 6784
rect 74442 6750 74458 6767
rect 73870 6734 74458 6750
rect 74888 6750 74904 6767
rect 75460 6767 75662 6784
rect 75720 6784 76680 6822
rect 75720 6767 75922 6784
rect 75460 6750 75476 6767
rect 74888 6734 75476 6750
rect 75906 6750 75922 6767
rect 76478 6767 76680 6784
rect 76738 6784 77698 6822
rect 76738 6767 76940 6784
rect 76478 6750 76494 6767
rect 75906 6734 76494 6750
rect 76924 6750 76940 6767
rect 77496 6767 77698 6784
rect 77756 6784 78716 6822
rect 77756 6767 77958 6784
rect 77496 6750 77512 6767
rect 76924 6734 77512 6750
rect 77942 6750 77958 6767
rect 78514 6767 78716 6784
rect 78774 6784 79734 6822
rect 78774 6767 78976 6784
rect 78514 6750 78530 6767
rect 77942 6734 78530 6750
rect 78960 6750 78976 6767
rect 79532 6767 79734 6784
rect 79792 6784 80752 6822
rect 79792 6767 79994 6784
rect 79532 6750 79548 6767
rect 78960 6734 79548 6750
rect 79978 6750 79994 6767
rect 80550 6767 80752 6784
rect 80810 6784 81770 6822
rect 80810 6767 81012 6784
rect 80550 6750 80566 6767
rect 79978 6734 80566 6750
rect 80996 6750 81012 6767
rect 81568 6767 81770 6784
rect 81828 6784 82788 6822
rect 81828 6767 82030 6784
rect 81568 6750 81584 6767
rect 80996 6734 81584 6750
rect 82014 6750 82030 6767
rect 82586 6767 82788 6784
rect 82846 6784 83806 6822
rect 82846 6767 83048 6784
rect 82586 6750 82602 6767
rect 82014 6734 82602 6750
rect 83032 6750 83048 6767
rect 83604 6767 83806 6784
rect 83864 6784 84824 6822
rect 83864 6767 84066 6784
rect 83604 6750 83620 6767
rect 83032 6734 83620 6750
rect 84050 6750 84066 6767
rect 84622 6767 84824 6784
rect 84882 6784 85842 6822
rect 84882 6767 85084 6784
rect 84622 6750 84638 6767
rect 84050 6734 84638 6750
rect 85068 6750 85084 6767
rect 85640 6767 85842 6784
rect 85900 6784 86860 6822
rect 85900 6767 86102 6784
rect 85640 6750 85656 6767
rect 85068 6734 85656 6750
rect 86086 6750 86102 6767
rect 86658 6767 86860 6784
rect 86918 6784 87878 6822
rect 86918 6767 87120 6784
rect 86658 6750 86674 6767
rect 86086 6734 86674 6750
rect 87104 6750 87120 6767
rect 87676 6767 87878 6784
rect 87676 6750 87692 6767
rect 87104 6734 87692 6750
rect 62672 6680 62832 6718
rect 62672 6663 62714 6680
rect 62698 6646 62714 6663
rect 62790 6663 62832 6680
rect 62890 6680 63050 6718
rect 62890 6663 62932 6680
rect 62790 6646 62806 6663
rect 62698 6630 62806 6646
rect 62916 6646 62932 6663
rect 63008 6663 63050 6680
rect 63108 6680 63268 6718
rect 63108 6663 63150 6680
rect 63008 6646 63024 6663
rect 62916 6630 63024 6646
rect 63134 6646 63150 6663
rect 63226 6663 63268 6680
rect 63326 6680 63486 6718
rect 63326 6663 63368 6680
rect 63226 6646 63242 6663
rect 63134 6630 63242 6646
rect 63352 6646 63368 6663
rect 63444 6663 63486 6680
rect 63544 6680 63704 6718
rect 63544 6663 63586 6680
rect 63444 6646 63460 6663
rect 63352 6630 63460 6646
rect 63570 6646 63586 6663
rect 63662 6663 63704 6680
rect 63762 6680 63922 6718
rect 63762 6663 63804 6680
rect 63662 6646 63678 6663
rect 63570 6630 63678 6646
rect 63788 6646 63804 6663
rect 63880 6663 63922 6680
rect 63980 6680 64140 6718
rect 63980 6663 64022 6680
rect 63880 6646 63896 6663
rect 63788 6630 63896 6646
rect 64006 6646 64022 6663
rect 64098 6663 64140 6680
rect 64198 6680 64358 6718
rect 64198 6663 64240 6680
rect 64098 6646 64114 6663
rect 64006 6630 64114 6646
rect 64224 6646 64240 6663
rect 64316 6663 64358 6680
rect 64416 6680 64576 6718
rect 64416 6663 64458 6680
rect 64316 6646 64332 6663
rect 64224 6630 64332 6646
rect 64442 6646 64458 6663
rect 64534 6663 64576 6680
rect 64634 6680 64794 6718
rect 64634 6663 64676 6680
rect 64534 6646 64550 6663
rect 64442 6630 64550 6646
rect 64660 6646 64676 6663
rect 64752 6663 64794 6680
rect 64752 6646 64768 6663
rect 64660 6630 64768 6646
rect 67762 6260 68350 6276
rect 67762 6243 67778 6260
rect 67576 6226 67778 6243
rect 68334 6243 68350 6260
rect 68780 6260 69368 6276
rect 68780 6243 68796 6260
rect 68334 6226 68536 6243
rect 67576 6188 68536 6226
rect 68594 6226 68796 6243
rect 69352 6243 69368 6260
rect 69798 6260 70386 6276
rect 69798 6243 69814 6260
rect 69352 6226 69554 6243
rect 68594 6188 69554 6226
rect 69612 6226 69814 6243
rect 70370 6243 70386 6260
rect 70816 6260 71404 6276
rect 70816 6243 70832 6260
rect 70370 6226 70572 6243
rect 69612 6188 70572 6226
rect 70630 6226 70832 6243
rect 71388 6243 71404 6260
rect 71834 6260 72422 6276
rect 71834 6243 71850 6260
rect 71388 6226 71590 6243
rect 70630 6188 71590 6226
rect 71648 6226 71850 6243
rect 72406 6243 72422 6260
rect 72852 6260 73440 6276
rect 72852 6243 72868 6260
rect 72406 6226 72608 6243
rect 71648 6188 72608 6226
rect 72666 6226 72868 6243
rect 73424 6243 73440 6260
rect 73870 6260 74458 6276
rect 73870 6243 73886 6260
rect 73424 6226 73626 6243
rect 72666 6188 73626 6226
rect 73684 6226 73886 6243
rect 74442 6243 74458 6260
rect 74888 6260 75476 6276
rect 74888 6243 74904 6260
rect 74442 6226 74644 6243
rect 73684 6188 74644 6226
rect 74702 6226 74904 6243
rect 75460 6243 75476 6260
rect 75906 6260 76494 6276
rect 75906 6243 75922 6260
rect 75460 6226 75662 6243
rect 74702 6188 75662 6226
rect 75720 6226 75922 6243
rect 76478 6243 76494 6260
rect 76924 6260 77512 6276
rect 76924 6243 76940 6260
rect 76478 6226 76680 6243
rect 75720 6188 76680 6226
rect 76738 6226 76940 6243
rect 77496 6243 77512 6260
rect 77942 6260 78530 6276
rect 77942 6243 77958 6260
rect 77496 6226 77698 6243
rect 76738 6188 77698 6226
rect 77756 6226 77958 6243
rect 78514 6243 78530 6260
rect 78960 6260 79548 6276
rect 78960 6243 78976 6260
rect 78514 6226 78716 6243
rect 77756 6188 78716 6226
rect 78774 6226 78976 6243
rect 79532 6243 79548 6260
rect 79978 6260 80566 6276
rect 79978 6243 79994 6260
rect 79532 6226 79734 6243
rect 78774 6188 79734 6226
rect 79792 6226 79994 6243
rect 80550 6243 80566 6260
rect 80996 6260 81584 6276
rect 80996 6243 81012 6260
rect 80550 6226 80752 6243
rect 79792 6188 80752 6226
rect 80810 6226 81012 6243
rect 81568 6243 81584 6260
rect 82014 6260 82602 6276
rect 82014 6243 82030 6260
rect 81568 6226 81770 6243
rect 80810 6188 81770 6226
rect 81828 6226 82030 6243
rect 82586 6243 82602 6260
rect 83032 6260 83620 6276
rect 83032 6243 83048 6260
rect 82586 6226 82788 6243
rect 81828 6188 82788 6226
rect 82846 6226 83048 6243
rect 83604 6243 83620 6260
rect 84050 6260 84638 6276
rect 84050 6243 84066 6260
rect 83604 6226 83806 6243
rect 82846 6188 83806 6226
rect 83864 6226 84066 6243
rect 84622 6243 84638 6260
rect 85068 6260 85656 6276
rect 85068 6243 85084 6260
rect 84622 6226 84824 6243
rect 83864 6188 84824 6226
rect 84882 6226 85084 6243
rect 85640 6243 85656 6260
rect 86086 6260 86674 6276
rect 86086 6243 86102 6260
rect 85640 6226 85842 6243
rect 84882 6188 85842 6226
rect 85900 6226 86102 6243
rect 86658 6243 86674 6260
rect 87104 6260 87692 6276
rect 87104 6243 87120 6260
rect 86658 6226 86860 6243
rect 85900 6188 86860 6226
rect 86918 6226 87120 6243
rect 87676 6243 87692 6260
rect 87676 6226 87878 6243
rect 86918 6188 87878 6226
rect 62698 6158 62806 6174
rect 62698 6141 62714 6158
rect 62672 6124 62714 6141
rect 62790 6141 62806 6158
rect 62916 6158 63024 6174
rect 62916 6141 62932 6158
rect 62790 6124 62832 6141
rect 62672 6086 62832 6124
rect 62890 6124 62932 6141
rect 63008 6141 63024 6158
rect 63134 6158 63242 6174
rect 63134 6141 63150 6158
rect 63008 6124 63050 6141
rect 62890 6086 63050 6124
rect 63108 6124 63150 6141
rect 63226 6141 63242 6158
rect 63352 6158 63460 6174
rect 63352 6141 63368 6158
rect 63226 6124 63268 6141
rect 63108 6086 63268 6124
rect 63326 6124 63368 6141
rect 63444 6141 63460 6158
rect 63570 6158 63678 6174
rect 63570 6141 63586 6158
rect 63444 6124 63486 6141
rect 63326 6086 63486 6124
rect 63544 6124 63586 6141
rect 63662 6141 63678 6158
rect 63788 6158 63896 6174
rect 63788 6141 63804 6158
rect 63662 6124 63704 6141
rect 63544 6086 63704 6124
rect 63762 6124 63804 6141
rect 63880 6141 63896 6158
rect 64006 6158 64114 6174
rect 64006 6141 64022 6158
rect 63880 6124 63922 6141
rect 63762 6086 63922 6124
rect 63980 6124 64022 6141
rect 64098 6141 64114 6158
rect 64224 6158 64332 6174
rect 64224 6141 64240 6158
rect 64098 6124 64140 6141
rect 63980 6086 64140 6124
rect 64198 6124 64240 6141
rect 64316 6141 64332 6158
rect 64442 6158 64550 6174
rect 64442 6141 64458 6158
rect 64316 6124 64358 6141
rect 64198 6086 64358 6124
rect 64416 6124 64458 6141
rect 64534 6141 64550 6158
rect 64660 6158 64768 6174
rect 64660 6141 64676 6158
rect 64534 6124 64576 6141
rect 64416 6086 64576 6124
rect 64634 6124 64676 6141
rect 64752 6141 64768 6158
rect 64752 6124 64794 6141
rect 64634 6086 64794 6124
rect 62672 5848 62832 5886
rect 62672 5831 62714 5848
rect 62698 5814 62714 5831
rect 62790 5831 62832 5848
rect 62890 5848 63050 5886
rect 62890 5831 62932 5848
rect 62790 5814 62806 5831
rect 62698 5798 62806 5814
rect 62916 5814 62932 5831
rect 63008 5831 63050 5848
rect 63108 5848 63268 5886
rect 63108 5831 63150 5848
rect 63008 5814 63024 5831
rect 62916 5798 63024 5814
rect 63134 5814 63150 5831
rect 63226 5831 63268 5848
rect 63326 5848 63486 5886
rect 63326 5831 63368 5848
rect 63226 5814 63242 5831
rect 63134 5798 63242 5814
rect 63352 5814 63368 5831
rect 63444 5831 63486 5848
rect 63544 5848 63704 5886
rect 63544 5831 63586 5848
rect 63444 5814 63460 5831
rect 63352 5798 63460 5814
rect 63570 5814 63586 5831
rect 63662 5831 63704 5848
rect 63762 5848 63922 5886
rect 63762 5831 63804 5848
rect 63662 5814 63678 5831
rect 63570 5798 63678 5814
rect 63788 5814 63804 5831
rect 63880 5831 63922 5848
rect 63980 5848 64140 5886
rect 63980 5831 64022 5848
rect 63880 5814 63896 5831
rect 63788 5798 63896 5814
rect 64006 5814 64022 5831
rect 64098 5831 64140 5848
rect 64198 5848 64358 5886
rect 64198 5831 64240 5848
rect 64098 5814 64114 5831
rect 64006 5798 64114 5814
rect 64224 5814 64240 5831
rect 64316 5831 64358 5848
rect 64416 5848 64576 5886
rect 64416 5831 64458 5848
rect 64316 5814 64332 5831
rect 64224 5798 64332 5814
rect 64442 5814 64458 5831
rect 64534 5831 64576 5848
rect 64634 5848 64794 5886
rect 64634 5831 64676 5848
rect 64534 5814 64550 5831
rect 64442 5798 64550 5814
rect 64660 5814 64676 5831
rect 64752 5831 64794 5848
rect 64752 5814 64768 5831
rect 64660 5798 64768 5814
rect 67576 5550 68536 5588
rect 67576 5533 67778 5550
rect 67762 5516 67778 5533
rect 68334 5533 68536 5550
rect 68594 5550 69554 5588
rect 68594 5533 68796 5550
rect 68334 5516 68350 5533
rect 67762 5500 68350 5516
rect 68780 5516 68796 5533
rect 69352 5533 69554 5550
rect 69612 5550 70572 5588
rect 69612 5533 69814 5550
rect 69352 5516 69368 5533
rect 68780 5500 69368 5516
rect 69798 5516 69814 5533
rect 70370 5533 70572 5550
rect 70630 5550 71590 5588
rect 70630 5533 70832 5550
rect 70370 5516 70386 5533
rect 69798 5500 70386 5516
rect 70816 5516 70832 5533
rect 71388 5533 71590 5550
rect 71648 5550 72608 5588
rect 71648 5533 71850 5550
rect 71388 5516 71404 5533
rect 70816 5500 71404 5516
rect 71834 5516 71850 5533
rect 72406 5533 72608 5550
rect 72666 5550 73626 5588
rect 72666 5533 72868 5550
rect 72406 5516 72422 5533
rect 71834 5500 72422 5516
rect 72852 5516 72868 5533
rect 73424 5533 73626 5550
rect 73684 5550 74644 5588
rect 73684 5533 73886 5550
rect 73424 5516 73440 5533
rect 72852 5500 73440 5516
rect 73870 5516 73886 5533
rect 74442 5533 74644 5550
rect 74702 5550 75662 5588
rect 74702 5533 74904 5550
rect 74442 5516 74458 5533
rect 73870 5500 74458 5516
rect 74888 5516 74904 5533
rect 75460 5533 75662 5550
rect 75720 5550 76680 5588
rect 75720 5533 75922 5550
rect 75460 5516 75476 5533
rect 74888 5500 75476 5516
rect 75906 5516 75922 5533
rect 76478 5533 76680 5550
rect 76738 5550 77698 5588
rect 76738 5533 76940 5550
rect 76478 5516 76494 5533
rect 75906 5500 76494 5516
rect 76924 5516 76940 5533
rect 77496 5533 77698 5550
rect 77756 5550 78716 5588
rect 77756 5533 77958 5550
rect 77496 5516 77512 5533
rect 76924 5500 77512 5516
rect 77942 5516 77958 5533
rect 78514 5533 78716 5550
rect 78774 5550 79734 5588
rect 78774 5533 78976 5550
rect 78514 5516 78530 5533
rect 77942 5500 78530 5516
rect 78960 5516 78976 5533
rect 79532 5533 79734 5550
rect 79792 5550 80752 5588
rect 79792 5533 79994 5550
rect 79532 5516 79548 5533
rect 78960 5500 79548 5516
rect 79978 5516 79994 5533
rect 80550 5533 80752 5550
rect 80810 5550 81770 5588
rect 80810 5533 81012 5550
rect 80550 5516 80566 5533
rect 79978 5500 80566 5516
rect 80996 5516 81012 5533
rect 81568 5533 81770 5550
rect 81828 5550 82788 5588
rect 81828 5533 82030 5550
rect 81568 5516 81584 5533
rect 80996 5500 81584 5516
rect 82014 5516 82030 5533
rect 82586 5533 82788 5550
rect 82846 5550 83806 5588
rect 82846 5533 83048 5550
rect 82586 5516 82602 5533
rect 82014 5500 82602 5516
rect 83032 5516 83048 5533
rect 83604 5533 83806 5550
rect 83864 5550 84824 5588
rect 83864 5533 84066 5550
rect 83604 5516 83620 5533
rect 83032 5500 83620 5516
rect 84050 5516 84066 5533
rect 84622 5533 84824 5550
rect 84882 5550 85842 5588
rect 84882 5533 85084 5550
rect 84622 5516 84638 5533
rect 84050 5500 84638 5516
rect 85068 5516 85084 5533
rect 85640 5533 85842 5550
rect 85900 5550 86860 5588
rect 85900 5533 86102 5550
rect 85640 5516 85656 5533
rect 85068 5500 85656 5516
rect 86086 5516 86102 5533
rect 86658 5533 86860 5550
rect 86918 5550 87878 5588
rect 86918 5533 87120 5550
rect 86658 5516 86674 5533
rect 86086 5500 86674 5516
rect 87104 5516 87120 5533
rect 87676 5533 87878 5550
rect 87676 5516 87692 5533
rect 87104 5500 87692 5516
rect 67762 5028 68350 5044
rect 67762 5011 67778 5028
rect 67576 4994 67778 5011
rect 68334 5011 68350 5028
rect 68780 5028 69368 5044
rect 68780 5011 68796 5028
rect 68334 4994 68536 5011
rect 67576 4956 68536 4994
rect 68594 4994 68796 5011
rect 69352 5011 69368 5028
rect 69798 5028 70386 5044
rect 69798 5011 69814 5028
rect 69352 4994 69554 5011
rect 68594 4956 69554 4994
rect 69612 4994 69814 5011
rect 70370 5011 70386 5028
rect 70816 5028 71404 5044
rect 70816 5011 70832 5028
rect 70370 4994 70572 5011
rect 69612 4956 70572 4994
rect 70630 4994 70832 5011
rect 71388 5011 71404 5028
rect 71834 5028 72422 5044
rect 71834 5011 71850 5028
rect 71388 4994 71590 5011
rect 70630 4956 71590 4994
rect 71648 4994 71850 5011
rect 72406 5011 72422 5028
rect 72852 5028 73440 5044
rect 72852 5011 72868 5028
rect 72406 4994 72608 5011
rect 71648 4956 72608 4994
rect 72666 4994 72868 5011
rect 73424 5011 73440 5028
rect 73870 5028 74458 5044
rect 73870 5011 73886 5028
rect 73424 4994 73626 5011
rect 72666 4956 73626 4994
rect 73684 4994 73886 5011
rect 74442 5011 74458 5028
rect 74888 5028 75476 5044
rect 74888 5011 74904 5028
rect 74442 4994 74644 5011
rect 73684 4956 74644 4994
rect 74702 4994 74904 5011
rect 75460 5011 75476 5028
rect 75906 5028 76494 5044
rect 75906 5011 75922 5028
rect 75460 4994 75662 5011
rect 74702 4956 75662 4994
rect 75720 4994 75922 5011
rect 76478 5011 76494 5028
rect 76924 5028 77512 5044
rect 76924 5011 76940 5028
rect 76478 4994 76680 5011
rect 75720 4956 76680 4994
rect 76738 4994 76940 5011
rect 77496 5011 77512 5028
rect 77942 5028 78530 5044
rect 77942 5011 77958 5028
rect 77496 4994 77698 5011
rect 76738 4956 77698 4994
rect 77756 4994 77958 5011
rect 78514 5011 78530 5028
rect 78960 5028 79548 5044
rect 78960 5011 78976 5028
rect 78514 4994 78716 5011
rect 77756 4956 78716 4994
rect 78774 4994 78976 5011
rect 79532 5011 79548 5028
rect 79978 5028 80566 5044
rect 79978 5011 79994 5028
rect 79532 4994 79734 5011
rect 78774 4956 79734 4994
rect 79792 4994 79994 5011
rect 80550 5011 80566 5028
rect 80996 5028 81584 5044
rect 80996 5011 81012 5028
rect 80550 4994 80752 5011
rect 79792 4956 80752 4994
rect 80810 4994 81012 5011
rect 81568 5011 81584 5028
rect 82014 5028 82602 5044
rect 82014 5011 82030 5028
rect 81568 4994 81770 5011
rect 80810 4956 81770 4994
rect 81828 4994 82030 5011
rect 82586 5011 82602 5028
rect 83032 5028 83620 5044
rect 83032 5011 83048 5028
rect 82586 4994 82788 5011
rect 81828 4956 82788 4994
rect 82846 4994 83048 5011
rect 83604 5011 83620 5028
rect 84050 5028 84638 5044
rect 84050 5011 84066 5028
rect 83604 4994 83806 5011
rect 82846 4956 83806 4994
rect 83864 4994 84066 5011
rect 84622 5011 84638 5028
rect 85068 5028 85656 5044
rect 85068 5011 85084 5028
rect 84622 4994 84824 5011
rect 83864 4956 84824 4994
rect 84882 4994 85084 5011
rect 85640 5011 85656 5028
rect 86086 5028 86674 5044
rect 86086 5011 86102 5028
rect 85640 4994 85842 5011
rect 84882 4956 85842 4994
rect 85900 4994 86102 5011
rect 86658 5011 86674 5028
rect 87104 5028 87692 5044
rect 87104 5011 87120 5028
rect 86658 4994 86860 5011
rect 85900 4956 86860 4994
rect 86918 4994 87120 5011
rect 87676 5011 87692 5028
rect 87676 4994 87878 5011
rect 86918 4956 87878 4994
rect 55777 4831 56365 4847
rect 55777 4814 55793 4831
rect 55591 4797 55793 4814
rect 56349 4814 56365 4831
rect 56795 4831 57383 4847
rect 56795 4814 56811 4831
rect 56349 4797 56551 4814
rect 55591 4759 56551 4797
rect 56609 4797 56811 4814
rect 57367 4814 57383 4831
rect 57813 4831 58401 4847
rect 57813 4814 57829 4831
rect 57367 4797 57569 4814
rect 56609 4759 57569 4797
rect 57627 4797 57829 4814
rect 58385 4814 58401 4831
rect 58831 4831 59419 4847
rect 58831 4814 58847 4831
rect 58385 4797 58587 4814
rect 57627 4759 58587 4797
rect 58645 4797 58847 4814
rect 59403 4814 59419 4831
rect 59849 4831 60437 4847
rect 59849 4814 59865 4831
rect 59403 4797 59605 4814
rect 58645 4759 59605 4797
rect 59663 4797 59865 4814
rect 60421 4814 60437 4831
rect 60867 4831 61455 4847
rect 60867 4814 60883 4831
rect 60421 4797 60623 4814
rect 59663 4759 60623 4797
rect 60681 4797 60883 4814
rect 61439 4814 61455 4831
rect 62628 4832 62784 4848
rect 62628 4815 62644 4832
rect 61439 4797 61641 4814
rect 60681 4759 61641 4797
rect 62586 4798 62644 4815
rect 62768 4815 62784 4832
rect 62926 4832 63082 4848
rect 62926 4815 62942 4832
rect 62768 4798 62826 4815
rect 62586 4760 62826 4798
rect 62884 4798 62942 4815
rect 63066 4815 63082 4832
rect 63224 4832 63380 4848
rect 63224 4815 63240 4832
rect 63066 4798 63124 4815
rect 62884 4760 63124 4798
rect 63182 4798 63240 4815
rect 63364 4815 63380 4832
rect 63522 4832 63678 4848
rect 63522 4815 63538 4832
rect 63364 4798 63422 4815
rect 63182 4760 63422 4798
rect 63480 4798 63538 4815
rect 63662 4815 63678 4832
rect 63820 4832 63976 4848
rect 63820 4815 63836 4832
rect 63662 4798 63720 4815
rect 63480 4760 63720 4798
rect 63778 4798 63836 4815
rect 63960 4815 63976 4832
rect 64118 4832 64274 4848
rect 64118 4815 64134 4832
rect 63960 4798 64018 4815
rect 63778 4760 64018 4798
rect 64076 4798 64134 4815
rect 64258 4815 64274 4832
rect 64416 4832 64572 4848
rect 64416 4815 64432 4832
rect 64258 4798 64316 4815
rect 64076 4760 64316 4798
rect 64374 4798 64432 4815
rect 64556 4815 64572 4832
rect 64714 4832 64870 4848
rect 64714 4815 64730 4832
rect 64556 4798 64614 4815
rect 64374 4760 64614 4798
rect 64672 4798 64730 4815
rect 64854 4815 64870 4832
rect 65012 4832 65168 4848
rect 65012 4815 65028 4832
rect 64854 4798 64912 4815
rect 64672 4760 64912 4798
rect 64970 4798 65028 4815
rect 65152 4815 65168 4832
rect 65310 4832 65466 4848
rect 65310 4815 65326 4832
rect 65152 4798 65210 4815
rect 64970 4760 65210 4798
rect 65268 4798 65326 4815
rect 65450 4815 65466 4832
rect 65608 4832 65764 4848
rect 65608 4815 65624 4832
rect 65450 4798 65508 4815
rect 65268 4760 65508 4798
rect 65566 4798 65624 4815
rect 65748 4815 65764 4832
rect 65748 4798 65806 4815
rect 65566 4760 65806 4798
rect 67576 4318 68536 4356
rect 67576 4301 67778 4318
rect 67762 4284 67778 4301
rect 68334 4301 68536 4318
rect 68594 4318 69554 4356
rect 68594 4301 68796 4318
rect 68334 4284 68350 4301
rect 67762 4268 68350 4284
rect 68780 4284 68796 4301
rect 69352 4301 69554 4318
rect 69612 4318 70572 4356
rect 69612 4301 69814 4318
rect 69352 4284 69368 4301
rect 68780 4268 69368 4284
rect 69798 4284 69814 4301
rect 70370 4301 70572 4318
rect 70630 4318 71590 4356
rect 70630 4301 70832 4318
rect 70370 4284 70386 4301
rect 69798 4268 70386 4284
rect 70816 4284 70832 4301
rect 71388 4301 71590 4318
rect 71648 4318 72608 4356
rect 71648 4301 71850 4318
rect 71388 4284 71404 4301
rect 70816 4268 71404 4284
rect 71834 4284 71850 4301
rect 72406 4301 72608 4318
rect 72666 4318 73626 4356
rect 72666 4301 72868 4318
rect 72406 4284 72422 4301
rect 71834 4268 72422 4284
rect 72852 4284 72868 4301
rect 73424 4301 73626 4318
rect 73684 4318 74644 4356
rect 73684 4301 73886 4318
rect 73424 4284 73440 4301
rect 72852 4268 73440 4284
rect 73870 4284 73886 4301
rect 74442 4301 74644 4318
rect 74702 4318 75662 4356
rect 74702 4301 74904 4318
rect 74442 4284 74458 4301
rect 73870 4268 74458 4284
rect 74888 4284 74904 4301
rect 75460 4301 75662 4318
rect 75720 4318 76680 4356
rect 75720 4301 75922 4318
rect 75460 4284 75476 4301
rect 74888 4268 75476 4284
rect 75906 4284 75922 4301
rect 76478 4301 76680 4318
rect 76738 4318 77698 4356
rect 76738 4301 76940 4318
rect 76478 4284 76494 4301
rect 75906 4268 76494 4284
rect 76924 4284 76940 4301
rect 77496 4301 77698 4318
rect 77756 4318 78716 4356
rect 77756 4301 77958 4318
rect 77496 4284 77512 4301
rect 76924 4268 77512 4284
rect 77942 4284 77958 4301
rect 78514 4301 78716 4318
rect 78774 4318 79734 4356
rect 78774 4301 78976 4318
rect 78514 4284 78530 4301
rect 77942 4268 78530 4284
rect 78960 4284 78976 4301
rect 79532 4301 79734 4318
rect 79792 4318 80752 4356
rect 79792 4301 79994 4318
rect 79532 4284 79548 4301
rect 78960 4268 79548 4284
rect 79978 4284 79994 4301
rect 80550 4301 80752 4318
rect 80810 4318 81770 4356
rect 80810 4301 81012 4318
rect 80550 4284 80566 4301
rect 79978 4268 80566 4284
rect 80996 4284 81012 4301
rect 81568 4301 81770 4318
rect 81828 4318 82788 4356
rect 81828 4301 82030 4318
rect 81568 4284 81584 4301
rect 80996 4268 81584 4284
rect 82014 4284 82030 4301
rect 82586 4301 82788 4318
rect 82846 4318 83806 4356
rect 82846 4301 83048 4318
rect 82586 4284 82602 4301
rect 82014 4268 82602 4284
rect 83032 4284 83048 4301
rect 83604 4301 83806 4318
rect 83864 4318 84824 4356
rect 83864 4301 84066 4318
rect 83604 4284 83620 4301
rect 83032 4268 83620 4284
rect 84050 4284 84066 4301
rect 84622 4301 84824 4318
rect 84882 4318 85842 4356
rect 84882 4301 85084 4318
rect 84622 4284 84638 4301
rect 84050 4268 84638 4284
rect 85068 4284 85084 4301
rect 85640 4301 85842 4318
rect 85900 4318 86860 4356
rect 85900 4301 86102 4318
rect 85640 4284 85656 4301
rect 85068 4268 85656 4284
rect 86086 4284 86102 4301
rect 86658 4301 86860 4318
rect 86918 4318 87878 4356
rect 86918 4301 87120 4318
rect 86658 4284 86674 4301
rect 86086 4268 86674 4284
rect 87104 4284 87120 4301
rect 87676 4301 87878 4318
rect 87676 4284 87692 4301
rect 87104 4268 87692 4284
rect 55591 4121 56551 4159
rect 55591 4104 55793 4121
rect 55777 4087 55793 4104
rect 56349 4104 56551 4121
rect 56609 4121 57569 4159
rect 56609 4104 56811 4121
rect 56349 4087 56365 4104
rect 55777 4071 56365 4087
rect 56795 4087 56811 4104
rect 57367 4104 57569 4121
rect 57627 4121 58587 4159
rect 57627 4104 57829 4121
rect 57367 4087 57383 4104
rect 56795 4071 57383 4087
rect 57813 4087 57829 4104
rect 58385 4104 58587 4121
rect 58645 4121 59605 4159
rect 58645 4104 58847 4121
rect 58385 4087 58401 4104
rect 57813 4071 58401 4087
rect 58831 4087 58847 4104
rect 59403 4104 59605 4121
rect 59663 4121 60623 4159
rect 59663 4104 59865 4121
rect 59403 4087 59419 4104
rect 58831 4071 59419 4087
rect 59849 4087 59865 4104
rect 60421 4104 60623 4121
rect 60681 4121 61641 4159
rect 60681 4104 60883 4121
rect 60421 4087 60437 4104
rect 59849 4071 60437 4087
rect 60867 4087 60883 4104
rect 61439 4104 61641 4121
rect 62586 4122 62826 4160
rect 62586 4105 62644 4122
rect 61439 4087 61455 4104
rect 60867 4071 61455 4087
rect 62628 4088 62644 4105
rect 62768 4105 62826 4122
rect 62884 4122 63124 4160
rect 62884 4105 62942 4122
rect 62768 4088 62784 4105
rect 62628 4072 62784 4088
rect 62926 4088 62942 4105
rect 63066 4105 63124 4122
rect 63182 4122 63422 4160
rect 63182 4105 63240 4122
rect 63066 4088 63082 4105
rect 62926 4072 63082 4088
rect 63224 4088 63240 4105
rect 63364 4105 63422 4122
rect 63480 4122 63720 4160
rect 63480 4105 63538 4122
rect 63364 4088 63380 4105
rect 63224 4072 63380 4088
rect 63522 4088 63538 4105
rect 63662 4105 63720 4122
rect 63778 4122 64018 4160
rect 63778 4105 63836 4122
rect 63662 4088 63678 4105
rect 63522 4072 63678 4088
rect 63820 4088 63836 4105
rect 63960 4105 64018 4122
rect 64076 4122 64316 4160
rect 64076 4105 64134 4122
rect 63960 4088 63976 4105
rect 63820 4072 63976 4088
rect 64118 4088 64134 4105
rect 64258 4105 64316 4122
rect 64374 4122 64614 4160
rect 64374 4105 64432 4122
rect 64258 4088 64274 4105
rect 64118 4072 64274 4088
rect 64416 4088 64432 4105
rect 64556 4105 64614 4122
rect 64672 4122 64912 4160
rect 64672 4105 64730 4122
rect 64556 4088 64572 4105
rect 64416 4072 64572 4088
rect 64714 4088 64730 4105
rect 64854 4105 64912 4122
rect 64970 4122 65210 4160
rect 64970 4105 65028 4122
rect 64854 4088 64870 4105
rect 64714 4072 64870 4088
rect 65012 4088 65028 4105
rect 65152 4105 65210 4122
rect 65268 4122 65508 4160
rect 65268 4105 65326 4122
rect 65152 4088 65168 4105
rect 65012 4072 65168 4088
rect 65310 4088 65326 4105
rect 65450 4105 65508 4122
rect 65566 4122 65806 4160
rect 65566 4105 65624 4122
rect 65450 4088 65466 4105
rect 65310 4072 65466 4088
rect 65608 4088 65624 4105
rect 65748 4105 65806 4122
rect 65748 4088 65764 4105
rect 65608 4072 65764 4088
rect 67762 3794 68350 3810
rect 67762 3777 67778 3794
rect 67576 3760 67778 3777
rect 68334 3777 68350 3794
rect 68780 3794 69368 3810
rect 68780 3777 68796 3794
rect 68334 3760 68536 3777
rect 55776 3718 56364 3734
rect 55776 3701 55792 3718
rect 55590 3684 55792 3701
rect 56348 3701 56364 3718
rect 56794 3718 57382 3734
rect 56794 3701 56810 3718
rect 56348 3684 56550 3701
rect 55590 3646 56550 3684
rect 56608 3684 56810 3701
rect 57366 3701 57382 3718
rect 57812 3718 58400 3734
rect 57812 3701 57828 3718
rect 57366 3684 57568 3701
rect 56608 3646 57568 3684
rect 57626 3684 57828 3701
rect 58384 3701 58400 3718
rect 58830 3718 59418 3734
rect 58830 3701 58846 3718
rect 58384 3684 58586 3701
rect 57626 3646 58586 3684
rect 58644 3684 58846 3701
rect 59402 3701 59418 3718
rect 59848 3718 60436 3734
rect 59848 3701 59864 3718
rect 59402 3684 59604 3701
rect 58644 3646 59604 3684
rect 59662 3684 59864 3701
rect 60420 3701 60436 3718
rect 60866 3718 61454 3734
rect 60866 3701 60882 3718
rect 60420 3684 60622 3701
rect 59662 3646 60622 3684
rect 60680 3684 60882 3701
rect 61438 3701 61454 3718
rect 62628 3720 62784 3736
rect 62628 3703 62644 3720
rect 61438 3684 61640 3701
rect 60680 3646 61640 3684
rect 62586 3686 62644 3703
rect 62768 3703 62784 3720
rect 62926 3720 63082 3736
rect 62926 3703 62942 3720
rect 62768 3686 62826 3703
rect 62586 3648 62826 3686
rect 62884 3686 62942 3703
rect 63066 3703 63082 3720
rect 63224 3720 63380 3736
rect 63224 3703 63240 3720
rect 63066 3686 63124 3703
rect 62884 3648 63124 3686
rect 63182 3686 63240 3703
rect 63364 3703 63380 3720
rect 63522 3720 63678 3736
rect 63522 3703 63538 3720
rect 63364 3686 63422 3703
rect 63182 3648 63422 3686
rect 63480 3686 63538 3703
rect 63662 3703 63678 3720
rect 63820 3720 63976 3736
rect 63820 3703 63836 3720
rect 63662 3686 63720 3703
rect 63480 3648 63720 3686
rect 63778 3686 63836 3703
rect 63960 3703 63976 3720
rect 64118 3720 64274 3736
rect 64118 3703 64134 3720
rect 63960 3686 64018 3703
rect 63778 3648 64018 3686
rect 64076 3686 64134 3703
rect 64258 3703 64274 3720
rect 64416 3720 64572 3736
rect 64416 3703 64432 3720
rect 64258 3686 64316 3703
rect 64076 3648 64316 3686
rect 64374 3686 64432 3703
rect 64556 3703 64572 3720
rect 64714 3720 64870 3736
rect 64714 3703 64730 3720
rect 64556 3686 64614 3703
rect 64374 3648 64614 3686
rect 64672 3686 64730 3703
rect 64854 3703 64870 3720
rect 65012 3720 65168 3736
rect 65012 3703 65028 3720
rect 64854 3686 64912 3703
rect 64672 3648 64912 3686
rect 64970 3686 65028 3703
rect 65152 3703 65168 3720
rect 65310 3720 65466 3736
rect 65310 3703 65326 3720
rect 65152 3686 65210 3703
rect 64970 3648 65210 3686
rect 65268 3686 65326 3703
rect 65450 3703 65466 3720
rect 65608 3720 65764 3736
rect 67576 3722 68536 3760
rect 68594 3760 68796 3777
rect 69352 3777 69368 3794
rect 69798 3794 70386 3810
rect 69798 3777 69814 3794
rect 69352 3760 69554 3777
rect 68594 3722 69554 3760
rect 69612 3760 69814 3777
rect 70370 3777 70386 3794
rect 70816 3794 71404 3810
rect 70816 3777 70832 3794
rect 70370 3760 70572 3777
rect 69612 3722 70572 3760
rect 70630 3760 70832 3777
rect 71388 3777 71404 3794
rect 71834 3794 72422 3810
rect 71834 3777 71850 3794
rect 71388 3760 71590 3777
rect 70630 3722 71590 3760
rect 71648 3760 71850 3777
rect 72406 3777 72422 3794
rect 72852 3794 73440 3810
rect 72852 3777 72868 3794
rect 72406 3760 72608 3777
rect 71648 3722 72608 3760
rect 72666 3760 72868 3777
rect 73424 3777 73440 3794
rect 73870 3794 74458 3810
rect 73870 3777 73886 3794
rect 73424 3760 73626 3777
rect 72666 3722 73626 3760
rect 73684 3760 73886 3777
rect 74442 3777 74458 3794
rect 74888 3794 75476 3810
rect 74888 3777 74904 3794
rect 74442 3760 74644 3777
rect 73684 3722 74644 3760
rect 74702 3760 74904 3777
rect 75460 3777 75476 3794
rect 75906 3794 76494 3810
rect 75906 3777 75922 3794
rect 75460 3760 75662 3777
rect 74702 3722 75662 3760
rect 75720 3760 75922 3777
rect 76478 3777 76494 3794
rect 76924 3794 77512 3810
rect 76924 3777 76940 3794
rect 76478 3760 76680 3777
rect 75720 3722 76680 3760
rect 76738 3760 76940 3777
rect 77496 3777 77512 3794
rect 77942 3794 78530 3810
rect 77942 3777 77958 3794
rect 77496 3760 77698 3777
rect 76738 3722 77698 3760
rect 77756 3760 77958 3777
rect 78514 3777 78530 3794
rect 78960 3794 79548 3810
rect 78960 3777 78976 3794
rect 78514 3760 78716 3777
rect 77756 3722 78716 3760
rect 78774 3760 78976 3777
rect 79532 3777 79548 3794
rect 79978 3794 80566 3810
rect 79978 3777 79994 3794
rect 79532 3760 79734 3777
rect 78774 3722 79734 3760
rect 79792 3760 79994 3777
rect 80550 3777 80566 3794
rect 80996 3794 81584 3810
rect 80996 3777 81012 3794
rect 80550 3760 80752 3777
rect 79792 3722 80752 3760
rect 80810 3760 81012 3777
rect 81568 3777 81584 3794
rect 82014 3794 82602 3810
rect 82014 3777 82030 3794
rect 81568 3760 81770 3777
rect 80810 3722 81770 3760
rect 81828 3760 82030 3777
rect 82586 3777 82602 3794
rect 83032 3794 83620 3810
rect 83032 3777 83048 3794
rect 82586 3760 82788 3777
rect 81828 3722 82788 3760
rect 82846 3760 83048 3777
rect 83604 3777 83620 3794
rect 84050 3794 84638 3810
rect 84050 3777 84066 3794
rect 83604 3760 83806 3777
rect 82846 3722 83806 3760
rect 83864 3760 84066 3777
rect 84622 3777 84638 3794
rect 85068 3794 85656 3810
rect 85068 3777 85084 3794
rect 84622 3760 84824 3777
rect 83864 3722 84824 3760
rect 84882 3760 85084 3777
rect 85640 3777 85656 3794
rect 86086 3794 86674 3810
rect 86086 3777 86102 3794
rect 85640 3760 85842 3777
rect 84882 3722 85842 3760
rect 85900 3760 86102 3777
rect 86658 3777 86674 3794
rect 87104 3794 87692 3810
rect 87104 3777 87120 3794
rect 86658 3760 86860 3777
rect 85900 3722 86860 3760
rect 86918 3760 87120 3777
rect 87676 3777 87692 3794
rect 87676 3760 87878 3777
rect 86918 3722 87878 3760
rect 65608 3703 65624 3720
rect 65450 3686 65508 3703
rect 65268 3648 65508 3686
rect 65566 3686 65624 3703
rect 65748 3703 65764 3720
rect 65748 3686 65806 3703
rect 65566 3648 65806 3686
rect 67576 3084 68536 3122
rect 67576 3067 67778 3084
rect 67762 3050 67778 3067
rect 68334 3067 68536 3084
rect 68594 3084 69554 3122
rect 68594 3067 68796 3084
rect 68334 3050 68350 3067
rect 55590 3008 56550 3046
rect 55590 2991 55792 3008
rect 55776 2974 55792 2991
rect 56348 2991 56550 3008
rect 56608 3008 57568 3046
rect 56608 2991 56810 3008
rect 56348 2974 56364 2991
rect 55776 2958 56364 2974
rect 56794 2974 56810 2991
rect 57366 2991 57568 3008
rect 57626 3008 58586 3046
rect 57626 2991 57828 3008
rect 57366 2974 57382 2991
rect 56794 2958 57382 2974
rect 57812 2974 57828 2991
rect 58384 2991 58586 3008
rect 58644 3008 59604 3046
rect 58644 2991 58846 3008
rect 58384 2974 58400 2991
rect 57812 2958 58400 2974
rect 58830 2974 58846 2991
rect 59402 2991 59604 3008
rect 59662 3008 60622 3046
rect 59662 2991 59864 3008
rect 59402 2974 59418 2991
rect 58830 2958 59418 2974
rect 59848 2974 59864 2991
rect 60420 2991 60622 3008
rect 60680 3008 61640 3046
rect 60680 2991 60882 3008
rect 60420 2974 60436 2991
rect 59848 2958 60436 2974
rect 60866 2974 60882 2991
rect 61438 2991 61640 3008
rect 62586 3010 62826 3048
rect 62586 2993 62644 3010
rect 61438 2974 61454 2991
rect 60866 2958 61454 2974
rect 62628 2976 62644 2993
rect 62768 2993 62826 3010
rect 62884 3010 63124 3048
rect 62884 2993 62942 3010
rect 62768 2976 62784 2993
rect 62628 2960 62784 2976
rect 62926 2976 62942 2993
rect 63066 2993 63124 3010
rect 63182 3010 63422 3048
rect 63182 2993 63240 3010
rect 63066 2976 63082 2993
rect 62926 2960 63082 2976
rect 63224 2976 63240 2993
rect 63364 2993 63422 3010
rect 63480 3010 63720 3048
rect 63480 2993 63538 3010
rect 63364 2976 63380 2993
rect 63224 2960 63380 2976
rect 63522 2976 63538 2993
rect 63662 2993 63720 3010
rect 63778 3010 64018 3048
rect 63778 2993 63836 3010
rect 63662 2976 63678 2993
rect 63522 2960 63678 2976
rect 63820 2976 63836 2993
rect 63960 2993 64018 3010
rect 64076 3010 64316 3048
rect 64076 2993 64134 3010
rect 63960 2976 63976 2993
rect 63820 2960 63976 2976
rect 64118 2976 64134 2993
rect 64258 2993 64316 3010
rect 64374 3010 64614 3048
rect 64374 2993 64432 3010
rect 64258 2976 64274 2993
rect 64118 2960 64274 2976
rect 64416 2976 64432 2993
rect 64556 2993 64614 3010
rect 64672 3010 64912 3048
rect 64672 2993 64730 3010
rect 64556 2976 64572 2993
rect 64416 2960 64572 2976
rect 64714 2976 64730 2993
rect 64854 2993 64912 3010
rect 64970 3010 65210 3048
rect 64970 2993 65028 3010
rect 64854 2976 64870 2993
rect 64714 2960 64870 2976
rect 65012 2976 65028 2993
rect 65152 2993 65210 3010
rect 65268 3010 65508 3048
rect 65268 2993 65326 3010
rect 65152 2976 65168 2993
rect 65012 2960 65168 2976
rect 65310 2976 65326 2993
rect 65450 2993 65508 3010
rect 65566 3010 65806 3048
rect 67762 3034 68350 3050
rect 68780 3050 68796 3067
rect 69352 3067 69554 3084
rect 69612 3084 70572 3122
rect 69612 3067 69814 3084
rect 69352 3050 69368 3067
rect 68780 3034 69368 3050
rect 69798 3050 69814 3067
rect 70370 3067 70572 3084
rect 70630 3084 71590 3122
rect 70630 3067 70832 3084
rect 70370 3050 70386 3067
rect 69798 3034 70386 3050
rect 70816 3050 70832 3067
rect 71388 3067 71590 3084
rect 71648 3084 72608 3122
rect 71648 3067 71850 3084
rect 71388 3050 71404 3067
rect 70816 3034 71404 3050
rect 71834 3050 71850 3067
rect 72406 3067 72608 3084
rect 72666 3084 73626 3122
rect 72666 3067 72868 3084
rect 72406 3050 72422 3067
rect 71834 3034 72422 3050
rect 72852 3050 72868 3067
rect 73424 3067 73626 3084
rect 73684 3084 74644 3122
rect 73684 3067 73886 3084
rect 73424 3050 73440 3067
rect 72852 3034 73440 3050
rect 73870 3050 73886 3067
rect 74442 3067 74644 3084
rect 74702 3084 75662 3122
rect 74702 3067 74904 3084
rect 74442 3050 74458 3067
rect 73870 3034 74458 3050
rect 74888 3050 74904 3067
rect 75460 3067 75662 3084
rect 75720 3084 76680 3122
rect 75720 3067 75922 3084
rect 75460 3050 75476 3067
rect 74888 3034 75476 3050
rect 75906 3050 75922 3067
rect 76478 3067 76680 3084
rect 76738 3084 77698 3122
rect 76738 3067 76940 3084
rect 76478 3050 76494 3067
rect 75906 3034 76494 3050
rect 76924 3050 76940 3067
rect 77496 3067 77698 3084
rect 77756 3084 78716 3122
rect 77756 3067 77958 3084
rect 77496 3050 77512 3067
rect 76924 3034 77512 3050
rect 77942 3050 77958 3067
rect 78514 3067 78716 3084
rect 78774 3084 79734 3122
rect 78774 3067 78976 3084
rect 78514 3050 78530 3067
rect 77942 3034 78530 3050
rect 78960 3050 78976 3067
rect 79532 3067 79734 3084
rect 79792 3084 80752 3122
rect 79792 3067 79994 3084
rect 79532 3050 79548 3067
rect 78960 3034 79548 3050
rect 79978 3050 79994 3067
rect 80550 3067 80752 3084
rect 80810 3084 81770 3122
rect 80810 3067 81012 3084
rect 80550 3050 80566 3067
rect 79978 3034 80566 3050
rect 80996 3050 81012 3067
rect 81568 3067 81770 3084
rect 81828 3084 82788 3122
rect 81828 3067 82030 3084
rect 81568 3050 81584 3067
rect 80996 3034 81584 3050
rect 82014 3050 82030 3067
rect 82586 3067 82788 3084
rect 82846 3084 83806 3122
rect 82846 3067 83048 3084
rect 82586 3050 82602 3067
rect 82014 3034 82602 3050
rect 83032 3050 83048 3067
rect 83604 3067 83806 3084
rect 83864 3084 84824 3122
rect 83864 3067 84066 3084
rect 83604 3050 83620 3067
rect 83032 3034 83620 3050
rect 84050 3050 84066 3067
rect 84622 3067 84824 3084
rect 84882 3084 85842 3122
rect 84882 3067 85084 3084
rect 84622 3050 84638 3067
rect 84050 3034 84638 3050
rect 85068 3050 85084 3067
rect 85640 3067 85842 3084
rect 85900 3084 86860 3122
rect 85900 3067 86102 3084
rect 85640 3050 85656 3067
rect 85068 3034 85656 3050
rect 86086 3050 86102 3067
rect 86658 3067 86860 3084
rect 86918 3084 87878 3122
rect 86918 3067 87120 3084
rect 86658 3050 86674 3067
rect 86086 3034 86674 3050
rect 87104 3050 87120 3067
rect 87676 3067 87878 3084
rect 87676 3050 87692 3067
rect 87104 3034 87692 3050
rect 65566 2993 65624 3010
rect 65450 2976 65466 2993
rect 65310 2960 65466 2976
rect 65608 2976 65624 2993
rect 65748 2993 65806 3010
rect 65748 2976 65764 2993
rect 65608 2960 65764 2976
rect 55777 2607 56365 2623
rect 55777 2590 55793 2607
rect 55591 2573 55793 2590
rect 56349 2590 56365 2607
rect 56795 2607 57383 2623
rect 56795 2590 56811 2607
rect 56349 2573 56551 2590
rect 55591 2535 56551 2573
rect 56609 2573 56811 2590
rect 57367 2590 57383 2607
rect 57813 2607 58401 2623
rect 57813 2590 57829 2607
rect 57367 2573 57569 2590
rect 56609 2535 57569 2573
rect 57627 2573 57829 2590
rect 58385 2590 58401 2607
rect 58831 2607 59419 2623
rect 58831 2590 58847 2607
rect 58385 2573 58587 2590
rect 57627 2535 58587 2573
rect 58645 2573 58847 2590
rect 59403 2590 59419 2607
rect 59849 2607 60437 2623
rect 59849 2590 59865 2607
rect 59403 2573 59605 2590
rect 58645 2535 59605 2573
rect 59663 2573 59865 2590
rect 60421 2590 60437 2607
rect 60867 2607 61455 2623
rect 60867 2590 60883 2607
rect 60421 2573 60623 2590
rect 59663 2535 60623 2573
rect 60681 2573 60883 2590
rect 61439 2590 61455 2607
rect 62626 2608 62782 2624
rect 62626 2591 62642 2608
rect 61439 2573 61641 2590
rect 60681 2535 61641 2573
rect 62584 2574 62642 2591
rect 62766 2591 62782 2608
rect 62924 2608 63080 2624
rect 62924 2591 62940 2608
rect 62766 2574 62824 2591
rect 62584 2536 62824 2574
rect 62882 2574 62940 2591
rect 63064 2591 63080 2608
rect 63222 2608 63378 2624
rect 63222 2591 63238 2608
rect 63064 2574 63122 2591
rect 62882 2536 63122 2574
rect 63180 2574 63238 2591
rect 63362 2591 63378 2608
rect 63520 2608 63676 2624
rect 63520 2591 63536 2608
rect 63362 2574 63420 2591
rect 63180 2536 63420 2574
rect 63478 2574 63536 2591
rect 63660 2591 63676 2608
rect 63818 2608 63974 2624
rect 63818 2591 63834 2608
rect 63660 2574 63718 2591
rect 63478 2536 63718 2574
rect 63776 2574 63834 2591
rect 63958 2591 63974 2608
rect 64116 2608 64272 2624
rect 64116 2591 64132 2608
rect 63958 2574 64016 2591
rect 63776 2536 64016 2574
rect 64074 2574 64132 2591
rect 64256 2591 64272 2608
rect 64414 2608 64570 2624
rect 64414 2591 64430 2608
rect 64256 2574 64314 2591
rect 64074 2536 64314 2574
rect 64372 2574 64430 2591
rect 64554 2591 64570 2608
rect 64712 2608 64868 2624
rect 64712 2591 64728 2608
rect 64554 2574 64612 2591
rect 64372 2536 64612 2574
rect 64670 2574 64728 2591
rect 64852 2591 64868 2608
rect 65010 2608 65166 2624
rect 65010 2591 65026 2608
rect 64852 2574 64910 2591
rect 64670 2536 64910 2574
rect 64968 2574 65026 2591
rect 65150 2591 65166 2608
rect 65308 2608 65464 2624
rect 65308 2591 65324 2608
rect 65150 2574 65208 2591
rect 64968 2536 65208 2574
rect 65266 2574 65324 2591
rect 65448 2591 65464 2608
rect 65606 2608 65762 2624
rect 65606 2591 65622 2608
rect 65448 2574 65506 2591
rect 65266 2536 65506 2574
rect 65564 2574 65622 2591
rect 65746 2591 65762 2608
rect 65746 2574 65804 2591
rect 65564 2536 65804 2574
rect 67762 2560 68350 2576
rect 67762 2543 67778 2560
rect 67576 2526 67778 2543
rect 68334 2543 68350 2560
rect 68780 2560 69368 2576
rect 68780 2543 68796 2560
rect 68334 2526 68536 2543
rect 67576 2488 68536 2526
rect 68594 2526 68796 2543
rect 69352 2543 69368 2560
rect 69798 2560 70386 2576
rect 69798 2543 69814 2560
rect 69352 2526 69554 2543
rect 68594 2488 69554 2526
rect 69612 2526 69814 2543
rect 70370 2543 70386 2560
rect 70816 2560 71404 2576
rect 70816 2543 70832 2560
rect 70370 2526 70572 2543
rect 69612 2488 70572 2526
rect 70630 2526 70832 2543
rect 71388 2543 71404 2560
rect 71834 2560 72422 2576
rect 71834 2543 71850 2560
rect 71388 2526 71590 2543
rect 70630 2488 71590 2526
rect 71648 2526 71850 2543
rect 72406 2543 72422 2560
rect 72852 2560 73440 2576
rect 72852 2543 72868 2560
rect 72406 2526 72608 2543
rect 71648 2488 72608 2526
rect 72666 2526 72868 2543
rect 73424 2543 73440 2560
rect 73870 2560 74458 2576
rect 73870 2543 73886 2560
rect 73424 2526 73626 2543
rect 72666 2488 73626 2526
rect 73684 2526 73886 2543
rect 74442 2543 74458 2560
rect 74888 2560 75476 2576
rect 74888 2543 74904 2560
rect 74442 2526 74644 2543
rect 73684 2488 74644 2526
rect 74702 2526 74904 2543
rect 75460 2543 75476 2560
rect 75906 2560 76494 2576
rect 75906 2543 75922 2560
rect 75460 2526 75662 2543
rect 74702 2488 75662 2526
rect 75720 2526 75922 2543
rect 76478 2543 76494 2560
rect 76924 2560 77512 2576
rect 76924 2543 76940 2560
rect 76478 2526 76680 2543
rect 75720 2488 76680 2526
rect 76738 2526 76940 2543
rect 77496 2543 77512 2560
rect 77942 2560 78530 2576
rect 77942 2543 77958 2560
rect 77496 2526 77698 2543
rect 76738 2488 77698 2526
rect 77756 2526 77958 2543
rect 78514 2543 78530 2560
rect 78960 2560 79548 2576
rect 78960 2543 78976 2560
rect 78514 2526 78716 2543
rect 77756 2488 78716 2526
rect 78774 2526 78976 2543
rect 79532 2543 79548 2560
rect 79978 2560 80566 2576
rect 79978 2543 79994 2560
rect 79532 2526 79734 2543
rect 78774 2488 79734 2526
rect 79792 2526 79994 2543
rect 80550 2543 80566 2560
rect 80996 2560 81584 2576
rect 80996 2543 81012 2560
rect 80550 2526 80752 2543
rect 79792 2488 80752 2526
rect 80810 2526 81012 2543
rect 81568 2543 81584 2560
rect 82014 2560 82602 2576
rect 82014 2543 82030 2560
rect 81568 2526 81770 2543
rect 80810 2488 81770 2526
rect 81828 2526 82030 2543
rect 82586 2543 82602 2560
rect 83032 2560 83620 2576
rect 83032 2543 83048 2560
rect 82586 2526 82788 2543
rect 81828 2488 82788 2526
rect 82846 2526 83048 2543
rect 83604 2543 83620 2560
rect 84050 2560 84638 2576
rect 84050 2543 84066 2560
rect 83604 2526 83806 2543
rect 82846 2488 83806 2526
rect 83864 2526 84066 2543
rect 84622 2543 84638 2560
rect 85068 2560 85656 2576
rect 85068 2543 85084 2560
rect 84622 2526 84824 2543
rect 83864 2488 84824 2526
rect 84882 2526 85084 2543
rect 85640 2543 85656 2560
rect 86086 2560 86674 2576
rect 86086 2543 86102 2560
rect 85640 2526 85842 2543
rect 84882 2488 85842 2526
rect 85900 2526 86102 2543
rect 86658 2543 86674 2560
rect 87104 2560 87692 2576
rect 87104 2543 87120 2560
rect 86658 2526 86860 2543
rect 85900 2488 86860 2526
rect 86918 2526 87120 2543
rect 87676 2543 87692 2560
rect 87676 2526 87878 2543
rect 86918 2488 87878 2526
rect 55591 1897 56551 1935
rect 55591 1880 55793 1897
rect 55777 1863 55793 1880
rect 56349 1880 56551 1897
rect 56609 1897 57569 1935
rect 56609 1880 56811 1897
rect 56349 1863 56365 1880
rect 55777 1847 56365 1863
rect 56795 1863 56811 1880
rect 57367 1880 57569 1897
rect 57627 1897 58587 1935
rect 57627 1880 57829 1897
rect 57367 1863 57383 1880
rect 56795 1847 57383 1863
rect 57813 1863 57829 1880
rect 58385 1880 58587 1897
rect 58645 1897 59605 1935
rect 58645 1880 58847 1897
rect 58385 1863 58401 1880
rect 57813 1847 58401 1863
rect 58831 1863 58847 1880
rect 59403 1880 59605 1897
rect 59663 1897 60623 1935
rect 59663 1880 59865 1897
rect 59403 1863 59419 1880
rect 58831 1847 59419 1863
rect 59849 1863 59865 1880
rect 60421 1880 60623 1897
rect 60681 1897 61641 1935
rect 60681 1880 60883 1897
rect 60421 1863 60437 1880
rect 59849 1847 60437 1863
rect 60867 1863 60883 1880
rect 61439 1880 61641 1897
rect 62584 1898 62824 1936
rect 62584 1881 62642 1898
rect 61439 1863 61455 1880
rect 60867 1847 61455 1863
rect 62626 1864 62642 1881
rect 62766 1881 62824 1898
rect 62882 1898 63122 1936
rect 62882 1881 62940 1898
rect 62766 1864 62782 1881
rect 62626 1848 62782 1864
rect 62924 1864 62940 1881
rect 63064 1881 63122 1898
rect 63180 1898 63420 1936
rect 63180 1881 63238 1898
rect 63064 1864 63080 1881
rect 62924 1848 63080 1864
rect 63222 1864 63238 1881
rect 63362 1881 63420 1898
rect 63478 1898 63718 1936
rect 63478 1881 63536 1898
rect 63362 1864 63378 1881
rect 63222 1848 63378 1864
rect 63520 1864 63536 1881
rect 63660 1881 63718 1898
rect 63776 1898 64016 1936
rect 63776 1881 63834 1898
rect 63660 1864 63676 1881
rect 63520 1848 63676 1864
rect 63818 1864 63834 1881
rect 63958 1881 64016 1898
rect 64074 1898 64314 1936
rect 64074 1881 64132 1898
rect 63958 1864 63974 1881
rect 63818 1848 63974 1864
rect 64116 1864 64132 1881
rect 64256 1881 64314 1898
rect 64372 1898 64612 1936
rect 64372 1881 64430 1898
rect 64256 1864 64272 1881
rect 64116 1848 64272 1864
rect 64414 1864 64430 1881
rect 64554 1881 64612 1898
rect 64670 1898 64910 1936
rect 64670 1881 64728 1898
rect 64554 1864 64570 1881
rect 64414 1848 64570 1864
rect 64712 1864 64728 1881
rect 64852 1881 64910 1898
rect 64968 1898 65208 1936
rect 64968 1881 65026 1898
rect 64852 1864 64868 1881
rect 64712 1848 64868 1864
rect 65010 1864 65026 1881
rect 65150 1881 65208 1898
rect 65266 1898 65506 1936
rect 65266 1881 65324 1898
rect 65150 1864 65166 1881
rect 65010 1848 65166 1864
rect 65308 1864 65324 1881
rect 65448 1881 65506 1898
rect 65564 1898 65804 1936
rect 65564 1881 65622 1898
rect 65448 1864 65464 1881
rect 65308 1848 65464 1864
rect 65606 1864 65622 1881
rect 65746 1881 65804 1898
rect 65746 1864 65762 1881
rect 65606 1848 65762 1864
rect 67576 1850 68536 1888
rect 67576 1833 67778 1850
rect 67762 1816 67778 1833
rect 68334 1833 68536 1850
rect 68594 1850 69554 1888
rect 68594 1833 68796 1850
rect 68334 1816 68350 1833
rect 67762 1800 68350 1816
rect 68780 1816 68796 1833
rect 69352 1833 69554 1850
rect 69612 1850 70572 1888
rect 69612 1833 69814 1850
rect 69352 1816 69368 1833
rect 68780 1800 69368 1816
rect 69798 1816 69814 1833
rect 70370 1833 70572 1850
rect 70630 1850 71590 1888
rect 70630 1833 70832 1850
rect 70370 1816 70386 1833
rect 69798 1800 70386 1816
rect 70816 1816 70832 1833
rect 71388 1833 71590 1850
rect 71648 1850 72608 1888
rect 71648 1833 71850 1850
rect 71388 1816 71404 1833
rect 70816 1800 71404 1816
rect 71834 1816 71850 1833
rect 72406 1833 72608 1850
rect 72666 1850 73626 1888
rect 72666 1833 72868 1850
rect 72406 1816 72422 1833
rect 71834 1800 72422 1816
rect 72852 1816 72868 1833
rect 73424 1833 73626 1850
rect 73684 1850 74644 1888
rect 73684 1833 73886 1850
rect 73424 1816 73440 1833
rect 72852 1800 73440 1816
rect 73870 1816 73886 1833
rect 74442 1833 74644 1850
rect 74702 1850 75662 1888
rect 74702 1833 74904 1850
rect 74442 1816 74458 1833
rect 73870 1800 74458 1816
rect 74888 1816 74904 1833
rect 75460 1833 75662 1850
rect 75720 1850 76680 1888
rect 75720 1833 75922 1850
rect 75460 1816 75476 1833
rect 74888 1800 75476 1816
rect 75906 1816 75922 1833
rect 76478 1833 76680 1850
rect 76738 1850 77698 1888
rect 76738 1833 76940 1850
rect 76478 1816 76494 1833
rect 75906 1800 76494 1816
rect 76924 1816 76940 1833
rect 77496 1833 77698 1850
rect 77756 1850 78716 1888
rect 77756 1833 77958 1850
rect 77496 1816 77512 1833
rect 76924 1800 77512 1816
rect 77942 1816 77958 1833
rect 78514 1833 78716 1850
rect 78774 1850 79734 1888
rect 78774 1833 78976 1850
rect 78514 1816 78530 1833
rect 77942 1800 78530 1816
rect 78960 1816 78976 1833
rect 79532 1833 79734 1850
rect 79792 1850 80752 1888
rect 79792 1833 79994 1850
rect 79532 1816 79548 1833
rect 78960 1800 79548 1816
rect 79978 1816 79994 1833
rect 80550 1833 80752 1850
rect 80810 1850 81770 1888
rect 80810 1833 81012 1850
rect 80550 1816 80566 1833
rect 79978 1800 80566 1816
rect 80996 1816 81012 1833
rect 81568 1833 81770 1850
rect 81828 1850 82788 1888
rect 81828 1833 82030 1850
rect 81568 1816 81584 1833
rect 80996 1800 81584 1816
rect 82014 1816 82030 1833
rect 82586 1833 82788 1850
rect 82846 1850 83806 1888
rect 82846 1833 83048 1850
rect 82586 1816 82602 1833
rect 82014 1800 82602 1816
rect 83032 1816 83048 1833
rect 83604 1833 83806 1850
rect 83864 1850 84824 1888
rect 83864 1833 84066 1850
rect 83604 1816 83620 1833
rect 83032 1800 83620 1816
rect 84050 1816 84066 1833
rect 84622 1833 84824 1850
rect 84882 1850 85842 1888
rect 84882 1833 85084 1850
rect 84622 1816 84638 1833
rect 84050 1800 84638 1816
rect 85068 1816 85084 1833
rect 85640 1833 85842 1850
rect 85900 1850 86860 1888
rect 85900 1833 86102 1850
rect 85640 1816 85656 1833
rect 85068 1800 85656 1816
rect 86086 1816 86102 1833
rect 86658 1833 86860 1850
rect 86918 1850 87878 1888
rect 86918 1833 87120 1850
rect 86658 1816 86674 1833
rect 86086 1800 86674 1816
rect 87104 1816 87120 1833
rect 87676 1833 87878 1850
rect 87676 1816 87692 1833
rect 87104 1800 87692 1816
rect 55776 1494 56364 1510
rect 55776 1477 55792 1494
rect 55590 1460 55792 1477
rect 56348 1477 56364 1494
rect 56794 1494 57382 1510
rect 56794 1477 56810 1494
rect 56348 1460 56550 1477
rect 55590 1422 56550 1460
rect 56608 1460 56810 1477
rect 57366 1477 57382 1494
rect 57812 1494 58400 1510
rect 57812 1477 57828 1494
rect 57366 1460 57568 1477
rect 56608 1422 57568 1460
rect 57626 1460 57828 1477
rect 58384 1477 58400 1494
rect 58830 1494 59418 1510
rect 58830 1477 58846 1494
rect 58384 1460 58586 1477
rect 57626 1422 58586 1460
rect 58644 1460 58846 1477
rect 59402 1477 59418 1494
rect 59848 1494 60436 1510
rect 59848 1477 59864 1494
rect 59402 1460 59604 1477
rect 58644 1422 59604 1460
rect 59662 1460 59864 1477
rect 60420 1477 60436 1494
rect 60866 1494 61454 1510
rect 60866 1477 60882 1494
rect 60420 1460 60622 1477
rect 59662 1422 60622 1460
rect 60680 1460 60882 1477
rect 61438 1477 61454 1494
rect 62626 1498 62782 1514
rect 62626 1481 62642 1498
rect 61438 1460 61640 1477
rect 60680 1422 61640 1460
rect 62584 1464 62642 1481
rect 62766 1481 62782 1498
rect 62924 1498 63080 1514
rect 62924 1481 62940 1498
rect 62766 1464 62824 1481
rect 62584 1426 62824 1464
rect 62882 1464 62940 1481
rect 63064 1481 63080 1498
rect 63222 1498 63378 1514
rect 63222 1481 63238 1498
rect 63064 1464 63122 1481
rect 62882 1426 63122 1464
rect 63180 1464 63238 1481
rect 63362 1481 63378 1498
rect 63520 1498 63676 1514
rect 63520 1481 63536 1498
rect 63362 1464 63420 1481
rect 63180 1426 63420 1464
rect 63478 1464 63536 1481
rect 63660 1481 63676 1498
rect 63818 1498 63974 1514
rect 63818 1481 63834 1498
rect 63660 1464 63718 1481
rect 63478 1426 63718 1464
rect 63776 1464 63834 1481
rect 63958 1481 63974 1498
rect 64116 1498 64272 1514
rect 64116 1481 64132 1498
rect 63958 1464 64016 1481
rect 63776 1426 64016 1464
rect 64074 1464 64132 1481
rect 64256 1481 64272 1498
rect 64414 1498 64570 1514
rect 64414 1481 64430 1498
rect 64256 1464 64314 1481
rect 64074 1426 64314 1464
rect 64372 1464 64430 1481
rect 64554 1481 64570 1498
rect 64712 1498 64868 1514
rect 64712 1481 64728 1498
rect 64554 1464 64612 1481
rect 64372 1426 64612 1464
rect 64670 1464 64728 1481
rect 64852 1481 64868 1498
rect 65010 1498 65166 1514
rect 65010 1481 65026 1498
rect 64852 1464 64910 1481
rect 64670 1426 64910 1464
rect 64968 1464 65026 1481
rect 65150 1481 65166 1498
rect 65308 1498 65464 1514
rect 65308 1481 65324 1498
rect 65150 1464 65208 1481
rect 64968 1426 65208 1464
rect 65266 1464 65324 1481
rect 65448 1481 65464 1498
rect 65606 1498 65762 1514
rect 65606 1481 65622 1498
rect 65448 1464 65506 1481
rect 65266 1426 65506 1464
rect 65564 1464 65622 1481
rect 65746 1481 65762 1498
rect 65746 1464 65804 1481
rect 65564 1426 65804 1464
rect 67762 1328 68350 1344
rect 67762 1311 67778 1328
rect 67576 1294 67778 1311
rect 68334 1311 68350 1328
rect 68780 1328 69368 1344
rect 68780 1311 68796 1328
rect 68334 1294 68536 1311
rect 67576 1256 68536 1294
rect 68594 1294 68796 1311
rect 69352 1311 69368 1328
rect 69798 1328 70386 1344
rect 69798 1311 69814 1328
rect 69352 1294 69554 1311
rect 68594 1256 69554 1294
rect 69612 1294 69814 1311
rect 70370 1311 70386 1328
rect 70816 1328 71404 1344
rect 70816 1311 70832 1328
rect 70370 1294 70572 1311
rect 69612 1256 70572 1294
rect 70630 1294 70832 1311
rect 71388 1311 71404 1328
rect 71834 1328 72422 1344
rect 71834 1311 71850 1328
rect 71388 1294 71590 1311
rect 70630 1256 71590 1294
rect 71648 1294 71850 1311
rect 72406 1311 72422 1328
rect 72852 1328 73440 1344
rect 72852 1311 72868 1328
rect 72406 1294 72608 1311
rect 71648 1256 72608 1294
rect 72666 1294 72868 1311
rect 73424 1311 73440 1328
rect 73870 1328 74458 1344
rect 73870 1311 73886 1328
rect 73424 1294 73626 1311
rect 72666 1256 73626 1294
rect 73684 1294 73886 1311
rect 74442 1311 74458 1328
rect 74888 1328 75476 1344
rect 74888 1311 74904 1328
rect 74442 1294 74644 1311
rect 73684 1256 74644 1294
rect 74702 1294 74904 1311
rect 75460 1311 75476 1328
rect 75906 1328 76494 1344
rect 75906 1311 75922 1328
rect 75460 1294 75662 1311
rect 74702 1256 75662 1294
rect 75720 1294 75922 1311
rect 76478 1311 76494 1328
rect 76924 1328 77512 1344
rect 76924 1311 76940 1328
rect 76478 1294 76680 1311
rect 75720 1256 76680 1294
rect 76738 1294 76940 1311
rect 77496 1311 77512 1328
rect 77942 1328 78530 1344
rect 77942 1311 77958 1328
rect 77496 1294 77698 1311
rect 76738 1256 77698 1294
rect 77756 1294 77958 1311
rect 78514 1311 78530 1328
rect 78960 1328 79548 1344
rect 78960 1311 78976 1328
rect 78514 1294 78716 1311
rect 77756 1256 78716 1294
rect 78774 1294 78976 1311
rect 79532 1311 79548 1328
rect 79978 1328 80566 1344
rect 79978 1311 79994 1328
rect 79532 1294 79734 1311
rect 78774 1256 79734 1294
rect 79792 1294 79994 1311
rect 80550 1311 80566 1328
rect 80996 1328 81584 1344
rect 80996 1311 81012 1328
rect 80550 1294 80752 1311
rect 79792 1256 80752 1294
rect 80810 1294 81012 1311
rect 81568 1311 81584 1328
rect 82014 1328 82602 1344
rect 82014 1311 82030 1328
rect 81568 1294 81770 1311
rect 80810 1256 81770 1294
rect 81828 1294 82030 1311
rect 82586 1311 82602 1328
rect 83032 1328 83620 1344
rect 83032 1311 83048 1328
rect 82586 1294 82788 1311
rect 81828 1256 82788 1294
rect 82846 1294 83048 1311
rect 83604 1311 83620 1328
rect 84050 1328 84638 1344
rect 84050 1311 84066 1328
rect 83604 1294 83806 1311
rect 82846 1256 83806 1294
rect 83864 1294 84066 1311
rect 84622 1311 84638 1328
rect 85068 1328 85656 1344
rect 85068 1311 85084 1328
rect 84622 1294 84824 1311
rect 83864 1256 84824 1294
rect 84882 1294 85084 1311
rect 85640 1311 85656 1328
rect 86086 1328 86674 1344
rect 86086 1311 86102 1328
rect 85640 1294 85842 1311
rect 84882 1256 85842 1294
rect 85900 1294 86102 1311
rect 86658 1311 86674 1328
rect 87104 1328 87692 1344
rect 87104 1311 87120 1328
rect 86658 1294 86860 1311
rect 85900 1256 86860 1294
rect 86918 1294 87120 1311
rect 87676 1311 87692 1328
rect 87676 1294 87878 1311
rect 86918 1256 87878 1294
rect 55590 784 56550 822
rect 55590 767 55792 784
rect 55776 750 55792 767
rect 56348 767 56550 784
rect 56608 784 57568 822
rect 56608 767 56810 784
rect 56348 750 56364 767
rect 55776 734 56364 750
rect 56794 750 56810 767
rect 57366 767 57568 784
rect 57626 784 58586 822
rect 57626 767 57828 784
rect 57366 750 57382 767
rect 56794 734 57382 750
rect 57812 750 57828 767
rect 58384 767 58586 784
rect 58644 784 59604 822
rect 58644 767 58846 784
rect 58384 750 58400 767
rect 57812 734 58400 750
rect 58830 750 58846 767
rect 59402 767 59604 784
rect 59662 784 60622 822
rect 59662 767 59864 784
rect 59402 750 59418 767
rect 58830 734 59418 750
rect 59848 750 59864 767
rect 60420 767 60622 784
rect 60680 784 61640 822
rect 60680 767 60882 784
rect 60420 750 60436 767
rect 59848 734 60436 750
rect 60866 750 60882 767
rect 61438 767 61640 784
rect 62584 788 62824 826
rect 62584 771 62642 788
rect 61438 750 61454 767
rect 60866 734 61454 750
rect 62626 754 62642 771
rect 62766 771 62824 788
rect 62882 788 63122 826
rect 62882 771 62940 788
rect 62766 754 62782 771
rect 62626 738 62782 754
rect 62924 754 62940 771
rect 63064 771 63122 788
rect 63180 788 63420 826
rect 63180 771 63238 788
rect 63064 754 63080 771
rect 62924 738 63080 754
rect 63222 754 63238 771
rect 63362 771 63420 788
rect 63478 788 63718 826
rect 63478 771 63536 788
rect 63362 754 63378 771
rect 63222 738 63378 754
rect 63520 754 63536 771
rect 63660 771 63718 788
rect 63776 788 64016 826
rect 63776 771 63834 788
rect 63660 754 63676 771
rect 63520 738 63676 754
rect 63818 754 63834 771
rect 63958 771 64016 788
rect 64074 788 64314 826
rect 64074 771 64132 788
rect 63958 754 63974 771
rect 63818 738 63974 754
rect 64116 754 64132 771
rect 64256 771 64314 788
rect 64372 788 64612 826
rect 64372 771 64430 788
rect 64256 754 64272 771
rect 64116 738 64272 754
rect 64414 754 64430 771
rect 64554 771 64612 788
rect 64670 788 64910 826
rect 64670 771 64728 788
rect 64554 754 64570 771
rect 64414 738 64570 754
rect 64712 754 64728 771
rect 64852 771 64910 788
rect 64968 788 65208 826
rect 64968 771 65026 788
rect 64852 754 64868 771
rect 64712 738 64868 754
rect 65010 754 65026 771
rect 65150 771 65208 788
rect 65266 788 65506 826
rect 65266 771 65324 788
rect 65150 754 65166 771
rect 65010 738 65166 754
rect 65308 754 65324 771
rect 65448 771 65506 788
rect 65564 788 65804 826
rect 65564 771 65622 788
rect 65448 754 65464 771
rect 65308 738 65464 754
rect 65606 754 65622 771
rect 65746 771 65804 788
rect 65746 754 65762 771
rect 65606 738 65762 754
rect 67576 618 68536 656
rect 67576 601 67778 618
rect 67762 584 67778 601
rect 68334 601 68536 618
rect 68594 618 69554 656
rect 68594 601 68796 618
rect 68334 584 68350 601
rect 67762 568 68350 584
rect 68780 584 68796 601
rect 69352 601 69554 618
rect 69612 618 70572 656
rect 69612 601 69814 618
rect 69352 584 69368 601
rect 68780 568 69368 584
rect 69798 584 69814 601
rect 70370 601 70572 618
rect 70630 618 71590 656
rect 70630 601 70832 618
rect 70370 584 70386 601
rect 69798 568 70386 584
rect 70816 584 70832 601
rect 71388 601 71590 618
rect 71648 618 72608 656
rect 71648 601 71850 618
rect 71388 584 71404 601
rect 70816 568 71404 584
rect 71834 584 71850 601
rect 72406 601 72608 618
rect 72666 618 73626 656
rect 72666 601 72868 618
rect 72406 584 72422 601
rect 71834 568 72422 584
rect 72852 584 72868 601
rect 73424 601 73626 618
rect 73684 618 74644 656
rect 73684 601 73886 618
rect 73424 584 73440 601
rect 72852 568 73440 584
rect 73870 584 73886 601
rect 74442 601 74644 618
rect 74702 618 75662 656
rect 74702 601 74904 618
rect 74442 584 74458 601
rect 73870 568 74458 584
rect 74888 584 74904 601
rect 75460 601 75662 618
rect 75720 618 76680 656
rect 75720 601 75922 618
rect 75460 584 75476 601
rect 74888 568 75476 584
rect 75906 584 75922 601
rect 76478 601 76680 618
rect 76738 618 77698 656
rect 76738 601 76940 618
rect 76478 584 76494 601
rect 75906 568 76494 584
rect 76924 584 76940 601
rect 77496 601 77698 618
rect 77756 618 78716 656
rect 77756 601 77958 618
rect 77496 584 77512 601
rect 76924 568 77512 584
rect 77942 584 77958 601
rect 78514 601 78716 618
rect 78774 618 79734 656
rect 78774 601 78976 618
rect 78514 584 78530 601
rect 77942 568 78530 584
rect 78960 584 78976 601
rect 79532 601 79734 618
rect 79792 618 80752 656
rect 79792 601 79994 618
rect 79532 584 79548 601
rect 78960 568 79548 584
rect 79978 584 79994 601
rect 80550 601 80752 618
rect 80810 618 81770 656
rect 80810 601 81012 618
rect 80550 584 80566 601
rect 79978 568 80566 584
rect 80996 584 81012 601
rect 81568 601 81770 618
rect 81828 618 82788 656
rect 81828 601 82030 618
rect 81568 584 81584 601
rect 80996 568 81584 584
rect 82014 584 82030 601
rect 82586 601 82788 618
rect 82846 618 83806 656
rect 82846 601 83048 618
rect 82586 584 82602 601
rect 82014 568 82602 584
rect 83032 584 83048 601
rect 83604 601 83806 618
rect 83864 618 84824 656
rect 83864 601 84066 618
rect 83604 584 83620 601
rect 83032 568 83620 584
rect 84050 584 84066 601
rect 84622 601 84824 618
rect 84882 618 85842 656
rect 84882 601 85084 618
rect 84622 584 84638 601
rect 84050 568 84638 584
rect 85068 584 85084 601
rect 85640 601 85842 618
rect 85900 618 86860 656
rect 85900 601 86102 618
rect 85640 584 85656 601
rect 85068 568 85656 584
rect 86086 584 86102 601
rect 86658 601 86860 618
rect 86918 618 87878 656
rect 86918 601 87120 618
rect 86658 584 86674 601
rect 86086 568 86674 584
rect 87104 584 87120 601
rect 87676 601 87878 618
rect 87676 584 87692 601
rect 87104 568 87692 584
<< polycont >>
rect 17686 27027 18242 27061
rect 18704 27027 19260 27061
rect 19722 27027 20278 27061
rect 20740 27027 21296 27061
rect 21758 27027 22314 27061
rect 22776 27027 23332 27061
rect 23794 27027 24350 27061
rect 24812 27027 25368 27061
rect 25830 27027 26386 27061
rect 26848 27027 27404 27061
rect 27866 27027 28422 27061
rect 28884 27027 29440 27061
rect 29902 27027 30458 27061
rect 30920 27027 31476 27061
rect 31938 27027 32494 27061
rect 32956 27027 33512 27061
rect 17686 26299 18242 26333
rect 18704 26299 19260 26333
rect 19722 26299 20278 26333
rect 20740 26299 21296 26333
rect 21758 26299 22314 26333
rect 22776 26299 23332 26333
rect 23794 26299 24350 26333
rect 24812 26299 25368 26333
rect 25830 26299 26386 26333
rect 26848 26299 27404 26333
rect 27866 26299 28422 26333
rect 28884 26299 29440 26333
rect 29902 26299 30458 26333
rect 30920 26299 31476 26333
rect 31938 26299 32494 26333
rect 32956 26299 33512 26333
rect 17686 25891 18242 25925
rect 18704 25891 19260 25925
rect 19722 25891 20278 25925
rect 20740 25891 21296 25925
rect 21758 25891 22314 25925
rect 22776 25891 23332 25925
rect 23794 25891 24350 25925
rect 24812 25891 25368 25925
rect 25830 25891 26386 25925
rect 26848 25891 27404 25925
rect 27866 25891 28422 25925
rect 28884 25891 29440 25925
rect 29902 25891 30458 25925
rect 30920 25891 31476 25925
rect 31938 25891 32494 25925
rect 32956 25891 33512 25925
rect 17686 25163 18242 25197
rect 18704 25163 19260 25197
rect 19722 25163 20278 25197
rect 20740 25163 21296 25197
rect 21758 25163 22314 25197
rect 22776 25163 23332 25197
rect 23794 25163 24350 25197
rect 24812 25163 25368 25197
rect 25830 25163 26386 25197
rect 26848 25163 27404 25197
rect 27866 25163 28422 25197
rect 28884 25163 29440 25197
rect 29902 25163 30458 25197
rect 30920 25163 31476 25197
rect 31938 25163 32494 25197
rect 32956 25163 33512 25197
rect 17686 24755 18242 24789
rect 18704 24755 19260 24789
rect 19722 24755 20278 24789
rect 20740 24755 21296 24789
rect 21758 24755 22314 24789
rect 22776 24755 23332 24789
rect 23794 24755 24350 24789
rect 24812 24755 25368 24789
rect 25830 24755 26386 24789
rect 26848 24755 27404 24789
rect 27866 24755 28422 24789
rect 28884 24755 29440 24789
rect 29902 24755 30458 24789
rect 30920 24755 31476 24789
rect 31938 24755 32494 24789
rect 32956 24755 33512 24789
rect 17686 24027 18242 24061
rect 18704 24027 19260 24061
rect 19722 24027 20278 24061
rect 20740 24027 21296 24061
rect 21758 24027 22314 24061
rect 22776 24027 23332 24061
rect 23794 24027 24350 24061
rect 24812 24027 25368 24061
rect 25830 24027 26386 24061
rect 26848 24027 27404 24061
rect 27866 24027 28422 24061
rect 28884 24027 29440 24061
rect 29902 24027 30458 24061
rect 30920 24027 31476 24061
rect 31938 24027 32494 24061
rect 32956 24027 33512 24061
rect 18672 22981 19228 23015
rect 19690 22981 20246 23015
rect 20708 22981 21264 23015
rect 21726 22981 22282 23015
rect 22744 22981 23300 23015
rect 23762 22981 24318 23015
rect 24780 22981 25336 23015
rect 25798 22981 26354 23015
rect 26816 22981 27372 23015
rect 27834 22981 28390 23015
rect 28852 22981 29408 23015
rect 29870 22981 30426 23015
rect 30888 22981 31444 23015
rect 31906 22981 32462 23015
rect 32924 22981 33480 23015
rect 18672 22253 19228 22287
rect 19690 22253 20246 22287
rect 20708 22253 21264 22287
rect 21726 22253 22282 22287
rect 22744 22253 23300 22287
rect 23762 22253 24318 22287
rect 24780 22253 25336 22287
rect 25798 22253 26354 22287
rect 26816 22253 27372 22287
rect 27834 22253 28390 22287
rect 28852 22253 29408 22287
rect 29870 22253 30426 22287
rect 30888 22253 31444 22287
rect 31906 22253 32462 22287
rect 32924 22253 33480 22287
rect 14664 21897 14740 21931
rect 14882 21897 14958 21931
rect 15100 21897 15176 21931
rect 15318 21897 15394 21931
rect 15536 21897 15612 21931
rect 15754 21897 15830 21931
rect 15972 21897 16048 21931
rect 16190 21897 16266 21931
rect 16408 21897 16484 21931
rect 16626 21897 16702 21931
rect 18672 21725 19228 21759
rect 19690 21725 20246 21759
rect 20708 21725 21264 21759
rect 21726 21725 22282 21759
rect 22744 21725 23300 21759
rect 23762 21725 24318 21759
rect 24780 21725 25336 21759
rect 25798 21725 26354 21759
rect 26816 21725 27372 21759
rect 27834 21725 28390 21759
rect 28852 21725 29408 21759
rect 29870 21725 30426 21759
rect 30888 21725 31444 21759
rect 31906 21725 32462 21759
rect 32924 21725 33480 21759
rect 14664 21369 14740 21403
rect 14882 21369 14958 21403
rect 15100 21369 15176 21403
rect 15318 21369 15394 21403
rect 15536 21369 15612 21403
rect 15754 21369 15830 21403
rect 15972 21369 16048 21403
rect 16190 21369 16266 21403
rect 16408 21369 16484 21403
rect 16626 21369 16702 21403
rect 14664 20959 14740 20993
rect 14882 20959 14958 20993
rect 15100 20959 15176 20993
rect 15318 20959 15394 20993
rect 15536 20959 15612 20993
rect 15754 20959 15830 20993
rect 15972 20959 16048 20993
rect 16190 20959 16266 20993
rect 16408 20959 16484 20993
rect 16626 20959 16702 20993
rect 18672 20997 19228 21031
rect 19690 20997 20246 21031
rect 20708 20997 21264 21031
rect 21726 20997 22282 21031
rect 22744 20997 23300 21031
rect 23762 20997 24318 21031
rect 24780 20997 25336 21031
rect 25798 20997 26354 21031
rect 26816 20997 27372 21031
rect 27834 20997 28390 21031
rect 28852 20997 29408 21031
rect 29870 20997 30426 21031
rect 30888 20997 31444 21031
rect 31906 20997 32462 21031
rect 32924 20997 33480 21031
rect 14664 20431 14740 20465
rect 14882 20431 14958 20465
rect 15100 20431 15176 20465
rect 15318 20431 15394 20465
rect 15536 20431 15612 20465
rect 15754 20431 15830 20465
rect 15972 20431 16048 20465
rect 16190 20431 16266 20465
rect 16408 20431 16484 20465
rect 16626 20431 16702 20465
rect 18672 20469 19228 20503
rect 19690 20469 20246 20503
rect 20708 20469 21264 20503
rect 21726 20469 22282 20503
rect 22744 20469 23300 20503
rect 23762 20469 24318 20503
rect 24780 20469 25336 20503
rect 25798 20469 26354 20503
rect 26816 20469 27372 20503
rect 27834 20469 28390 20503
rect 28852 20469 29408 20503
rect 29870 20469 30426 20503
rect 30888 20469 31444 20503
rect 31906 20469 32462 20503
rect 32924 20469 33480 20503
rect 14664 20021 14740 20055
rect 14882 20021 14958 20055
rect 15100 20021 15176 20055
rect 15318 20021 15394 20055
rect 15536 20021 15612 20055
rect 15754 20021 15830 20055
rect 15972 20021 16048 20055
rect 16190 20021 16266 20055
rect 16408 20021 16484 20055
rect 16626 20021 16702 20055
rect 18672 19741 19228 19775
rect 19690 19741 20246 19775
rect 20708 19741 21264 19775
rect 21726 19741 22282 19775
rect 22744 19741 23300 19775
rect 23762 19741 24318 19775
rect 24780 19741 25336 19775
rect 25798 19741 26354 19775
rect 26816 19741 27372 19775
rect 27834 19741 28390 19775
rect 28852 19741 29408 19775
rect 29870 19741 30426 19775
rect 30888 19741 31444 19775
rect 31906 19741 32462 19775
rect 32924 19741 33480 19775
rect 14664 19493 14740 19527
rect 14882 19493 14958 19527
rect 15100 19493 15176 19527
rect 15318 19493 15394 19527
rect 15536 19493 15612 19527
rect 15754 19493 15830 19527
rect 15972 19493 16048 19527
rect 16190 19493 16266 19527
rect 16408 19493 16484 19527
rect 16626 19493 16702 19527
rect 18672 19213 19228 19247
rect 19690 19213 20246 19247
rect 20708 19213 21264 19247
rect 21726 19213 22282 19247
rect 22744 19213 23300 19247
rect 23762 19213 24318 19247
rect 24780 19213 25336 19247
rect 25798 19213 26354 19247
rect 26816 19213 27372 19247
rect 27834 19213 28390 19247
rect 28852 19213 29408 19247
rect 29870 19213 30426 19247
rect 30888 19213 31444 19247
rect 31906 19213 32462 19247
rect 32924 19213 33480 19247
rect 14664 19083 14740 19117
rect 14882 19083 14958 19117
rect 15100 19083 15176 19117
rect 15318 19083 15394 19117
rect 15536 19083 15612 19117
rect 15754 19083 15830 19117
rect 15972 19083 16048 19117
rect 16190 19083 16266 19117
rect 16408 19083 16484 19117
rect 16626 19083 16702 19117
rect 14664 18555 14740 18589
rect 14882 18555 14958 18589
rect 15100 18555 15176 18589
rect 15318 18555 15394 18589
rect 15536 18555 15612 18589
rect 15754 18555 15830 18589
rect 15972 18555 16048 18589
rect 16190 18555 16266 18589
rect 16408 18555 16484 18589
rect 16626 18555 16702 18589
rect 18672 18485 19228 18519
rect 19690 18485 20246 18519
rect 20708 18485 21264 18519
rect 21726 18485 22282 18519
rect 22744 18485 23300 18519
rect 23762 18485 24318 18519
rect 24780 18485 25336 18519
rect 25798 18485 26354 18519
rect 26816 18485 27372 18519
rect 27834 18485 28390 18519
rect 28852 18485 29408 18519
rect 29870 18485 30426 18519
rect 30888 18485 31444 18519
rect 31906 18485 32462 18519
rect 32924 18485 33480 18519
rect 47474 25275 47574 25309
rect 47732 25275 47832 25309
rect 47990 25275 48090 25309
rect 48248 25275 48348 25309
rect 48506 25275 48606 25309
rect 48764 25275 48864 25309
rect 47474 24747 47574 24781
rect 47732 24747 47832 24781
rect 47990 24747 48090 24781
rect 48248 24747 48348 24781
rect 48506 24747 48606 24781
rect 48764 24747 48864 24781
rect 49310 24563 49344 24597
rect 47474 24342 47574 24376
rect 47732 24342 47832 24376
rect 47990 24342 48090 24376
rect 48248 24342 48348 24376
rect 48506 24342 48606 24376
rect 48764 24342 48864 24376
rect 47474 24032 47574 24066
rect 47732 24032 47832 24066
rect 47990 24032 48090 24066
rect 48248 24032 48348 24066
rect 48506 24032 48606 24066
rect 48764 24032 48864 24066
rect 47474 23275 47574 23309
rect 47732 23275 47832 23309
rect 47990 23275 48090 23309
rect 48248 23275 48348 23309
rect 48506 23275 48606 23309
rect 48764 23275 48864 23309
rect 47474 22747 47574 22781
rect 47732 22747 47832 22781
rect 47990 22747 48090 22781
rect 48248 22747 48348 22781
rect 48506 22747 48606 22781
rect 48764 22747 48864 22781
rect 49310 22563 49344 22597
rect 47474 22342 47574 22376
rect 47732 22342 47832 22376
rect 47990 22342 48090 22376
rect 48248 22342 48348 22376
rect 48506 22342 48606 22376
rect 48764 22342 48864 22376
rect 47474 22032 47574 22066
rect 47732 22032 47832 22066
rect 47990 22032 48090 22066
rect 48248 22032 48348 22066
rect 48506 22032 48606 22066
rect 48764 22032 48864 22066
rect 71686 27027 72242 27061
rect 72704 27027 73260 27061
rect 73722 27027 74278 27061
rect 74740 27027 75296 27061
rect 75758 27027 76314 27061
rect 76776 27027 77332 27061
rect 77794 27027 78350 27061
rect 78812 27027 79368 27061
rect 79830 27027 80386 27061
rect 80848 27027 81404 27061
rect 81866 27027 82422 27061
rect 82884 27027 83440 27061
rect 83902 27027 84458 27061
rect 84920 27027 85476 27061
rect 85938 27027 86494 27061
rect 86956 27027 87512 27061
rect 71686 26299 72242 26333
rect 72704 26299 73260 26333
rect 73722 26299 74278 26333
rect 74740 26299 75296 26333
rect 75758 26299 76314 26333
rect 76776 26299 77332 26333
rect 77794 26299 78350 26333
rect 78812 26299 79368 26333
rect 79830 26299 80386 26333
rect 80848 26299 81404 26333
rect 81866 26299 82422 26333
rect 82884 26299 83440 26333
rect 83902 26299 84458 26333
rect 84920 26299 85476 26333
rect 85938 26299 86494 26333
rect 86956 26299 87512 26333
rect 71686 25891 72242 25925
rect 72704 25891 73260 25925
rect 73722 25891 74278 25925
rect 74740 25891 75296 25925
rect 75758 25891 76314 25925
rect 76776 25891 77332 25925
rect 77794 25891 78350 25925
rect 78812 25891 79368 25925
rect 79830 25891 80386 25925
rect 80848 25891 81404 25925
rect 81866 25891 82422 25925
rect 82884 25891 83440 25925
rect 83902 25891 84458 25925
rect 84920 25891 85476 25925
rect 85938 25891 86494 25925
rect 86956 25891 87512 25925
rect 71686 25163 72242 25197
rect 72704 25163 73260 25197
rect 73722 25163 74278 25197
rect 74740 25163 75296 25197
rect 75758 25163 76314 25197
rect 76776 25163 77332 25197
rect 77794 25163 78350 25197
rect 78812 25163 79368 25197
rect 79830 25163 80386 25197
rect 80848 25163 81404 25197
rect 81866 25163 82422 25197
rect 82884 25163 83440 25197
rect 83902 25163 84458 25197
rect 84920 25163 85476 25197
rect 85938 25163 86494 25197
rect 86956 25163 87512 25197
rect 71686 24755 72242 24789
rect 72704 24755 73260 24789
rect 73722 24755 74278 24789
rect 74740 24755 75296 24789
rect 75758 24755 76314 24789
rect 76776 24755 77332 24789
rect 77794 24755 78350 24789
rect 78812 24755 79368 24789
rect 79830 24755 80386 24789
rect 80848 24755 81404 24789
rect 81866 24755 82422 24789
rect 82884 24755 83440 24789
rect 83902 24755 84458 24789
rect 84920 24755 85476 24789
rect 85938 24755 86494 24789
rect 86956 24755 87512 24789
rect 71686 24027 72242 24061
rect 72704 24027 73260 24061
rect 73722 24027 74278 24061
rect 74740 24027 75296 24061
rect 75758 24027 76314 24061
rect 76776 24027 77332 24061
rect 77794 24027 78350 24061
rect 78812 24027 79368 24061
rect 79830 24027 80386 24061
rect 80848 24027 81404 24061
rect 81866 24027 82422 24061
rect 82884 24027 83440 24061
rect 83902 24027 84458 24061
rect 84920 24027 85476 24061
rect 85938 24027 86494 24061
rect 86956 24027 87512 24061
rect 72672 22981 73228 23015
rect 73690 22981 74246 23015
rect 74708 22981 75264 23015
rect 75726 22981 76282 23015
rect 76744 22981 77300 23015
rect 77762 22981 78318 23015
rect 78780 22981 79336 23015
rect 79798 22981 80354 23015
rect 80816 22981 81372 23015
rect 81834 22981 82390 23015
rect 82852 22981 83408 23015
rect 83870 22981 84426 23015
rect 84888 22981 85444 23015
rect 85906 22981 86462 23015
rect 86924 22981 87480 23015
rect 72672 22253 73228 22287
rect 73690 22253 74246 22287
rect 74708 22253 75264 22287
rect 75726 22253 76282 22287
rect 76744 22253 77300 22287
rect 77762 22253 78318 22287
rect 78780 22253 79336 22287
rect 79798 22253 80354 22287
rect 80816 22253 81372 22287
rect 81834 22253 82390 22287
rect 82852 22253 83408 22287
rect 83870 22253 84426 22287
rect 84888 22253 85444 22287
rect 85906 22253 86462 22287
rect 86924 22253 87480 22287
rect 68664 21897 68740 21931
rect 68882 21897 68958 21931
rect 69100 21897 69176 21931
rect 69318 21897 69394 21931
rect 69536 21897 69612 21931
rect 69754 21897 69830 21931
rect 69972 21897 70048 21931
rect 70190 21897 70266 21931
rect 70408 21897 70484 21931
rect 70626 21897 70702 21931
rect 72672 21725 73228 21759
rect 73690 21725 74246 21759
rect 74708 21725 75264 21759
rect 75726 21725 76282 21759
rect 76744 21725 77300 21759
rect 77762 21725 78318 21759
rect 78780 21725 79336 21759
rect 79798 21725 80354 21759
rect 80816 21725 81372 21759
rect 81834 21725 82390 21759
rect 82852 21725 83408 21759
rect 83870 21725 84426 21759
rect 84888 21725 85444 21759
rect 85906 21725 86462 21759
rect 86924 21725 87480 21759
rect 68664 21369 68740 21403
rect 68882 21369 68958 21403
rect 69100 21369 69176 21403
rect 69318 21369 69394 21403
rect 69536 21369 69612 21403
rect 69754 21369 69830 21403
rect 69972 21369 70048 21403
rect 70190 21369 70266 21403
rect 70408 21369 70484 21403
rect 70626 21369 70702 21403
rect 68664 20959 68740 20993
rect 68882 20959 68958 20993
rect 69100 20959 69176 20993
rect 69318 20959 69394 20993
rect 69536 20959 69612 20993
rect 69754 20959 69830 20993
rect 69972 20959 70048 20993
rect 70190 20959 70266 20993
rect 70408 20959 70484 20993
rect 70626 20959 70702 20993
rect 72672 20997 73228 21031
rect 73690 20997 74246 21031
rect 74708 20997 75264 21031
rect 75726 20997 76282 21031
rect 76744 20997 77300 21031
rect 77762 20997 78318 21031
rect 78780 20997 79336 21031
rect 79798 20997 80354 21031
rect 80816 20997 81372 21031
rect 81834 20997 82390 21031
rect 82852 20997 83408 21031
rect 83870 20997 84426 21031
rect 84888 20997 85444 21031
rect 85906 20997 86462 21031
rect 86924 20997 87480 21031
rect 68664 20431 68740 20465
rect 68882 20431 68958 20465
rect 69100 20431 69176 20465
rect 69318 20431 69394 20465
rect 69536 20431 69612 20465
rect 69754 20431 69830 20465
rect 69972 20431 70048 20465
rect 70190 20431 70266 20465
rect 70408 20431 70484 20465
rect 70626 20431 70702 20465
rect 72672 20469 73228 20503
rect 73690 20469 74246 20503
rect 74708 20469 75264 20503
rect 75726 20469 76282 20503
rect 76744 20469 77300 20503
rect 77762 20469 78318 20503
rect 78780 20469 79336 20503
rect 79798 20469 80354 20503
rect 80816 20469 81372 20503
rect 81834 20469 82390 20503
rect 82852 20469 83408 20503
rect 83870 20469 84426 20503
rect 84888 20469 85444 20503
rect 85906 20469 86462 20503
rect 86924 20469 87480 20503
rect 68664 20021 68740 20055
rect 68882 20021 68958 20055
rect 69100 20021 69176 20055
rect 69318 20021 69394 20055
rect 69536 20021 69612 20055
rect 69754 20021 69830 20055
rect 69972 20021 70048 20055
rect 70190 20021 70266 20055
rect 70408 20021 70484 20055
rect 70626 20021 70702 20055
rect 72672 19741 73228 19775
rect 73690 19741 74246 19775
rect 74708 19741 75264 19775
rect 75726 19741 76282 19775
rect 76744 19741 77300 19775
rect 77762 19741 78318 19775
rect 78780 19741 79336 19775
rect 79798 19741 80354 19775
rect 80816 19741 81372 19775
rect 81834 19741 82390 19775
rect 82852 19741 83408 19775
rect 83870 19741 84426 19775
rect 84888 19741 85444 19775
rect 85906 19741 86462 19775
rect 86924 19741 87480 19775
rect 68664 19493 68740 19527
rect 68882 19493 68958 19527
rect 69100 19493 69176 19527
rect 69318 19493 69394 19527
rect 69536 19493 69612 19527
rect 69754 19493 69830 19527
rect 69972 19493 70048 19527
rect 70190 19493 70266 19527
rect 70408 19493 70484 19527
rect 70626 19493 70702 19527
rect 72672 19213 73228 19247
rect 73690 19213 74246 19247
rect 74708 19213 75264 19247
rect 75726 19213 76282 19247
rect 76744 19213 77300 19247
rect 77762 19213 78318 19247
rect 78780 19213 79336 19247
rect 79798 19213 80354 19247
rect 80816 19213 81372 19247
rect 81834 19213 82390 19247
rect 82852 19213 83408 19247
rect 83870 19213 84426 19247
rect 84888 19213 85444 19247
rect 85906 19213 86462 19247
rect 86924 19213 87480 19247
rect 68664 19083 68740 19117
rect 68882 19083 68958 19117
rect 69100 19083 69176 19117
rect 69318 19083 69394 19117
rect 69536 19083 69612 19117
rect 69754 19083 69830 19117
rect 69972 19083 70048 19117
rect 70190 19083 70266 19117
rect 70408 19083 70484 19117
rect 70626 19083 70702 19117
rect 68664 18555 68740 18589
rect 68882 18555 68958 18589
rect 69100 18555 69176 18589
rect 69318 18555 69394 18589
rect 69536 18555 69612 18589
rect 69754 18555 69830 18589
rect 69972 18555 70048 18589
rect 70190 18555 70266 18589
rect 70408 18555 70484 18589
rect 70626 18555 70702 18589
rect 72672 18485 73228 18519
rect 73690 18485 74246 18519
rect 74708 18485 75264 18519
rect 75726 18485 76282 18519
rect 76744 18485 77300 18519
rect 77762 18485 78318 18519
rect 78780 18485 79336 18519
rect 79798 18485 80354 18519
rect 80816 18485 81372 18519
rect 81834 18485 82390 18519
rect 82852 18485 83408 18519
rect 83870 18485 84426 18519
rect 84888 18485 85444 18519
rect 85906 18485 86462 18519
rect 86924 18485 87480 18519
rect -12884 16145 -12784 16179
rect -12626 16145 -12526 16179
rect -12368 16145 -12268 16179
rect -12110 16145 -12010 16179
rect -11852 16145 -11752 16179
rect -11594 16145 -11494 16179
rect -12884 15617 -12784 15651
rect -12626 15617 -12526 15651
rect -12368 15617 -12268 15651
rect -12110 15617 -12010 15651
rect -11852 15617 -11752 15651
rect -11594 15617 -11494 15651
rect -10284 16145 -10184 16179
rect -10026 16145 -9926 16179
rect -9768 16145 -9668 16179
rect -9510 16145 -9410 16179
rect -9252 16145 -9152 16179
rect -8994 16145 -8894 16179
rect -10284 15617 -10184 15651
rect -10026 15617 -9926 15651
rect -9768 15617 -9668 15651
rect -9510 15617 -9410 15651
rect -9252 15617 -9152 15651
rect -8994 15617 -8894 15651
rect -11048 15433 -11014 15467
rect -8448 15433 -8414 15467
rect -7948 15433 -7914 15467
rect -12884 15212 -12784 15246
rect -12626 15212 -12526 15246
rect -12368 15212 -12268 15246
rect -12110 15212 -12010 15246
rect -11852 15212 -11752 15246
rect -11594 15212 -11494 15246
rect -12884 14902 -12784 14936
rect -12626 14902 -12526 14936
rect -12368 14902 -12268 14936
rect -12110 14902 -12010 14936
rect -11852 14902 -11752 14936
rect -11594 14902 -11494 14936
rect -10284 15212 -10184 15246
rect -10026 15212 -9926 15246
rect -9768 15212 -9668 15246
rect -9510 15212 -9410 15246
rect -9252 15212 -9152 15246
rect -8994 15212 -8894 15246
rect -10284 14902 -10184 14936
rect -10026 14902 -9926 14936
rect -9768 14902 -9668 14936
rect -9510 14902 -9410 14936
rect -9252 14902 -9152 14936
rect -8994 14902 -8894 14936
rect 13780 14860 14336 14894
rect 14798 14860 15354 14894
rect 15816 14860 16372 14894
rect 16834 14860 17390 14894
rect 17852 14860 18408 14894
rect 18870 14860 19426 14894
rect 19888 14860 20444 14894
rect 20906 14860 21462 14894
rect 21924 14860 22480 14894
rect 22942 14860 23498 14894
rect 23960 14860 24516 14894
rect 24978 14860 25534 14894
rect 25996 14860 26552 14894
rect 27014 14860 27570 14894
rect 28032 14860 28588 14894
rect 29050 14860 29606 14894
rect 30068 14860 30624 14894
rect 31086 14860 31642 14894
rect 32104 14860 32660 14894
rect 33122 14860 33678 14894
rect 13780 14150 14336 14184
rect 14798 14150 15354 14184
rect 15816 14150 16372 14184
rect 16834 14150 17390 14184
rect 17852 14150 18408 14184
rect 18870 14150 19426 14184
rect 19888 14150 20444 14184
rect 20906 14150 21462 14184
rect 21924 14150 22480 14184
rect 22942 14150 23498 14184
rect 23960 14150 24516 14184
rect 24978 14150 25534 14184
rect 25996 14150 26552 14184
rect 27014 14150 27570 14184
rect 28032 14150 28588 14184
rect 29050 14150 29606 14184
rect 30068 14150 30624 14184
rect 31086 14150 31642 14184
rect 32104 14150 32660 14184
rect 33122 14150 33678 14184
rect 2014 14066 2570 14100
rect 3032 14066 3588 14100
rect 4050 14066 4606 14100
rect 5068 14066 5624 14100
rect 6086 14066 6642 14100
rect 7104 14066 7660 14100
rect 8122 14066 8678 14100
rect 9140 14066 9696 14100
rect 10158 14066 10714 14100
rect 13780 13626 14336 13660
rect 14798 13626 15354 13660
rect 15816 13626 16372 13660
rect 16834 13626 17390 13660
rect 17852 13626 18408 13660
rect 18870 13626 19426 13660
rect 19888 13626 20444 13660
rect 20906 13626 21462 13660
rect 21924 13626 22480 13660
rect 22942 13626 23498 13660
rect 23960 13626 24516 13660
rect 24978 13626 25534 13660
rect 25996 13626 26552 13660
rect 27014 13626 27570 13660
rect 28032 13626 28588 13660
rect 29050 13626 29606 13660
rect 30068 13626 30624 13660
rect 31086 13626 31642 13660
rect 32104 13626 32660 13660
rect 33122 13626 33678 13660
rect 2014 13356 2570 13390
rect 3032 13356 3588 13390
rect 2014 13248 2570 13282
rect 4050 13356 4606 13390
rect 3032 13248 3588 13282
rect 5068 13356 5624 13390
rect 4050 13248 4606 13282
rect 6086 13356 6642 13390
rect 5068 13248 5624 13282
rect 7104 13356 7660 13390
rect 6086 13248 6642 13282
rect 8122 13356 8678 13390
rect 7104 13248 7660 13282
rect 9140 13356 9696 13390
rect 8122 13248 8678 13282
rect 10158 13356 10714 13390
rect 9140 13248 9696 13282
rect 10158 13248 10714 13282
rect 13780 12916 14336 12950
rect 14798 12916 15354 12950
rect 15816 12916 16372 12950
rect 16834 12916 17390 12950
rect 17852 12916 18408 12950
rect 18870 12916 19426 12950
rect 19888 12916 20444 12950
rect 20906 12916 21462 12950
rect 21924 12916 22480 12950
rect 22942 12916 23498 12950
rect 23960 12916 24516 12950
rect 24978 12916 25534 12950
rect 25996 12916 26552 12950
rect 27014 12916 27570 12950
rect 28032 12916 28588 12950
rect 29050 12916 29606 12950
rect 30068 12916 30624 12950
rect 31086 12916 31642 12950
rect 32104 12916 32660 12950
rect 33122 12916 33678 12950
rect 2014 12538 2570 12572
rect 3032 12538 3588 12572
rect 2014 12430 2570 12464
rect 4050 12538 4606 12572
rect 3032 12430 3588 12464
rect 5068 12538 5624 12572
rect 4050 12430 4606 12464
rect 6086 12538 6642 12572
rect 5068 12430 5624 12464
rect 7104 12538 7660 12572
rect 6086 12430 6642 12464
rect 8122 12538 8678 12572
rect 7104 12430 7660 12464
rect 9140 12538 9696 12572
rect 8122 12430 8678 12464
rect 10158 12538 10714 12572
rect 9140 12430 9696 12464
rect 10158 12430 10714 12464
rect 13780 12394 14336 12428
rect 14798 12394 15354 12428
rect 15816 12394 16372 12428
rect 16834 12394 17390 12428
rect 17852 12394 18408 12428
rect 18870 12394 19426 12428
rect 19888 12394 20444 12428
rect 20906 12394 21462 12428
rect 21924 12394 22480 12428
rect 22942 12394 23498 12428
rect 23960 12394 24516 12428
rect 24978 12394 25534 12428
rect 25996 12394 26552 12428
rect 27014 12394 27570 12428
rect 28032 12394 28588 12428
rect 29050 12394 29606 12428
rect 30068 12394 30624 12428
rect 31086 12394 31642 12428
rect 32104 12394 32660 12428
rect 33122 12394 33678 12428
rect 2014 11720 2570 11754
rect 3032 11720 3588 11754
rect 2014 11612 2570 11646
rect 4050 11720 4606 11754
rect 3032 11612 3588 11646
rect 5068 11720 5624 11754
rect 4050 11612 4606 11646
rect 6086 11720 6642 11754
rect 5068 11612 5624 11646
rect 7104 11720 7660 11754
rect 6086 11612 6642 11646
rect 8122 11720 8678 11754
rect 7104 11612 7660 11646
rect 9140 11720 9696 11754
rect 8122 11612 8678 11646
rect 10158 11720 10714 11754
rect 9140 11612 9696 11646
rect 13780 11684 14336 11718
rect 14798 11684 15354 11718
rect 15816 11684 16372 11718
rect 16834 11684 17390 11718
rect 17852 11684 18408 11718
rect 18870 11684 19426 11718
rect 19888 11684 20444 11718
rect 20906 11684 21462 11718
rect 21924 11684 22480 11718
rect 22942 11684 23498 11718
rect 23960 11684 24516 11718
rect 24978 11684 25534 11718
rect 25996 11684 26552 11718
rect 27014 11684 27570 11718
rect 28032 11684 28588 11718
rect 29050 11684 29606 11718
rect 30068 11684 30624 11718
rect 31086 11684 31642 11718
rect 32104 11684 32660 11718
rect 33122 11684 33678 11718
rect 10158 11612 10714 11646
rect 13778 11160 14334 11194
rect 14796 11160 15352 11194
rect 15814 11160 16370 11194
rect 16832 11160 17388 11194
rect 17850 11160 18406 11194
rect 18868 11160 19424 11194
rect 19886 11160 20442 11194
rect 20904 11160 21460 11194
rect 21922 11160 22478 11194
rect 22940 11160 23496 11194
rect 23958 11160 24514 11194
rect 24976 11160 25532 11194
rect 25994 11160 26550 11194
rect 27012 11160 27568 11194
rect 28030 11160 28586 11194
rect 29048 11160 29604 11194
rect 30066 11160 30622 11194
rect 31084 11160 31640 11194
rect 32102 11160 32658 11194
rect 33120 11160 33676 11194
rect 2014 10902 2570 10936
rect 3032 10902 3588 10936
rect 2014 10794 2570 10828
rect 4050 10902 4606 10936
rect 3032 10794 3588 10828
rect 5068 10902 5624 10936
rect 4050 10794 4606 10828
rect 6086 10902 6642 10936
rect 5068 10794 5624 10828
rect 7104 10902 7660 10936
rect 6086 10794 6642 10828
rect 8122 10902 8678 10936
rect 7104 10794 7660 10828
rect 9140 10902 9696 10936
rect 8122 10794 8678 10828
rect 10158 10902 10714 10936
rect 9140 10794 9696 10828
rect 10158 10794 10714 10828
rect 13778 10450 14334 10484
rect 14796 10450 15352 10484
rect 15814 10450 16370 10484
rect 16832 10450 17388 10484
rect 17850 10450 18406 10484
rect 18868 10450 19424 10484
rect 19886 10450 20442 10484
rect 20904 10450 21460 10484
rect 21922 10450 22478 10484
rect 22940 10450 23496 10484
rect 23958 10450 24514 10484
rect 24976 10450 25532 10484
rect 25994 10450 26550 10484
rect 27012 10450 27568 10484
rect 28030 10450 28586 10484
rect 29048 10450 29604 10484
rect 30066 10450 30622 10484
rect 31084 10450 31640 10484
rect 32102 10450 32658 10484
rect 33120 10450 33676 10484
rect 2014 10084 2570 10118
rect 3032 10084 3588 10118
rect 2014 9976 2570 10010
rect 4050 10084 4606 10118
rect 3032 9976 3588 10010
rect 5068 10084 5624 10118
rect 4050 9976 4606 10010
rect 6086 10084 6642 10118
rect 5068 9976 5624 10010
rect 7104 10084 7660 10118
rect 6086 9976 6642 10010
rect 8122 10084 8678 10118
rect 7104 9976 7660 10010
rect 9140 10084 9696 10118
rect 8122 9976 8678 10010
rect 10158 10084 10714 10118
rect 9140 9976 9696 10010
rect 10158 9976 10714 10010
rect 13778 9926 14334 9960
rect 14796 9926 15352 9960
rect 15814 9926 16370 9960
rect 16832 9926 17388 9960
rect 17850 9926 18406 9960
rect 18868 9926 19424 9960
rect 19886 9926 20442 9960
rect 20904 9926 21460 9960
rect 21922 9926 22478 9960
rect 22940 9926 23496 9960
rect 23958 9926 24514 9960
rect 24976 9926 25532 9960
rect 25994 9926 26550 9960
rect 27012 9926 27568 9960
rect 28030 9926 28586 9960
rect 29048 9926 29604 9960
rect 30066 9926 30622 9960
rect 31084 9926 31640 9960
rect 32102 9926 32658 9960
rect 33120 9926 33676 9960
rect 2014 9266 2570 9300
rect 3032 9266 3588 9300
rect 2014 9158 2570 9192
rect 4050 9266 4606 9300
rect 3032 9158 3588 9192
rect 5068 9266 5624 9300
rect 4050 9158 4606 9192
rect 6086 9266 6642 9300
rect 5068 9158 5624 9192
rect 7104 9266 7660 9300
rect 6086 9158 6642 9192
rect 8122 9266 8678 9300
rect 7104 9158 7660 9192
rect 9140 9266 9696 9300
rect 8122 9158 8678 9192
rect 10158 9266 10714 9300
rect 9140 9158 9696 9192
rect 10158 9158 10714 9192
rect 13778 9216 14334 9250
rect 14796 9216 15352 9250
rect 15814 9216 16370 9250
rect 16832 9216 17388 9250
rect 17850 9216 18406 9250
rect 18868 9216 19424 9250
rect 19886 9216 20442 9250
rect 20904 9216 21460 9250
rect 21922 9216 22478 9250
rect 22940 9216 23496 9250
rect 23958 9216 24514 9250
rect 24976 9216 25532 9250
rect 25994 9216 26550 9250
rect 27012 9216 27568 9250
rect 28030 9216 28586 9250
rect 29048 9216 29604 9250
rect 30066 9216 30622 9250
rect 31084 9216 31640 9250
rect 32102 9216 32658 9250
rect 33120 9216 33676 9250
rect 13778 8694 14334 8728
rect 14796 8694 15352 8728
rect 15814 8694 16370 8728
rect 16832 8694 17388 8728
rect 17850 8694 18406 8728
rect 18868 8694 19424 8728
rect 19886 8694 20442 8728
rect 20904 8694 21460 8728
rect 21922 8694 22478 8728
rect 22940 8694 23496 8728
rect 23958 8694 24514 8728
rect 24976 8694 25532 8728
rect 25994 8694 26550 8728
rect 27012 8694 27568 8728
rect 28030 8694 28586 8728
rect 29048 8694 29604 8728
rect 30066 8694 30622 8728
rect 31084 8694 31640 8728
rect 32102 8694 32658 8728
rect 33120 8694 33676 8728
rect 2014 8448 2570 8482
rect 3032 8448 3588 8482
rect 2014 8340 2570 8374
rect 4050 8448 4606 8482
rect 3032 8340 3588 8374
rect 5068 8448 5624 8482
rect 4050 8340 4606 8374
rect 6086 8448 6642 8482
rect 5068 8340 5624 8374
rect 7104 8448 7660 8482
rect 6086 8340 6642 8374
rect 8122 8448 8678 8482
rect 7104 8340 7660 8374
rect 9140 8448 9696 8482
rect 8122 8340 8678 8374
rect 10158 8448 10714 8482
rect 9140 8340 9696 8374
rect 10158 8340 10714 8374
rect 13778 7984 14334 8018
rect 14796 7984 15352 8018
rect 15814 7984 16370 8018
rect 16832 7984 17388 8018
rect 17850 7984 18406 8018
rect 18868 7984 19424 8018
rect 19886 7984 20442 8018
rect 20904 7984 21460 8018
rect 21922 7984 22478 8018
rect 22940 7984 23496 8018
rect 23958 7984 24514 8018
rect 24976 7984 25532 8018
rect 25994 7984 26550 8018
rect 27012 7984 27568 8018
rect 28030 7984 28586 8018
rect 29048 7984 29604 8018
rect 30066 7984 30622 8018
rect 31084 7984 31640 8018
rect 32102 7984 32658 8018
rect 33120 7984 33676 8018
rect 2014 7630 2570 7664
rect 3032 7630 3588 7664
rect 4050 7630 4606 7664
rect 5068 7630 5624 7664
rect 6086 7630 6642 7664
rect 7104 7630 7660 7664
rect 8122 7630 8678 7664
rect 9140 7630 9696 7664
rect 10158 7630 10714 7664
rect 13778 7460 14334 7494
rect 14796 7460 15352 7494
rect 15814 7460 16370 7494
rect 16832 7460 17388 7494
rect 17850 7460 18406 7494
rect 18868 7460 19424 7494
rect 19886 7460 20442 7494
rect 20904 7460 21460 7494
rect 21922 7460 22478 7494
rect 22940 7460 23496 7494
rect 23958 7460 24514 7494
rect 24976 7460 25532 7494
rect 25994 7460 26550 7494
rect 27012 7460 27568 7494
rect 28030 7460 28586 7494
rect 29048 7460 29604 7494
rect 30066 7460 30622 7494
rect 31084 7460 31640 7494
rect 32102 7460 32658 7494
rect 33120 7460 33676 7494
rect 8714 6956 8790 6990
rect 8932 6956 9008 6990
rect 9150 6956 9226 6990
rect 9368 6956 9444 6990
rect 9586 6956 9662 6990
rect 9804 6956 9880 6990
rect 10022 6956 10098 6990
rect 10240 6956 10316 6990
rect 10458 6956 10534 6990
rect 10676 6956 10752 6990
rect 13778 6750 14334 6784
rect 14796 6750 15352 6784
rect 15814 6750 16370 6784
rect 16832 6750 17388 6784
rect 17850 6750 18406 6784
rect 18868 6750 19424 6784
rect 19886 6750 20442 6784
rect 20904 6750 21460 6784
rect 21922 6750 22478 6784
rect 22940 6750 23496 6784
rect 23958 6750 24514 6784
rect 24976 6750 25532 6784
rect 25994 6750 26550 6784
rect 27012 6750 27568 6784
rect 28030 6750 28586 6784
rect 29048 6750 29604 6784
rect 30066 6750 30622 6784
rect 31084 6750 31640 6784
rect 32102 6750 32658 6784
rect 33120 6750 33676 6784
rect 8714 6646 8790 6680
rect 8932 6646 9008 6680
rect 9150 6646 9226 6680
rect 9368 6646 9444 6680
rect 9586 6646 9662 6680
rect 9804 6646 9880 6680
rect 10022 6646 10098 6680
rect 10240 6646 10316 6680
rect 10458 6646 10534 6680
rect 10676 6646 10752 6680
rect 13778 6226 14334 6260
rect 14796 6226 15352 6260
rect 15814 6226 16370 6260
rect 16832 6226 17388 6260
rect 17850 6226 18406 6260
rect 18868 6226 19424 6260
rect 19886 6226 20442 6260
rect 20904 6226 21460 6260
rect 21922 6226 22478 6260
rect 22940 6226 23496 6260
rect 23958 6226 24514 6260
rect 24976 6226 25532 6260
rect 25994 6226 26550 6260
rect 27012 6226 27568 6260
rect 28030 6226 28586 6260
rect 29048 6226 29604 6260
rect 30066 6226 30622 6260
rect 31084 6226 31640 6260
rect 32102 6226 32658 6260
rect 33120 6226 33676 6260
rect 8714 6124 8790 6158
rect 8932 6124 9008 6158
rect 9150 6124 9226 6158
rect 9368 6124 9444 6158
rect 9586 6124 9662 6158
rect 9804 6124 9880 6158
rect 10022 6124 10098 6158
rect 10240 6124 10316 6158
rect 10458 6124 10534 6158
rect 10676 6124 10752 6158
rect 8714 5814 8790 5848
rect 8932 5814 9008 5848
rect 9150 5814 9226 5848
rect 9368 5814 9444 5848
rect 9586 5814 9662 5848
rect 9804 5814 9880 5848
rect 10022 5814 10098 5848
rect 10240 5814 10316 5848
rect 10458 5814 10534 5848
rect 10676 5814 10752 5848
rect 13778 5516 14334 5550
rect 14796 5516 15352 5550
rect 15814 5516 16370 5550
rect 16832 5516 17388 5550
rect 17850 5516 18406 5550
rect 18868 5516 19424 5550
rect 19886 5516 20442 5550
rect 20904 5516 21460 5550
rect 21922 5516 22478 5550
rect 22940 5516 23496 5550
rect 23958 5516 24514 5550
rect 24976 5516 25532 5550
rect 25994 5516 26550 5550
rect 27012 5516 27568 5550
rect 28030 5516 28586 5550
rect 29048 5516 29604 5550
rect 30066 5516 30622 5550
rect 31084 5516 31640 5550
rect 32102 5516 32658 5550
rect 33120 5516 33676 5550
rect 13778 4994 14334 5028
rect 14796 4994 15352 5028
rect 15814 4994 16370 5028
rect 16832 4994 17388 5028
rect 17850 4994 18406 5028
rect 18868 4994 19424 5028
rect 19886 4994 20442 5028
rect 20904 4994 21460 5028
rect 21922 4994 22478 5028
rect 22940 4994 23496 5028
rect 23958 4994 24514 5028
rect 24976 4994 25532 5028
rect 25994 4994 26550 5028
rect 27012 4994 27568 5028
rect 28030 4994 28586 5028
rect 29048 4994 29604 5028
rect 30066 4994 30622 5028
rect 31084 4994 31640 5028
rect 32102 4994 32658 5028
rect 33120 4994 33676 5028
rect 1793 4797 2349 4831
rect 2811 4797 3367 4831
rect 3829 4797 4385 4831
rect 4847 4797 5403 4831
rect 5865 4797 6421 4831
rect 6883 4797 7439 4831
rect 8644 4798 8768 4832
rect 8942 4798 9066 4832
rect 9240 4798 9364 4832
rect 9538 4798 9662 4832
rect 9836 4798 9960 4832
rect 10134 4798 10258 4832
rect 10432 4798 10556 4832
rect 10730 4798 10854 4832
rect 11028 4798 11152 4832
rect 11326 4798 11450 4832
rect 11624 4798 11748 4832
rect 13778 4284 14334 4318
rect 14796 4284 15352 4318
rect 15814 4284 16370 4318
rect 16832 4284 17388 4318
rect 17850 4284 18406 4318
rect 18868 4284 19424 4318
rect 19886 4284 20442 4318
rect 20904 4284 21460 4318
rect 21922 4284 22478 4318
rect 22940 4284 23496 4318
rect 23958 4284 24514 4318
rect 24976 4284 25532 4318
rect 25994 4284 26550 4318
rect 27012 4284 27568 4318
rect 28030 4284 28586 4318
rect 29048 4284 29604 4318
rect 30066 4284 30622 4318
rect 31084 4284 31640 4318
rect 32102 4284 32658 4318
rect 33120 4284 33676 4318
rect 1793 4087 2349 4121
rect 2811 4087 3367 4121
rect 3829 4087 4385 4121
rect 4847 4087 5403 4121
rect 5865 4087 6421 4121
rect 6883 4087 7439 4121
rect 8644 4088 8768 4122
rect 8942 4088 9066 4122
rect 9240 4088 9364 4122
rect 9538 4088 9662 4122
rect 9836 4088 9960 4122
rect 10134 4088 10258 4122
rect 10432 4088 10556 4122
rect 10730 4088 10854 4122
rect 11028 4088 11152 4122
rect 11326 4088 11450 4122
rect 11624 4088 11748 4122
rect 13778 3760 14334 3794
rect 1792 3684 2348 3718
rect 2810 3684 3366 3718
rect 3828 3684 4384 3718
rect 4846 3684 5402 3718
rect 5864 3684 6420 3718
rect 6882 3684 7438 3718
rect 8644 3686 8768 3720
rect 8942 3686 9066 3720
rect 9240 3686 9364 3720
rect 9538 3686 9662 3720
rect 9836 3686 9960 3720
rect 10134 3686 10258 3720
rect 10432 3686 10556 3720
rect 10730 3686 10854 3720
rect 11028 3686 11152 3720
rect 11326 3686 11450 3720
rect 14796 3760 15352 3794
rect 15814 3760 16370 3794
rect 16832 3760 17388 3794
rect 17850 3760 18406 3794
rect 18868 3760 19424 3794
rect 19886 3760 20442 3794
rect 20904 3760 21460 3794
rect 21922 3760 22478 3794
rect 22940 3760 23496 3794
rect 23958 3760 24514 3794
rect 24976 3760 25532 3794
rect 25994 3760 26550 3794
rect 27012 3760 27568 3794
rect 28030 3760 28586 3794
rect 29048 3760 29604 3794
rect 30066 3760 30622 3794
rect 31084 3760 31640 3794
rect 32102 3760 32658 3794
rect 33120 3760 33676 3794
rect 11624 3686 11748 3720
rect 13778 3050 14334 3084
rect 1792 2974 2348 3008
rect 2810 2974 3366 3008
rect 3828 2974 4384 3008
rect 4846 2974 5402 3008
rect 5864 2974 6420 3008
rect 6882 2974 7438 3008
rect 8644 2976 8768 3010
rect 8942 2976 9066 3010
rect 9240 2976 9364 3010
rect 9538 2976 9662 3010
rect 9836 2976 9960 3010
rect 10134 2976 10258 3010
rect 10432 2976 10556 3010
rect 10730 2976 10854 3010
rect 11028 2976 11152 3010
rect 11326 2976 11450 3010
rect 14796 3050 15352 3084
rect 15814 3050 16370 3084
rect 16832 3050 17388 3084
rect 17850 3050 18406 3084
rect 18868 3050 19424 3084
rect 19886 3050 20442 3084
rect 20904 3050 21460 3084
rect 21922 3050 22478 3084
rect 22940 3050 23496 3084
rect 23958 3050 24514 3084
rect 24976 3050 25532 3084
rect 25994 3050 26550 3084
rect 27012 3050 27568 3084
rect 28030 3050 28586 3084
rect 29048 3050 29604 3084
rect 30066 3050 30622 3084
rect 31084 3050 31640 3084
rect 32102 3050 32658 3084
rect 33120 3050 33676 3084
rect 11624 2976 11748 3010
rect 1793 2573 2349 2607
rect 2811 2573 3367 2607
rect 3829 2573 4385 2607
rect 4847 2573 5403 2607
rect 5865 2573 6421 2607
rect 6883 2573 7439 2607
rect 8642 2574 8766 2608
rect 8940 2574 9064 2608
rect 9238 2574 9362 2608
rect 9536 2574 9660 2608
rect 9834 2574 9958 2608
rect 10132 2574 10256 2608
rect 10430 2574 10554 2608
rect 10728 2574 10852 2608
rect 11026 2574 11150 2608
rect 11324 2574 11448 2608
rect 11622 2574 11746 2608
rect 13778 2526 14334 2560
rect 14796 2526 15352 2560
rect 15814 2526 16370 2560
rect 16832 2526 17388 2560
rect 17850 2526 18406 2560
rect 18868 2526 19424 2560
rect 19886 2526 20442 2560
rect 20904 2526 21460 2560
rect 21922 2526 22478 2560
rect 22940 2526 23496 2560
rect 23958 2526 24514 2560
rect 24976 2526 25532 2560
rect 25994 2526 26550 2560
rect 27012 2526 27568 2560
rect 28030 2526 28586 2560
rect 29048 2526 29604 2560
rect 30066 2526 30622 2560
rect 31084 2526 31640 2560
rect 32102 2526 32658 2560
rect 33120 2526 33676 2560
rect 1793 1863 2349 1897
rect 2811 1863 3367 1897
rect 3829 1863 4385 1897
rect 4847 1863 5403 1897
rect 5865 1863 6421 1897
rect 6883 1863 7439 1897
rect 8642 1864 8766 1898
rect 8940 1864 9064 1898
rect 9238 1864 9362 1898
rect 9536 1864 9660 1898
rect 9834 1864 9958 1898
rect 10132 1864 10256 1898
rect 10430 1864 10554 1898
rect 10728 1864 10852 1898
rect 11026 1864 11150 1898
rect 11324 1864 11448 1898
rect 11622 1864 11746 1898
rect 13778 1816 14334 1850
rect 14796 1816 15352 1850
rect 15814 1816 16370 1850
rect 16832 1816 17388 1850
rect 17850 1816 18406 1850
rect 18868 1816 19424 1850
rect 19886 1816 20442 1850
rect 20904 1816 21460 1850
rect 21922 1816 22478 1850
rect 22940 1816 23496 1850
rect 23958 1816 24514 1850
rect 24976 1816 25532 1850
rect 25994 1816 26550 1850
rect 27012 1816 27568 1850
rect 28030 1816 28586 1850
rect 29048 1816 29604 1850
rect 30066 1816 30622 1850
rect 31084 1816 31640 1850
rect 32102 1816 32658 1850
rect 33120 1816 33676 1850
rect 1792 1460 2348 1494
rect 2810 1460 3366 1494
rect 3828 1460 4384 1494
rect 4846 1460 5402 1494
rect 5864 1460 6420 1494
rect 6882 1460 7438 1494
rect 8642 1464 8766 1498
rect 8940 1464 9064 1498
rect 9238 1464 9362 1498
rect 9536 1464 9660 1498
rect 9834 1464 9958 1498
rect 10132 1464 10256 1498
rect 10430 1464 10554 1498
rect 10728 1464 10852 1498
rect 11026 1464 11150 1498
rect 11324 1464 11448 1498
rect 11622 1464 11746 1498
rect 13778 1294 14334 1328
rect 14796 1294 15352 1328
rect 15814 1294 16370 1328
rect 16832 1294 17388 1328
rect 17850 1294 18406 1328
rect 18868 1294 19424 1328
rect 19886 1294 20442 1328
rect 20904 1294 21460 1328
rect 21922 1294 22478 1328
rect 22940 1294 23496 1328
rect 23958 1294 24514 1328
rect 24976 1294 25532 1328
rect 25994 1294 26550 1328
rect 27012 1294 27568 1328
rect 28030 1294 28586 1328
rect 29048 1294 29604 1328
rect 30066 1294 30622 1328
rect 31084 1294 31640 1328
rect 32102 1294 32658 1328
rect 33120 1294 33676 1328
rect 1792 750 2348 784
rect 2810 750 3366 784
rect 3828 750 4384 784
rect 4846 750 5402 784
rect 5864 750 6420 784
rect 6882 750 7438 784
rect 8642 754 8766 788
rect 8940 754 9064 788
rect 9238 754 9362 788
rect 9536 754 9660 788
rect 9834 754 9958 788
rect 10132 754 10256 788
rect 10430 754 10554 788
rect 10728 754 10852 788
rect 11026 754 11150 788
rect 11324 754 11448 788
rect 11622 754 11746 788
rect 13778 584 14334 618
rect 14796 584 15352 618
rect 15814 584 16370 618
rect 16832 584 17388 618
rect 17850 584 18406 618
rect 18868 584 19424 618
rect 19886 584 20442 618
rect 20904 584 21460 618
rect 21922 584 22478 618
rect 22940 584 23496 618
rect 23958 584 24514 618
rect 24976 584 25532 618
rect 25994 584 26550 618
rect 27012 584 27568 618
rect 28030 584 28586 618
rect 29048 584 29604 618
rect 30066 584 30622 618
rect 31084 584 31640 618
rect 32102 584 32658 618
rect 33120 584 33676 618
rect 48900 8311 49000 8345
rect 49158 8311 49258 8345
rect 49416 8311 49516 8345
rect 49674 8311 49774 8345
rect 49932 8311 50032 8345
rect 50190 8311 50290 8345
rect 48900 7783 49000 7817
rect 49158 7783 49258 7817
rect 49416 7783 49516 7817
rect 49674 7783 49774 7817
rect 49932 7783 50032 7817
rect 50190 7783 50290 7817
rect 50736 7599 50770 7633
rect 48900 7378 49000 7412
rect 49158 7378 49258 7412
rect 49416 7378 49516 7412
rect 49674 7378 49774 7412
rect 49932 7378 50032 7412
rect 50190 7378 50290 7412
rect 48900 7068 49000 7102
rect 49158 7068 49258 7102
rect 49416 7068 49516 7102
rect 49674 7068 49774 7102
rect 49932 7068 50032 7102
rect 50190 7068 50290 7102
rect 48900 6347 49000 6381
rect 49158 6347 49258 6381
rect 49416 6347 49516 6381
rect 49674 6347 49774 6381
rect 49932 6347 50032 6381
rect 50190 6347 50290 6381
rect 48900 5819 49000 5853
rect 49158 5819 49258 5853
rect 49416 5819 49516 5853
rect 49674 5819 49774 5853
rect 49932 5819 50032 5853
rect 50190 5819 50290 5853
rect 50736 5635 50770 5669
rect 48900 5414 49000 5448
rect 49158 5414 49258 5448
rect 49416 5414 49516 5448
rect 49674 5414 49774 5448
rect 49932 5414 50032 5448
rect 50190 5414 50290 5448
rect 48900 5104 49000 5138
rect 49158 5104 49258 5138
rect 49416 5104 49516 5138
rect 49674 5104 49774 5138
rect 49932 5104 50032 5138
rect 50190 5104 50290 5138
rect 48900 4347 49000 4381
rect 49158 4347 49258 4381
rect 49416 4347 49516 4381
rect 49674 4347 49774 4381
rect 49932 4347 50032 4381
rect 50190 4347 50290 4381
rect 48900 3819 49000 3853
rect 49158 3819 49258 3853
rect 49416 3819 49516 3853
rect 49674 3819 49774 3853
rect 49932 3819 50032 3853
rect 50190 3819 50290 3853
rect 50736 3635 50770 3669
rect 48900 3414 49000 3448
rect 49158 3414 49258 3448
rect 49416 3414 49516 3448
rect 49674 3414 49774 3448
rect 49932 3414 50032 3448
rect 50190 3414 50290 3448
rect 48900 3104 49000 3138
rect 49158 3104 49258 3138
rect 49416 3104 49516 3138
rect 49674 3104 49774 3138
rect 49932 3104 50032 3138
rect 50190 3104 50290 3138
rect 48900 2257 49000 2291
rect 49158 2257 49258 2291
rect 49416 2257 49516 2291
rect 49674 2257 49774 2291
rect 49932 2257 50032 2291
rect 50190 2257 50290 2291
rect 48900 1729 49000 1763
rect 49158 1729 49258 1763
rect 49416 1729 49516 1763
rect 49674 1729 49774 1763
rect 49932 1729 50032 1763
rect 50190 1729 50290 1763
rect 50736 1545 50770 1579
rect 48900 1324 49000 1358
rect 49158 1324 49258 1358
rect 49416 1324 49516 1358
rect 49674 1324 49774 1358
rect 49932 1324 50032 1358
rect 50190 1324 50290 1358
rect 48900 1014 49000 1048
rect 49158 1014 49258 1048
rect 49416 1014 49516 1048
rect 49674 1014 49774 1048
rect 49932 1014 50032 1048
rect 50190 1014 50290 1048
rect 67780 14860 68336 14894
rect 68798 14860 69354 14894
rect 69816 14860 70372 14894
rect 70834 14860 71390 14894
rect 71852 14860 72408 14894
rect 72870 14860 73426 14894
rect 73888 14860 74444 14894
rect 74906 14860 75462 14894
rect 75924 14860 76480 14894
rect 76942 14860 77498 14894
rect 77960 14860 78516 14894
rect 78978 14860 79534 14894
rect 79996 14860 80552 14894
rect 81014 14860 81570 14894
rect 82032 14860 82588 14894
rect 83050 14860 83606 14894
rect 84068 14860 84624 14894
rect 85086 14860 85642 14894
rect 86104 14860 86660 14894
rect 87122 14860 87678 14894
rect 67780 14150 68336 14184
rect 68798 14150 69354 14184
rect 69816 14150 70372 14184
rect 70834 14150 71390 14184
rect 71852 14150 72408 14184
rect 72870 14150 73426 14184
rect 73888 14150 74444 14184
rect 74906 14150 75462 14184
rect 75924 14150 76480 14184
rect 76942 14150 77498 14184
rect 77960 14150 78516 14184
rect 78978 14150 79534 14184
rect 79996 14150 80552 14184
rect 81014 14150 81570 14184
rect 82032 14150 82588 14184
rect 83050 14150 83606 14184
rect 84068 14150 84624 14184
rect 85086 14150 85642 14184
rect 86104 14150 86660 14184
rect 87122 14150 87678 14184
rect 56014 14066 56570 14100
rect 57032 14066 57588 14100
rect 58050 14066 58606 14100
rect 59068 14066 59624 14100
rect 60086 14066 60642 14100
rect 61104 14066 61660 14100
rect 62122 14066 62678 14100
rect 63140 14066 63696 14100
rect 64158 14066 64714 14100
rect 67780 13626 68336 13660
rect 68798 13626 69354 13660
rect 69816 13626 70372 13660
rect 70834 13626 71390 13660
rect 71852 13626 72408 13660
rect 72870 13626 73426 13660
rect 73888 13626 74444 13660
rect 74906 13626 75462 13660
rect 75924 13626 76480 13660
rect 76942 13626 77498 13660
rect 77960 13626 78516 13660
rect 78978 13626 79534 13660
rect 79996 13626 80552 13660
rect 81014 13626 81570 13660
rect 82032 13626 82588 13660
rect 83050 13626 83606 13660
rect 84068 13626 84624 13660
rect 85086 13626 85642 13660
rect 86104 13626 86660 13660
rect 87122 13626 87678 13660
rect 56014 13356 56570 13390
rect 57032 13356 57588 13390
rect 56014 13248 56570 13282
rect 58050 13356 58606 13390
rect 57032 13248 57588 13282
rect 59068 13356 59624 13390
rect 58050 13248 58606 13282
rect 60086 13356 60642 13390
rect 59068 13248 59624 13282
rect 61104 13356 61660 13390
rect 60086 13248 60642 13282
rect 62122 13356 62678 13390
rect 61104 13248 61660 13282
rect 63140 13356 63696 13390
rect 62122 13248 62678 13282
rect 64158 13356 64714 13390
rect 63140 13248 63696 13282
rect 64158 13248 64714 13282
rect 67780 12916 68336 12950
rect 68798 12916 69354 12950
rect 69816 12916 70372 12950
rect 70834 12916 71390 12950
rect 71852 12916 72408 12950
rect 72870 12916 73426 12950
rect 73888 12916 74444 12950
rect 74906 12916 75462 12950
rect 75924 12916 76480 12950
rect 76942 12916 77498 12950
rect 77960 12916 78516 12950
rect 78978 12916 79534 12950
rect 79996 12916 80552 12950
rect 81014 12916 81570 12950
rect 82032 12916 82588 12950
rect 83050 12916 83606 12950
rect 84068 12916 84624 12950
rect 85086 12916 85642 12950
rect 86104 12916 86660 12950
rect 87122 12916 87678 12950
rect 56014 12538 56570 12572
rect 57032 12538 57588 12572
rect 56014 12430 56570 12464
rect 58050 12538 58606 12572
rect 57032 12430 57588 12464
rect 59068 12538 59624 12572
rect 58050 12430 58606 12464
rect 60086 12538 60642 12572
rect 59068 12430 59624 12464
rect 61104 12538 61660 12572
rect 60086 12430 60642 12464
rect 62122 12538 62678 12572
rect 61104 12430 61660 12464
rect 63140 12538 63696 12572
rect 62122 12430 62678 12464
rect 64158 12538 64714 12572
rect 63140 12430 63696 12464
rect 64158 12430 64714 12464
rect 67780 12394 68336 12428
rect 68798 12394 69354 12428
rect 69816 12394 70372 12428
rect 70834 12394 71390 12428
rect 71852 12394 72408 12428
rect 72870 12394 73426 12428
rect 73888 12394 74444 12428
rect 74906 12394 75462 12428
rect 75924 12394 76480 12428
rect 76942 12394 77498 12428
rect 77960 12394 78516 12428
rect 78978 12394 79534 12428
rect 79996 12394 80552 12428
rect 81014 12394 81570 12428
rect 82032 12394 82588 12428
rect 83050 12394 83606 12428
rect 84068 12394 84624 12428
rect 85086 12394 85642 12428
rect 86104 12394 86660 12428
rect 87122 12394 87678 12428
rect 56014 11720 56570 11754
rect 57032 11720 57588 11754
rect 56014 11612 56570 11646
rect 58050 11720 58606 11754
rect 57032 11612 57588 11646
rect 59068 11720 59624 11754
rect 58050 11612 58606 11646
rect 60086 11720 60642 11754
rect 59068 11612 59624 11646
rect 61104 11720 61660 11754
rect 60086 11612 60642 11646
rect 62122 11720 62678 11754
rect 61104 11612 61660 11646
rect 63140 11720 63696 11754
rect 62122 11612 62678 11646
rect 64158 11720 64714 11754
rect 63140 11612 63696 11646
rect 67780 11684 68336 11718
rect 68798 11684 69354 11718
rect 69816 11684 70372 11718
rect 70834 11684 71390 11718
rect 71852 11684 72408 11718
rect 72870 11684 73426 11718
rect 73888 11684 74444 11718
rect 74906 11684 75462 11718
rect 75924 11684 76480 11718
rect 76942 11684 77498 11718
rect 77960 11684 78516 11718
rect 78978 11684 79534 11718
rect 79996 11684 80552 11718
rect 81014 11684 81570 11718
rect 82032 11684 82588 11718
rect 83050 11684 83606 11718
rect 84068 11684 84624 11718
rect 85086 11684 85642 11718
rect 86104 11684 86660 11718
rect 87122 11684 87678 11718
rect 64158 11612 64714 11646
rect 67778 11160 68334 11194
rect 68796 11160 69352 11194
rect 69814 11160 70370 11194
rect 70832 11160 71388 11194
rect 71850 11160 72406 11194
rect 72868 11160 73424 11194
rect 73886 11160 74442 11194
rect 74904 11160 75460 11194
rect 75922 11160 76478 11194
rect 76940 11160 77496 11194
rect 77958 11160 78514 11194
rect 78976 11160 79532 11194
rect 79994 11160 80550 11194
rect 81012 11160 81568 11194
rect 82030 11160 82586 11194
rect 83048 11160 83604 11194
rect 84066 11160 84622 11194
rect 85084 11160 85640 11194
rect 86102 11160 86658 11194
rect 87120 11160 87676 11194
rect 56014 10902 56570 10936
rect 57032 10902 57588 10936
rect 56014 10794 56570 10828
rect 58050 10902 58606 10936
rect 57032 10794 57588 10828
rect 59068 10902 59624 10936
rect 58050 10794 58606 10828
rect 60086 10902 60642 10936
rect 59068 10794 59624 10828
rect 61104 10902 61660 10936
rect 60086 10794 60642 10828
rect 62122 10902 62678 10936
rect 61104 10794 61660 10828
rect 63140 10902 63696 10936
rect 62122 10794 62678 10828
rect 64158 10902 64714 10936
rect 63140 10794 63696 10828
rect 64158 10794 64714 10828
rect 67778 10450 68334 10484
rect 68796 10450 69352 10484
rect 69814 10450 70370 10484
rect 70832 10450 71388 10484
rect 71850 10450 72406 10484
rect 72868 10450 73424 10484
rect 73886 10450 74442 10484
rect 74904 10450 75460 10484
rect 75922 10450 76478 10484
rect 76940 10450 77496 10484
rect 77958 10450 78514 10484
rect 78976 10450 79532 10484
rect 79994 10450 80550 10484
rect 81012 10450 81568 10484
rect 82030 10450 82586 10484
rect 83048 10450 83604 10484
rect 84066 10450 84622 10484
rect 85084 10450 85640 10484
rect 86102 10450 86658 10484
rect 87120 10450 87676 10484
rect 56014 10084 56570 10118
rect 57032 10084 57588 10118
rect 56014 9976 56570 10010
rect 58050 10084 58606 10118
rect 57032 9976 57588 10010
rect 59068 10084 59624 10118
rect 58050 9976 58606 10010
rect 60086 10084 60642 10118
rect 59068 9976 59624 10010
rect 61104 10084 61660 10118
rect 60086 9976 60642 10010
rect 62122 10084 62678 10118
rect 61104 9976 61660 10010
rect 63140 10084 63696 10118
rect 62122 9976 62678 10010
rect 64158 10084 64714 10118
rect 63140 9976 63696 10010
rect 64158 9976 64714 10010
rect 67778 9926 68334 9960
rect 68796 9926 69352 9960
rect 69814 9926 70370 9960
rect 70832 9926 71388 9960
rect 71850 9926 72406 9960
rect 72868 9926 73424 9960
rect 73886 9926 74442 9960
rect 74904 9926 75460 9960
rect 75922 9926 76478 9960
rect 76940 9926 77496 9960
rect 77958 9926 78514 9960
rect 78976 9926 79532 9960
rect 79994 9926 80550 9960
rect 81012 9926 81568 9960
rect 82030 9926 82586 9960
rect 83048 9926 83604 9960
rect 84066 9926 84622 9960
rect 85084 9926 85640 9960
rect 86102 9926 86658 9960
rect 87120 9926 87676 9960
rect 56014 9266 56570 9300
rect 57032 9266 57588 9300
rect 56014 9158 56570 9192
rect 58050 9266 58606 9300
rect 57032 9158 57588 9192
rect 59068 9266 59624 9300
rect 58050 9158 58606 9192
rect 60086 9266 60642 9300
rect 59068 9158 59624 9192
rect 61104 9266 61660 9300
rect 60086 9158 60642 9192
rect 62122 9266 62678 9300
rect 61104 9158 61660 9192
rect 63140 9266 63696 9300
rect 62122 9158 62678 9192
rect 64158 9266 64714 9300
rect 63140 9158 63696 9192
rect 64158 9158 64714 9192
rect 67778 9216 68334 9250
rect 68796 9216 69352 9250
rect 69814 9216 70370 9250
rect 70832 9216 71388 9250
rect 71850 9216 72406 9250
rect 72868 9216 73424 9250
rect 73886 9216 74442 9250
rect 74904 9216 75460 9250
rect 75922 9216 76478 9250
rect 76940 9216 77496 9250
rect 77958 9216 78514 9250
rect 78976 9216 79532 9250
rect 79994 9216 80550 9250
rect 81012 9216 81568 9250
rect 82030 9216 82586 9250
rect 83048 9216 83604 9250
rect 84066 9216 84622 9250
rect 85084 9216 85640 9250
rect 86102 9216 86658 9250
rect 87120 9216 87676 9250
rect 67778 8694 68334 8728
rect 68796 8694 69352 8728
rect 69814 8694 70370 8728
rect 70832 8694 71388 8728
rect 71850 8694 72406 8728
rect 72868 8694 73424 8728
rect 73886 8694 74442 8728
rect 74904 8694 75460 8728
rect 75922 8694 76478 8728
rect 76940 8694 77496 8728
rect 77958 8694 78514 8728
rect 78976 8694 79532 8728
rect 79994 8694 80550 8728
rect 81012 8694 81568 8728
rect 82030 8694 82586 8728
rect 83048 8694 83604 8728
rect 84066 8694 84622 8728
rect 85084 8694 85640 8728
rect 86102 8694 86658 8728
rect 87120 8694 87676 8728
rect 56014 8448 56570 8482
rect 57032 8448 57588 8482
rect 56014 8340 56570 8374
rect 58050 8448 58606 8482
rect 57032 8340 57588 8374
rect 59068 8448 59624 8482
rect 58050 8340 58606 8374
rect 60086 8448 60642 8482
rect 59068 8340 59624 8374
rect 61104 8448 61660 8482
rect 60086 8340 60642 8374
rect 62122 8448 62678 8482
rect 61104 8340 61660 8374
rect 63140 8448 63696 8482
rect 62122 8340 62678 8374
rect 64158 8448 64714 8482
rect 63140 8340 63696 8374
rect 64158 8340 64714 8374
rect 67778 7984 68334 8018
rect 68796 7984 69352 8018
rect 69814 7984 70370 8018
rect 70832 7984 71388 8018
rect 71850 7984 72406 8018
rect 72868 7984 73424 8018
rect 73886 7984 74442 8018
rect 74904 7984 75460 8018
rect 75922 7984 76478 8018
rect 76940 7984 77496 8018
rect 77958 7984 78514 8018
rect 78976 7984 79532 8018
rect 79994 7984 80550 8018
rect 81012 7984 81568 8018
rect 82030 7984 82586 8018
rect 83048 7984 83604 8018
rect 84066 7984 84622 8018
rect 85084 7984 85640 8018
rect 86102 7984 86658 8018
rect 87120 7984 87676 8018
rect 56014 7630 56570 7664
rect 57032 7630 57588 7664
rect 58050 7630 58606 7664
rect 59068 7630 59624 7664
rect 60086 7630 60642 7664
rect 61104 7630 61660 7664
rect 62122 7630 62678 7664
rect 63140 7630 63696 7664
rect 64158 7630 64714 7664
rect 67778 7460 68334 7494
rect 68796 7460 69352 7494
rect 69814 7460 70370 7494
rect 70832 7460 71388 7494
rect 71850 7460 72406 7494
rect 72868 7460 73424 7494
rect 73886 7460 74442 7494
rect 74904 7460 75460 7494
rect 75922 7460 76478 7494
rect 76940 7460 77496 7494
rect 77958 7460 78514 7494
rect 78976 7460 79532 7494
rect 79994 7460 80550 7494
rect 81012 7460 81568 7494
rect 82030 7460 82586 7494
rect 83048 7460 83604 7494
rect 84066 7460 84622 7494
rect 85084 7460 85640 7494
rect 86102 7460 86658 7494
rect 87120 7460 87676 7494
rect 62714 6956 62790 6990
rect 62932 6956 63008 6990
rect 63150 6956 63226 6990
rect 63368 6956 63444 6990
rect 63586 6956 63662 6990
rect 63804 6956 63880 6990
rect 64022 6956 64098 6990
rect 64240 6956 64316 6990
rect 64458 6956 64534 6990
rect 64676 6956 64752 6990
rect 67778 6750 68334 6784
rect 68796 6750 69352 6784
rect 69814 6750 70370 6784
rect 70832 6750 71388 6784
rect 71850 6750 72406 6784
rect 72868 6750 73424 6784
rect 73886 6750 74442 6784
rect 74904 6750 75460 6784
rect 75922 6750 76478 6784
rect 76940 6750 77496 6784
rect 77958 6750 78514 6784
rect 78976 6750 79532 6784
rect 79994 6750 80550 6784
rect 81012 6750 81568 6784
rect 82030 6750 82586 6784
rect 83048 6750 83604 6784
rect 84066 6750 84622 6784
rect 85084 6750 85640 6784
rect 86102 6750 86658 6784
rect 87120 6750 87676 6784
rect 62714 6646 62790 6680
rect 62932 6646 63008 6680
rect 63150 6646 63226 6680
rect 63368 6646 63444 6680
rect 63586 6646 63662 6680
rect 63804 6646 63880 6680
rect 64022 6646 64098 6680
rect 64240 6646 64316 6680
rect 64458 6646 64534 6680
rect 64676 6646 64752 6680
rect 67778 6226 68334 6260
rect 68796 6226 69352 6260
rect 69814 6226 70370 6260
rect 70832 6226 71388 6260
rect 71850 6226 72406 6260
rect 72868 6226 73424 6260
rect 73886 6226 74442 6260
rect 74904 6226 75460 6260
rect 75922 6226 76478 6260
rect 76940 6226 77496 6260
rect 77958 6226 78514 6260
rect 78976 6226 79532 6260
rect 79994 6226 80550 6260
rect 81012 6226 81568 6260
rect 82030 6226 82586 6260
rect 83048 6226 83604 6260
rect 84066 6226 84622 6260
rect 85084 6226 85640 6260
rect 86102 6226 86658 6260
rect 87120 6226 87676 6260
rect 62714 6124 62790 6158
rect 62932 6124 63008 6158
rect 63150 6124 63226 6158
rect 63368 6124 63444 6158
rect 63586 6124 63662 6158
rect 63804 6124 63880 6158
rect 64022 6124 64098 6158
rect 64240 6124 64316 6158
rect 64458 6124 64534 6158
rect 64676 6124 64752 6158
rect 62714 5814 62790 5848
rect 62932 5814 63008 5848
rect 63150 5814 63226 5848
rect 63368 5814 63444 5848
rect 63586 5814 63662 5848
rect 63804 5814 63880 5848
rect 64022 5814 64098 5848
rect 64240 5814 64316 5848
rect 64458 5814 64534 5848
rect 64676 5814 64752 5848
rect 67778 5516 68334 5550
rect 68796 5516 69352 5550
rect 69814 5516 70370 5550
rect 70832 5516 71388 5550
rect 71850 5516 72406 5550
rect 72868 5516 73424 5550
rect 73886 5516 74442 5550
rect 74904 5516 75460 5550
rect 75922 5516 76478 5550
rect 76940 5516 77496 5550
rect 77958 5516 78514 5550
rect 78976 5516 79532 5550
rect 79994 5516 80550 5550
rect 81012 5516 81568 5550
rect 82030 5516 82586 5550
rect 83048 5516 83604 5550
rect 84066 5516 84622 5550
rect 85084 5516 85640 5550
rect 86102 5516 86658 5550
rect 87120 5516 87676 5550
rect 67778 4994 68334 5028
rect 68796 4994 69352 5028
rect 69814 4994 70370 5028
rect 70832 4994 71388 5028
rect 71850 4994 72406 5028
rect 72868 4994 73424 5028
rect 73886 4994 74442 5028
rect 74904 4994 75460 5028
rect 75922 4994 76478 5028
rect 76940 4994 77496 5028
rect 77958 4994 78514 5028
rect 78976 4994 79532 5028
rect 79994 4994 80550 5028
rect 81012 4994 81568 5028
rect 82030 4994 82586 5028
rect 83048 4994 83604 5028
rect 84066 4994 84622 5028
rect 85084 4994 85640 5028
rect 86102 4994 86658 5028
rect 87120 4994 87676 5028
rect 55793 4797 56349 4831
rect 56811 4797 57367 4831
rect 57829 4797 58385 4831
rect 58847 4797 59403 4831
rect 59865 4797 60421 4831
rect 60883 4797 61439 4831
rect 62644 4798 62768 4832
rect 62942 4798 63066 4832
rect 63240 4798 63364 4832
rect 63538 4798 63662 4832
rect 63836 4798 63960 4832
rect 64134 4798 64258 4832
rect 64432 4798 64556 4832
rect 64730 4798 64854 4832
rect 65028 4798 65152 4832
rect 65326 4798 65450 4832
rect 65624 4798 65748 4832
rect 67778 4284 68334 4318
rect 68796 4284 69352 4318
rect 69814 4284 70370 4318
rect 70832 4284 71388 4318
rect 71850 4284 72406 4318
rect 72868 4284 73424 4318
rect 73886 4284 74442 4318
rect 74904 4284 75460 4318
rect 75922 4284 76478 4318
rect 76940 4284 77496 4318
rect 77958 4284 78514 4318
rect 78976 4284 79532 4318
rect 79994 4284 80550 4318
rect 81012 4284 81568 4318
rect 82030 4284 82586 4318
rect 83048 4284 83604 4318
rect 84066 4284 84622 4318
rect 85084 4284 85640 4318
rect 86102 4284 86658 4318
rect 87120 4284 87676 4318
rect 55793 4087 56349 4121
rect 56811 4087 57367 4121
rect 57829 4087 58385 4121
rect 58847 4087 59403 4121
rect 59865 4087 60421 4121
rect 60883 4087 61439 4121
rect 62644 4088 62768 4122
rect 62942 4088 63066 4122
rect 63240 4088 63364 4122
rect 63538 4088 63662 4122
rect 63836 4088 63960 4122
rect 64134 4088 64258 4122
rect 64432 4088 64556 4122
rect 64730 4088 64854 4122
rect 65028 4088 65152 4122
rect 65326 4088 65450 4122
rect 65624 4088 65748 4122
rect 67778 3760 68334 3794
rect 55792 3684 56348 3718
rect 56810 3684 57366 3718
rect 57828 3684 58384 3718
rect 58846 3684 59402 3718
rect 59864 3684 60420 3718
rect 60882 3684 61438 3718
rect 62644 3686 62768 3720
rect 62942 3686 63066 3720
rect 63240 3686 63364 3720
rect 63538 3686 63662 3720
rect 63836 3686 63960 3720
rect 64134 3686 64258 3720
rect 64432 3686 64556 3720
rect 64730 3686 64854 3720
rect 65028 3686 65152 3720
rect 65326 3686 65450 3720
rect 68796 3760 69352 3794
rect 69814 3760 70370 3794
rect 70832 3760 71388 3794
rect 71850 3760 72406 3794
rect 72868 3760 73424 3794
rect 73886 3760 74442 3794
rect 74904 3760 75460 3794
rect 75922 3760 76478 3794
rect 76940 3760 77496 3794
rect 77958 3760 78514 3794
rect 78976 3760 79532 3794
rect 79994 3760 80550 3794
rect 81012 3760 81568 3794
rect 82030 3760 82586 3794
rect 83048 3760 83604 3794
rect 84066 3760 84622 3794
rect 85084 3760 85640 3794
rect 86102 3760 86658 3794
rect 87120 3760 87676 3794
rect 65624 3686 65748 3720
rect 67778 3050 68334 3084
rect 55792 2974 56348 3008
rect 56810 2974 57366 3008
rect 57828 2974 58384 3008
rect 58846 2974 59402 3008
rect 59864 2974 60420 3008
rect 60882 2974 61438 3008
rect 62644 2976 62768 3010
rect 62942 2976 63066 3010
rect 63240 2976 63364 3010
rect 63538 2976 63662 3010
rect 63836 2976 63960 3010
rect 64134 2976 64258 3010
rect 64432 2976 64556 3010
rect 64730 2976 64854 3010
rect 65028 2976 65152 3010
rect 65326 2976 65450 3010
rect 68796 3050 69352 3084
rect 69814 3050 70370 3084
rect 70832 3050 71388 3084
rect 71850 3050 72406 3084
rect 72868 3050 73424 3084
rect 73886 3050 74442 3084
rect 74904 3050 75460 3084
rect 75922 3050 76478 3084
rect 76940 3050 77496 3084
rect 77958 3050 78514 3084
rect 78976 3050 79532 3084
rect 79994 3050 80550 3084
rect 81012 3050 81568 3084
rect 82030 3050 82586 3084
rect 83048 3050 83604 3084
rect 84066 3050 84622 3084
rect 85084 3050 85640 3084
rect 86102 3050 86658 3084
rect 87120 3050 87676 3084
rect 65624 2976 65748 3010
rect 55793 2573 56349 2607
rect 56811 2573 57367 2607
rect 57829 2573 58385 2607
rect 58847 2573 59403 2607
rect 59865 2573 60421 2607
rect 60883 2573 61439 2607
rect 62642 2574 62766 2608
rect 62940 2574 63064 2608
rect 63238 2574 63362 2608
rect 63536 2574 63660 2608
rect 63834 2574 63958 2608
rect 64132 2574 64256 2608
rect 64430 2574 64554 2608
rect 64728 2574 64852 2608
rect 65026 2574 65150 2608
rect 65324 2574 65448 2608
rect 65622 2574 65746 2608
rect 67778 2526 68334 2560
rect 68796 2526 69352 2560
rect 69814 2526 70370 2560
rect 70832 2526 71388 2560
rect 71850 2526 72406 2560
rect 72868 2526 73424 2560
rect 73886 2526 74442 2560
rect 74904 2526 75460 2560
rect 75922 2526 76478 2560
rect 76940 2526 77496 2560
rect 77958 2526 78514 2560
rect 78976 2526 79532 2560
rect 79994 2526 80550 2560
rect 81012 2526 81568 2560
rect 82030 2526 82586 2560
rect 83048 2526 83604 2560
rect 84066 2526 84622 2560
rect 85084 2526 85640 2560
rect 86102 2526 86658 2560
rect 87120 2526 87676 2560
rect 55793 1863 56349 1897
rect 56811 1863 57367 1897
rect 57829 1863 58385 1897
rect 58847 1863 59403 1897
rect 59865 1863 60421 1897
rect 60883 1863 61439 1897
rect 62642 1864 62766 1898
rect 62940 1864 63064 1898
rect 63238 1864 63362 1898
rect 63536 1864 63660 1898
rect 63834 1864 63958 1898
rect 64132 1864 64256 1898
rect 64430 1864 64554 1898
rect 64728 1864 64852 1898
rect 65026 1864 65150 1898
rect 65324 1864 65448 1898
rect 65622 1864 65746 1898
rect 67778 1816 68334 1850
rect 68796 1816 69352 1850
rect 69814 1816 70370 1850
rect 70832 1816 71388 1850
rect 71850 1816 72406 1850
rect 72868 1816 73424 1850
rect 73886 1816 74442 1850
rect 74904 1816 75460 1850
rect 75922 1816 76478 1850
rect 76940 1816 77496 1850
rect 77958 1816 78514 1850
rect 78976 1816 79532 1850
rect 79994 1816 80550 1850
rect 81012 1816 81568 1850
rect 82030 1816 82586 1850
rect 83048 1816 83604 1850
rect 84066 1816 84622 1850
rect 85084 1816 85640 1850
rect 86102 1816 86658 1850
rect 87120 1816 87676 1850
rect 55792 1460 56348 1494
rect 56810 1460 57366 1494
rect 57828 1460 58384 1494
rect 58846 1460 59402 1494
rect 59864 1460 60420 1494
rect 60882 1460 61438 1494
rect 62642 1464 62766 1498
rect 62940 1464 63064 1498
rect 63238 1464 63362 1498
rect 63536 1464 63660 1498
rect 63834 1464 63958 1498
rect 64132 1464 64256 1498
rect 64430 1464 64554 1498
rect 64728 1464 64852 1498
rect 65026 1464 65150 1498
rect 65324 1464 65448 1498
rect 65622 1464 65746 1498
rect 67778 1294 68334 1328
rect 68796 1294 69352 1328
rect 69814 1294 70370 1328
rect 70832 1294 71388 1328
rect 71850 1294 72406 1328
rect 72868 1294 73424 1328
rect 73886 1294 74442 1328
rect 74904 1294 75460 1328
rect 75922 1294 76478 1328
rect 76940 1294 77496 1328
rect 77958 1294 78514 1328
rect 78976 1294 79532 1328
rect 79994 1294 80550 1328
rect 81012 1294 81568 1328
rect 82030 1294 82586 1328
rect 83048 1294 83604 1328
rect 84066 1294 84622 1328
rect 85084 1294 85640 1328
rect 86102 1294 86658 1328
rect 87120 1294 87676 1328
rect 55792 750 56348 784
rect 56810 750 57366 784
rect 57828 750 58384 784
rect 58846 750 59402 784
rect 59864 750 60420 784
rect 60882 750 61438 784
rect 62642 754 62766 788
rect 62940 754 63064 788
rect 63238 754 63362 788
rect 63536 754 63660 788
rect 63834 754 63958 788
rect 64132 754 64256 788
rect 64430 754 64554 788
rect 64728 754 64852 788
rect 65026 754 65150 788
rect 65324 754 65448 788
rect 65622 754 65746 788
rect 67778 584 68334 618
rect 68796 584 69352 618
rect 69814 584 70370 618
rect 70832 584 71388 618
rect 71850 584 72406 618
rect 72868 584 73424 618
rect 73886 584 74442 618
rect 74904 584 75460 618
rect 75922 584 76478 618
rect 76940 584 77496 618
rect 77958 584 78514 618
rect 78976 584 79532 618
rect 79994 584 80550 618
rect 81012 584 81568 618
rect 82030 584 82586 618
rect 83048 584 83604 618
rect 84066 584 84622 618
rect 85084 584 85640 618
rect 86102 584 86658 618
rect 87120 584 87676 618
<< locali >>
rect 11328 28100 11428 28262
rect 35672 28100 35772 28262
rect 17670 27027 17686 27061
rect 18242 27027 18258 27061
rect 18688 27027 18704 27061
rect 19260 27027 19276 27061
rect 19706 27027 19722 27061
rect 20278 27027 20294 27061
rect 20724 27027 20740 27061
rect 21296 27027 21312 27061
rect 21742 27027 21758 27061
rect 22314 27027 22330 27061
rect 22760 27027 22776 27061
rect 23332 27027 23348 27061
rect 23778 27027 23794 27061
rect 24350 27027 24366 27061
rect 24796 27027 24812 27061
rect 25368 27027 25384 27061
rect 25814 27027 25830 27061
rect 26386 27027 26402 27061
rect 26832 27027 26848 27061
rect 27404 27027 27420 27061
rect 27850 27027 27866 27061
rect 28422 27027 28438 27061
rect 28868 27027 28884 27061
rect 29440 27027 29456 27061
rect 29886 27027 29902 27061
rect 30458 27027 30474 27061
rect 30904 27027 30920 27061
rect 31476 27027 31492 27061
rect 31922 27027 31938 27061
rect 32494 27027 32510 27061
rect 32940 27027 32956 27061
rect 33512 27027 33528 27061
rect 17438 26968 17472 26984
rect 17438 26376 17472 26392
rect 18456 26968 18490 26984
rect 18456 26376 18490 26392
rect 19474 26968 19508 26984
rect 19474 26376 19508 26392
rect 20492 26968 20526 26984
rect 20492 26376 20526 26392
rect 21510 26968 21544 26984
rect 21510 26376 21544 26392
rect 22528 26968 22562 26984
rect 22528 26376 22562 26392
rect 23546 26968 23580 26984
rect 23546 26376 23580 26392
rect 24564 26968 24598 26984
rect 24564 26376 24598 26392
rect 25582 26968 25616 26984
rect 25582 26376 25616 26392
rect 26600 26968 26634 26984
rect 26600 26376 26634 26392
rect 27618 26968 27652 26984
rect 27618 26376 27652 26392
rect 28636 26968 28670 26984
rect 28636 26376 28670 26392
rect 29654 26968 29688 26984
rect 29654 26376 29688 26392
rect 30672 26968 30706 26984
rect 30672 26376 30706 26392
rect 31690 26968 31724 26984
rect 31690 26376 31724 26392
rect 32708 26968 32742 26984
rect 32708 26376 32742 26392
rect 33726 26968 33760 26984
rect 33726 26376 33760 26392
rect 17670 26299 17686 26333
rect 18242 26299 18258 26333
rect 18688 26299 18704 26333
rect 19260 26299 19276 26333
rect 19706 26299 19722 26333
rect 20278 26299 20294 26333
rect 20724 26299 20740 26333
rect 21296 26299 21312 26333
rect 21742 26299 21758 26333
rect 22314 26299 22330 26333
rect 22760 26299 22776 26333
rect 23332 26299 23348 26333
rect 23778 26299 23794 26333
rect 24350 26299 24366 26333
rect 24796 26299 24812 26333
rect 25368 26299 25384 26333
rect 25814 26299 25830 26333
rect 26386 26299 26402 26333
rect 26832 26299 26848 26333
rect 27404 26299 27420 26333
rect 27850 26299 27866 26333
rect 28422 26299 28438 26333
rect 28868 26299 28884 26333
rect 29440 26299 29456 26333
rect 29886 26299 29902 26333
rect 30458 26299 30474 26333
rect 30904 26299 30920 26333
rect 31476 26299 31492 26333
rect 31922 26299 31938 26333
rect 32494 26299 32510 26333
rect 32940 26299 32956 26333
rect 33512 26299 33528 26333
rect 18936 26142 19026 26172
rect 18936 26108 18964 26142
rect 18998 26108 19026 26142
rect 18936 26080 19026 26108
rect 19954 26142 20044 26172
rect 19954 26108 19982 26142
rect 20016 26108 20044 26142
rect 19954 26080 20044 26108
rect 20972 26142 21062 26172
rect 20972 26108 21000 26142
rect 21034 26108 21062 26142
rect 20972 26080 21062 26108
rect 21990 26142 22080 26172
rect 21990 26108 22018 26142
rect 22052 26108 22080 26142
rect 21990 26080 22080 26108
rect 23008 26142 23098 26172
rect 23008 26108 23036 26142
rect 23070 26108 23098 26142
rect 23008 26080 23098 26108
rect 24026 26142 24116 26172
rect 24026 26108 24054 26142
rect 24088 26108 24116 26142
rect 24026 26080 24116 26108
rect 25044 26142 25134 26172
rect 25044 26108 25072 26142
rect 25106 26108 25134 26142
rect 25044 26080 25134 26108
rect 26062 26142 26152 26172
rect 26062 26108 26090 26142
rect 26124 26108 26152 26142
rect 26062 26080 26152 26108
rect 27080 26142 27170 26172
rect 27080 26108 27108 26142
rect 27142 26108 27170 26142
rect 27080 26080 27170 26108
rect 28098 26142 28188 26172
rect 28098 26108 28126 26142
rect 28160 26108 28188 26142
rect 28098 26080 28188 26108
rect 29116 26142 29206 26172
rect 29116 26108 29144 26142
rect 29178 26108 29206 26142
rect 29116 26080 29206 26108
rect 30134 26142 30224 26172
rect 30134 26108 30162 26142
rect 30196 26108 30224 26142
rect 30134 26080 30224 26108
rect 31152 26142 31242 26172
rect 31152 26108 31180 26142
rect 31214 26108 31242 26142
rect 31152 26080 31242 26108
rect 32170 26142 32260 26172
rect 32170 26108 32198 26142
rect 32232 26108 32260 26142
rect 32170 26080 32260 26108
rect 33188 26142 33278 26172
rect 33188 26108 33216 26142
rect 33250 26108 33278 26142
rect 33188 26080 33278 26108
rect 17670 25891 17686 25925
rect 18242 25891 18258 25925
rect 18688 25891 18704 25925
rect 19260 25891 19276 25925
rect 19706 25891 19722 25925
rect 20278 25891 20294 25925
rect 20724 25891 20740 25925
rect 21296 25891 21312 25925
rect 21742 25891 21758 25925
rect 22314 25891 22330 25925
rect 22760 25891 22776 25925
rect 23332 25891 23348 25925
rect 23778 25891 23794 25925
rect 24350 25891 24366 25925
rect 24796 25891 24812 25925
rect 25368 25891 25384 25925
rect 25814 25891 25830 25925
rect 26386 25891 26402 25925
rect 26832 25891 26848 25925
rect 27404 25891 27420 25925
rect 27850 25891 27866 25925
rect 28422 25891 28438 25925
rect 28868 25891 28884 25925
rect 29440 25891 29456 25925
rect 29886 25891 29902 25925
rect 30458 25891 30474 25925
rect 30904 25891 30920 25925
rect 31476 25891 31492 25925
rect 31922 25891 31938 25925
rect 32494 25891 32510 25925
rect 32940 25891 32956 25925
rect 33512 25891 33528 25925
rect 17438 25832 17472 25848
rect 17438 25240 17472 25256
rect 18456 25832 18490 25848
rect 18456 25240 18490 25256
rect 19474 25832 19508 25848
rect 19474 25240 19508 25256
rect 20492 25832 20526 25848
rect 20492 25240 20526 25256
rect 21510 25832 21544 25848
rect 21510 25240 21544 25256
rect 22528 25832 22562 25848
rect 22528 25240 22562 25256
rect 23546 25832 23580 25848
rect 23546 25240 23580 25256
rect 24564 25832 24598 25848
rect 24564 25240 24598 25256
rect 25582 25832 25616 25848
rect 25582 25240 25616 25256
rect 26600 25832 26634 25848
rect 26600 25240 26634 25256
rect 27618 25832 27652 25848
rect 27618 25240 27652 25256
rect 28636 25832 28670 25848
rect 28636 25240 28670 25256
rect 29654 25832 29688 25848
rect 29654 25240 29688 25256
rect 30672 25832 30706 25848
rect 30672 25240 30706 25256
rect 31690 25832 31724 25848
rect 31690 25240 31724 25256
rect 32708 25832 32742 25848
rect 32708 25240 32742 25256
rect 33726 25832 33760 25848
rect 33726 25240 33760 25256
rect 17670 25163 17686 25197
rect 18242 25163 18258 25197
rect 18688 25163 18704 25197
rect 19260 25163 19276 25197
rect 19706 25163 19722 25197
rect 20278 25163 20294 25197
rect 20724 25163 20740 25197
rect 21296 25163 21312 25197
rect 21742 25163 21758 25197
rect 22314 25163 22330 25197
rect 22760 25163 22776 25197
rect 23332 25163 23348 25197
rect 23778 25163 23794 25197
rect 24350 25163 24366 25197
rect 24796 25163 24812 25197
rect 25368 25163 25384 25197
rect 25814 25163 25830 25197
rect 26386 25163 26402 25197
rect 26832 25163 26848 25197
rect 27404 25163 27420 25197
rect 27850 25163 27866 25197
rect 28422 25163 28438 25197
rect 28868 25163 28884 25197
rect 29440 25163 29456 25197
rect 29886 25163 29902 25197
rect 30458 25163 30474 25197
rect 30904 25163 30920 25197
rect 31476 25163 31492 25197
rect 31922 25163 31938 25197
rect 32494 25163 32510 25197
rect 32940 25163 32956 25197
rect 33512 25163 33528 25197
rect 17918 24990 18008 25020
rect 17918 24956 17946 24990
rect 17980 24956 18008 24990
rect 17918 24928 18008 24956
rect 18936 24990 19026 25020
rect 18936 24956 18964 24990
rect 18998 24956 19026 24990
rect 18936 24928 19026 24956
rect 19954 24990 20044 25020
rect 19954 24956 19982 24990
rect 20016 24956 20044 24990
rect 19954 24928 20044 24956
rect 20972 24990 21062 25020
rect 20972 24956 21000 24990
rect 21034 24956 21062 24990
rect 20972 24928 21062 24956
rect 21990 24990 22080 25020
rect 21990 24956 22018 24990
rect 22052 24956 22080 24990
rect 21990 24928 22080 24956
rect 23008 24990 23098 25020
rect 23008 24956 23036 24990
rect 23070 24956 23098 24990
rect 23008 24928 23098 24956
rect 24026 24990 24116 25020
rect 24026 24956 24054 24990
rect 24088 24956 24116 24990
rect 24026 24928 24116 24956
rect 25044 24990 25134 25020
rect 25044 24956 25072 24990
rect 25106 24956 25134 24990
rect 25044 24928 25134 24956
rect 26062 24990 26152 25020
rect 26062 24956 26090 24990
rect 26124 24956 26152 24990
rect 26062 24928 26152 24956
rect 27080 24990 27170 25020
rect 27080 24956 27108 24990
rect 27142 24956 27170 24990
rect 27080 24928 27170 24956
rect 28098 24990 28188 25020
rect 28098 24956 28126 24990
rect 28160 24956 28188 24990
rect 28098 24928 28188 24956
rect 29116 24990 29206 25020
rect 29116 24956 29144 24990
rect 29178 24956 29206 24990
rect 29116 24928 29206 24956
rect 30134 24990 30224 25020
rect 30134 24956 30162 24990
rect 30196 24956 30224 24990
rect 30134 24928 30224 24956
rect 31152 24990 31242 25020
rect 31152 24956 31180 24990
rect 31214 24956 31242 24990
rect 31152 24928 31242 24956
rect 32170 24990 32260 25020
rect 32170 24956 32198 24990
rect 32232 24956 32260 24990
rect 32170 24928 32260 24956
rect 33188 24990 33278 25020
rect 33188 24956 33216 24990
rect 33250 24956 33278 24990
rect 33188 24928 33278 24956
rect 17670 24755 17686 24789
rect 18242 24755 18258 24789
rect 18688 24755 18704 24789
rect 19260 24755 19276 24789
rect 19706 24755 19722 24789
rect 20278 24755 20294 24789
rect 20724 24755 20740 24789
rect 21296 24755 21312 24789
rect 21742 24755 21758 24789
rect 22314 24755 22330 24789
rect 22760 24755 22776 24789
rect 23332 24755 23348 24789
rect 23778 24755 23794 24789
rect 24350 24755 24366 24789
rect 24796 24755 24812 24789
rect 25368 24755 25384 24789
rect 25814 24755 25830 24789
rect 26386 24755 26402 24789
rect 26832 24755 26848 24789
rect 27404 24755 27420 24789
rect 27850 24755 27866 24789
rect 28422 24755 28438 24789
rect 28868 24755 28884 24789
rect 29440 24755 29456 24789
rect 29886 24755 29902 24789
rect 30458 24755 30474 24789
rect 30904 24755 30920 24789
rect 31476 24755 31492 24789
rect 31922 24755 31938 24789
rect 32494 24755 32510 24789
rect 32940 24755 32956 24789
rect 33512 24755 33528 24789
rect 17438 24696 17472 24712
rect 17438 24104 17472 24120
rect 18456 24696 18490 24712
rect 18456 24104 18490 24120
rect 19474 24696 19508 24712
rect 19474 24104 19508 24120
rect 20492 24696 20526 24712
rect 20492 24104 20526 24120
rect 21510 24696 21544 24712
rect 21510 24104 21544 24120
rect 22528 24696 22562 24712
rect 22528 24104 22562 24120
rect 23546 24696 23580 24712
rect 23546 24104 23580 24120
rect 24564 24696 24598 24712
rect 24564 24104 24598 24120
rect 25582 24696 25616 24712
rect 25582 24104 25616 24120
rect 26600 24696 26634 24712
rect 26600 24104 26634 24120
rect 27618 24696 27652 24712
rect 27618 24104 27652 24120
rect 28636 24696 28670 24712
rect 28636 24104 28670 24120
rect 29654 24696 29688 24712
rect 29654 24104 29688 24120
rect 30672 24696 30706 24712
rect 30672 24104 30706 24120
rect 31690 24696 31724 24712
rect 31690 24104 31724 24120
rect 32708 24696 32742 24712
rect 32708 24104 32742 24120
rect 33726 24696 33760 24712
rect 33726 24104 33760 24120
rect 17670 24027 17686 24061
rect 18242 24027 18258 24061
rect 18688 24027 18704 24061
rect 19260 24027 19276 24061
rect 19706 24027 19722 24061
rect 20278 24027 20294 24061
rect 20724 24027 20740 24061
rect 21296 24027 21312 24061
rect 21742 24027 21758 24061
rect 22314 24027 22330 24061
rect 22760 24027 22776 24061
rect 23332 24027 23348 24061
rect 23778 24027 23794 24061
rect 24350 24027 24366 24061
rect 24796 24027 24812 24061
rect 25368 24027 25384 24061
rect 25814 24027 25830 24061
rect 26386 24027 26402 24061
rect 26832 24027 26848 24061
rect 27404 24027 27420 24061
rect 27850 24027 27866 24061
rect 28422 24027 28438 24061
rect 28868 24027 28884 24061
rect 29440 24027 29456 24061
rect 29886 24027 29902 24061
rect 30458 24027 30474 24061
rect 30904 24027 30920 24061
rect 31476 24027 31492 24061
rect 31922 24027 31938 24061
rect 32494 24027 32510 24061
rect 32940 24027 32956 24061
rect 33512 24027 33528 24061
rect 18936 23546 19026 23576
rect 18936 23512 18964 23546
rect 18998 23512 19026 23546
rect 18936 23484 19026 23512
rect 19954 23546 20044 23576
rect 19954 23512 19982 23546
rect 20016 23512 20044 23546
rect 19954 23484 20044 23512
rect 20972 23546 21062 23576
rect 20972 23512 21000 23546
rect 21034 23512 21062 23546
rect 20972 23484 21062 23512
rect 21990 23546 22080 23576
rect 21990 23512 22018 23546
rect 22052 23512 22080 23546
rect 21990 23484 22080 23512
rect 23008 23546 23098 23576
rect 23008 23512 23036 23546
rect 23070 23512 23098 23546
rect 23008 23484 23098 23512
rect 24026 23546 24116 23576
rect 24026 23512 24054 23546
rect 24088 23512 24116 23546
rect 24026 23484 24116 23512
rect 25044 23546 25134 23576
rect 25044 23512 25072 23546
rect 25106 23512 25134 23546
rect 25044 23484 25134 23512
rect 26062 23546 26152 23576
rect 26062 23512 26090 23546
rect 26124 23512 26152 23546
rect 26062 23484 26152 23512
rect 27080 23546 27170 23576
rect 27080 23512 27108 23546
rect 27142 23512 27170 23546
rect 27080 23484 27170 23512
rect 28098 23546 28188 23576
rect 28098 23512 28126 23546
rect 28160 23512 28188 23546
rect 28098 23484 28188 23512
rect 29116 23546 29206 23576
rect 29116 23512 29144 23546
rect 29178 23512 29206 23546
rect 29116 23484 29206 23512
rect 30134 23546 30224 23576
rect 30134 23512 30162 23546
rect 30196 23512 30224 23546
rect 30134 23484 30224 23512
rect 31152 23546 31242 23576
rect 31152 23512 31180 23546
rect 31214 23512 31242 23546
rect 31152 23484 31242 23512
rect 32170 23546 32260 23576
rect 32170 23512 32198 23546
rect 32232 23512 32260 23546
rect 32170 23484 32260 23512
rect 33188 23546 33278 23576
rect 33188 23512 33216 23546
rect 33250 23512 33278 23546
rect 33188 23484 33278 23512
rect 18656 22981 18672 23015
rect 19228 22981 19244 23015
rect 19674 22981 19690 23015
rect 20246 22981 20262 23015
rect 20692 22981 20708 23015
rect 21264 22981 21280 23015
rect 21710 22981 21726 23015
rect 22282 22981 22298 23015
rect 22728 22981 22744 23015
rect 23300 22981 23316 23015
rect 23746 22981 23762 23015
rect 24318 22981 24334 23015
rect 24764 22981 24780 23015
rect 25336 22981 25352 23015
rect 25782 22981 25798 23015
rect 26354 22981 26370 23015
rect 26800 22981 26816 23015
rect 27372 22981 27388 23015
rect 27818 22981 27834 23015
rect 28390 22981 28406 23015
rect 28836 22981 28852 23015
rect 29408 22981 29424 23015
rect 29854 22981 29870 23015
rect 30426 22981 30442 23015
rect 30872 22981 30888 23015
rect 31444 22981 31460 23015
rect 31890 22981 31906 23015
rect 32462 22981 32478 23015
rect 32908 22981 32924 23015
rect 33480 22981 33496 23015
rect 18424 22922 18458 22938
rect 18424 22330 18458 22346
rect 19442 22922 19476 22938
rect 19442 22330 19476 22346
rect 20460 22922 20494 22938
rect 20460 22330 20494 22346
rect 21478 22922 21512 22938
rect 21478 22330 21512 22346
rect 22496 22922 22530 22938
rect 22496 22330 22530 22346
rect 23514 22922 23548 22938
rect 23514 22330 23548 22346
rect 24532 22922 24566 22938
rect 24532 22330 24566 22346
rect 25550 22922 25584 22938
rect 25550 22330 25584 22346
rect 26568 22922 26602 22938
rect 26568 22330 26602 22346
rect 27586 22922 27620 22938
rect 27586 22330 27620 22346
rect 28604 22922 28638 22938
rect 28604 22330 28638 22346
rect 29622 22922 29656 22938
rect 29622 22330 29656 22346
rect 30640 22922 30674 22938
rect 30640 22330 30674 22346
rect 31658 22922 31692 22938
rect 31658 22330 31692 22346
rect 32676 22922 32710 22938
rect 32676 22330 32710 22346
rect 33694 22922 33728 22938
rect 33694 22330 33728 22346
rect 14662 22274 14752 22304
rect 14662 22240 14690 22274
rect 14724 22240 14752 22274
rect 14662 22212 14752 22240
rect 15680 22274 15770 22304
rect 15680 22240 15708 22274
rect 15742 22240 15770 22274
rect 15680 22212 15770 22240
rect 16698 22274 16788 22304
rect 16698 22240 16726 22274
rect 16760 22240 16788 22274
rect 18656 22253 18672 22287
rect 19228 22253 19244 22287
rect 19674 22253 19690 22287
rect 20246 22253 20262 22287
rect 20692 22253 20708 22287
rect 21264 22253 21280 22287
rect 21710 22253 21726 22287
rect 22282 22253 22298 22287
rect 22728 22253 22744 22287
rect 23300 22253 23316 22287
rect 23746 22253 23762 22287
rect 24318 22253 24334 22287
rect 24764 22253 24780 22287
rect 25336 22253 25352 22287
rect 25782 22253 25798 22287
rect 26354 22253 26370 22287
rect 26800 22253 26816 22287
rect 27372 22253 27388 22287
rect 27818 22253 27834 22287
rect 28390 22253 28406 22287
rect 28836 22253 28852 22287
rect 29408 22253 29424 22287
rect 29854 22253 29870 22287
rect 30426 22253 30442 22287
rect 30872 22253 30888 22287
rect 31444 22253 31460 22287
rect 31890 22253 31906 22287
rect 32462 22253 32478 22287
rect 32908 22253 32924 22287
rect 33480 22253 33496 22287
rect 16698 22212 16788 22240
rect 18936 22034 19026 22064
rect 18936 22000 18964 22034
rect 18998 22000 19026 22034
rect 18936 21972 19026 22000
rect 19954 22034 20044 22064
rect 19954 22000 19982 22034
rect 20016 22000 20044 22034
rect 19954 21972 20044 22000
rect 20972 22034 21062 22064
rect 20972 22000 21000 22034
rect 21034 22000 21062 22034
rect 20972 21972 21062 22000
rect 21990 22034 22080 22064
rect 21990 22000 22018 22034
rect 22052 22000 22080 22034
rect 21990 21972 22080 22000
rect 23008 22034 23098 22064
rect 23008 22000 23036 22034
rect 23070 22000 23098 22034
rect 23008 21972 23098 22000
rect 24026 22034 24116 22064
rect 24026 22000 24054 22034
rect 24088 22000 24116 22034
rect 24026 21972 24116 22000
rect 25044 22034 25134 22064
rect 25044 22000 25072 22034
rect 25106 22000 25134 22034
rect 25044 21972 25134 22000
rect 26062 22034 26152 22064
rect 26062 22000 26090 22034
rect 26124 22000 26152 22034
rect 26062 21972 26152 22000
rect 27080 22034 27170 22064
rect 27080 22000 27108 22034
rect 27142 22000 27170 22034
rect 27080 21972 27170 22000
rect 28098 22034 28188 22064
rect 28098 22000 28126 22034
rect 28160 22000 28188 22034
rect 28098 21972 28188 22000
rect 29116 22034 29206 22064
rect 29116 22000 29144 22034
rect 29178 22000 29206 22034
rect 29116 21972 29206 22000
rect 30134 22034 30224 22064
rect 30134 22000 30162 22034
rect 30196 22000 30224 22034
rect 30134 21972 30224 22000
rect 31152 22034 31242 22064
rect 31152 22000 31180 22034
rect 31214 22000 31242 22034
rect 31152 21972 31242 22000
rect 32170 22034 32260 22064
rect 32170 22000 32198 22034
rect 32232 22000 32260 22034
rect 32170 21972 32260 22000
rect 33188 22034 33278 22064
rect 33188 22000 33216 22034
rect 33250 22000 33278 22034
rect 33188 21972 33278 22000
rect 14648 21897 14664 21931
rect 14740 21897 14756 21931
rect 14866 21897 14882 21931
rect 14958 21897 14974 21931
rect 15084 21897 15100 21931
rect 15176 21897 15192 21931
rect 15302 21897 15318 21931
rect 15394 21897 15410 21931
rect 15520 21897 15536 21931
rect 15612 21897 15628 21931
rect 15738 21897 15754 21931
rect 15830 21897 15846 21931
rect 15956 21897 15972 21931
rect 16048 21897 16064 21931
rect 16174 21897 16190 21931
rect 16266 21897 16282 21931
rect 16392 21897 16408 21931
rect 16484 21897 16500 21931
rect 16610 21897 16626 21931
rect 16702 21897 16718 21931
rect 14576 21838 14610 21854
rect 14576 21446 14610 21462
rect 14794 21838 14828 21854
rect 14794 21446 14828 21462
rect 15012 21838 15046 21854
rect 15012 21446 15046 21462
rect 15230 21838 15264 21854
rect 15230 21446 15264 21462
rect 15448 21838 15482 21854
rect 15448 21446 15482 21462
rect 15666 21838 15700 21854
rect 15666 21446 15700 21462
rect 15884 21838 15918 21854
rect 15884 21446 15918 21462
rect 16102 21838 16136 21854
rect 16102 21446 16136 21462
rect 16320 21838 16354 21854
rect 16320 21446 16354 21462
rect 16538 21838 16572 21854
rect 16538 21446 16572 21462
rect 16756 21838 16790 21854
rect 18656 21725 18672 21759
rect 19228 21725 19244 21759
rect 19674 21725 19690 21759
rect 20246 21725 20262 21759
rect 20692 21725 20708 21759
rect 21264 21725 21280 21759
rect 21710 21725 21726 21759
rect 22282 21725 22298 21759
rect 22728 21725 22744 21759
rect 23300 21725 23316 21759
rect 23746 21725 23762 21759
rect 24318 21725 24334 21759
rect 24764 21725 24780 21759
rect 25336 21725 25352 21759
rect 25782 21725 25798 21759
rect 26354 21725 26370 21759
rect 26800 21725 26816 21759
rect 27372 21725 27388 21759
rect 27818 21725 27834 21759
rect 28390 21725 28406 21759
rect 28836 21725 28852 21759
rect 29408 21725 29424 21759
rect 29854 21725 29870 21759
rect 30426 21725 30442 21759
rect 30872 21725 30888 21759
rect 31444 21725 31460 21759
rect 31890 21725 31906 21759
rect 32462 21725 32478 21759
rect 32908 21725 32924 21759
rect 33480 21725 33496 21759
rect 16756 21446 16790 21462
rect 18424 21666 18458 21682
rect 14894 21403 14954 21404
rect 14648 21369 14664 21403
rect 14740 21369 14756 21403
rect 14866 21369 14882 21403
rect 14958 21369 14974 21403
rect 15084 21369 15100 21403
rect 15176 21369 15192 21403
rect 15302 21369 15318 21403
rect 15394 21369 15410 21403
rect 15520 21369 15536 21403
rect 15612 21369 15628 21403
rect 15738 21369 15754 21403
rect 15830 21369 15846 21403
rect 15956 21369 15972 21403
rect 16048 21369 16064 21403
rect 16174 21369 16190 21403
rect 16266 21369 16282 21403
rect 16392 21369 16408 21403
rect 16484 21369 16500 21403
rect 16610 21369 16626 21403
rect 16702 21369 16718 21403
rect 14620 21190 14710 21220
rect 14620 21156 14648 21190
rect 14682 21156 14710 21190
rect 14620 21128 14710 21156
rect 15638 21190 15728 21220
rect 15638 21156 15666 21190
rect 15700 21156 15728 21190
rect 15638 21128 15728 21156
rect 16656 21190 16746 21220
rect 16656 21156 16684 21190
rect 16718 21156 16746 21190
rect 16656 21128 16746 21156
rect 18424 21074 18458 21090
rect 19442 21666 19476 21682
rect 19442 21074 19476 21090
rect 20460 21666 20494 21682
rect 20460 21074 20494 21090
rect 21478 21666 21512 21682
rect 21478 21074 21512 21090
rect 22496 21666 22530 21682
rect 22496 21074 22530 21090
rect 23514 21666 23548 21682
rect 23514 21074 23548 21090
rect 24532 21666 24566 21682
rect 24532 21074 24566 21090
rect 25550 21666 25584 21682
rect 25550 21074 25584 21090
rect 26568 21666 26602 21682
rect 26568 21074 26602 21090
rect 27586 21666 27620 21682
rect 27586 21074 27620 21090
rect 28604 21666 28638 21682
rect 28604 21074 28638 21090
rect 29622 21666 29656 21682
rect 29622 21074 29656 21090
rect 30640 21666 30674 21682
rect 30640 21074 30674 21090
rect 31658 21666 31692 21682
rect 31658 21074 31692 21090
rect 32676 21666 32710 21682
rect 32676 21074 32710 21090
rect 33694 21666 33728 21682
rect 33694 21074 33728 21090
rect 18656 20997 18672 21031
rect 19228 20997 19244 21031
rect 19674 20997 19690 21031
rect 20246 20997 20262 21031
rect 20692 20997 20708 21031
rect 21264 20997 21280 21031
rect 21710 20997 21726 21031
rect 22282 20997 22298 21031
rect 22728 20997 22744 21031
rect 23300 20997 23316 21031
rect 23746 20997 23762 21031
rect 24318 20997 24334 21031
rect 24764 20997 24780 21031
rect 25336 20997 25352 21031
rect 25782 20997 25798 21031
rect 26354 20997 26370 21031
rect 26800 20997 26816 21031
rect 27372 20997 27388 21031
rect 27818 20997 27834 21031
rect 28390 20997 28406 21031
rect 28836 20997 28852 21031
rect 29408 20997 29424 21031
rect 29854 20997 29870 21031
rect 30426 20997 30442 21031
rect 30872 20997 30888 21031
rect 31444 20997 31460 21031
rect 31890 20997 31906 21031
rect 32462 20997 32478 21031
rect 32908 20997 32924 21031
rect 33480 20997 33496 21031
rect 14648 20959 14664 20993
rect 14740 20959 14756 20993
rect 14866 20959 14882 20993
rect 14958 20959 14974 20993
rect 15084 20959 15100 20993
rect 15176 20959 15192 20993
rect 15302 20959 15318 20993
rect 15394 20959 15410 20993
rect 15520 20959 15536 20993
rect 15612 20959 15628 20993
rect 15738 20959 15754 20993
rect 15830 20959 15846 20993
rect 15956 20959 15972 20993
rect 16048 20959 16064 20993
rect 16174 20959 16190 20993
rect 16266 20959 16282 20993
rect 16392 20959 16408 20993
rect 16484 20959 16500 20993
rect 16610 20959 16626 20993
rect 16702 20959 16718 20993
rect 14576 20900 14610 20916
rect 14576 20508 14610 20524
rect 14794 20900 14828 20916
rect 14794 20508 14828 20524
rect 15012 20900 15046 20916
rect 15012 20508 15046 20524
rect 15230 20900 15264 20916
rect 15230 20508 15264 20524
rect 15448 20900 15482 20916
rect 15448 20508 15482 20524
rect 15666 20900 15700 20916
rect 15666 20508 15700 20524
rect 15884 20900 15918 20916
rect 15884 20508 15918 20524
rect 16102 20900 16136 20916
rect 16102 20508 16136 20524
rect 16320 20900 16354 20916
rect 16320 20508 16354 20524
rect 16538 20900 16572 20916
rect 16538 20508 16572 20524
rect 16756 20900 16790 20916
rect 18894 20766 18984 20796
rect 18894 20732 18922 20766
rect 18956 20732 18984 20766
rect 18894 20704 18984 20732
rect 19912 20766 20002 20796
rect 19912 20732 19940 20766
rect 19974 20732 20002 20766
rect 19912 20704 20002 20732
rect 20930 20766 21020 20796
rect 20930 20732 20958 20766
rect 20992 20732 21020 20766
rect 20930 20704 21020 20732
rect 21948 20766 22038 20796
rect 21948 20732 21976 20766
rect 22010 20732 22038 20766
rect 21948 20704 22038 20732
rect 22966 20766 23056 20796
rect 22966 20732 22994 20766
rect 23028 20732 23056 20766
rect 22966 20704 23056 20732
rect 23984 20766 24074 20796
rect 23984 20732 24012 20766
rect 24046 20732 24074 20766
rect 23984 20704 24074 20732
rect 25002 20766 25092 20796
rect 25002 20732 25030 20766
rect 25064 20732 25092 20766
rect 25002 20704 25092 20732
rect 26020 20766 26110 20796
rect 26020 20732 26048 20766
rect 26082 20732 26110 20766
rect 26020 20704 26110 20732
rect 27038 20766 27128 20796
rect 27038 20732 27066 20766
rect 27100 20732 27128 20766
rect 27038 20704 27128 20732
rect 28056 20766 28146 20796
rect 28056 20732 28084 20766
rect 28118 20732 28146 20766
rect 28056 20704 28146 20732
rect 29074 20766 29164 20796
rect 29074 20732 29102 20766
rect 29136 20732 29164 20766
rect 29074 20704 29164 20732
rect 30092 20766 30182 20796
rect 30092 20732 30120 20766
rect 30154 20732 30182 20766
rect 30092 20704 30182 20732
rect 31110 20766 31200 20796
rect 31110 20732 31138 20766
rect 31172 20732 31200 20766
rect 31110 20704 31200 20732
rect 32128 20766 32218 20796
rect 32128 20732 32156 20766
rect 32190 20732 32218 20766
rect 32128 20704 32218 20732
rect 33146 20766 33236 20796
rect 33146 20732 33174 20766
rect 33208 20732 33236 20766
rect 33146 20704 33236 20732
rect 16756 20508 16790 20524
rect 18656 20469 18672 20503
rect 19228 20469 19244 20503
rect 19674 20469 19690 20503
rect 20246 20469 20262 20503
rect 20692 20469 20708 20503
rect 21264 20469 21280 20503
rect 21710 20469 21726 20503
rect 22282 20469 22298 20503
rect 22728 20469 22744 20503
rect 23300 20469 23316 20503
rect 23746 20469 23762 20503
rect 24318 20469 24334 20503
rect 24764 20469 24780 20503
rect 25336 20469 25352 20503
rect 25782 20469 25798 20503
rect 26354 20469 26370 20503
rect 26800 20469 26816 20503
rect 27372 20469 27388 20503
rect 27818 20469 27834 20503
rect 28390 20469 28406 20503
rect 28836 20469 28852 20503
rect 29408 20469 29424 20503
rect 29854 20469 29870 20503
rect 30426 20469 30442 20503
rect 30872 20469 30888 20503
rect 31444 20469 31460 20503
rect 31890 20469 31906 20503
rect 32462 20469 32478 20503
rect 32908 20469 32924 20503
rect 33480 20469 33496 20503
rect 15326 20465 15386 20466
rect 16198 20465 16258 20466
rect 14648 20431 14664 20465
rect 14740 20431 14756 20465
rect 14866 20431 14882 20465
rect 14958 20431 14974 20465
rect 15084 20431 15100 20465
rect 15176 20431 15192 20465
rect 15302 20431 15318 20465
rect 15394 20431 15410 20465
rect 15520 20431 15536 20465
rect 15612 20431 15628 20465
rect 15738 20431 15754 20465
rect 15830 20431 15846 20465
rect 15956 20431 15972 20465
rect 16048 20431 16064 20465
rect 16174 20431 16190 20465
rect 16266 20431 16282 20465
rect 16392 20431 16408 20465
rect 16484 20431 16500 20465
rect 16610 20431 16626 20465
rect 16702 20431 16718 20465
rect 18424 20410 18458 20426
rect 14592 20248 14682 20278
rect 14592 20214 14620 20248
rect 14654 20214 14682 20248
rect 14592 20186 14682 20214
rect 15610 20248 15700 20278
rect 15610 20214 15638 20248
rect 15672 20214 15700 20248
rect 15610 20186 15700 20214
rect 16628 20248 16718 20278
rect 16628 20214 16656 20248
rect 16690 20214 16718 20248
rect 16628 20186 16718 20214
rect 14648 20021 14664 20055
rect 14740 20021 14756 20055
rect 14866 20021 14882 20055
rect 14958 20021 14974 20055
rect 15084 20021 15100 20055
rect 15176 20021 15192 20055
rect 15302 20021 15318 20055
rect 15394 20021 15410 20055
rect 15520 20021 15536 20055
rect 15612 20021 15628 20055
rect 15738 20021 15754 20055
rect 15830 20021 15846 20055
rect 15956 20021 15972 20055
rect 16048 20021 16064 20055
rect 16174 20021 16190 20055
rect 16266 20021 16282 20055
rect 16392 20021 16408 20055
rect 16484 20021 16500 20055
rect 16610 20021 16626 20055
rect 16702 20021 16718 20055
rect 14888 20020 14948 20021
rect 15326 20020 15386 20021
rect 14576 19962 14610 19978
rect 14576 19570 14610 19586
rect 14794 19962 14828 19978
rect 14794 19570 14828 19586
rect 15012 19962 15046 19978
rect 15012 19570 15046 19586
rect 15230 19962 15264 19978
rect 15230 19570 15264 19586
rect 15448 19962 15482 19978
rect 15448 19570 15482 19586
rect 15666 19962 15700 19978
rect 15666 19570 15700 19586
rect 15884 19962 15918 19978
rect 15884 19570 15918 19586
rect 16102 19962 16136 19978
rect 16102 19570 16136 19586
rect 16320 19962 16354 19978
rect 16320 19570 16354 19586
rect 16538 19962 16572 19978
rect 16538 19570 16572 19586
rect 16756 19962 16790 19978
rect 18424 19818 18458 19834
rect 19442 20410 19476 20426
rect 19442 19818 19476 19834
rect 20460 20410 20494 20426
rect 20460 19818 20494 19834
rect 21478 20410 21512 20426
rect 21478 19818 21512 19834
rect 22496 20410 22530 20426
rect 22496 19818 22530 19834
rect 23514 20410 23548 20426
rect 23514 19818 23548 19834
rect 24532 20410 24566 20426
rect 24532 19818 24566 19834
rect 25550 20410 25584 20426
rect 25550 19818 25584 19834
rect 26568 20410 26602 20426
rect 26568 19818 26602 19834
rect 27586 20410 27620 20426
rect 27586 19818 27620 19834
rect 28604 20410 28638 20426
rect 28604 19818 28638 19834
rect 29622 20410 29656 20426
rect 29622 19818 29656 19834
rect 30640 20410 30674 20426
rect 30640 19818 30674 19834
rect 31658 20410 31692 20426
rect 31658 19818 31692 19834
rect 32676 20410 32710 20426
rect 32676 19818 32710 19834
rect 33694 20410 33728 20426
rect 33694 19818 33728 19834
rect 18656 19741 18672 19775
rect 19228 19741 19244 19775
rect 19674 19741 19690 19775
rect 20246 19741 20262 19775
rect 20692 19741 20708 19775
rect 21264 19741 21280 19775
rect 21710 19741 21726 19775
rect 22282 19741 22298 19775
rect 22728 19741 22744 19775
rect 23300 19741 23316 19775
rect 23746 19741 23762 19775
rect 24318 19741 24334 19775
rect 24764 19741 24780 19775
rect 25336 19741 25352 19775
rect 25782 19741 25798 19775
rect 26354 19741 26370 19775
rect 26800 19741 26816 19775
rect 27372 19741 27388 19775
rect 27818 19741 27834 19775
rect 28390 19741 28406 19775
rect 28836 19741 28852 19775
rect 29408 19741 29424 19775
rect 29854 19741 29870 19775
rect 30426 19741 30442 19775
rect 30872 19741 30888 19775
rect 31444 19741 31460 19775
rect 31890 19741 31906 19775
rect 32462 19741 32478 19775
rect 32908 19741 32924 19775
rect 33480 19741 33496 19775
rect 16756 19570 16790 19586
rect 18894 19528 18984 19558
rect 14648 19493 14664 19527
rect 14740 19493 14756 19527
rect 14866 19493 14882 19527
rect 14958 19493 14974 19527
rect 15084 19493 15100 19527
rect 15176 19493 15192 19527
rect 15302 19493 15318 19527
rect 15394 19493 15410 19527
rect 15520 19493 15536 19527
rect 15612 19493 15628 19527
rect 15738 19493 15754 19527
rect 15830 19493 15846 19527
rect 15956 19493 15972 19527
rect 16048 19493 16064 19527
rect 16174 19493 16190 19527
rect 16266 19493 16282 19527
rect 16392 19493 16408 19527
rect 16484 19493 16500 19527
rect 16610 19493 16626 19527
rect 16702 19493 16718 19527
rect 18894 19494 18922 19528
rect 18956 19494 18984 19528
rect 18894 19466 18984 19494
rect 19912 19528 20002 19558
rect 19912 19494 19940 19528
rect 19974 19494 20002 19528
rect 19912 19466 20002 19494
rect 20930 19528 21020 19558
rect 20930 19494 20958 19528
rect 20992 19494 21020 19528
rect 20930 19466 21020 19494
rect 21948 19528 22038 19558
rect 21948 19494 21976 19528
rect 22010 19494 22038 19528
rect 21948 19466 22038 19494
rect 22966 19528 23056 19558
rect 22966 19494 22994 19528
rect 23028 19494 23056 19528
rect 22966 19466 23056 19494
rect 23984 19528 24074 19558
rect 23984 19494 24012 19528
rect 24046 19494 24074 19528
rect 23984 19466 24074 19494
rect 25002 19528 25092 19558
rect 25002 19494 25030 19528
rect 25064 19494 25092 19528
rect 25002 19466 25092 19494
rect 26020 19528 26110 19558
rect 26020 19494 26048 19528
rect 26082 19494 26110 19528
rect 26020 19466 26110 19494
rect 27038 19528 27128 19558
rect 27038 19494 27066 19528
rect 27100 19494 27128 19528
rect 27038 19466 27128 19494
rect 28056 19528 28146 19558
rect 28056 19494 28084 19528
rect 28118 19494 28146 19528
rect 28056 19466 28146 19494
rect 29074 19528 29164 19558
rect 29074 19494 29102 19528
rect 29136 19494 29164 19528
rect 29074 19466 29164 19494
rect 30092 19528 30182 19558
rect 30092 19494 30120 19528
rect 30154 19494 30182 19528
rect 30092 19466 30182 19494
rect 31110 19528 31200 19558
rect 31110 19494 31138 19528
rect 31172 19494 31200 19528
rect 31110 19466 31200 19494
rect 32128 19528 32218 19558
rect 32128 19494 32156 19528
rect 32190 19494 32218 19528
rect 32128 19466 32218 19494
rect 33146 19528 33236 19558
rect 33146 19494 33174 19528
rect 33208 19494 33236 19528
rect 33146 19466 33236 19494
rect 14592 19334 14682 19364
rect 14592 19300 14620 19334
rect 14654 19300 14682 19334
rect 14592 19272 14682 19300
rect 15610 19334 15700 19364
rect 15610 19300 15638 19334
rect 15672 19300 15700 19334
rect 15610 19272 15700 19300
rect 16628 19334 16718 19364
rect 16628 19300 16656 19334
rect 16690 19300 16718 19334
rect 16628 19272 16718 19300
rect 18656 19213 18672 19247
rect 19228 19213 19244 19247
rect 19674 19213 19690 19247
rect 20246 19213 20262 19247
rect 20692 19213 20708 19247
rect 21264 19213 21280 19247
rect 21710 19213 21726 19247
rect 22282 19213 22298 19247
rect 22728 19213 22744 19247
rect 23300 19213 23316 19247
rect 23746 19213 23762 19247
rect 24318 19213 24334 19247
rect 24764 19213 24780 19247
rect 25336 19213 25352 19247
rect 25782 19213 25798 19247
rect 26354 19213 26370 19247
rect 26800 19213 26816 19247
rect 27372 19213 27388 19247
rect 27818 19213 27834 19247
rect 28390 19213 28406 19247
rect 28836 19213 28852 19247
rect 29408 19213 29424 19247
rect 29854 19213 29870 19247
rect 30426 19213 30442 19247
rect 30872 19213 30888 19247
rect 31444 19213 31460 19247
rect 31890 19213 31906 19247
rect 32462 19213 32478 19247
rect 32908 19213 32924 19247
rect 33480 19213 33496 19247
rect 18424 19154 18458 19170
rect 14648 19083 14664 19117
rect 14740 19083 14756 19117
rect 14866 19083 14882 19117
rect 14958 19083 14974 19117
rect 15084 19083 15100 19117
rect 15176 19083 15192 19117
rect 15302 19083 15318 19117
rect 15394 19083 15410 19117
rect 15520 19083 15536 19117
rect 15612 19083 15628 19117
rect 15738 19083 15754 19117
rect 15830 19083 15846 19117
rect 15956 19083 15972 19117
rect 16048 19083 16064 19117
rect 16174 19083 16190 19117
rect 16266 19083 16282 19117
rect 16392 19083 16408 19117
rect 16484 19083 16500 19117
rect 16610 19083 16626 19117
rect 16702 19083 16718 19117
rect 15330 19082 15390 19083
rect 14576 19024 14610 19040
rect 14576 18632 14610 18648
rect 14794 19024 14828 19040
rect 14794 18632 14828 18648
rect 15012 19024 15046 19040
rect 15012 18632 15046 18648
rect 15230 19024 15264 19040
rect 15230 18632 15264 18648
rect 15448 19024 15482 19040
rect 15448 18632 15482 18648
rect 15666 19024 15700 19040
rect 15666 18632 15700 18648
rect 15884 19024 15918 19040
rect 15884 18632 15918 18648
rect 16102 19024 16136 19040
rect 16102 18632 16136 18648
rect 16320 19024 16354 19040
rect 16320 18632 16354 18648
rect 16538 19024 16572 19040
rect 16538 18632 16572 18648
rect 16756 19024 16790 19040
rect 16756 18632 16790 18648
rect 14648 18555 14664 18589
rect 14740 18555 14756 18589
rect 14866 18555 14882 18589
rect 14958 18555 14974 18589
rect 15084 18555 15100 18589
rect 15176 18555 15192 18589
rect 15302 18555 15318 18589
rect 15394 18555 15410 18589
rect 15520 18555 15536 18589
rect 15612 18555 15628 18589
rect 15738 18555 15754 18589
rect 15830 18555 15846 18589
rect 15956 18555 15972 18589
rect 16048 18555 16064 18589
rect 16174 18555 16190 18589
rect 16266 18555 16282 18589
rect 16392 18555 16408 18589
rect 16484 18555 16500 18589
rect 16610 18555 16626 18589
rect 16702 18555 16718 18589
rect 18424 18562 18458 18578
rect 19442 19154 19476 19170
rect 19442 18562 19476 18578
rect 20460 19154 20494 19170
rect 20460 18562 20494 18578
rect 21478 19154 21512 19170
rect 21478 18562 21512 18578
rect 22496 19154 22530 19170
rect 22496 18562 22530 18578
rect 23514 19154 23548 19170
rect 23514 18562 23548 18578
rect 24532 19154 24566 19170
rect 24532 18562 24566 18578
rect 25550 19154 25584 19170
rect 25550 18562 25584 18578
rect 26568 19154 26602 19170
rect 26568 18562 26602 18578
rect 27586 19154 27620 19170
rect 27586 18562 27620 18578
rect 28604 19154 28638 19170
rect 28604 18562 28638 18578
rect 29622 19154 29656 19170
rect 29622 18562 29656 18578
rect 30640 19154 30674 19170
rect 30640 18562 30674 18578
rect 31658 19154 31692 19170
rect 31658 18562 31692 18578
rect 32676 19154 32710 19170
rect 32676 18562 32710 18578
rect 33694 19154 33728 19170
rect 33694 18562 33728 18578
rect 18656 18485 18672 18519
rect 19228 18485 19244 18519
rect 19674 18485 19690 18519
rect 20246 18485 20262 18519
rect 20692 18485 20708 18519
rect 21264 18485 21280 18519
rect 21710 18485 21726 18519
rect 22282 18485 22298 18519
rect 22728 18485 22744 18519
rect 23300 18485 23316 18519
rect 23746 18485 23762 18519
rect 24318 18485 24334 18519
rect 24764 18485 24780 18519
rect 25336 18485 25352 18519
rect 25782 18485 25798 18519
rect 26354 18485 26370 18519
rect 26800 18485 26816 18519
rect 27372 18485 27388 18519
rect 27818 18485 27834 18519
rect 28390 18485 28406 18519
rect 28836 18485 28852 18519
rect 29408 18485 29424 18519
rect 29854 18485 29870 18519
rect 30426 18485 30442 18519
rect 30872 18485 30888 18519
rect 31444 18485 31460 18519
rect 31890 18485 31906 18519
rect 32462 18485 32478 18519
rect 32908 18485 32924 18519
rect 33480 18485 33496 18519
rect 11328 17658 11428 17820
rect 65328 28100 65428 28262
rect 47264 25378 47310 25411
rect 49004 25378 49074 25411
rect 47264 25377 47360 25378
rect 48978 25377 49074 25378
rect 47264 25315 47298 25377
rect 49040 25316 49074 25377
rect 47458 25275 47474 25309
rect 47574 25275 47590 25309
rect 47716 25275 47732 25309
rect 47832 25275 47848 25309
rect 47974 25275 47990 25309
rect 48090 25275 48106 25309
rect 48232 25275 48248 25309
rect 48348 25275 48364 25309
rect 48490 25275 48506 25309
rect 48606 25275 48622 25309
rect 48748 25275 48764 25309
rect 48864 25275 48880 25309
rect 47378 25216 47412 25232
rect 47378 24824 47412 24840
rect 47636 25216 47670 25232
rect 47636 24824 47670 24840
rect 47894 25216 47928 25232
rect 47894 24824 47928 24840
rect 48152 25216 48186 25232
rect 48152 24824 48186 24840
rect 48410 25216 48444 25232
rect 48410 24824 48444 24840
rect 48668 25216 48702 25232
rect 48668 24824 48702 24840
rect 48926 25216 48960 25232
rect 48926 24824 48960 24840
rect 47458 24747 47474 24781
rect 47574 24747 47590 24781
rect 47716 24747 47732 24781
rect 47832 24747 47848 24781
rect 47974 24747 47990 24781
rect 48090 24747 48106 24781
rect 48232 24747 48248 24781
rect 48348 24747 48364 24781
rect 48490 24747 48506 24781
rect 48606 24747 48622 24781
rect 48748 24747 48764 24781
rect 48864 24747 48880 24781
rect 47264 24679 47298 24741
rect 49148 24875 49177 24909
rect 49211 24875 49269 24909
rect 49303 24875 49361 24909
rect 49395 24875 49424 24909
rect 49040 24679 49074 24740
rect 47264 24678 47360 24679
rect 47264 24645 47310 24678
rect 49004 24646 49074 24679
rect 48978 24645 49074 24646
rect 49214 24833 49280 24841
rect 49214 24799 49230 24833
rect 49264 24799 49280 24833
rect 49214 24765 49280 24799
rect 49214 24731 49230 24765
rect 49264 24731 49280 24765
rect 49214 24697 49280 24731
rect 49214 24663 49230 24697
rect 49264 24663 49280 24697
rect 49214 24645 49280 24663
rect 49314 24833 49356 24875
rect 49348 24799 49356 24833
rect 49314 24765 49356 24799
rect 49348 24731 49356 24765
rect 49314 24697 49356 24731
rect 49348 24663 49356 24697
rect 49314 24647 49356 24663
rect 49214 24586 49260 24645
rect 49255 24538 49260 24586
rect 49294 24608 49360 24611
rect 49294 24597 49311 24608
rect 49294 24563 49310 24597
rect 49357 24568 49360 24608
rect 49344 24563 49360 24568
rect 49214 24525 49260 24538
rect 49214 24513 49280 24525
rect 49214 24479 49230 24513
rect 49264 24479 49280 24513
rect 47264 24444 47334 24478
rect 49004 24444 49074 24478
rect 47264 24382 47298 24444
rect 49040 24382 49074 24444
rect 49214 24445 49280 24479
rect 49214 24411 49230 24445
rect 49264 24411 49280 24445
rect 49214 24399 49280 24411
rect 49314 24513 49360 24529
rect 49348 24479 49360 24513
rect 49314 24445 49360 24479
rect 49348 24411 49360 24445
rect 47458 24342 47474 24376
rect 47574 24342 47590 24376
rect 47716 24342 47732 24376
rect 47832 24342 47848 24376
rect 47974 24342 47990 24376
rect 48090 24342 48106 24376
rect 48232 24342 48248 24376
rect 48348 24342 48364 24376
rect 48490 24342 48506 24376
rect 48606 24342 48622 24376
rect 48748 24342 48764 24376
rect 48864 24342 48880 24376
rect 47378 24292 47412 24308
rect 47378 24100 47412 24116
rect 47636 24292 47670 24308
rect 47636 24100 47670 24116
rect 47894 24292 47928 24308
rect 47894 24100 47928 24116
rect 48152 24292 48186 24308
rect 48152 24100 48186 24116
rect 48410 24292 48444 24308
rect 48410 24100 48444 24116
rect 48668 24292 48702 24308
rect 48668 24100 48702 24116
rect 48926 24292 48960 24308
rect 48926 24100 48960 24116
rect 47458 24032 47474 24066
rect 47574 24032 47590 24066
rect 47716 24032 47732 24066
rect 47832 24032 47848 24066
rect 47974 24032 47990 24066
rect 48090 24032 48106 24066
rect 48232 24032 48248 24066
rect 48348 24032 48364 24066
rect 48490 24032 48506 24066
rect 48606 24032 48622 24066
rect 48748 24032 48764 24066
rect 48864 24032 48880 24066
rect 49314 24365 49360 24411
rect 49148 24331 49177 24365
rect 49211 24331 49269 24365
rect 49303 24331 49361 24365
rect 49395 24331 49424 24365
rect 47264 23964 47298 24026
rect 49040 23964 49074 24026
rect 47264 23930 47332 23964
rect 49006 23930 49074 23964
rect 47264 23378 47310 23411
rect 49004 23378 49074 23411
rect 47264 23377 47360 23378
rect 48978 23377 49074 23378
rect 47264 23315 47298 23377
rect 49040 23316 49074 23377
rect 47458 23275 47474 23309
rect 47574 23275 47590 23309
rect 47716 23275 47732 23309
rect 47832 23275 47848 23309
rect 47974 23275 47990 23309
rect 48090 23275 48106 23309
rect 48232 23275 48248 23309
rect 48348 23275 48364 23309
rect 48490 23275 48506 23309
rect 48606 23275 48622 23309
rect 48748 23275 48764 23309
rect 48864 23275 48880 23309
rect 47378 23216 47412 23232
rect 47378 22824 47412 22840
rect 47636 23216 47670 23232
rect 47636 22824 47670 22840
rect 47894 23216 47928 23232
rect 47894 22824 47928 22840
rect 48152 23216 48186 23232
rect 48152 22824 48186 22840
rect 48410 23216 48444 23232
rect 48410 22824 48444 22840
rect 48668 23216 48702 23232
rect 48668 22824 48702 22840
rect 48926 23216 48960 23232
rect 48926 22824 48960 22840
rect 47458 22747 47474 22781
rect 47574 22747 47590 22781
rect 47716 22747 47732 22781
rect 47832 22747 47848 22781
rect 47974 22747 47990 22781
rect 48090 22747 48106 22781
rect 48232 22747 48248 22781
rect 48348 22747 48364 22781
rect 48490 22747 48506 22781
rect 48606 22747 48622 22781
rect 48748 22747 48764 22781
rect 48864 22747 48880 22781
rect 47264 22679 47298 22741
rect 49148 22875 49177 22909
rect 49211 22875 49269 22909
rect 49303 22875 49361 22909
rect 49395 22875 49424 22909
rect 49040 22679 49074 22740
rect 47264 22678 47360 22679
rect 47264 22645 47310 22678
rect 49004 22646 49074 22679
rect 48978 22645 49074 22646
rect 49214 22833 49280 22841
rect 49214 22799 49230 22833
rect 49264 22799 49280 22833
rect 49214 22765 49280 22799
rect 49214 22731 49230 22765
rect 49264 22731 49280 22765
rect 49214 22697 49280 22731
rect 49214 22663 49230 22697
rect 49264 22663 49280 22697
rect 49214 22645 49280 22663
rect 49314 22833 49356 22875
rect 49348 22799 49356 22833
rect 49314 22765 49356 22799
rect 49348 22731 49356 22765
rect 49314 22697 49356 22731
rect 49348 22663 49356 22697
rect 49314 22647 49356 22663
rect 49214 22586 49260 22645
rect 49255 22538 49260 22586
rect 49294 22608 49360 22611
rect 49294 22597 49311 22608
rect 49294 22563 49310 22597
rect 49357 22568 49360 22608
rect 49344 22563 49360 22568
rect 49214 22525 49260 22538
rect 49214 22513 49280 22525
rect 49214 22479 49230 22513
rect 49264 22479 49280 22513
rect 47264 22444 47334 22478
rect 49004 22444 49074 22478
rect 47264 22382 47298 22444
rect 49040 22382 49074 22444
rect 49214 22445 49280 22479
rect 49214 22411 49230 22445
rect 49264 22411 49280 22445
rect 49214 22399 49280 22411
rect 49314 22513 49360 22529
rect 49348 22479 49360 22513
rect 49314 22445 49360 22479
rect 49348 22411 49360 22445
rect 47458 22342 47474 22376
rect 47574 22342 47590 22376
rect 47716 22342 47732 22376
rect 47832 22342 47848 22376
rect 47974 22342 47990 22376
rect 48090 22342 48106 22376
rect 48232 22342 48248 22376
rect 48348 22342 48364 22376
rect 48490 22342 48506 22376
rect 48606 22342 48622 22376
rect 48748 22342 48764 22376
rect 48864 22342 48880 22376
rect 47378 22292 47412 22308
rect 47378 22100 47412 22116
rect 47636 22292 47670 22308
rect 47636 22100 47670 22116
rect 47894 22292 47928 22308
rect 47894 22100 47928 22116
rect 48152 22292 48186 22308
rect 48152 22100 48186 22116
rect 48410 22292 48444 22308
rect 48410 22100 48444 22116
rect 48668 22292 48702 22308
rect 48668 22100 48702 22116
rect 48926 22292 48960 22308
rect 48926 22100 48960 22116
rect 47458 22032 47474 22066
rect 47574 22032 47590 22066
rect 47716 22032 47732 22066
rect 47832 22032 47848 22066
rect 47974 22032 47990 22066
rect 48090 22032 48106 22066
rect 48232 22032 48248 22066
rect 48348 22032 48364 22066
rect 48490 22032 48506 22066
rect 48606 22032 48622 22066
rect 48748 22032 48764 22066
rect 48864 22032 48880 22066
rect 49314 22365 49360 22411
rect 49148 22331 49177 22365
rect 49211 22331 49269 22365
rect 49303 22331 49361 22365
rect 49395 22331 49424 22365
rect 47264 21964 47298 22026
rect 49040 21964 49074 22026
rect 47264 21930 47332 21964
rect 49006 21930 49074 21964
rect 35672 17658 35772 17820
rect 89672 28100 89772 28262
rect 71670 27027 71686 27061
rect 72242 27027 72258 27061
rect 72688 27027 72704 27061
rect 73260 27027 73276 27061
rect 73706 27027 73722 27061
rect 74278 27027 74294 27061
rect 74724 27027 74740 27061
rect 75296 27027 75312 27061
rect 75742 27027 75758 27061
rect 76314 27027 76330 27061
rect 76760 27027 76776 27061
rect 77332 27027 77348 27061
rect 77778 27027 77794 27061
rect 78350 27027 78366 27061
rect 78796 27027 78812 27061
rect 79368 27027 79384 27061
rect 79814 27027 79830 27061
rect 80386 27027 80402 27061
rect 80832 27027 80848 27061
rect 81404 27027 81420 27061
rect 81850 27027 81866 27061
rect 82422 27027 82438 27061
rect 82868 27027 82884 27061
rect 83440 27027 83456 27061
rect 83886 27027 83902 27061
rect 84458 27027 84474 27061
rect 84904 27027 84920 27061
rect 85476 27027 85492 27061
rect 85922 27027 85938 27061
rect 86494 27027 86510 27061
rect 86940 27027 86956 27061
rect 87512 27027 87528 27061
rect 71438 26968 71472 26984
rect 71438 26376 71472 26392
rect 72456 26968 72490 26984
rect 72456 26376 72490 26392
rect 73474 26968 73508 26984
rect 73474 26376 73508 26392
rect 74492 26968 74526 26984
rect 74492 26376 74526 26392
rect 75510 26968 75544 26984
rect 75510 26376 75544 26392
rect 76528 26968 76562 26984
rect 76528 26376 76562 26392
rect 77546 26968 77580 26984
rect 77546 26376 77580 26392
rect 78564 26968 78598 26984
rect 78564 26376 78598 26392
rect 79582 26968 79616 26984
rect 79582 26376 79616 26392
rect 80600 26968 80634 26984
rect 80600 26376 80634 26392
rect 81618 26968 81652 26984
rect 81618 26376 81652 26392
rect 82636 26968 82670 26984
rect 82636 26376 82670 26392
rect 83654 26968 83688 26984
rect 83654 26376 83688 26392
rect 84672 26968 84706 26984
rect 84672 26376 84706 26392
rect 85690 26968 85724 26984
rect 85690 26376 85724 26392
rect 86708 26968 86742 26984
rect 86708 26376 86742 26392
rect 87726 26968 87760 26984
rect 87726 26376 87760 26392
rect 71670 26299 71686 26333
rect 72242 26299 72258 26333
rect 72688 26299 72704 26333
rect 73260 26299 73276 26333
rect 73706 26299 73722 26333
rect 74278 26299 74294 26333
rect 74724 26299 74740 26333
rect 75296 26299 75312 26333
rect 75742 26299 75758 26333
rect 76314 26299 76330 26333
rect 76760 26299 76776 26333
rect 77332 26299 77348 26333
rect 77778 26299 77794 26333
rect 78350 26299 78366 26333
rect 78796 26299 78812 26333
rect 79368 26299 79384 26333
rect 79814 26299 79830 26333
rect 80386 26299 80402 26333
rect 80832 26299 80848 26333
rect 81404 26299 81420 26333
rect 81850 26299 81866 26333
rect 82422 26299 82438 26333
rect 82868 26299 82884 26333
rect 83440 26299 83456 26333
rect 83886 26299 83902 26333
rect 84458 26299 84474 26333
rect 84904 26299 84920 26333
rect 85476 26299 85492 26333
rect 85922 26299 85938 26333
rect 86494 26299 86510 26333
rect 86940 26299 86956 26333
rect 87512 26299 87528 26333
rect 72936 26142 73026 26172
rect 72936 26108 72964 26142
rect 72998 26108 73026 26142
rect 72936 26080 73026 26108
rect 73954 26142 74044 26172
rect 73954 26108 73982 26142
rect 74016 26108 74044 26142
rect 73954 26080 74044 26108
rect 74972 26142 75062 26172
rect 74972 26108 75000 26142
rect 75034 26108 75062 26142
rect 74972 26080 75062 26108
rect 75990 26142 76080 26172
rect 75990 26108 76018 26142
rect 76052 26108 76080 26142
rect 75990 26080 76080 26108
rect 77008 26142 77098 26172
rect 77008 26108 77036 26142
rect 77070 26108 77098 26142
rect 77008 26080 77098 26108
rect 78026 26142 78116 26172
rect 78026 26108 78054 26142
rect 78088 26108 78116 26142
rect 78026 26080 78116 26108
rect 79044 26142 79134 26172
rect 79044 26108 79072 26142
rect 79106 26108 79134 26142
rect 79044 26080 79134 26108
rect 80062 26142 80152 26172
rect 80062 26108 80090 26142
rect 80124 26108 80152 26142
rect 80062 26080 80152 26108
rect 81080 26142 81170 26172
rect 81080 26108 81108 26142
rect 81142 26108 81170 26142
rect 81080 26080 81170 26108
rect 82098 26142 82188 26172
rect 82098 26108 82126 26142
rect 82160 26108 82188 26142
rect 82098 26080 82188 26108
rect 83116 26142 83206 26172
rect 83116 26108 83144 26142
rect 83178 26108 83206 26142
rect 83116 26080 83206 26108
rect 84134 26142 84224 26172
rect 84134 26108 84162 26142
rect 84196 26108 84224 26142
rect 84134 26080 84224 26108
rect 85152 26142 85242 26172
rect 85152 26108 85180 26142
rect 85214 26108 85242 26142
rect 85152 26080 85242 26108
rect 86170 26142 86260 26172
rect 86170 26108 86198 26142
rect 86232 26108 86260 26142
rect 86170 26080 86260 26108
rect 87188 26142 87278 26172
rect 87188 26108 87216 26142
rect 87250 26108 87278 26142
rect 87188 26080 87278 26108
rect 71670 25891 71686 25925
rect 72242 25891 72258 25925
rect 72688 25891 72704 25925
rect 73260 25891 73276 25925
rect 73706 25891 73722 25925
rect 74278 25891 74294 25925
rect 74724 25891 74740 25925
rect 75296 25891 75312 25925
rect 75742 25891 75758 25925
rect 76314 25891 76330 25925
rect 76760 25891 76776 25925
rect 77332 25891 77348 25925
rect 77778 25891 77794 25925
rect 78350 25891 78366 25925
rect 78796 25891 78812 25925
rect 79368 25891 79384 25925
rect 79814 25891 79830 25925
rect 80386 25891 80402 25925
rect 80832 25891 80848 25925
rect 81404 25891 81420 25925
rect 81850 25891 81866 25925
rect 82422 25891 82438 25925
rect 82868 25891 82884 25925
rect 83440 25891 83456 25925
rect 83886 25891 83902 25925
rect 84458 25891 84474 25925
rect 84904 25891 84920 25925
rect 85476 25891 85492 25925
rect 85922 25891 85938 25925
rect 86494 25891 86510 25925
rect 86940 25891 86956 25925
rect 87512 25891 87528 25925
rect 71438 25832 71472 25848
rect 71438 25240 71472 25256
rect 72456 25832 72490 25848
rect 72456 25240 72490 25256
rect 73474 25832 73508 25848
rect 73474 25240 73508 25256
rect 74492 25832 74526 25848
rect 74492 25240 74526 25256
rect 75510 25832 75544 25848
rect 75510 25240 75544 25256
rect 76528 25832 76562 25848
rect 76528 25240 76562 25256
rect 77546 25832 77580 25848
rect 77546 25240 77580 25256
rect 78564 25832 78598 25848
rect 78564 25240 78598 25256
rect 79582 25832 79616 25848
rect 79582 25240 79616 25256
rect 80600 25832 80634 25848
rect 80600 25240 80634 25256
rect 81618 25832 81652 25848
rect 81618 25240 81652 25256
rect 82636 25832 82670 25848
rect 82636 25240 82670 25256
rect 83654 25832 83688 25848
rect 83654 25240 83688 25256
rect 84672 25832 84706 25848
rect 84672 25240 84706 25256
rect 85690 25832 85724 25848
rect 85690 25240 85724 25256
rect 86708 25832 86742 25848
rect 86708 25240 86742 25256
rect 87726 25832 87760 25848
rect 87726 25240 87760 25256
rect 71670 25163 71686 25197
rect 72242 25163 72258 25197
rect 72688 25163 72704 25197
rect 73260 25163 73276 25197
rect 73706 25163 73722 25197
rect 74278 25163 74294 25197
rect 74724 25163 74740 25197
rect 75296 25163 75312 25197
rect 75742 25163 75758 25197
rect 76314 25163 76330 25197
rect 76760 25163 76776 25197
rect 77332 25163 77348 25197
rect 77778 25163 77794 25197
rect 78350 25163 78366 25197
rect 78796 25163 78812 25197
rect 79368 25163 79384 25197
rect 79814 25163 79830 25197
rect 80386 25163 80402 25197
rect 80832 25163 80848 25197
rect 81404 25163 81420 25197
rect 81850 25163 81866 25197
rect 82422 25163 82438 25197
rect 82868 25163 82884 25197
rect 83440 25163 83456 25197
rect 83886 25163 83902 25197
rect 84458 25163 84474 25197
rect 84904 25163 84920 25197
rect 85476 25163 85492 25197
rect 85922 25163 85938 25197
rect 86494 25163 86510 25197
rect 86940 25163 86956 25197
rect 87512 25163 87528 25197
rect 71918 24990 72008 25020
rect 71918 24956 71946 24990
rect 71980 24956 72008 24990
rect 71918 24928 72008 24956
rect 72936 24990 73026 25020
rect 72936 24956 72964 24990
rect 72998 24956 73026 24990
rect 72936 24928 73026 24956
rect 73954 24990 74044 25020
rect 73954 24956 73982 24990
rect 74016 24956 74044 24990
rect 73954 24928 74044 24956
rect 74972 24990 75062 25020
rect 74972 24956 75000 24990
rect 75034 24956 75062 24990
rect 74972 24928 75062 24956
rect 75990 24990 76080 25020
rect 75990 24956 76018 24990
rect 76052 24956 76080 24990
rect 75990 24928 76080 24956
rect 77008 24990 77098 25020
rect 77008 24956 77036 24990
rect 77070 24956 77098 24990
rect 77008 24928 77098 24956
rect 78026 24990 78116 25020
rect 78026 24956 78054 24990
rect 78088 24956 78116 24990
rect 78026 24928 78116 24956
rect 79044 24990 79134 25020
rect 79044 24956 79072 24990
rect 79106 24956 79134 24990
rect 79044 24928 79134 24956
rect 80062 24990 80152 25020
rect 80062 24956 80090 24990
rect 80124 24956 80152 24990
rect 80062 24928 80152 24956
rect 81080 24990 81170 25020
rect 81080 24956 81108 24990
rect 81142 24956 81170 24990
rect 81080 24928 81170 24956
rect 82098 24990 82188 25020
rect 82098 24956 82126 24990
rect 82160 24956 82188 24990
rect 82098 24928 82188 24956
rect 83116 24990 83206 25020
rect 83116 24956 83144 24990
rect 83178 24956 83206 24990
rect 83116 24928 83206 24956
rect 84134 24990 84224 25020
rect 84134 24956 84162 24990
rect 84196 24956 84224 24990
rect 84134 24928 84224 24956
rect 85152 24990 85242 25020
rect 85152 24956 85180 24990
rect 85214 24956 85242 24990
rect 85152 24928 85242 24956
rect 86170 24990 86260 25020
rect 86170 24956 86198 24990
rect 86232 24956 86260 24990
rect 86170 24928 86260 24956
rect 87188 24990 87278 25020
rect 87188 24956 87216 24990
rect 87250 24956 87278 24990
rect 87188 24928 87278 24956
rect 71670 24755 71686 24789
rect 72242 24755 72258 24789
rect 72688 24755 72704 24789
rect 73260 24755 73276 24789
rect 73706 24755 73722 24789
rect 74278 24755 74294 24789
rect 74724 24755 74740 24789
rect 75296 24755 75312 24789
rect 75742 24755 75758 24789
rect 76314 24755 76330 24789
rect 76760 24755 76776 24789
rect 77332 24755 77348 24789
rect 77778 24755 77794 24789
rect 78350 24755 78366 24789
rect 78796 24755 78812 24789
rect 79368 24755 79384 24789
rect 79814 24755 79830 24789
rect 80386 24755 80402 24789
rect 80832 24755 80848 24789
rect 81404 24755 81420 24789
rect 81850 24755 81866 24789
rect 82422 24755 82438 24789
rect 82868 24755 82884 24789
rect 83440 24755 83456 24789
rect 83886 24755 83902 24789
rect 84458 24755 84474 24789
rect 84904 24755 84920 24789
rect 85476 24755 85492 24789
rect 85922 24755 85938 24789
rect 86494 24755 86510 24789
rect 86940 24755 86956 24789
rect 87512 24755 87528 24789
rect 71438 24696 71472 24712
rect 71438 24104 71472 24120
rect 72456 24696 72490 24712
rect 72456 24104 72490 24120
rect 73474 24696 73508 24712
rect 73474 24104 73508 24120
rect 74492 24696 74526 24712
rect 74492 24104 74526 24120
rect 75510 24696 75544 24712
rect 75510 24104 75544 24120
rect 76528 24696 76562 24712
rect 76528 24104 76562 24120
rect 77546 24696 77580 24712
rect 77546 24104 77580 24120
rect 78564 24696 78598 24712
rect 78564 24104 78598 24120
rect 79582 24696 79616 24712
rect 79582 24104 79616 24120
rect 80600 24696 80634 24712
rect 80600 24104 80634 24120
rect 81618 24696 81652 24712
rect 81618 24104 81652 24120
rect 82636 24696 82670 24712
rect 82636 24104 82670 24120
rect 83654 24696 83688 24712
rect 83654 24104 83688 24120
rect 84672 24696 84706 24712
rect 84672 24104 84706 24120
rect 85690 24696 85724 24712
rect 85690 24104 85724 24120
rect 86708 24696 86742 24712
rect 86708 24104 86742 24120
rect 87726 24696 87760 24712
rect 87726 24104 87760 24120
rect 71670 24027 71686 24061
rect 72242 24027 72258 24061
rect 72688 24027 72704 24061
rect 73260 24027 73276 24061
rect 73706 24027 73722 24061
rect 74278 24027 74294 24061
rect 74724 24027 74740 24061
rect 75296 24027 75312 24061
rect 75742 24027 75758 24061
rect 76314 24027 76330 24061
rect 76760 24027 76776 24061
rect 77332 24027 77348 24061
rect 77778 24027 77794 24061
rect 78350 24027 78366 24061
rect 78796 24027 78812 24061
rect 79368 24027 79384 24061
rect 79814 24027 79830 24061
rect 80386 24027 80402 24061
rect 80832 24027 80848 24061
rect 81404 24027 81420 24061
rect 81850 24027 81866 24061
rect 82422 24027 82438 24061
rect 82868 24027 82884 24061
rect 83440 24027 83456 24061
rect 83886 24027 83902 24061
rect 84458 24027 84474 24061
rect 84904 24027 84920 24061
rect 85476 24027 85492 24061
rect 85922 24027 85938 24061
rect 86494 24027 86510 24061
rect 86940 24027 86956 24061
rect 87512 24027 87528 24061
rect 72936 23546 73026 23576
rect 72936 23512 72964 23546
rect 72998 23512 73026 23546
rect 72936 23484 73026 23512
rect 73954 23546 74044 23576
rect 73954 23512 73982 23546
rect 74016 23512 74044 23546
rect 73954 23484 74044 23512
rect 74972 23546 75062 23576
rect 74972 23512 75000 23546
rect 75034 23512 75062 23546
rect 74972 23484 75062 23512
rect 75990 23546 76080 23576
rect 75990 23512 76018 23546
rect 76052 23512 76080 23546
rect 75990 23484 76080 23512
rect 77008 23546 77098 23576
rect 77008 23512 77036 23546
rect 77070 23512 77098 23546
rect 77008 23484 77098 23512
rect 78026 23546 78116 23576
rect 78026 23512 78054 23546
rect 78088 23512 78116 23546
rect 78026 23484 78116 23512
rect 79044 23546 79134 23576
rect 79044 23512 79072 23546
rect 79106 23512 79134 23546
rect 79044 23484 79134 23512
rect 80062 23546 80152 23576
rect 80062 23512 80090 23546
rect 80124 23512 80152 23546
rect 80062 23484 80152 23512
rect 81080 23546 81170 23576
rect 81080 23512 81108 23546
rect 81142 23512 81170 23546
rect 81080 23484 81170 23512
rect 82098 23546 82188 23576
rect 82098 23512 82126 23546
rect 82160 23512 82188 23546
rect 82098 23484 82188 23512
rect 83116 23546 83206 23576
rect 83116 23512 83144 23546
rect 83178 23512 83206 23546
rect 83116 23484 83206 23512
rect 84134 23546 84224 23576
rect 84134 23512 84162 23546
rect 84196 23512 84224 23546
rect 84134 23484 84224 23512
rect 85152 23546 85242 23576
rect 85152 23512 85180 23546
rect 85214 23512 85242 23546
rect 85152 23484 85242 23512
rect 86170 23546 86260 23576
rect 86170 23512 86198 23546
rect 86232 23512 86260 23546
rect 86170 23484 86260 23512
rect 87188 23546 87278 23576
rect 87188 23512 87216 23546
rect 87250 23512 87278 23546
rect 87188 23484 87278 23512
rect 72656 22981 72672 23015
rect 73228 22981 73244 23015
rect 73674 22981 73690 23015
rect 74246 22981 74262 23015
rect 74692 22981 74708 23015
rect 75264 22981 75280 23015
rect 75710 22981 75726 23015
rect 76282 22981 76298 23015
rect 76728 22981 76744 23015
rect 77300 22981 77316 23015
rect 77746 22981 77762 23015
rect 78318 22981 78334 23015
rect 78764 22981 78780 23015
rect 79336 22981 79352 23015
rect 79782 22981 79798 23015
rect 80354 22981 80370 23015
rect 80800 22981 80816 23015
rect 81372 22981 81388 23015
rect 81818 22981 81834 23015
rect 82390 22981 82406 23015
rect 82836 22981 82852 23015
rect 83408 22981 83424 23015
rect 83854 22981 83870 23015
rect 84426 22981 84442 23015
rect 84872 22981 84888 23015
rect 85444 22981 85460 23015
rect 85890 22981 85906 23015
rect 86462 22981 86478 23015
rect 86908 22981 86924 23015
rect 87480 22981 87496 23015
rect 72424 22922 72458 22938
rect 72424 22330 72458 22346
rect 73442 22922 73476 22938
rect 73442 22330 73476 22346
rect 74460 22922 74494 22938
rect 74460 22330 74494 22346
rect 75478 22922 75512 22938
rect 75478 22330 75512 22346
rect 76496 22922 76530 22938
rect 76496 22330 76530 22346
rect 77514 22922 77548 22938
rect 77514 22330 77548 22346
rect 78532 22922 78566 22938
rect 78532 22330 78566 22346
rect 79550 22922 79584 22938
rect 79550 22330 79584 22346
rect 80568 22922 80602 22938
rect 80568 22330 80602 22346
rect 81586 22922 81620 22938
rect 81586 22330 81620 22346
rect 82604 22922 82638 22938
rect 82604 22330 82638 22346
rect 83622 22922 83656 22938
rect 83622 22330 83656 22346
rect 84640 22922 84674 22938
rect 84640 22330 84674 22346
rect 85658 22922 85692 22938
rect 85658 22330 85692 22346
rect 86676 22922 86710 22938
rect 86676 22330 86710 22346
rect 87694 22922 87728 22938
rect 87694 22330 87728 22346
rect 68662 22274 68752 22304
rect 68662 22240 68690 22274
rect 68724 22240 68752 22274
rect 68662 22212 68752 22240
rect 69680 22274 69770 22304
rect 69680 22240 69708 22274
rect 69742 22240 69770 22274
rect 69680 22212 69770 22240
rect 70698 22274 70788 22304
rect 70698 22240 70726 22274
rect 70760 22240 70788 22274
rect 72656 22253 72672 22287
rect 73228 22253 73244 22287
rect 73674 22253 73690 22287
rect 74246 22253 74262 22287
rect 74692 22253 74708 22287
rect 75264 22253 75280 22287
rect 75710 22253 75726 22287
rect 76282 22253 76298 22287
rect 76728 22253 76744 22287
rect 77300 22253 77316 22287
rect 77746 22253 77762 22287
rect 78318 22253 78334 22287
rect 78764 22253 78780 22287
rect 79336 22253 79352 22287
rect 79782 22253 79798 22287
rect 80354 22253 80370 22287
rect 80800 22253 80816 22287
rect 81372 22253 81388 22287
rect 81818 22253 81834 22287
rect 82390 22253 82406 22287
rect 82836 22253 82852 22287
rect 83408 22253 83424 22287
rect 83854 22253 83870 22287
rect 84426 22253 84442 22287
rect 84872 22253 84888 22287
rect 85444 22253 85460 22287
rect 85890 22253 85906 22287
rect 86462 22253 86478 22287
rect 86908 22253 86924 22287
rect 87480 22253 87496 22287
rect 70698 22212 70788 22240
rect 72936 22034 73026 22064
rect 72936 22000 72964 22034
rect 72998 22000 73026 22034
rect 72936 21972 73026 22000
rect 73954 22034 74044 22064
rect 73954 22000 73982 22034
rect 74016 22000 74044 22034
rect 73954 21972 74044 22000
rect 74972 22034 75062 22064
rect 74972 22000 75000 22034
rect 75034 22000 75062 22034
rect 74972 21972 75062 22000
rect 75990 22034 76080 22064
rect 75990 22000 76018 22034
rect 76052 22000 76080 22034
rect 75990 21972 76080 22000
rect 77008 22034 77098 22064
rect 77008 22000 77036 22034
rect 77070 22000 77098 22034
rect 77008 21972 77098 22000
rect 78026 22034 78116 22064
rect 78026 22000 78054 22034
rect 78088 22000 78116 22034
rect 78026 21972 78116 22000
rect 79044 22034 79134 22064
rect 79044 22000 79072 22034
rect 79106 22000 79134 22034
rect 79044 21972 79134 22000
rect 80062 22034 80152 22064
rect 80062 22000 80090 22034
rect 80124 22000 80152 22034
rect 80062 21972 80152 22000
rect 81080 22034 81170 22064
rect 81080 22000 81108 22034
rect 81142 22000 81170 22034
rect 81080 21972 81170 22000
rect 82098 22034 82188 22064
rect 82098 22000 82126 22034
rect 82160 22000 82188 22034
rect 82098 21972 82188 22000
rect 83116 22034 83206 22064
rect 83116 22000 83144 22034
rect 83178 22000 83206 22034
rect 83116 21972 83206 22000
rect 84134 22034 84224 22064
rect 84134 22000 84162 22034
rect 84196 22000 84224 22034
rect 84134 21972 84224 22000
rect 85152 22034 85242 22064
rect 85152 22000 85180 22034
rect 85214 22000 85242 22034
rect 85152 21972 85242 22000
rect 86170 22034 86260 22064
rect 86170 22000 86198 22034
rect 86232 22000 86260 22034
rect 86170 21972 86260 22000
rect 87188 22034 87278 22064
rect 87188 22000 87216 22034
rect 87250 22000 87278 22034
rect 87188 21972 87278 22000
rect 68648 21897 68664 21931
rect 68740 21897 68756 21931
rect 68866 21897 68882 21931
rect 68958 21897 68974 21931
rect 69084 21897 69100 21931
rect 69176 21897 69192 21931
rect 69302 21897 69318 21931
rect 69394 21897 69410 21931
rect 69520 21897 69536 21931
rect 69612 21897 69628 21931
rect 69738 21897 69754 21931
rect 69830 21897 69846 21931
rect 69956 21897 69972 21931
rect 70048 21897 70064 21931
rect 70174 21897 70190 21931
rect 70266 21897 70282 21931
rect 70392 21897 70408 21931
rect 70484 21897 70500 21931
rect 70610 21897 70626 21931
rect 70702 21897 70718 21931
rect 68576 21838 68610 21854
rect 68576 21446 68610 21462
rect 68794 21838 68828 21854
rect 68794 21446 68828 21462
rect 69012 21838 69046 21854
rect 69012 21446 69046 21462
rect 69230 21838 69264 21854
rect 69230 21446 69264 21462
rect 69448 21838 69482 21854
rect 69448 21446 69482 21462
rect 69666 21838 69700 21854
rect 69666 21446 69700 21462
rect 69884 21838 69918 21854
rect 69884 21446 69918 21462
rect 70102 21838 70136 21854
rect 70102 21446 70136 21462
rect 70320 21838 70354 21854
rect 70320 21446 70354 21462
rect 70538 21838 70572 21854
rect 70538 21446 70572 21462
rect 70756 21838 70790 21854
rect 72656 21725 72672 21759
rect 73228 21725 73244 21759
rect 73674 21725 73690 21759
rect 74246 21725 74262 21759
rect 74692 21725 74708 21759
rect 75264 21725 75280 21759
rect 75710 21725 75726 21759
rect 76282 21725 76298 21759
rect 76728 21725 76744 21759
rect 77300 21725 77316 21759
rect 77746 21725 77762 21759
rect 78318 21725 78334 21759
rect 78764 21725 78780 21759
rect 79336 21725 79352 21759
rect 79782 21725 79798 21759
rect 80354 21725 80370 21759
rect 80800 21725 80816 21759
rect 81372 21725 81388 21759
rect 81818 21725 81834 21759
rect 82390 21725 82406 21759
rect 82836 21725 82852 21759
rect 83408 21725 83424 21759
rect 83854 21725 83870 21759
rect 84426 21725 84442 21759
rect 84872 21725 84888 21759
rect 85444 21725 85460 21759
rect 85890 21725 85906 21759
rect 86462 21725 86478 21759
rect 86908 21725 86924 21759
rect 87480 21725 87496 21759
rect 70756 21446 70790 21462
rect 72424 21666 72458 21682
rect 68894 21403 68954 21404
rect 68648 21369 68664 21403
rect 68740 21369 68756 21403
rect 68866 21369 68882 21403
rect 68958 21369 68974 21403
rect 69084 21369 69100 21403
rect 69176 21369 69192 21403
rect 69302 21369 69318 21403
rect 69394 21369 69410 21403
rect 69520 21369 69536 21403
rect 69612 21369 69628 21403
rect 69738 21369 69754 21403
rect 69830 21369 69846 21403
rect 69956 21369 69972 21403
rect 70048 21369 70064 21403
rect 70174 21369 70190 21403
rect 70266 21369 70282 21403
rect 70392 21369 70408 21403
rect 70484 21369 70500 21403
rect 70610 21369 70626 21403
rect 70702 21369 70718 21403
rect 68620 21190 68710 21220
rect 68620 21156 68648 21190
rect 68682 21156 68710 21190
rect 68620 21128 68710 21156
rect 69638 21190 69728 21220
rect 69638 21156 69666 21190
rect 69700 21156 69728 21190
rect 69638 21128 69728 21156
rect 70656 21190 70746 21220
rect 70656 21156 70684 21190
rect 70718 21156 70746 21190
rect 70656 21128 70746 21156
rect 72424 21074 72458 21090
rect 73442 21666 73476 21682
rect 73442 21074 73476 21090
rect 74460 21666 74494 21682
rect 74460 21074 74494 21090
rect 75478 21666 75512 21682
rect 75478 21074 75512 21090
rect 76496 21666 76530 21682
rect 76496 21074 76530 21090
rect 77514 21666 77548 21682
rect 77514 21074 77548 21090
rect 78532 21666 78566 21682
rect 78532 21074 78566 21090
rect 79550 21666 79584 21682
rect 79550 21074 79584 21090
rect 80568 21666 80602 21682
rect 80568 21074 80602 21090
rect 81586 21666 81620 21682
rect 81586 21074 81620 21090
rect 82604 21666 82638 21682
rect 82604 21074 82638 21090
rect 83622 21666 83656 21682
rect 83622 21074 83656 21090
rect 84640 21666 84674 21682
rect 84640 21074 84674 21090
rect 85658 21666 85692 21682
rect 85658 21074 85692 21090
rect 86676 21666 86710 21682
rect 86676 21074 86710 21090
rect 87694 21666 87728 21682
rect 87694 21074 87728 21090
rect 72656 20997 72672 21031
rect 73228 20997 73244 21031
rect 73674 20997 73690 21031
rect 74246 20997 74262 21031
rect 74692 20997 74708 21031
rect 75264 20997 75280 21031
rect 75710 20997 75726 21031
rect 76282 20997 76298 21031
rect 76728 20997 76744 21031
rect 77300 20997 77316 21031
rect 77746 20997 77762 21031
rect 78318 20997 78334 21031
rect 78764 20997 78780 21031
rect 79336 20997 79352 21031
rect 79782 20997 79798 21031
rect 80354 20997 80370 21031
rect 80800 20997 80816 21031
rect 81372 20997 81388 21031
rect 81818 20997 81834 21031
rect 82390 20997 82406 21031
rect 82836 20997 82852 21031
rect 83408 20997 83424 21031
rect 83854 20997 83870 21031
rect 84426 20997 84442 21031
rect 84872 20997 84888 21031
rect 85444 20997 85460 21031
rect 85890 20997 85906 21031
rect 86462 20997 86478 21031
rect 86908 20997 86924 21031
rect 87480 20997 87496 21031
rect 68648 20959 68664 20993
rect 68740 20959 68756 20993
rect 68866 20959 68882 20993
rect 68958 20959 68974 20993
rect 69084 20959 69100 20993
rect 69176 20959 69192 20993
rect 69302 20959 69318 20993
rect 69394 20959 69410 20993
rect 69520 20959 69536 20993
rect 69612 20959 69628 20993
rect 69738 20959 69754 20993
rect 69830 20959 69846 20993
rect 69956 20959 69972 20993
rect 70048 20959 70064 20993
rect 70174 20959 70190 20993
rect 70266 20959 70282 20993
rect 70392 20959 70408 20993
rect 70484 20959 70500 20993
rect 70610 20959 70626 20993
rect 70702 20959 70718 20993
rect 68576 20900 68610 20916
rect 68576 20508 68610 20524
rect 68794 20900 68828 20916
rect 68794 20508 68828 20524
rect 69012 20900 69046 20916
rect 69012 20508 69046 20524
rect 69230 20900 69264 20916
rect 69230 20508 69264 20524
rect 69448 20900 69482 20916
rect 69448 20508 69482 20524
rect 69666 20900 69700 20916
rect 69666 20508 69700 20524
rect 69884 20900 69918 20916
rect 69884 20508 69918 20524
rect 70102 20900 70136 20916
rect 70102 20508 70136 20524
rect 70320 20900 70354 20916
rect 70320 20508 70354 20524
rect 70538 20900 70572 20916
rect 70538 20508 70572 20524
rect 70756 20900 70790 20916
rect 72894 20766 72984 20796
rect 72894 20732 72922 20766
rect 72956 20732 72984 20766
rect 72894 20704 72984 20732
rect 73912 20766 74002 20796
rect 73912 20732 73940 20766
rect 73974 20732 74002 20766
rect 73912 20704 74002 20732
rect 74930 20766 75020 20796
rect 74930 20732 74958 20766
rect 74992 20732 75020 20766
rect 74930 20704 75020 20732
rect 75948 20766 76038 20796
rect 75948 20732 75976 20766
rect 76010 20732 76038 20766
rect 75948 20704 76038 20732
rect 76966 20766 77056 20796
rect 76966 20732 76994 20766
rect 77028 20732 77056 20766
rect 76966 20704 77056 20732
rect 77984 20766 78074 20796
rect 77984 20732 78012 20766
rect 78046 20732 78074 20766
rect 77984 20704 78074 20732
rect 79002 20766 79092 20796
rect 79002 20732 79030 20766
rect 79064 20732 79092 20766
rect 79002 20704 79092 20732
rect 80020 20766 80110 20796
rect 80020 20732 80048 20766
rect 80082 20732 80110 20766
rect 80020 20704 80110 20732
rect 81038 20766 81128 20796
rect 81038 20732 81066 20766
rect 81100 20732 81128 20766
rect 81038 20704 81128 20732
rect 82056 20766 82146 20796
rect 82056 20732 82084 20766
rect 82118 20732 82146 20766
rect 82056 20704 82146 20732
rect 83074 20766 83164 20796
rect 83074 20732 83102 20766
rect 83136 20732 83164 20766
rect 83074 20704 83164 20732
rect 84092 20766 84182 20796
rect 84092 20732 84120 20766
rect 84154 20732 84182 20766
rect 84092 20704 84182 20732
rect 85110 20766 85200 20796
rect 85110 20732 85138 20766
rect 85172 20732 85200 20766
rect 85110 20704 85200 20732
rect 86128 20766 86218 20796
rect 86128 20732 86156 20766
rect 86190 20732 86218 20766
rect 86128 20704 86218 20732
rect 87146 20766 87236 20796
rect 87146 20732 87174 20766
rect 87208 20732 87236 20766
rect 87146 20704 87236 20732
rect 70756 20508 70790 20524
rect 72656 20469 72672 20503
rect 73228 20469 73244 20503
rect 73674 20469 73690 20503
rect 74246 20469 74262 20503
rect 74692 20469 74708 20503
rect 75264 20469 75280 20503
rect 75710 20469 75726 20503
rect 76282 20469 76298 20503
rect 76728 20469 76744 20503
rect 77300 20469 77316 20503
rect 77746 20469 77762 20503
rect 78318 20469 78334 20503
rect 78764 20469 78780 20503
rect 79336 20469 79352 20503
rect 79782 20469 79798 20503
rect 80354 20469 80370 20503
rect 80800 20469 80816 20503
rect 81372 20469 81388 20503
rect 81818 20469 81834 20503
rect 82390 20469 82406 20503
rect 82836 20469 82852 20503
rect 83408 20469 83424 20503
rect 83854 20469 83870 20503
rect 84426 20469 84442 20503
rect 84872 20469 84888 20503
rect 85444 20469 85460 20503
rect 85890 20469 85906 20503
rect 86462 20469 86478 20503
rect 86908 20469 86924 20503
rect 87480 20469 87496 20503
rect 69326 20465 69386 20466
rect 70198 20465 70258 20466
rect 68648 20431 68664 20465
rect 68740 20431 68756 20465
rect 68866 20431 68882 20465
rect 68958 20431 68974 20465
rect 69084 20431 69100 20465
rect 69176 20431 69192 20465
rect 69302 20431 69318 20465
rect 69394 20431 69410 20465
rect 69520 20431 69536 20465
rect 69612 20431 69628 20465
rect 69738 20431 69754 20465
rect 69830 20431 69846 20465
rect 69956 20431 69972 20465
rect 70048 20431 70064 20465
rect 70174 20431 70190 20465
rect 70266 20431 70282 20465
rect 70392 20431 70408 20465
rect 70484 20431 70500 20465
rect 70610 20431 70626 20465
rect 70702 20431 70718 20465
rect 72424 20410 72458 20426
rect 68592 20248 68682 20278
rect 68592 20214 68620 20248
rect 68654 20214 68682 20248
rect 68592 20186 68682 20214
rect 69610 20248 69700 20278
rect 69610 20214 69638 20248
rect 69672 20214 69700 20248
rect 69610 20186 69700 20214
rect 70628 20248 70718 20278
rect 70628 20214 70656 20248
rect 70690 20214 70718 20248
rect 70628 20186 70718 20214
rect 68648 20021 68664 20055
rect 68740 20021 68756 20055
rect 68866 20021 68882 20055
rect 68958 20021 68974 20055
rect 69084 20021 69100 20055
rect 69176 20021 69192 20055
rect 69302 20021 69318 20055
rect 69394 20021 69410 20055
rect 69520 20021 69536 20055
rect 69612 20021 69628 20055
rect 69738 20021 69754 20055
rect 69830 20021 69846 20055
rect 69956 20021 69972 20055
rect 70048 20021 70064 20055
rect 70174 20021 70190 20055
rect 70266 20021 70282 20055
rect 70392 20021 70408 20055
rect 70484 20021 70500 20055
rect 70610 20021 70626 20055
rect 70702 20021 70718 20055
rect 68888 20020 68948 20021
rect 69326 20020 69386 20021
rect 68576 19962 68610 19978
rect 68576 19570 68610 19586
rect 68794 19962 68828 19978
rect 68794 19570 68828 19586
rect 69012 19962 69046 19978
rect 69012 19570 69046 19586
rect 69230 19962 69264 19978
rect 69230 19570 69264 19586
rect 69448 19962 69482 19978
rect 69448 19570 69482 19586
rect 69666 19962 69700 19978
rect 69666 19570 69700 19586
rect 69884 19962 69918 19978
rect 69884 19570 69918 19586
rect 70102 19962 70136 19978
rect 70102 19570 70136 19586
rect 70320 19962 70354 19978
rect 70320 19570 70354 19586
rect 70538 19962 70572 19978
rect 70538 19570 70572 19586
rect 70756 19962 70790 19978
rect 72424 19818 72458 19834
rect 73442 20410 73476 20426
rect 73442 19818 73476 19834
rect 74460 20410 74494 20426
rect 74460 19818 74494 19834
rect 75478 20410 75512 20426
rect 75478 19818 75512 19834
rect 76496 20410 76530 20426
rect 76496 19818 76530 19834
rect 77514 20410 77548 20426
rect 77514 19818 77548 19834
rect 78532 20410 78566 20426
rect 78532 19818 78566 19834
rect 79550 20410 79584 20426
rect 79550 19818 79584 19834
rect 80568 20410 80602 20426
rect 80568 19818 80602 19834
rect 81586 20410 81620 20426
rect 81586 19818 81620 19834
rect 82604 20410 82638 20426
rect 82604 19818 82638 19834
rect 83622 20410 83656 20426
rect 83622 19818 83656 19834
rect 84640 20410 84674 20426
rect 84640 19818 84674 19834
rect 85658 20410 85692 20426
rect 85658 19818 85692 19834
rect 86676 20410 86710 20426
rect 86676 19818 86710 19834
rect 87694 20410 87728 20426
rect 87694 19818 87728 19834
rect 72656 19741 72672 19775
rect 73228 19741 73244 19775
rect 73674 19741 73690 19775
rect 74246 19741 74262 19775
rect 74692 19741 74708 19775
rect 75264 19741 75280 19775
rect 75710 19741 75726 19775
rect 76282 19741 76298 19775
rect 76728 19741 76744 19775
rect 77300 19741 77316 19775
rect 77746 19741 77762 19775
rect 78318 19741 78334 19775
rect 78764 19741 78780 19775
rect 79336 19741 79352 19775
rect 79782 19741 79798 19775
rect 80354 19741 80370 19775
rect 80800 19741 80816 19775
rect 81372 19741 81388 19775
rect 81818 19741 81834 19775
rect 82390 19741 82406 19775
rect 82836 19741 82852 19775
rect 83408 19741 83424 19775
rect 83854 19741 83870 19775
rect 84426 19741 84442 19775
rect 84872 19741 84888 19775
rect 85444 19741 85460 19775
rect 85890 19741 85906 19775
rect 86462 19741 86478 19775
rect 86908 19741 86924 19775
rect 87480 19741 87496 19775
rect 70756 19570 70790 19586
rect 72894 19528 72984 19558
rect 68648 19493 68664 19527
rect 68740 19493 68756 19527
rect 68866 19493 68882 19527
rect 68958 19493 68974 19527
rect 69084 19493 69100 19527
rect 69176 19493 69192 19527
rect 69302 19493 69318 19527
rect 69394 19493 69410 19527
rect 69520 19493 69536 19527
rect 69612 19493 69628 19527
rect 69738 19493 69754 19527
rect 69830 19493 69846 19527
rect 69956 19493 69972 19527
rect 70048 19493 70064 19527
rect 70174 19493 70190 19527
rect 70266 19493 70282 19527
rect 70392 19493 70408 19527
rect 70484 19493 70500 19527
rect 70610 19493 70626 19527
rect 70702 19493 70718 19527
rect 72894 19494 72922 19528
rect 72956 19494 72984 19528
rect 72894 19466 72984 19494
rect 73912 19528 74002 19558
rect 73912 19494 73940 19528
rect 73974 19494 74002 19528
rect 73912 19466 74002 19494
rect 74930 19528 75020 19558
rect 74930 19494 74958 19528
rect 74992 19494 75020 19528
rect 74930 19466 75020 19494
rect 75948 19528 76038 19558
rect 75948 19494 75976 19528
rect 76010 19494 76038 19528
rect 75948 19466 76038 19494
rect 76966 19528 77056 19558
rect 76966 19494 76994 19528
rect 77028 19494 77056 19528
rect 76966 19466 77056 19494
rect 77984 19528 78074 19558
rect 77984 19494 78012 19528
rect 78046 19494 78074 19528
rect 77984 19466 78074 19494
rect 79002 19528 79092 19558
rect 79002 19494 79030 19528
rect 79064 19494 79092 19528
rect 79002 19466 79092 19494
rect 80020 19528 80110 19558
rect 80020 19494 80048 19528
rect 80082 19494 80110 19528
rect 80020 19466 80110 19494
rect 81038 19528 81128 19558
rect 81038 19494 81066 19528
rect 81100 19494 81128 19528
rect 81038 19466 81128 19494
rect 82056 19528 82146 19558
rect 82056 19494 82084 19528
rect 82118 19494 82146 19528
rect 82056 19466 82146 19494
rect 83074 19528 83164 19558
rect 83074 19494 83102 19528
rect 83136 19494 83164 19528
rect 83074 19466 83164 19494
rect 84092 19528 84182 19558
rect 84092 19494 84120 19528
rect 84154 19494 84182 19528
rect 84092 19466 84182 19494
rect 85110 19528 85200 19558
rect 85110 19494 85138 19528
rect 85172 19494 85200 19528
rect 85110 19466 85200 19494
rect 86128 19528 86218 19558
rect 86128 19494 86156 19528
rect 86190 19494 86218 19528
rect 86128 19466 86218 19494
rect 87146 19528 87236 19558
rect 87146 19494 87174 19528
rect 87208 19494 87236 19528
rect 87146 19466 87236 19494
rect 68592 19334 68682 19364
rect 68592 19300 68620 19334
rect 68654 19300 68682 19334
rect 68592 19272 68682 19300
rect 69610 19334 69700 19364
rect 69610 19300 69638 19334
rect 69672 19300 69700 19334
rect 69610 19272 69700 19300
rect 70628 19334 70718 19364
rect 70628 19300 70656 19334
rect 70690 19300 70718 19334
rect 70628 19272 70718 19300
rect 72656 19213 72672 19247
rect 73228 19213 73244 19247
rect 73674 19213 73690 19247
rect 74246 19213 74262 19247
rect 74692 19213 74708 19247
rect 75264 19213 75280 19247
rect 75710 19213 75726 19247
rect 76282 19213 76298 19247
rect 76728 19213 76744 19247
rect 77300 19213 77316 19247
rect 77746 19213 77762 19247
rect 78318 19213 78334 19247
rect 78764 19213 78780 19247
rect 79336 19213 79352 19247
rect 79782 19213 79798 19247
rect 80354 19213 80370 19247
rect 80800 19213 80816 19247
rect 81372 19213 81388 19247
rect 81818 19213 81834 19247
rect 82390 19213 82406 19247
rect 82836 19213 82852 19247
rect 83408 19213 83424 19247
rect 83854 19213 83870 19247
rect 84426 19213 84442 19247
rect 84872 19213 84888 19247
rect 85444 19213 85460 19247
rect 85890 19213 85906 19247
rect 86462 19213 86478 19247
rect 86908 19213 86924 19247
rect 87480 19213 87496 19247
rect 72424 19154 72458 19170
rect 68648 19083 68664 19117
rect 68740 19083 68756 19117
rect 68866 19083 68882 19117
rect 68958 19083 68974 19117
rect 69084 19083 69100 19117
rect 69176 19083 69192 19117
rect 69302 19083 69318 19117
rect 69394 19083 69410 19117
rect 69520 19083 69536 19117
rect 69612 19083 69628 19117
rect 69738 19083 69754 19117
rect 69830 19083 69846 19117
rect 69956 19083 69972 19117
rect 70048 19083 70064 19117
rect 70174 19083 70190 19117
rect 70266 19083 70282 19117
rect 70392 19083 70408 19117
rect 70484 19083 70500 19117
rect 70610 19083 70626 19117
rect 70702 19083 70718 19117
rect 69330 19082 69390 19083
rect 68576 19024 68610 19040
rect 68576 18632 68610 18648
rect 68794 19024 68828 19040
rect 68794 18632 68828 18648
rect 69012 19024 69046 19040
rect 69012 18632 69046 18648
rect 69230 19024 69264 19040
rect 69230 18632 69264 18648
rect 69448 19024 69482 19040
rect 69448 18632 69482 18648
rect 69666 19024 69700 19040
rect 69666 18632 69700 18648
rect 69884 19024 69918 19040
rect 69884 18632 69918 18648
rect 70102 19024 70136 19040
rect 70102 18632 70136 18648
rect 70320 19024 70354 19040
rect 70320 18632 70354 18648
rect 70538 19024 70572 19040
rect 70538 18632 70572 18648
rect 70756 19024 70790 19040
rect 70756 18632 70790 18648
rect 68648 18555 68664 18589
rect 68740 18555 68756 18589
rect 68866 18555 68882 18589
rect 68958 18555 68974 18589
rect 69084 18555 69100 18589
rect 69176 18555 69192 18589
rect 69302 18555 69318 18589
rect 69394 18555 69410 18589
rect 69520 18555 69536 18589
rect 69612 18555 69628 18589
rect 69738 18555 69754 18589
rect 69830 18555 69846 18589
rect 69956 18555 69972 18589
rect 70048 18555 70064 18589
rect 70174 18555 70190 18589
rect 70266 18555 70282 18589
rect 70392 18555 70408 18589
rect 70484 18555 70500 18589
rect 70610 18555 70626 18589
rect 70702 18555 70718 18589
rect 72424 18562 72458 18578
rect 73442 19154 73476 19170
rect 73442 18562 73476 18578
rect 74460 19154 74494 19170
rect 74460 18562 74494 18578
rect 75478 19154 75512 19170
rect 75478 18562 75512 18578
rect 76496 19154 76530 19170
rect 76496 18562 76530 18578
rect 77514 19154 77548 19170
rect 77514 18562 77548 18578
rect 78532 19154 78566 19170
rect 78532 18562 78566 18578
rect 79550 19154 79584 19170
rect 79550 18562 79584 18578
rect 80568 19154 80602 19170
rect 80568 18562 80602 18578
rect 81586 19154 81620 19170
rect 81586 18562 81620 18578
rect 82604 19154 82638 19170
rect 82604 18562 82638 18578
rect 83622 19154 83656 19170
rect 83622 18562 83656 18578
rect 84640 19154 84674 19170
rect 84640 18562 84674 18578
rect 85658 19154 85692 19170
rect 85658 18562 85692 18578
rect 86676 19154 86710 19170
rect 86676 18562 86710 18578
rect 87694 19154 87728 19170
rect 87694 18562 87728 18578
rect 72656 18485 72672 18519
rect 73228 18485 73244 18519
rect 73674 18485 73690 18519
rect 74246 18485 74262 18519
rect 74692 18485 74708 18519
rect 75264 18485 75280 18519
rect 75710 18485 75726 18519
rect 76282 18485 76298 18519
rect 76728 18485 76744 18519
rect 77300 18485 77316 18519
rect 77746 18485 77762 18519
rect 78318 18485 78334 18519
rect 78764 18485 78780 18519
rect 79336 18485 79352 18519
rect 79782 18485 79798 18519
rect 80354 18485 80370 18519
rect 80800 18485 80816 18519
rect 81372 18485 81388 18519
rect 81818 18485 81834 18519
rect 82390 18485 82406 18519
rect 82836 18485 82852 18519
rect 83408 18485 83424 18519
rect 83854 18485 83870 18519
rect 84426 18485 84442 18519
rect 84872 18485 84888 18519
rect 85444 18485 85460 18519
rect 85890 18485 85906 18519
rect 86462 18485 86478 18519
rect 86908 18485 86924 18519
rect 87480 18485 87496 18519
rect 65328 17658 65428 17820
rect 89672 17658 89772 17820
rect -13094 16248 -13048 16281
rect -11354 16248 -11284 16281
rect -13094 16247 -12998 16248
rect -11380 16247 -11284 16248
rect -13094 16185 -13060 16247
rect -11318 16186 -11284 16247
rect -12900 16145 -12884 16179
rect -12784 16145 -12768 16179
rect -12642 16145 -12626 16179
rect -12526 16145 -12510 16179
rect -12384 16145 -12368 16179
rect -12268 16145 -12252 16179
rect -12126 16145 -12110 16179
rect -12010 16145 -11994 16179
rect -11868 16145 -11852 16179
rect -11752 16145 -11736 16179
rect -11610 16145 -11594 16179
rect -11494 16145 -11478 16179
rect -12980 16086 -12946 16102
rect -12980 15694 -12946 15710
rect -12722 16086 -12688 16102
rect -12722 15694 -12688 15710
rect -12464 16086 -12430 16102
rect -12464 15694 -12430 15710
rect -12206 16086 -12172 16102
rect -12206 15694 -12172 15710
rect -11948 16086 -11914 16102
rect -11948 15694 -11914 15710
rect -11690 16086 -11656 16102
rect -11690 15694 -11656 15710
rect -11432 16086 -11398 16102
rect -11432 15694 -11398 15710
rect -12900 15617 -12884 15651
rect -12784 15617 -12768 15651
rect -12642 15617 -12626 15651
rect -12526 15617 -12510 15651
rect -12384 15617 -12368 15651
rect -12268 15617 -12252 15651
rect -12126 15617 -12110 15651
rect -12010 15617 -11994 15651
rect -11868 15617 -11852 15651
rect -11752 15617 -11736 15651
rect -11610 15617 -11594 15651
rect -11494 15617 -11478 15651
rect -13094 15549 -13060 15611
rect -10494 16248 -10448 16281
rect -8754 16248 -8684 16281
rect -10494 16247 -10398 16248
rect -8780 16247 -8684 16248
rect -10494 16185 -10460 16247
rect -8718 16186 -8684 16247
rect -11210 15745 -11181 15779
rect -11147 15745 -11089 15779
rect -11055 15745 -10997 15779
rect -10963 15745 -10934 15779
rect -11318 15549 -11284 15610
rect -13094 15548 -12998 15549
rect -13094 15515 -13048 15548
rect -11354 15516 -11284 15549
rect -11380 15515 -11284 15516
rect -11144 15703 -11078 15711
rect -11144 15669 -11128 15703
rect -11094 15669 -11078 15703
rect -11144 15635 -11078 15669
rect -11144 15601 -11128 15635
rect -11094 15601 -11078 15635
rect -11144 15567 -11078 15601
rect -11144 15533 -11128 15567
rect -11094 15533 -11078 15567
rect -11144 15515 -11078 15533
rect -11044 15703 -11002 15745
rect -11010 15669 -11002 15703
rect -11044 15635 -11002 15669
rect -11010 15601 -11002 15635
rect -10300 16145 -10284 16179
rect -10184 16145 -10168 16179
rect -10042 16145 -10026 16179
rect -9926 16145 -9910 16179
rect -9784 16145 -9768 16179
rect -9668 16145 -9652 16179
rect -9526 16145 -9510 16179
rect -9410 16145 -9394 16179
rect -9268 16145 -9252 16179
rect -9152 16145 -9136 16179
rect -9010 16145 -8994 16179
rect -8894 16145 -8878 16179
rect -10380 16086 -10346 16102
rect -10380 15694 -10346 15710
rect -10122 16086 -10088 16102
rect -10122 15694 -10088 15710
rect -9864 16086 -9830 16102
rect -9864 15694 -9830 15710
rect -9606 16086 -9572 16102
rect -9606 15694 -9572 15710
rect -9348 16086 -9314 16102
rect -9348 15694 -9314 15710
rect -9090 16086 -9056 16102
rect -9090 15694 -9056 15710
rect -8832 16086 -8798 16102
rect -8832 15694 -8798 15710
rect -10300 15617 -10284 15651
rect -10184 15617 -10168 15651
rect -10042 15617 -10026 15651
rect -9926 15617 -9910 15651
rect -9784 15617 -9768 15651
rect -9668 15617 -9652 15651
rect -9526 15617 -9510 15651
rect -9410 15617 -9394 15651
rect -9268 15617 -9252 15651
rect -9152 15617 -9136 15651
rect -9010 15617 -8994 15651
rect -8894 15617 -8878 15651
rect -11044 15567 -11002 15601
rect -11010 15533 -11002 15567
rect -11044 15517 -11002 15533
rect -10494 15549 -10460 15611
rect -8610 15745 -8581 15779
rect -8547 15745 -8489 15779
rect -8455 15745 -8397 15779
rect -8363 15745 -8334 15779
rect -8110 15745 -8081 15779
rect -8047 15745 -7989 15779
rect -7955 15745 -7897 15779
rect -7863 15745 -7834 15779
rect -8718 15549 -8684 15610
rect -10494 15548 -10398 15549
rect -10494 15515 -10448 15548
rect -8754 15516 -8684 15549
rect -8780 15515 -8684 15516
rect -8544 15703 -8478 15711
rect -8544 15669 -8528 15703
rect -8494 15669 -8478 15703
rect -8544 15635 -8478 15669
rect -8544 15601 -8528 15635
rect -8494 15601 -8478 15635
rect -8544 15567 -8478 15601
rect -8544 15533 -8528 15567
rect -8494 15533 -8478 15567
rect -8544 15515 -8478 15533
rect -8444 15703 -8402 15745
rect -8410 15669 -8402 15703
rect -8444 15635 -8402 15669
rect -8410 15601 -8402 15635
rect -8444 15567 -8402 15601
rect -8410 15533 -8402 15567
rect -8444 15517 -8402 15533
rect -8044 15703 -7978 15711
rect -8044 15669 -8028 15703
rect -7994 15669 -7978 15703
rect -8044 15635 -7978 15669
rect -8044 15601 -8028 15635
rect -7994 15601 -7978 15635
rect -8044 15567 -7978 15601
rect -8044 15533 -8028 15567
rect -7994 15533 -7978 15567
rect -8044 15515 -7978 15533
rect -7944 15703 -7902 15745
rect -7910 15669 -7902 15703
rect -7944 15635 -7902 15669
rect -7910 15601 -7902 15635
rect -7944 15567 -7902 15601
rect -7910 15533 -7902 15567
rect -7944 15517 -7902 15533
rect -11144 15456 -11098 15515
rect -11103 15408 -11098 15456
rect -11064 15478 -10998 15481
rect -11064 15467 -11047 15478
rect -11064 15433 -11048 15467
rect -11001 15438 -10998 15478
rect -8544 15456 -8498 15515
rect -11014 15433 -10998 15438
rect -8503 15408 -8498 15456
rect -8464 15478 -8398 15481
rect -8044 15478 -7998 15515
rect -8464 15467 -8447 15478
rect -8464 15433 -8448 15467
rect -8401 15438 -8398 15478
rect -8414 15433 -8398 15438
rect -8004 15430 -7998 15478
rect -7964 15434 -7950 15481
rect -7902 15434 -7898 15481
rect -7964 15433 -7948 15434
rect -7914 15433 -7898 15434
rect -11144 15395 -11098 15408
rect -11144 15383 -11078 15395
rect -11144 15349 -11128 15383
rect -11094 15349 -11078 15383
rect -13094 15314 -13024 15348
rect -11354 15314 -11284 15348
rect -13094 15252 -13060 15314
rect -11318 15252 -11284 15314
rect -11144 15315 -11078 15349
rect -11144 15281 -11128 15315
rect -11094 15281 -11078 15315
rect -11144 15269 -11078 15281
rect -11044 15383 -10998 15399
rect -11010 15349 -10998 15383
rect -8544 15395 -8498 15408
rect -8544 15383 -8478 15395
rect -11044 15315 -10998 15349
rect -8544 15349 -8528 15383
rect -8494 15349 -8478 15383
rect -11010 15281 -10998 15315
rect -12900 15212 -12884 15246
rect -12784 15212 -12768 15246
rect -12642 15212 -12626 15246
rect -12526 15212 -12510 15246
rect -12384 15212 -12368 15246
rect -12268 15212 -12252 15246
rect -12126 15212 -12110 15246
rect -12010 15212 -11994 15246
rect -11868 15212 -11852 15246
rect -11752 15212 -11736 15246
rect -11610 15212 -11594 15246
rect -11494 15212 -11478 15246
rect -12980 15162 -12946 15178
rect -12980 14970 -12946 14986
rect -12722 15162 -12688 15178
rect -12722 14970 -12688 14986
rect -12464 15162 -12430 15178
rect -12464 14970 -12430 14986
rect -12206 15162 -12172 15178
rect -12206 14970 -12172 14986
rect -11948 15162 -11914 15178
rect -11948 14970 -11914 14986
rect -11690 15162 -11656 15178
rect -11690 14970 -11656 14986
rect -11432 15162 -11398 15178
rect -11432 14970 -11398 14986
rect -12900 14902 -12884 14936
rect -12784 14902 -12768 14936
rect -12642 14902 -12626 14936
rect -12526 14902 -12510 14936
rect -12384 14902 -12368 14936
rect -12268 14902 -12252 14936
rect -12126 14902 -12110 14936
rect -12010 14902 -11994 14936
rect -11868 14902 -11852 14936
rect -11752 14902 -11736 14936
rect -11610 14902 -11594 14936
rect -11494 14902 -11478 14936
rect -11044 15235 -10998 15281
rect -10494 15314 -10424 15348
rect -8754 15314 -8684 15348
rect -10494 15252 -10460 15314
rect -8718 15252 -8684 15314
rect -8544 15315 -8478 15349
rect -8544 15281 -8528 15315
rect -8494 15281 -8478 15315
rect -8544 15269 -8478 15281
rect -8444 15383 -8398 15399
rect -8410 15349 -8398 15383
rect -8444 15315 -8398 15349
rect -8410 15281 -8398 15315
rect -11210 15201 -11181 15235
rect -11147 15201 -11089 15235
rect -11055 15201 -10997 15235
rect -10963 15201 -10934 15235
rect -10300 15212 -10284 15246
rect -10184 15212 -10168 15246
rect -10042 15212 -10026 15246
rect -9926 15212 -9910 15246
rect -9784 15212 -9768 15246
rect -9668 15212 -9652 15246
rect -9526 15212 -9510 15246
rect -9410 15212 -9394 15246
rect -9268 15212 -9252 15246
rect -9152 15212 -9136 15246
rect -9010 15212 -8994 15246
rect -8894 15212 -8878 15246
rect -10380 15162 -10346 15178
rect -10380 14970 -10346 14986
rect -10122 15162 -10088 15178
rect -10122 14970 -10088 14986
rect -9864 15162 -9830 15178
rect -9864 14970 -9830 14986
rect -9606 15162 -9572 15178
rect -9606 14970 -9572 14986
rect -9348 15162 -9314 15178
rect -9348 14970 -9314 14986
rect -9090 15162 -9056 15178
rect -9090 14970 -9056 14986
rect -8832 15162 -8798 15178
rect -8832 14970 -8798 14986
rect -10300 14902 -10284 14936
rect -10184 14902 -10168 14936
rect -10042 14902 -10026 14936
rect -9926 14902 -9910 14936
rect -9784 14902 -9768 14936
rect -9668 14902 -9652 14936
rect -9526 14902 -9510 14936
rect -9410 14902 -9394 14936
rect -9268 14902 -9252 14936
rect -9152 14902 -9136 14936
rect -9010 14902 -8994 14936
rect -8894 14902 -8878 14936
rect -8444 15235 -8398 15281
rect -8044 15395 -7998 15430
rect -8044 15383 -7978 15395
rect -8044 15349 -8028 15383
rect -7994 15349 -7978 15383
rect -8044 15315 -7978 15349
rect -8044 15281 -8028 15315
rect -7994 15281 -7978 15315
rect -8044 15269 -7978 15281
rect -7944 15383 -7898 15399
rect -7910 15349 -7898 15383
rect -7944 15315 -7898 15349
rect -7910 15281 -7898 15315
rect -7944 15235 -7898 15281
rect -8610 15201 -8581 15235
rect -8547 15201 -8489 15235
rect -8455 15201 -8397 15235
rect -8363 15201 -8334 15235
rect -8110 15201 -8081 15235
rect -8047 15201 -7989 15235
rect -7955 15201 -7897 15235
rect -7863 15201 -7834 15235
rect -1372 15200 -1272 15362
rect -13094 14834 -13060 14896
rect -11318 14834 -11284 14896
rect -13094 14800 -13026 14834
rect -11352 14800 -11284 14834
rect -10494 14834 -10460 14896
rect -8718 14834 -8684 14896
rect -10494 14800 -10426 14834
rect -8752 14800 -8684 14834
rect 35772 15200 35872 15362
rect 13764 14860 13780 14894
rect 14336 14860 14352 14894
rect 14782 14860 14798 14894
rect 15354 14860 15370 14894
rect 15800 14860 15816 14894
rect 16372 14860 16388 14894
rect 16818 14860 16834 14894
rect 17390 14860 17406 14894
rect 17836 14860 17852 14894
rect 18408 14860 18424 14894
rect 18854 14860 18870 14894
rect 19426 14860 19442 14894
rect 19872 14860 19888 14894
rect 20444 14860 20460 14894
rect 20890 14860 20906 14894
rect 21462 14860 21478 14894
rect 21908 14860 21924 14894
rect 22480 14860 22496 14894
rect 22926 14860 22942 14894
rect 23498 14860 23514 14894
rect 23944 14860 23960 14894
rect 24516 14860 24532 14894
rect 24962 14860 24978 14894
rect 25534 14860 25550 14894
rect 25980 14860 25996 14894
rect 26552 14860 26568 14894
rect 26998 14860 27014 14894
rect 27570 14860 27586 14894
rect 28016 14860 28032 14894
rect 28588 14860 28604 14894
rect 29034 14860 29050 14894
rect 29606 14860 29622 14894
rect 30052 14860 30068 14894
rect 30624 14860 30640 14894
rect 31070 14860 31086 14894
rect 31642 14860 31658 14894
rect 32088 14860 32104 14894
rect 32660 14860 32676 14894
rect 33106 14860 33122 14894
rect 33678 14860 33694 14894
rect 13532 14810 13566 14826
rect 2282 14318 2364 14342
rect 2282 14284 2306 14318
rect 2340 14284 2364 14318
rect 2282 14260 2364 14284
rect 3300 14318 3382 14342
rect 3300 14284 3324 14318
rect 3358 14284 3382 14318
rect 3300 14260 3382 14284
rect 4318 14318 4400 14342
rect 4318 14284 4342 14318
rect 4376 14284 4400 14318
rect 4318 14260 4400 14284
rect 5336 14318 5418 14342
rect 5336 14284 5360 14318
rect 5394 14284 5418 14318
rect 5336 14260 5418 14284
rect 6354 14318 6436 14342
rect 6354 14284 6378 14318
rect 6412 14284 6436 14318
rect 6354 14260 6436 14284
rect 7372 14318 7454 14342
rect 7372 14284 7396 14318
rect 7430 14284 7454 14318
rect 7372 14260 7454 14284
rect 8390 14318 8472 14342
rect 8390 14284 8414 14318
rect 8448 14284 8472 14318
rect 8390 14260 8472 14284
rect 9408 14318 9490 14342
rect 9408 14284 9432 14318
rect 9466 14284 9490 14318
rect 9408 14260 9490 14284
rect 10426 14318 10508 14342
rect 10426 14284 10450 14318
rect 10484 14284 10508 14318
rect 10426 14260 10508 14284
rect 13532 14218 13566 14234
rect 14550 14810 14584 14826
rect 14550 14218 14584 14234
rect 15568 14810 15602 14826
rect 15568 14218 15602 14234
rect 16586 14810 16620 14826
rect 16586 14218 16620 14234
rect 17604 14810 17638 14826
rect 17604 14218 17638 14234
rect 18622 14810 18656 14826
rect 18622 14218 18656 14234
rect 19640 14810 19674 14826
rect 19640 14218 19674 14234
rect 20658 14810 20692 14826
rect 20658 14218 20692 14234
rect 21676 14810 21710 14826
rect 21676 14218 21710 14234
rect 22694 14810 22728 14826
rect 22694 14218 22728 14234
rect 23712 14810 23746 14826
rect 23712 14218 23746 14234
rect 24730 14810 24764 14826
rect 24730 14218 24764 14234
rect 25748 14810 25782 14826
rect 25748 14218 25782 14234
rect 26766 14810 26800 14826
rect 26766 14218 26800 14234
rect 27784 14810 27818 14826
rect 27784 14218 27818 14234
rect 28802 14810 28836 14826
rect 28802 14218 28836 14234
rect 29820 14810 29854 14826
rect 29820 14218 29854 14234
rect 30838 14810 30872 14826
rect 30838 14218 30872 14234
rect 31856 14810 31890 14826
rect 31856 14218 31890 14234
rect 32874 14810 32908 14826
rect 32874 14218 32908 14234
rect 33892 14810 33926 14826
rect 33892 14218 33926 14234
rect 15050 14184 15110 14186
rect 16064 14184 16124 14192
rect 17068 14184 17128 14198
rect 18094 14184 18154 14186
rect 19118 14184 19178 14192
rect 20138 14184 20198 14186
rect 22164 14184 22224 14192
rect 23188 14184 23248 14186
rect 24198 14184 24258 14186
rect 25218 14184 25278 14192
rect 26248 14184 26308 14186
rect 27252 14184 27312 14192
rect 28268 14184 28328 14192
rect 29298 14184 29358 14186
rect 30312 14184 30372 14186
rect 31328 14184 31388 14186
rect 32354 14184 32414 14186
rect 33376 14184 33436 14186
rect 13764 14150 13780 14184
rect 14336 14150 14352 14184
rect 14782 14150 14798 14184
rect 15354 14150 15370 14184
rect 15800 14150 15816 14184
rect 16372 14150 16388 14184
rect 16818 14150 16834 14184
rect 17390 14150 17406 14184
rect 17836 14150 17852 14184
rect 18408 14150 18424 14184
rect 18854 14150 18870 14184
rect 19426 14150 19442 14184
rect 19872 14150 19888 14184
rect 20444 14150 20460 14184
rect 20890 14150 20906 14184
rect 21462 14150 21478 14184
rect 21908 14150 21924 14184
rect 22480 14150 22496 14184
rect 22926 14150 22942 14184
rect 23498 14150 23514 14184
rect 23944 14150 23960 14184
rect 24516 14150 24532 14184
rect 24962 14150 24978 14184
rect 25534 14150 25550 14184
rect 25980 14150 25996 14184
rect 26552 14150 26568 14184
rect 26998 14150 27014 14184
rect 27570 14150 27586 14184
rect 28016 14150 28032 14184
rect 28588 14150 28604 14184
rect 29034 14150 29050 14184
rect 29606 14150 29622 14184
rect 30052 14150 30068 14184
rect 30624 14150 30640 14184
rect 31070 14150 31086 14184
rect 31642 14150 31658 14184
rect 32088 14150 32104 14184
rect 32660 14150 32676 14184
rect 33106 14150 33122 14184
rect 33678 14150 33694 14184
rect 1998 14066 2014 14100
rect 2570 14066 2586 14100
rect 3016 14066 3032 14100
rect 3588 14066 3604 14100
rect 4034 14066 4050 14100
rect 4606 14066 4622 14100
rect 5052 14066 5068 14100
rect 5624 14066 5640 14100
rect 6070 14066 6086 14100
rect 6642 14066 6658 14100
rect 7088 14066 7104 14100
rect 7660 14066 7676 14100
rect 8106 14066 8122 14100
rect 8678 14066 8694 14100
rect 9124 14066 9140 14100
rect 9696 14066 9712 14100
rect 10142 14066 10158 14100
rect 10714 14066 10730 14100
rect 1766 14016 1800 14032
rect 1766 13424 1800 13440
rect 2784 14016 2818 14032
rect 2784 13424 2818 13440
rect 3802 14016 3836 14032
rect 3802 13424 3836 13440
rect 4820 14016 4854 14032
rect 4820 13424 4854 13440
rect 5838 14016 5872 14032
rect 5838 13424 5872 13440
rect 6856 14016 6890 14032
rect 6856 13424 6890 13440
rect 7874 14016 7908 14032
rect 7874 13424 7908 13440
rect 8892 14016 8926 14032
rect 8892 13424 8926 13440
rect 9910 14016 9944 14032
rect 9910 13424 9944 13440
rect 10928 14016 10962 14032
rect 14016 13926 14098 13950
rect 14016 13892 14040 13926
rect 14074 13892 14098 13926
rect 14016 13868 14098 13892
rect 15034 13926 15116 13950
rect 15034 13892 15058 13926
rect 15092 13892 15116 13926
rect 15034 13868 15116 13892
rect 16052 13926 16134 13950
rect 16052 13892 16076 13926
rect 16110 13892 16134 13926
rect 16052 13868 16134 13892
rect 17070 13926 17152 13950
rect 17070 13892 17094 13926
rect 17128 13892 17152 13926
rect 17070 13868 17152 13892
rect 18088 13926 18170 13950
rect 18088 13892 18112 13926
rect 18146 13892 18170 13926
rect 18088 13868 18170 13892
rect 19106 13926 19188 13950
rect 19106 13892 19130 13926
rect 19164 13892 19188 13926
rect 19106 13868 19188 13892
rect 20124 13926 20206 13950
rect 20124 13892 20148 13926
rect 20182 13892 20206 13926
rect 20124 13868 20206 13892
rect 21142 13926 21224 13950
rect 21142 13892 21166 13926
rect 21200 13892 21224 13926
rect 21142 13868 21224 13892
rect 22160 13926 22242 13950
rect 22160 13892 22184 13926
rect 22218 13892 22242 13926
rect 22160 13868 22242 13892
rect 23178 13926 23260 13950
rect 23178 13892 23202 13926
rect 23236 13892 23260 13926
rect 23178 13868 23260 13892
rect 24196 13926 24278 13950
rect 24196 13892 24220 13926
rect 24254 13892 24278 13926
rect 24196 13868 24278 13892
rect 25214 13926 25296 13950
rect 25214 13892 25238 13926
rect 25272 13892 25296 13926
rect 25214 13868 25296 13892
rect 26232 13926 26314 13950
rect 26232 13892 26256 13926
rect 26290 13892 26314 13926
rect 26232 13868 26314 13892
rect 27250 13926 27332 13950
rect 27250 13892 27274 13926
rect 27308 13892 27332 13926
rect 27250 13868 27332 13892
rect 28268 13926 28350 13950
rect 28268 13892 28292 13926
rect 28326 13892 28350 13926
rect 28268 13868 28350 13892
rect 29286 13926 29368 13950
rect 29286 13892 29310 13926
rect 29344 13892 29368 13926
rect 29286 13868 29368 13892
rect 30304 13926 30386 13950
rect 30304 13892 30328 13926
rect 30362 13892 30386 13926
rect 30304 13868 30386 13892
rect 31322 13926 31404 13950
rect 31322 13892 31346 13926
rect 31380 13892 31404 13926
rect 31322 13868 31404 13892
rect 32340 13926 32422 13950
rect 32340 13892 32364 13926
rect 32398 13892 32422 13926
rect 32340 13868 32422 13892
rect 33358 13926 33440 13950
rect 33358 13892 33382 13926
rect 33416 13892 33440 13926
rect 33358 13868 33440 13892
rect 13764 13626 13780 13660
rect 14336 13626 14352 13660
rect 14782 13626 14798 13660
rect 15354 13626 15370 13660
rect 15800 13626 15816 13660
rect 16372 13626 16388 13660
rect 16818 13626 16834 13660
rect 17390 13626 17406 13660
rect 17836 13626 17852 13660
rect 18408 13626 18424 13660
rect 18854 13626 18870 13660
rect 19426 13626 19442 13660
rect 19872 13626 19888 13660
rect 20444 13626 20460 13660
rect 20890 13626 20906 13660
rect 21462 13626 21478 13660
rect 21908 13626 21924 13660
rect 22480 13626 22496 13660
rect 22926 13626 22942 13660
rect 23498 13626 23514 13660
rect 23944 13626 23960 13660
rect 24516 13626 24532 13660
rect 24962 13626 24978 13660
rect 25534 13626 25550 13660
rect 25980 13626 25996 13660
rect 26552 13626 26568 13660
rect 26998 13626 27014 13660
rect 27570 13626 27586 13660
rect 28016 13626 28032 13660
rect 28588 13626 28604 13660
rect 29034 13626 29050 13660
rect 29606 13626 29622 13660
rect 30052 13626 30068 13660
rect 30624 13626 30640 13660
rect 31070 13626 31086 13660
rect 31642 13626 31658 13660
rect 32088 13626 32104 13660
rect 32660 13626 32676 13660
rect 33106 13626 33122 13660
rect 33678 13626 33694 13660
rect 23188 13620 23248 13626
rect 10928 13424 10962 13440
rect 13532 13576 13566 13592
rect 1744 13336 1826 13360
rect 1998 13356 2014 13390
rect 2570 13356 2586 13390
rect 1744 13302 1768 13336
rect 1802 13302 1826 13336
rect 1744 13278 1826 13302
rect 2762 13336 2844 13360
rect 3016 13356 3032 13390
rect 3588 13356 3604 13390
rect 2762 13302 2786 13336
rect 2820 13302 2844 13336
rect 1998 13248 2014 13282
rect 2570 13248 2586 13282
rect 2762 13278 2844 13302
rect 3780 13336 3862 13360
rect 4034 13356 4050 13390
rect 4606 13356 4622 13390
rect 3780 13302 3804 13336
rect 3838 13302 3862 13336
rect 3016 13248 3032 13282
rect 3588 13248 3604 13282
rect 3780 13278 3862 13302
rect 4798 13336 4880 13360
rect 5052 13356 5068 13390
rect 5624 13356 5640 13390
rect 4798 13302 4822 13336
rect 4856 13302 4880 13336
rect 4034 13248 4050 13282
rect 4606 13248 4622 13282
rect 4798 13278 4880 13302
rect 5816 13336 5898 13360
rect 6070 13356 6086 13390
rect 6642 13356 6658 13390
rect 5816 13302 5840 13336
rect 5874 13302 5898 13336
rect 5052 13248 5068 13282
rect 5624 13248 5640 13282
rect 5816 13278 5898 13302
rect 6834 13336 6916 13360
rect 7088 13356 7104 13390
rect 7660 13356 7676 13390
rect 6834 13302 6858 13336
rect 6892 13302 6916 13336
rect 6070 13248 6086 13282
rect 6642 13248 6658 13282
rect 6834 13278 6916 13302
rect 7852 13336 7934 13360
rect 8106 13356 8122 13390
rect 8678 13356 8694 13390
rect 7852 13302 7876 13336
rect 7910 13302 7934 13336
rect 7088 13248 7104 13282
rect 7660 13248 7676 13282
rect 7852 13278 7934 13302
rect 8870 13336 8952 13360
rect 9124 13356 9140 13390
rect 9696 13356 9712 13390
rect 8870 13302 8894 13336
rect 8928 13302 8952 13336
rect 8106 13248 8122 13282
rect 8678 13248 8694 13282
rect 8870 13278 8952 13302
rect 9888 13336 9970 13360
rect 10142 13356 10158 13390
rect 10714 13356 10730 13390
rect 9888 13302 9912 13336
rect 9946 13302 9970 13336
rect 9124 13248 9140 13282
rect 9696 13248 9712 13282
rect 9888 13278 9970 13302
rect 10906 13336 10988 13360
rect 10906 13302 10930 13336
rect 10964 13302 10988 13336
rect 10142 13248 10158 13282
rect 10714 13248 10730 13282
rect 10906 13278 10988 13302
rect 7358 13246 7418 13248
rect 1766 13198 1800 13214
rect 1766 12606 1800 12622
rect 2784 13198 2818 13214
rect 2784 12606 2818 12622
rect 3802 13198 3836 13214
rect 3802 12606 3836 12622
rect 4820 13198 4854 13214
rect 4820 12606 4854 12622
rect 5838 13198 5872 13214
rect 5838 12606 5872 12622
rect 6856 13198 6890 13214
rect 6856 12606 6890 12622
rect 7874 13198 7908 13214
rect 7874 12606 7908 12622
rect 8892 13198 8926 13214
rect 8892 12606 8926 12622
rect 9910 13198 9944 13214
rect 9910 12606 9944 12622
rect 10928 13198 10962 13214
rect 13532 12984 13566 13000
rect 14550 13576 14584 13592
rect 14550 12984 14584 13000
rect 15568 13576 15602 13592
rect 15568 12984 15602 13000
rect 16586 13576 16620 13592
rect 16586 12984 16620 13000
rect 17604 13576 17638 13592
rect 17604 12984 17638 13000
rect 18622 13576 18656 13592
rect 18622 12984 18656 13000
rect 19640 13576 19674 13592
rect 19640 12984 19674 13000
rect 20658 13576 20692 13592
rect 20658 12984 20692 13000
rect 21676 13576 21710 13592
rect 21676 12984 21710 13000
rect 22694 13576 22728 13592
rect 22694 12984 22728 13000
rect 23712 13576 23746 13592
rect 23712 12984 23746 13000
rect 24730 13576 24764 13592
rect 24730 12984 24764 13000
rect 25748 13576 25782 13592
rect 25748 12984 25782 13000
rect 26766 13576 26800 13592
rect 26766 12984 26800 13000
rect 27784 13576 27818 13592
rect 27784 12984 27818 13000
rect 28802 13576 28836 13592
rect 28802 12984 28836 13000
rect 29820 13576 29854 13592
rect 29820 12984 29854 13000
rect 30838 13576 30872 13592
rect 30838 12984 30872 13000
rect 31856 13576 31890 13592
rect 31856 12984 31890 13000
rect 32874 13576 32908 13592
rect 32874 12984 32908 13000
rect 33892 13576 33926 13592
rect 33892 12984 33926 13000
rect 19116 12950 19176 12956
rect 21152 12950 21212 12956
rect 22172 12950 22232 12956
rect 27244 12950 27304 12956
rect 13764 12916 13780 12950
rect 14336 12916 14352 12950
rect 14782 12916 14798 12950
rect 15354 12916 15370 12950
rect 15800 12916 15816 12950
rect 16372 12916 16388 12950
rect 16818 12916 16834 12950
rect 17390 12916 17406 12950
rect 17836 12916 17852 12950
rect 18408 12916 18424 12950
rect 18854 12916 18870 12950
rect 19426 12916 19442 12950
rect 19872 12916 19888 12950
rect 20444 12916 20460 12950
rect 20890 12916 20906 12950
rect 21462 12916 21478 12950
rect 21908 12916 21924 12950
rect 22480 12916 22496 12950
rect 22926 12916 22942 12950
rect 23498 12916 23514 12950
rect 23944 12916 23960 12950
rect 24516 12916 24532 12950
rect 24962 12916 24978 12950
rect 25534 12916 25550 12950
rect 25980 12916 25996 12950
rect 26552 12916 26568 12950
rect 26998 12916 27014 12950
rect 27570 12916 27586 12950
rect 28016 12916 28032 12950
rect 28588 12916 28604 12950
rect 29034 12916 29050 12950
rect 29606 12916 29622 12950
rect 30052 12916 30068 12950
rect 30624 12916 30640 12950
rect 31070 12916 31086 12950
rect 31642 12916 31658 12950
rect 32088 12916 32104 12950
rect 32660 12916 32676 12950
rect 33106 12916 33122 12950
rect 33678 12916 33694 12950
rect 14004 12690 14086 12714
rect 14004 12656 14028 12690
rect 14062 12656 14086 12690
rect 14004 12632 14086 12656
rect 15022 12690 15104 12714
rect 15022 12656 15046 12690
rect 15080 12656 15104 12690
rect 15022 12632 15104 12656
rect 16040 12690 16122 12714
rect 16040 12656 16064 12690
rect 16098 12656 16122 12690
rect 16040 12632 16122 12656
rect 17058 12690 17140 12714
rect 17058 12656 17082 12690
rect 17116 12656 17140 12690
rect 17058 12632 17140 12656
rect 18076 12690 18158 12714
rect 18076 12656 18100 12690
rect 18134 12656 18158 12690
rect 18076 12632 18158 12656
rect 19094 12690 19176 12714
rect 19094 12656 19118 12690
rect 19152 12656 19176 12690
rect 19094 12632 19176 12656
rect 20112 12690 20194 12714
rect 20112 12656 20136 12690
rect 20170 12656 20194 12690
rect 20112 12632 20194 12656
rect 21130 12690 21212 12714
rect 21130 12656 21154 12690
rect 21188 12656 21212 12690
rect 21130 12632 21212 12656
rect 22148 12690 22230 12714
rect 22148 12656 22172 12690
rect 22206 12656 22230 12690
rect 22148 12632 22230 12656
rect 23166 12690 23248 12714
rect 23166 12656 23190 12690
rect 23224 12656 23248 12690
rect 23166 12632 23248 12656
rect 24184 12690 24266 12714
rect 24184 12656 24208 12690
rect 24242 12656 24266 12690
rect 24184 12632 24266 12656
rect 25202 12690 25284 12714
rect 25202 12656 25226 12690
rect 25260 12656 25284 12690
rect 25202 12632 25284 12656
rect 26220 12690 26302 12714
rect 26220 12656 26244 12690
rect 26278 12656 26302 12690
rect 26220 12632 26302 12656
rect 27238 12690 27320 12714
rect 27238 12656 27262 12690
rect 27296 12656 27320 12690
rect 27238 12632 27320 12656
rect 28256 12690 28338 12714
rect 28256 12656 28280 12690
rect 28314 12656 28338 12690
rect 28256 12632 28338 12656
rect 29274 12690 29356 12714
rect 29274 12656 29298 12690
rect 29332 12656 29356 12690
rect 29274 12632 29356 12656
rect 30292 12690 30374 12714
rect 30292 12656 30316 12690
rect 30350 12656 30374 12690
rect 30292 12632 30374 12656
rect 31310 12690 31392 12714
rect 31310 12656 31334 12690
rect 31368 12656 31392 12690
rect 31310 12632 31392 12656
rect 32328 12690 32410 12714
rect 32328 12656 32352 12690
rect 32386 12656 32410 12690
rect 32328 12632 32410 12656
rect 33346 12690 33428 12714
rect 33346 12656 33370 12690
rect 33404 12656 33428 12690
rect 33346 12632 33428 12656
rect 10928 12606 10962 12622
rect 3290 12572 3350 12574
rect 4304 12572 4364 12574
rect 8378 12572 8438 12574
rect 9394 12572 9454 12574
rect 1744 12518 1826 12542
rect 1998 12538 2014 12572
rect 2570 12538 2586 12572
rect 1744 12484 1768 12518
rect 1802 12484 1826 12518
rect 1744 12460 1826 12484
rect 2762 12518 2844 12542
rect 3016 12538 3032 12572
rect 3588 12538 3604 12572
rect 2762 12484 2786 12518
rect 2820 12484 2844 12518
rect 1998 12430 2014 12464
rect 2570 12430 2586 12464
rect 2762 12460 2844 12484
rect 3780 12518 3862 12542
rect 4034 12538 4050 12572
rect 4606 12538 4622 12572
rect 3780 12484 3804 12518
rect 3838 12484 3862 12518
rect 3016 12430 3032 12464
rect 3588 12430 3604 12464
rect 3780 12460 3862 12484
rect 4798 12518 4880 12542
rect 5052 12538 5068 12572
rect 5624 12538 5640 12572
rect 4798 12484 4822 12518
rect 4856 12484 4880 12518
rect 4034 12430 4050 12464
rect 4606 12430 4622 12464
rect 4798 12460 4880 12484
rect 5816 12518 5898 12542
rect 6070 12538 6086 12572
rect 6642 12538 6658 12572
rect 5816 12484 5840 12518
rect 5874 12484 5898 12518
rect 5052 12430 5068 12464
rect 5624 12430 5640 12464
rect 5816 12460 5898 12484
rect 6834 12518 6916 12542
rect 7088 12538 7104 12572
rect 7660 12538 7676 12572
rect 6834 12484 6858 12518
rect 6892 12484 6916 12518
rect 6070 12430 6086 12464
rect 6642 12430 6658 12464
rect 6834 12460 6916 12484
rect 7852 12518 7934 12542
rect 8106 12538 8122 12572
rect 8678 12538 8694 12572
rect 7852 12484 7876 12518
rect 7910 12484 7934 12518
rect 7088 12430 7104 12464
rect 7660 12430 7676 12464
rect 7852 12460 7934 12484
rect 8870 12518 8952 12542
rect 9124 12538 9140 12572
rect 9696 12538 9712 12572
rect 8870 12484 8894 12518
rect 8928 12484 8952 12518
rect 8106 12430 8122 12464
rect 8678 12430 8694 12464
rect 8870 12460 8952 12484
rect 9888 12518 9970 12542
rect 10142 12538 10158 12572
rect 10714 12538 10730 12572
rect 9888 12484 9912 12518
rect 9946 12484 9970 12518
rect 9124 12430 9140 12464
rect 9696 12430 9712 12464
rect 9888 12460 9970 12484
rect 10906 12518 10988 12542
rect 10906 12484 10930 12518
rect 10964 12484 10988 12518
rect 10142 12430 10158 12464
rect 10714 12430 10730 12464
rect 10906 12460 10988 12484
rect 1766 12380 1800 12396
rect 1766 11788 1800 11804
rect 2784 12380 2818 12396
rect 2784 11788 2818 11804
rect 3802 12380 3836 12396
rect 3802 11788 3836 11804
rect 4820 12380 4854 12396
rect 4820 11788 4854 11804
rect 5838 12380 5872 12396
rect 5838 11788 5872 11804
rect 6856 12380 6890 12396
rect 6856 11788 6890 11804
rect 7874 12380 7908 12396
rect 7874 11788 7908 11804
rect 8892 12380 8926 12396
rect 8892 11788 8926 11804
rect 9910 12380 9944 12396
rect 9910 11788 9944 11804
rect 10928 12380 10962 12396
rect 13764 12394 13780 12428
rect 14336 12394 14352 12428
rect 14782 12394 14798 12428
rect 15354 12394 15370 12428
rect 15800 12394 15816 12428
rect 16372 12394 16388 12428
rect 16818 12394 16834 12428
rect 17390 12394 17406 12428
rect 17836 12394 17852 12428
rect 18408 12394 18424 12428
rect 18854 12394 18870 12428
rect 19426 12394 19442 12428
rect 19872 12394 19888 12428
rect 20444 12394 20460 12428
rect 20890 12394 20906 12428
rect 21462 12394 21478 12428
rect 21908 12394 21924 12428
rect 22480 12394 22496 12428
rect 22926 12394 22942 12428
rect 23498 12394 23514 12428
rect 23944 12394 23960 12428
rect 24516 12394 24532 12428
rect 24962 12394 24978 12428
rect 25534 12394 25550 12428
rect 25980 12394 25996 12428
rect 26552 12394 26568 12428
rect 26998 12394 27014 12428
rect 27570 12394 27586 12428
rect 28016 12394 28032 12428
rect 28588 12394 28604 12428
rect 29034 12394 29050 12428
rect 29606 12394 29622 12428
rect 30052 12394 30068 12428
rect 30624 12394 30640 12428
rect 31070 12394 31086 12428
rect 31642 12394 31658 12428
rect 32088 12394 32104 12428
rect 32660 12394 32676 12428
rect 33106 12394 33122 12428
rect 33678 12394 33694 12428
rect 15050 12390 15110 12394
rect 16066 12390 16126 12394
rect 20142 12386 20202 12394
rect 24208 12390 24268 12394
rect 26242 12390 26302 12394
rect 32354 12390 32414 12394
rect 10928 11788 10962 11804
rect 13532 12344 13566 12360
rect 3294 11754 3354 11756
rect 4308 11754 4368 11756
rect 8382 11754 8442 11756
rect 9398 11754 9458 11756
rect 1744 11700 1826 11724
rect 1998 11720 2014 11754
rect 2570 11720 2586 11754
rect 1744 11666 1768 11700
rect 1802 11666 1826 11700
rect 1744 11642 1826 11666
rect 2762 11700 2844 11724
rect 3016 11720 3032 11754
rect 3588 11720 3604 11754
rect 2762 11666 2786 11700
rect 2820 11666 2844 11700
rect 1998 11612 2014 11646
rect 2570 11612 2586 11646
rect 2762 11642 2844 11666
rect 3780 11700 3862 11724
rect 4034 11720 4050 11754
rect 4606 11720 4622 11754
rect 3780 11666 3804 11700
rect 3838 11666 3862 11700
rect 3016 11612 3032 11646
rect 3588 11612 3604 11646
rect 3780 11642 3862 11666
rect 4798 11700 4880 11724
rect 5052 11720 5068 11754
rect 5624 11720 5640 11754
rect 4798 11666 4822 11700
rect 4856 11666 4880 11700
rect 4034 11612 4050 11646
rect 4606 11612 4622 11646
rect 4798 11642 4880 11666
rect 5816 11700 5898 11724
rect 6070 11720 6086 11754
rect 6642 11720 6658 11754
rect 5816 11666 5840 11700
rect 5874 11666 5898 11700
rect 5052 11612 5068 11646
rect 5624 11612 5640 11646
rect 5816 11642 5898 11666
rect 6834 11700 6916 11724
rect 7088 11720 7104 11754
rect 7660 11720 7676 11754
rect 6834 11666 6858 11700
rect 6892 11666 6916 11700
rect 6070 11612 6086 11646
rect 6642 11612 6658 11646
rect 6834 11642 6916 11666
rect 7852 11700 7934 11724
rect 8106 11720 8122 11754
rect 8678 11720 8694 11754
rect 7852 11666 7876 11700
rect 7910 11666 7934 11700
rect 7088 11612 7104 11646
rect 7660 11612 7676 11646
rect 7852 11642 7934 11666
rect 8870 11700 8952 11724
rect 9124 11720 9140 11754
rect 9696 11720 9712 11754
rect 8870 11666 8894 11700
rect 8928 11666 8952 11700
rect 8106 11612 8122 11646
rect 8678 11612 8694 11646
rect 8870 11642 8952 11666
rect 9888 11700 9970 11724
rect 10142 11720 10158 11754
rect 10714 11720 10730 11754
rect 13532 11752 13566 11768
rect 14550 12344 14584 12360
rect 14550 11752 14584 11768
rect 15568 12344 15602 12360
rect 15568 11752 15602 11768
rect 16586 12344 16620 12360
rect 16586 11752 16620 11768
rect 17604 12344 17638 12360
rect 17604 11752 17638 11768
rect 18622 12344 18656 12360
rect 18622 11752 18656 11768
rect 19640 12344 19674 12360
rect 19640 11752 19674 11768
rect 20658 12344 20692 12360
rect 20658 11752 20692 11768
rect 21676 12344 21710 12360
rect 21676 11752 21710 11768
rect 22694 12344 22728 12360
rect 22694 11752 22728 11768
rect 23712 12344 23746 12360
rect 23712 11752 23746 11768
rect 24730 12344 24764 12360
rect 24730 11752 24764 11768
rect 25748 12344 25782 12360
rect 25748 11752 25782 11768
rect 26766 12344 26800 12360
rect 26766 11752 26800 11768
rect 27784 12344 27818 12360
rect 27784 11752 27818 11768
rect 28802 12344 28836 12360
rect 28802 11752 28836 11768
rect 29820 12344 29854 12360
rect 29820 11752 29854 11768
rect 30838 12344 30872 12360
rect 30838 11752 30872 11768
rect 31856 12344 31890 12360
rect 31856 11752 31890 11768
rect 32874 12344 32908 12360
rect 32874 11752 32908 11768
rect 33892 12344 33926 12360
rect 33892 11752 33926 11768
rect 9888 11666 9912 11700
rect 9946 11666 9970 11700
rect 9124 11612 9140 11646
rect 9696 11612 9712 11646
rect 9888 11642 9970 11666
rect 10906 11700 10988 11724
rect 17076 11718 17136 11720
rect 10906 11666 10930 11700
rect 10964 11666 10988 11700
rect 13764 11684 13780 11718
rect 14336 11684 14352 11718
rect 14782 11684 14798 11718
rect 15354 11684 15370 11718
rect 15800 11684 15816 11718
rect 16372 11684 16388 11718
rect 16818 11684 16834 11718
rect 17390 11684 17406 11718
rect 17836 11684 17852 11718
rect 18408 11684 18424 11718
rect 18854 11684 18870 11718
rect 19426 11684 19442 11718
rect 19872 11684 19888 11718
rect 20444 11684 20460 11718
rect 20890 11684 20906 11718
rect 21462 11684 21478 11718
rect 21908 11684 21924 11718
rect 22480 11684 22496 11718
rect 22926 11684 22942 11718
rect 23498 11684 23514 11718
rect 23944 11684 23960 11718
rect 24516 11684 24532 11718
rect 24962 11684 24978 11718
rect 25534 11684 25550 11718
rect 25980 11684 25996 11718
rect 26552 11684 26568 11718
rect 26998 11684 27014 11718
rect 27570 11684 27586 11718
rect 28016 11684 28032 11718
rect 28588 11684 28604 11718
rect 29034 11684 29050 11718
rect 29606 11684 29622 11718
rect 30052 11684 30068 11718
rect 30624 11684 30640 11718
rect 31070 11684 31086 11718
rect 31642 11684 31658 11718
rect 32088 11684 32104 11718
rect 32660 11684 32676 11718
rect 33106 11684 33122 11718
rect 33678 11684 33694 11718
rect 19110 11680 19170 11684
rect 28268 11670 28328 11684
rect 29302 11670 29362 11684
rect 10142 11612 10158 11646
rect 10714 11612 10730 11646
rect 10906 11642 10988 11666
rect 1766 11562 1800 11578
rect 1766 10970 1800 10986
rect 2784 11562 2818 11578
rect 2784 10970 2818 10986
rect 3802 11562 3836 11578
rect 3802 10970 3836 10986
rect 4820 11562 4854 11578
rect 4820 10970 4854 10986
rect 5838 11562 5872 11578
rect 5838 10970 5872 10986
rect 6856 11562 6890 11578
rect 6856 10970 6890 10986
rect 7874 11562 7908 11578
rect 7874 10970 7908 10986
rect 8892 11562 8926 11578
rect 8892 10970 8926 10986
rect 9910 11562 9944 11578
rect 9910 10970 9944 10986
rect 10928 11562 10962 11578
rect 14016 11456 14098 11480
rect 14016 11422 14040 11456
rect 14074 11422 14098 11456
rect 14016 11398 14098 11422
rect 15034 11456 15116 11480
rect 15034 11422 15058 11456
rect 15092 11422 15116 11456
rect 15034 11398 15116 11422
rect 16052 11456 16134 11480
rect 16052 11422 16076 11456
rect 16110 11422 16134 11456
rect 16052 11398 16134 11422
rect 17070 11456 17152 11480
rect 17070 11422 17094 11456
rect 17128 11422 17152 11456
rect 17070 11398 17152 11422
rect 18088 11456 18170 11480
rect 18088 11422 18112 11456
rect 18146 11422 18170 11456
rect 18088 11398 18170 11422
rect 19106 11456 19188 11480
rect 19106 11422 19130 11456
rect 19164 11422 19188 11456
rect 19106 11398 19188 11422
rect 20124 11456 20206 11480
rect 20124 11422 20148 11456
rect 20182 11422 20206 11456
rect 20124 11398 20206 11422
rect 21142 11456 21224 11480
rect 21142 11422 21166 11456
rect 21200 11422 21224 11456
rect 21142 11398 21224 11422
rect 22160 11456 22242 11480
rect 22160 11422 22184 11456
rect 22218 11422 22242 11456
rect 22160 11398 22242 11422
rect 23178 11456 23260 11480
rect 23178 11422 23202 11456
rect 23236 11422 23260 11456
rect 23178 11398 23260 11422
rect 24196 11456 24278 11480
rect 24196 11422 24220 11456
rect 24254 11422 24278 11456
rect 24196 11398 24278 11422
rect 25214 11456 25296 11480
rect 25214 11422 25238 11456
rect 25272 11422 25296 11456
rect 25214 11398 25296 11422
rect 26232 11456 26314 11480
rect 26232 11422 26256 11456
rect 26290 11422 26314 11456
rect 26232 11398 26314 11422
rect 27250 11456 27332 11480
rect 27250 11422 27274 11456
rect 27308 11422 27332 11456
rect 27250 11398 27332 11422
rect 28268 11456 28350 11480
rect 28268 11422 28292 11456
rect 28326 11422 28350 11456
rect 28268 11398 28350 11422
rect 29286 11456 29368 11480
rect 29286 11422 29310 11456
rect 29344 11422 29368 11456
rect 29286 11398 29368 11422
rect 30304 11456 30386 11480
rect 30304 11422 30328 11456
rect 30362 11422 30386 11456
rect 30304 11398 30386 11422
rect 31322 11456 31404 11480
rect 31322 11422 31346 11456
rect 31380 11422 31404 11456
rect 31322 11398 31404 11422
rect 32340 11456 32422 11480
rect 32340 11422 32364 11456
rect 32398 11422 32422 11456
rect 32340 11398 32422 11422
rect 33358 11456 33440 11480
rect 33358 11422 33382 11456
rect 33416 11422 33440 11456
rect 33358 11398 33440 11422
rect 13762 11160 13778 11194
rect 14334 11160 14350 11194
rect 14780 11160 14796 11194
rect 15352 11160 15368 11194
rect 15798 11160 15814 11194
rect 16370 11160 16386 11194
rect 16816 11160 16832 11194
rect 17388 11160 17404 11194
rect 17834 11160 17850 11194
rect 18406 11160 18422 11194
rect 18852 11160 18868 11194
rect 19424 11160 19440 11194
rect 19870 11160 19886 11194
rect 20442 11160 20458 11194
rect 20888 11160 20904 11194
rect 21460 11160 21476 11194
rect 21906 11160 21922 11194
rect 22478 11160 22494 11194
rect 22924 11160 22940 11194
rect 23496 11160 23512 11194
rect 23942 11160 23958 11194
rect 24514 11160 24530 11194
rect 24960 11160 24976 11194
rect 25532 11160 25548 11194
rect 25978 11160 25994 11194
rect 26550 11160 26566 11194
rect 26996 11160 27012 11194
rect 27568 11160 27584 11194
rect 28014 11160 28030 11194
rect 28586 11160 28602 11194
rect 29032 11160 29048 11194
rect 29604 11160 29620 11194
rect 30050 11160 30066 11194
rect 30622 11160 30638 11194
rect 31068 11160 31084 11194
rect 31640 11160 31656 11194
rect 32086 11160 32102 11194
rect 32658 11160 32674 11194
rect 33104 11160 33120 11194
rect 33676 11160 33692 11194
rect 16072 11156 16132 11160
rect 10928 10970 10962 10986
rect 13530 11110 13564 11126
rect 1744 10882 1826 10906
rect 1998 10902 2014 10936
rect 2570 10902 2586 10936
rect 1744 10848 1768 10882
rect 1802 10848 1826 10882
rect 1744 10824 1826 10848
rect 2762 10882 2844 10906
rect 3016 10902 3032 10936
rect 3588 10902 3604 10936
rect 2762 10848 2786 10882
rect 2820 10848 2844 10882
rect 1998 10794 2014 10828
rect 2570 10794 2586 10828
rect 2762 10824 2844 10848
rect 3780 10882 3862 10906
rect 4034 10902 4050 10936
rect 4606 10902 4622 10936
rect 3780 10848 3804 10882
rect 3838 10848 3862 10882
rect 3016 10794 3032 10828
rect 3588 10794 3604 10828
rect 3780 10824 3862 10848
rect 4798 10882 4880 10906
rect 5052 10902 5068 10936
rect 5624 10902 5640 10936
rect 4798 10848 4822 10882
rect 4856 10848 4880 10882
rect 4034 10794 4050 10828
rect 4606 10794 4622 10828
rect 4798 10824 4880 10848
rect 5816 10882 5898 10906
rect 6070 10902 6086 10936
rect 6642 10902 6658 10936
rect 5816 10848 5840 10882
rect 5874 10848 5898 10882
rect 5052 10794 5068 10828
rect 5624 10794 5640 10828
rect 5816 10824 5898 10848
rect 6834 10882 6916 10906
rect 7088 10902 7104 10936
rect 7660 10902 7676 10936
rect 6834 10848 6858 10882
rect 6892 10848 6916 10882
rect 6070 10794 6086 10828
rect 6642 10794 6658 10828
rect 6834 10824 6916 10848
rect 7852 10882 7934 10906
rect 8106 10902 8122 10936
rect 8678 10902 8694 10936
rect 7852 10848 7876 10882
rect 7910 10848 7934 10882
rect 7088 10794 7104 10828
rect 7660 10794 7676 10828
rect 7852 10824 7934 10848
rect 8870 10882 8952 10906
rect 9124 10902 9140 10936
rect 9696 10902 9712 10936
rect 8870 10848 8894 10882
rect 8928 10848 8952 10882
rect 8106 10794 8122 10828
rect 8678 10794 8694 10828
rect 8870 10824 8952 10848
rect 9888 10882 9970 10906
rect 10142 10902 10158 10936
rect 10714 10902 10730 10936
rect 9888 10848 9912 10882
rect 9946 10848 9970 10882
rect 9124 10794 9140 10828
rect 9696 10794 9712 10828
rect 9888 10824 9970 10848
rect 10906 10882 10988 10906
rect 10906 10848 10930 10882
rect 10964 10848 10988 10882
rect 10142 10794 10158 10828
rect 10714 10794 10730 10828
rect 10906 10824 10988 10848
rect 7354 10792 7414 10794
rect 1766 10744 1800 10760
rect 1766 10152 1800 10168
rect 2784 10744 2818 10760
rect 2784 10152 2818 10168
rect 3802 10744 3836 10760
rect 3802 10152 3836 10168
rect 4820 10744 4854 10760
rect 4820 10152 4854 10168
rect 5838 10744 5872 10760
rect 5838 10152 5872 10168
rect 6856 10744 6890 10760
rect 6856 10152 6890 10168
rect 7874 10744 7908 10760
rect 7874 10152 7908 10168
rect 8892 10744 8926 10760
rect 8892 10152 8926 10168
rect 9910 10744 9944 10760
rect 9910 10152 9944 10168
rect 10928 10744 10962 10760
rect 13530 10518 13564 10534
rect 14548 11110 14582 11126
rect 14548 10518 14582 10534
rect 15566 11110 15600 11126
rect 15566 10518 15600 10534
rect 16584 11110 16618 11126
rect 16584 10518 16618 10534
rect 17602 11110 17636 11126
rect 17602 10518 17636 10534
rect 18620 11110 18654 11126
rect 18620 10518 18654 10534
rect 19638 11110 19672 11126
rect 19638 10518 19672 10534
rect 20656 11110 20690 11126
rect 20656 10518 20690 10534
rect 21674 11110 21708 11126
rect 21674 10518 21708 10534
rect 22692 11110 22726 11126
rect 22692 10518 22726 10534
rect 23710 11110 23744 11126
rect 23710 10518 23744 10534
rect 24728 11110 24762 11126
rect 24728 10518 24762 10534
rect 25746 11110 25780 11126
rect 25746 10518 25780 10534
rect 26764 11110 26798 11126
rect 26764 10518 26798 10534
rect 27782 11110 27816 11126
rect 27782 10518 27816 10534
rect 28800 11110 28834 11126
rect 28800 10518 28834 10534
rect 29818 11110 29852 11126
rect 29818 10518 29852 10534
rect 30836 11110 30870 11126
rect 30836 10518 30870 10534
rect 31854 11110 31888 11126
rect 31854 10518 31888 10534
rect 32872 11110 32906 11126
rect 32872 10518 32906 10534
rect 33890 11110 33924 11126
rect 33890 10518 33924 10534
rect 21140 10484 21200 10488
rect 22168 10484 22228 10486
rect 24212 10484 24272 10488
rect 13762 10450 13778 10484
rect 14334 10450 14350 10484
rect 14780 10450 14796 10484
rect 15352 10450 15368 10484
rect 15798 10450 15814 10484
rect 16370 10450 16386 10484
rect 16816 10450 16832 10484
rect 17388 10450 17404 10484
rect 17834 10450 17850 10484
rect 18406 10450 18422 10484
rect 18852 10450 18868 10484
rect 19424 10450 19440 10484
rect 19870 10450 19886 10484
rect 20442 10450 20458 10484
rect 20888 10450 20904 10484
rect 21460 10450 21476 10484
rect 21906 10450 21922 10484
rect 22478 10450 22494 10484
rect 22924 10450 22940 10484
rect 23496 10450 23512 10484
rect 23942 10450 23958 10484
rect 24514 10450 24530 10484
rect 24960 10450 24976 10484
rect 25532 10450 25548 10484
rect 25978 10450 25994 10484
rect 26550 10450 26566 10484
rect 26996 10450 27012 10484
rect 27568 10450 27584 10484
rect 28014 10450 28030 10484
rect 28586 10450 28602 10484
rect 29032 10450 29048 10484
rect 29604 10450 29620 10484
rect 30050 10450 30066 10484
rect 30622 10450 30638 10484
rect 31068 10450 31084 10484
rect 31640 10450 31656 10484
rect 32086 10450 32102 10484
rect 32658 10450 32674 10484
rect 33104 10450 33120 10484
rect 33676 10450 33692 10484
rect 14016 10236 14098 10260
rect 14016 10202 14040 10236
rect 14074 10202 14098 10236
rect 14016 10178 14098 10202
rect 15034 10236 15116 10260
rect 15034 10202 15058 10236
rect 15092 10202 15116 10236
rect 15034 10178 15116 10202
rect 16052 10236 16134 10260
rect 16052 10202 16076 10236
rect 16110 10202 16134 10236
rect 16052 10178 16134 10202
rect 17070 10236 17152 10260
rect 17070 10202 17094 10236
rect 17128 10202 17152 10236
rect 17070 10178 17152 10202
rect 18088 10236 18170 10260
rect 18088 10202 18112 10236
rect 18146 10202 18170 10236
rect 18088 10178 18170 10202
rect 19106 10236 19188 10260
rect 19106 10202 19130 10236
rect 19164 10202 19188 10236
rect 19106 10178 19188 10202
rect 20124 10236 20206 10260
rect 20124 10202 20148 10236
rect 20182 10202 20206 10236
rect 20124 10178 20206 10202
rect 21142 10236 21224 10260
rect 21142 10202 21166 10236
rect 21200 10202 21224 10236
rect 21142 10178 21224 10202
rect 22160 10236 22242 10260
rect 22160 10202 22184 10236
rect 22218 10202 22242 10236
rect 22160 10178 22242 10202
rect 23178 10236 23260 10260
rect 23178 10202 23202 10236
rect 23236 10202 23260 10236
rect 23178 10178 23260 10202
rect 24196 10236 24278 10260
rect 24196 10202 24220 10236
rect 24254 10202 24278 10236
rect 24196 10178 24278 10202
rect 25214 10236 25296 10260
rect 25214 10202 25238 10236
rect 25272 10202 25296 10236
rect 25214 10178 25296 10202
rect 26232 10236 26314 10260
rect 26232 10202 26256 10236
rect 26290 10202 26314 10236
rect 26232 10178 26314 10202
rect 27250 10236 27332 10260
rect 27250 10202 27274 10236
rect 27308 10202 27332 10236
rect 27250 10178 27332 10202
rect 28268 10236 28350 10260
rect 28268 10202 28292 10236
rect 28326 10202 28350 10236
rect 28268 10178 28350 10202
rect 29286 10236 29368 10260
rect 29286 10202 29310 10236
rect 29344 10202 29368 10236
rect 29286 10178 29368 10202
rect 30304 10236 30386 10260
rect 30304 10202 30328 10236
rect 30362 10202 30386 10236
rect 30304 10178 30386 10202
rect 31322 10236 31404 10260
rect 31322 10202 31346 10236
rect 31380 10202 31404 10236
rect 31322 10178 31404 10202
rect 32340 10236 32422 10260
rect 32340 10202 32364 10236
rect 32398 10202 32422 10236
rect 32340 10178 32422 10202
rect 33358 10236 33440 10260
rect 33358 10202 33382 10236
rect 33416 10202 33440 10236
rect 33358 10178 33440 10202
rect 10928 10152 10962 10168
rect 3280 10118 3340 10120
rect 4294 10118 4354 10120
rect 8368 10118 8428 10120
rect 9384 10118 9444 10120
rect 1744 10064 1826 10088
rect 1998 10084 2014 10118
rect 2570 10084 2586 10118
rect 1744 10030 1768 10064
rect 1802 10030 1826 10064
rect 1744 10006 1826 10030
rect 2762 10064 2844 10088
rect 3016 10084 3032 10118
rect 3588 10084 3604 10118
rect 2762 10030 2786 10064
rect 2820 10030 2844 10064
rect 1998 9976 2014 10010
rect 2570 9976 2586 10010
rect 2762 10006 2844 10030
rect 3780 10064 3862 10088
rect 4034 10084 4050 10118
rect 4606 10084 4622 10118
rect 3780 10030 3804 10064
rect 3838 10030 3862 10064
rect 3016 9976 3032 10010
rect 3588 9976 3604 10010
rect 3780 10006 3862 10030
rect 4798 10064 4880 10088
rect 5052 10084 5068 10118
rect 5624 10084 5640 10118
rect 4798 10030 4822 10064
rect 4856 10030 4880 10064
rect 4034 9976 4050 10010
rect 4606 9976 4622 10010
rect 4798 10006 4880 10030
rect 5816 10064 5898 10088
rect 6070 10084 6086 10118
rect 6642 10084 6658 10118
rect 5816 10030 5840 10064
rect 5874 10030 5898 10064
rect 5052 9976 5068 10010
rect 5624 9976 5640 10010
rect 5816 10006 5898 10030
rect 6834 10064 6916 10088
rect 7088 10084 7104 10118
rect 7660 10084 7676 10118
rect 6834 10030 6858 10064
rect 6892 10030 6916 10064
rect 6070 9976 6086 10010
rect 6642 9976 6658 10010
rect 6834 10006 6916 10030
rect 7852 10064 7934 10088
rect 8106 10084 8122 10118
rect 8678 10084 8694 10118
rect 7852 10030 7876 10064
rect 7910 10030 7934 10064
rect 7088 9976 7104 10010
rect 7660 9976 7676 10010
rect 7852 10006 7934 10030
rect 8870 10064 8952 10088
rect 9124 10084 9140 10118
rect 9696 10084 9712 10118
rect 8870 10030 8894 10064
rect 8928 10030 8952 10064
rect 8106 9976 8122 10010
rect 8678 9976 8694 10010
rect 8870 10006 8952 10030
rect 9888 10064 9970 10088
rect 10142 10084 10158 10118
rect 10714 10084 10730 10118
rect 9888 10030 9912 10064
rect 9946 10030 9970 10064
rect 9124 9976 9140 10010
rect 9696 9976 9712 10010
rect 9888 10006 9970 10030
rect 10906 10064 10988 10088
rect 10906 10030 10930 10064
rect 10964 10030 10988 10064
rect 10142 9976 10158 10010
rect 10714 9976 10730 10010
rect 10906 10006 10988 10030
rect 1766 9926 1800 9942
rect 1766 9334 1800 9350
rect 2784 9926 2818 9942
rect 2784 9334 2818 9350
rect 3802 9926 3836 9942
rect 3802 9334 3836 9350
rect 4820 9926 4854 9942
rect 4820 9334 4854 9350
rect 5838 9926 5872 9942
rect 5838 9334 5872 9350
rect 6856 9926 6890 9942
rect 6856 9334 6890 9350
rect 7874 9926 7908 9942
rect 7874 9334 7908 9350
rect 8892 9926 8926 9942
rect 8892 9334 8926 9350
rect 9910 9926 9944 9942
rect 9910 9334 9944 9350
rect 10928 9926 10962 9942
rect 13762 9926 13778 9960
rect 14334 9926 14350 9960
rect 14780 9926 14796 9960
rect 15352 9926 15368 9960
rect 15798 9926 15814 9960
rect 16370 9926 16386 9960
rect 16816 9926 16832 9960
rect 17388 9926 17404 9960
rect 17834 9926 17850 9960
rect 18406 9926 18422 9960
rect 18852 9926 18868 9960
rect 19424 9926 19440 9960
rect 19870 9926 19886 9960
rect 20442 9926 20458 9960
rect 20888 9926 20904 9960
rect 21460 9926 21476 9960
rect 21906 9926 21922 9960
rect 22478 9926 22494 9960
rect 22924 9926 22940 9960
rect 23496 9926 23512 9960
rect 23942 9926 23958 9960
rect 24514 9926 24530 9960
rect 24960 9926 24976 9960
rect 25532 9926 25548 9960
rect 25978 9926 25994 9960
rect 26550 9926 26566 9960
rect 26996 9926 27012 9960
rect 27568 9926 27584 9960
rect 28014 9926 28030 9960
rect 28586 9926 28602 9960
rect 29032 9926 29048 9960
rect 29604 9926 29620 9960
rect 30050 9926 30066 9960
rect 30622 9926 30638 9960
rect 31068 9926 31084 9960
rect 31640 9926 31656 9960
rect 32086 9926 32102 9960
rect 32658 9926 32674 9960
rect 33104 9926 33120 9960
rect 33676 9926 33692 9960
rect 10928 9334 10962 9350
rect 13530 9876 13564 9892
rect 3284 9300 3344 9302
rect 4298 9300 4358 9302
rect 8372 9300 8432 9302
rect 9388 9300 9448 9302
rect 1744 9246 1826 9270
rect 1998 9266 2014 9300
rect 2570 9266 2586 9300
rect 1744 9212 1768 9246
rect 1802 9212 1826 9246
rect 1744 9188 1826 9212
rect 2762 9246 2844 9270
rect 3016 9266 3032 9300
rect 3588 9266 3604 9300
rect 2762 9212 2786 9246
rect 2820 9212 2844 9246
rect 1998 9158 2014 9192
rect 2570 9158 2586 9192
rect 2762 9188 2844 9212
rect 3780 9246 3862 9270
rect 4034 9266 4050 9300
rect 4606 9266 4622 9300
rect 3780 9212 3804 9246
rect 3838 9212 3862 9246
rect 3016 9158 3032 9192
rect 3588 9158 3604 9192
rect 3780 9188 3862 9212
rect 4798 9246 4880 9270
rect 5052 9266 5068 9300
rect 5624 9266 5640 9300
rect 4798 9212 4822 9246
rect 4856 9212 4880 9246
rect 4034 9158 4050 9192
rect 4606 9158 4622 9192
rect 4798 9188 4880 9212
rect 5816 9246 5898 9270
rect 6070 9266 6086 9300
rect 6642 9266 6658 9300
rect 5816 9212 5840 9246
rect 5874 9212 5898 9246
rect 5052 9158 5068 9192
rect 5624 9158 5640 9192
rect 5816 9188 5898 9212
rect 6834 9246 6916 9270
rect 7088 9266 7104 9300
rect 7660 9266 7676 9300
rect 6834 9212 6858 9246
rect 6892 9212 6916 9246
rect 6070 9158 6086 9192
rect 6642 9158 6658 9192
rect 6834 9188 6916 9212
rect 7852 9246 7934 9270
rect 8106 9266 8122 9300
rect 8678 9266 8694 9300
rect 7852 9212 7876 9246
rect 7910 9212 7934 9246
rect 7088 9158 7104 9192
rect 7660 9158 7676 9192
rect 7852 9188 7934 9212
rect 8870 9246 8952 9270
rect 9124 9266 9140 9300
rect 9696 9266 9712 9300
rect 8870 9212 8894 9246
rect 8928 9212 8952 9246
rect 8106 9158 8122 9192
rect 8678 9158 8694 9192
rect 8870 9188 8952 9212
rect 9888 9246 9970 9270
rect 10142 9266 10158 9300
rect 10714 9266 10730 9300
rect 13530 9284 13564 9300
rect 14548 9876 14582 9892
rect 14548 9284 14582 9300
rect 15566 9876 15600 9892
rect 15566 9284 15600 9300
rect 16584 9876 16618 9892
rect 16584 9284 16618 9300
rect 17602 9876 17636 9892
rect 17602 9284 17636 9300
rect 18620 9876 18654 9892
rect 18620 9284 18654 9300
rect 19638 9876 19672 9892
rect 19638 9284 19672 9300
rect 20656 9876 20690 9892
rect 20656 9284 20690 9300
rect 21674 9876 21708 9892
rect 21674 9284 21708 9300
rect 22692 9876 22726 9892
rect 22692 9284 22726 9300
rect 23710 9876 23744 9892
rect 23710 9284 23744 9300
rect 24728 9876 24762 9892
rect 24728 9284 24762 9300
rect 25746 9876 25780 9892
rect 25746 9284 25780 9300
rect 26764 9876 26798 9892
rect 26764 9284 26798 9300
rect 27782 9876 27816 9892
rect 27782 9284 27816 9300
rect 28800 9876 28834 9892
rect 28800 9284 28834 9300
rect 29818 9876 29852 9892
rect 29818 9284 29852 9300
rect 30836 9876 30870 9892
rect 30836 9284 30870 9300
rect 31854 9876 31888 9892
rect 31854 9284 31888 9300
rect 32872 9876 32906 9892
rect 32872 9284 32906 9300
rect 33890 9876 33924 9892
rect 33890 9284 33924 9300
rect 9888 9212 9912 9246
rect 9946 9212 9970 9246
rect 9124 9158 9140 9192
rect 9696 9158 9712 9192
rect 9888 9188 9970 9212
rect 10906 9246 10988 9270
rect 10906 9212 10930 9246
rect 10964 9212 10988 9246
rect 13762 9216 13778 9250
rect 14334 9216 14350 9250
rect 14780 9216 14796 9250
rect 15352 9216 15368 9250
rect 15798 9216 15814 9250
rect 16370 9216 16386 9250
rect 16816 9216 16832 9250
rect 17388 9216 17404 9250
rect 17834 9216 17850 9250
rect 18406 9216 18422 9250
rect 18852 9216 18868 9250
rect 19424 9216 19440 9250
rect 19870 9216 19886 9250
rect 20442 9216 20458 9250
rect 20888 9216 20904 9250
rect 21460 9216 21476 9250
rect 21906 9216 21922 9250
rect 22478 9216 22494 9250
rect 22924 9216 22940 9250
rect 23496 9216 23512 9250
rect 23942 9216 23958 9250
rect 24514 9216 24530 9250
rect 24960 9216 24976 9250
rect 25532 9216 25548 9250
rect 25978 9216 25994 9250
rect 26550 9216 26566 9250
rect 26996 9216 27012 9250
rect 27568 9216 27584 9250
rect 28014 9216 28030 9250
rect 28586 9216 28602 9250
rect 29032 9216 29048 9250
rect 29604 9216 29620 9250
rect 30050 9216 30066 9250
rect 30622 9216 30638 9250
rect 31068 9216 31084 9250
rect 31640 9216 31656 9250
rect 32086 9216 32102 9250
rect 32658 9216 32674 9250
rect 33104 9216 33120 9250
rect 33676 9216 33692 9250
rect 10142 9158 10158 9192
rect 10714 9158 10730 9192
rect 10906 9188 10988 9212
rect 1766 9108 1800 9124
rect 1766 8516 1800 8532
rect 2784 9108 2818 9124
rect 2784 8516 2818 8532
rect 3802 9108 3836 9124
rect 3802 8516 3836 8532
rect 4820 9108 4854 9124
rect 4820 8516 4854 8532
rect 5838 9108 5872 9124
rect 5838 8516 5872 8532
rect 6856 9108 6890 9124
rect 6856 8516 6890 8532
rect 7874 9108 7908 9124
rect 7874 8516 7908 8532
rect 8892 9108 8926 9124
rect 8892 8516 8926 8532
rect 9910 9108 9944 9124
rect 9910 8516 9944 8532
rect 10928 9108 10962 9124
rect 14030 8988 14112 9012
rect 14030 8954 14054 8988
rect 14088 8954 14112 8988
rect 14030 8930 14112 8954
rect 15048 8988 15130 9012
rect 15048 8954 15072 8988
rect 15106 8954 15130 8988
rect 15048 8930 15130 8954
rect 16066 8988 16148 9012
rect 16066 8954 16090 8988
rect 16124 8954 16148 8988
rect 16066 8930 16148 8954
rect 17084 8988 17166 9012
rect 17084 8954 17108 8988
rect 17142 8954 17166 8988
rect 17084 8930 17166 8954
rect 18102 8988 18184 9012
rect 18102 8954 18126 8988
rect 18160 8954 18184 8988
rect 18102 8930 18184 8954
rect 19120 8988 19202 9012
rect 19120 8954 19144 8988
rect 19178 8954 19202 8988
rect 19120 8930 19202 8954
rect 20138 8988 20220 9012
rect 20138 8954 20162 8988
rect 20196 8954 20220 8988
rect 20138 8930 20220 8954
rect 21156 8988 21238 9012
rect 21156 8954 21180 8988
rect 21214 8954 21238 8988
rect 21156 8930 21238 8954
rect 22174 8988 22256 9012
rect 22174 8954 22198 8988
rect 22232 8954 22256 8988
rect 22174 8930 22256 8954
rect 23192 8988 23274 9012
rect 23192 8954 23216 8988
rect 23250 8954 23274 8988
rect 23192 8930 23274 8954
rect 24210 8988 24292 9012
rect 24210 8954 24234 8988
rect 24268 8954 24292 8988
rect 24210 8930 24292 8954
rect 25228 8988 25310 9012
rect 25228 8954 25252 8988
rect 25286 8954 25310 8988
rect 25228 8930 25310 8954
rect 26246 8988 26328 9012
rect 26246 8954 26270 8988
rect 26304 8954 26328 8988
rect 26246 8930 26328 8954
rect 27264 8988 27346 9012
rect 27264 8954 27288 8988
rect 27322 8954 27346 8988
rect 27264 8930 27346 8954
rect 28282 8988 28364 9012
rect 28282 8954 28306 8988
rect 28340 8954 28364 8988
rect 28282 8930 28364 8954
rect 29300 8988 29382 9012
rect 29300 8954 29324 8988
rect 29358 8954 29382 8988
rect 29300 8930 29382 8954
rect 30318 8988 30400 9012
rect 30318 8954 30342 8988
rect 30376 8954 30400 8988
rect 30318 8930 30400 8954
rect 31336 8988 31418 9012
rect 31336 8954 31360 8988
rect 31394 8954 31418 8988
rect 31336 8930 31418 8954
rect 32354 8988 32436 9012
rect 32354 8954 32378 8988
rect 32412 8954 32436 8988
rect 32354 8930 32436 8954
rect 33372 8988 33454 9012
rect 33372 8954 33396 8988
rect 33430 8954 33454 8988
rect 33372 8930 33454 8954
rect 13762 8694 13778 8728
rect 14334 8694 14350 8728
rect 14780 8694 14796 8728
rect 15352 8694 15368 8728
rect 15798 8694 15814 8728
rect 16370 8694 16386 8728
rect 16816 8694 16832 8728
rect 17388 8694 17404 8728
rect 17834 8694 17850 8728
rect 18406 8694 18422 8728
rect 18852 8694 18868 8728
rect 19424 8694 19440 8728
rect 19870 8694 19886 8728
rect 20442 8694 20458 8728
rect 20888 8694 20904 8728
rect 21460 8694 21476 8728
rect 21906 8694 21922 8728
rect 22478 8694 22494 8728
rect 22924 8694 22940 8728
rect 23496 8694 23512 8728
rect 23942 8694 23958 8728
rect 24514 8694 24530 8728
rect 24960 8694 24976 8728
rect 25532 8694 25548 8728
rect 25978 8694 25994 8728
rect 26550 8694 26566 8728
rect 26996 8694 27012 8728
rect 27568 8694 27584 8728
rect 28014 8694 28030 8728
rect 28586 8694 28602 8728
rect 29032 8694 29048 8728
rect 29604 8694 29620 8728
rect 30050 8694 30066 8728
rect 30622 8694 30638 8728
rect 31068 8694 31084 8728
rect 31640 8694 31656 8728
rect 32086 8694 32102 8728
rect 32658 8694 32674 8728
rect 33104 8694 33120 8728
rect 33676 8694 33692 8728
rect 10928 8516 10962 8532
rect 13530 8644 13564 8660
rect 2258 8482 2318 8484
rect 3284 8482 3344 8486
rect 4298 8482 4358 8486
rect 5318 8482 5378 8484
rect 6340 8482 6400 8484
rect 8372 8482 8432 8486
rect 9388 8482 9448 8486
rect 10408 8482 10468 8484
rect 1744 8428 1826 8452
rect 1998 8448 2014 8482
rect 2570 8448 2586 8482
rect 1744 8394 1768 8428
rect 1802 8394 1826 8428
rect 1744 8370 1826 8394
rect 2762 8428 2844 8452
rect 3016 8448 3032 8482
rect 3588 8448 3604 8482
rect 2762 8394 2786 8428
rect 2820 8394 2844 8428
rect 1998 8340 2014 8374
rect 2570 8340 2586 8374
rect 2762 8370 2844 8394
rect 3780 8428 3862 8452
rect 4034 8448 4050 8482
rect 4606 8448 4622 8482
rect 3780 8394 3804 8428
rect 3838 8394 3862 8428
rect 3016 8340 3032 8374
rect 3588 8340 3604 8374
rect 3780 8370 3862 8394
rect 4798 8428 4880 8452
rect 5052 8448 5068 8482
rect 5624 8448 5640 8482
rect 4798 8394 4822 8428
rect 4856 8394 4880 8428
rect 4034 8340 4050 8374
rect 4606 8340 4622 8374
rect 4798 8370 4880 8394
rect 5816 8428 5898 8452
rect 6070 8448 6086 8482
rect 6642 8448 6658 8482
rect 5816 8394 5840 8428
rect 5874 8394 5898 8428
rect 5052 8340 5068 8374
rect 5624 8340 5640 8374
rect 5816 8370 5898 8394
rect 6834 8428 6916 8452
rect 7088 8448 7104 8482
rect 7660 8448 7676 8482
rect 6834 8394 6858 8428
rect 6892 8394 6916 8428
rect 6070 8340 6086 8374
rect 6642 8340 6658 8374
rect 6834 8370 6916 8394
rect 7852 8428 7934 8452
rect 8106 8448 8122 8482
rect 8678 8448 8694 8482
rect 7852 8394 7876 8428
rect 7910 8394 7934 8428
rect 7088 8340 7104 8374
rect 7660 8340 7676 8374
rect 7852 8370 7934 8394
rect 8870 8428 8952 8452
rect 9124 8448 9140 8482
rect 9696 8448 9712 8482
rect 8870 8394 8894 8428
rect 8928 8394 8952 8428
rect 8106 8340 8122 8374
rect 8678 8340 8694 8374
rect 8870 8370 8952 8394
rect 9888 8428 9970 8452
rect 10142 8448 10158 8482
rect 10714 8448 10730 8482
rect 9888 8394 9912 8428
rect 9946 8394 9970 8428
rect 9124 8340 9140 8374
rect 9696 8340 9712 8374
rect 9888 8370 9970 8394
rect 10906 8428 10988 8452
rect 10906 8394 10930 8428
rect 10964 8394 10988 8428
rect 10142 8340 10158 8374
rect 10714 8340 10730 8374
rect 10906 8370 10988 8394
rect 1766 8290 1800 8306
rect 1766 7698 1800 7714
rect 2784 8290 2818 8306
rect 2784 7698 2818 7714
rect 3802 8290 3836 8306
rect 3802 7698 3836 7714
rect 4820 8290 4854 8306
rect 4820 7698 4854 7714
rect 5838 8290 5872 8306
rect 5838 7698 5872 7714
rect 6856 8290 6890 8306
rect 6856 7698 6890 7714
rect 7874 8290 7908 8306
rect 7874 7698 7908 7714
rect 8892 8290 8926 8306
rect 8892 7698 8926 7714
rect 9910 8290 9944 8306
rect 9910 7698 9944 7714
rect 10928 8290 10962 8306
rect 13530 8052 13564 8068
rect 14548 8644 14582 8660
rect 14548 8052 14582 8068
rect 15566 8644 15600 8660
rect 15566 8052 15600 8068
rect 16584 8644 16618 8660
rect 16584 8052 16618 8068
rect 17602 8644 17636 8660
rect 17602 8052 17636 8068
rect 18620 8644 18654 8660
rect 18620 8052 18654 8068
rect 19638 8644 19672 8660
rect 19638 8052 19672 8068
rect 20656 8644 20690 8660
rect 20656 8052 20690 8068
rect 21674 8644 21708 8660
rect 21674 8052 21708 8068
rect 22692 8644 22726 8660
rect 22692 8052 22726 8068
rect 23710 8644 23744 8660
rect 23710 8052 23744 8068
rect 24728 8644 24762 8660
rect 24728 8052 24762 8068
rect 25746 8644 25780 8660
rect 25746 8052 25780 8068
rect 26764 8644 26798 8660
rect 26764 8052 26798 8068
rect 27782 8644 27816 8660
rect 27782 8052 27816 8068
rect 28800 8644 28834 8660
rect 28800 8052 28834 8068
rect 29818 8644 29852 8660
rect 29818 8052 29852 8068
rect 30836 8644 30870 8660
rect 30836 8052 30870 8068
rect 31854 8644 31888 8660
rect 31854 8052 31888 8068
rect 32872 8644 32906 8660
rect 32872 8052 32906 8068
rect 33890 8644 33924 8660
rect 33890 8052 33924 8068
rect 22180 8018 22240 8020
rect 24224 8018 24284 8022
rect 32358 8018 32418 8020
rect 13762 7984 13778 8018
rect 14334 7984 14350 8018
rect 14780 7984 14796 8018
rect 15352 7984 15368 8018
rect 15798 7984 15814 8018
rect 16370 7984 16386 8018
rect 16816 7984 16832 8018
rect 17388 7984 17404 8018
rect 17834 7984 17850 8018
rect 18406 7984 18422 8018
rect 18852 7984 18868 8018
rect 19424 7984 19440 8018
rect 19870 7984 19886 8018
rect 20442 7984 20458 8018
rect 20888 7984 20904 8018
rect 21460 7984 21476 8018
rect 21906 7984 21922 8018
rect 22478 7984 22494 8018
rect 22924 7984 22940 8018
rect 23496 7984 23512 8018
rect 23942 7984 23958 8018
rect 24514 7984 24530 8018
rect 24960 7984 24976 8018
rect 25532 7984 25548 8018
rect 25978 7984 25994 8018
rect 26550 7984 26566 8018
rect 26996 7984 27012 8018
rect 27568 7984 27584 8018
rect 28014 7984 28030 8018
rect 28586 7984 28602 8018
rect 29032 7984 29048 8018
rect 29604 7984 29620 8018
rect 30050 7984 30066 8018
rect 30622 7984 30638 8018
rect 31068 7984 31084 8018
rect 31640 7984 31656 8018
rect 32086 7984 32102 8018
rect 32658 7984 32674 8018
rect 33104 7984 33120 8018
rect 33676 7984 33692 8018
rect 10928 7698 10962 7714
rect 14016 7766 14098 7790
rect 14016 7732 14040 7766
rect 14074 7732 14098 7766
rect 14016 7708 14098 7732
rect 15034 7766 15116 7790
rect 15034 7732 15058 7766
rect 15092 7732 15116 7766
rect 15034 7708 15116 7732
rect 16052 7766 16134 7790
rect 16052 7732 16076 7766
rect 16110 7732 16134 7766
rect 16052 7708 16134 7732
rect 17070 7766 17152 7790
rect 17070 7732 17094 7766
rect 17128 7732 17152 7766
rect 17070 7708 17152 7732
rect 18088 7766 18170 7790
rect 18088 7732 18112 7766
rect 18146 7732 18170 7766
rect 18088 7708 18170 7732
rect 19106 7766 19188 7790
rect 19106 7732 19130 7766
rect 19164 7732 19188 7766
rect 19106 7708 19188 7732
rect 20124 7766 20206 7790
rect 20124 7732 20148 7766
rect 20182 7732 20206 7766
rect 20124 7708 20206 7732
rect 21142 7766 21224 7790
rect 21142 7732 21166 7766
rect 21200 7732 21224 7766
rect 21142 7708 21224 7732
rect 22160 7766 22242 7790
rect 22160 7732 22184 7766
rect 22218 7732 22242 7766
rect 22160 7708 22242 7732
rect 23178 7766 23260 7790
rect 23178 7732 23202 7766
rect 23236 7732 23260 7766
rect 23178 7708 23260 7732
rect 24196 7766 24278 7790
rect 24196 7732 24220 7766
rect 24254 7732 24278 7766
rect 24196 7708 24278 7732
rect 25214 7766 25296 7790
rect 25214 7732 25238 7766
rect 25272 7732 25296 7766
rect 25214 7708 25296 7732
rect 26232 7766 26314 7790
rect 26232 7732 26256 7766
rect 26290 7732 26314 7766
rect 26232 7708 26314 7732
rect 27250 7766 27332 7790
rect 27250 7732 27274 7766
rect 27308 7732 27332 7766
rect 27250 7708 27332 7732
rect 28268 7766 28350 7790
rect 28268 7732 28292 7766
rect 28326 7732 28350 7766
rect 28268 7708 28350 7732
rect 29286 7766 29368 7790
rect 29286 7732 29310 7766
rect 29344 7732 29368 7766
rect 29286 7708 29368 7732
rect 30304 7766 30386 7790
rect 30304 7732 30328 7766
rect 30362 7732 30386 7766
rect 30304 7708 30386 7732
rect 31322 7766 31404 7790
rect 31322 7732 31346 7766
rect 31380 7732 31404 7766
rect 31322 7708 31404 7732
rect 32340 7766 32422 7790
rect 32340 7732 32364 7766
rect 32398 7732 32422 7766
rect 32340 7708 32422 7732
rect 33358 7766 33440 7790
rect 33358 7732 33382 7766
rect 33416 7732 33440 7766
rect 33358 7708 33440 7732
rect 1998 7630 2014 7664
rect 2570 7630 2586 7664
rect 3016 7630 3032 7664
rect 3588 7630 3604 7664
rect 4034 7630 4050 7664
rect 4606 7630 4622 7664
rect 5052 7630 5068 7664
rect 5624 7630 5640 7664
rect 6070 7630 6086 7664
rect 6642 7630 6658 7664
rect 7088 7630 7104 7664
rect 7660 7630 7676 7664
rect 8106 7630 8122 7664
rect 8678 7630 8694 7664
rect 9124 7630 9140 7664
rect 9696 7630 9712 7664
rect 10142 7630 10158 7664
rect 10714 7630 10730 7664
rect 13762 7460 13778 7494
rect 14334 7460 14350 7494
rect 14780 7460 14796 7494
rect 15352 7460 15368 7494
rect 15798 7460 15814 7494
rect 16370 7460 16386 7494
rect 16816 7460 16832 7494
rect 17388 7460 17404 7494
rect 17834 7460 17850 7494
rect 18406 7460 18422 7494
rect 18852 7460 18868 7494
rect 19424 7460 19440 7494
rect 19870 7460 19886 7494
rect 20442 7460 20458 7494
rect 20888 7460 20904 7494
rect 21460 7460 21476 7494
rect 21906 7460 21922 7494
rect 22478 7460 22494 7494
rect 22924 7460 22940 7494
rect 23496 7460 23512 7494
rect 23942 7460 23958 7494
rect 24514 7460 24530 7494
rect 24960 7460 24976 7494
rect 25532 7460 25548 7494
rect 25978 7460 25994 7494
rect 26550 7460 26566 7494
rect 26996 7460 27012 7494
rect 27568 7460 27584 7494
rect 28014 7460 28030 7494
rect 28586 7460 28602 7494
rect 29032 7460 29048 7494
rect 29604 7460 29620 7494
rect 30050 7460 30066 7494
rect 30622 7460 30638 7494
rect 31068 7460 31084 7494
rect 31640 7460 31656 7494
rect 32086 7460 32102 7494
rect 32658 7460 32674 7494
rect 33104 7460 33120 7494
rect 33676 7460 33692 7494
rect 13530 7410 13564 7426
rect 2254 7386 2336 7410
rect 2254 7352 2278 7386
rect 2312 7352 2336 7386
rect 2254 7328 2336 7352
rect 3272 7386 3354 7410
rect 3272 7352 3296 7386
rect 3330 7352 3354 7386
rect 3272 7328 3354 7352
rect 4290 7386 4372 7410
rect 4290 7352 4314 7386
rect 4348 7352 4372 7386
rect 4290 7328 4372 7352
rect 5308 7386 5390 7410
rect 5308 7352 5332 7386
rect 5366 7352 5390 7386
rect 5308 7328 5390 7352
rect 6326 7386 6408 7410
rect 6326 7352 6350 7386
rect 6384 7352 6408 7386
rect 6326 7328 6408 7352
rect 7344 7386 7426 7410
rect 7344 7352 7368 7386
rect 7402 7352 7426 7386
rect 7344 7328 7426 7352
rect 8362 7386 8444 7410
rect 8362 7352 8386 7386
rect 8420 7352 8444 7386
rect 8362 7328 8444 7352
rect 9380 7386 9462 7410
rect 9380 7352 9404 7386
rect 9438 7352 9462 7386
rect 9380 7328 9462 7352
rect 10398 7386 10480 7410
rect 10398 7352 10422 7386
rect 10456 7352 10480 7386
rect 10398 7328 10480 7352
rect 8698 6956 8714 6990
rect 8790 6956 8806 6990
rect 8916 6956 8932 6990
rect 9008 6956 9024 6990
rect 9134 6956 9150 6990
rect 9226 6956 9242 6990
rect 9352 6956 9368 6990
rect 9444 6956 9460 6990
rect 9570 6956 9586 6990
rect 9662 6956 9678 6990
rect 9788 6956 9804 6990
rect 9880 6956 9896 6990
rect 10006 6956 10022 6990
rect 10098 6956 10114 6990
rect 10224 6956 10240 6990
rect 10316 6956 10332 6990
rect 10442 6956 10458 6990
rect 10534 6956 10550 6990
rect 10660 6956 10676 6990
rect 10752 6956 10768 6990
rect 8626 6906 8660 6922
rect 8626 6714 8660 6730
rect 8844 6906 8878 6922
rect 8844 6714 8878 6730
rect 9062 6906 9096 6922
rect 9062 6714 9096 6730
rect 9280 6906 9314 6922
rect 9280 6714 9314 6730
rect 9498 6906 9532 6922
rect 9498 6714 9532 6730
rect 9716 6906 9750 6922
rect 9716 6714 9750 6730
rect 9934 6906 9968 6922
rect 9934 6714 9968 6730
rect 10152 6906 10186 6922
rect 10152 6714 10186 6730
rect 10370 6906 10404 6922
rect 10370 6714 10404 6730
rect 10588 6906 10622 6922
rect 10588 6714 10622 6730
rect 10806 6906 10840 6922
rect 13530 6818 13564 6834
rect 14548 7410 14582 7426
rect 14548 6818 14582 6834
rect 15566 7410 15600 7426
rect 15566 6818 15600 6834
rect 16584 7410 16618 7426
rect 16584 6818 16618 6834
rect 17602 7410 17636 7426
rect 17602 6818 17636 6834
rect 18620 7410 18654 7426
rect 18620 6818 18654 6834
rect 19638 7410 19672 7426
rect 19638 6818 19672 6834
rect 20656 7410 20690 7426
rect 20656 6818 20690 6834
rect 21674 7410 21708 7426
rect 21674 6818 21708 6834
rect 22692 7410 22726 7426
rect 22692 6818 22726 6834
rect 23710 7410 23744 7426
rect 23710 6818 23744 6834
rect 24728 7410 24762 7426
rect 24728 6818 24762 6834
rect 25746 7410 25780 7426
rect 25746 6818 25780 6834
rect 26764 7410 26798 7426
rect 26764 6818 26798 6834
rect 27782 7410 27816 7426
rect 27782 6818 27816 6834
rect 28800 7410 28834 7426
rect 28800 6818 28834 6834
rect 29818 7410 29852 7426
rect 29818 6818 29852 6834
rect 30836 7410 30870 7426
rect 30836 6818 30870 6834
rect 31854 7410 31888 7426
rect 31854 6818 31888 6834
rect 32872 7410 32906 7426
rect 32872 6818 32906 6834
rect 33890 7410 33924 7426
rect 33890 6818 33924 6834
rect 16056 6784 16116 6788
rect 13762 6750 13778 6784
rect 14334 6750 14350 6784
rect 14780 6750 14796 6784
rect 15352 6750 15368 6784
rect 15798 6750 15814 6784
rect 16370 6750 16386 6784
rect 16816 6750 16832 6784
rect 17388 6750 17404 6784
rect 17834 6750 17850 6784
rect 18406 6750 18422 6784
rect 18852 6750 18868 6784
rect 19424 6750 19440 6784
rect 19870 6750 19886 6784
rect 20442 6750 20458 6784
rect 20888 6750 20904 6784
rect 21460 6750 21476 6784
rect 21906 6750 21922 6784
rect 22478 6750 22494 6784
rect 22924 6750 22940 6784
rect 23496 6750 23512 6784
rect 23942 6750 23958 6784
rect 24514 6750 24530 6784
rect 24960 6750 24976 6784
rect 25532 6750 25548 6784
rect 25978 6750 25994 6784
rect 26550 6750 26566 6784
rect 26996 6750 27012 6784
rect 27568 6750 27584 6784
rect 28014 6750 28030 6784
rect 28586 6750 28602 6784
rect 29032 6750 29048 6784
rect 29604 6750 29620 6784
rect 30050 6750 30066 6784
rect 30622 6750 30638 6784
rect 31068 6750 31084 6784
rect 31640 6750 31656 6784
rect 32086 6750 32102 6784
rect 32658 6750 32674 6784
rect 33104 6750 33120 6784
rect 33676 6750 33692 6784
rect 10806 6714 10840 6730
rect 8698 6646 8714 6680
rect 8790 6646 8806 6680
rect 8916 6646 8932 6680
rect 9008 6646 9024 6680
rect 9134 6646 9150 6680
rect 9226 6646 9242 6680
rect 9352 6646 9368 6680
rect 9444 6646 9460 6680
rect 9570 6646 9586 6680
rect 9662 6646 9678 6680
rect 9788 6646 9804 6680
rect 9880 6646 9896 6680
rect 10006 6646 10022 6680
rect 10098 6646 10114 6680
rect 10224 6646 10240 6680
rect 10316 6646 10332 6680
rect 10442 6646 10458 6680
rect 10534 6646 10550 6680
rect 10660 6646 10676 6680
rect 10752 6646 10768 6680
rect 14016 6518 14098 6542
rect 14016 6484 14040 6518
rect 14074 6484 14098 6518
rect 14016 6460 14098 6484
rect 15034 6518 15116 6542
rect 15034 6484 15058 6518
rect 15092 6484 15116 6518
rect 15034 6460 15116 6484
rect 16052 6518 16134 6542
rect 16052 6484 16076 6518
rect 16110 6484 16134 6518
rect 16052 6460 16134 6484
rect 17070 6518 17152 6542
rect 17070 6484 17094 6518
rect 17128 6484 17152 6518
rect 17070 6460 17152 6484
rect 18088 6518 18170 6542
rect 18088 6484 18112 6518
rect 18146 6484 18170 6518
rect 18088 6460 18170 6484
rect 19106 6518 19188 6542
rect 19106 6484 19130 6518
rect 19164 6484 19188 6518
rect 19106 6460 19188 6484
rect 20124 6518 20206 6542
rect 20124 6484 20148 6518
rect 20182 6484 20206 6518
rect 20124 6460 20206 6484
rect 21142 6518 21224 6542
rect 21142 6484 21166 6518
rect 21200 6484 21224 6518
rect 21142 6460 21224 6484
rect 22160 6518 22242 6542
rect 22160 6484 22184 6518
rect 22218 6484 22242 6518
rect 22160 6460 22242 6484
rect 23178 6518 23260 6542
rect 23178 6484 23202 6518
rect 23236 6484 23260 6518
rect 23178 6460 23260 6484
rect 24196 6518 24278 6542
rect 24196 6484 24220 6518
rect 24254 6484 24278 6518
rect 24196 6460 24278 6484
rect 25214 6518 25296 6542
rect 25214 6484 25238 6518
rect 25272 6484 25296 6518
rect 25214 6460 25296 6484
rect 26232 6518 26314 6542
rect 26232 6484 26256 6518
rect 26290 6484 26314 6518
rect 26232 6460 26314 6484
rect 27250 6518 27332 6542
rect 27250 6484 27274 6518
rect 27308 6484 27332 6518
rect 27250 6460 27332 6484
rect 28268 6518 28350 6542
rect 28268 6484 28292 6518
rect 28326 6484 28350 6518
rect 28268 6460 28350 6484
rect 29286 6518 29368 6542
rect 29286 6484 29310 6518
rect 29344 6484 29368 6518
rect 29286 6460 29368 6484
rect 30304 6518 30386 6542
rect 30304 6484 30328 6518
rect 30362 6484 30386 6518
rect 30304 6460 30386 6484
rect 31322 6518 31404 6542
rect 31322 6484 31346 6518
rect 31380 6484 31404 6518
rect 31322 6460 31404 6484
rect 32340 6518 32422 6542
rect 32340 6484 32364 6518
rect 32398 6484 32422 6518
rect 32340 6460 32422 6484
rect 33358 6518 33440 6542
rect 33358 6484 33382 6518
rect 33416 6484 33440 6518
rect 33358 6460 33440 6484
rect 8332 6410 8414 6434
rect 8332 6376 8356 6410
rect 8390 6376 8414 6410
rect 8332 6352 8414 6376
rect 9350 6410 9432 6434
rect 9350 6376 9374 6410
rect 9408 6376 9432 6410
rect 9350 6352 9432 6376
rect 10368 6410 10450 6434
rect 10368 6376 10392 6410
rect 10426 6376 10450 6410
rect 10368 6352 10450 6376
rect 11386 6410 11468 6434
rect 11386 6376 11410 6410
rect 11444 6376 11468 6410
rect 11386 6352 11468 6376
rect 13762 6226 13778 6260
rect 14334 6226 14350 6260
rect 14780 6226 14796 6260
rect 15352 6226 15368 6260
rect 15798 6226 15814 6260
rect 16370 6226 16386 6260
rect 16816 6226 16832 6260
rect 17388 6226 17404 6260
rect 17834 6226 17850 6260
rect 18406 6226 18422 6260
rect 18852 6226 18868 6260
rect 19424 6226 19440 6260
rect 19870 6226 19886 6260
rect 20442 6226 20458 6260
rect 20888 6226 20904 6260
rect 21460 6226 21476 6260
rect 21906 6226 21922 6260
rect 22478 6226 22494 6260
rect 22924 6226 22940 6260
rect 23496 6226 23512 6260
rect 23942 6226 23958 6260
rect 24514 6226 24530 6260
rect 24960 6226 24976 6260
rect 25532 6226 25548 6260
rect 25978 6226 25994 6260
rect 26550 6226 26566 6260
rect 26996 6226 27012 6260
rect 27568 6226 27584 6260
rect 28014 6226 28030 6260
rect 28586 6226 28602 6260
rect 29032 6226 29048 6260
rect 29604 6226 29620 6260
rect 30050 6226 30066 6260
rect 30622 6226 30638 6260
rect 31068 6226 31084 6260
rect 31640 6226 31656 6260
rect 32086 6226 32102 6260
rect 32658 6226 32674 6260
rect 33104 6226 33120 6260
rect 33676 6226 33692 6260
rect 13530 6176 13564 6192
rect 8698 6124 8714 6158
rect 8790 6124 8806 6158
rect 8916 6124 8932 6158
rect 9008 6124 9024 6158
rect 9134 6124 9150 6158
rect 9226 6124 9242 6158
rect 9352 6124 9368 6158
rect 9444 6124 9460 6158
rect 9570 6124 9586 6158
rect 9662 6124 9678 6158
rect 9788 6124 9804 6158
rect 9880 6124 9896 6158
rect 10006 6124 10022 6158
rect 10098 6124 10114 6158
rect 10224 6124 10240 6158
rect 10316 6124 10332 6158
rect 10442 6124 10458 6158
rect 10534 6124 10550 6158
rect 10660 6124 10676 6158
rect 10752 6124 10768 6158
rect 8626 6074 8660 6090
rect 8626 5882 8660 5898
rect 8844 6074 8878 6090
rect 8844 5882 8878 5898
rect 9062 6074 9096 6090
rect 9062 5882 9096 5898
rect 9280 6074 9314 6090
rect 9280 5882 9314 5898
rect 9498 6074 9532 6090
rect 9498 5882 9532 5898
rect 9716 6074 9750 6090
rect 9716 5882 9750 5898
rect 9934 6074 9968 6090
rect 9934 5882 9968 5898
rect 10152 6074 10186 6090
rect 10152 5882 10186 5898
rect 10370 6074 10404 6090
rect 10370 5882 10404 5898
rect 10588 6074 10622 6090
rect 10588 5882 10622 5898
rect 10806 6074 10840 6090
rect 10806 5882 10840 5898
rect 8698 5814 8714 5848
rect 8790 5814 8806 5848
rect 8916 5814 8932 5848
rect 9008 5814 9024 5848
rect 9134 5814 9150 5848
rect 9226 5814 9242 5848
rect 9352 5814 9368 5848
rect 9444 5814 9460 5848
rect 9570 5814 9586 5848
rect 9662 5814 9678 5848
rect 9788 5814 9804 5848
rect 9880 5814 9896 5848
rect 10006 5814 10022 5848
rect 10098 5814 10114 5848
rect 10224 5814 10240 5848
rect 10316 5814 10332 5848
rect 10442 5814 10458 5848
rect 10534 5814 10550 5848
rect 10660 5814 10676 5848
rect 10752 5814 10768 5848
rect 13530 5584 13564 5600
rect 14548 6176 14582 6192
rect 14548 5584 14582 5600
rect 15566 6176 15600 6192
rect 15566 5584 15600 5600
rect 16584 6176 16618 6192
rect 16584 5584 16618 5600
rect 17602 6176 17636 6192
rect 17602 5584 17636 5600
rect 18620 6176 18654 6192
rect 18620 5584 18654 5600
rect 19638 6176 19672 6192
rect 19638 5584 19672 5600
rect 20656 6176 20690 6192
rect 20656 5584 20690 5600
rect 21674 6176 21708 6192
rect 21674 5584 21708 5600
rect 22692 6176 22726 6192
rect 22692 5584 22726 5600
rect 23710 6176 23744 6192
rect 23710 5584 23744 5600
rect 24728 6176 24762 6192
rect 24728 5584 24762 5600
rect 25746 6176 25780 6192
rect 25746 5584 25780 5600
rect 26764 6176 26798 6192
rect 26764 5584 26798 5600
rect 27782 6176 27816 6192
rect 27782 5584 27816 5600
rect 28800 6176 28834 6192
rect 28800 5584 28834 5600
rect 29818 6176 29852 6192
rect 29818 5584 29852 5600
rect 30836 6176 30870 6192
rect 30836 5584 30870 5600
rect 31854 6176 31888 6192
rect 31854 5584 31888 5600
rect 32872 6176 32906 6192
rect 32872 5584 32906 5600
rect 33890 6176 33924 6192
rect 33890 5584 33924 5600
rect 22180 5550 22240 5552
rect 24224 5550 24284 5554
rect 27262 5550 27322 5554
rect 13762 5516 13778 5550
rect 14334 5516 14350 5550
rect 14780 5516 14796 5550
rect 15352 5516 15368 5550
rect 15798 5516 15814 5550
rect 16370 5516 16386 5550
rect 16816 5516 16832 5550
rect 17388 5516 17404 5550
rect 17834 5516 17850 5550
rect 18406 5516 18422 5550
rect 18852 5516 18868 5550
rect 19424 5516 19440 5550
rect 19870 5516 19886 5550
rect 20442 5516 20458 5550
rect 20888 5516 20904 5550
rect 21460 5516 21476 5550
rect 21906 5516 21922 5550
rect 22478 5516 22494 5550
rect 22924 5516 22940 5550
rect 23496 5516 23512 5550
rect 23942 5516 23958 5550
rect 24514 5516 24530 5550
rect 24960 5516 24976 5550
rect 25532 5516 25548 5550
rect 25978 5516 25994 5550
rect 26550 5516 26566 5550
rect 26996 5516 27012 5550
rect 27568 5516 27584 5550
rect 28014 5516 28030 5550
rect 28586 5516 28602 5550
rect 29032 5516 29048 5550
rect 29604 5516 29620 5550
rect 30050 5516 30066 5550
rect 30622 5516 30638 5550
rect 31068 5516 31084 5550
rect 31640 5516 31656 5550
rect 32086 5516 32102 5550
rect 32658 5516 32674 5550
rect 33104 5516 33120 5550
rect 33676 5516 33692 5550
rect 14030 5298 14112 5322
rect 14030 5264 14054 5298
rect 14088 5264 14112 5298
rect 14030 5240 14112 5264
rect 15048 5298 15130 5322
rect 15048 5264 15072 5298
rect 15106 5264 15130 5298
rect 15048 5240 15130 5264
rect 16066 5298 16148 5322
rect 16066 5264 16090 5298
rect 16124 5264 16148 5298
rect 16066 5240 16148 5264
rect 17084 5298 17166 5322
rect 17084 5264 17108 5298
rect 17142 5264 17166 5298
rect 17084 5240 17166 5264
rect 18102 5298 18184 5322
rect 18102 5264 18126 5298
rect 18160 5264 18184 5298
rect 18102 5240 18184 5264
rect 19120 5298 19202 5322
rect 19120 5264 19144 5298
rect 19178 5264 19202 5298
rect 19120 5240 19202 5264
rect 20138 5298 20220 5322
rect 20138 5264 20162 5298
rect 20196 5264 20220 5298
rect 20138 5240 20220 5264
rect 21156 5298 21238 5322
rect 21156 5264 21180 5298
rect 21214 5264 21238 5298
rect 21156 5240 21238 5264
rect 22174 5298 22256 5322
rect 22174 5264 22198 5298
rect 22232 5264 22256 5298
rect 22174 5240 22256 5264
rect 23192 5298 23274 5322
rect 23192 5264 23216 5298
rect 23250 5264 23274 5298
rect 23192 5240 23274 5264
rect 24210 5298 24292 5322
rect 24210 5264 24234 5298
rect 24268 5264 24292 5298
rect 24210 5240 24292 5264
rect 25228 5298 25310 5322
rect 25228 5264 25252 5298
rect 25286 5264 25310 5298
rect 25228 5240 25310 5264
rect 26246 5298 26328 5322
rect 26246 5264 26270 5298
rect 26304 5264 26328 5298
rect 26246 5240 26328 5264
rect 27264 5298 27346 5322
rect 27264 5264 27288 5298
rect 27322 5264 27346 5298
rect 27264 5240 27346 5264
rect 28282 5298 28364 5322
rect 28282 5264 28306 5298
rect 28340 5264 28364 5298
rect 28282 5240 28364 5264
rect 29300 5298 29382 5322
rect 29300 5264 29324 5298
rect 29358 5264 29382 5298
rect 29300 5240 29382 5264
rect 30318 5298 30400 5322
rect 30318 5264 30342 5298
rect 30376 5264 30400 5298
rect 30318 5240 30400 5264
rect 31336 5298 31418 5322
rect 31336 5264 31360 5298
rect 31394 5264 31418 5298
rect 31336 5240 31418 5264
rect 32354 5298 32436 5322
rect 32354 5264 32378 5298
rect 32412 5264 32436 5298
rect 32354 5240 32436 5264
rect 33372 5298 33454 5322
rect 33372 5264 33396 5298
rect 33430 5264 33454 5298
rect 33372 5240 33454 5264
rect 8630 5122 8712 5146
rect 2038 5066 2120 5090
rect 2038 5032 2062 5066
rect 2096 5032 2120 5066
rect 2038 5008 2120 5032
rect 3056 5066 3138 5090
rect 3056 5032 3080 5066
rect 3114 5032 3138 5066
rect 3056 5008 3138 5032
rect 4074 5066 4156 5090
rect 4074 5032 4098 5066
rect 4132 5032 4156 5066
rect 4074 5008 4156 5032
rect 5092 5066 5174 5090
rect 5092 5032 5116 5066
rect 5150 5032 5174 5066
rect 5092 5008 5174 5032
rect 6110 5066 6192 5090
rect 6110 5032 6134 5066
rect 6168 5032 6192 5066
rect 6110 5008 6192 5032
rect 7128 5066 7210 5090
rect 7128 5032 7152 5066
rect 7186 5032 7210 5066
rect 8630 5088 8654 5122
rect 8688 5088 8712 5122
rect 8630 5064 8712 5088
rect 9648 5122 9730 5146
rect 9648 5088 9672 5122
rect 9706 5088 9730 5122
rect 9648 5064 9730 5088
rect 10666 5122 10748 5146
rect 10666 5088 10690 5122
rect 10724 5088 10748 5122
rect 10666 5064 10748 5088
rect 11684 5122 11766 5146
rect 11684 5088 11708 5122
rect 11742 5088 11766 5122
rect 11684 5064 11766 5088
rect 7128 5008 7210 5032
rect 13762 4994 13778 5028
rect 14334 4994 14350 5028
rect 14780 4994 14796 5028
rect 15352 4994 15368 5028
rect 15798 4994 15814 5028
rect 16370 4994 16386 5028
rect 16816 4994 16832 5028
rect 17388 4994 17404 5028
rect 17834 4994 17850 5028
rect 18406 4994 18422 5028
rect 18852 4994 18868 5028
rect 19424 4994 19440 5028
rect 19870 4994 19886 5028
rect 20442 4994 20458 5028
rect 20888 4994 20904 5028
rect 21460 4994 21476 5028
rect 21906 4994 21922 5028
rect 22478 4994 22494 5028
rect 22924 4994 22940 5028
rect 23496 4994 23512 5028
rect 23942 4994 23958 5028
rect 24514 4994 24530 5028
rect 24960 4994 24976 5028
rect 25532 4994 25548 5028
rect 25978 4994 25994 5028
rect 26550 4994 26566 5028
rect 26996 4994 27012 5028
rect 27568 4994 27584 5028
rect 28014 4994 28030 5028
rect 28586 4994 28602 5028
rect 29032 4994 29048 5028
rect 29604 4994 29620 5028
rect 30050 4994 30066 5028
rect 30622 4994 30638 5028
rect 31068 4994 31084 5028
rect 31640 4994 31656 5028
rect 32086 4994 32102 5028
rect 32658 4994 32674 5028
rect 33104 4994 33120 5028
rect 33676 4994 33692 5028
rect 17084 4992 17144 4994
rect 13530 4944 13564 4960
rect 1777 4797 1793 4831
rect 2349 4797 2365 4831
rect 2795 4797 2811 4831
rect 3367 4797 3383 4831
rect 3813 4797 3829 4831
rect 4385 4797 4401 4831
rect 4831 4797 4847 4831
rect 5403 4797 5419 4831
rect 5849 4797 5865 4831
rect 6421 4797 6437 4831
rect 6867 4797 6883 4831
rect 7439 4797 7455 4831
rect 8628 4798 8644 4832
rect 8768 4798 8784 4832
rect 8926 4798 8942 4832
rect 9066 4798 9082 4832
rect 9224 4798 9240 4832
rect 9364 4798 9380 4832
rect 9522 4798 9538 4832
rect 9662 4798 9678 4832
rect 9820 4798 9836 4832
rect 9960 4798 9976 4832
rect 10118 4798 10134 4832
rect 10258 4798 10274 4832
rect 10416 4798 10432 4832
rect 10556 4798 10572 4832
rect 10714 4798 10730 4832
rect 10854 4798 10870 4832
rect 11012 4798 11028 4832
rect 11152 4798 11168 4832
rect 11310 4798 11326 4832
rect 11450 4798 11466 4832
rect 11608 4798 11624 4832
rect 11748 4798 11764 4832
rect 1545 4747 1579 4763
rect 1545 4155 1579 4171
rect 2563 4747 2597 4763
rect 2563 4155 2597 4171
rect 3581 4747 3615 4763
rect 3581 4155 3615 4171
rect 4599 4747 4633 4763
rect 4599 4155 4633 4171
rect 5617 4747 5651 4763
rect 5617 4155 5651 4171
rect 6635 4747 6669 4763
rect 6635 4155 6669 4171
rect 7653 4747 7687 4763
rect 7653 4155 7687 4171
rect 8540 4748 8574 4764
rect 8540 4156 8574 4172
rect 8838 4748 8872 4764
rect 8838 4156 8872 4172
rect 9136 4748 9170 4764
rect 9136 4156 9170 4172
rect 9434 4748 9468 4764
rect 9434 4156 9468 4172
rect 9732 4748 9766 4764
rect 9732 4156 9766 4172
rect 10030 4748 10064 4764
rect 10030 4156 10064 4172
rect 10328 4748 10362 4764
rect 10328 4156 10362 4172
rect 10626 4748 10660 4764
rect 10626 4156 10660 4172
rect 10924 4748 10958 4764
rect 10924 4156 10958 4172
rect 11222 4748 11256 4764
rect 11222 4156 11256 4172
rect 11520 4748 11554 4764
rect 11520 4156 11554 4172
rect 11818 4748 11852 4764
rect 13530 4352 13564 4368
rect 14548 4944 14582 4960
rect 14548 4352 14582 4368
rect 15566 4944 15600 4960
rect 15566 4352 15600 4368
rect 16584 4944 16618 4960
rect 16584 4352 16618 4368
rect 17602 4944 17636 4960
rect 17602 4352 17636 4368
rect 18620 4944 18654 4960
rect 18620 4352 18654 4368
rect 19638 4944 19672 4960
rect 19638 4352 19672 4368
rect 20656 4944 20690 4960
rect 20656 4352 20690 4368
rect 21674 4944 21708 4960
rect 21674 4352 21708 4368
rect 22692 4944 22726 4960
rect 22692 4352 22726 4368
rect 23710 4944 23744 4960
rect 23710 4352 23744 4368
rect 24728 4944 24762 4960
rect 24728 4352 24762 4368
rect 25746 4944 25780 4960
rect 25746 4352 25780 4368
rect 26764 4944 26798 4960
rect 26764 4352 26798 4368
rect 27782 4944 27816 4960
rect 27782 4352 27816 4368
rect 28800 4944 28834 4960
rect 28800 4352 28834 4368
rect 29818 4944 29852 4960
rect 29818 4352 29852 4368
rect 30836 4944 30870 4960
rect 30836 4352 30870 4368
rect 31854 4944 31888 4960
rect 31854 4352 31888 4368
rect 32872 4944 32906 4960
rect 32872 4352 32906 4368
rect 33890 4944 33924 4960
rect 33890 4352 33924 4368
rect 21156 4318 21216 4328
rect 13762 4284 13778 4318
rect 14334 4284 14350 4318
rect 14780 4284 14796 4318
rect 15352 4284 15368 4318
rect 15798 4284 15814 4318
rect 16370 4284 16386 4318
rect 16816 4284 16832 4318
rect 17388 4284 17404 4318
rect 17834 4284 17850 4318
rect 18406 4284 18422 4318
rect 18852 4284 18868 4318
rect 19424 4284 19440 4318
rect 19870 4284 19886 4318
rect 20442 4284 20458 4318
rect 20888 4284 20904 4318
rect 21460 4284 21476 4318
rect 21906 4284 21922 4318
rect 22478 4284 22494 4318
rect 22924 4284 22940 4318
rect 23496 4284 23512 4318
rect 23942 4284 23958 4318
rect 24514 4284 24530 4318
rect 24960 4284 24976 4318
rect 25532 4284 25548 4318
rect 25978 4284 25994 4318
rect 26550 4284 26566 4318
rect 26996 4284 27012 4318
rect 27568 4284 27584 4318
rect 28014 4284 28030 4318
rect 28586 4284 28602 4318
rect 29032 4284 29048 4318
rect 29604 4284 29620 4318
rect 30050 4284 30066 4318
rect 30622 4284 30638 4318
rect 31068 4284 31084 4318
rect 31640 4284 31656 4318
rect 32086 4284 32102 4318
rect 32658 4284 32674 4318
rect 33104 4284 33120 4318
rect 33676 4284 33692 4318
rect 11818 4156 11852 4172
rect 3058 4121 3118 4122
rect 4068 4121 4128 4122
rect 6116 4121 6176 4122
rect 1777 4087 1793 4121
rect 2349 4087 2365 4121
rect 2795 4087 2811 4121
rect 3367 4087 3383 4121
rect 3813 4087 3829 4121
rect 4385 4087 4401 4121
rect 4831 4087 4847 4121
rect 5403 4087 5419 4121
rect 5849 4087 5865 4121
rect 6421 4087 6437 4121
rect 6867 4087 6883 4121
rect 7439 4087 7455 4121
rect 8628 4088 8644 4122
rect 8768 4088 8784 4122
rect 8926 4088 8942 4122
rect 9066 4088 9082 4122
rect 9224 4088 9240 4122
rect 9364 4088 9380 4122
rect 9522 4088 9538 4122
rect 9662 4088 9678 4122
rect 9820 4088 9836 4122
rect 9960 4088 9976 4122
rect 10118 4088 10134 4122
rect 10258 4088 10274 4122
rect 10416 4088 10432 4122
rect 10556 4088 10572 4122
rect 10714 4088 10730 4122
rect 10854 4088 10870 4122
rect 11012 4088 11028 4122
rect 11152 4088 11168 4122
rect 11310 4088 11326 4122
rect 11450 4088 11466 4122
rect 11608 4088 11624 4122
rect 11748 4088 11764 4122
rect 8976 4068 9036 4088
rect 14030 4050 14112 4074
rect 14030 4016 14054 4050
rect 14088 4016 14112 4050
rect 14030 3992 14112 4016
rect 15048 4050 15130 4074
rect 15048 4016 15072 4050
rect 15106 4016 15130 4050
rect 15048 3992 15130 4016
rect 16066 4050 16148 4074
rect 16066 4016 16090 4050
rect 16124 4016 16148 4050
rect 16066 3992 16148 4016
rect 17084 4050 17166 4074
rect 17084 4016 17108 4050
rect 17142 4016 17166 4050
rect 17084 3992 17166 4016
rect 18102 4050 18184 4074
rect 18102 4016 18126 4050
rect 18160 4016 18184 4050
rect 18102 3992 18184 4016
rect 19120 4050 19202 4074
rect 19120 4016 19144 4050
rect 19178 4016 19202 4050
rect 19120 3992 19202 4016
rect 20138 4050 20220 4074
rect 20138 4016 20162 4050
rect 20196 4016 20220 4050
rect 20138 3992 20220 4016
rect 21156 4050 21238 4074
rect 21156 4016 21180 4050
rect 21214 4016 21238 4050
rect 21156 3992 21238 4016
rect 22174 4050 22256 4074
rect 22174 4016 22198 4050
rect 22232 4016 22256 4050
rect 22174 3992 22256 4016
rect 23192 4050 23274 4074
rect 23192 4016 23216 4050
rect 23250 4016 23274 4050
rect 23192 3992 23274 4016
rect 24210 4050 24292 4074
rect 24210 4016 24234 4050
rect 24268 4016 24292 4050
rect 24210 3992 24292 4016
rect 25228 4050 25310 4074
rect 25228 4016 25252 4050
rect 25286 4016 25310 4050
rect 25228 3992 25310 4016
rect 26246 4050 26328 4074
rect 26246 4016 26270 4050
rect 26304 4016 26328 4050
rect 26246 3992 26328 4016
rect 27264 4050 27346 4074
rect 27264 4016 27288 4050
rect 27322 4016 27346 4050
rect 27264 3992 27346 4016
rect 28282 4050 28364 4074
rect 28282 4016 28306 4050
rect 28340 4016 28364 4050
rect 28282 3992 28364 4016
rect 29300 4050 29382 4074
rect 29300 4016 29324 4050
rect 29358 4016 29382 4050
rect 29300 3992 29382 4016
rect 30318 4050 30400 4074
rect 30318 4016 30342 4050
rect 30376 4016 30400 4050
rect 30318 3992 30400 4016
rect 31336 4050 31418 4074
rect 31336 4016 31360 4050
rect 31394 4016 31418 4050
rect 31336 3992 31418 4016
rect 32354 4050 32436 4074
rect 32354 4016 32378 4050
rect 32412 4016 32436 4050
rect 32354 3992 32436 4016
rect 33372 4050 33454 4074
rect 33372 4016 33396 4050
rect 33430 4016 33454 4050
rect 33372 3992 33454 4016
rect 2052 3940 2134 3964
rect 2052 3906 2076 3940
rect 2110 3906 2134 3940
rect 2052 3882 2134 3906
rect 3070 3940 3152 3964
rect 3070 3906 3094 3940
rect 3128 3906 3152 3940
rect 3070 3882 3152 3906
rect 4088 3940 4170 3964
rect 4088 3906 4112 3940
rect 4146 3906 4170 3940
rect 4088 3882 4170 3906
rect 5106 3940 5188 3964
rect 5106 3906 5130 3940
rect 5164 3906 5188 3940
rect 5106 3882 5188 3906
rect 6124 3940 6206 3964
rect 6124 3906 6148 3940
rect 6182 3906 6206 3940
rect 6124 3882 6206 3906
rect 7142 3940 7224 3964
rect 7142 3906 7166 3940
rect 7200 3906 7224 3940
rect 7142 3882 7224 3906
rect 8590 3928 8672 3952
rect 8590 3894 8614 3928
rect 8648 3894 8672 3928
rect 8590 3870 8672 3894
rect 9608 3928 9690 3952
rect 9608 3894 9632 3928
rect 9666 3894 9690 3928
rect 9608 3870 9690 3894
rect 10626 3928 10708 3952
rect 10626 3894 10650 3928
rect 10684 3894 10708 3928
rect 10626 3870 10708 3894
rect 11644 3928 11726 3952
rect 11644 3894 11668 3928
rect 11702 3894 11726 3928
rect 11644 3870 11726 3894
rect 13762 3760 13778 3794
rect 14334 3760 14350 3794
rect 14780 3760 14796 3794
rect 15352 3760 15368 3794
rect 15798 3760 15814 3794
rect 16370 3760 16386 3794
rect 16816 3760 16832 3794
rect 17388 3760 17404 3794
rect 17834 3760 17850 3794
rect 18406 3760 18422 3794
rect 18852 3760 18868 3794
rect 19424 3760 19440 3794
rect 19870 3760 19886 3794
rect 20442 3760 20458 3794
rect 20888 3760 20904 3794
rect 21460 3760 21476 3794
rect 21906 3760 21922 3794
rect 22478 3760 22494 3794
rect 22924 3760 22940 3794
rect 23496 3760 23512 3794
rect 23942 3760 23958 3794
rect 24514 3760 24530 3794
rect 24960 3760 24976 3794
rect 25532 3760 25548 3794
rect 25978 3760 25994 3794
rect 26550 3760 26566 3794
rect 26996 3760 27012 3794
rect 27568 3760 27584 3794
rect 28014 3760 28030 3794
rect 28586 3760 28602 3794
rect 29032 3760 29048 3794
rect 29604 3760 29620 3794
rect 30050 3760 30066 3794
rect 30622 3760 30638 3794
rect 31068 3760 31084 3794
rect 31640 3760 31656 3794
rect 32086 3760 32102 3794
rect 32658 3760 32674 3794
rect 33104 3760 33120 3794
rect 33676 3760 33692 3794
rect 17070 3758 17130 3760
rect 1776 3684 1792 3718
rect 2348 3684 2364 3718
rect 2794 3684 2810 3718
rect 3366 3684 3382 3718
rect 3812 3684 3828 3718
rect 4384 3684 4400 3718
rect 4830 3684 4846 3718
rect 5402 3684 5418 3718
rect 5848 3684 5864 3718
rect 6420 3684 6436 3718
rect 6866 3684 6882 3718
rect 7438 3684 7454 3718
rect 8628 3686 8644 3720
rect 8768 3686 8784 3720
rect 8926 3686 8942 3720
rect 9066 3686 9082 3720
rect 9224 3686 9240 3720
rect 9364 3686 9380 3720
rect 9522 3686 9538 3720
rect 9662 3686 9678 3720
rect 9820 3686 9836 3720
rect 9960 3686 9976 3720
rect 10118 3686 10134 3720
rect 10258 3686 10274 3720
rect 10416 3686 10432 3720
rect 10556 3686 10572 3720
rect 10714 3686 10730 3720
rect 10854 3686 10870 3720
rect 11012 3686 11028 3720
rect 11152 3686 11168 3720
rect 11310 3686 11326 3720
rect 11450 3686 11466 3720
rect 11608 3686 11624 3720
rect 11748 3686 11764 3720
rect 13530 3710 13564 3726
rect 3058 3682 3118 3684
rect 5094 3682 5154 3684
rect 6116 3682 6176 3684
rect 1544 3634 1578 3650
rect 1544 3042 1578 3058
rect 2562 3634 2596 3650
rect 2562 3042 2596 3058
rect 3580 3634 3614 3650
rect 3580 3042 3614 3058
rect 4598 3634 4632 3650
rect 4598 3042 4632 3058
rect 5616 3634 5650 3650
rect 5616 3042 5650 3058
rect 6634 3634 6668 3650
rect 6634 3042 6668 3058
rect 7652 3634 7686 3650
rect 7652 3042 7686 3058
rect 8540 3636 8574 3652
rect 8540 3044 8574 3060
rect 8838 3636 8872 3652
rect 8838 3044 8872 3060
rect 9136 3636 9170 3652
rect 9136 3044 9170 3060
rect 9434 3636 9468 3652
rect 9434 3044 9468 3060
rect 9732 3636 9766 3652
rect 9732 3044 9766 3060
rect 10030 3636 10064 3652
rect 10030 3044 10064 3060
rect 10328 3636 10362 3652
rect 10328 3044 10362 3060
rect 10626 3636 10660 3652
rect 10626 3044 10660 3060
rect 10924 3636 10958 3652
rect 10924 3044 10958 3060
rect 11222 3636 11256 3652
rect 11222 3044 11256 3060
rect 11520 3636 11554 3652
rect 11520 3044 11554 3060
rect 11818 3636 11852 3652
rect 13530 3118 13564 3134
rect 14548 3710 14582 3726
rect 14548 3118 14582 3134
rect 15566 3710 15600 3726
rect 15566 3118 15600 3134
rect 16584 3710 16618 3726
rect 16584 3118 16618 3134
rect 17602 3710 17636 3726
rect 17602 3118 17636 3134
rect 18620 3710 18654 3726
rect 18620 3118 18654 3134
rect 19638 3710 19672 3726
rect 19638 3118 19672 3134
rect 20656 3710 20690 3726
rect 20656 3118 20690 3134
rect 21674 3710 21708 3726
rect 21674 3118 21708 3134
rect 22692 3710 22726 3726
rect 22692 3118 22726 3134
rect 23710 3710 23744 3726
rect 23710 3118 23744 3134
rect 24728 3710 24762 3726
rect 24728 3118 24762 3134
rect 25746 3710 25780 3726
rect 25746 3118 25780 3134
rect 26764 3710 26798 3726
rect 26764 3118 26798 3134
rect 27782 3710 27816 3726
rect 27782 3118 27816 3134
rect 28800 3710 28834 3726
rect 28800 3118 28834 3134
rect 29818 3710 29852 3726
rect 29818 3118 29852 3134
rect 30836 3710 30870 3726
rect 30836 3118 30870 3134
rect 31854 3710 31888 3726
rect 31854 3118 31888 3134
rect 32872 3710 32906 3726
rect 32872 3118 32906 3134
rect 33890 3710 33924 3726
rect 33890 3118 33924 3134
rect 15038 3084 15098 3086
rect 21150 3084 21210 3086
rect 23184 3084 23244 3086
rect 27250 3084 27310 3090
rect 31326 3084 31386 3086
rect 32342 3084 32402 3086
rect 11818 3044 11852 3060
rect 13762 3050 13778 3084
rect 14334 3050 14350 3084
rect 14780 3050 14796 3084
rect 15352 3050 15368 3084
rect 15798 3050 15814 3084
rect 16370 3050 16386 3084
rect 16816 3050 16832 3084
rect 17388 3050 17404 3084
rect 17834 3050 17850 3084
rect 18406 3050 18422 3084
rect 18852 3050 18868 3084
rect 19424 3050 19440 3084
rect 19870 3050 19886 3084
rect 20442 3050 20458 3084
rect 20888 3050 20904 3084
rect 21460 3050 21476 3084
rect 21906 3050 21922 3084
rect 22478 3050 22494 3084
rect 22924 3050 22940 3084
rect 23496 3050 23512 3084
rect 23942 3050 23958 3084
rect 24514 3050 24530 3084
rect 24960 3050 24976 3084
rect 25532 3050 25548 3084
rect 25978 3050 25994 3084
rect 26550 3050 26566 3084
rect 26996 3050 27012 3084
rect 27568 3050 27584 3084
rect 28014 3050 28030 3084
rect 28586 3050 28602 3084
rect 29032 3050 29048 3084
rect 29604 3050 29620 3084
rect 30050 3050 30066 3084
rect 30622 3050 30638 3084
rect 31068 3050 31084 3084
rect 31640 3050 31656 3084
rect 32086 3050 32102 3084
rect 32658 3050 32674 3084
rect 33104 3050 33120 3084
rect 33676 3050 33692 3084
rect 3060 3008 3120 3012
rect 4070 3008 4130 3012
rect 6118 3008 6178 3012
rect 1776 2974 1792 3008
rect 2348 2974 2364 3008
rect 2794 2974 2810 3008
rect 3366 2974 3382 3008
rect 3812 2974 3828 3008
rect 4384 2974 4400 3008
rect 4830 2974 4846 3008
rect 5402 2974 5418 3008
rect 5848 2974 5864 3008
rect 6420 2974 6436 3008
rect 6866 2974 6882 3008
rect 7438 2974 7454 3008
rect 8628 2976 8644 3010
rect 8768 2976 8784 3010
rect 8926 2976 8942 3010
rect 9066 2976 9082 3010
rect 9224 2976 9240 3010
rect 9364 2976 9380 3010
rect 9522 2976 9538 3010
rect 9662 2976 9678 3010
rect 9820 2976 9836 3010
rect 9960 2976 9976 3010
rect 10118 2976 10134 3010
rect 10258 2976 10274 3010
rect 10416 2976 10432 3010
rect 10556 2976 10572 3010
rect 10714 2976 10730 3010
rect 10854 2976 10870 3010
rect 11012 2976 11028 3010
rect 11152 2976 11168 3010
rect 11310 2976 11326 3010
rect 11450 2976 11466 3010
rect 11608 2976 11624 3010
rect 11748 2976 11764 3010
rect 2026 2814 2108 2838
rect 2026 2780 2050 2814
rect 2084 2780 2108 2814
rect 2026 2756 2108 2780
rect 3044 2814 3126 2838
rect 3044 2780 3068 2814
rect 3102 2780 3126 2814
rect 3044 2756 3126 2780
rect 4062 2814 4144 2838
rect 4062 2780 4086 2814
rect 4120 2780 4144 2814
rect 4062 2756 4144 2780
rect 5080 2814 5162 2838
rect 5080 2780 5104 2814
rect 5138 2780 5162 2814
rect 5080 2756 5162 2780
rect 6098 2814 6180 2838
rect 6098 2780 6122 2814
rect 6156 2780 6180 2814
rect 6098 2756 6180 2780
rect 7116 2814 7198 2838
rect 7116 2780 7140 2814
rect 7174 2780 7198 2814
rect 7116 2756 7198 2780
rect 8590 2814 8672 2838
rect 8590 2780 8614 2814
rect 8648 2780 8672 2814
rect 8590 2756 8672 2780
rect 9608 2814 9690 2838
rect 9608 2780 9632 2814
rect 9666 2780 9690 2814
rect 9608 2756 9690 2780
rect 10626 2814 10708 2838
rect 10626 2780 10650 2814
rect 10684 2780 10708 2814
rect 10626 2756 10708 2780
rect 11644 2814 11726 2838
rect 11644 2780 11668 2814
rect 11702 2780 11726 2814
rect 11644 2756 11726 2780
rect 14016 2828 14098 2852
rect 14016 2794 14040 2828
rect 14074 2794 14098 2828
rect 14016 2770 14098 2794
rect 15034 2828 15116 2852
rect 15034 2794 15058 2828
rect 15092 2794 15116 2828
rect 15034 2770 15116 2794
rect 16052 2828 16134 2852
rect 16052 2794 16076 2828
rect 16110 2794 16134 2828
rect 16052 2770 16134 2794
rect 17070 2828 17152 2852
rect 17070 2794 17094 2828
rect 17128 2794 17152 2828
rect 17070 2770 17152 2794
rect 18088 2828 18170 2852
rect 18088 2794 18112 2828
rect 18146 2794 18170 2828
rect 18088 2770 18170 2794
rect 19106 2828 19188 2852
rect 19106 2794 19130 2828
rect 19164 2794 19188 2828
rect 19106 2770 19188 2794
rect 20124 2828 20206 2852
rect 20124 2794 20148 2828
rect 20182 2794 20206 2828
rect 20124 2770 20206 2794
rect 21142 2828 21224 2852
rect 21142 2794 21166 2828
rect 21200 2794 21224 2828
rect 21142 2770 21224 2794
rect 22160 2828 22242 2852
rect 22160 2794 22184 2828
rect 22218 2794 22242 2828
rect 22160 2770 22242 2794
rect 23178 2828 23260 2852
rect 23178 2794 23202 2828
rect 23236 2794 23260 2828
rect 23178 2770 23260 2794
rect 24196 2828 24278 2852
rect 24196 2794 24220 2828
rect 24254 2794 24278 2828
rect 24196 2770 24278 2794
rect 25214 2828 25296 2852
rect 25214 2794 25238 2828
rect 25272 2794 25296 2828
rect 25214 2770 25296 2794
rect 26232 2828 26314 2852
rect 26232 2794 26256 2828
rect 26290 2794 26314 2828
rect 26232 2770 26314 2794
rect 27250 2828 27332 2852
rect 27250 2794 27274 2828
rect 27308 2794 27332 2828
rect 27250 2770 27332 2794
rect 28268 2828 28350 2852
rect 28268 2794 28292 2828
rect 28326 2794 28350 2828
rect 28268 2770 28350 2794
rect 29286 2828 29368 2852
rect 29286 2794 29310 2828
rect 29344 2794 29368 2828
rect 29286 2770 29368 2794
rect 30304 2828 30386 2852
rect 30304 2794 30328 2828
rect 30362 2794 30386 2828
rect 30304 2770 30386 2794
rect 31322 2828 31404 2852
rect 31322 2794 31346 2828
rect 31380 2794 31404 2828
rect 31322 2770 31404 2794
rect 32340 2828 32422 2852
rect 32340 2794 32364 2828
rect 32398 2794 32422 2828
rect 32340 2770 32422 2794
rect 33358 2828 33440 2852
rect 33358 2794 33382 2828
rect 33416 2794 33440 2828
rect 33358 2770 33440 2794
rect 1777 2573 1793 2607
rect 2349 2573 2365 2607
rect 2795 2573 2811 2607
rect 3367 2573 3383 2607
rect 3813 2573 3829 2607
rect 4385 2573 4401 2607
rect 4831 2573 4847 2607
rect 5403 2573 5419 2607
rect 5849 2573 5865 2607
rect 6421 2573 6437 2607
rect 6867 2573 6883 2607
rect 7439 2573 7455 2607
rect 8626 2574 8642 2608
rect 8766 2574 8782 2608
rect 8924 2574 8940 2608
rect 9064 2574 9080 2608
rect 9222 2574 9238 2608
rect 9362 2574 9378 2608
rect 9520 2574 9536 2608
rect 9660 2574 9676 2608
rect 9818 2574 9834 2608
rect 9958 2574 9974 2608
rect 10116 2574 10132 2608
rect 10256 2574 10272 2608
rect 10414 2574 10430 2608
rect 10554 2574 10570 2608
rect 10712 2574 10728 2608
rect 10852 2574 10868 2608
rect 11010 2574 11026 2608
rect 11150 2574 11166 2608
rect 11308 2574 11324 2608
rect 11448 2574 11464 2608
rect 11606 2574 11622 2608
rect 11746 2574 11762 2608
rect 3060 2572 3120 2573
rect 5096 2572 5156 2573
rect 6118 2572 6178 2573
rect 1545 2523 1579 2539
rect 1545 1931 1579 1947
rect 2563 2523 2597 2539
rect 2563 1931 2597 1947
rect 3581 2523 3615 2539
rect 3581 1931 3615 1947
rect 4599 2523 4633 2539
rect 4599 1931 4633 1947
rect 5617 2523 5651 2539
rect 5617 1931 5651 1947
rect 6635 2523 6669 2539
rect 6635 1931 6669 1947
rect 7653 2523 7687 2539
rect 7653 1931 7687 1947
rect 8538 2524 8572 2540
rect 8538 1932 8572 1948
rect 8836 2524 8870 2540
rect 8836 1932 8870 1948
rect 9134 2524 9168 2540
rect 9134 1932 9168 1948
rect 9432 2524 9466 2540
rect 9432 1932 9466 1948
rect 9730 2524 9764 2540
rect 9730 1932 9764 1948
rect 10028 2524 10062 2540
rect 10028 1932 10062 1948
rect 10326 2524 10360 2540
rect 10326 1932 10360 1948
rect 10624 2524 10658 2540
rect 10624 1932 10658 1948
rect 10922 2524 10956 2540
rect 10922 1932 10956 1948
rect 11220 2524 11254 2540
rect 11220 1932 11254 1948
rect 11518 2524 11552 2540
rect 11518 1932 11552 1948
rect 11816 2524 11850 2540
rect 13762 2526 13778 2560
rect 14334 2526 14350 2560
rect 14780 2526 14796 2560
rect 15352 2526 15368 2560
rect 15798 2526 15814 2560
rect 16370 2526 16386 2560
rect 16816 2526 16832 2560
rect 17388 2526 17404 2560
rect 17834 2526 17850 2560
rect 18406 2526 18422 2560
rect 18852 2526 18868 2560
rect 19424 2526 19440 2560
rect 19870 2526 19886 2560
rect 20442 2526 20458 2560
rect 20888 2526 20904 2560
rect 21460 2526 21476 2560
rect 21906 2526 21922 2560
rect 22478 2526 22494 2560
rect 22924 2526 22940 2560
rect 23496 2526 23512 2560
rect 23942 2526 23958 2560
rect 24514 2526 24530 2560
rect 24960 2526 24976 2560
rect 25532 2526 25548 2560
rect 25978 2526 25994 2560
rect 26550 2526 26566 2560
rect 26996 2526 27012 2560
rect 27568 2526 27584 2560
rect 28014 2526 28030 2560
rect 28586 2526 28602 2560
rect 29032 2526 29048 2560
rect 29604 2526 29620 2560
rect 30050 2526 30066 2560
rect 30622 2526 30638 2560
rect 31068 2526 31084 2560
rect 31640 2526 31656 2560
rect 32086 2526 32102 2560
rect 32658 2526 32674 2560
rect 33104 2526 33120 2560
rect 33676 2526 33692 2560
rect 20148 2520 20208 2526
rect 25220 2520 25280 2526
rect 26240 2520 26300 2526
rect 28276 2520 28336 2526
rect 11816 1932 11850 1948
rect 13530 2476 13564 2492
rect 3062 1897 3122 1902
rect 4072 1897 4132 1902
rect 5098 1897 5158 1898
rect 6120 1897 6180 1902
rect 1777 1863 1793 1897
rect 2349 1863 2365 1897
rect 2795 1863 2811 1897
rect 3367 1863 3383 1897
rect 3813 1863 3829 1897
rect 4385 1863 4401 1897
rect 4831 1863 4847 1897
rect 5403 1863 5419 1897
rect 5849 1863 5865 1897
rect 6421 1863 6437 1897
rect 6867 1863 6883 1897
rect 7439 1863 7455 1897
rect 8626 1864 8642 1898
rect 8766 1864 8782 1898
rect 8924 1864 8940 1898
rect 9064 1864 9080 1898
rect 9222 1864 9238 1898
rect 9362 1864 9378 1898
rect 9520 1864 9536 1898
rect 9660 1864 9676 1898
rect 9818 1864 9834 1898
rect 9958 1864 9974 1898
rect 10116 1864 10132 1898
rect 10256 1864 10272 1898
rect 10414 1864 10430 1898
rect 10554 1864 10570 1898
rect 10712 1864 10728 1898
rect 10852 1864 10868 1898
rect 11010 1864 11026 1898
rect 11150 1864 11166 1898
rect 11308 1864 11324 1898
rect 11448 1864 11464 1898
rect 11606 1864 11622 1898
rect 11746 1864 11762 1898
rect 13530 1884 13564 1900
rect 14548 2476 14582 2492
rect 14548 1884 14582 1900
rect 15566 2476 15600 2492
rect 15566 1884 15600 1900
rect 16584 2476 16618 2492
rect 16584 1884 16618 1900
rect 17602 2476 17636 2492
rect 17602 1884 17636 1900
rect 18620 2476 18654 2492
rect 18620 1884 18654 1900
rect 19638 2476 19672 2492
rect 19638 1884 19672 1900
rect 20656 2476 20690 2492
rect 20656 1884 20690 1900
rect 21674 2476 21708 2492
rect 21674 1884 21708 1900
rect 22692 2476 22726 2492
rect 22692 1884 22726 1900
rect 23710 2476 23744 2492
rect 23710 1884 23744 1900
rect 24728 2476 24762 2492
rect 24728 1884 24762 1900
rect 25746 2476 25780 2492
rect 25746 1884 25780 1900
rect 26764 2476 26798 2492
rect 26764 1884 26798 1900
rect 27782 2476 27816 2492
rect 27782 1884 27816 1900
rect 28800 2476 28834 2492
rect 28800 1884 28834 1900
rect 29818 2476 29852 2492
rect 29818 1884 29852 1900
rect 30836 2476 30870 2492
rect 30836 1884 30870 1900
rect 31854 2476 31888 2492
rect 31854 1884 31888 1900
rect 32872 2476 32906 2492
rect 32872 1884 32906 1900
rect 33890 2476 33924 2492
rect 33890 1884 33924 1900
rect 24204 1850 24264 1856
rect 13762 1816 13778 1850
rect 14334 1816 14350 1850
rect 14780 1816 14796 1850
rect 15352 1816 15368 1850
rect 15798 1816 15814 1850
rect 16370 1816 16386 1850
rect 16816 1816 16832 1850
rect 17388 1816 17404 1850
rect 17834 1816 17850 1850
rect 18406 1816 18422 1850
rect 18852 1816 18868 1850
rect 19424 1816 19440 1850
rect 19870 1816 19886 1850
rect 20442 1816 20458 1850
rect 20888 1816 20904 1850
rect 21460 1816 21476 1850
rect 21906 1816 21922 1850
rect 22478 1816 22494 1850
rect 22924 1816 22940 1850
rect 23496 1816 23512 1850
rect 23942 1816 23958 1850
rect 24514 1816 24530 1850
rect 24960 1816 24976 1850
rect 25532 1816 25548 1850
rect 25978 1816 25994 1850
rect 26550 1816 26566 1850
rect 26996 1816 27012 1850
rect 27568 1816 27584 1850
rect 28014 1816 28030 1850
rect 28586 1816 28602 1850
rect 29032 1816 29048 1850
rect 29604 1816 29620 1850
rect 30050 1816 30066 1850
rect 30622 1816 30638 1850
rect 31068 1816 31084 1850
rect 31640 1816 31656 1850
rect 32086 1816 32102 1850
rect 32658 1816 32674 1850
rect 33104 1816 33120 1850
rect 33676 1816 33692 1850
rect 2052 1716 2134 1740
rect 2052 1682 2076 1716
rect 2110 1682 2134 1716
rect 2052 1658 2134 1682
rect 3070 1716 3152 1740
rect 3070 1682 3094 1716
rect 3128 1682 3152 1716
rect 3070 1658 3152 1682
rect 4088 1716 4170 1740
rect 4088 1682 4112 1716
rect 4146 1682 4170 1716
rect 4088 1658 4170 1682
rect 5106 1716 5188 1740
rect 5106 1682 5130 1716
rect 5164 1682 5188 1716
rect 5106 1658 5188 1682
rect 6124 1716 6206 1740
rect 6124 1682 6148 1716
rect 6182 1682 6206 1716
rect 6124 1658 6206 1682
rect 7142 1716 7224 1740
rect 7142 1682 7166 1716
rect 7200 1682 7224 1716
rect 7142 1658 7224 1682
rect 8644 1702 8726 1726
rect 8644 1668 8668 1702
rect 8702 1668 8726 1702
rect 8644 1644 8726 1668
rect 9662 1702 9744 1726
rect 9662 1668 9686 1702
rect 9720 1668 9744 1702
rect 9662 1644 9744 1668
rect 10680 1702 10762 1726
rect 10680 1668 10704 1702
rect 10738 1668 10762 1702
rect 10680 1644 10762 1668
rect 11698 1702 11780 1726
rect 11698 1668 11722 1702
rect 11756 1668 11780 1702
rect 11698 1644 11780 1668
rect 14016 1608 14098 1632
rect 14016 1574 14040 1608
rect 14074 1574 14098 1608
rect 14016 1550 14098 1574
rect 15034 1608 15116 1632
rect 15034 1574 15058 1608
rect 15092 1574 15116 1608
rect 15034 1550 15116 1574
rect 16052 1608 16134 1632
rect 16052 1574 16076 1608
rect 16110 1574 16134 1608
rect 16052 1550 16134 1574
rect 17070 1608 17152 1632
rect 17070 1574 17094 1608
rect 17128 1574 17152 1608
rect 17070 1550 17152 1574
rect 18088 1608 18170 1632
rect 18088 1574 18112 1608
rect 18146 1574 18170 1608
rect 18088 1550 18170 1574
rect 19106 1608 19188 1632
rect 19106 1574 19130 1608
rect 19164 1574 19188 1608
rect 19106 1550 19188 1574
rect 20124 1608 20206 1632
rect 20124 1574 20148 1608
rect 20182 1574 20206 1608
rect 20124 1550 20206 1574
rect 21142 1608 21224 1632
rect 21142 1574 21166 1608
rect 21200 1574 21224 1608
rect 21142 1550 21224 1574
rect 22160 1608 22242 1632
rect 22160 1574 22184 1608
rect 22218 1574 22242 1608
rect 22160 1550 22242 1574
rect 23178 1608 23260 1632
rect 23178 1574 23202 1608
rect 23236 1574 23260 1608
rect 23178 1550 23260 1574
rect 24196 1608 24278 1632
rect 24196 1574 24220 1608
rect 24254 1574 24278 1608
rect 24196 1550 24278 1574
rect 25214 1608 25296 1632
rect 25214 1574 25238 1608
rect 25272 1574 25296 1608
rect 25214 1550 25296 1574
rect 26232 1608 26314 1632
rect 26232 1574 26256 1608
rect 26290 1574 26314 1608
rect 26232 1550 26314 1574
rect 27250 1608 27332 1632
rect 27250 1574 27274 1608
rect 27308 1574 27332 1608
rect 27250 1550 27332 1574
rect 28268 1608 28350 1632
rect 28268 1574 28292 1608
rect 28326 1574 28350 1608
rect 28268 1550 28350 1574
rect 29286 1608 29368 1632
rect 29286 1574 29310 1608
rect 29344 1574 29368 1608
rect 29286 1550 29368 1574
rect 30304 1608 30386 1632
rect 30304 1574 30328 1608
rect 30362 1574 30386 1608
rect 30304 1550 30386 1574
rect 31322 1608 31404 1632
rect 31322 1574 31346 1608
rect 31380 1574 31404 1608
rect 31322 1550 31404 1574
rect 32340 1608 32422 1632
rect 32340 1574 32364 1608
rect 32398 1574 32422 1608
rect 32340 1550 32422 1574
rect 33358 1608 33440 1632
rect 33358 1574 33382 1608
rect 33416 1574 33440 1608
rect 33358 1550 33440 1574
rect 1776 1460 1792 1494
rect 2348 1460 2364 1494
rect 2794 1460 2810 1494
rect 3366 1460 3382 1494
rect 3812 1460 3828 1494
rect 4384 1460 4400 1494
rect 4830 1460 4846 1494
rect 5402 1460 5418 1494
rect 5848 1460 5864 1494
rect 6420 1460 6436 1494
rect 6866 1460 6882 1494
rect 7438 1460 7454 1494
rect 8626 1464 8642 1498
rect 8766 1464 8782 1498
rect 8924 1464 8940 1498
rect 9064 1464 9080 1498
rect 9222 1464 9238 1498
rect 9362 1464 9378 1498
rect 9520 1464 9536 1498
rect 9660 1464 9676 1498
rect 9818 1464 9834 1498
rect 9958 1464 9974 1498
rect 10116 1464 10132 1498
rect 10256 1464 10272 1498
rect 10414 1464 10430 1498
rect 10554 1464 10570 1498
rect 10712 1464 10728 1498
rect 10852 1464 10868 1498
rect 11010 1464 11026 1498
rect 11150 1464 11166 1498
rect 11308 1464 11324 1498
rect 11448 1464 11464 1498
rect 11606 1464 11622 1498
rect 11746 1464 11762 1498
rect 1544 1410 1578 1426
rect 1544 818 1578 834
rect 2562 1410 2596 1426
rect 2562 818 2596 834
rect 3580 1410 3614 1426
rect 3580 818 3614 834
rect 4598 1410 4632 1426
rect 4598 818 4632 834
rect 5616 1410 5650 1426
rect 5616 818 5650 834
rect 6634 1410 6668 1426
rect 6634 818 6668 834
rect 7652 1410 7686 1426
rect 7652 818 7686 834
rect 8538 1414 8572 1430
rect 8538 822 8572 838
rect 8836 1414 8870 1430
rect 8836 822 8870 838
rect 9134 1414 9168 1430
rect 9134 822 9168 838
rect 9432 1414 9466 1430
rect 9432 822 9466 838
rect 9730 1414 9764 1430
rect 9730 822 9764 838
rect 10028 1414 10062 1430
rect 10028 822 10062 838
rect 10326 1414 10360 1430
rect 10326 822 10360 838
rect 10624 1414 10658 1430
rect 10624 822 10658 838
rect 10922 1414 10956 1430
rect 10922 822 10956 838
rect 11220 1414 11254 1430
rect 11220 822 11254 838
rect 11518 1414 11552 1430
rect 11518 822 11552 838
rect 11816 1414 11850 1430
rect 13762 1294 13778 1328
rect 14334 1294 14350 1328
rect 14780 1294 14796 1328
rect 15352 1294 15368 1328
rect 15798 1294 15814 1328
rect 16370 1294 16386 1328
rect 16816 1294 16832 1328
rect 17388 1294 17404 1328
rect 17834 1294 17850 1328
rect 18406 1294 18422 1328
rect 18852 1294 18868 1328
rect 19424 1294 19440 1328
rect 19870 1294 19886 1328
rect 20442 1294 20458 1328
rect 20888 1294 20904 1328
rect 21460 1294 21476 1328
rect 21906 1294 21922 1328
rect 22478 1294 22494 1328
rect 22924 1294 22940 1328
rect 23496 1294 23512 1328
rect 23942 1294 23958 1328
rect 24514 1294 24530 1328
rect 24960 1294 24976 1328
rect 25532 1294 25548 1328
rect 25978 1294 25994 1328
rect 26550 1294 26566 1328
rect 26996 1294 27012 1328
rect 27568 1294 27584 1328
rect 28014 1294 28030 1328
rect 28586 1294 28602 1328
rect 29032 1294 29048 1328
rect 29604 1294 29620 1328
rect 30050 1294 30066 1328
rect 30622 1294 30638 1328
rect 31068 1294 31084 1328
rect 31640 1294 31656 1328
rect 32086 1294 32102 1328
rect 32658 1294 32674 1328
rect 33104 1294 33120 1328
rect 33676 1294 33692 1328
rect 14016 1290 14076 1294
rect 15038 1290 15098 1294
rect 16064 1290 16124 1294
rect 17080 1290 17140 1294
rect 18094 1290 18154 1294
rect 19124 1284 19184 1294
rect 20140 1284 20200 1294
rect 21144 1290 21204 1294
rect 22174 1284 22234 1294
rect 23194 1290 23254 1294
rect 24204 1290 24264 1294
rect 25228 1284 25288 1294
rect 27254 1290 27314 1294
rect 28274 1284 28334 1294
rect 29298 1290 29358 1294
rect 32342 1290 32402 1294
rect 33364 1292 33424 1294
rect 11816 822 11850 838
rect 13530 1244 13564 1260
rect 1776 750 1792 784
rect 2348 750 2364 784
rect 2794 750 2810 784
rect 3366 750 3382 784
rect 3812 750 3828 784
rect 4384 750 4400 784
rect 4830 750 4846 784
rect 5402 750 5418 784
rect 5848 750 5864 784
rect 6420 750 6436 784
rect 6866 750 6882 784
rect 7438 750 7454 784
rect 8626 754 8642 788
rect 8766 754 8782 788
rect 8924 754 8940 788
rect 9064 754 9080 788
rect 9222 754 9238 788
rect 9362 754 9378 788
rect 9520 754 9536 788
rect 9660 754 9676 788
rect 9818 754 9834 788
rect 9958 754 9974 788
rect 10116 754 10132 788
rect 10256 754 10272 788
rect 10414 754 10430 788
rect 10554 754 10570 788
rect 10712 754 10728 788
rect 10852 754 10868 788
rect 11010 754 11026 788
rect 11150 754 11166 788
rect 11308 754 11324 788
rect 11448 754 11464 788
rect 11606 754 11622 788
rect 11746 754 11762 788
rect 14548 1244 14582 1260
rect 14532 668 14548 708
rect 15566 1244 15600 1260
rect 14582 668 14592 708
rect 13530 652 13564 668
rect 14548 652 14582 668
rect 15566 652 15600 668
rect 16584 1244 16618 1260
rect 16584 652 16618 668
rect 17602 1244 17636 1260
rect 18620 1244 18654 1260
rect 18606 668 18620 712
rect 19638 1244 19672 1260
rect 18654 668 18666 712
rect 17602 652 17636 668
rect 18620 652 18654 668
rect 19638 652 19672 668
rect 20656 1244 20690 1260
rect 20656 652 20690 668
rect 21674 1244 21708 1260
rect 21674 652 21708 668
rect 22692 1244 22726 1260
rect 22692 652 22726 668
rect 23710 1244 23744 1260
rect 24728 1244 24762 1260
rect 24714 668 24728 714
rect 25746 1244 25780 1260
rect 24762 668 24774 714
rect 23710 652 23744 668
rect 24728 652 24762 668
rect 25746 652 25780 668
rect 26764 1244 26798 1260
rect 26764 652 26798 668
rect 27782 1244 27816 1260
rect 28800 1244 28834 1260
rect 28786 668 28800 704
rect 29818 1244 29852 1260
rect 28834 668 28846 704
rect 27782 652 27816 668
rect 28800 652 28834 668
rect 29818 652 29852 668
rect 30836 1244 30870 1260
rect 30836 652 30870 668
rect 31854 1244 31888 1260
rect 32872 1244 32906 1260
rect 32856 668 32872 706
rect 33890 1244 33924 1260
rect 32906 668 32916 706
rect 31854 652 31888 668
rect 32872 652 32906 668
rect 33890 652 33924 668
rect 20136 618 20196 620
rect 26248 618 26308 620
rect 31334 618 31394 620
rect 13762 584 13778 618
rect 14334 584 14350 618
rect 14780 584 14796 618
rect 15352 584 15368 618
rect 15798 584 15814 618
rect 16370 584 16386 618
rect 16816 584 16832 618
rect 17388 584 17404 618
rect 17834 584 17850 618
rect 18406 584 18422 618
rect 18852 584 18868 618
rect 19424 584 19440 618
rect 19870 584 19886 618
rect 20442 584 20458 618
rect 20888 584 20904 618
rect 21460 584 21476 618
rect 21906 584 21922 618
rect 22478 584 22494 618
rect 22924 584 22940 618
rect 23496 584 23512 618
rect 23942 584 23958 618
rect 24514 584 24530 618
rect 24960 584 24976 618
rect 25532 584 25548 618
rect 25978 584 25994 618
rect 26550 584 26566 618
rect 26996 584 27012 618
rect 27568 584 27584 618
rect 28014 584 28030 618
rect 28586 584 28602 618
rect 29032 584 29048 618
rect 29604 584 29620 618
rect 30050 584 30066 618
rect 30622 584 30638 618
rect 31068 584 31084 618
rect 31640 584 31656 618
rect 32086 584 32102 618
rect 32658 584 32674 618
rect 33104 584 33120 618
rect 33676 584 33692 618
rect 2026 522 2108 546
rect 2026 488 2050 522
rect 2084 488 2108 522
rect 2026 464 2108 488
rect 3044 522 3126 546
rect 3044 488 3068 522
rect 3102 488 3126 522
rect 3044 464 3126 488
rect 4062 522 4144 546
rect 4062 488 4086 522
rect 4120 488 4144 522
rect 4062 464 4144 488
rect 5080 522 5162 546
rect 5080 488 5104 522
rect 5138 488 5162 522
rect 5080 464 5162 488
rect 6098 522 6180 546
rect 6098 488 6122 522
rect 6156 488 6180 522
rect 6098 464 6180 488
rect 7116 522 7198 546
rect 7116 488 7140 522
rect 7174 488 7198 522
rect 7116 464 7198 488
rect 8618 468 8700 492
rect 8618 434 8642 468
rect 8676 434 8700 468
rect 8618 410 8700 434
rect 9636 468 9718 492
rect 9636 434 9660 468
rect 9694 434 9718 468
rect 9636 410 9718 434
rect 10654 468 10736 492
rect 10654 434 10678 468
rect 10712 434 10736 468
rect 10654 410 10736 434
rect 11672 468 11754 492
rect 11672 434 11696 468
rect 11730 434 11754 468
rect 11672 410 11754 434
rect -1372 -682 -1272 -520
rect 52628 15200 52728 15362
rect 89772 15200 89872 15362
rect 67764 14860 67780 14894
rect 68336 14860 68352 14894
rect 68782 14860 68798 14894
rect 69354 14860 69370 14894
rect 69800 14860 69816 14894
rect 70372 14860 70388 14894
rect 70818 14860 70834 14894
rect 71390 14860 71406 14894
rect 71836 14860 71852 14894
rect 72408 14860 72424 14894
rect 72854 14860 72870 14894
rect 73426 14860 73442 14894
rect 73872 14860 73888 14894
rect 74444 14860 74460 14894
rect 74890 14860 74906 14894
rect 75462 14860 75478 14894
rect 75908 14860 75924 14894
rect 76480 14860 76496 14894
rect 76926 14860 76942 14894
rect 77498 14860 77514 14894
rect 77944 14860 77960 14894
rect 78516 14860 78532 14894
rect 78962 14860 78978 14894
rect 79534 14860 79550 14894
rect 79980 14860 79996 14894
rect 80552 14860 80568 14894
rect 80998 14860 81014 14894
rect 81570 14860 81586 14894
rect 82016 14860 82032 14894
rect 82588 14860 82604 14894
rect 83034 14860 83050 14894
rect 83606 14860 83622 14894
rect 84052 14860 84068 14894
rect 84624 14860 84640 14894
rect 85070 14860 85086 14894
rect 85642 14860 85658 14894
rect 86088 14860 86104 14894
rect 86660 14860 86676 14894
rect 87106 14860 87122 14894
rect 87678 14860 87694 14894
rect 48690 8414 48736 8447
rect 50430 8414 50500 8447
rect 48690 8413 48786 8414
rect 50404 8413 50500 8414
rect 48690 8351 48724 8413
rect 50466 8352 50500 8413
rect 48884 8311 48900 8345
rect 49000 8311 49016 8345
rect 49142 8311 49158 8345
rect 49258 8311 49274 8345
rect 49400 8311 49416 8345
rect 49516 8311 49532 8345
rect 49658 8311 49674 8345
rect 49774 8311 49790 8345
rect 49916 8311 49932 8345
rect 50032 8311 50048 8345
rect 50174 8311 50190 8345
rect 50290 8311 50306 8345
rect 48804 8252 48838 8268
rect 48804 7860 48838 7876
rect 49062 8252 49096 8268
rect 49062 7860 49096 7876
rect 49320 8252 49354 8268
rect 49320 7860 49354 7876
rect 49578 8252 49612 8268
rect 49578 7860 49612 7876
rect 49836 8252 49870 8268
rect 49836 7860 49870 7876
rect 50094 8252 50128 8268
rect 50094 7860 50128 7876
rect 50352 8252 50386 8268
rect 50352 7860 50386 7876
rect 48884 7783 48900 7817
rect 49000 7783 49016 7817
rect 49142 7783 49158 7817
rect 49258 7783 49274 7817
rect 49400 7783 49416 7817
rect 49516 7783 49532 7817
rect 49658 7783 49674 7817
rect 49774 7783 49790 7817
rect 49916 7783 49932 7817
rect 50032 7783 50048 7817
rect 50174 7783 50190 7817
rect 50290 7783 50306 7817
rect 48690 7715 48724 7777
rect 50574 7911 50603 7945
rect 50637 7911 50695 7945
rect 50729 7911 50787 7945
rect 50821 7911 50850 7945
rect 50466 7715 50500 7776
rect 48690 7714 48786 7715
rect 48690 7681 48736 7714
rect 50430 7682 50500 7715
rect 50404 7681 50500 7682
rect 50640 7869 50706 7877
rect 50640 7835 50656 7869
rect 50690 7835 50706 7869
rect 50640 7801 50706 7835
rect 50640 7767 50656 7801
rect 50690 7767 50706 7801
rect 50640 7733 50706 7767
rect 50640 7699 50656 7733
rect 50690 7699 50706 7733
rect 50640 7681 50706 7699
rect 50740 7869 50782 7911
rect 50774 7835 50782 7869
rect 50740 7801 50782 7835
rect 50774 7767 50782 7801
rect 50740 7733 50782 7767
rect 50774 7699 50782 7733
rect 50740 7683 50782 7699
rect 50640 7622 50686 7681
rect 50681 7574 50686 7622
rect 50720 7644 50786 7647
rect 50720 7633 50737 7644
rect 50720 7599 50736 7633
rect 50783 7604 50786 7644
rect 50770 7599 50786 7604
rect 50640 7561 50686 7574
rect 50640 7549 50706 7561
rect 50640 7515 50656 7549
rect 50690 7515 50706 7549
rect 48690 7480 48760 7514
rect 50430 7480 50500 7514
rect 48690 7418 48724 7480
rect 50466 7418 50500 7480
rect 50640 7481 50706 7515
rect 50640 7447 50656 7481
rect 50690 7447 50706 7481
rect 50640 7435 50706 7447
rect 50740 7549 50786 7565
rect 50774 7515 50786 7549
rect 50740 7481 50786 7515
rect 50774 7447 50786 7481
rect 48884 7378 48900 7412
rect 49000 7378 49016 7412
rect 49142 7378 49158 7412
rect 49258 7378 49274 7412
rect 49400 7378 49416 7412
rect 49516 7378 49532 7412
rect 49658 7378 49674 7412
rect 49774 7378 49790 7412
rect 49916 7378 49932 7412
rect 50032 7378 50048 7412
rect 50174 7378 50190 7412
rect 50290 7378 50306 7412
rect 48804 7328 48838 7344
rect 48804 7136 48838 7152
rect 49062 7328 49096 7344
rect 49062 7136 49096 7152
rect 49320 7328 49354 7344
rect 49320 7136 49354 7152
rect 49578 7328 49612 7344
rect 49578 7136 49612 7152
rect 49836 7328 49870 7344
rect 49836 7136 49870 7152
rect 50094 7328 50128 7344
rect 50094 7136 50128 7152
rect 50352 7328 50386 7344
rect 50352 7136 50386 7152
rect 48884 7068 48900 7102
rect 49000 7068 49016 7102
rect 49142 7068 49158 7102
rect 49258 7068 49274 7102
rect 49400 7068 49416 7102
rect 49516 7068 49532 7102
rect 49658 7068 49674 7102
rect 49774 7068 49790 7102
rect 49916 7068 49932 7102
rect 50032 7068 50048 7102
rect 50174 7068 50190 7102
rect 50290 7068 50306 7102
rect 50740 7401 50786 7447
rect 50574 7367 50603 7401
rect 50637 7367 50695 7401
rect 50729 7367 50787 7401
rect 50821 7367 50850 7401
rect 48690 7000 48724 7062
rect 50466 7000 50500 7062
rect 48690 6966 48758 7000
rect 50432 6966 50500 7000
rect 48690 6450 48736 6483
rect 50430 6450 50500 6483
rect 48690 6449 48786 6450
rect 50404 6449 50500 6450
rect 48690 6387 48724 6449
rect 50466 6388 50500 6449
rect 48884 6347 48900 6381
rect 49000 6347 49016 6381
rect 49142 6347 49158 6381
rect 49258 6347 49274 6381
rect 49400 6347 49416 6381
rect 49516 6347 49532 6381
rect 49658 6347 49674 6381
rect 49774 6347 49790 6381
rect 49916 6347 49932 6381
rect 50032 6347 50048 6381
rect 50174 6347 50190 6381
rect 50290 6347 50306 6381
rect 48804 6288 48838 6304
rect 48804 5896 48838 5912
rect 49062 6288 49096 6304
rect 49062 5896 49096 5912
rect 49320 6288 49354 6304
rect 49320 5896 49354 5912
rect 49578 6288 49612 6304
rect 49578 5896 49612 5912
rect 49836 6288 49870 6304
rect 49836 5896 49870 5912
rect 50094 6288 50128 6304
rect 50094 5896 50128 5912
rect 50352 6288 50386 6304
rect 50352 5896 50386 5912
rect 48884 5819 48900 5853
rect 49000 5819 49016 5853
rect 49142 5819 49158 5853
rect 49258 5819 49274 5853
rect 49400 5819 49416 5853
rect 49516 5819 49532 5853
rect 49658 5819 49674 5853
rect 49774 5819 49790 5853
rect 49916 5819 49932 5853
rect 50032 5819 50048 5853
rect 50174 5819 50190 5853
rect 50290 5819 50306 5853
rect 48690 5751 48724 5813
rect 50574 5947 50603 5981
rect 50637 5947 50695 5981
rect 50729 5947 50787 5981
rect 50821 5947 50850 5981
rect 50466 5751 50500 5812
rect 48690 5750 48786 5751
rect 48690 5717 48736 5750
rect 50430 5718 50500 5751
rect 50404 5717 50500 5718
rect 50640 5905 50706 5913
rect 50640 5871 50656 5905
rect 50690 5871 50706 5905
rect 50640 5837 50706 5871
rect 50640 5803 50656 5837
rect 50690 5803 50706 5837
rect 50640 5769 50706 5803
rect 50640 5735 50656 5769
rect 50690 5735 50706 5769
rect 50640 5717 50706 5735
rect 50740 5905 50782 5947
rect 50774 5871 50782 5905
rect 50740 5837 50782 5871
rect 50774 5803 50782 5837
rect 50740 5769 50782 5803
rect 50774 5735 50782 5769
rect 50740 5719 50782 5735
rect 50640 5658 50686 5717
rect 50681 5610 50686 5658
rect 50720 5680 50786 5683
rect 50720 5669 50737 5680
rect 50720 5635 50736 5669
rect 50783 5640 50786 5680
rect 50770 5635 50786 5640
rect 50640 5597 50686 5610
rect 50640 5585 50706 5597
rect 50640 5551 50656 5585
rect 50690 5551 50706 5585
rect 48690 5516 48760 5550
rect 50430 5516 50500 5550
rect 48690 5454 48724 5516
rect 50466 5454 50500 5516
rect 50640 5517 50706 5551
rect 50640 5483 50656 5517
rect 50690 5483 50706 5517
rect 50640 5471 50706 5483
rect 50740 5585 50786 5601
rect 50774 5551 50786 5585
rect 50740 5517 50786 5551
rect 50774 5483 50786 5517
rect 48884 5414 48900 5448
rect 49000 5414 49016 5448
rect 49142 5414 49158 5448
rect 49258 5414 49274 5448
rect 49400 5414 49416 5448
rect 49516 5414 49532 5448
rect 49658 5414 49674 5448
rect 49774 5414 49790 5448
rect 49916 5414 49932 5448
rect 50032 5414 50048 5448
rect 50174 5414 50190 5448
rect 50290 5414 50306 5448
rect 48804 5364 48838 5380
rect 48804 5172 48838 5188
rect 49062 5364 49096 5380
rect 49062 5172 49096 5188
rect 49320 5364 49354 5380
rect 49320 5172 49354 5188
rect 49578 5364 49612 5380
rect 49578 5172 49612 5188
rect 49836 5364 49870 5380
rect 49836 5172 49870 5188
rect 50094 5364 50128 5380
rect 50094 5172 50128 5188
rect 50352 5364 50386 5380
rect 50352 5172 50386 5188
rect 48884 5104 48900 5138
rect 49000 5104 49016 5138
rect 49142 5104 49158 5138
rect 49258 5104 49274 5138
rect 49400 5104 49416 5138
rect 49516 5104 49532 5138
rect 49658 5104 49674 5138
rect 49774 5104 49790 5138
rect 49916 5104 49932 5138
rect 50032 5104 50048 5138
rect 50174 5104 50190 5138
rect 50290 5104 50306 5138
rect 50740 5437 50786 5483
rect 50574 5403 50603 5437
rect 50637 5403 50695 5437
rect 50729 5403 50787 5437
rect 50821 5403 50850 5437
rect 48690 5036 48724 5098
rect 50466 5036 50500 5098
rect 48690 5002 48758 5036
rect 50432 5002 50500 5036
rect 48690 4450 48736 4483
rect 50430 4450 50500 4483
rect 48690 4449 48786 4450
rect 50404 4449 50500 4450
rect 48690 4387 48724 4449
rect 50466 4388 50500 4449
rect 48884 4347 48900 4381
rect 49000 4347 49016 4381
rect 49142 4347 49158 4381
rect 49258 4347 49274 4381
rect 49400 4347 49416 4381
rect 49516 4347 49532 4381
rect 49658 4347 49674 4381
rect 49774 4347 49790 4381
rect 49916 4347 49932 4381
rect 50032 4347 50048 4381
rect 50174 4347 50190 4381
rect 50290 4347 50306 4381
rect 48804 4288 48838 4304
rect 48804 3896 48838 3912
rect 49062 4288 49096 4304
rect 49062 3896 49096 3912
rect 49320 4288 49354 4304
rect 49320 3896 49354 3912
rect 49578 4288 49612 4304
rect 49578 3896 49612 3912
rect 49836 4288 49870 4304
rect 49836 3896 49870 3912
rect 50094 4288 50128 4304
rect 50094 3896 50128 3912
rect 50352 4288 50386 4304
rect 50352 3896 50386 3912
rect 48884 3819 48900 3853
rect 49000 3819 49016 3853
rect 49142 3819 49158 3853
rect 49258 3819 49274 3853
rect 49400 3819 49416 3853
rect 49516 3819 49532 3853
rect 49658 3819 49674 3853
rect 49774 3819 49790 3853
rect 49916 3819 49932 3853
rect 50032 3819 50048 3853
rect 50174 3819 50190 3853
rect 50290 3819 50306 3853
rect 48690 3751 48724 3813
rect 50574 3947 50603 3981
rect 50637 3947 50695 3981
rect 50729 3947 50787 3981
rect 50821 3947 50850 3981
rect 50466 3751 50500 3812
rect 48690 3750 48786 3751
rect 48690 3717 48736 3750
rect 50430 3718 50500 3751
rect 50404 3717 50500 3718
rect 50640 3905 50706 3913
rect 50640 3871 50656 3905
rect 50690 3871 50706 3905
rect 50640 3837 50706 3871
rect 50640 3803 50656 3837
rect 50690 3803 50706 3837
rect 50640 3769 50706 3803
rect 50640 3735 50656 3769
rect 50690 3735 50706 3769
rect 50640 3717 50706 3735
rect 50740 3905 50782 3947
rect 50774 3871 50782 3905
rect 50740 3837 50782 3871
rect 50774 3803 50782 3837
rect 50740 3769 50782 3803
rect 50774 3735 50782 3769
rect 50740 3719 50782 3735
rect 50640 3658 50686 3717
rect 50681 3610 50686 3658
rect 50720 3680 50786 3683
rect 50720 3669 50737 3680
rect 50720 3635 50736 3669
rect 50783 3640 50786 3680
rect 50770 3635 50786 3640
rect 50640 3597 50686 3610
rect 50640 3585 50706 3597
rect 50640 3551 50656 3585
rect 50690 3551 50706 3585
rect 48690 3516 48760 3550
rect 50430 3516 50500 3550
rect 48690 3454 48724 3516
rect 50466 3454 50500 3516
rect 50640 3517 50706 3551
rect 50640 3483 50656 3517
rect 50690 3483 50706 3517
rect 50640 3471 50706 3483
rect 50740 3585 50786 3601
rect 50774 3551 50786 3585
rect 50740 3517 50786 3551
rect 50774 3483 50786 3517
rect 48884 3414 48900 3448
rect 49000 3414 49016 3448
rect 49142 3414 49158 3448
rect 49258 3414 49274 3448
rect 49400 3414 49416 3448
rect 49516 3414 49532 3448
rect 49658 3414 49674 3448
rect 49774 3414 49790 3448
rect 49916 3414 49932 3448
rect 50032 3414 50048 3448
rect 50174 3414 50190 3448
rect 50290 3414 50306 3448
rect 48804 3364 48838 3380
rect 48804 3172 48838 3188
rect 49062 3364 49096 3380
rect 49062 3172 49096 3188
rect 49320 3364 49354 3380
rect 49320 3172 49354 3188
rect 49578 3364 49612 3380
rect 49578 3172 49612 3188
rect 49836 3364 49870 3380
rect 49836 3172 49870 3188
rect 50094 3364 50128 3380
rect 50094 3172 50128 3188
rect 50352 3364 50386 3380
rect 50352 3172 50386 3188
rect 48884 3104 48900 3138
rect 49000 3104 49016 3138
rect 49142 3104 49158 3138
rect 49258 3104 49274 3138
rect 49400 3104 49416 3138
rect 49516 3104 49532 3138
rect 49658 3104 49674 3138
rect 49774 3104 49790 3138
rect 49916 3104 49932 3138
rect 50032 3104 50048 3138
rect 50174 3104 50190 3138
rect 50290 3104 50306 3138
rect 50740 3437 50786 3483
rect 50574 3403 50603 3437
rect 50637 3403 50695 3437
rect 50729 3403 50787 3437
rect 50821 3403 50850 3437
rect 48690 3036 48724 3098
rect 50466 3036 50500 3098
rect 48690 3002 48758 3036
rect 50432 3002 50500 3036
rect 48690 2360 48736 2393
rect 50430 2360 50500 2393
rect 48690 2359 48786 2360
rect 50404 2359 50500 2360
rect 48690 2297 48724 2359
rect 50466 2298 50500 2359
rect 48884 2257 48900 2291
rect 49000 2257 49016 2291
rect 49142 2257 49158 2291
rect 49258 2257 49274 2291
rect 49400 2257 49416 2291
rect 49516 2257 49532 2291
rect 49658 2257 49674 2291
rect 49774 2257 49790 2291
rect 49916 2257 49932 2291
rect 50032 2257 50048 2291
rect 50174 2257 50190 2291
rect 50290 2257 50306 2291
rect 48804 2198 48838 2214
rect 48804 1806 48838 1822
rect 49062 2198 49096 2214
rect 49062 1806 49096 1822
rect 49320 2198 49354 2214
rect 49320 1806 49354 1822
rect 49578 2198 49612 2214
rect 49578 1806 49612 1822
rect 49836 2198 49870 2214
rect 49836 1806 49870 1822
rect 50094 2198 50128 2214
rect 50094 1806 50128 1822
rect 50352 2198 50386 2214
rect 50352 1806 50386 1822
rect 48884 1729 48900 1763
rect 49000 1729 49016 1763
rect 49142 1729 49158 1763
rect 49258 1729 49274 1763
rect 49400 1729 49416 1763
rect 49516 1729 49532 1763
rect 49658 1729 49674 1763
rect 49774 1729 49790 1763
rect 49916 1729 49932 1763
rect 50032 1729 50048 1763
rect 50174 1729 50190 1763
rect 50290 1729 50306 1763
rect 48690 1661 48724 1723
rect 50574 1857 50603 1891
rect 50637 1857 50695 1891
rect 50729 1857 50787 1891
rect 50821 1857 50850 1891
rect 50466 1661 50500 1722
rect 48690 1660 48786 1661
rect 48690 1627 48736 1660
rect 50430 1628 50500 1661
rect 50404 1627 50500 1628
rect 50640 1815 50706 1823
rect 50640 1781 50656 1815
rect 50690 1781 50706 1815
rect 50640 1747 50706 1781
rect 50640 1713 50656 1747
rect 50690 1713 50706 1747
rect 50640 1679 50706 1713
rect 50640 1645 50656 1679
rect 50690 1645 50706 1679
rect 50640 1627 50706 1645
rect 50740 1815 50782 1857
rect 50774 1781 50782 1815
rect 50740 1747 50782 1781
rect 50774 1713 50782 1747
rect 50740 1679 50782 1713
rect 50774 1645 50782 1679
rect 50740 1629 50782 1645
rect 50640 1568 50686 1627
rect 50681 1520 50686 1568
rect 50720 1590 50786 1593
rect 50720 1579 50737 1590
rect 50720 1545 50736 1579
rect 50783 1550 50786 1590
rect 50770 1545 50786 1550
rect 50640 1507 50686 1520
rect 50640 1495 50706 1507
rect 50640 1461 50656 1495
rect 50690 1461 50706 1495
rect 48690 1426 48760 1460
rect 50430 1426 50500 1460
rect 48690 1364 48724 1426
rect 50466 1364 50500 1426
rect 50640 1427 50706 1461
rect 50640 1393 50656 1427
rect 50690 1393 50706 1427
rect 50640 1381 50706 1393
rect 50740 1495 50786 1511
rect 50774 1461 50786 1495
rect 50740 1427 50786 1461
rect 50774 1393 50786 1427
rect 48884 1324 48900 1358
rect 49000 1324 49016 1358
rect 49142 1324 49158 1358
rect 49258 1324 49274 1358
rect 49400 1324 49416 1358
rect 49516 1324 49532 1358
rect 49658 1324 49674 1358
rect 49774 1324 49790 1358
rect 49916 1324 49932 1358
rect 50032 1324 50048 1358
rect 50174 1324 50190 1358
rect 50290 1324 50306 1358
rect 48804 1274 48838 1290
rect 48804 1082 48838 1098
rect 49062 1274 49096 1290
rect 49062 1082 49096 1098
rect 49320 1274 49354 1290
rect 49320 1082 49354 1098
rect 49578 1274 49612 1290
rect 49578 1082 49612 1098
rect 49836 1274 49870 1290
rect 49836 1082 49870 1098
rect 50094 1274 50128 1290
rect 50094 1082 50128 1098
rect 50352 1274 50386 1290
rect 50352 1082 50386 1098
rect 48884 1014 48900 1048
rect 49000 1014 49016 1048
rect 49142 1014 49158 1048
rect 49258 1014 49274 1048
rect 49400 1014 49416 1048
rect 49516 1014 49532 1048
rect 49658 1014 49674 1048
rect 49774 1014 49790 1048
rect 49916 1014 49932 1048
rect 50032 1014 50048 1048
rect 50174 1014 50190 1048
rect 50290 1014 50306 1048
rect 50740 1347 50786 1393
rect 50574 1313 50603 1347
rect 50637 1313 50695 1347
rect 50729 1313 50787 1347
rect 50821 1313 50850 1347
rect 48690 946 48724 1008
rect 50466 946 50500 1008
rect 48690 912 48758 946
rect 50432 912 50500 946
rect 35772 -682 35872 -520
rect 67532 14810 67566 14826
rect 56282 14318 56364 14342
rect 56282 14284 56306 14318
rect 56340 14284 56364 14318
rect 56282 14260 56364 14284
rect 57300 14318 57382 14342
rect 57300 14284 57324 14318
rect 57358 14284 57382 14318
rect 57300 14260 57382 14284
rect 58318 14318 58400 14342
rect 58318 14284 58342 14318
rect 58376 14284 58400 14318
rect 58318 14260 58400 14284
rect 59336 14318 59418 14342
rect 59336 14284 59360 14318
rect 59394 14284 59418 14318
rect 59336 14260 59418 14284
rect 60354 14318 60436 14342
rect 60354 14284 60378 14318
rect 60412 14284 60436 14318
rect 60354 14260 60436 14284
rect 61372 14318 61454 14342
rect 61372 14284 61396 14318
rect 61430 14284 61454 14318
rect 61372 14260 61454 14284
rect 62390 14318 62472 14342
rect 62390 14284 62414 14318
rect 62448 14284 62472 14318
rect 62390 14260 62472 14284
rect 63408 14318 63490 14342
rect 63408 14284 63432 14318
rect 63466 14284 63490 14318
rect 63408 14260 63490 14284
rect 64426 14318 64508 14342
rect 64426 14284 64450 14318
rect 64484 14284 64508 14318
rect 64426 14260 64508 14284
rect 67532 14218 67566 14234
rect 68550 14810 68584 14826
rect 68550 14218 68584 14234
rect 69568 14810 69602 14826
rect 69568 14218 69602 14234
rect 70586 14810 70620 14826
rect 70586 14218 70620 14234
rect 71604 14810 71638 14826
rect 71604 14218 71638 14234
rect 72622 14810 72656 14826
rect 72622 14218 72656 14234
rect 73640 14810 73674 14826
rect 73640 14218 73674 14234
rect 74658 14810 74692 14826
rect 74658 14218 74692 14234
rect 75676 14810 75710 14826
rect 75676 14218 75710 14234
rect 76694 14810 76728 14826
rect 76694 14218 76728 14234
rect 77712 14810 77746 14826
rect 77712 14218 77746 14234
rect 78730 14810 78764 14826
rect 78730 14218 78764 14234
rect 79748 14810 79782 14826
rect 79748 14218 79782 14234
rect 80766 14810 80800 14826
rect 80766 14218 80800 14234
rect 81784 14810 81818 14826
rect 81784 14218 81818 14234
rect 82802 14810 82836 14826
rect 82802 14218 82836 14234
rect 83820 14810 83854 14826
rect 83820 14218 83854 14234
rect 84838 14810 84872 14826
rect 84838 14218 84872 14234
rect 85856 14810 85890 14826
rect 85856 14218 85890 14234
rect 86874 14810 86908 14826
rect 86874 14218 86908 14234
rect 87892 14810 87926 14826
rect 87892 14218 87926 14234
rect 69050 14184 69110 14186
rect 70064 14184 70124 14192
rect 71068 14184 71128 14198
rect 72094 14184 72154 14186
rect 73118 14184 73178 14192
rect 74138 14184 74198 14186
rect 76164 14184 76224 14192
rect 77188 14184 77248 14186
rect 78198 14184 78258 14186
rect 79218 14184 79278 14192
rect 80248 14184 80308 14186
rect 81252 14184 81312 14192
rect 82268 14184 82328 14192
rect 83298 14184 83358 14186
rect 84312 14184 84372 14186
rect 85328 14184 85388 14186
rect 86354 14184 86414 14186
rect 87376 14184 87436 14186
rect 67764 14150 67780 14184
rect 68336 14150 68352 14184
rect 68782 14150 68798 14184
rect 69354 14150 69370 14184
rect 69800 14150 69816 14184
rect 70372 14150 70388 14184
rect 70818 14150 70834 14184
rect 71390 14150 71406 14184
rect 71836 14150 71852 14184
rect 72408 14150 72424 14184
rect 72854 14150 72870 14184
rect 73426 14150 73442 14184
rect 73872 14150 73888 14184
rect 74444 14150 74460 14184
rect 74890 14150 74906 14184
rect 75462 14150 75478 14184
rect 75908 14150 75924 14184
rect 76480 14150 76496 14184
rect 76926 14150 76942 14184
rect 77498 14150 77514 14184
rect 77944 14150 77960 14184
rect 78516 14150 78532 14184
rect 78962 14150 78978 14184
rect 79534 14150 79550 14184
rect 79980 14150 79996 14184
rect 80552 14150 80568 14184
rect 80998 14150 81014 14184
rect 81570 14150 81586 14184
rect 82016 14150 82032 14184
rect 82588 14150 82604 14184
rect 83034 14150 83050 14184
rect 83606 14150 83622 14184
rect 84052 14150 84068 14184
rect 84624 14150 84640 14184
rect 85070 14150 85086 14184
rect 85642 14150 85658 14184
rect 86088 14150 86104 14184
rect 86660 14150 86676 14184
rect 87106 14150 87122 14184
rect 87678 14150 87694 14184
rect 55998 14066 56014 14100
rect 56570 14066 56586 14100
rect 57016 14066 57032 14100
rect 57588 14066 57604 14100
rect 58034 14066 58050 14100
rect 58606 14066 58622 14100
rect 59052 14066 59068 14100
rect 59624 14066 59640 14100
rect 60070 14066 60086 14100
rect 60642 14066 60658 14100
rect 61088 14066 61104 14100
rect 61660 14066 61676 14100
rect 62106 14066 62122 14100
rect 62678 14066 62694 14100
rect 63124 14066 63140 14100
rect 63696 14066 63712 14100
rect 64142 14066 64158 14100
rect 64714 14066 64730 14100
rect 55766 14016 55800 14032
rect 55766 13424 55800 13440
rect 56784 14016 56818 14032
rect 56784 13424 56818 13440
rect 57802 14016 57836 14032
rect 57802 13424 57836 13440
rect 58820 14016 58854 14032
rect 58820 13424 58854 13440
rect 59838 14016 59872 14032
rect 59838 13424 59872 13440
rect 60856 14016 60890 14032
rect 60856 13424 60890 13440
rect 61874 14016 61908 14032
rect 61874 13424 61908 13440
rect 62892 14016 62926 14032
rect 62892 13424 62926 13440
rect 63910 14016 63944 14032
rect 63910 13424 63944 13440
rect 64928 14016 64962 14032
rect 68016 13926 68098 13950
rect 68016 13892 68040 13926
rect 68074 13892 68098 13926
rect 68016 13868 68098 13892
rect 69034 13926 69116 13950
rect 69034 13892 69058 13926
rect 69092 13892 69116 13926
rect 69034 13868 69116 13892
rect 70052 13926 70134 13950
rect 70052 13892 70076 13926
rect 70110 13892 70134 13926
rect 70052 13868 70134 13892
rect 71070 13926 71152 13950
rect 71070 13892 71094 13926
rect 71128 13892 71152 13926
rect 71070 13868 71152 13892
rect 72088 13926 72170 13950
rect 72088 13892 72112 13926
rect 72146 13892 72170 13926
rect 72088 13868 72170 13892
rect 73106 13926 73188 13950
rect 73106 13892 73130 13926
rect 73164 13892 73188 13926
rect 73106 13868 73188 13892
rect 74124 13926 74206 13950
rect 74124 13892 74148 13926
rect 74182 13892 74206 13926
rect 74124 13868 74206 13892
rect 75142 13926 75224 13950
rect 75142 13892 75166 13926
rect 75200 13892 75224 13926
rect 75142 13868 75224 13892
rect 76160 13926 76242 13950
rect 76160 13892 76184 13926
rect 76218 13892 76242 13926
rect 76160 13868 76242 13892
rect 77178 13926 77260 13950
rect 77178 13892 77202 13926
rect 77236 13892 77260 13926
rect 77178 13868 77260 13892
rect 78196 13926 78278 13950
rect 78196 13892 78220 13926
rect 78254 13892 78278 13926
rect 78196 13868 78278 13892
rect 79214 13926 79296 13950
rect 79214 13892 79238 13926
rect 79272 13892 79296 13926
rect 79214 13868 79296 13892
rect 80232 13926 80314 13950
rect 80232 13892 80256 13926
rect 80290 13892 80314 13926
rect 80232 13868 80314 13892
rect 81250 13926 81332 13950
rect 81250 13892 81274 13926
rect 81308 13892 81332 13926
rect 81250 13868 81332 13892
rect 82268 13926 82350 13950
rect 82268 13892 82292 13926
rect 82326 13892 82350 13926
rect 82268 13868 82350 13892
rect 83286 13926 83368 13950
rect 83286 13892 83310 13926
rect 83344 13892 83368 13926
rect 83286 13868 83368 13892
rect 84304 13926 84386 13950
rect 84304 13892 84328 13926
rect 84362 13892 84386 13926
rect 84304 13868 84386 13892
rect 85322 13926 85404 13950
rect 85322 13892 85346 13926
rect 85380 13892 85404 13926
rect 85322 13868 85404 13892
rect 86340 13926 86422 13950
rect 86340 13892 86364 13926
rect 86398 13892 86422 13926
rect 86340 13868 86422 13892
rect 87358 13926 87440 13950
rect 87358 13892 87382 13926
rect 87416 13892 87440 13926
rect 87358 13868 87440 13892
rect 67764 13626 67780 13660
rect 68336 13626 68352 13660
rect 68782 13626 68798 13660
rect 69354 13626 69370 13660
rect 69800 13626 69816 13660
rect 70372 13626 70388 13660
rect 70818 13626 70834 13660
rect 71390 13626 71406 13660
rect 71836 13626 71852 13660
rect 72408 13626 72424 13660
rect 72854 13626 72870 13660
rect 73426 13626 73442 13660
rect 73872 13626 73888 13660
rect 74444 13626 74460 13660
rect 74890 13626 74906 13660
rect 75462 13626 75478 13660
rect 75908 13626 75924 13660
rect 76480 13626 76496 13660
rect 76926 13626 76942 13660
rect 77498 13626 77514 13660
rect 77944 13626 77960 13660
rect 78516 13626 78532 13660
rect 78962 13626 78978 13660
rect 79534 13626 79550 13660
rect 79980 13626 79996 13660
rect 80552 13626 80568 13660
rect 80998 13626 81014 13660
rect 81570 13626 81586 13660
rect 82016 13626 82032 13660
rect 82588 13626 82604 13660
rect 83034 13626 83050 13660
rect 83606 13626 83622 13660
rect 84052 13626 84068 13660
rect 84624 13626 84640 13660
rect 85070 13626 85086 13660
rect 85642 13626 85658 13660
rect 86088 13626 86104 13660
rect 86660 13626 86676 13660
rect 87106 13626 87122 13660
rect 87678 13626 87694 13660
rect 77188 13620 77248 13626
rect 64928 13424 64962 13440
rect 67532 13576 67566 13592
rect 55744 13336 55826 13360
rect 55998 13356 56014 13390
rect 56570 13356 56586 13390
rect 55744 13302 55768 13336
rect 55802 13302 55826 13336
rect 55744 13278 55826 13302
rect 56762 13336 56844 13360
rect 57016 13356 57032 13390
rect 57588 13356 57604 13390
rect 56762 13302 56786 13336
rect 56820 13302 56844 13336
rect 55998 13248 56014 13282
rect 56570 13248 56586 13282
rect 56762 13278 56844 13302
rect 57780 13336 57862 13360
rect 58034 13356 58050 13390
rect 58606 13356 58622 13390
rect 57780 13302 57804 13336
rect 57838 13302 57862 13336
rect 57016 13248 57032 13282
rect 57588 13248 57604 13282
rect 57780 13278 57862 13302
rect 58798 13336 58880 13360
rect 59052 13356 59068 13390
rect 59624 13356 59640 13390
rect 58798 13302 58822 13336
rect 58856 13302 58880 13336
rect 58034 13248 58050 13282
rect 58606 13248 58622 13282
rect 58798 13278 58880 13302
rect 59816 13336 59898 13360
rect 60070 13356 60086 13390
rect 60642 13356 60658 13390
rect 59816 13302 59840 13336
rect 59874 13302 59898 13336
rect 59052 13248 59068 13282
rect 59624 13248 59640 13282
rect 59816 13278 59898 13302
rect 60834 13336 60916 13360
rect 61088 13356 61104 13390
rect 61660 13356 61676 13390
rect 60834 13302 60858 13336
rect 60892 13302 60916 13336
rect 60070 13248 60086 13282
rect 60642 13248 60658 13282
rect 60834 13278 60916 13302
rect 61852 13336 61934 13360
rect 62106 13356 62122 13390
rect 62678 13356 62694 13390
rect 61852 13302 61876 13336
rect 61910 13302 61934 13336
rect 61088 13248 61104 13282
rect 61660 13248 61676 13282
rect 61852 13278 61934 13302
rect 62870 13336 62952 13360
rect 63124 13356 63140 13390
rect 63696 13356 63712 13390
rect 62870 13302 62894 13336
rect 62928 13302 62952 13336
rect 62106 13248 62122 13282
rect 62678 13248 62694 13282
rect 62870 13278 62952 13302
rect 63888 13336 63970 13360
rect 64142 13356 64158 13390
rect 64714 13356 64730 13390
rect 63888 13302 63912 13336
rect 63946 13302 63970 13336
rect 63124 13248 63140 13282
rect 63696 13248 63712 13282
rect 63888 13278 63970 13302
rect 64906 13336 64988 13360
rect 64906 13302 64930 13336
rect 64964 13302 64988 13336
rect 64142 13248 64158 13282
rect 64714 13248 64730 13282
rect 64906 13278 64988 13302
rect 61358 13246 61418 13248
rect 55766 13198 55800 13214
rect 55766 12606 55800 12622
rect 56784 13198 56818 13214
rect 56784 12606 56818 12622
rect 57802 13198 57836 13214
rect 57802 12606 57836 12622
rect 58820 13198 58854 13214
rect 58820 12606 58854 12622
rect 59838 13198 59872 13214
rect 59838 12606 59872 12622
rect 60856 13198 60890 13214
rect 60856 12606 60890 12622
rect 61874 13198 61908 13214
rect 61874 12606 61908 12622
rect 62892 13198 62926 13214
rect 62892 12606 62926 12622
rect 63910 13198 63944 13214
rect 63910 12606 63944 12622
rect 64928 13198 64962 13214
rect 67532 12984 67566 13000
rect 68550 13576 68584 13592
rect 68550 12984 68584 13000
rect 69568 13576 69602 13592
rect 69568 12984 69602 13000
rect 70586 13576 70620 13592
rect 70586 12984 70620 13000
rect 71604 13576 71638 13592
rect 71604 12984 71638 13000
rect 72622 13576 72656 13592
rect 72622 12984 72656 13000
rect 73640 13576 73674 13592
rect 73640 12984 73674 13000
rect 74658 13576 74692 13592
rect 74658 12984 74692 13000
rect 75676 13576 75710 13592
rect 75676 12984 75710 13000
rect 76694 13576 76728 13592
rect 76694 12984 76728 13000
rect 77712 13576 77746 13592
rect 77712 12984 77746 13000
rect 78730 13576 78764 13592
rect 78730 12984 78764 13000
rect 79748 13576 79782 13592
rect 79748 12984 79782 13000
rect 80766 13576 80800 13592
rect 80766 12984 80800 13000
rect 81784 13576 81818 13592
rect 81784 12984 81818 13000
rect 82802 13576 82836 13592
rect 82802 12984 82836 13000
rect 83820 13576 83854 13592
rect 83820 12984 83854 13000
rect 84838 13576 84872 13592
rect 84838 12984 84872 13000
rect 85856 13576 85890 13592
rect 85856 12984 85890 13000
rect 86874 13576 86908 13592
rect 86874 12984 86908 13000
rect 87892 13576 87926 13592
rect 87892 12984 87926 13000
rect 73116 12950 73176 12956
rect 75152 12950 75212 12956
rect 76172 12950 76232 12956
rect 81244 12950 81304 12956
rect 67764 12916 67780 12950
rect 68336 12916 68352 12950
rect 68782 12916 68798 12950
rect 69354 12916 69370 12950
rect 69800 12916 69816 12950
rect 70372 12916 70388 12950
rect 70818 12916 70834 12950
rect 71390 12916 71406 12950
rect 71836 12916 71852 12950
rect 72408 12916 72424 12950
rect 72854 12916 72870 12950
rect 73426 12916 73442 12950
rect 73872 12916 73888 12950
rect 74444 12916 74460 12950
rect 74890 12916 74906 12950
rect 75462 12916 75478 12950
rect 75908 12916 75924 12950
rect 76480 12916 76496 12950
rect 76926 12916 76942 12950
rect 77498 12916 77514 12950
rect 77944 12916 77960 12950
rect 78516 12916 78532 12950
rect 78962 12916 78978 12950
rect 79534 12916 79550 12950
rect 79980 12916 79996 12950
rect 80552 12916 80568 12950
rect 80998 12916 81014 12950
rect 81570 12916 81586 12950
rect 82016 12916 82032 12950
rect 82588 12916 82604 12950
rect 83034 12916 83050 12950
rect 83606 12916 83622 12950
rect 84052 12916 84068 12950
rect 84624 12916 84640 12950
rect 85070 12916 85086 12950
rect 85642 12916 85658 12950
rect 86088 12916 86104 12950
rect 86660 12916 86676 12950
rect 87106 12916 87122 12950
rect 87678 12916 87694 12950
rect 68004 12690 68086 12714
rect 68004 12656 68028 12690
rect 68062 12656 68086 12690
rect 68004 12632 68086 12656
rect 69022 12690 69104 12714
rect 69022 12656 69046 12690
rect 69080 12656 69104 12690
rect 69022 12632 69104 12656
rect 70040 12690 70122 12714
rect 70040 12656 70064 12690
rect 70098 12656 70122 12690
rect 70040 12632 70122 12656
rect 71058 12690 71140 12714
rect 71058 12656 71082 12690
rect 71116 12656 71140 12690
rect 71058 12632 71140 12656
rect 72076 12690 72158 12714
rect 72076 12656 72100 12690
rect 72134 12656 72158 12690
rect 72076 12632 72158 12656
rect 73094 12690 73176 12714
rect 73094 12656 73118 12690
rect 73152 12656 73176 12690
rect 73094 12632 73176 12656
rect 74112 12690 74194 12714
rect 74112 12656 74136 12690
rect 74170 12656 74194 12690
rect 74112 12632 74194 12656
rect 75130 12690 75212 12714
rect 75130 12656 75154 12690
rect 75188 12656 75212 12690
rect 75130 12632 75212 12656
rect 76148 12690 76230 12714
rect 76148 12656 76172 12690
rect 76206 12656 76230 12690
rect 76148 12632 76230 12656
rect 77166 12690 77248 12714
rect 77166 12656 77190 12690
rect 77224 12656 77248 12690
rect 77166 12632 77248 12656
rect 78184 12690 78266 12714
rect 78184 12656 78208 12690
rect 78242 12656 78266 12690
rect 78184 12632 78266 12656
rect 79202 12690 79284 12714
rect 79202 12656 79226 12690
rect 79260 12656 79284 12690
rect 79202 12632 79284 12656
rect 80220 12690 80302 12714
rect 80220 12656 80244 12690
rect 80278 12656 80302 12690
rect 80220 12632 80302 12656
rect 81238 12690 81320 12714
rect 81238 12656 81262 12690
rect 81296 12656 81320 12690
rect 81238 12632 81320 12656
rect 82256 12690 82338 12714
rect 82256 12656 82280 12690
rect 82314 12656 82338 12690
rect 82256 12632 82338 12656
rect 83274 12690 83356 12714
rect 83274 12656 83298 12690
rect 83332 12656 83356 12690
rect 83274 12632 83356 12656
rect 84292 12690 84374 12714
rect 84292 12656 84316 12690
rect 84350 12656 84374 12690
rect 84292 12632 84374 12656
rect 85310 12690 85392 12714
rect 85310 12656 85334 12690
rect 85368 12656 85392 12690
rect 85310 12632 85392 12656
rect 86328 12690 86410 12714
rect 86328 12656 86352 12690
rect 86386 12656 86410 12690
rect 86328 12632 86410 12656
rect 87346 12690 87428 12714
rect 87346 12656 87370 12690
rect 87404 12656 87428 12690
rect 87346 12632 87428 12656
rect 64928 12606 64962 12622
rect 57290 12572 57350 12574
rect 58304 12572 58364 12574
rect 62378 12572 62438 12574
rect 63394 12572 63454 12574
rect 55744 12518 55826 12542
rect 55998 12538 56014 12572
rect 56570 12538 56586 12572
rect 55744 12484 55768 12518
rect 55802 12484 55826 12518
rect 55744 12460 55826 12484
rect 56762 12518 56844 12542
rect 57016 12538 57032 12572
rect 57588 12538 57604 12572
rect 56762 12484 56786 12518
rect 56820 12484 56844 12518
rect 55998 12430 56014 12464
rect 56570 12430 56586 12464
rect 56762 12460 56844 12484
rect 57780 12518 57862 12542
rect 58034 12538 58050 12572
rect 58606 12538 58622 12572
rect 57780 12484 57804 12518
rect 57838 12484 57862 12518
rect 57016 12430 57032 12464
rect 57588 12430 57604 12464
rect 57780 12460 57862 12484
rect 58798 12518 58880 12542
rect 59052 12538 59068 12572
rect 59624 12538 59640 12572
rect 58798 12484 58822 12518
rect 58856 12484 58880 12518
rect 58034 12430 58050 12464
rect 58606 12430 58622 12464
rect 58798 12460 58880 12484
rect 59816 12518 59898 12542
rect 60070 12538 60086 12572
rect 60642 12538 60658 12572
rect 59816 12484 59840 12518
rect 59874 12484 59898 12518
rect 59052 12430 59068 12464
rect 59624 12430 59640 12464
rect 59816 12460 59898 12484
rect 60834 12518 60916 12542
rect 61088 12538 61104 12572
rect 61660 12538 61676 12572
rect 60834 12484 60858 12518
rect 60892 12484 60916 12518
rect 60070 12430 60086 12464
rect 60642 12430 60658 12464
rect 60834 12460 60916 12484
rect 61852 12518 61934 12542
rect 62106 12538 62122 12572
rect 62678 12538 62694 12572
rect 61852 12484 61876 12518
rect 61910 12484 61934 12518
rect 61088 12430 61104 12464
rect 61660 12430 61676 12464
rect 61852 12460 61934 12484
rect 62870 12518 62952 12542
rect 63124 12538 63140 12572
rect 63696 12538 63712 12572
rect 62870 12484 62894 12518
rect 62928 12484 62952 12518
rect 62106 12430 62122 12464
rect 62678 12430 62694 12464
rect 62870 12460 62952 12484
rect 63888 12518 63970 12542
rect 64142 12538 64158 12572
rect 64714 12538 64730 12572
rect 63888 12484 63912 12518
rect 63946 12484 63970 12518
rect 63124 12430 63140 12464
rect 63696 12430 63712 12464
rect 63888 12460 63970 12484
rect 64906 12518 64988 12542
rect 64906 12484 64930 12518
rect 64964 12484 64988 12518
rect 64142 12430 64158 12464
rect 64714 12430 64730 12464
rect 64906 12460 64988 12484
rect 55766 12380 55800 12396
rect 55766 11788 55800 11804
rect 56784 12380 56818 12396
rect 56784 11788 56818 11804
rect 57802 12380 57836 12396
rect 57802 11788 57836 11804
rect 58820 12380 58854 12396
rect 58820 11788 58854 11804
rect 59838 12380 59872 12396
rect 59838 11788 59872 11804
rect 60856 12380 60890 12396
rect 60856 11788 60890 11804
rect 61874 12380 61908 12396
rect 61874 11788 61908 11804
rect 62892 12380 62926 12396
rect 62892 11788 62926 11804
rect 63910 12380 63944 12396
rect 63910 11788 63944 11804
rect 64928 12380 64962 12396
rect 67764 12394 67780 12428
rect 68336 12394 68352 12428
rect 68782 12394 68798 12428
rect 69354 12394 69370 12428
rect 69800 12394 69816 12428
rect 70372 12394 70388 12428
rect 70818 12394 70834 12428
rect 71390 12394 71406 12428
rect 71836 12394 71852 12428
rect 72408 12394 72424 12428
rect 72854 12394 72870 12428
rect 73426 12394 73442 12428
rect 73872 12394 73888 12428
rect 74444 12394 74460 12428
rect 74890 12394 74906 12428
rect 75462 12394 75478 12428
rect 75908 12394 75924 12428
rect 76480 12394 76496 12428
rect 76926 12394 76942 12428
rect 77498 12394 77514 12428
rect 77944 12394 77960 12428
rect 78516 12394 78532 12428
rect 78962 12394 78978 12428
rect 79534 12394 79550 12428
rect 79980 12394 79996 12428
rect 80552 12394 80568 12428
rect 80998 12394 81014 12428
rect 81570 12394 81586 12428
rect 82016 12394 82032 12428
rect 82588 12394 82604 12428
rect 83034 12394 83050 12428
rect 83606 12394 83622 12428
rect 84052 12394 84068 12428
rect 84624 12394 84640 12428
rect 85070 12394 85086 12428
rect 85642 12394 85658 12428
rect 86088 12394 86104 12428
rect 86660 12394 86676 12428
rect 87106 12394 87122 12428
rect 87678 12394 87694 12428
rect 69050 12390 69110 12394
rect 70066 12390 70126 12394
rect 74142 12386 74202 12394
rect 78208 12390 78268 12394
rect 80242 12390 80302 12394
rect 86354 12390 86414 12394
rect 64928 11788 64962 11804
rect 67532 12344 67566 12360
rect 57294 11754 57354 11756
rect 58308 11754 58368 11756
rect 62382 11754 62442 11756
rect 63398 11754 63458 11756
rect 55744 11700 55826 11724
rect 55998 11720 56014 11754
rect 56570 11720 56586 11754
rect 55744 11666 55768 11700
rect 55802 11666 55826 11700
rect 55744 11642 55826 11666
rect 56762 11700 56844 11724
rect 57016 11720 57032 11754
rect 57588 11720 57604 11754
rect 56762 11666 56786 11700
rect 56820 11666 56844 11700
rect 55998 11612 56014 11646
rect 56570 11612 56586 11646
rect 56762 11642 56844 11666
rect 57780 11700 57862 11724
rect 58034 11720 58050 11754
rect 58606 11720 58622 11754
rect 57780 11666 57804 11700
rect 57838 11666 57862 11700
rect 57016 11612 57032 11646
rect 57588 11612 57604 11646
rect 57780 11642 57862 11666
rect 58798 11700 58880 11724
rect 59052 11720 59068 11754
rect 59624 11720 59640 11754
rect 58798 11666 58822 11700
rect 58856 11666 58880 11700
rect 58034 11612 58050 11646
rect 58606 11612 58622 11646
rect 58798 11642 58880 11666
rect 59816 11700 59898 11724
rect 60070 11720 60086 11754
rect 60642 11720 60658 11754
rect 59816 11666 59840 11700
rect 59874 11666 59898 11700
rect 59052 11612 59068 11646
rect 59624 11612 59640 11646
rect 59816 11642 59898 11666
rect 60834 11700 60916 11724
rect 61088 11720 61104 11754
rect 61660 11720 61676 11754
rect 60834 11666 60858 11700
rect 60892 11666 60916 11700
rect 60070 11612 60086 11646
rect 60642 11612 60658 11646
rect 60834 11642 60916 11666
rect 61852 11700 61934 11724
rect 62106 11720 62122 11754
rect 62678 11720 62694 11754
rect 61852 11666 61876 11700
rect 61910 11666 61934 11700
rect 61088 11612 61104 11646
rect 61660 11612 61676 11646
rect 61852 11642 61934 11666
rect 62870 11700 62952 11724
rect 63124 11720 63140 11754
rect 63696 11720 63712 11754
rect 62870 11666 62894 11700
rect 62928 11666 62952 11700
rect 62106 11612 62122 11646
rect 62678 11612 62694 11646
rect 62870 11642 62952 11666
rect 63888 11700 63970 11724
rect 64142 11720 64158 11754
rect 64714 11720 64730 11754
rect 67532 11752 67566 11768
rect 68550 12344 68584 12360
rect 68550 11752 68584 11768
rect 69568 12344 69602 12360
rect 69568 11752 69602 11768
rect 70586 12344 70620 12360
rect 70586 11752 70620 11768
rect 71604 12344 71638 12360
rect 71604 11752 71638 11768
rect 72622 12344 72656 12360
rect 72622 11752 72656 11768
rect 73640 12344 73674 12360
rect 73640 11752 73674 11768
rect 74658 12344 74692 12360
rect 74658 11752 74692 11768
rect 75676 12344 75710 12360
rect 75676 11752 75710 11768
rect 76694 12344 76728 12360
rect 76694 11752 76728 11768
rect 77712 12344 77746 12360
rect 77712 11752 77746 11768
rect 78730 12344 78764 12360
rect 78730 11752 78764 11768
rect 79748 12344 79782 12360
rect 79748 11752 79782 11768
rect 80766 12344 80800 12360
rect 80766 11752 80800 11768
rect 81784 12344 81818 12360
rect 81784 11752 81818 11768
rect 82802 12344 82836 12360
rect 82802 11752 82836 11768
rect 83820 12344 83854 12360
rect 83820 11752 83854 11768
rect 84838 12344 84872 12360
rect 84838 11752 84872 11768
rect 85856 12344 85890 12360
rect 85856 11752 85890 11768
rect 86874 12344 86908 12360
rect 86874 11752 86908 11768
rect 87892 12344 87926 12360
rect 87892 11752 87926 11768
rect 63888 11666 63912 11700
rect 63946 11666 63970 11700
rect 63124 11612 63140 11646
rect 63696 11612 63712 11646
rect 63888 11642 63970 11666
rect 64906 11700 64988 11724
rect 71076 11718 71136 11720
rect 64906 11666 64930 11700
rect 64964 11666 64988 11700
rect 67764 11684 67780 11718
rect 68336 11684 68352 11718
rect 68782 11684 68798 11718
rect 69354 11684 69370 11718
rect 69800 11684 69816 11718
rect 70372 11684 70388 11718
rect 70818 11684 70834 11718
rect 71390 11684 71406 11718
rect 71836 11684 71852 11718
rect 72408 11684 72424 11718
rect 72854 11684 72870 11718
rect 73426 11684 73442 11718
rect 73872 11684 73888 11718
rect 74444 11684 74460 11718
rect 74890 11684 74906 11718
rect 75462 11684 75478 11718
rect 75908 11684 75924 11718
rect 76480 11684 76496 11718
rect 76926 11684 76942 11718
rect 77498 11684 77514 11718
rect 77944 11684 77960 11718
rect 78516 11684 78532 11718
rect 78962 11684 78978 11718
rect 79534 11684 79550 11718
rect 79980 11684 79996 11718
rect 80552 11684 80568 11718
rect 80998 11684 81014 11718
rect 81570 11684 81586 11718
rect 82016 11684 82032 11718
rect 82588 11684 82604 11718
rect 83034 11684 83050 11718
rect 83606 11684 83622 11718
rect 84052 11684 84068 11718
rect 84624 11684 84640 11718
rect 85070 11684 85086 11718
rect 85642 11684 85658 11718
rect 86088 11684 86104 11718
rect 86660 11684 86676 11718
rect 87106 11684 87122 11718
rect 87678 11684 87694 11718
rect 73110 11680 73170 11684
rect 82268 11670 82328 11684
rect 83302 11670 83362 11684
rect 64142 11612 64158 11646
rect 64714 11612 64730 11646
rect 64906 11642 64988 11666
rect 55766 11562 55800 11578
rect 55766 10970 55800 10986
rect 56784 11562 56818 11578
rect 56784 10970 56818 10986
rect 57802 11562 57836 11578
rect 57802 10970 57836 10986
rect 58820 11562 58854 11578
rect 58820 10970 58854 10986
rect 59838 11562 59872 11578
rect 59838 10970 59872 10986
rect 60856 11562 60890 11578
rect 60856 10970 60890 10986
rect 61874 11562 61908 11578
rect 61874 10970 61908 10986
rect 62892 11562 62926 11578
rect 62892 10970 62926 10986
rect 63910 11562 63944 11578
rect 63910 10970 63944 10986
rect 64928 11562 64962 11578
rect 68016 11456 68098 11480
rect 68016 11422 68040 11456
rect 68074 11422 68098 11456
rect 68016 11398 68098 11422
rect 69034 11456 69116 11480
rect 69034 11422 69058 11456
rect 69092 11422 69116 11456
rect 69034 11398 69116 11422
rect 70052 11456 70134 11480
rect 70052 11422 70076 11456
rect 70110 11422 70134 11456
rect 70052 11398 70134 11422
rect 71070 11456 71152 11480
rect 71070 11422 71094 11456
rect 71128 11422 71152 11456
rect 71070 11398 71152 11422
rect 72088 11456 72170 11480
rect 72088 11422 72112 11456
rect 72146 11422 72170 11456
rect 72088 11398 72170 11422
rect 73106 11456 73188 11480
rect 73106 11422 73130 11456
rect 73164 11422 73188 11456
rect 73106 11398 73188 11422
rect 74124 11456 74206 11480
rect 74124 11422 74148 11456
rect 74182 11422 74206 11456
rect 74124 11398 74206 11422
rect 75142 11456 75224 11480
rect 75142 11422 75166 11456
rect 75200 11422 75224 11456
rect 75142 11398 75224 11422
rect 76160 11456 76242 11480
rect 76160 11422 76184 11456
rect 76218 11422 76242 11456
rect 76160 11398 76242 11422
rect 77178 11456 77260 11480
rect 77178 11422 77202 11456
rect 77236 11422 77260 11456
rect 77178 11398 77260 11422
rect 78196 11456 78278 11480
rect 78196 11422 78220 11456
rect 78254 11422 78278 11456
rect 78196 11398 78278 11422
rect 79214 11456 79296 11480
rect 79214 11422 79238 11456
rect 79272 11422 79296 11456
rect 79214 11398 79296 11422
rect 80232 11456 80314 11480
rect 80232 11422 80256 11456
rect 80290 11422 80314 11456
rect 80232 11398 80314 11422
rect 81250 11456 81332 11480
rect 81250 11422 81274 11456
rect 81308 11422 81332 11456
rect 81250 11398 81332 11422
rect 82268 11456 82350 11480
rect 82268 11422 82292 11456
rect 82326 11422 82350 11456
rect 82268 11398 82350 11422
rect 83286 11456 83368 11480
rect 83286 11422 83310 11456
rect 83344 11422 83368 11456
rect 83286 11398 83368 11422
rect 84304 11456 84386 11480
rect 84304 11422 84328 11456
rect 84362 11422 84386 11456
rect 84304 11398 84386 11422
rect 85322 11456 85404 11480
rect 85322 11422 85346 11456
rect 85380 11422 85404 11456
rect 85322 11398 85404 11422
rect 86340 11456 86422 11480
rect 86340 11422 86364 11456
rect 86398 11422 86422 11456
rect 86340 11398 86422 11422
rect 87358 11456 87440 11480
rect 87358 11422 87382 11456
rect 87416 11422 87440 11456
rect 87358 11398 87440 11422
rect 67762 11160 67778 11194
rect 68334 11160 68350 11194
rect 68780 11160 68796 11194
rect 69352 11160 69368 11194
rect 69798 11160 69814 11194
rect 70370 11160 70386 11194
rect 70816 11160 70832 11194
rect 71388 11160 71404 11194
rect 71834 11160 71850 11194
rect 72406 11160 72422 11194
rect 72852 11160 72868 11194
rect 73424 11160 73440 11194
rect 73870 11160 73886 11194
rect 74442 11160 74458 11194
rect 74888 11160 74904 11194
rect 75460 11160 75476 11194
rect 75906 11160 75922 11194
rect 76478 11160 76494 11194
rect 76924 11160 76940 11194
rect 77496 11160 77512 11194
rect 77942 11160 77958 11194
rect 78514 11160 78530 11194
rect 78960 11160 78976 11194
rect 79532 11160 79548 11194
rect 79978 11160 79994 11194
rect 80550 11160 80566 11194
rect 80996 11160 81012 11194
rect 81568 11160 81584 11194
rect 82014 11160 82030 11194
rect 82586 11160 82602 11194
rect 83032 11160 83048 11194
rect 83604 11160 83620 11194
rect 84050 11160 84066 11194
rect 84622 11160 84638 11194
rect 85068 11160 85084 11194
rect 85640 11160 85656 11194
rect 86086 11160 86102 11194
rect 86658 11160 86674 11194
rect 87104 11160 87120 11194
rect 87676 11160 87692 11194
rect 70072 11156 70132 11160
rect 64928 10970 64962 10986
rect 67530 11110 67564 11126
rect 55744 10882 55826 10906
rect 55998 10902 56014 10936
rect 56570 10902 56586 10936
rect 55744 10848 55768 10882
rect 55802 10848 55826 10882
rect 55744 10824 55826 10848
rect 56762 10882 56844 10906
rect 57016 10902 57032 10936
rect 57588 10902 57604 10936
rect 56762 10848 56786 10882
rect 56820 10848 56844 10882
rect 55998 10794 56014 10828
rect 56570 10794 56586 10828
rect 56762 10824 56844 10848
rect 57780 10882 57862 10906
rect 58034 10902 58050 10936
rect 58606 10902 58622 10936
rect 57780 10848 57804 10882
rect 57838 10848 57862 10882
rect 57016 10794 57032 10828
rect 57588 10794 57604 10828
rect 57780 10824 57862 10848
rect 58798 10882 58880 10906
rect 59052 10902 59068 10936
rect 59624 10902 59640 10936
rect 58798 10848 58822 10882
rect 58856 10848 58880 10882
rect 58034 10794 58050 10828
rect 58606 10794 58622 10828
rect 58798 10824 58880 10848
rect 59816 10882 59898 10906
rect 60070 10902 60086 10936
rect 60642 10902 60658 10936
rect 59816 10848 59840 10882
rect 59874 10848 59898 10882
rect 59052 10794 59068 10828
rect 59624 10794 59640 10828
rect 59816 10824 59898 10848
rect 60834 10882 60916 10906
rect 61088 10902 61104 10936
rect 61660 10902 61676 10936
rect 60834 10848 60858 10882
rect 60892 10848 60916 10882
rect 60070 10794 60086 10828
rect 60642 10794 60658 10828
rect 60834 10824 60916 10848
rect 61852 10882 61934 10906
rect 62106 10902 62122 10936
rect 62678 10902 62694 10936
rect 61852 10848 61876 10882
rect 61910 10848 61934 10882
rect 61088 10794 61104 10828
rect 61660 10794 61676 10828
rect 61852 10824 61934 10848
rect 62870 10882 62952 10906
rect 63124 10902 63140 10936
rect 63696 10902 63712 10936
rect 62870 10848 62894 10882
rect 62928 10848 62952 10882
rect 62106 10794 62122 10828
rect 62678 10794 62694 10828
rect 62870 10824 62952 10848
rect 63888 10882 63970 10906
rect 64142 10902 64158 10936
rect 64714 10902 64730 10936
rect 63888 10848 63912 10882
rect 63946 10848 63970 10882
rect 63124 10794 63140 10828
rect 63696 10794 63712 10828
rect 63888 10824 63970 10848
rect 64906 10882 64988 10906
rect 64906 10848 64930 10882
rect 64964 10848 64988 10882
rect 64142 10794 64158 10828
rect 64714 10794 64730 10828
rect 64906 10824 64988 10848
rect 61354 10792 61414 10794
rect 55766 10744 55800 10760
rect 55766 10152 55800 10168
rect 56784 10744 56818 10760
rect 56784 10152 56818 10168
rect 57802 10744 57836 10760
rect 57802 10152 57836 10168
rect 58820 10744 58854 10760
rect 58820 10152 58854 10168
rect 59838 10744 59872 10760
rect 59838 10152 59872 10168
rect 60856 10744 60890 10760
rect 60856 10152 60890 10168
rect 61874 10744 61908 10760
rect 61874 10152 61908 10168
rect 62892 10744 62926 10760
rect 62892 10152 62926 10168
rect 63910 10744 63944 10760
rect 63910 10152 63944 10168
rect 64928 10744 64962 10760
rect 67530 10518 67564 10534
rect 68548 11110 68582 11126
rect 68548 10518 68582 10534
rect 69566 11110 69600 11126
rect 69566 10518 69600 10534
rect 70584 11110 70618 11126
rect 70584 10518 70618 10534
rect 71602 11110 71636 11126
rect 71602 10518 71636 10534
rect 72620 11110 72654 11126
rect 72620 10518 72654 10534
rect 73638 11110 73672 11126
rect 73638 10518 73672 10534
rect 74656 11110 74690 11126
rect 74656 10518 74690 10534
rect 75674 11110 75708 11126
rect 75674 10518 75708 10534
rect 76692 11110 76726 11126
rect 76692 10518 76726 10534
rect 77710 11110 77744 11126
rect 77710 10518 77744 10534
rect 78728 11110 78762 11126
rect 78728 10518 78762 10534
rect 79746 11110 79780 11126
rect 79746 10518 79780 10534
rect 80764 11110 80798 11126
rect 80764 10518 80798 10534
rect 81782 11110 81816 11126
rect 81782 10518 81816 10534
rect 82800 11110 82834 11126
rect 82800 10518 82834 10534
rect 83818 11110 83852 11126
rect 83818 10518 83852 10534
rect 84836 11110 84870 11126
rect 84836 10518 84870 10534
rect 85854 11110 85888 11126
rect 85854 10518 85888 10534
rect 86872 11110 86906 11126
rect 86872 10518 86906 10534
rect 87890 11110 87924 11126
rect 87890 10518 87924 10534
rect 75140 10484 75200 10488
rect 76168 10484 76228 10486
rect 78212 10484 78272 10488
rect 67762 10450 67778 10484
rect 68334 10450 68350 10484
rect 68780 10450 68796 10484
rect 69352 10450 69368 10484
rect 69798 10450 69814 10484
rect 70370 10450 70386 10484
rect 70816 10450 70832 10484
rect 71388 10450 71404 10484
rect 71834 10450 71850 10484
rect 72406 10450 72422 10484
rect 72852 10450 72868 10484
rect 73424 10450 73440 10484
rect 73870 10450 73886 10484
rect 74442 10450 74458 10484
rect 74888 10450 74904 10484
rect 75460 10450 75476 10484
rect 75906 10450 75922 10484
rect 76478 10450 76494 10484
rect 76924 10450 76940 10484
rect 77496 10450 77512 10484
rect 77942 10450 77958 10484
rect 78514 10450 78530 10484
rect 78960 10450 78976 10484
rect 79532 10450 79548 10484
rect 79978 10450 79994 10484
rect 80550 10450 80566 10484
rect 80996 10450 81012 10484
rect 81568 10450 81584 10484
rect 82014 10450 82030 10484
rect 82586 10450 82602 10484
rect 83032 10450 83048 10484
rect 83604 10450 83620 10484
rect 84050 10450 84066 10484
rect 84622 10450 84638 10484
rect 85068 10450 85084 10484
rect 85640 10450 85656 10484
rect 86086 10450 86102 10484
rect 86658 10450 86674 10484
rect 87104 10450 87120 10484
rect 87676 10450 87692 10484
rect 68016 10236 68098 10260
rect 68016 10202 68040 10236
rect 68074 10202 68098 10236
rect 68016 10178 68098 10202
rect 69034 10236 69116 10260
rect 69034 10202 69058 10236
rect 69092 10202 69116 10236
rect 69034 10178 69116 10202
rect 70052 10236 70134 10260
rect 70052 10202 70076 10236
rect 70110 10202 70134 10236
rect 70052 10178 70134 10202
rect 71070 10236 71152 10260
rect 71070 10202 71094 10236
rect 71128 10202 71152 10236
rect 71070 10178 71152 10202
rect 72088 10236 72170 10260
rect 72088 10202 72112 10236
rect 72146 10202 72170 10236
rect 72088 10178 72170 10202
rect 73106 10236 73188 10260
rect 73106 10202 73130 10236
rect 73164 10202 73188 10236
rect 73106 10178 73188 10202
rect 74124 10236 74206 10260
rect 74124 10202 74148 10236
rect 74182 10202 74206 10236
rect 74124 10178 74206 10202
rect 75142 10236 75224 10260
rect 75142 10202 75166 10236
rect 75200 10202 75224 10236
rect 75142 10178 75224 10202
rect 76160 10236 76242 10260
rect 76160 10202 76184 10236
rect 76218 10202 76242 10236
rect 76160 10178 76242 10202
rect 77178 10236 77260 10260
rect 77178 10202 77202 10236
rect 77236 10202 77260 10236
rect 77178 10178 77260 10202
rect 78196 10236 78278 10260
rect 78196 10202 78220 10236
rect 78254 10202 78278 10236
rect 78196 10178 78278 10202
rect 79214 10236 79296 10260
rect 79214 10202 79238 10236
rect 79272 10202 79296 10236
rect 79214 10178 79296 10202
rect 80232 10236 80314 10260
rect 80232 10202 80256 10236
rect 80290 10202 80314 10236
rect 80232 10178 80314 10202
rect 81250 10236 81332 10260
rect 81250 10202 81274 10236
rect 81308 10202 81332 10236
rect 81250 10178 81332 10202
rect 82268 10236 82350 10260
rect 82268 10202 82292 10236
rect 82326 10202 82350 10236
rect 82268 10178 82350 10202
rect 83286 10236 83368 10260
rect 83286 10202 83310 10236
rect 83344 10202 83368 10236
rect 83286 10178 83368 10202
rect 84304 10236 84386 10260
rect 84304 10202 84328 10236
rect 84362 10202 84386 10236
rect 84304 10178 84386 10202
rect 85322 10236 85404 10260
rect 85322 10202 85346 10236
rect 85380 10202 85404 10236
rect 85322 10178 85404 10202
rect 86340 10236 86422 10260
rect 86340 10202 86364 10236
rect 86398 10202 86422 10236
rect 86340 10178 86422 10202
rect 87358 10236 87440 10260
rect 87358 10202 87382 10236
rect 87416 10202 87440 10236
rect 87358 10178 87440 10202
rect 64928 10152 64962 10168
rect 57280 10118 57340 10120
rect 58294 10118 58354 10120
rect 62368 10118 62428 10120
rect 63384 10118 63444 10120
rect 55744 10064 55826 10088
rect 55998 10084 56014 10118
rect 56570 10084 56586 10118
rect 55744 10030 55768 10064
rect 55802 10030 55826 10064
rect 55744 10006 55826 10030
rect 56762 10064 56844 10088
rect 57016 10084 57032 10118
rect 57588 10084 57604 10118
rect 56762 10030 56786 10064
rect 56820 10030 56844 10064
rect 55998 9976 56014 10010
rect 56570 9976 56586 10010
rect 56762 10006 56844 10030
rect 57780 10064 57862 10088
rect 58034 10084 58050 10118
rect 58606 10084 58622 10118
rect 57780 10030 57804 10064
rect 57838 10030 57862 10064
rect 57016 9976 57032 10010
rect 57588 9976 57604 10010
rect 57780 10006 57862 10030
rect 58798 10064 58880 10088
rect 59052 10084 59068 10118
rect 59624 10084 59640 10118
rect 58798 10030 58822 10064
rect 58856 10030 58880 10064
rect 58034 9976 58050 10010
rect 58606 9976 58622 10010
rect 58798 10006 58880 10030
rect 59816 10064 59898 10088
rect 60070 10084 60086 10118
rect 60642 10084 60658 10118
rect 59816 10030 59840 10064
rect 59874 10030 59898 10064
rect 59052 9976 59068 10010
rect 59624 9976 59640 10010
rect 59816 10006 59898 10030
rect 60834 10064 60916 10088
rect 61088 10084 61104 10118
rect 61660 10084 61676 10118
rect 60834 10030 60858 10064
rect 60892 10030 60916 10064
rect 60070 9976 60086 10010
rect 60642 9976 60658 10010
rect 60834 10006 60916 10030
rect 61852 10064 61934 10088
rect 62106 10084 62122 10118
rect 62678 10084 62694 10118
rect 61852 10030 61876 10064
rect 61910 10030 61934 10064
rect 61088 9976 61104 10010
rect 61660 9976 61676 10010
rect 61852 10006 61934 10030
rect 62870 10064 62952 10088
rect 63124 10084 63140 10118
rect 63696 10084 63712 10118
rect 62870 10030 62894 10064
rect 62928 10030 62952 10064
rect 62106 9976 62122 10010
rect 62678 9976 62694 10010
rect 62870 10006 62952 10030
rect 63888 10064 63970 10088
rect 64142 10084 64158 10118
rect 64714 10084 64730 10118
rect 63888 10030 63912 10064
rect 63946 10030 63970 10064
rect 63124 9976 63140 10010
rect 63696 9976 63712 10010
rect 63888 10006 63970 10030
rect 64906 10064 64988 10088
rect 64906 10030 64930 10064
rect 64964 10030 64988 10064
rect 64142 9976 64158 10010
rect 64714 9976 64730 10010
rect 64906 10006 64988 10030
rect 55766 9926 55800 9942
rect 55766 9334 55800 9350
rect 56784 9926 56818 9942
rect 56784 9334 56818 9350
rect 57802 9926 57836 9942
rect 57802 9334 57836 9350
rect 58820 9926 58854 9942
rect 58820 9334 58854 9350
rect 59838 9926 59872 9942
rect 59838 9334 59872 9350
rect 60856 9926 60890 9942
rect 60856 9334 60890 9350
rect 61874 9926 61908 9942
rect 61874 9334 61908 9350
rect 62892 9926 62926 9942
rect 62892 9334 62926 9350
rect 63910 9926 63944 9942
rect 63910 9334 63944 9350
rect 64928 9926 64962 9942
rect 67762 9926 67778 9960
rect 68334 9926 68350 9960
rect 68780 9926 68796 9960
rect 69352 9926 69368 9960
rect 69798 9926 69814 9960
rect 70370 9926 70386 9960
rect 70816 9926 70832 9960
rect 71388 9926 71404 9960
rect 71834 9926 71850 9960
rect 72406 9926 72422 9960
rect 72852 9926 72868 9960
rect 73424 9926 73440 9960
rect 73870 9926 73886 9960
rect 74442 9926 74458 9960
rect 74888 9926 74904 9960
rect 75460 9926 75476 9960
rect 75906 9926 75922 9960
rect 76478 9926 76494 9960
rect 76924 9926 76940 9960
rect 77496 9926 77512 9960
rect 77942 9926 77958 9960
rect 78514 9926 78530 9960
rect 78960 9926 78976 9960
rect 79532 9926 79548 9960
rect 79978 9926 79994 9960
rect 80550 9926 80566 9960
rect 80996 9926 81012 9960
rect 81568 9926 81584 9960
rect 82014 9926 82030 9960
rect 82586 9926 82602 9960
rect 83032 9926 83048 9960
rect 83604 9926 83620 9960
rect 84050 9926 84066 9960
rect 84622 9926 84638 9960
rect 85068 9926 85084 9960
rect 85640 9926 85656 9960
rect 86086 9926 86102 9960
rect 86658 9926 86674 9960
rect 87104 9926 87120 9960
rect 87676 9926 87692 9960
rect 64928 9334 64962 9350
rect 67530 9876 67564 9892
rect 57284 9300 57344 9302
rect 58298 9300 58358 9302
rect 62372 9300 62432 9302
rect 63388 9300 63448 9302
rect 55744 9246 55826 9270
rect 55998 9266 56014 9300
rect 56570 9266 56586 9300
rect 55744 9212 55768 9246
rect 55802 9212 55826 9246
rect 55744 9188 55826 9212
rect 56762 9246 56844 9270
rect 57016 9266 57032 9300
rect 57588 9266 57604 9300
rect 56762 9212 56786 9246
rect 56820 9212 56844 9246
rect 55998 9158 56014 9192
rect 56570 9158 56586 9192
rect 56762 9188 56844 9212
rect 57780 9246 57862 9270
rect 58034 9266 58050 9300
rect 58606 9266 58622 9300
rect 57780 9212 57804 9246
rect 57838 9212 57862 9246
rect 57016 9158 57032 9192
rect 57588 9158 57604 9192
rect 57780 9188 57862 9212
rect 58798 9246 58880 9270
rect 59052 9266 59068 9300
rect 59624 9266 59640 9300
rect 58798 9212 58822 9246
rect 58856 9212 58880 9246
rect 58034 9158 58050 9192
rect 58606 9158 58622 9192
rect 58798 9188 58880 9212
rect 59816 9246 59898 9270
rect 60070 9266 60086 9300
rect 60642 9266 60658 9300
rect 59816 9212 59840 9246
rect 59874 9212 59898 9246
rect 59052 9158 59068 9192
rect 59624 9158 59640 9192
rect 59816 9188 59898 9212
rect 60834 9246 60916 9270
rect 61088 9266 61104 9300
rect 61660 9266 61676 9300
rect 60834 9212 60858 9246
rect 60892 9212 60916 9246
rect 60070 9158 60086 9192
rect 60642 9158 60658 9192
rect 60834 9188 60916 9212
rect 61852 9246 61934 9270
rect 62106 9266 62122 9300
rect 62678 9266 62694 9300
rect 61852 9212 61876 9246
rect 61910 9212 61934 9246
rect 61088 9158 61104 9192
rect 61660 9158 61676 9192
rect 61852 9188 61934 9212
rect 62870 9246 62952 9270
rect 63124 9266 63140 9300
rect 63696 9266 63712 9300
rect 62870 9212 62894 9246
rect 62928 9212 62952 9246
rect 62106 9158 62122 9192
rect 62678 9158 62694 9192
rect 62870 9188 62952 9212
rect 63888 9246 63970 9270
rect 64142 9266 64158 9300
rect 64714 9266 64730 9300
rect 67530 9284 67564 9300
rect 68548 9876 68582 9892
rect 68548 9284 68582 9300
rect 69566 9876 69600 9892
rect 69566 9284 69600 9300
rect 70584 9876 70618 9892
rect 70584 9284 70618 9300
rect 71602 9876 71636 9892
rect 71602 9284 71636 9300
rect 72620 9876 72654 9892
rect 72620 9284 72654 9300
rect 73638 9876 73672 9892
rect 73638 9284 73672 9300
rect 74656 9876 74690 9892
rect 74656 9284 74690 9300
rect 75674 9876 75708 9892
rect 75674 9284 75708 9300
rect 76692 9876 76726 9892
rect 76692 9284 76726 9300
rect 77710 9876 77744 9892
rect 77710 9284 77744 9300
rect 78728 9876 78762 9892
rect 78728 9284 78762 9300
rect 79746 9876 79780 9892
rect 79746 9284 79780 9300
rect 80764 9876 80798 9892
rect 80764 9284 80798 9300
rect 81782 9876 81816 9892
rect 81782 9284 81816 9300
rect 82800 9876 82834 9892
rect 82800 9284 82834 9300
rect 83818 9876 83852 9892
rect 83818 9284 83852 9300
rect 84836 9876 84870 9892
rect 84836 9284 84870 9300
rect 85854 9876 85888 9892
rect 85854 9284 85888 9300
rect 86872 9876 86906 9892
rect 86872 9284 86906 9300
rect 87890 9876 87924 9892
rect 87890 9284 87924 9300
rect 63888 9212 63912 9246
rect 63946 9212 63970 9246
rect 63124 9158 63140 9192
rect 63696 9158 63712 9192
rect 63888 9188 63970 9212
rect 64906 9246 64988 9270
rect 64906 9212 64930 9246
rect 64964 9212 64988 9246
rect 67762 9216 67778 9250
rect 68334 9216 68350 9250
rect 68780 9216 68796 9250
rect 69352 9216 69368 9250
rect 69798 9216 69814 9250
rect 70370 9216 70386 9250
rect 70816 9216 70832 9250
rect 71388 9216 71404 9250
rect 71834 9216 71850 9250
rect 72406 9216 72422 9250
rect 72852 9216 72868 9250
rect 73424 9216 73440 9250
rect 73870 9216 73886 9250
rect 74442 9216 74458 9250
rect 74888 9216 74904 9250
rect 75460 9216 75476 9250
rect 75906 9216 75922 9250
rect 76478 9216 76494 9250
rect 76924 9216 76940 9250
rect 77496 9216 77512 9250
rect 77942 9216 77958 9250
rect 78514 9216 78530 9250
rect 78960 9216 78976 9250
rect 79532 9216 79548 9250
rect 79978 9216 79994 9250
rect 80550 9216 80566 9250
rect 80996 9216 81012 9250
rect 81568 9216 81584 9250
rect 82014 9216 82030 9250
rect 82586 9216 82602 9250
rect 83032 9216 83048 9250
rect 83604 9216 83620 9250
rect 84050 9216 84066 9250
rect 84622 9216 84638 9250
rect 85068 9216 85084 9250
rect 85640 9216 85656 9250
rect 86086 9216 86102 9250
rect 86658 9216 86674 9250
rect 87104 9216 87120 9250
rect 87676 9216 87692 9250
rect 64142 9158 64158 9192
rect 64714 9158 64730 9192
rect 64906 9188 64988 9212
rect 55766 9108 55800 9124
rect 55766 8516 55800 8532
rect 56784 9108 56818 9124
rect 56784 8516 56818 8532
rect 57802 9108 57836 9124
rect 57802 8516 57836 8532
rect 58820 9108 58854 9124
rect 58820 8516 58854 8532
rect 59838 9108 59872 9124
rect 59838 8516 59872 8532
rect 60856 9108 60890 9124
rect 60856 8516 60890 8532
rect 61874 9108 61908 9124
rect 61874 8516 61908 8532
rect 62892 9108 62926 9124
rect 62892 8516 62926 8532
rect 63910 9108 63944 9124
rect 63910 8516 63944 8532
rect 64928 9108 64962 9124
rect 68030 8988 68112 9012
rect 68030 8954 68054 8988
rect 68088 8954 68112 8988
rect 68030 8930 68112 8954
rect 69048 8988 69130 9012
rect 69048 8954 69072 8988
rect 69106 8954 69130 8988
rect 69048 8930 69130 8954
rect 70066 8988 70148 9012
rect 70066 8954 70090 8988
rect 70124 8954 70148 8988
rect 70066 8930 70148 8954
rect 71084 8988 71166 9012
rect 71084 8954 71108 8988
rect 71142 8954 71166 8988
rect 71084 8930 71166 8954
rect 72102 8988 72184 9012
rect 72102 8954 72126 8988
rect 72160 8954 72184 8988
rect 72102 8930 72184 8954
rect 73120 8988 73202 9012
rect 73120 8954 73144 8988
rect 73178 8954 73202 8988
rect 73120 8930 73202 8954
rect 74138 8988 74220 9012
rect 74138 8954 74162 8988
rect 74196 8954 74220 8988
rect 74138 8930 74220 8954
rect 75156 8988 75238 9012
rect 75156 8954 75180 8988
rect 75214 8954 75238 8988
rect 75156 8930 75238 8954
rect 76174 8988 76256 9012
rect 76174 8954 76198 8988
rect 76232 8954 76256 8988
rect 76174 8930 76256 8954
rect 77192 8988 77274 9012
rect 77192 8954 77216 8988
rect 77250 8954 77274 8988
rect 77192 8930 77274 8954
rect 78210 8988 78292 9012
rect 78210 8954 78234 8988
rect 78268 8954 78292 8988
rect 78210 8930 78292 8954
rect 79228 8988 79310 9012
rect 79228 8954 79252 8988
rect 79286 8954 79310 8988
rect 79228 8930 79310 8954
rect 80246 8988 80328 9012
rect 80246 8954 80270 8988
rect 80304 8954 80328 8988
rect 80246 8930 80328 8954
rect 81264 8988 81346 9012
rect 81264 8954 81288 8988
rect 81322 8954 81346 8988
rect 81264 8930 81346 8954
rect 82282 8988 82364 9012
rect 82282 8954 82306 8988
rect 82340 8954 82364 8988
rect 82282 8930 82364 8954
rect 83300 8988 83382 9012
rect 83300 8954 83324 8988
rect 83358 8954 83382 8988
rect 83300 8930 83382 8954
rect 84318 8988 84400 9012
rect 84318 8954 84342 8988
rect 84376 8954 84400 8988
rect 84318 8930 84400 8954
rect 85336 8988 85418 9012
rect 85336 8954 85360 8988
rect 85394 8954 85418 8988
rect 85336 8930 85418 8954
rect 86354 8988 86436 9012
rect 86354 8954 86378 8988
rect 86412 8954 86436 8988
rect 86354 8930 86436 8954
rect 87372 8988 87454 9012
rect 87372 8954 87396 8988
rect 87430 8954 87454 8988
rect 87372 8930 87454 8954
rect 67762 8694 67778 8728
rect 68334 8694 68350 8728
rect 68780 8694 68796 8728
rect 69352 8694 69368 8728
rect 69798 8694 69814 8728
rect 70370 8694 70386 8728
rect 70816 8694 70832 8728
rect 71388 8694 71404 8728
rect 71834 8694 71850 8728
rect 72406 8694 72422 8728
rect 72852 8694 72868 8728
rect 73424 8694 73440 8728
rect 73870 8694 73886 8728
rect 74442 8694 74458 8728
rect 74888 8694 74904 8728
rect 75460 8694 75476 8728
rect 75906 8694 75922 8728
rect 76478 8694 76494 8728
rect 76924 8694 76940 8728
rect 77496 8694 77512 8728
rect 77942 8694 77958 8728
rect 78514 8694 78530 8728
rect 78960 8694 78976 8728
rect 79532 8694 79548 8728
rect 79978 8694 79994 8728
rect 80550 8694 80566 8728
rect 80996 8694 81012 8728
rect 81568 8694 81584 8728
rect 82014 8694 82030 8728
rect 82586 8694 82602 8728
rect 83032 8694 83048 8728
rect 83604 8694 83620 8728
rect 84050 8694 84066 8728
rect 84622 8694 84638 8728
rect 85068 8694 85084 8728
rect 85640 8694 85656 8728
rect 86086 8694 86102 8728
rect 86658 8694 86674 8728
rect 87104 8694 87120 8728
rect 87676 8694 87692 8728
rect 64928 8516 64962 8532
rect 67530 8644 67564 8660
rect 56258 8482 56318 8484
rect 57284 8482 57344 8486
rect 58298 8482 58358 8486
rect 59318 8482 59378 8484
rect 60340 8482 60400 8484
rect 62372 8482 62432 8486
rect 63388 8482 63448 8486
rect 64408 8482 64468 8484
rect 55744 8428 55826 8452
rect 55998 8448 56014 8482
rect 56570 8448 56586 8482
rect 55744 8394 55768 8428
rect 55802 8394 55826 8428
rect 55744 8370 55826 8394
rect 56762 8428 56844 8452
rect 57016 8448 57032 8482
rect 57588 8448 57604 8482
rect 56762 8394 56786 8428
rect 56820 8394 56844 8428
rect 55998 8340 56014 8374
rect 56570 8340 56586 8374
rect 56762 8370 56844 8394
rect 57780 8428 57862 8452
rect 58034 8448 58050 8482
rect 58606 8448 58622 8482
rect 57780 8394 57804 8428
rect 57838 8394 57862 8428
rect 57016 8340 57032 8374
rect 57588 8340 57604 8374
rect 57780 8370 57862 8394
rect 58798 8428 58880 8452
rect 59052 8448 59068 8482
rect 59624 8448 59640 8482
rect 58798 8394 58822 8428
rect 58856 8394 58880 8428
rect 58034 8340 58050 8374
rect 58606 8340 58622 8374
rect 58798 8370 58880 8394
rect 59816 8428 59898 8452
rect 60070 8448 60086 8482
rect 60642 8448 60658 8482
rect 59816 8394 59840 8428
rect 59874 8394 59898 8428
rect 59052 8340 59068 8374
rect 59624 8340 59640 8374
rect 59816 8370 59898 8394
rect 60834 8428 60916 8452
rect 61088 8448 61104 8482
rect 61660 8448 61676 8482
rect 60834 8394 60858 8428
rect 60892 8394 60916 8428
rect 60070 8340 60086 8374
rect 60642 8340 60658 8374
rect 60834 8370 60916 8394
rect 61852 8428 61934 8452
rect 62106 8448 62122 8482
rect 62678 8448 62694 8482
rect 61852 8394 61876 8428
rect 61910 8394 61934 8428
rect 61088 8340 61104 8374
rect 61660 8340 61676 8374
rect 61852 8370 61934 8394
rect 62870 8428 62952 8452
rect 63124 8448 63140 8482
rect 63696 8448 63712 8482
rect 62870 8394 62894 8428
rect 62928 8394 62952 8428
rect 62106 8340 62122 8374
rect 62678 8340 62694 8374
rect 62870 8370 62952 8394
rect 63888 8428 63970 8452
rect 64142 8448 64158 8482
rect 64714 8448 64730 8482
rect 63888 8394 63912 8428
rect 63946 8394 63970 8428
rect 63124 8340 63140 8374
rect 63696 8340 63712 8374
rect 63888 8370 63970 8394
rect 64906 8428 64988 8452
rect 64906 8394 64930 8428
rect 64964 8394 64988 8428
rect 64142 8340 64158 8374
rect 64714 8340 64730 8374
rect 64906 8370 64988 8394
rect 55766 8290 55800 8306
rect 55766 7698 55800 7714
rect 56784 8290 56818 8306
rect 56784 7698 56818 7714
rect 57802 8290 57836 8306
rect 57802 7698 57836 7714
rect 58820 8290 58854 8306
rect 58820 7698 58854 7714
rect 59838 8290 59872 8306
rect 59838 7698 59872 7714
rect 60856 8290 60890 8306
rect 60856 7698 60890 7714
rect 61874 8290 61908 8306
rect 61874 7698 61908 7714
rect 62892 8290 62926 8306
rect 62892 7698 62926 7714
rect 63910 8290 63944 8306
rect 63910 7698 63944 7714
rect 64928 8290 64962 8306
rect 67530 8052 67564 8068
rect 68548 8644 68582 8660
rect 68548 8052 68582 8068
rect 69566 8644 69600 8660
rect 69566 8052 69600 8068
rect 70584 8644 70618 8660
rect 70584 8052 70618 8068
rect 71602 8644 71636 8660
rect 71602 8052 71636 8068
rect 72620 8644 72654 8660
rect 72620 8052 72654 8068
rect 73638 8644 73672 8660
rect 73638 8052 73672 8068
rect 74656 8644 74690 8660
rect 74656 8052 74690 8068
rect 75674 8644 75708 8660
rect 75674 8052 75708 8068
rect 76692 8644 76726 8660
rect 76692 8052 76726 8068
rect 77710 8644 77744 8660
rect 77710 8052 77744 8068
rect 78728 8644 78762 8660
rect 78728 8052 78762 8068
rect 79746 8644 79780 8660
rect 79746 8052 79780 8068
rect 80764 8644 80798 8660
rect 80764 8052 80798 8068
rect 81782 8644 81816 8660
rect 81782 8052 81816 8068
rect 82800 8644 82834 8660
rect 82800 8052 82834 8068
rect 83818 8644 83852 8660
rect 83818 8052 83852 8068
rect 84836 8644 84870 8660
rect 84836 8052 84870 8068
rect 85854 8644 85888 8660
rect 85854 8052 85888 8068
rect 86872 8644 86906 8660
rect 86872 8052 86906 8068
rect 87890 8644 87924 8660
rect 87890 8052 87924 8068
rect 76180 8018 76240 8020
rect 78224 8018 78284 8022
rect 86358 8018 86418 8020
rect 67762 7984 67778 8018
rect 68334 7984 68350 8018
rect 68780 7984 68796 8018
rect 69352 7984 69368 8018
rect 69798 7984 69814 8018
rect 70370 7984 70386 8018
rect 70816 7984 70832 8018
rect 71388 7984 71404 8018
rect 71834 7984 71850 8018
rect 72406 7984 72422 8018
rect 72852 7984 72868 8018
rect 73424 7984 73440 8018
rect 73870 7984 73886 8018
rect 74442 7984 74458 8018
rect 74888 7984 74904 8018
rect 75460 7984 75476 8018
rect 75906 7984 75922 8018
rect 76478 7984 76494 8018
rect 76924 7984 76940 8018
rect 77496 7984 77512 8018
rect 77942 7984 77958 8018
rect 78514 7984 78530 8018
rect 78960 7984 78976 8018
rect 79532 7984 79548 8018
rect 79978 7984 79994 8018
rect 80550 7984 80566 8018
rect 80996 7984 81012 8018
rect 81568 7984 81584 8018
rect 82014 7984 82030 8018
rect 82586 7984 82602 8018
rect 83032 7984 83048 8018
rect 83604 7984 83620 8018
rect 84050 7984 84066 8018
rect 84622 7984 84638 8018
rect 85068 7984 85084 8018
rect 85640 7984 85656 8018
rect 86086 7984 86102 8018
rect 86658 7984 86674 8018
rect 87104 7984 87120 8018
rect 87676 7984 87692 8018
rect 64928 7698 64962 7714
rect 68016 7766 68098 7790
rect 68016 7732 68040 7766
rect 68074 7732 68098 7766
rect 68016 7708 68098 7732
rect 69034 7766 69116 7790
rect 69034 7732 69058 7766
rect 69092 7732 69116 7766
rect 69034 7708 69116 7732
rect 70052 7766 70134 7790
rect 70052 7732 70076 7766
rect 70110 7732 70134 7766
rect 70052 7708 70134 7732
rect 71070 7766 71152 7790
rect 71070 7732 71094 7766
rect 71128 7732 71152 7766
rect 71070 7708 71152 7732
rect 72088 7766 72170 7790
rect 72088 7732 72112 7766
rect 72146 7732 72170 7766
rect 72088 7708 72170 7732
rect 73106 7766 73188 7790
rect 73106 7732 73130 7766
rect 73164 7732 73188 7766
rect 73106 7708 73188 7732
rect 74124 7766 74206 7790
rect 74124 7732 74148 7766
rect 74182 7732 74206 7766
rect 74124 7708 74206 7732
rect 75142 7766 75224 7790
rect 75142 7732 75166 7766
rect 75200 7732 75224 7766
rect 75142 7708 75224 7732
rect 76160 7766 76242 7790
rect 76160 7732 76184 7766
rect 76218 7732 76242 7766
rect 76160 7708 76242 7732
rect 77178 7766 77260 7790
rect 77178 7732 77202 7766
rect 77236 7732 77260 7766
rect 77178 7708 77260 7732
rect 78196 7766 78278 7790
rect 78196 7732 78220 7766
rect 78254 7732 78278 7766
rect 78196 7708 78278 7732
rect 79214 7766 79296 7790
rect 79214 7732 79238 7766
rect 79272 7732 79296 7766
rect 79214 7708 79296 7732
rect 80232 7766 80314 7790
rect 80232 7732 80256 7766
rect 80290 7732 80314 7766
rect 80232 7708 80314 7732
rect 81250 7766 81332 7790
rect 81250 7732 81274 7766
rect 81308 7732 81332 7766
rect 81250 7708 81332 7732
rect 82268 7766 82350 7790
rect 82268 7732 82292 7766
rect 82326 7732 82350 7766
rect 82268 7708 82350 7732
rect 83286 7766 83368 7790
rect 83286 7732 83310 7766
rect 83344 7732 83368 7766
rect 83286 7708 83368 7732
rect 84304 7766 84386 7790
rect 84304 7732 84328 7766
rect 84362 7732 84386 7766
rect 84304 7708 84386 7732
rect 85322 7766 85404 7790
rect 85322 7732 85346 7766
rect 85380 7732 85404 7766
rect 85322 7708 85404 7732
rect 86340 7766 86422 7790
rect 86340 7732 86364 7766
rect 86398 7732 86422 7766
rect 86340 7708 86422 7732
rect 87358 7766 87440 7790
rect 87358 7732 87382 7766
rect 87416 7732 87440 7766
rect 87358 7708 87440 7732
rect 55998 7630 56014 7664
rect 56570 7630 56586 7664
rect 57016 7630 57032 7664
rect 57588 7630 57604 7664
rect 58034 7630 58050 7664
rect 58606 7630 58622 7664
rect 59052 7630 59068 7664
rect 59624 7630 59640 7664
rect 60070 7630 60086 7664
rect 60642 7630 60658 7664
rect 61088 7630 61104 7664
rect 61660 7630 61676 7664
rect 62106 7630 62122 7664
rect 62678 7630 62694 7664
rect 63124 7630 63140 7664
rect 63696 7630 63712 7664
rect 64142 7630 64158 7664
rect 64714 7630 64730 7664
rect 67762 7460 67778 7494
rect 68334 7460 68350 7494
rect 68780 7460 68796 7494
rect 69352 7460 69368 7494
rect 69798 7460 69814 7494
rect 70370 7460 70386 7494
rect 70816 7460 70832 7494
rect 71388 7460 71404 7494
rect 71834 7460 71850 7494
rect 72406 7460 72422 7494
rect 72852 7460 72868 7494
rect 73424 7460 73440 7494
rect 73870 7460 73886 7494
rect 74442 7460 74458 7494
rect 74888 7460 74904 7494
rect 75460 7460 75476 7494
rect 75906 7460 75922 7494
rect 76478 7460 76494 7494
rect 76924 7460 76940 7494
rect 77496 7460 77512 7494
rect 77942 7460 77958 7494
rect 78514 7460 78530 7494
rect 78960 7460 78976 7494
rect 79532 7460 79548 7494
rect 79978 7460 79994 7494
rect 80550 7460 80566 7494
rect 80996 7460 81012 7494
rect 81568 7460 81584 7494
rect 82014 7460 82030 7494
rect 82586 7460 82602 7494
rect 83032 7460 83048 7494
rect 83604 7460 83620 7494
rect 84050 7460 84066 7494
rect 84622 7460 84638 7494
rect 85068 7460 85084 7494
rect 85640 7460 85656 7494
rect 86086 7460 86102 7494
rect 86658 7460 86674 7494
rect 87104 7460 87120 7494
rect 87676 7460 87692 7494
rect 67530 7410 67564 7426
rect 56254 7386 56336 7410
rect 56254 7352 56278 7386
rect 56312 7352 56336 7386
rect 56254 7328 56336 7352
rect 57272 7386 57354 7410
rect 57272 7352 57296 7386
rect 57330 7352 57354 7386
rect 57272 7328 57354 7352
rect 58290 7386 58372 7410
rect 58290 7352 58314 7386
rect 58348 7352 58372 7386
rect 58290 7328 58372 7352
rect 59308 7386 59390 7410
rect 59308 7352 59332 7386
rect 59366 7352 59390 7386
rect 59308 7328 59390 7352
rect 60326 7386 60408 7410
rect 60326 7352 60350 7386
rect 60384 7352 60408 7386
rect 60326 7328 60408 7352
rect 61344 7386 61426 7410
rect 61344 7352 61368 7386
rect 61402 7352 61426 7386
rect 61344 7328 61426 7352
rect 62362 7386 62444 7410
rect 62362 7352 62386 7386
rect 62420 7352 62444 7386
rect 62362 7328 62444 7352
rect 63380 7386 63462 7410
rect 63380 7352 63404 7386
rect 63438 7352 63462 7386
rect 63380 7328 63462 7352
rect 64398 7386 64480 7410
rect 64398 7352 64422 7386
rect 64456 7352 64480 7386
rect 64398 7328 64480 7352
rect 62698 6956 62714 6990
rect 62790 6956 62806 6990
rect 62916 6956 62932 6990
rect 63008 6956 63024 6990
rect 63134 6956 63150 6990
rect 63226 6956 63242 6990
rect 63352 6956 63368 6990
rect 63444 6956 63460 6990
rect 63570 6956 63586 6990
rect 63662 6956 63678 6990
rect 63788 6956 63804 6990
rect 63880 6956 63896 6990
rect 64006 6956 64022 6990
rect 64098 6956 64114 6990
rect 64224 6956 64240 6990
rect 64316 6956 64332 6990
rect 64442 6956 64458 6990
rect 64534 6956 64550 6990
rect 64660 6956 64676 6990
rect 64752 6956 64768 6990
rect 62626 6906 62660 6922
rect 62626 6714 62660 6730
rect 62844 6906 62878 6922
rect 62844 6714 62878 6730
rect 63062 6906 63096 6922
rect 63062 6714 63096 6730
rect 63280 6906 63314 6922
rect 63280 6714 63314 6730
rect 63498 6906 63532 6922
rect 63498 6714 63532 6730
rect 63716 6906 63750 6922
rect 63716 6714 63750 6730
rect 63934 6906 63968 6922
rect 63934 6714 63968 6730
rect 64152 6906 64186 6922
rect 64152 6714 64186 6730
rect 64370 6906 64404 6922
rect 64370 6714 64404 6730
rect 64588 6906 64622 6922
rect 64588 6714 64622 6730
rect 64806 6906 64840 6922
rect 67530 6818 67564 6834
rect 68548 7410 68582 7426
rect 68548 6818 68582 6834
rect 69566 7410 69600 7426
rect 69566 6818 69600 6834
rect 70584 7410 70618 7426
rect 70584 6818 70618 6834
rect 71602 7410 71636 7426
rect 71602 6818 71636 6834
rect 72620 7410 72654 7426
rect 72620 6818 72654 6834
rect 73638 7410 73672 7426
rect 73638 6818 73672 6834
rect 74656 7410 74690 7426
rect 74656 6818 74690 6834
rect 75674 7410 75708 7426
rect 75674 6818 75708 6834
rect 76692 7410 76726 7426
rect 76692 6818 76726 6834
rect 77710 7410 77744 7426
rect 77710 6818 77744 6834
rect 78728 7410 78762 7426
rect 78728 6818 78762 6834
rect 79746 7410 79780 7426
rect 79746 6818 79780 6834
rect 80764 7410 80798 7426
rect 80764 6818 80798 6834
rect 81782 7410 81816 7426
rect 81782 6818 81816 6834
rect 82800 7410 82834 7426
rect 82800 6818 82834 6834
rect 83818 7410 83852 7426
rect 83818 6818 83852 6834
rect 84836 7410 84870 7426
rect 84836 6818 84870 6834
rect 85854 7410 85888 7426
rect 85854 6818 85888 6834
rect 86872 7410 86906 7426
rect 86872 6818 86906 6834
rect 87890 7410 87924 7426
rect 87890 6818 87924 6834
rect 70056 6784 70116 6788
rect 67762 6750 67778 6784
rect 68334 6750 68350 6784
rect 68780 6750 68796 6784
rect 69352 6750 69368 6784
rect 69798 6750 69814 6784
rect 70370 6750 70386 6784
rect 70816 6750 70832 6784
rect 71388 6750 71404 6784
rect 71834 6750 71850 6784
rect 72406 6750 72422 6784
rect 72852 6750 72868 6784
rect 73424 6750 73440 6784
rect 73870 6750 73886 6784
rect 74442 6750 74458 6784
rect 74888 6750 74904 6784
rect 75460 6750 75476 6784
rect 75906 6750 75922 6784
rect 76478 6750 76494 6784
rect 76924 6750 76940 6784
rect 77496 6750 77512 6784
rect 77942 6750 77958 6784
rect 78514 6750 78530 6784
rect 78960 6750 78976 6784
rect 79532 6750 79548 6784
rect 79978 6750 79994 6784
rect 80550 6750 80566 6784
rect 80996 6750 81012 6784
rect 81568 6750 81584 6784
rect 82014 6750 82030 6784
rect 82586 6750 82602 6784
rect 83032 6750 83048 6784
rect 83604 6750 83620 6784
rect 84050 6750 84066 6784
rect 84622 6750 84638 6784
rect 85068 6750 85084 6784
rect 85640 6750 85656 6784
rect 86086 6750 86102 6784
rect 86658 6750 86674 6784
rect 87104 6750 87120 6784
rect 87676 6750 87692 6784
rect 64806 6714 64840 6730
rect 62698 6646 62714 6680
rect 62790 6646 62806 6680
rect 62916 6646 62932 6680
rect 63008 6646 63024 6680
rect 63134 6646 63150 6680
rect 63226 6646 63242 6680
rect 63352 6646 63368 6680
rect 63444 6646 63460 6680
rect 63570 6646 63586 6680
rect 63662 6646 63678 6680
rect 63788 6646 63804 6680
rect 63880 6646 63896 6680
rect 64006 6646 64022 6680
rect 64098 6646 64114 6680
rect 64224 6646 64240 6680
rect 64316 6646 64332 6680
rect 64442 6646 64458 6680
rect 64534 6646 64550 6680
rect 64660 6646 64676 6680
rect 64752 6646 64768 6680
rect 68016 6518 68098 6542
rect 68016 6484 68040 6518
rect 68074 6484 68098 6518
rect 68016 6460 68098 6484
rect 69034 6518 69116 6542
rect 69034 6484 69058 6518
rect 69092 6484 69116 6518
rect 69034 6460 69116 6484
rect 70052 6518 70134 6542
rect 70052 6484 70076 6518
rect 70110 6484 70134 6518
rect 70052 6460 70134 6484
rect 71070 6518 71152 6542
rect 71070 6484 71094 6518
rect 71128 6484 71152 6518
rect 71070 6460 71152 6484
rect 72088 6518 72170 6542
rect 72088 6484 72112 6518
rect 72146 6484 72170 6518
rect 72088 6460 72170 6484
rect 73106 6518 73188 6542
rect 73106 6484 73130 6518
rect 73164 6484 73188 6518
rect 73106 6460 73188 6484
rect 74124 6518 74206 6542
rect 74124 6484 74148 6518
rect 74182 6484 74206 6518
rect 74124 6460 74206 6484
rect 75142 6518 75224 6542
rect 75142 6484 75166 6518
rect 75200 6484 75224 6518
rect 75142 6460 75224 6484
rect 76160 6518 76242 6542
rect 76160 6484 76184 6518
rect 76218 6484 76242 6518
rect 76160 6460 76242 6484
rect 77178 6518 77260 6542
rect 77178 6484 77202 6518
rect 77236 6484 77260 6518
rect 77178 6460 77260 6484
rect 78196 6518 78278 6542
rect 78196 6484 78220 6518
rect 78254 6484 78278 6518
rect 78196 6460 78278 6484
rect 79214 6518 79296 6542
rect 79214 6484 79238 6518
rect 79272 6484 79296 6518
rect 79214 6460 79296 6484
rect 80232 6518 80314 6542
rect 80232 6484 80256 6518
rect 80290 6484 80314 6518
rect 80232 6460 80314 6484
rect 81250 6518 81332 6542
rect 81250 6484 81274 6518
rect 81308 6484 81332 6518
rect 81250 6460 81332 6484
rect 82268 6518 82350 6542
rect 82268 6484 82292 6518
rect 82326 6484 82350 6518
rect 82268 6460 82350 6484
rect 83286 6518 83368 6542
rect 83286 6484 83310 6518
rect 83344 6484 83368 6518
rect 83286 6460 83368 6484
rect 84304 6518 84386 6542
rect 84304 6484 84328 6518
rect 84362 6484 84386 6518
rect 84304 6460 84386 6484
rect 85322 6518 85404 6542
rect 85322 6484 85346 6518
rect 85380 6484 85404 6518
rect 85322 6460 85404 6484
rect 86340 6518 86422 6542
rect 86340 6484 86364 6518
rect 86398 6484 86422 6518
rect 86340 6460 86422 6484
rect 87358 6518 87440 6542
rect 87358 6484 87382 6518
rect 87416 6484 87440 6518
rect 87358 6460 87440 6484
rect 62332 6410 62414 6434
rect 62332 6376 62356 6410
rect 62390 6376 62414 6410
rect 62332 6352 62414 6376
rect 63350 6410 63432 6434
rect 63350 6376 63374 6410
rect 63408 6376 63432 6410
rect 63350 6352 63432 6376
rect 64368 6410 64450 6434
rect 64368 6376 64392 6410
rect 64426 6376 64450 6410
rect 64368 6352 64450 6376
rect 65386 6410 65468 6434
rect 65386 6376 65410 6410
rect 65444 6376 65468 6410
rect 65386 6352 65468 6376
rect 67762 6226 67778 6260
rect 68334 6226 68350 6260
rect 68780 6226 68796 6260
rect 69352 6226 69368 6260
rect 69798 6226 69814 6260
rect 70370 6226 70386 6260
rect 70816 6226 70832 6260
rect 71388 6226 71404 6260
rect 71834 6226 71850 6260
rect 72406 6226 72422 6260
rect 72852 6226 72868 6260
rect 73424 6226 73440 6260
rect 73870 6226 73886 6260
rect 74442 6226 74458 6260
rect 74888 6226 74904 6260
rect 75460 6226 75476 6260
rect 75906 6226 75922 6260
rect 76478 6226 76494 6260
rect 76924 6226 76940 6260
rect 77496 6226 77512 6260
rect 77942 6226 77958 6260
rect 78514 6226 78530 6260
rect 78960 6226 78976 6260
rect 79532 6226 79548 6260
rect 79978 6226 79994 6260
rect 80550 6226 80566 6260
rect 80996 6226 81012 6260
rect 81568 6226 81584 6260
rect 82014 6226 82030 6260
rect 82586 6226 82602 6260
rect 83032 6226 83048 6260
rect 83604 6226 83620 6260
rect 84050 6226 84066 6260
rect 84622 6226 84638 6260
rect 85068 6226 85084 6260
rect 85640 6226 85656 6260
rect 86086 6226 86102 6260
rect 86658 6226 86674 6260
rect 87104 6226 87120 6260
rect 87676 6226 87692 6260
rect 67530 6176 67564 6192
rect 62698 6124 62714 6158
rect 62790 6124 62806 6158
rect 62916 6124 62932 6158
rect 63008 6124 63024 6158
rect 63134 6124 63150 6158
rect 63226 6124 63242 6158
rect 63352 6124 63368 6158
rect 63444 6124 63460 6158
rect 63570 6124 63586 6158
rect 63662 6124 63678 6158
rect 63788 6124 63804 6158
rect 63880 6124 63896 6158
rect 64006 6124 64022 6158
rect 64098 6124 64114 6158
rect 64224 6124 64240 6158
rect 64316 6124 64332 6158
rect 64442 6124 64458 6158
rect 64534 6124 64550 6158
rect 64660 6124 64676 6158
rect 64752 6124 64768 6158
rect 62626 6074 62660 6090
rect 62626 5882 62660 5898
rect 62844 6074 62878 6090
rect 62844 5882 62878 5898
rect 63062 6074 63096 6090
rect 63062 5882 63096 5898
rect 63280 6074 63314 6090
rect 63280 5882 63314 5898
rect 63498 6074 63532 6090
rect 63498 5882 63532 5898
rect 63716 6074 63750 6090
rect 63716 5882 63750 5898
rect 63934 6074 63968 6090
rect 63934 5882 63968 5898
rect 64152 6074 64186 6090
rect 64152 5882 64186 5898
rect 64370 6074 64404 6090
rect 64370 5882 64404 5898
rect 64588 6074 64622 6090
rect 64588 5882 64622 5898
rect 64806 6074 64840 6090
rect 64806 5882 64840 5898
rect 62698 5814 62714 5848
rect 62790 5814 62806 5848
rect 62916 5814 62932 5848
rect 63008 5814 63024 5848
rect 63134 5814 63150 5848
rect 63226 5814 63242 5848
rect 63352 5814 63368 5848
rect 63444 5814 63460 5848
rect 63570 5814 63586 5848
rect 63662 5814 63678 5848
rect 63788 5814 63804 5848
rect 63880 5814 63896 5848
rect 64006 5814 64022 5848
rect 64098 5814 64114 5848
rect 64224 5814 64240 5848
rect 64316 5814 64332 5848
rect 64442 5814 64458 5848
rect 64534 5814 64550 5848
rect 64660 5814 64676 5848
rect 64752 5814 64768 5848
rect 67530 5584 67564 5600
rect 68548 6176 68582 6192
rect 68548 5584 68582 5600
rect 69566 6176 69600 6192
rect 69566 5584 69600 5600
rect 70584 6176 70618 6192
rect 70584 5584 70618 5600
rect 71602 6176 71636 6192
rect 71602 5584 71636 5600
rect 72620 6176 72654 6192
rect 72620 5584 72654 5600
rect 73638 6176 73672 6192
rect 73638 5584 73672 5600
rect 74656 6176 74690 6192
rect 74656 5584 74690 5600
rect 75674 6176 75708 6192
rect 75674 5584 75708 5600
rect 76692 6176 76726 6192
rect 76692 5584 76726 5600
rect 77710 6176 77744 6192
rect 77710 5584 77744 5600
rect 78728 6176 78762 6192
rect 78728 5584 78762 5600
rect 79746 6176 79780 6192
rect 79746 5584 79780 5600
rect 80764 6176 80798 6192
rect 80764 5584 80798 5600
rect 81782 6176 81816 6192
rect 81782 5584 81816 5600
rect 82800 6176 82834 6192
rect 82800 5584 82834 5600
rect 83818 6176 83852 6192
rect 83818 5584 83852 5600
rect 84836 6176 84870 6192
rect 84836 5584 84870 5600
rect 85854 6176 85888 6192
rect 85854 5584 85888 5600
rect 86872 6176 86906 6192
rect 86872 5584 86906 5600
rect 87890 6176 87924 6192
rect 87890 5584 87924 5600
rect 76180 5550 76240 5552
rect 78224 5550 78284 5554
rect 81262 5550 81322 5554
rect 67762 5516 67778 5550
rect 68334 5516 68350 5550
rect 68780 5516 68796 5550
rect 69352 5516 69368 5550
rect 69798 5516 69814 5550
rect 70370 5516 70386 5550
rect 70816 5516 70832 5550
rect 71388 5516 71404 5550
rect 71834 5516 71850 5550
rect 72406 5516 72422 5550
rect 72852 5516 72868 5550
rect 73424 5516 73440 5550
rect 73870 5516 73886 5550
rect 74442 5516 74458 5550
rect 74888 5516 74904 5550
rect 75460 5516 75476 5550
rect 75906 5516 75922 5550
rect 76478 5516 76494 5550
rect 76924 5516 76940 5550
rect 77496 5516 77512 5550
rect 77942 5516 77958 5550
rect 78514 5516 78530 5550
rect 78960 5516 78976 5550
rect 79532 5516 79548 5550
rect 79978 5516 79994 5550
rect 80550 5516 80566 5550
rect 80996 5516 81012 5550
rect 81568 5516 81584 5550
rect 82014 5516 82030 5550
rect 82586 5516 82602 5550
rect 83032 5516 83048 5550
rect 83604 5516 83620 5550
rect 84050 5516 84066 5550
rect 84622 5516 84638 5550
rect 85068 5516 85084 5550
rect 85640 5516 85656 5550
rect 86086 5516 86102 5550
rect 86658 5516 86674 5550
rect 87104 5516 87120 5550
rect 87676 5516 87692 5550
rect 68030 5298 68112 5322
rect 68030 5264 68054 5298
rect 68088 5264 68112 5298
rect 68030 5240 68112 5264
rect 69048 5298 69130 5322
rect 69048 5264 69072 5298
rect 69106 5264 69130 5298
rect 69048 5240 69130 5264
rect 70066 5298 70148 5322
rect 70066 5264 70090 5298
rect 70124 5264 70148 5298
rect 70066 5240 70148 5264
rect 71084 5298 71166 5322
rect 71084 5264 71108 5298
rect 71142 5264 71166 5298
rect 71084 5240 71166 5264
rect 72102 5298 72184 5322
rect 72102 5264 72126 5298
rect 72160 5264 72184 5298
rect 72102 5240 72184 5264
rect 73120 5298 73202 5322
rect 73120 5264 73144 5298
rect 73178 5264 73202 5298
rect 73120 5240 73202 5264
rect 74138 5298 74220 5322
rect 74138 5264 74162 5298
rect 74196 5264 74220 5298
rect 74138 5240 74220 5264
rect 75156 5298 75238 5322
rect 75156 5264 75180 5298
rect 75214 5264 75238 5298
rect 75156 5240 75238 5264
rect 76174 5298 76256 5322
rect 76174 5264 76198 5298
rect 76232 5264 76256 5298
rect 76174 5240 76256 5264
rect 77192 5298 77274 5322
rect 77192 5264 77216 5298
rect 77250 5264 77274 5298
rect 77192 5240 77274 5264
rect 78210 5298 78292 5322
rect 78210 5264 78234 5298
rect 78268 5264 78292 5298
rect 78210 5240 78292 5264
rect 79228 5298 79310 5322
rect 79228 5264 79252 5298
rect 79286 5264 79310 5298
rect 79228 5240 79310 5264
rect 80246 5298 80328 5322
rect 80246 5264 80270 5298
rect 80304 5264 80328 5298
rect 80246 5240 80328 5264
rect 81264 5298 81346 5322
rect 81264 5264 81288 5298
rect 81322 5264 81346 5298
rect 81264 5240 81346 5264
rect 82282 5298 82364 5322
rect 82282 5264 82306 5298
rect 82340 5264 82364 5298
rect 82282 5240 82364 5264
rect 83300 5298 83382 5322
rect 83300 5264 83324 5298
rect 83358 5264 83382 5298
rect 83300 5240 83382 5264
rect 84318 5298 84400 5322
rect 84318 5264 84342 5298
rect 84376 5264 84400 5298
rect 84318 5240 84400 5264
rect 85336 5298 85418 5322
rect 85336 5264 85360 5298
rect 85394 5264 85418 5298
rect 85336 5240 85418 5264
rect 86354 5298 86436 5322
rect 86354 5264 86378 5298
rect 86412 5264 86436 5298
rect 86354 5240 86436 5264
rect 87372 5298 87454 5322
rect 87372 5264 87396 5298
rect 87430 5264 87454 5298
rect 87372 5240 87454 5264
rect 62630 5122 62712 5146
rect 56038 5066 56120 5090
rect 56038 5032 56062 5066
rect 56096 5032 56120 5066
rect 56038 5008 56120 5032
rect 57056 5066 57138 5090
rect 57056 5032 57080 5066
rect 57114 5032 57138 5066
rect 57056 5008 57138 5032
rect 58074 5066 58156 5090
rect 58074 5032 58098 5066
rect 58132 5032 58156 5066
rect 58074 5008 58156 5032
rect 59092 5066 59174 5090
rect 59092 5032 59116 5066
rect 59150 5032 59174 5066
rect 59092 5008 59174 5032
rect 60110 5066 60192 5090
rect 60110 5032 60134 5066
rect 60168 5032 60192 5066
rect 60110 5008 60192 5032
rect 61128 5066 61210 5090
rect 61128 5032 61152 5066
rect 61186 5032 61210 5066
rect 62630 5088 62654 5122
rect 62688 5088 62712 5122
rect 62630 5064 62712 5088
rect 63648 5122 63730 5146
rect 63648 5088 63672 5122
rect 63706 5088 63730 5122
rect 63648 5064 63730 5088
rect 64666 5122 64748 5146
rect 64666 5088 64690 5122
rect 64724 5088 64748 5122
rect 64666 5064 64748 5088
rect 65684 5122 65766 5146
rect 65684 5088 65708 5122
rect 65742 5088 65766 5122
rect 65684 5064 65766 5088
rect 61128 5008 61210 5032
rect 67762 4994 67778 5028
rect 68334 4994 68350 5028
rect 68780 4994 68796 5028
rect 69352 4994 69368 5028
rect 69798 4994 69814 5028
rect 70370 4994 70386 5028
rect 70816 4994 70832 5028
rect 71388 4994 71404 5028
rect 71834 4994 71850 5028
rect 72406 4994 72422 5028
rect 72852 4994 72868 5028
rect 73424 4994 73440 5028
rect 73870 4994 73886 5028
rect 74442 4994 74458 5028
rect 74888 4994 74904 5028
rect 75460 4994 75476 5028
rect 75906 4994 75922 5028
rect 76478 4994 76494 5028
rect 76924 4994 76940 5028
rect 77496 4994 77512 5028
rect 77942 4994 77958 5028
rect 78514 4994 78530 5028
rect 78960 4994 78976 5028
rect 79532 4994 79548 5028
rect 79978 4994 79994 5028
rect 80550 4994 80566 5028
rect 80996 4994 81012 5028
rect 81568 4994 81584 5028
rect 82014 4994 82030 5028
rect 82586 4994 82602 5028
rect 83032 4994 83048 5028
rect 83604 4994 83620 5028
rect 84050 4994 84066 5028
rect 84622 4994 84638 5028
rect 85068 4994 85084 5028
rect 85640 4994 85656 5028
rect 86086 4994 86102 5028
rect 86658 4994 86674 5028
rect 87104 4994 87120 5028
rect 87676 4994 87692 5028
rect 71084 4992 71144 4994
rect 67530 4944 67564 4960
rect 55777 4797 55793 4831
rect 56349 4797 56365 4831
rect 56795 4797 56811 4831
rect 57367 4797 57383 4831
rect 57813 4797 57829 4831
rect 58385 4797 58401 4831
rect 58831 4797 58847 4831
rect 59403 4797 59419 4831
rect 59849 4797 59865 4831
rect 60421 4797 60437 4831
rect 60867 4797 60883 4831
rect 61439 4797 61455 4831
rect 62628 4798 62644 4832
rect 62768 4798 62784 4832
rect 62926 4798 62942 4832
rect 63066 4798 63082 4832
rect 63224 4798 63240 4832
rect 63364 4798 63380 4832
rect 63522 4798 63538 4832
rect 63662 4798 63678 4832
rect 63820 4798 63836 4832
rect 63960 4798 63976 4832
rect 64118 4798 64134 4832
rect 64258 4798 64274 4832
rect 64416 4798 64432 4832
rect 64556 4798 64572 4832
rect 64714 4798 64730 4832
rect 64854 4798 64870 4832
rect 65012 4798 65028 4832
rect 65152 4798 65168 4832
rect 65310 4798 65326 4832
rect 65450 4798 65466 4832
rect 65608 4798 65624 4832
rect 65748 4798 65764 4832
rect 55545 4747 55579 4763
rect 55545 4155 55579 4171
rect 56563 4747 56597 4763
rect 56563 4155 56597 4171
rect 57581 4747 57615 4763
rect 57581 4155 57615 4171
rect 58599 4747 58633 4763
rect 58599 4155 58633 4171
rect 59617 4747 59651 4763
rect 59617 4155 59651 4171
rect 60635 4747 60669 4763
rect 60635 4155 60669 4171
rect 61653 4747 61687 4763
rect 61653 4155 61687 4171
rect 62540 4748 62574 4764
rect 62540 4156 62574 4172
rect 62838 4748 62872 4764
rect 62838 4156 62872 4172
rect 63136 4748 63170 4764
rect 63136 4156 63170 4172
rect 63434 4748 63468 4764
rect 63434 4156 63468 4172
rect 63732 4748 63766 4764
rect 63732 4156 63766 4172
rect 64030 4748 64064 4764
rect 64030 4156 64064 4172
rect 64328 4748 64362 4764
rect 64328 4156 64362 4172
rect 64626 4748 64660 4764
rect 64626 4156 64660 4172
rect 64924 4748 64958 4764
rect 64924 4156 64958 4172
rect 65222 4748 65256 4764
rect 65222 4156 65256 4172
rect 65520 4748 65554 4764
rect 65520 4156 65554 4172
rect 65818 4748 65852 4764
rect 67530 4352 67564 4368
rect 68548 4944 68582 4960
rect 68548 4352 68582 4368
rect 69566 4944 69600 4960
rect 69566 4352 69600 4368
rect 70584 4944 70618 4960
rect 70584 4352 70618 4368
rect 71602 4944 71636 4960
rect 71602 4352 71636 4368
rect 72620 4944 72654 4960
rect 72620 4352 72654 4368
rect 73638 4944 73672 4960
rect 73638 4352 73672 4368
rect 74656 4944 74690 4960
rect 74656 4352 74690 4368
rect 75674 4944 75708 4960
rect 75674 4352 75708 4368
rect 76692 4944 76726 4960
rect 76692 4352 76726 4368
rect 77710 4944 77744 4960
rect 77710 4352 77744 4368
rect 78728 4944 78762 4960
rect 78728 4352 78762 4368
rect 79746 4944 79780 4960
rect 79746 4352 79780 4368
rect 80764 4944 80798 4960
rect 80764 4352 80798 4368
rect 81782 4944 81816 4960
rect 81782 4352 81816 4368
rect 82800 4944 82834 4960
rect 82800 4352 82834 4368
rect 83818 4944 83852 4960
rect 83818 4352 83852 4368
rect 84836 4944 84870 4960
rect 84836 4352 84870 4368
rect 85854 4944 85888 4960
rect 85854 4352 85888 4368
rect 86872 4944 86906 4960
rect 86872 4352 86906 4368
rect 87890 4944 87924 4960
rect 87890 4352 87924 4368
rect 75156 4318 75216 4328
rect 67762 4284 67778 4318
rect 68334 4284 68350 4318
rect 68780 4284 68796 4318
rect 69352 4284 69368 4318
rect 69798 4284 69814 4318
rect 70370 4284 70386 4318
rect 70816 4284 70832 4318
rect 71388 4284 71404 4318
rect 71834 4284 71850 4318
rect 72406 4284 72422 4318
rect 72852 4284 72868 4318
rect 73424 4284 73440 4318
rect 73870 4284 73886 4318
rect 74442 4284 74458 4318
rect 74888 4284 74904 4318
rect 75460 4284 75476 4318
rect 75906 4284 75922 4318
rect 76478 4284 76494 4318
rect 76924 4284 76940 4318
rect 77496 4284 77512 4318
rect 77942 4284 77958 4318
rect 78514 4284 78530 4318
rect 78960 4284 78976 4318
rect 79532 4284 79548 4318
rect 79978 4284 79994 4318
rect 80550 4284 80566 4318
rect 80996 4284 81012 4318
rect 81568 4284 81584 4318
rect 82014 4284 82030 4318
rect 82586 4284 82602 4318
rect 83032 4284 83048 4318
rect 83604 4284 83620 4318
rect 84050 4284 84066 4318
rect 84622 4284 84638 4318
rect 85068 4284 85084 4318
rect 85640 4284 85656 4318
rect 86086 4284 86102 4318
rect 86658 4284 86674 4318
rect 87104 4284 87120 4318
rect 87676 4284 87692 4318
rect 65818 4156 65852 4172
rect 57058 4121 57118 4122
rect 58068 4121 58128 4122
rect 60116 4121 60176 4122
rect 55777 4087 55793 4121
rect 56349 4087 56365 4121
rect 56795 4087 56811 4121
rect 57367 4087 57383 4121
rect 57813 4087 57829 4121
rect 58385 4087 58401 4121
rect 58831 4087 58847 4121
rect 59403 4087 59419 4121
rect 59849 4087 59865 4121
rect 60421 4087 60437 4121
rect 60867 4087 60883 4121
rect 61439 4087 61455 4121
rect 62628 4088 62644 4122
rect 62768 4088 62784 4122
rect 62926 4088 62942 4122
rect 63066 4088 63082 4122
rect 63224 4088 63240 4122
rect 63364 4088 63380 4122
rect 63522 4088 63538 4122
rect 63662 4088 63678 4122
rect 63820 4088 63836 4122
rect 63960 4088 63976 4122
rect 64118 4088 64134 4122
rect 64258 4088 64274 4122
rect 64416 4088 64432 4122
rect 64556 4088 64572 4122
rect 64714 4088 64730 4122
rect 64854 4088 64870 4122
rect 65012 4088 65028 4122
rect 65152 4088 65168 4122
rect 65310 4088 65326 4122
rect 65450 4088 65466 4122
rect 65608 4088 65624 4122
rect 65748 4088 65764 4122
rect 62976 4068 63036 4088
rect 68030 4050 68112 4074
rect 68030 4016 68054 4050
rect 68088 4016 68112 4050
rect 68030 3992 68112 4016
rect 69048 4050 69130 4074
rect 69048 4016 69072 4050
rect 69106 4016 69130 4050
rect 69048 3992 69130 4016
rect 70066 4050 70148 4074
rect 70066 4016 70090 4050
rect 70124 4016 70148 4050
rect 70066 3992 70148 4016
rect 71084 4050 71166 4074
rect 71084 4016 71108 4050
rect 71142 4016 71166 4050
rect 71084 3992 71166 4016
rect 72102 4050 72184 4074
rect 72102 4016 72126 4050
rect 72160 4016 72184 4050
rect 72102 3992 72184 4016
rect 73120 4050 73202 4074
rect 73120 4016 73144 4050
rect 73178 4016 73202 4050
rect 73120 3992 73202 4016
rect 74138 4050 74220 4074
rect 74138 4016 74162 4050
rect 74196 4016 74220 4050
rect 74138 3992 74220 4016
rect 75156 4050 75238 4074
rect 75156 4016 75180 4050
rect 75214 4016 75238 4050
rect 75156 3992 75238 4016
rect 76174 4050 76256 4074
rect 76174 4016 76198 4050
rect 76232 4016 76256 4050
rect 76174 3992 76256 4016
rect 77192 4050 77274 4074
rect 77192 4016 77216 4050
rect 77250 4016 77274 4050
rect 77192 3992 77274 4016
rect 78210 4050 78292 4074
rect 78210 4016 78234 4050
rect 78268 4016 78292 4050
rect 78210 3992 78292 4016
rect 79228 4050 79310 4074
rect 79228 4016 79252 4050
rect 79286 4016 79310 4050
rect 79228 3992 79310 4016
rect 80246 4050 80328 4074
rect 80246 4016 80270 4050
rect 80304 4016 80328 4050
rect 80246 3992 80328 4016
rect 81264 4050 81346 4074
rect 81264 4016 81288 4050
rect 81322 4016 81346 4050
rect 81264 3992 81346 4016
rect 82282 4050 82364 4074
rect 82282 4016 82306 4050
rect 82340 4016 82364 4050
rect 82282 3992 82364 4016
rect 83300 4050 83382 4074
rect 83300 4016 83324 4050
rect 83358 4016 83382 4050
rect 83300 3992 83382 4016
rect 84318 4050 84400 4074
rect 84318 4016 84342 4050
rect 84376 4016 84400 4050
rect 84318 3992 84400 4016
rect 85336 4050 85418 4074
rect 85336 4016 85360 4050
rect 85394 4016 85418 4050
rect 85336 3992 85418 4016
rect 86354 4050 86436 4074
rect 86354 4016 86378 4050
rect 86412 4016 86436 4050
rect 86354 3992 86436 4016
rect 87372 4050 87454 4074
rect 87372 4016 87396 4050
rect 87430 4016 87454 4050
rect 87372 3992 87454 4016
rect 56052 3940 56134 3964
rect 56052 3906 56076 3940
rect 56110 3906 56134 3940
rect 56052 3882 56134 3906
rect 57070 3940 57152 3964
rect 57070 3906 57094 3940
rect 57128 3906 57152 3940
rect 57070 3882 57152 3906
rect 58088 3940 58170 3964
rect 58088 3906 58112 3940
rect 58146 3906 58170 3940
rect 58088 3882 58170 3906
rect 59106 3940 59188 3964
rect 59106 3906 59130 3940
rect 59164 3906 59188 3940
rect 59106 3882 59188 3906
rect 60124 3940 60206 3964
rect 60124 3906 60148 3940
rect 60182 3906 60206 3940
rect 60124 3882 60206 3906
rect 61142 3940 61224 3964
rect 61142 3906 61166 3940
rect 61200 3906 61224 3940
rect 61142 3882 61224 3906
rect 62590 3928 62672 3952
rect 62590 3894 62614 3928
rect 62648 3894 62672 3928
rect 62590 3870 62672 3894
rect 63608 3928 63690 3952
rect 63608 3894 63632 3928
rect 63666 3894 63690 3928
rect 63608 3870 63690 3894
rect 64626 3928 64708 3952
rect 64626 3894 64650 3928
rect 64684 3894 64708 3928
rect 64626 3870 64708 3894
rect 65644 3928 65726 3952
rect 65644 3894 65668 3928
rect 65702 3894 65726 3928
rect 65644 3870 65726 3894
rect 67762 3760 67778 3794
rect 68334 3760 68350 3794
rect 68780 3760 68796 3794
rect 69352 3760 69368 3794
rect 69798 3760 69814 3794
rect 70370 3760 70386 3794
rect 70816 3760 70832 3794
rect 71388 3760 71404 3794
rect 71834 3760 71850 3794
rect 72406 3760 72422 3794
rect 72852 3760 72868 3794
rect 73424 3760 73440 3794
rect 73870 3760 73886 3794
rect 74442 3760 74458 3794
rect 74888 3760 74904 3794
rect 75460 3760 75476 3794
rect 75906 3760 75922 3794
rect 76478 3760 76494 3794
rect 76924 3760 76940 3794
rect 77496 3760 77512 3794
rect 77942 3760 77958 3794
rect 78514 3760 78530 3794
rect 78960 3760 78976 3794
rect 79532 3760 79548 3794
rect 79978 3760 79994 3794
rect 80550 3760 80566 3794
rect 80996 3760 81012 3794
rect 81568 3760 81584 3794
rect 82014 3760 82030 3794
rect 82586 3760 82602 3794
rect 83032 3760 83048 3794
rect 83604 3760 83620 3794
rect 84050 3760 84066 3794
rect 84622 3760 84638 3794
rect 85068 3760 85084 3794
rect 85640 3760 85656 3794
rect 86086 3760 86102 3794
rect 86658 3760 86674 3794
rect 87104 3760 87120 3794
rect 87676 3760 87692 3794
rect 71070 3758 71130 3760
rect 55776 3684 55792 3718
rect 56348 3684 56364 3718
rect 56794 3684 56810 3718
rect 57366 3684 57382 3718
rect 57812 3684 57828 3718
rect 58384 3684 58400 3718
rect 58830 3684 58846 3718
rect 59402 3684 59418 3718
rect 59848 3684 59864 3718
rect 60420 3684 60436 3718
rect 60866 3684 60882 3718
rect 61438 3684 61454 3718
rect 62628 3686 62644 3720
rect 62768 3686 62784 3720
rect 62926 3686 62942 3720
rect 63066 3686 63082 3720
rect 63224 3686 63240 3720
rect 63364 3686 63380 3720
rect 63522 3686 63538 3720
rect 63662 3686 63678 3720
rect 63820 3686 63836 3720
rect 63960 3686 63976 3720
rect 64118 3686 64134 3720
rect 64258 3686 64274 3720
rect 64416 3686 64432 3720
rect 64556 3686 64572 3720
rect 64714 3686 64730 3720
rect 64854 3686 64870 3720
rect 65012 3686 65028 3720
rect 65152 3686 65168 3720
rect 65310 3686 65326 3720
rect 65450 3686 65466 3720
rect 65608 3686 65624 3720
rect 65748 3686 65764 3720
rect 67530 3710 67564 3726
rect 57058 3682 57118 3684
rect 59094 3682 59154 3684
rect 60116 3682 60176 3684
rect 55544 3634 55578 3650
rect 55544 3042 55578 3058
rect 56562 3634 56596 3650
rect 56562 3042 56596 3058
rect 57580 3634 57614 3650
rect 57580 3042 57614 3058
rect 58598 3634 58632 3650
rect 58598 3042 58632 3058
rect 59616 3634 59650 3650
rect 59616 3042 59650 3058
rect 60634 3634 60668 3650
rect 60634 3042 60668 3058
rect 61652 3634 61686 3650
rect 61652 3042 61686 3058
rect 62540 3636 62574 3652
rect 62540 3044 62574 3060
rect 62838 3636 62872 3652
rect 62838 3044 62872 3060
rect 63136 3636 63170 3652
rect 63136 3044 63170 3060
rect 63434 3636 63468 3652
rect 63434 3044 63468 3060
rect 63732 3636 63766 3652
rect 63732 3044 63766 3060
rect 64030 3636 64064 3652
rect 64030 3044 64064 3060
rect 64328 3636 64362 3652
rect 64328 3044 64362 3060
rect 64626 3636 64660 3652
rect 64626 3044 64660 3060
rect 64924 3636 64958 3652
rect 64924 3044 64958 3060
rect 65222 3636 65256 3652
rect 65222 3044 65256 3060
rect 65520 3636 65554 3652
rect 65520 3044 65554 3060
rect 65818 3636 65852 3652
rect 67530 3118 67564 3134
rect 68548 3710 68582 3726
rect 68548 3118 68582 3134
rect 69566 3710 69600 3726
rect 69566 3118 69600 3134
rect 70584 3710 70618 3726
rect 70584 3118 70618 3134
rect 71602 3710 71636 3726
rect 71602 3118 71636 3134
rect 72620 3710 72654 3726
rect 72620 3118 72654 3134
rect 73638 3710 73672 3726
rect 73638 3118 73672 3134
rect 74656 3710 74690 3726
rect 74656 3118 74690 3134
rect 75674 3710 75708 3726
rect 75674 3118 75708 3134
rect 76692 3710 76726 3726
rect 76692 3118 76726 3134
rect 77710 3710 77744 3726
rect 77710 3118 77744 3134
rect 78728 3710 78762 3726
rect 78728 3118 78762 3134
rect 79746 3710 79780 3726
rect 79746 3118 79780 3134
rect 80764 3710 80798 3726
rect 80764 3118 80798 3134
rect 81782 3710 81816 3726
rect 81782 3118 81816 3134
rect 82800 3710 82834 3726
rect 82800 3118 82834 3134
rect 83818 3710 83852 3726
rect 83818 3118 83852 3134
rect 84836 3710 84870 3726
rect 84836 3118 84870 3134
rect 85854 3710 85888 3726
rect 85854 3118 85888 3134
rect 86872 3710 86906 3726
rect 86872 3118 86906 3134
rect 87890 3710 87924 3726
rect 87890 3118 87924 3134
rect 69038 3084 69098 3086
rect 75150 3084 75210 3086
rect 77184 3084 77244 3086
rect 81250 3084 81310 3090
rect 85326 3084 85386 3086
rect 86342 3084 86402 3086
rect 65818 3044 65852 3060
rect 67762 3050 67778 3084
rect 68334 3050 68350 3084
rect 68780 3050 68796 3084
rect 69352 3050 69368 3084
rect 69798 3050 69814 3084
rect 70370 3050 70386 3084
rect 70816 3050 70832 3084
rect 71388 3050 71404 3084
rect 71834 3050 71850 3084
rect 72406 3050 72422 3084
rect 72852 3050 72868 3084
rect 73424 3050 73440 3084
rect 73870 3050 73886 3084
rect 74442 3050 74458 3084
rect 74888 3050 74904 3084
rect 75460 3050 75476 3084
rect 75906 3050 75922 3084
rect 76478 3050 76494 3084
rect 76924 3050 76940 3084
rect 77496 3050 77512 3084
rect 77942 3050 77958 3084
rect 78514 3050 78530 3084
rect 78960 3050 78976 3084
rect 79532 3050 79548 3084
rect 79978 3050 79994 3084
rect 80550 3050 80566 3084
rect 80996 3050 81012 3084
rect 81568 3050 81584 3084
rect 82014 3050 82030 3084
rect 82586 3050 82602 3084
rect 83032 3050 83048 3084
rect 83604 3050 83620 3084
rect 84050 3050 84066 3084
rect 84622 3050 84638 3084
rect 85068 3050 85084 3084
rect 85640 3050 85656 3084
rect 86086 3050 86102 3084
rect 86658 3050 86674 3084
rect 87104 3050 87120 3084
rect 87676 3050 87692 3084
rect 57060 3008 57120 3012
rect 58070 3008 58130 3012
rect 60118 3008 60178 3012
rect 55776 2974 55792 3008
rect 56348 2974 56364 3008
rect 56794 2974 56810 3008
rect 57366 2974 57382 3008
rect 57812 2974 57828 3008
rect 58384 2974 58400 3008
rect 58830 2974 58846 3008
rect 59402 2974 59418 3008
rect 59848 2974 59864 3008
rect 60420 2974 60436 3008
rect 60866 2974 60882 3008
rect 61438 2974 61454 3008
rect 62628 2976 62644 3010
rect 62768 2976 62784 3010
rect 62926 2976 62942 3010
rect 63066 2976 63082 3010
rect 63224 2976 63240 3010
rect 63364 2976 63380 3010
rect 63522 2976 63538 3010
rect 63662 2976 63678 3010
rect 63820 2976 63836 3010
rect 63960 2976 63976 3010
rect 64118 2976 64134 3010
rect 64258 2976 64274 3010
rect 64416 2976 64432 3010
rect 64556 2976 64572 3010
rect 64714 2976 64730 3010
rect 64854 2976 64870 3010
rect 65012 2976 65028 3010
rect 65152 2976 65168 3010
rect 65310 2976 65326 3010
rect 65450 2976 65466 3010
rect 65608 2976 65624 3010
rect 65748 2976 65764 3010
rect 56026 2814 56108 2838
rect 56026 2780 56050 2814
rect 56084 2780 56108 2814
rect 56026 2756 56108 2780
rect 57044 2814 57126 2838
rect 57044 2780 57068 2814
rect 57102 2780 57126 2814
rect 57044 2756 57126 2780
rect 58062 2814 58144 2838
rect 58062 2780 58086 2814
rect 58120 2780 58144 2814
rect 58062 2756 58144 2780
rect 59080 2814 59162 2838
rect 59080 2780 59104 2814
rect 59138 2780 59162 2814
rect 59080 2756 59162 2780
rect 60098 2814 60180 2838
rect 60098 2780 60122 2814
rect 60156 2780 60180 2814
rect 60098 2756 60180 2780
rect 61116 2814 61198 2838
rect 61116 2780 61140 2814
rect 61174 2780 61198 2814
rect 61116 2756 61198 2780
rect 62590 2814 62672 2838
rect 62590 2780 62614 2814
rect 62648 2780 62672 2814
rect 62590 2756 62672 2780
rect 63608 2814 63690 2838
rect 63608 2780 63632 2814
rect 63666 2780 63690 2814
rect 63608 2756 63690 2780
rect 64626 2814 64708 2838
rect 64626 2780 64650 2814
rect 64684 2780 64708 2814
rect 64626 2756 64708 2780
rect 65644 2814 65726 2838
rect 65644 2780 65668 2814
rect 65702 2780 65726 2814
rect 65644 2756 65726 2780
rect 68016 2828 68098 2852
rect 68016 2794 68040 2828
rect 68074 2794 68098 2828
rect 68016 2770 68098 2794
rect 69034 2828 69116 2852
rect 69034 2794 69058 2828
rect 69092 2794 69116 2828
rect 69034 2770 69116 2794
rect 70052 2828 70134 2852
rect 70052 2794 70076 2828
rect 70110 2794 70134 2828
rect 70052 2770 70134 2794
rect 71070 2828 71152 2852
rect 71070 2794 71094 2828
rect 71128 2794 71152 2828
rect 71070 2770 71152 2794
rect 72088 2828 72170 2852
rect 72088 2794 72112 2828
rect 72146 2794 72170 2828
rect 72088 2770 72170 2794
rect 73106 2828 73188 2852
rect 73106 2794 73130 2828
rect 73164 2794 73188 2828
rect 73106 2770 73188 2794
rect 74124 2828 74206 2852
rect 74124 2794 74148 2828
rect 74182 2794 74206 2828
rect 74124 2770 74206 2794
rect 75142 2828 75224 2852
rect 75142 2794 75166 2828
rect 75200 2794 75224 2828
rect 75142 2770 75224 2794
rect 76160 2828 76242 2852
rect 76160 2794 76184 2828
rect 76218 2794 76242 2828
rect 76160 2770 76242 2794
rect 77178 2828 77260 2852
rect 77178 2794 77202 2828
rect 77236 2794 77260 2828
rect 77178 2770 77260 2794
rect 78196 2828 78278 2852
rect 78196 2794 78220 2828
rect 78254 2794 78278 2828
rect 78196 2770 78278 2794
rect 79214 2828 79296 2852
rect 79214 2794 79238 2828
rect 79272 2794 79296 2828
rect 79214 2770 79296 2794
rect 80232 2828 80314 2852
rect 80232 2794 80256 2828
rect 80290 2794 80314 2828
rect 80232 2770 80314 2794
rect 81250 2828 81332 2852
rect 81250 2794 81274 2828
rect 81308 2794 81332 2828
rect 81250 2770 81332 2794
rect 82268 2828 82350 2852
rect 82268 2794 82292 2828
rect 82326 2794 82350 2828
rect 82268 2770 82350 2794
rect 83286 2828 83368 2852
rect 83286 2794 83310 2828
rect 83344 2794 83368 2828
rect 83286 2770 83368 2794
rect 84304 2828 84386 2852
rect 84304 2794 84328 2828
rect 84362 2794 84386 2828
rect 84304 2770 84386 2794
rect 85322 2828 85404 2852
rect 85322 2794 85346 2828
rect 85380 2794 85404 2828
rect 85322 2770 85404 2794
rect 86340 2828 86422 2852
rect 86340 2794 86364 2828
rect 86398 2794 86422 2828
rect 86340 2770 86422 2794
rect 87358 2828 87440 2852
rect 87358 2794 87382 2828
rect 87416 2794 87440 2828
rect 87358 2770 87440 2794
rect 55777 2573 55793 2607
rect 56349 2573 56365 2607
rect 56795 2573 56811 2607
rect 57367 2573 57383 2607
rect 57813 2573 57829 2607
rect 58385 2573 58401 2607
rect 58831 2573 58847 2607
rect 59403 2573 59419 2607
rect 59849 2573 59865 2607
rect 60421 2573 60437 2607
rect 60867 2573 60883 2607
rect 61439 2573 61455 2607
rect 62626 2574 62642 2608
rect 62766 2574 62782 2608
rect 62924 2574 62940 2608
rect 63064 2574 63080 2608
rect 63222 2574 63238 2608
rect 63362 2574 63378 2608
rect 63520 2574 63536 2608
rect 63660 2574 63676 2608
rect 63818 2574 63834 2608
rect 63958 2574 63974 2608
rect 64116 2574 64132 2608
rect 64256 2574 64272 2608
rect 64414 2574 64430 2608
rect 64554 2574 64570 2608
rect 64712 2574 64728 2608
rect 64852 2574 64868 2608
rect 65010 2574 65026 2608
rect 65150 2574 65166 2608
rect 65308 2574 65324 2608
rect 65448 2574 65464 2608
rect 65606 2574 65622 2608
rect 65746 2574 65762 2608
rect 57060 2572 57120 2573
rect 59096 2572 59156 2573
rect 60118 2572 60178 2573
rect 55545 2523 55579 2539
rect 55545 1931 55579 1947
rect 56563 2523 56597 2539
rect 56563 1931 56597 1947
rect 57581 2523 57615 2539
rect 57581 1931 57615 1947
rect 58599 2523 58633 2539
rect 58599 1931 58633 1947
rect 59617 2523 59651 2539
rect 59617 1931 59651 1947
rect 60635 2523 60669 2539
rect 60635 1931 60669 1947
rect 61653 2523 61687 2539
rect 61653 1931 61687 1947
rect 62538 2524 62572 2540
rect 62538 1932 62572 1948
rect 62836 2524 62870 2540
rect 62836 1932 62870 1948
rect 63134 2524 63168 2540
rect 63134 1932 63168 1948
rect 63432 2524 63466 2540
rect 63432 1932 63466 1948
rect 63730 2524 63764 2540
rect 63730 1932 63764 1948
rect 64028 2524 64062 2540
rect 64028 1932 64062 1948
rect 64326 2524 64360 2540
rect 64326 1932 64360 1948
rect 64624 2524 64658 2540
rect 64624 1932 64658 1948
rect 64922 2524 64956 2540
rect 64922 1932 64956 1948
rect 65220 2524 65254 2540
rect 65220 1932 65254 1948
rect 65518 2524 65552 2540
rect 65518 1932 65552 1948
rect 65816 2524 65850 2540
rect 67762 2526 67778 2560
rect 68334 2526 68350 2560
rect 68780 2526 68796 2560
rect 69352 2526 69368 2560
rect 69798 2526 69814 2560
rect 70370 2526 70386 2560
rect 70816 2526 70832 2560
rect 71388 2526 71404 2560
rect 71834 2526 71850 2560
rect 72406 2526 72422 2560
rect 72852 2526 72868 2560
rect 73424 2526 73440 2560
rect 73870 2526 73886 2560
rect 74442 2526 74458 2560
rect 74888 2526 74904 2560
rect 75460 2526 75476 2560
rect 75906 2526 75922 2560
rect 76478 2526 76494 2560
rect 76924 2526 76940 2560
rect 77496 2526 77512 2560
rect 77942 2526 77958 2560
rect 78514 2526 78530 2560
rect 78960 2526 78976 2560
rect 79532 2526 79548 2560
rect 79978 2526 79994 2560
rect 80550 2526 80566 2560
rect 80996 2526 81012 2560
rect 81568 2526 81584 2560
rect 82014 2526 82030 2560
rect 82586 2526 82602 2560
rect 83032 2526 83048 2560
rect 83604 2526 83620 2560
rect 84050 2526 84066 2560
rect 84622 2526 84638 2560
rect 85068 2526 85084 2560
rect 85640 2526 85656 2560
rect 86086 2526 86102 2560
rect 86658 2526 86674 2560
rect 87104 2526 87120 2560
rect 87676 2526 87692 2560
rect 74148 2520 74208 2526
rect 79220 2520 79280 2526
rect 80240 2520 80300 2526
rect 82276 2520 82336 2526
rect 65816 1932 65850 1948
rect 67530 2476 67564 2492
rect 57062 1897 57122 1902
rect 58072 1897 58132 1902
rect 59098 1897 59158 1898
rect 60120 1897 60180 1902
rect 55777 1863 55793 1897
rect 56349 1863 56365 1897
rect 56795 1863 56811 1897
rect 57367 1863 57383 1897
rect 57813 1863 57829 1897
rect 58385 1863 58401 1897
rect 58831 1863 58847 1897
rect 59403 1863 59419 1897
rect 59849 1863 59865 1897
rect 60421 1863 60437 1897
rect 60867 1863 60883 1897
rect 61439 1863 61455 1897
rect 62626 1864 62642 1898
rect 62766 1864 62782 1898
rect 62924 1864 62940 1898
rect 63064 1864 63080 1898
rect 63222 1864 63238 1898
rect 63362 1864 63378 1898
rect 63520 1864 63536 1898
rect 63660 1864 63676 1898
rect 63818 1864 63834 1898
rect 63958 1864 63974 1898
rect 64116 1864 64132 1898
rect 64256 1864 64272 1898
rect 64414 1864 64430 1898
rect 64554 1864 64570 1898
rect 64712 1864 64728 1898
rect 64852 1864 64868 1898
rect 65010 1864 65026 1898
rect 65150 1864 65166 1898
rect 65308 1864 65324 1898
rect 65448 1864 65464 1898
rect 65606 1864 65622 1898
rect 65746 1864 65762 1898
rect 67530 1884 67564 1900
rect 68548 2476 68582 2492
rect 68548 1884 68582 1900
rect 69566 2476 69600 2492
rect 69566 1884 69600 1900
rect 70584 2476 70618 2492
rect 70584 1884 70618 1900
rect 71602 2476 71636 2492
rect 71602 1884 71636 1900
rect 72620 2476 72654 2492
rect 72620 1884 72654 1900
rect 73638 2476 73672 2492
rect 73638 1884 73672 1900
rect 74656 2476 74690 2492
rect 74656 1884 74690 1900
rect 75674 2476 75708 2492
rect 75674 1884 75708 1900
rect 76692 2476 76726 2492
rect 76692 1884 76726 1900
rect 77710 2476 77744 2492
rect 77710 1884 77744 1900
rect 78728 2476 78762 2492
rect 78728 1884 78762 1900
rect 79746 2476 79780 2492
rect 79746 1884 79780 1900
rect 80764 2476 80798 2492
rect 80764 1884 80798 1900
rect 81782 2476 81816 2492
rect 81782 1884 81816 1900
rect 82800 2476 82834 2492
rect 82800 1884 82834 1900
rect 83818 2476 83852 2492
rect 83818 1884 83852 1900
rect 84836 2476 84870 2492
rect 84836 1884 84870 1900
rect 85854 2476 85888 2492
rect 85854 1884 85888 1900
rect 86872 2476 86906 2492
rect 86872 1884 86906 1900
rect 87890 2476 87924 2492
rect 87890 1884 87924 1900
rect 78204 1850 78264 1856
rect 67762 1816 67778 1850
rect 68334 1816 68350 1850
rect 68780 1816 68796 1850
rect 69352 1816 69368 1850
rect 69798 1816 69814 1850
rect 70370 1816 70386 1850
rect 70816 1816 70832 1850
rect 71388 1816 71404 1850
rect 71834 1816 71850 1850
rect 72406 1816 72422 1850
rect 72852 1816 72868 1850
rect 73424 1816 73440 1850
rect 73870 1816 73886 1850
rect 74442 1816 74458 1850
rect 74888 1816 74904 1850
rect 75460 1816 75476 1850
rect 75906 1816 75922 1850
rect 76478 1816 76494 1850
rect 76924 1816 76940 1850
rect 77496 1816 77512 1850
rect 77942 1816 77958 1850
rect 78514 1816 78530 1850
rect 78960 1816 78976 1850
rect 79532 1816 79548 1850
rect 79978 1816 79994 1850
rect 80550 1816 80566 1850
rect 80996 1816 81012 1850
rect 81568 1816 81584 1850
rect 82014 1816 82030 1850
rect 82586 1816 82602 1850
rect 83032 1816 83048 1850
rect 83604 1816 83620 1850
rect 84050 1816 84066 1850
rect 84622 1816 84638 1850
rect 85068 1816 85084 1850
rect 85640 1816 85656 1850
rect 86086 1816 86102 1850
rect 86658 1816 86674 1850
rect 87104 1816 87120 1850
rect 87676 1816 87692 1850
rect 56052 1716 56134 1740
rect 56052 1682 56076 1716
rect 56110 1682 56134 1716
rect 56052 1658 56134 1682
rect 57070 1716 57152 1740
rect 57070 1682 57094 1716
rect 57128 1682 57152 1716
rect 57070 1658 57152 1682
rect 58088 1716 58170 1740
rect 58088 1682 58112 1716
rect 58146 1682 58170 1716
rect 58088 1658 58170 1682
rect 59106 1716 59188 1740
rect 59106 1682 59130 1716
rect 59164 1682 59188 1716
rect 59106 1658 59188 1682
rect 60124 1716 60206 1740
rect 60124 1682 60148 1716
rect 60182 1682 60206 1716
rect 60124 1658 60206 1682
rect 61142 1716 61224 1740
rect 61142 1682 61166 1716
rect 61200 1682 61224 1716
rect 61142 1658 61224 1682
rect 62644 1702 62726 1726
rect 62644 1668 62668 1702
rect 62702 1668 62726 1702
rect 62644 1644 62726 1668
rect 63662 1702 63744 1726
rect 63662 1668 63686 1702
rect 63720 1668 63744 1702
rect 63662 1644 63744 1668
rect 64680 1702 64762 1726
rect 64680 1668 64704 1702
rect 64738 1668 64762 1702
rect 64680 1644 64762 1668
rect 65698 1702 65780 1726
rect 65698 1668 65722 1702
rect 65756 1668 65780 1702
rect 65698 1644 65780 1668
rect 68016 1608 68098 1632
rect 68016 1574 68040 1608
rect 68074 1574 68098 1608
rect 68016 1550 68098 1574
rect 69034 1608 69116 1632
rect 69034 1574 69058 1608
rect 69092 1574 69116 1608
rect 69034 1550 69116 1574
rect 70052 1608 70134 1632
rect 70052 1574 70076 1608
rect 70110 1574 70134 1608
rect 70052 1550 70134 1574
rect 71070 1608 71152 1632
rect 71070 1574 71094 1608
rect 71128 1574 71152 1608
rect 71070 1550 71152 1574
rect 72088 1608 72170 1632
rect 72088 1574 72112 1608
rect 72146 1574 72170 1608
rect 72088 1550 72170 1574
rect 73106 1608 73188 1632
rect 73106 1574 73130 1608
rect 73164 1574 73188 1608
rect 73106 1550 73188 1574
rect 74124 1608 74206 1632
rect 74124 1574 74148 1608
rect 74182 1574 74206 1608
rect 74124 1550 74206 1574
rect 75142 1608 75224 1632
rect 75142 1574 75166 1608
rect 75200 1574 75224 1608
rect 75142 1550 75224 1574
rect 76160 1608 76242 1632
rect 76160 1574 76184 1608
rect 76218 1574 76242 1608
rect 76160 1550 76242 1574
rect 77178 1608 77260 1632
rect 77178 1574 77202 1608
rect 77236 1574 77260 1608
rect 77178 1550 77260 1574
rect 78196 1608 78278 1632
rect 78196 1574 78220 1608
rect 78254 1574 78278 1608
rect 78196 1550 78278 1574
rect 79214 1608 79296 1632
rect 79214 1574 79238 1608
rect 79272 1574 79296 1608
rect 79214 1550 79296 1574
rect 80232 1608 80314 1632
rect 80232 1574 80256 1608
rect 80290 1574 80314 1608
rect 80232 1550 80314 1574
rect 81250 1608 81332 1632
rect 81250 1574 81274 1608
rect 81308 1574 81332 1608
rect 81250 1550 81332 1574
rect 82268 1608 82350 1632
rect 82268 1574 82292 1608
rect 82326 1574 82350 1608
rect 82268 1550 82350 1574
rect 83286 1608 83368 1632
rect 83286 1574 83310 1608
rect 83344 1574 83368 1608
rect 83286 1550 83368 1574
rect 84304 1608 84386 1632
rect 84304 1574 84328 1608
rect 84362 1574 84386 1608
rect 84304 1550 84386 1574
rect 85322 1608 85404 1632
rect 85322 1574 85346 1608
rect 85380 1574 85404 1608
rect 85322 1550 85404 1574
rect 86340 1608 86422 1632
rect 86340 1574 86364 1608
rect 86398 1574 86422 1608
rect 86340 1550 86422 1574
rect 87358 1608 87440 1632
rect 87358 1574 87382 1608
rect 87416 1574 87440 1608
rect 87358 1550 87440 1574
rect 55776 1460 55792 1494
rect 56348 1460 56364 1494
rect 56794 1460 56810 1494
rect 57366 1460 57382 1494
rect 57812 1460 57828 1494
rect 58384 1460 58400 1494
rect 58830 1460 58846 1494
rect 59402 1460 59418 1494
rect 59848 1460 59864 1494
rect 60420 1460 60436 1494
rect 60866 1460 60882 1494
rect 61438 1460 61454 1494
rect 62626 1464 62642 1498
rect 62766 1464 62782 1498
rect 62924 1464 62940 1498
rect 63064 1464 63080 1498
rect 63222 1464 63238 1498
rect 63362 1464 63378 1498
rect 63520 1464 63536 1498
rect 63660 1464 63676 1498
rect 63818 1464 63834 1498
rect 63958 1464 63974 1498
rect 64116 1464 64132 1498
rect 64256 1464 64272 1498
rect 64414 1464 64430 1498
rect 64554 1464 64570 1498
rect 64712 1464 64728 1498
rect 64852 1464 64868 1498
rect 65010 1464 65026 1498
rect 65150 1464 65166 1498
rect 65308 1464 65324 1498
rect 65448 1464 65464 1498
rect 65606 1464 65622 1498
rect 65746 1464 65762 1498
rect 55544 1410 55578 1426
rect 55544 818 55578 834
rect 56562 1410 56596 1426
rect 56562 818 56596 834
rect 57580 1410 57614 1426
rect 57580 818 57614 834
rect 58598 1410 58632 1426
rect 58598 818 58632 834
rect 59616 1410 59650 1426
rect 59616 818 59650 834
rect 60634 1410 60668 1426
rect 60634 818 60668 834
rect 61652 1410 61686 1426
rect 61652 818 61686 834
rect 62538 1414 62572 1430
rect 62538 822 62572 838
rect 62836 1414 62870 1430
rect 62836 822 62870 838
rect 63134 1414 63168 1430
rect 63134 822 63168 838
rect 63432 1414 63466 1430
rect 63432 822 63466 838
rect 63730 1414 63764 1430
rect 63730 822 63764 838
rect 64028 1414 64062 1430
rect 64028 822 64062 838
rect 64326 1414 64360 1430
rect 64326 822 64360 838
rect 64624 1414 64658 1430
rect 64624 822 64658 838
rect 64922 1414 64956 1430
rect 64922 822 64956 838
rect 65220 1414 65254 1430
rect 65220 822 65254 838
rect 65518 1414 65552 1430
rect 65518 822 65552 838
rect 65816 1414 65850 1430
rect 67762 1294 67778 1328
rect 68334 1294 68350 1328
rect 68780 1294 68796 1328
rect 69352 1294 69368 1328
rect 69798 1294 69814 1328
rect 70370 1294 70386 1328
rect 70816 1294 70832 1328
rect 71388 1294 71404 1328
rect 71834 1294 71850 1328
rect 72406 1294 72422 1328
rect 72852 1294 72868 1328
rect 73424 1294 73440 1328
rect 73870 1294 73886 1328
rect 74442 1294 74458 1328
rect 74888 1294 74904 1328
rect 75460 1294 75476 1328
rect 75906 1294 75922 1328
rect 76478 1294 76494 1328
rect 76924 1294 76940 1328
rect 77496 1294 77512 1328
rect 77942 1294 77958 1328
rect 78514 1294 78530 1328
rect 78960 1294 78976 1328
rect 79532 1294 79548 1328
rect 79978 1294 79994 1328
rect 80550 1294 80566 1328
rect 80996 1294 81012 1328
rect 81568 1294 81584 1328
rect 82014 1294 82030 1328
rect 82586 1294 82602 1328
rect 83032 1294 83048 1328
rect 83604 1294 83620 1328
rect 84050 1294 84066 1328
rect 84622 1294 84638 1328
rect 85068 1294 85084 1328
rect 85640 1294 85656 1328
rect 86086 1294 86102 1328
rect 86658 1294 86674 1328
rect 87104 1294 87120 1328
rect 87676 1294 87692 1328
rect 68016 1290 68076 1294
rect 69038 1290 69098 1294
rect 70064 1290 70124 1294
rect 71080 1290 71140 1294
rect 72094 1290 72154 1294
rect 73124 1284 73184 1294
rect 74140 1284 74200 1294
rect 75144 1290 75204 1294
rect 76174 1284 76234 1294
rect 77194 1290 77254 1294
rect 78204 1290 78264 1294
rect 79228 1284 79288 1294
rect 81254 1290 81314 1294
rect 82274 1284 82334 1294
rect 83298 1290 83358 1294
rect 86342 1290 86402 1294
rect 87364 1292 87424 1294
rect 65816 822 65850 838
rect 67530 1244 67564 1260
rect 55776 750 55792 784
rect 56348 750 56364 784
rect 56794 750 56810 784
rect 57366 750 57382 784
rect 57812 750 57828 784
rect 58384 750 58400 784
rect 58830 750 58846 784
rect 59402 750 59418 784
rect 59848 750 59864 784
rect 60420 750 60436 784
rect 60866 750 60882 784
rect 61438 750 61454 784
rect 62626 754 62642 788
rect 62766 754 62782 788
rect 62924 754 62940 788
rect 63064 754 63080 788
rect 63222 754 63238 788
rect 63362 754 63378 788
rect 63520 754 63536 788
rect 63660 754 63676 788
rect 63818 754 63834 788
rect 63958 754 63974 788
rect 64116 754 64132 788
rect 64256 754 64272 788
rect 64414 754 64430 788
rect 64554 754 64570 788
rect 64712 754 64728 788
rect 64852 754 64868 788
rect 65010 754 65026 788
rect 65150 754 65166 788
rect 65308 754 65324 788
rect 65448 754 65464 788
rect 65606 754 65622 788
rect 65746 754 65762 788
rect 68548 1244 68582 1260
rect 68532 668 68548 708
rect 69566 1244 69600 1260
rect 68582 668 68592 708
rect 67530 652 67564 668
rect 68548 652 68582 668
rect 69566 652 69600 668
rect 70584 1244 70618 1260
rect 70584 652 70618 668
rect 71602 1244 71636 1260
rect 72620 1244 72654 1260
rect 72606 668 72620 712
rect 73638 1244 73672 1260
rect 72654 668 72666 712
rect 71602 652 71636 668
rect 72620 652 72654 668
rect 73638 652 73672 668
rect 74656 1244 74690 1260
rect 74656 652 74690 668
rect 75674 1244 75708 1260
rect 75674 652 75708 668
rect 76692 1244 76726 1260
rect 76692 652 76726 668
rect 77710 1244 77744 1260
rect 78728 1244 78762 1260
rect 78714 668 78728 714
rect 79746 1244 79780 1260
rect 78762 668 78774 714
rect 77710 652 77744 668
rect 78728 652 78762 668
rect 79746 652 79780 668
rect 80764 1244 80798 1260
rect 80764 652 80798 668
rect 81782 1244 81816 1260
rect 82800 1244 82834 1260
rect 82786 668 82800 704
rect 83818 1244 83852 1260
rect 82834 668 82846 704
rect 81782 652 81816 668
rect 82800 652 82834 668
rect 83818 652 83852 668
rect 84836 1244 84870 1260
rect 84836 652 84870 668
rect 85854 1244 85888 1260
rect 86872 1244 86906 1260
rect 86856 668 86872 706
rect 87890 1244 87924 1260
rect 86906 668 86916 706
rect 85854 652 85888 668
rect 86872 652 86906 668
rect 87890 652 87924 668
rect 74136 618 74196 620
rect 80248 618 80308 620
rect 85334 618 85394 620
rect 67762 584 67778 618
rect 68334 584 68350 618
rect 68780 584 68796 618
rect 69352 584 69368 618
rect 69798 584 69814 618
rect 70370 584 70386 618
rect 70816 584 70832 618
rect 71388 584 71404 618
rect 71834 584 71850 618
rect 72406 584 72422 618
rect 72852 584 72868 618
rect 73424 584 73440 618
rect 73870 584 73886 618
rect 74442 584 74458 618
rect 74888 584 74904 618
rect 75460 584 75476 618
rect 75906 584 75922 618
rect 76478 584 76494 618
rect 76924 584 76940 618
rect 77496 584 77512 618
rect 77942 584 77958 618
rect 78514 584 78530 618
rect 78960 584 78976 618
rect 79532 584 79548 618
rect 79978 584 79994 618
rect 80550 584 80566 618
rect 80996 584 81012 618
rect 81568 584 81584 618
rect 82014 584 82030 618
rect 82586 584 82602 618
rect 83032 584 83048 618
rect 83604 584 83620 618
rect 84050 584 84066 618
rect 84622 584 84638 618
rect 85068 584 85084 618
rect 85640 584 85656 618
rect 86086 584 86102 618
rect 86658 584 86674 618
rect 87104 584 87120 618
rect 87676 584 87692 618
rect 56026 522 56108 546
rect 56026 488 56050 522
rect 56084 488 56108 522
rect 56026 464 56108 488
rect 57044 522 57126 546
rect 57044 488 57068 522
rect 57102 488 57126 522
rect 57044 464 57126 488
rect 58062 522 58144 546
rect 58062 488 58086 522
rect 58120 488 58144 522
rect 58062 464 58144 488
rect 59080 522 59162 546
rect 59080 488 59104 522
rect 59138 488 59162 522
rect 59080 464 59162 488
rect 60098 522 60180 546
rect 60098 488 60122 522
rect 60156 488 60180 522
rect 60098 464 60180 488
rect 61116 522 61198 546
rect 61116 488 61140 522
rect 61174 488 61198 522
rect 61116 464 61198 488
rect 62618 468 62700 492
rect 62618 434 62642 468
rect 62676 434 62700 468
rect 62618 410 62700 434
rect 63636 468 63718 492
rect 63636 434 63660 468
rect 63694 434 63718 468
rect 63636 410 63718 434
rect 64654 468 64736 492
rect 64654 434 64678 468
rect 64712 434 64736 468
rect 64654 410 64736 434
rect 65672 468 65754 492
rect 65672 434 65696 468
rect 65730 434 65754 468
rect 65672 410 65754 434
rect 52628 -682 52728 -520
rect 89772 -682 89872 -520
<< viali >>
rect 11428 28162 11490 28262
rect 11490 28162 35610 28262
rect 35610 28162 35672 28262
rect 11328 18278 11428 27642
rect 17732 27027 18196 27061
rect 18750 27027 19214 27061
rect 19768 27027 20232 27061
rect 20786 27027 21250 27061
rect 21804 27027 22268 27061
rect 22822 27027 23286 27061
rect 23840 27027 24304 27061
rect 24858 27027 25322 27061
rect 25876 27027 26340 27061
rect 26894 27027 27358 27061
rect 27912 27027 28376 27061
rect 28930 27027 29394 27061
rect 29948 27027 30412 27061
rect 30966 27027 31430 27061
rect 31984 27027 32448 27061
rect 33002 27027 33466 27061
rect 17438 26392 17472 26968
rect 18456 26392 18490 26968
rect 19474 26392 19508 26968
rect 20492 26392 20526 26968
rect 21510 26392 21544 26968
rect 22528 26392 22562 26968
rect 23546 26392 23580 26968
rect 24564 26392 24598 26968
rect 25582 26392 25616 26968
rect 26600 26392 26634 26968
rect 27618 26392 27652 26968
rect 28636 26392 28670 26968
rect 29654 26392 29688 26968
rect 30672 26392 30706 26968
rect 31690 26392 31724 26968
rect 32708 26392 32742 26968
rect 33726 26392 33760 26968
rect 17732 26299 18196 26333
rect 18750 26299 19214 26333
rect 19768 26299 20232 26333
rect 20786 26299 21250 26333
rect 21804 26299 22268 26333
rect 22822 26299 23286 26333
rect 23840 26299 24304 26333
rect 24858 26299 25322 26333
rect 25876 26299 26340 26333
rect 26894 26299 27358 26333
rect 27912 26299 28376 26333
rect 28930 26299 29394 26333
rect 29948 26299 30412 26333
rect 30966 26299 31430 26333
rect 31984 26299 32448 26333
rect 33002 26299 33466 26333
rect 17732 25891 18196 25925
rect 18750 25891 19214 25925
rect 19768 25891 20232 25925
rect 20786 25891 21250 25925
rect 21804 25891 22268 25925
rect 22822 25891 23286 25925
rect 23840 25891 24304 25925
rect 24858 25891 25322 25925
rect 25876 25891 26340 25925
rect 26894 25891 27358 25925
rect 27912 25891 28376 25925
rect 28930 25891 29394 25925
rect 29948 25891 30412 25925
rect 30966 25891 31430 25925
rect 31984 25891 32448 25925
rect 33002 25891 33466 25925
rect 17438 25256 17472 25832
rect 18456 25256 18490 25832
rect 19474 25256 19508 25832
rect 20492 25256 20526 25832
rect 21510 25256 21544 25832
rect 22528 25256 22562 25832
rect 23546 25256 23580 25832
rect 24564 25256 24598 25832
rect 25582 25256 25616 25832
rect 26600 25256 26634 25832
rect 27618 25256 27652 25832
rect 28636 25256 28670 25832
rect 29654 25256 29688 25832
rect 30672 25256 30706 25832
rect 31690 25256 31724 25832
rect 32708 25256 32742 25832
rect 33726 25256 33760 25832
rect 17732 25163 18196 25197
rect 18750 25163 19214 25197
rect 19768 25163 20232 25197
rect 20786 25163 21250 25197
rect 21804 25163 22268 25197
rect 22822 25163 23286 25197
rect 23840 25163 24304 25197
rect 24858 25163 25322 25197
rect 25876 25163 26340 25197
rect 26894 25163 27358 25197
rect 27912 25163 28376 25197
rect 28930 25163 29394 25197
rect 29948 25163 30412 25197
rect 30966 25163 31430 25197
rect 31984 25163 32448 25197
rect 33002 25163 33466 25197
rect 17732 24755 18196 24789
rect 18750 24755 19214 24789
rect 19768 24755 20232 24789
rect 20786 24755 21250 24789
rect 21804 24755 22268 24789
rect 22822 24755 23286 24789
rect 23840 24755 24304 24789
rect 24858 24755 25322 24789
rect 25876 24755 26340 24789
rect 26894 24755 27358 24789
rect 27912 24755 28376 24789
rect 28930 24755 29394 24789
rect 29948 24755 30412 24789
rect 30966 24755 31430 24789
rect 31984 24755 32448 24789
rect 33002 24755 33466 24789
rect 17438 24120 17472 24696
rect 18456 24120 18490 24696
rect 19474 24120 19508 24696
rect 20492 24120 20526 24696
rect 21510 24120 21544 24696
rect 22528 24120 22562 24696
rect 23546 24120 23580 24696
rect 24564 24120 24598 24696
rect 25582 24120 25616 24696
rect 26600 24120 26634 24696
rect 27618 24120 27652 24696
rect 28636 24120 28670 24696
rect 29654 24120 29688 24696
rect 30672 24120 30706 24696
rect 31690 24120 31724 24696
rect 32708 24120 32742 24696
rect 33726 24120 33760 24696
rect 17732 24027 18196 24061
rect 18750 24027 19214 24061
rect 19768 24027 20232 24061
rect 20786 24027 21250 24061
rect 21804 24027 22268 24061
rect 22822 24027 23286 24061
rect 23840 24027 24304 24061
rect 24858 24027 25322 24061
rect 25876 24027 26340 24061
rect 26894 24027 27358 24061
rect 27912 24027 28376 24061
rect 28930 24027 29394 24061
rect 29948 24027 30412 24061
rect 30966 24027 31430 24061
rect 31984 24027 32448 24061
rect 33002 24027 33466 24061
rect 18718 22981 19182 23015
rect 19736 22981 20200 23015
rect 20754 22981 21218 23015
rect 21772 22981 22236 23015
rect 22790 22981 23254 23015
rect 23808 22981 24272 23015
rect 24826 22981 25290 23015
rect 25844 22981 26308 23015
rect 26862 22981 27326 23015
rect 27880 22981 28344 23015
rect 28898 22981 29362 23015
rect 29916 22981 30380 23015
rect 30934 22981 31398 23015
rect 31952 22981 32416 23015
rect 32970 22981 33434 23015
rect 18424 22346 18458 22922
rect 19442 22346 19476 22922
rect 20460 22346 20494 22922
rect 21478 22346 21512 22922
rect 22496 22346 22530 22922
rect 23514 22346 23548 22922
rect 24532 22346 24566 22922
rect 25550 22346 25584 22922
rect 26568 22346 26602 22922
rect 27586 22346 27620 22922
rect 28604 22346 28638 22922
rect 29622 22346 29656 22922
rect 30640 22346 30674 22922
rect 31658 22346 31692 22922
rect 32676 22346 32710 22922
rect 33694 22346 33728 22922
rect 18718 22253 19182 22287
rect 19736 22253 20200 22287
rect 20754 22253 21218 22287
rect 21772 22253 22236 22287
rect 22790 22253 23254 22287
rect 23808 22253 24272 22287
rect 24826 22253 25290 22287
rect 25844 22253 26308 22287
rect 26862 22253 27326 22287
rect 27880 22253 28344 22287
rect 28898 22253 29362 22287
rect 29916 22253 30380 22287
rect 30934 22253 31398 22287
rect 31952 22253 32416 22287
rect 32970 22253 33434 22287
rect 14670 21897 14734 21931
rect 14888 21897 14952 21931
rect 15106 21897 15170 21931
rect 15324 21897 15388 21931
rect 15542 21897 15606 21931
rect 15760 21897 15824 21931
rect 15978 21897 16042 21931
rect 16196 21897 16260 21931
rect 16414 21897 16478 21931
rect 16632 21897 16696 21931
rect 14576 21462 14610 21838
rect 14794 21462 14828 21838
rect 15012 21462 15046 21838
rect 15230 21462 15264 21838
rect 15448 21462 15482 21838
rect 15666 21462 15700 21838
rect 15884 21462 15918 21838
rect 16102 21462 16136 21838
rect 16320 21462 16354 21838
rect 16538 21462 16572 21838
rect 16756 21462 16790 21838
rect 18718 21725 19182 21759
rect 19736 21725 20200 21759
rect 20754 21725 21218 21759
rect 21772 21725 22236 21759
rect 22790 21725 23254 21759
rect 23808 21725 24272 21759
rect 24826 21725 25290 21759
rect 25844 21725 26308 21759
rect 26862 21725 27326 21759
rect 27880 21725 28344 21759
rect 28898 21725 29362 21759
rect 29916 21725 30380 21759
rect 30934 21725 31398 21759
rect 31952 21725 32416 21759
rect 32970 21725 33434 21759
rect 14670 21369 14734 21403
rect 14888 21369 14952 21403
rect 15106 21369 15170 21403
rect 15324 21369 15388 21403
rect 15542 21369 15606 21403
rect 15760 21369 15824 21403
rect 15978 21369 16042 21403
rect 16196 21369 16260 21403
rect 16414 21369 16478 21403
rect 16632 21369 16696 21403
rect 18424 21090 18458 21666
rect 19442 21090 19476 21666
rect 20460 21090 20494 21666
rect 21478 21090 21512 21666
rect 22496 21090 22530 21666
rect 23514 21090 23548 21666
rect 24532 21090 24566 21666
rect 25550 21090 25584 21666
rect 26568 21090 26602 21666
rect 27586 21090 27620 21666
rect 28604 21090 28638 21666
rect 29622 21090 29656 21666
rect 30640 21090 30674 21666
rect 31658 21090 31692 21666
rect 32676 21090 32710 21666
rect 33694 21090 33728 21666
rect 18718 20997 19182 21031
rect 19736 20997 20200 21031
rect 20754 20997 21218 21031
rect 21772 20997 22236 21031
rect 22790 20997 23254 21031
rect 23808 20997 24272 21031
rect 24826 20997 25290 21031
rect 25844 20997 26308 21031
rect 26862 20997 27326 21031
rect 27880 20997 28344 21031
rect 28898 20997 29362 21031
rect 29916 20997 30380 21031
rect 30934 20997 31398 21031
rect 31952 20997 32416 21031
rect 32970 20997 33434 21031
rect 14670 20959 14734 20993
rect 14888 20959 14952 20993
rect 15106 20959 15170 20993
rect 15324 20959 15388 20993
rect 15542 20959 15606 20993
rect 15760 20959 15824 20993
rect 15978 20959 16042 20993
rect 16196 20959 16260 20993
rect 16414 20959 16478 20993
rect 16632 20959 16696 20993
rect 14576 20524 14610 20900
rect 14794 20524 14828 20900
rect 15012 20524 15046 20900
rect 15230 20524 15264 20900
rect 15448 20524 15482 20900
rect 15666 20524 15700 20900
rect 15884 20524 15918 20900
rect 16102 20524 16136 20900
rect 16320 20524 16354 20900
rect 16538 20524 16572 20900
rect 16756 20524 16790 20900
rect 18718 20469 19182 20503
rect 19736 20469 20200 20503
rect 20754 20469 21218 20503
rect 21772 20469 22236 20503
rect 22790 20469 23254 20503
rect 23808 20469 24272 20503
rect 24826 20469 25290 20503
rect 25844 20469 26308 20503
rect 26862 20469 27326 20503
rect 27880 20469 28344 20503
rect 28898 20469 29362 20503
rect 29916 20469 30380 20503
rect 30934 20469 31398 20503
rect 31952 20469 32416 20503
rect 32970 20469 33434 20503
rect 14670 20431 14734 20465
rect 14888 20431 14952 20465
rect 15106 20431 15170 20465
rect 15324 20431 15388 20465
rect 15542 20431 15606 20465
rect 15760 20431 15824 20465
rect 15978 20431 16042 20465
rect 16196 20431 16260 20465
rect 16414 20431 16478 20465
rect 16632 20431 16696 20465
rect 14670 20021 14734 20055
rect 14888 20021 14952 20055
rect 15106 20021 15170 20055
rect 15324 20021 15388 20055
rect 15542 20021 15606 20055
rect 15760 20021 15824 20055
rect 15978 20021 16042 20055
rect 16196 20021 16260 20055
rect 16414 20021 16478 20055
rect 16632 20021 16696 20055
rect 14576 19586 14610 19962
rect 14794 19586 14828 19962
rect 15012 19586 15046 19962
rect 15230 19586 15264 19962
rect 15448 19586 15482 19962
rect 15666 19586 15700 19962
rect 15884 19586 15918 19962
rect 16102 19586 16136 19962
rect 16320 19586 16354 19962
rect 16538 19586 16572 19962
rect 16756 19586 16790 19962
rect 18424 19834 18458 20410
rect 19442 19834 19476 20410
rect 20460 19834 20494 20410
rect 21478 19834 21512 20410
rect 22496 19834 22530 20410
rect 23514 19834 23548 20410
rect 24532 19834 24566 20410
rect 25550 19834 25584 20410
rect 26568 19834 26602 20410
rect 27586 19834 27620 20410
rect 28604 19834 28638 20410
rect 29622 19834 29656 20410
rect 30640 19834 30674 20410
rect 31658 19834 31692 20410
rect 32676 19834 32710 20410
rect 33694 19834 33728 20410
rect 18718 19741 19182 19775
rect 19736 19741 20200 19775
rect 20754 19741 21218 19775
rect 21772 19741 22236 19775
rect 22790 19741 23254 19775
rect 23808 19741 24272 19775
rect 24826 19741 25290 19775
rect 25844 19741 26308 19775
rect 26862 19741 27326 19775
rect 27880 19741 28344 19775
rect 28898 19741 29362 19775
rect 29916 19741 30380 19775
rect 30934 19741 31398 19775
rect 31952 19741 32416 19775
rect 32970 19741 33434 19775
rect 14670 19493 14734 19527
rect 14888 19493 14952 19527
rect 15106 19493 15170 19527
rect 15324 19493 15388 19527
rect 15542 19493 15606 19527
rect 15760 19493 15824 19527
rect 15978 19493 16042 19527
rect 16196 19493 16260 19527
rect 16414 19493 16478 19527
rect 16632 19493 16696 19527
rect 18718 19213 19182 19247
rect 19736 19213 20200 19247
rect 20754 19213 21218 19247
rect 21772 19213 22236 19247
rect 22790 19213 23254 19247
rect 23808 19213 24272 19247
rect 24826 19213 25290 19247
rect 25844 19213 26308 19247
rect 26862 19213 27326 19247
rect 27880 19213 28344 19247
rect 28898 19213 29362 19247
rect 29916 19213 30380 19247
rect 30934 19213 31398 19247
rect 31952 19213 32416 19247
rect 32970 19213 33434 19247
rect 14670 19083 14734 19117
rect 14888 19083 14952 19117
rect 15106 19083 15170 19117
rect 15324 19083 15388 19117
rect 15542 19083 15606 19117
rect 15760 19083 15824 19117
rect 15978 19083 16042 19117
rect 16196 19083 16260 19117
rect 16414 19083 16478 19117
rect 16632 19083 16696 19117
rect 14576 18648 14610 19024
rect 14794 18648 14828 19024
rect 15012 18648 15046 19024
rect 15230 18648 15264 19024
rect 15448 18648 15482 19024
rect 15666 18648 15700 19024
rect 15884 18648 15918 19024
rect 16102 18648 16136 19024
rect 16320 18648 16354 19024
rect 16538 18648 16572 19024
rect 16756 18648 16790 19024
rect 14670 18555 14734 18589
rect 14888 18555 14952 18589
rect 15106 18555 15170 18589
rect 15324 18555 15388 18589
rect 15542 18555 15606 18589
rect 15760 18555 15824 18589
rect 15978 18555 16042 18589
rect 16196 18555 16260 18589
rect 16414 18555 16478 18589
rect 16632 18555 16696 18589
rect 18424 18578 18458 19154
rect 19442 18578 19476 19154
rect 20460 18578 20494 19154
rect 21478 18578 21512 19154
rect 22496 18578 22530 19154
rect 23514 18578 23548 19154
rect 24532 18578 24566 19154
rect 25550 18578 25584 19154
rect 26568 18578 26602 19154
rect 27586 18578 27620 19154
rect 28604 18578 28638 19154
rect 29622 18578 29656 19154
rect 30640 18578 30674 19154
rect 31658 18578 31692 19154
rect 32676 18578 32710 19154
rect 33694 18578 33728 19154
rect 18718 18485 19182 18519
rect 19736 18485 20200 18519
rect 20754 18485 21218 18519
rect 21772 18485 22236 18519
rect 22790 18485 23254 18519
rect 23808 18485 24272 18519
rect 24826 18485 25290 18519
rect 25844 18485 26308 18519
rect 26862 18485 27326 18519
rect 27880 18485 28344 18519
rect 28898 18485 29362 18519
rect 29916 18485 30380 18519
rect 30934 18485 31398 18519
rect 31952 18485 32416 18519
rect 32970 18485 33434 18519
rect 35672 18278 35772 27642
rect 65428 28162 65490 28262
rect 65490 28162 89610 28262
rect 89610 28162 89672 28262
rect 47310 25411 47530 25412
rect 48802 25411 49004 25412
rect 47310 25378 47360 25411
rect 47360 25378 47530 25411
rect 48802 25378 48978 25411
rect 48978 25378 49004 25411
rect 49038 25315 49074 25316
rect 47262 24742 47264 25314
rect 47264 24742 47298 25314
rect 47298 24742 47300 25314
rect 47482 25275 47566 25309
rect 47740 25275 47824 25309
rect 47998 25275 48082 25309
rect 48256 25275 48340 25309
rect 48514 25275 48598 25309
rect 48772 25275 48856 25309
rect 47378 24840 47412 25216
rect 47636 24840 47670 25216
rect 47894 24840 47928 25216
rect 48152 24840 48186 25216
rect 48410 24840 48444 25216
rect 48668 24840 48702 25216
rect 48926 24840 48960 25216
rect 47482 24747 47566 24781
rect 47740 24747 47824 24781
rect 47998 24747 48082 24781
rect 48256 24747 48340 24781
rect 48514 24747 48598 24781
rect 48772 24747 48856 24781
rect 49038 24741 49040 25315
rect 49040 24741 49074 25315
rect 49177 24875 49211 24909
rect 49269 24875 49303 24909
rect 49361 24875 49395 24909
rect 49038 24740 49074 24741
rect 48802 24679 49004 24680
rect 47310 24645 47360 24678
rect 47360 24645 47530 24678
rect 48802 24646 48978 24679
rect 48978 24646 49004 24679
rect 47310 24644 47530 24645
rect 49207 24538 49255 24586
rect 49311 24597 49357 24608
rect 49311 24568 49344 24597
rect 49344 24568 49357 24597
rect 47334 24478 47542 24480
rect 48806 24478 49004 24482
rect 47334 24444 47360 24478
rect 47360 24444 47542 24478
rect 48806 24444 48978 24478
rect 48978 24444 49004 24478
rect 47334 24442 47542 24444
rect 47262 24026 47264 24382
rect 47264 24026 47298 24382
rect 47482 24342 47566 24376
rect 47740 24342 47824 24376
rect 47998 24342 48082 24376
rect 48256 24342 48340 24376
rect 48514 24342 48598 24376
rect 48772 24342 48856 24376
rect 47378 24116 47412 24292
rect 47636 24116 47670 24292
rect 47894 24116 47928 24292
rect 48152 24116 48186 24292
rect 48410 24116 48444 24292
rect 48668 24116 48702 24292
rect 48926 24116 48960 24292
rect 47482 24032 47566 24066
rect 47740 24032 47824 24066
rect 47998 24032 48082 24066
rect 48256 24032 48340 24066
rect 48514 24032 48598 24066
rect 48772 24032 48856 24066
rect 49038 24026 49040 24382
rect 49040 24026 49074 24382
rect 49074 24026 49076 24382
rect 49177 24331 49211 24365
rect 49269 24331 49303 24365
rect 49361 24331 49395 24365
rect 47332 23964 47540 23966
rect 47332 23930 47360 23964
rect 47360 23930 47540 23964
rect 48804 23930 48978 23964
rect 48978 23930 49006 23964
rect 48804 23928 49006 23930
rect 47310 23411 47530 23412
rect 48802 23411 49004 23412
rect 47310 23378 47360 23411
rect 47360 23378 47530 23411
rect 48802 23378 48978 23411
rect 48978 23378 49004 23411
rect 49038 23315 49074 23316
rect 47262 22742 47264 23314
rect 47264 22742 47298 23314
rect 47298 22742 47300 23314
rect 47482 23275 47566 23309
rect 47740 23275 47824 23309
rect 47998 23275 48082 23309
rect 48256 23275 48340 23309
rect 48514 23275 48598 23309
rect 48772 23275 48856 23309
rect 47378 22840 47412 23216
rect 47636 22840 47670 23216
rect 47894 22840 47928 23216
rect 48152 22840 48186 23216
rect 48410 22840 48444 23216
rect 48668 22840 48702 23216
rect 48926 22840 48960 23216
rect 47482 22747 47566 22781
rect 47740 22747 47824 22781
rect 47998 22747 48082 22781
rect 48256 22747 48340 22781
rect 48514 22747 48598 22781
rect 48772 22747 48856 22781
rect 49038 22741 49040 23315
rect 49040 22741 49074 23315
rect 49177 22875 49211 22909
rect 49269 22875 49303 22909
rect 49361 22875 49395 22909
rect 49038 22740 49074 22741
rect 48802 22679 49004 22680
rect 47310 22645 47360 22678
rect 47360 22645 47530 22678
rect 48802 22646 48978 22679
rect 48978 22646 49004 22679
rect 47310 22644 47530 22645
rect 49207 22538 49255 22586
rect 49311 22597 49357 22608
rect 49311 22568 49344 22597
rect 49344 22568 49357 22597
rect 47334 22478 47542 22480
rect 48806 22478 49004 22482
rect 47334 22444 47360 22478
rect 47360 22444 47542 22478
rect 48806 22444 48978 22478
rect 48978 22444 49004 22478
rect 47334 22442 47542 22444
rect 47262 22026 47264 22382
rect 47264 22026 47298 22382
rect 47482 22342 47566 22376
rect 47740 22342 47824 22376
rect 47998 22342 48082 22376
rect 48256 22342 48340 22376
rect 48514 22342 48598 22376
rect 48772 22342 48856 22376
rect 47378 22116 47412 22292
rect 47636 22116 47670 22292
rect 47894 22116 47928 22292
rect 48152 22116 48186 22292
rect 48410 22116 48444 22292
rect 48668 22116 48702 22292
rect 48926 22116 48960 22292
rect 47482 22032 47566 22066
rect 47740 22032 47824 22066
rect 47998 22032 48082 22066
rect 48256 22032 48340 22066
rect 48514 22032 48598 22066
rect 48772 22032 48856 22066
rect 49038 22026 49040 22382
rect 49040 22026 49074 22382
rect 49074 22026 49076 22382
rect 49177 22331 49211 22365
rect 49269 22331 49303 22365
rect 49361 22331 49395 22365
rect 47332 21964 47540 21966
rect 47332 21930 47360 21964
rect 47360 21930 47540 21964
rect 48804 21930 48978 21964
rect 48978 21930 49006 21964
rect 48804 21928 49006 21930
rect 11428 17658 11490 17758
rect 11490 17658 35610 17758
rect 35610 17658 35672 17758
rect 65328 18278 65428 27642
rect 71732 27027 72196 27061
rect 72750 27027 73214 27061
rect 73768 27027 74232 27061
rect 74786 27027 75250 27061
rect 75804 27027 76268 27061
rect 76822 27027 77286 27061
rect 77840 27027 78304 27061
rect 78858 27027 79322 27061
rect 79876 27027 80340 27061
rect 80894 27027 81358 27061
rect 81912 27027 82376 27061
rect 82930 27027 83394 27061
rect 83948 27027 84412 27061
rect 84966 27027 85430 27061
rect 85984 27027 86448 27061
rect 87002 27027 87466 27061
rect 71438 26392 71472 26968
rect 72456 26392 72490 26968
rect 73474 26392 73508 26968
rect 74492 26392 74526 26968
rect 75510 26392 75544 26968
rect 76528 26392 76562 26968
rect 77546 26392 77580 26968
rect 78564 26392 78598 26968
rect 79582 26392 79616 26968
rect 80600 26392 80634 26968
rect 81618 26392 81652 26968
rect 82636 26392 82670 26968
rect 83654 26392 83688 26968
rect 84672 26392 84706 26968
rect 85690 26392 85724 26968
rect 86708 26392 86742 26968
rect 87726 26392 87760 26968
rect 71732 26299 72196 26333
rect 72750 26299 73214 26333
rect 73768 26299 74232 26333
rect 74786 26299 75250 26333
rect 75804 26299 76268 26333
rect 76822 26299 77286 26333
rect 77840 26299 78304 26333
rect 78858 26299 79322 26333
rect 79876 26299 80340 26333
rect 80894 26299 81358 26333
rect 81912 26299 82376 26333
rect 82930 26299 83394 26333
rect 83948 26299 84412 26333
rect 84966 26299 85430 26333
rect 85984 26299 86448 26333
rect 87002 26299 87466 26333
rect 71732 25891 72196 25925
rect 72750 25891 73214 25925
rect 73768 25891 74232 25925
rect 74786 25891 75250 25925
rect 75804 25891 76268 25925
rect 76822 25891 77286 25925
rect 77840 25891 78304 25925
rect 78858 25891 79322 25925
rect 79876 25891 80340 25925
rect 80894 25891 81358 25925
rect 81912 25891 82376 25925
rect 82930 25891 83394 25925
rect 83948 25891 84412 25925
rect 84966 25891 85430 25925
rect 85984 25891 86448 25925
rect 87002 25891 87466 25925
rect 71438 25256 71472 25832
rect 72456 25256 72490 25832
rect 73474 25256 73508 25832
rect 74492 25256 74526 25832
rect 75510 25256 75544 25832
rect 76528 25256 76562 25832
rect 77546 25256 77580 25832
rect 78564 25256 78598 25832
rect 79582 25256 79616 25832
rect 80600 25256 80634 25832
rect 81618 25256 81652 25832
rect 82636 25256 82670 25832
rect 83654 25256 83688 25832
rect 84672 25256 84706 25832
rect 85690 25256 85724 25832
rect 86708 25256 86742 25832
rect 87726 25256 87760 25832
rect 71732 25163 72196 25197
rect 72750 25163 73214 25197
rect 73768 25163 74232 25197
rect 74786 25163 75250 25197
rect 75804 25163 76268 25197
rect 76822 25163 77286 25197
rect 77840 25163 78304 25197
rect 78858 25163 79322 25197
rect 79876 25163 80340 25197
rect 80894 25163 81358 25197
rect 81912 25163 82376 25197
rect 82930 25163 83394 25197
rect 83948 25163 84412 25197
rect 84966 25163 85430 25197
rect 85984 25163 86448 25197
rect 87002 25163 87466 25197
rect 71732 24755 72196 24789
rect 72750 24755 73214 24789
rect 73768 24755 74232 24789
rect 74786 24755 75250 24789
rect 75804 24755 76268 24789
rect 76822 24755 77286 24789
rect 77840 24755 78304 24789
rect 78858 24755 79322 24789
rect 79876 24755 80340 24789
rect 80894 24755 81358 24789
rect 81912 24755 82376 24789
rect 82930 24755 83394 24789
rect 83948 24755 84412 24789
rect 84966 24755 85430 24789
rect 85984 24755 86448 24789
rect 87002 24755 87466 24789
rect 71438 24120 71472 24696
rect 72456 24120 72490 24696
rect 73474 24120 73508 24696
rect 74492 24120 74526 24696
rect 75510 24120 75544 24696
rect 76528 24120 76562 24696
rect 77546 24120 77580 24696
rect 78564 24120 78598 24696
rect 79582 24120 79616 24696
rect 80600 24120 80634 24696
rect 81618 24120 81652 24696
rect 82636 24120 82670 24696
rect 83654 24120 83688 24696
rect 84672 24120 84706 24696
rect 85690 24120 85724 24696
rect 86708 24120 86742 24696
rect 87726 24120 87760 24696
rect 71732 24027 72196 24061
rect 72750 24027 73214 24061
rect 73768 24027 74232 24061
rect 74786 24027 75250 24061
rect 75804 24027 76268 24061
rect 76822 24027 77286 24061
rect 77840 24027 78304 24061
rect 78858 24027 79322 24061
rect 79876 24027 80340 24061
rect 80894 24027 81358 24061
rect 81912 24027 82376 24061
rect 82930 24027 83394 24061
rect 83948 24027 84412 24061
rect 84966 24027 85430 24061
rect 85984 24027 86448 24061
rect 87002 24027 87466 24061
rect 72718 22981 73182 23015
rect 73736 22981 74200 23015
rect 74754 22981 75218 23015
rect 75772 22981 76236 23015
rect 76790 22981 77254 23015
rect 77808 22981 78272 23015
rect 78826 22981 79290 23015
rect 79844 22981 80308 23015
rect 80862 22981 81326 23015
rect 81880 22981 82344 23015
rect 82898 22981 83362 23015
rect 83916 22981 84380 23015
rect 84934 22981 85398 23015
rect 85952 22981 86416 23015
rect 86970 22981 87434 23015
rect 72424 22346 72458 22922
rect 73442 22346 73476 22922
rect 74460 22346 74494 22922
rect 75478 22346 75512 22922
rect 76496 22346 76530 22922
rect 77514 22346 77548 22922
rect 78532 22346 78566 22922
rect 79550 22346 79584 22922
rect 80568 22346 80602 22922
rect 81586 22346 81620 22922
rect 82604 22346 82638 22922
rect 83622 22346 83656 22922
rect 84640 22346 84674 22922
rect 85658 22346 85692 22922
rect 86676 22346 86710 22922
rect 87694 22346 87728 22922
rect 72718 22253 73182 22287
rect 73736 22253 74200 22287
rect 74754 22253 75218 22287
rect 75772 22253 76236 22287
rect 76790 22253 77254 22287
rect 77808 22253 78272 22287
rect 78826 22253 79290 22287
rect 79844 22253 80308 22287
rect 80862 22253 81326 22287
rect 81880 22253 82344 22287
rect 82898 22253 83362 22287
rect 83916 22253 84380 22287
rect 84934 22253 85398 22287
rect 85952 22253 86416 22287
rect 86970 22253 87434 22287
rect 68670 21897 68734 21931
rect 68888 21897 68952 21931
rect 69106 21897 69170 21931
rect 69324 21897 69388 21931
rect 69542 21897 69606 21931
rect 69760 21897 69824 21931
rect 69978 21897 70042 21931
rect 70196 21897 70260 21931
rect 70414 21897 70478 21931
rect 70632 21897 70696 21931
rect 68576 21462 68610 21838
rect 68794 21462 68828 21838
rect 69012 21462 69046 21838
rect 69230 21462 69264 21838
rect 69448 21462 69482 21838
rect 69666 21462 69700 21838
rect 69884 21462 69918 21838
rect 70102 21462 70136 21838
rect 70320 21462 70354 21838
rect 70538 21462 70572 21838
rect 70756 21462 70790 21838
rect 72718 21725 73182 21759
rect 73736 21725 74200 21759
rect 74754 21725 75218 21759
rect 75772 21725 76236 21759
rect 76790 21725 77254 21759
rect 77808 21725 78272 21759
rect 78826 21725 79290 21759
rect 79844 21725 80308 21759
rect 80862 21725 81326 21759
rect 81880 21725 82344 21759
rect 82898 21725 83362 21759
rect 83916 21725 84380 21759
rect 84934 21725 85398 21759
rect 85952 21725 86416 21759
rect 86970 21725 87434 21759
rect 68670 21369 68734 21403
rect 68888 21369 68952 21403
rect 69106 21369 69170 21403
rect 69324 21369 69388 21403
rect 69542 21369 69606 21403
rect 69760 21369 69824 21403
rect 69978 21369 70042 21403
rect 70196 21369 70260 21403
rect 70414 21369 70478 21403
rect 70632 21369 70696 21403
rect 72424 21090 72458 21666
rect 73442 21090 73476 21666
rect 74460 21090 74494 21666
rect 75478 21090 75512 21666
rect 76496 21090 76530 21666
rect 77514 21090 77548 21666
rect 78532 21090 78566 21666
rect 79550 21090 79584 21666
rect 80568 21090 80602 21666
rect 81586 21090 81620 21666
rect 82604 21090 82638 21666
rect 83622 21090 83656 21666
rect 84640 21090 84674 21666
rect 85658 21090 85692 21666
rect 86676 21090 86710 21666
rect 87694 21090 87728 21666
rect 72718 20997 73182 21031
rect 73736 20997 74200 21031
rect 74754 20997 75218 21031
rect 75772 20997 76236 21031
rect 76790 20997 77254 21031
rect 77808 20997 78272 21031
rect 78826 20997 79290 21031
rect 79844 20997 80308 21031
rect 80862 20997 81326 21031
rect 81880 20997 82344 21031
rect 82898 20997 83362 21031
rect 83916 20997 84380 21031
rect 84934 20997 85398 21031
rect 85952 20997 86416 21031
rect 86970 20997 87434 21031
rect 68670 20959 68734 20993
rect 68888 20959 68952 20993
rect 69106 20959 69170 20993
rect 69324 20959 69388 20993
rect 69542 20959 69606 20993
rect 69760 20959 69824 20993
rect 69978 20959 70042 20993
rect 70196 20959 70260 20993
rect 70414 20959 70478 20993
rect 70632 20959 70696 20993
rect 68576 20524 68610 20900
rect 68794 20524 68828 20900
rect 69012 20524 69046 20900
rect 69230 20524 69264 20900
rect 69448 20524 69482 20900
rect 69666 20524 69700 20900
rect 69884 20524 69918 20900
rect 70102 20524 70136 20900
rect 70320 20524 70354 20900
rect 70538 20524 70572 20900
rect 70756 20524 70790 20900
rect 72718 20469 73182 20503
rect 73736 20469 74200 20503
rect 74754 20469 75218 20503
rect 75772 20469 76236 20503
rect 76790 20469 77254 20503
rect 77808 20469 78272 20503
rect 78826 20469 79290 20503
rect 79844 20469 80308 20503
rect 80862 20469 81326 20503
rect 81880 20469 82344 20503
rect 82898 20469 83362 20503
rect 83916 20469 84380 20503
rect 84934 20469 85398 20503
rect 85952 20469 86416 20503
rect 86970 20469 87434 20503
rect 68670 20431 68734 20465
rect 68888 20431 68952 20465
rect 69106 20431 69170 20465
rect 69324 20431 69388 20465
rect 69542 20431 69606 20465
rect 69760 20431 69824 20465
rect 69978 20431 70042 20465
rect 70196 20431 70260 20465
rect 70414 20431 70478 20465
rect 70632 20431 70696 20465
rect 68670 20021 68734 20055
rect 68888 20021 68952 20055
rect 69106 20021 69170 20055
rect 69324 20021 69388 20055
rect 69542 20021 69606 20055
rect 69760 20021 69824 20055
rect 69978 20021 70042 20055
rect 70196 20021 70260 20055
rect 70414 20021 70478 20055
rect 70632 20021 70696 20055
rect 68576 19586 68610 19962
rect 68794 19586 68828 19962
rect 69012 19586 69046 19962
rect 69230 19586 69264 19962
rect 69448 19586 69482 19962
rect 69666 19586 69700 19962
rect 69884 19586 69918 19962
rect 70102 19586 70136 19962
rect 70320 19586 70354 19962
rect 70538 19586 70572 19962
rect 70756 19586 70790 19962
rect 72424 19834 72458 20410
rect 73442 19834 73476 20410
rect 74460 19834 74494 20410
rect 75478 19834 75512 20410
rect 76496 19834 76530 20410
rect 77514 19834 77548 20410
rect 78532 19834 78566 20410
rect 79550 19834 79584 20410
rect 80568 19834 80602 20410
rect 81586 19834 81620 20410
rect 82604 19834 82638 20410
rect 83622 19834 83656 20410
rect 84640 19834 84674 20410
rect 85658 19834 85692 20410
rect 86676 19834 86710 20410
rect 87694 19834 87728 20410
rect 72718 19741 73182 19775
rect 73736 19741 74200 19775
rect 74754 19741 75218 19775
rect 75772 19741 76236 19775
rect 76790 19741 77254 19775
rect 77808 19741 78272 19775
rect 78826 19741 79290 19775
rect 79844 19741 80308 19775
rect 80862 19741 81326 19775
rect 81880 19741 82344 19775
rect 82898 19741 83362 19775
rect 83916 19741 84380 19775
rect 84934 19741 85398 19775
rect 85952 19741 86416 19775
rect 86970 19741 87434 19775
rect 68670 19493 68734 19527
rect 68888 19493 68952 19527
rect 69106 19493 69170 19527
rect 69324 19493 69388 19527
rect 69542 19493 69606 19527
rect 69760 19493 69824 19527
rect 69978 19493 70042 19527
rect 70196 19493 70260 19527
rect 70414 19493 70478 19527
rect 70632 19493 70696 19527
rect 72718 19213 73182 19247
rect 73736 19213 74200 19247
rect 74754 19213 75218 19247
rect 75772 19213 76236 19247
rect 76790 19213 77254 19247
rect 77808 19213 78272 19247
rect 78826 19213 79290 19247
rect 79844 19213 80308 19247
rect 80862 19213 81326 19247
rect 81880 19213 82344 19247
rect 82898 19213 83362 19247
rect 83916 19213 84380 19247
rect 84934 19213 85398 19247
rect 85952 19213 86416 19247
rect 86970 19213 87434 19247
rect 68670 19083 68734 19117
rect 68888 19083 68952 19117
rect 69106 19083 69170 19117
rect 69324 19083 69388 19117
rect 69542 19083 69606 19117
rect 69760 19083 69824 19117
rect 69978 19083 70042 19117
rect 70196 19083 70260 19117
rect 70414 19083 70478 19117
rect 70632 19083 70696 19117
rect 68576 18648 68610 19024
rect 68794 18648 68828 19024
rect 69012 18648 69046 19024
rect 69230 18648 69264 19024
rect 69448 18648 69482 19024
rect 69666 18648 69700 19024
rect 69884 18648 69918 19024
rect 70102 18648 70136 19024
rect 70320 18648 70354 19024
rect 70538 18648 70572 19024
rect 70756 18648 70790 19024
rect 68670 18555 68734 18589
rect 68888 18555 68952 18589
rect 69106 18555 69170 18589
rect 69324 18555 69388 18589
rect 69542 18555 69606 18589
rect 69760 18555 69824 18589
rect 69978 18555 70042 18589
rect 70196 18555 70260 18589
rect 70414 18555 70478 18589
rect 70632 18555 70696 18589
rect 72424 18578 72458 19154
rect 73442 18578 73476 19154
rect 74460 18578 74494 19154
rect 75478 18578 75512 19154
rect 76496 18578 76530 19154
rect 77514 18578 77548 19154
rect 78532 18578 78566 19154
rect 79550 18578 79584 19154
rect 80568 18578 80602 19154
rect 81586 18578 81620 19154
rect 82604 18578 82638 19154
rect 83622 18578 83656 19154
rect 84640 18578 84674 19154
rect 85658 18578 85692 19154
rect 86676 18578 86710 19154
rect 87694 18578 87728 19154
rect 72718 18485 73182 18519
rect 73736 18485 74200 18519
rect 74754 18485 75218 18519
rect 75772 18485 76236 18519
rect 76790 18485 77254 18519
rect 77808 18485 78272 18519
rect 78826 18485 79290 18519
rect 79844 18485 80308 18519
rect 80862 18485 81326 18519
rect 81880 18485 82344 18519
rect 82898 18485 83362 18519
rect 83916 18485 84380 18519
rect 84934 18485 85398 18519
rect 85952 18485 86416 18519
rect 86970 18485 87434 18519
rect 89672 18278 89772 27642
rect 65428 17658 65490 17758
rect 65490 17658 89610 17758
rect 89610 17658 89672 17758
rect -13048 16281 -12828 16282
rect -11556 16281 -11354 16282
rect -10448 16281 -10228 16282
rect -8956 16281 -8754 16282
rect -13048 16248 -12998 16281
rect -12998 16248 -12828 16281
rect -11556 16248 -11380 16281
rect -11380 16248 -11354 16281
rect -11320 16185 -11284 16186
rect -13096 15612 -13094 16184
rect -13094 15612 -13060 16184
rect -13060 15612 -13058 16184
rect -12876 16145 -12792 16179
rect -12618 16145 -12534 16179
rect -12360 16145 -12276 16179
rect -12102 16145 -12018 16179
rect -11844 16145 -11760 16179
rect -11586 16145 -11502 16179
rect -12980 15710 -12946 16086
rect -12722 15710 -12688 16086
rect -12464 15710 -12430 16086
rect -12206 15710 -12172 16086
rect -11948 15710 -11914 16086
rect -11690 15710 -11656 16086
rect -11432 15710 -11398 16086
rect -12876 15617 -12792 15651
rect -12618 15617 -12534 15651
rect -12360 15617 -12276 15651
rect -12102 15617 -12018 15651
rect -11844 15617 -11760 15651
rect -11586 15617 -11502 15651
rect -11320 15611 -11318 16185
rect -11318 15611 -11284 16185
rect -10448 16248 -10398 16281
rect -10398 16248 -10228 16281
rect -8956 16248 -8780 16281
rect -8780 16248 -8754 16281
rect -8720 16185 -8684 16186
rect -11181 15745 -11147 15779
rect -11089 15745 -11055 15779
rect -10997 15745 -10963 15779
rect -11320 15610 -11284 15611
rect -11556 15549 -11354 15550
rect -13048 15515 -12998 15548
rect -12998 15515 -12828 15548
rect -11556 15516 -11380 15549
rect -11380 15516 -11354 15549
rect -10496 15612 -10494 16184
rect -10494 15612 -10460 16184
rect -10460 15612 -10458 16184
rect -10276 16145 -10192 16179
rect -10018 16145 -9934 16179
rect -9760 16145 -9676 16179
rect -9502 16145 -9418 16179
rect -9244 16145 -9160 16179
rect -8986 16145 -8902 16179
rect -10380 15710 -10346 16086
rect -10122 15710 -10088 16086
rect -9864 15710 -9830 16086
rect -9606 15710 -9572 16086
rect -9348 15710 -9314 16086
rect -9090 15710 -9056 16086
rect -8832 15710 -8798 16086
rect -10276 15617 -10192 15651
rect -10018 15617 -9934 15651
rect -9760 15617 -9676 15651
rect -9502 15617 -9418 15651
rect -9244 15617 -9160 15651
rect -8986 15617 -8902 15651
rect -8720 15611 -8718 16185
rect -8718 15611 -8684 16185
rect -8581 15745 -8547 15779
rect -8489 15745 -8455 15779
rect -8397 15745 -8363 15779
rect -8081 15745 -8047 15779
rect -7989 15745 -7955 15779
rect -7897 15745 -7863 15779
rect -8720 15610 -8684 15611
rect -8956 15549 -8754 15550
rect -10448 15515 -10398 15548
rect -10398 15515 -10228 15548
rect -8956 15516 -8780 15549
rect -8780 15516 -8754 15549
rect -13048 15514 -12828 15515
rect -10448 15514 -10228 15515
rect -11151 15408 -11103 15456
rect -11047 15467 -11001 15478
rect -11047 15438 -11014 15467
rect -11014 15438 -11001 15467
rect -8551 15408 -8503 15456
rect -8447 15467 -8401 15478
rect -8447 15438 -8414 15467
rect -8414 15438 -8401 15467
rect -8052 15430 -8004 15478
rect -7950 15467 -7902 15482
rect -7950 15434 -7948 15467
rect -7948 15434 -7914 15467
rect -7914 15434 -7902 15467
rect -13024 15348 -12816 15350
rect -11552 15348 -11354 15352
rect -13024 15314 -12998 15348
rect -12998 15314 -12816 15348
rect -11552 15314 -11380 15348
rect -11380 15314 -11354 15348
rect -13024 15312 -12816 15314
rect -10424 15348 -10216 15350
rect -8952 15348 -8754 15352
rect -13096 14896 -13094 15252
rect -13094 14896 -13060 15252
rect -12876 15212 -12792 15246
rect -12618 15212 -12534 15246
rect -12360 15212 -12276 15246
rect -12102 15212 -12018 15246
rect -11844 15212 -11760 15246
rect -11586 15212 -11502 15246
rect -12980 14986 -12946 15162
rect -12722 14986 -12688 15162
rect -12464 14986 -12430 15162
rect -12206 14986 -12172 15162
rect -11948 14986 -11914 15162
rect -11690 14986 -11656 15162
rect -11432 14986 -11398 15162
rect -12876 14902 -12792 14936
rect -12618 14902 -12534 14936
rect -12360 14902 -12276 14936
rect -12102 14902 -12018 14936
rect -11844 14902 -11760 14936
rect -11586 14902 -11502 14936
rect -11320 14896 -11318 15252
rect -11318 14896 -11284 15252
rect -11284 14896 -11282 15252
rect -10424 15314 -10398 15348
rect -10398 15314 -10216 15348
rect -8952 15314 -8780 15348
rect -8780 15314 -8754 15348
rect -10424 15312 -10216 15314
rect -11181 15201 -11147 15235
rect -11089 15201 -11055 15235
rect -10997 15201 -10963 15235
rect -10496 14896 -10494 15252
rect -10494 14896 -10460 15252
rect -10276 15212 -10192 15246
rect -10018 15212 -9934 15246
rect -9760 15212 -9676 15246
rect -9502 15212 -9418 15246
rect -9244 15212 -9160 15246
rect -8986 15212 -8902 15246
rect -10380 14986 -10346 15162
rect -10122 14986 -10088 15162
rect -9864 14986 -9830 15162
rect -9606 14986 -9572 15162
rect -9348 14986 -9314 15162
rect -9090 14986 -9056 15162
rect -8832 14986 -8798 15162
rect -10276 14902 -10192 14936
rect -10018 14902 -9934 14936
rect -9760 14902 -9676 14936
rect -9502 14902 -9418 14936
rect -9244 14902 -9160 14936
rect -8986 14902 -8902 14936
rect -8720 14896 -8718 15252
rect -8718 14896 -8684 15252
rect -8684 14896 -8682 15252
rect -8581 15201 -8547 15235
rect -8489 15201 -8455 15235
rect -8397 15201 -8363 15235
rect -8081 15201 -8047 15235
rect -7989 15201 -7955 15235
rect -7897 15201 -7863 15235
rect -1272 15262 -1210 15362
rect -1210 15262 35710 15362
rect 35710 15262 35772 15362
rect -13026 14834 -12818 14836
rect -13026 14800 -12998 14834
rect -12998 14800 -12818 14834
rect -11554 14800 -11380 14834
rect -11380 14800 -11352 14834
rect -10426 14834 -10218 14836
rect -10426 14800 -10398 14834
rect -10398 14800 -10218 14834
rect -8954 14800 -8780 14834
rect -8780 14800 -8752 14834
rect -11554 14798 -11352 14800
rect -8954 14798 -8752 14800
rect 13826 14860 14290 14894
rect 14844 14860 15308 14894
rect 15862 14860 16326 14894
rect 16880 14860 17344 14894
rect 17898 14860 18362 14894
rect 18916 14860 19380 14894
rect 19934 14860 20398 14894
rect 20952 14860 21416 14894
rect 21970 14860 22434 14894
rect 22988 14860 23452 14894
rect 24006 14860 24470 14894
rect 25024 14860 25488 14894
rect 26042 14860 26506 14894
rect 27060 14860 27524 14894
rect 28078 14860 28542 14894
rect 29096 14860 29560 14894
rect 30114 14860 30578 14894
rect 31132 14860 31596 14894
rect 32150 14860 32614 14894
rect 33168 14860 33632 14894
rect -1372 210 -1272 14470
rect 13532 14234 13566 14810
rect 14550 14234 14584 14810
rect 15568 14234 15602 14810
rect 16586 14234 16620 14810
rect 17604 14234 17638 14810
rect 18622 14234 18656 14810
rect 19640 14234 19674 14810
rect 20658 14234 20692 14810
rect 21676 14234 21710 14810
rect 22694 14234 22728 14810
rect 23712 14234 23746 14810
rect 24730 14234 24764 14810
rect 25748 14234 25782 14810
rect 26766 14234 26800 14810
rect 27784 14234 27818 14810
rect 28802 14234 28836 14810
rect 29820 14234 29854 14810
rect 30838 14234 30872 14810
rect 31856 14234 31890 14810
rect 32874 14234 32908 14810
rect 33892 14234 33926 14810
rect 13826 14150 14290 14184
rect 14844 14150 15308 14184
rect 15862 14150 16326 14184
rect 16880 14150 17344 14184
rect 17898 14150 18362 14184
rect 18916 14150 19380 14184
rect 19934 14150 20398 14184
rect 20952 14150 21416 14184
rect 21970 14150 22434 14184
rect 22988 14150 23452 14184
rect 24006 14150 24470 14184
rect 25024 14150 25488 14184
rect 26042 14150 26506 14184
rect 27060 14150 27524 14184
rect 28078 14150 28542 14184
rect 29096 14150 29560 14184
rect 30114 14150 30578 14184
rect 31132 14150 31596 14184
rect 32150 14150 32614 14184
rect 33168 14150 33632 14184
rect 2060 14066 2524 14100
rect 3078 14066 3542 14100
rect 4096 14066 4560 14100
rect 5114 14066 5578 14100
rect 6132 14066 6596 14100
rect 7150 14066 7614 14100
rect 8168 14066 8632 14100
rect 9186 14066 9650 14100
rect 10204 14066 10668 14100
rect 1766 13440 1800 14016
rect 2784 13440 2818 14016
rect 3802 13440 3836 14016
rect 4820 13440 4854 14016
rect 5838 13440 5872 14016
rect 6856 13440 6890 14016
rect 7874 13440 7908 14016
rect 8892 13440 8926 14016
rect 9910 13440 9944 14016
rect 10928 13440 10962 14016
rect 13826 13626 14290 13660
rect 14844 13626 15308 13660
rect 15862 13626 16326 13660
rect 16880 13626 17344 13660
rect 17898 13626 18362 13660
rect 18916 13626 19380 13660
rect 19934 13626 20398 13660
rect 20952 13626 21416 13660
rect 21970 13626 22434 13660
rect 22988 13626 23452 13660
rect 24006 13626 24470 13660
rect 25024 13626 25488 13660
rect 26042 13626 26506 13660
rect 27060 13626 27524 13660
rect 28078 13626 28542 13660
rect 29096 13626 29560 13660
rect 30114 13626 30578 13660
rect 31132 13626 31596 13660
rect 32150 13626 32614 13660
rect 33168 13626 33632 13660
rect 2060 13356 2524 13390
rect 3078 13356 3542 13390
rect 2060 13248 2524 13282
rect 4096 13356 4560 13390
rect 3078 13248 3542 13282
rect 5114 13356 5578 13390
rect 4096 13248 4560 13282
rect 6132 13356 6596 13390
rect 5114 13248 5578 13282
rect 7150 13356 7614 13390
rect 6132 13248 6596 13282
rect 8168 13356 8632 13390
rect 7150 13248 7614 13282
rect 9186 13356 9650 13390
rect 8168 13248 8632 13282
rect 10204 13356 10668 13390
rect 9186 13248 9650 13282
rect 10204 13248 10668 13282
rect 1766 12622 1800 13198
rect 2784 12622 2818 13198
rect 3802 12622 3836 13198
rect 4820 12622 4854 13198
rect 5838 12622 5872 13198
rect 6856 12622 6890 13198
rect 7874 12622 7908 13198
rect 8892 12622 8926 13198
rect 9910 12622 9944 13198
rect 10928 12622 10962 13198
rect 13532 13000 13566 13576
rect 14550 13000 14584 13576
rect 15568 13000 15602 13576
rect 16586 13000 16620 13576
rect 17604 13000 17638 13576
rect 18622 13000 18656 13576
rect 19640 13000 19674 13576
rect 20658 13000 20692 13576
rect 21676 13000 21710 13576
rect 22694 13000 22728 13576
rect 23712 13000 23746 13576
rect 24730 13000 24764 13576
rect 25748 13000 25782 13576
rect 26766 13000 26800 13576
rect 27784 13000 27818 13576
rect 28802 13000 28836 13576
rect 29820 13000 29854 13576
rect 30838 13000 30872 13576
rect 31856 13000 31890 13576
rect 32874 13000 32908 13576
rect 33892 13000 33926 13576
rect 13826 12916 14290 12950
rect 14844 12916 15308 12950
rect 15862 12916 16326 12950
rect 16880 12916 17344 12950
rect 17898 12916 18362 12950
rect 18916 12916 19380 12950
rect 19934 12916 20398 12950
rect 20952 12916 21416 12950
rect 21970 12916 22434 12950
rect 22988 12916 23452 12950
rect 24006 12916 24470 12950
rect 25024 12916 25488 12950
rect 26042 12916 26506 12950
rect 27060 12916 27524 12950
rect 28078 12916 28542 12950
rect 29096 12916 29560 12950
rect 30114 12916 30578 12950
rect 31132 12916 31596 12950
rect 32150 12916 32614 12950
rect 33168 12916 33632 12950
rect 2060 12538 2524 12572
rect 3078 12538 3542 12572
rect 2060 12430 2524 12464
rect 4096 12538 4560 12572
rect 3078 12430 3542 12464
rect 5114 12538 5578 12572
rect 4096 12430 4560 12464
rect 6132 12538 6596 12572
rect 5114 12430 5578 12464
rect 7150 12538 7614 12572
rect 6132 12430 6596 12464
rect 8168 12538 8632 12572
rect 7150 12430 7614 12464
rect 9186 12538 9650 12572
rect 8168 12430 8632 12464
rect 10204 12538 10668 12572
rect 9186 12430 9650 12464
rect 10204 12430 10668 12464
rect 1766 11804 1800 12380
rect 2784 11804 2818 12380
rect 3802 11804 3836 12380
rect 4820 11804 4854 12380
rect 5838 11804 5872 12380
rect 6856 11804 6890 12380
rect 7874 11804 7908 12380
rect 8892 11804 8926 12380
rect 9910 11804 9944 12380
rect 13826 12394 14290 12428
rect 14844 12394 15308 12428
rect 15862 12394 16326 12428
rect 16880 12394 17344 12428
rect 17898 12394 18362 12428
rect 18916 12394 19380 12428
rect 19934 12394 20398 12428
rect 20952 12394 21416 12428
rect 21970 12394 22434 12428
rect 22988 12394 23452 12428
rect 24006 12394 24470 12428
rect 25024 12394 25488 12428
rect 26042 12394 26506 12428
rect 27060 12394 27524 12428
rect 28078 12394 28542 12428
rect 29096 12394 29560 12428
rect 30114 12394 30578 12428
rect 31132 12394 31596 12428
rect 32150 12394 32614 12428
rect 33168 12394 33632 12428
rect 10928 11804 10962 12380
rect 13532 11768 13566 12344
rect 2060 11720 2524 11754
rect 3078 11720 3542 11754
rect 2060 11612 2524 11646
rect 4096 11720 4560 11754
rect 3078 11612 3542 11646
rect 5114 11720 5578 11754
rect 4096 11612 4560 11646
rect 6132 11720 6596 11754
rect 5114 11612 5578 11646
rect 7150 11720 7614 11754
rect 6132 11612 6596 11646
rect 8168 11720 8632 11754
rect 7150 11612 7614 11646
rect 9186 11720 9650 11754
rect 8168 11612 8632 11646
rect 10204 11720 10668 11754
rect 14550 11768 14584 12344
rect 15568 11768 15602 12344
rect 16586 11768 16620 12344
rect 17604 11768 17638 12344
rect 18622 11768 18656 12344
rect 19640 11768 19674 12344
rect 20658 11768 20692 12344
rect 21676 11768 21710 12344
rect 22694 11768 22728 12344
rect 23712 11768 23746 12344
rect 24730 11768 24764 12344
rect 25748 11768 25782 12344
rect 26766 11768 26800 12344
rect 27784 11768 27818 12344
rect 28802 11768 28836 12344
rect 29820 11768 29854 12344
rect 30838 11768 30872 12344
rect 31856 11768 31890 12344
rect 32874 11768 32908 12344
rect 33892 11768 33926 12344
rect 9186 11612 9650 11646
rect 13826 11684 14290 11718
rect 14844 11684 15308 11718
rect 15862 11684 16326 11718
rect 16880 11684 17344 11718
rect 17898 11684 18362 11718
rect 18916 11684 19380 11718
rect 19934 11684 20398 11718
rect 20952 11684 21416 11718
rect 21970 11684 22434 11718
rect 22988 11684 23452 11718
rect 24006 11684 24470 11718
rect 25024 11684 25488 11718
rect 26042 11684 26506 11718
rect 27060 11684 27524 11718
rect 28078 11684 28542 11718
rect 29096 11684 29560 11718
rect 30114 11684 30578 11718
rect 31132 11684 31596 11718
rect 32150 11684 32614 11718
rect 33168 11684 33632 11718
rect 10204 11612 10668 11646
rect 1766 10986 1800 11562
rect 2784 10986 2818 11562
rect 3802 10986 3836 11562
rect 4820 10986 4854 11562
rect 5838 10986 5872 11562
rect 6856 10986 6890 11562
rect 7874 10986 7908 11562
rect 8892 10986 8926 11562
rect 9910 10986 9944 11562
rect 10928 10986 10962 11562
rect 13824 11160 14288 11194
rect 14842 11160 15306 11194
rect 15860 11160 16324 11194
rect 16878 11160 17342 11194
rect 17896 11160 18360 11194
rect 18914 11160 19378 11194
rect 19932 11160 20396 11194
rect 20950 11160 21414 11194
rect 21968 11160 22432 11194
rect 22986 11160 23450 11194
rect 24004 11160 24468 11194
rect 25022 11160 25486 11194
rect 26040 11160 26504 11194
rect 27058 11160 27522 11194
rect 28076 11160 28540 11194
rect 29094 11160 29558 11194
rect 30112 11160 30576 11194
rect 31130 11160 31594 11194
rect 32148 11160 32612 11194
rect 33166 11160 33630 11194
rect 2060 10902 2524 10936
rect 3078 10902 3542 10936
rect 2060 10794 2524 10828
rect 4096 10902 4560 10936
rect 3078 10794 3542 10828
rect 5114 10902 5578 10936
rect 4096 10794 4560 10828
rect 6132 10902 6596 10936
rect 5114 10794 5578 10828
rect 7150 10902 7614 10936
rect 6132 10794 6596 10828
rect 8168 10902 8632 10936
rect 7150 10794 7614 10828
rect 9186 10902 9650 10936
rect 8168 10794 8632 10828
rect 10204 10902 10668 10936
rect 9186 10794 9650 10828
rect 10204 10794 10668 10828
rect 1766 10168 1800 10744
rect 2784 10168 2818 10744
rect 3802 10168 3836 10744
rect 4820 10168 4854 10744
rect 5838 10168 5872 10744
rect 6856 10168 6890 10744
rect 7874 10168 7908 10744
rect 8892 10168 8926 10744
rect 9910 10168 9944 10744
rect 10928 10168 10962 10744
rect 13530 10534 13564 11110
rect 14548 10534 14582 11110
rect 15566 10534 15600 11110
rect 16584 10534 16618 11110
rect 17602 10534 17636 11110
rect 18620 10534 18654 11110
rect 19638 10534 19672 11110
rect 20656 10534 20690 11110
rect 21674 10534 21708 11110
rect 22692 10534 22726 11110
rect 23710 10534 23744 11110
rect 24728 10534 24762 11110
rect 25746 10534 25780 11110
rect 26764 10534 26798 11110
rect 27782 10534 27816 11110
rect 28800 10534 28834 11110
rect 29818 10534 29852 11110
rect 30836 10534 30870 11110
rect 31854 10534 31888 11110
rect 32872 10534 32906 11110
rect 33890 10534 33924 11110
rect 13824 10450 14288 10484
rect 14842 10450 15306 10484
rect 15860 10450 16324 10484
rect 16878 10450 17342 10484
rect 17896 10450 18360 10484
rect 18914 10450 19378 10484
rect 19932 10450 20396 10484
rect 20950 10450 21414 10484
rect 21968 10450 22432 10484
rect 22986 10450 23450 10484
rect 24004 10450 24468 10484
rect 25022 10450 25486 10484
rect 26040 10450 26504 10484
rect 27058 10450 27522 10484
rect 28076 10450 28540 10484
rect 29094 10450 29558 10484
rect 30112 10450 30576 10484
rect 31130 10450 31594 10484
rect 32148 10450 32612 10484
rect 33166 10450 33630 10484
rect 2060 10084 2524 10118
rect 3078 10084 3542 10118
rect 2060 9976 2524 10010
rect 4096 10084 4560 10118
rect 3078 9976 3542 10010
rect 5114 10084 5578 10118
rect 4096 9976 4560 10010
rect 6132 10084 6596 10118
rect 5114 9976 5578 10010
rect 7150 10084 7614 10118
rect 6132 9976 6596 10010
rect 8168 10084 8632 10118
rect 7150 9976 7614 10010
rect 9186 10084 9650 10118
rect 8168 9976 8632 10010
rect 10204 10084 10668 10118
rect 9186 9976 9650 10010
rect 10204 9976 10668 10010
rect 1766 9350 1800 9926
rect 2784 9350 2818 9926
rect 3802 9350 3836 9926
rect 4820 9350 4854 9926
rect 5838 9350 5872 9926
rect 6856 9350 6890 9926
rect 7874 9350 7908 9926
rect 8892 9350 8926 9926
rect 9910 9350 9944 9926
rect 13824 9926 14288 9960
rect 14842 9926 15306 9960
rect 15860 9926 16324 9960
rect 16878 9926 17342 9960
rect 17896 9926 18360 9960
rect 18914 9926 19378 9960
rect 19932 9926 20396 9960
rect 20950 9926 21414 9960
rect 21968 9926 22432 9960
rect 22986 9926 23450 9960
rect 24004 9926 24468 9960
rect 25022 9926 25486 9960
rect 26040 9926 26504 9960
rect 27058 9926 27522 9960
rect 28076 9926 28540 9960
rect 29094 9926 29558 9960
rect 30112 9926 30576 9960
rect 31130 9926 31594 9960
rect 32148 9926 32612 9960
rect 33166 9926 33630 9960
rect 10928 9350 10962 9926
rect 13530 9300 13564 9876
rect 2060 9266 2524 9300
rect 3078 9266 3542 9300
rect 2060 9158 2524 9192
rect 4096 9266 4560 9300
rect 3078 9158 3542 9192
rect 5114 9266 5578 9300
rect 4096 9158 4560 9192
rect 6132 9266 6596 9300
rect 5114 9158 5578 9192
rect 7150 9266 7614 9300
rect 6132 9158 6596 9192
rect 8168 9266 8632 9300
rect 7150 9158 7614 9192
rect 9186 9266 9650 9300
rect 8168 9158 8632 9192
rect 10204 9266 10668 9300
rect 14548 9300 14582 9876
rect 15566 9300 15600 9876
rect 16584 9300 16618 9876
rect 17602 9300 17636 9876
rect 18620 9300 18654 9876
rect 19638 9300 19672 9876
rect 20656 9300 20690 9876
rect 21674 9300 21708 9876
rect 22692 9300 22726 9876
rect 23710 9300 23744 9876
rect 24728 9300 24762 9876
rect 25746 9300 25780 9876
rect 26764 9300 26798 9876
rect 27782 9300 27816 9876
rect 28800 9300 28834 9876
rect 29818 9300 29852 9876
rect 30836 9300 30870 9876
rect 31854 9300 31888 9876
rect 32872 9300 32906 9876
rect 33890 9300 33924 9876
rect 9186 9158 9650 9192
rect 13824 9216 14288 9250
rect 14842 9216 15306 9250
rect 15860 9216 16324 9250
rect 16878 9216 17342 9250
rect 17896 9216 18360 9250
rect 18914 9216 19378 9250
rect 19932 9216 20396 9250
rect 20950 9216 21414 9250
rect 21968 9216 22432 9250
rect 22986 9216 23450 9250
rect 24004 9216 24468 9250
rect 25022 9216 25486 9250
rect 26040 9216 26504 9250
rect 27058 9216 27522 9250
rect 28076 9216 28540 9250
rect 29094 9216 29558 9250
rect 30112 9216 30576 9250
rect 31130 9216 31594 9250
rect 32148 9216 32612 9250
rect 33166 9216 33630 9250
rect 10204 9158 10668 9192
rect 1766 8532 1800 9108
rect 2784 8532 2818 9108
rect 3802 8532 3836 9108
rect 4820 8532 4854 9108
rect 5838 8532 5872 9108
rect 6856 8532 6890 9108
rect 7874 8532 7908 9108
rect 8892 8532 8926 9108
rect 9910 8532 9944 9108
rect 10928 8532 10962 9108
rect 13824 8694 14288 8728
rect 14842 8694 15306 8728
rect 15860 8694 16324 8728
rect 16878 8694 17342 8728
rect 17896 8694 18360 8728
rect 18914 8694 19378 8728
rect 19932 8694 20396 8728
rect 20950 8694 21414 8728
rect 21968 8694 22432 8728
rect 22986 8694 23450 8728
rect 24004 8694 24468 8728
rect 25022 8694 25486 8728
rect 26040 8694 26504 8728
rect 27058 8694 27522 8728
rect 28076 8694 28540 8728
rect 29094 8694 29558 8728
rect 30112 8694 30576 8728
rect 31130 8694 31594 8728
rect 32148 8694 32612 8728
rect 33166 8694 33630 8728
rect 2060 8448 2524 8482
rect 3078 8448 3542 8482
rect 2060 8340 2524 8374
rect 4096 8448 4560 8482
rect 3078 8340 3542 8374
rect 5114 8448 5578 8482
rect 4096 8340 4560 8374
rect 6132 8448 6596 8482
rect 5114 8340 5578 8374
rect 7150 8448 7614 8482
rect 6132 8340 6596 8374
rect 8168 8448 8632 8482
rect 7150 8340 7614 8374
rect 9186 8448 9650 8482
rect 8168 8340 8632 8374
rect 10204 8448 10668 8482
rect 9186 8340 9650 8374
rect 10204 8340 10668 8374
rect 1766 7714 1800 8290
rect 2784 7714 2818 8290
rect 3802 7714 3836 8290
rect 4820 7714 4854 8290
rect 5838 7714 5872 8290
rect 6856 7714 6890 8290
rect 7874 7714 7908 8290
rect 8892 7714 8926 8290
rect 9910 7714 9944 8290
rect 10928 7714 10962 8290
rect 13530 8068 13564 8644
rect 14548 8068 14582 8644
rect 15566 8068 15600 8644
rect 16584 8068 16618 8644
rect 17602 8068 17636 8644
rect 18620 8068 18654 8644
rect 19638 8068 19672 8644
rect 20656 8068 20690 8644
rect 21674 8068 21708 8644
rect 22692 8068 22726 8644
rect 23710 8068 23744 8644
rect 24728 8068 24762 8644
rect 25746 8068 25780 8644
rect 26764 8068 26798 8644
rect 27782 8068 27816 8644
rect 28800 8068 28834 8644
rect 29818 8068 29852 8644
rect 30836 8068 30870 8644
rect 31854 8068 31888 8644
rect 32872 8068 32906 8644
rect 33890 8068 33924 8644
rect 13824 7984 14288 8018
rect 14842 7984 15306 8018
rect 15860 7984 16324 8018
rect 16878 7984 17342 8018
rect 17896 7984 18360 8018
rect 18914 7984 19378 8018
rect 19932 7984 20396 8018
rect 20950 7984 21414 8018
rect 21968 7984 22432 8018
rect 22986 7984 23450 8018
rect 24004 7984 24468 8018
rect 25022 7984 25486 8018
rect 26040 7984 26504 8018
rect 27058 7984 27522 8018
rect 28076 7984 28540 8018
rect 29094 7984 29558 8018
rect 30112 7984 30576 8018
rect 31130 7984 31594 8018
rect 32148 7984 32612 8018
rect 33166 7984 33630 8018
rect 2060 7630 2524 7664
rect 3078 7630 3542 7664
rect 4096 7630 4560 7664
rect 5114 7630 5578 7664
rect 6132 7630 6596 7664
rect 7150 7630 7614 7664
rect 8168 7630 8632 7664
rect 9186 7630 9650 7664
rect 10204 7630 10668 7664
rect 13824 7460 14288 7494
rect 14842 7460 15306 7494
rect 15860 7460 16324 7494
rect 16878 7460 17342 7494
rect 17896 7460 18360 7494
rect 18914 7460 19378 7494
rect 19932 7460 20396 7494
rect 20950 7460 21414 7494
rect 21968 7460 22432 7494
rect 22986 7460 23450 7494
rect 24004 7460 24468 7494
rect 25022 7460 25486 7494
rect 26040 7460 26504 7494
rect 27058 7460 27522 7494
rect 28076 7460 28540 7494
rect 29094 7460 29558 7494
rect 30112 7460 30576 7494
rect 31130 7460 31594 7494
rect 32148 7460 32612 7494
rect 33166 7460 33630 7494
rect 8720 6956 8784 6990
rect 8938 6956 9002 6990
rect 9156 6956 9220 6990
rect 9374 6956 9438 6990
rect 9592 6956 9656 6990
rect 9810 6956 9874 6990
rect 10028 6956 10092 6990
rect 10246 6956 10310 6990
rect 10464 6956 10528 6990
rect 10682 6956 10746 6990
rect 8626 6730 8660 6906
rect 8844 6730 8878 6906
rect 9062 6730 9096 6906
rect 9280 6730 9314 6906
rect 9498 6730 9532 6906
rect 9716 6730 9750 6906
rect 9934 6730 9968 6906
rect 10152 6730 10186 6906
rect 10370 6730 10404 6906
rect 10588 6730 10622 6906
rect 10806 6730 10840 6906
rect 13530 6834 13564 7410
rect 14548 6834 14582 7410
rect 15566 6834 15600 7410
rect 16584 6834 16618 7410
rect 17602 6834 17636 7410
rect 18620 6834 18654 7410
rect 19638 6834 19672 7410
rect 20656 6834 20690 7410
rect 21674 6834 21708 7410
rect 22692 6834 22726 7410
rect 23710 6834 23744 7410
rect 24728 6834 24762 7410
rect 25746 6834 25780 7410
rect 26764 6834 26798 7410
rect 27782 6834 27816 7410
rect 28800 6834 28834 7410
rect 29818 6834 29852 7410
rect 30836 6834 30870 7410
rect 31854 6834 31888 7410
rect 32872 6834 32906 7410
rect 33890 6834 33924 7410
rect 13824 6750 14288 6784
rect 14842 6750 15306 6784
rect 15860 6750 16324 6784
rect 16878 6750 17342 6784
rect 17896 6750 18360 6784
rect 18914 6750 19378 6784
rect 19932 6750 20396 6784
rect 20950 6750 21414 6784
rect 21968 6750 22432 6784
rect 22986 6750 23450 6784
rect 24004 6750 24468 6784
rect 25022 6750 25486 6784
rect 26040 6750 26504 6784
rect 27058 6750 27522 6784
rect 28076 6750 28540 6784
rect 29094 6750 29558 6784
rect 30112 6750 30576 6784
rect 31130 6750 31594 6784
rect 32148 6750 32612 6784
rect 33166 6750 33630 6784
rect 8720 6646 8784 6680
rect 8938 6646 9002 6680
rect 9156 6646 9220 6680
rect 9374 6646 9438 6680
rect 9592 6646 9656 6680
rect 9810 6646 9874 6680
rect 10028 6646 10092 6680
rect 10246 6646 10310 6680
rect 10464 6646 10528 6680
rect 10682 6646 10746 6680
rect 13824 6226 14288 6260
rect 14842 6226 15306 6260
rect 15860 6226 16324 6260
rect 16878 6226 17342 6260
rect 17896 6226 18360 6260
rect 18914 6226 19378 6260
rect 19932 6226 20396 6260
rect 20950 6226 21414 6260
rect 21968 6226 22432 6260
rect 22986 6226 23450 6260
rect 24004 6226 24468 6260
rect 25022 6226 25486 6260
rect 26040 6226 26504 6260
rect 27058 6226 27522 6260
rect 28076 6226 28540 6260
rect 29094 6226 29558 6260
rect 30112 6226 30576 6260
rect 31130 6226 31594 6260
rect 32148 6226 32612 6260
rect 33166 6226 33630 6260
rect 8720 6124 8784 6158
rect 8938 6124 9002 6158
rect 9156 6124 9220 6158
rect 9374 6124 9438 6158
rect 9592 6124 9656 6158
rect 9810 6124 9874 6158
rect 10028 6124 10092 6158
rect 10246 6124 10310 6158
rect 10464 6124 10528 6158
rect 10682 6124 10746 6158
rect 8626 5898 8660 6074
rect 8844 5898 8878 6074
rect 9062 5898 9096 6074
rect 9280 5898 9314 6074
rect 9498 5898 9532 6074
rect 9716 5898 9750 6074
rect 9934 5898 9968 6074
rect 10152 5898 10186 6074
rect 10370 5898 10404 6074
rect 10588 5898 10622 6074
rect 10806 5898 10840 6074
rect 8720 5814 8784 5848
rect 8938 5814 9002 5848
rect 9156 5814 9220 5848
rect 9374 5814 9438 5848
rect 9592 5814 9656 5848
rect 9810 5814 9874 5848
rect 10028 5814 10092 5848
rect 10246 5814 10310 5848
rect 10464 5814 10528 5848
rect 10682 5814 10746 5848
rect 13530 5600 13564 6176
rect 14548 5600 14582 6176
rect 15566 5600 15600 6176
rect 16584 5600 16618 6176
rect 17602 5600 17636 6176
rect 18620 5600 18654 6176
rect 19638 5600 19672 6176
rect 20656 5600 20690 6176
rect 21674 5600 21708 6176
rect 22692 5600 22726 6176
rect 23710 5600 23744 6176
rect 24728 5600 24762 6176
rect 25746 5600 25780 6176
rect 26764 5600 26798 6176
rect 27782 5600 27816 6176
rect 28800 5600 28834 6176
rect 29818 5600 29852 6176
rect 30836 5600 30870 6176
rect 31854 5600 31888 6176
rect 32872 5600 32906 6176
rect 33890 5600 33924 6176
rect 13824 5516 14288 5550
rect 14842 5516 15306 5550
rect 15860 5516 16324 5550
rect 16878 5516 17342 5550
rect 17896 5516 18360 5550
rect 18914 5516 19378 5550
rect 19932 5516 20396 5550
rect 20950 5516 21414 5550
rect 21968 5516 22432 5550
rect 22986 5516 23450 5550
rect 24004 5516 24468 5550
rect 25022 5516 25486 5550
rect 26040 5516 26504 5550
rect 27058 5516 27522 5550
rect 28076 5516 28540 5550
rect 29094 5516 29558 5550
rect 30112 5516 30576 5550
rect 31130 5516 31594 5550
rect 32148 5516 32612 5550
rect 33166 5516 33630 5550
rect 13824 4994 14288 5028
rect 14842 4994 15306 5028
rect 15860 4994 16324 5028
rect 16878 4994 17342 5028
rect 17896 4994 18360 5028
rect 18914 4994 19378 5028
rect 19932 4994 20396 5028
rect 20950 4994 21414 5028
rect 21968 4994 22432 5028
rect 22986 4994 23450 5028
rect 24004 4994 24468 5028
rect 25022 4994 25486 5028
rect 26040 4994 26504 5028
rect 27058 4994 27522 5028
rect 28076 4994 28540 5028
rect 29094 4994 29558 5028
rect 30112 4994 30576 5028
rect 31130 4994 31594 5028
rect 32148 4994 32612 5028
rect 33166 4994 33630 5028
rect 1839 4797 2303 4831
rect 2857 4797 3321 4831
rect 3875 4797 4339 4831
rect 4893 4797 5357 4831
rect 5911 4797 6375 4831
rect 6929 4797 7393 4831
rect 8654 4798 8758 4832
rect 8952 4798 9056 4832
rect 9250 4798 9354 4832
rect 9548 4798 9652 4832
rect 9846 4798 9950 4832
rect 10144 4798 10248 4832
rect 10442 4798 10546 4832
rect 10740 4798 10844 4832
rect 11038 4798 11142 4832
rect 11336 4798 11440 4832
rect 11634 4798 11738 4832
rect 1545 4171 1579 4747
rect 2563 4171 2597 4747
rect 3581 4171 3615 4747
rect 4599 4171 4633 4747
rect 5617 4171 5651 4747
rect 6635 4171 6669 4747
rect 7653 4171 7687 4747
rect 8540 4172 8574 4748
rect 8838 4172 8872 4748
rect 9136 4172 9170 4748
rect 9434 4172 9468 4748
rect 9732 4172 9766 4748
rect 10030 4172 10064 4748
rect 10328 4172 10362 4748
rect 10626 4172 10660 4748
rect 10924 4172 10958 4748
rect 11222 4172 11256 4748
rect 11520 4172 11554 4748
rect 11818 4172 11852 4748
rect 13530 4368 13564 4944
rect 14548 4368 14582 4944
rect 15566 4368 15600 4944
rect 16584 4368 16618 4944
rect 17602 4368 17636 4944
rect 18620 4368 18654 4944
rect 19638 4368 19672 4944
rect 20656 4368 20690 4944
rect 21674 4368 21708 4944
rect 22692 4368 22726 4944
rect 23710 4368 23744 4944
rect 24728 4368 24762 4944
rect 25746 4368 25780 4944
rect 26764 4368 26798 4944
rect 27782 4368 27816 4944
rect 28800 4368 28834 4944
rect 29818 4368 29852 4944
rect 30836 4368 30870 4944
rect 31854 4368 31888 4944
rect 32872 4368 32906 4944
rect 33890 4368 33924 4944
rect 13824 4284 14288 4318
rect 14842 4284 15306 4318
rect 15860 4284 16324 4318
rect 16878 4284 17342 4318
rect 17896 4284 18360 4318
rect 18914 4284 19378 4318
rect 19932 4284 20396 4318
rect 20950 4284 21414 4318
rect 21968 4284 22432 4318
rect 22986 4284 23450 4318
rect 24004 4284 24468 4318
rect 25022 4284 25486 4318
rect 26040 4284 26504 4318
rect 27058 4284 27522 4318
rect 28076 4284 28540 4318
rect 29094 4284 29558 4318
rect 30112 4284 30576 4318
rect 31130 4284 31594 4318
rect 32148 4284 32612 4318
rect 33166 4284 33630 4318
rect 1839 4087 2303 4121
rect 2857 4087 3321 4121
rect 3875 4087 4339 4121
rect 4893 4087 5357 4121
rect 5911 4087 6375 4121
rect 6929 4087 7393 4121
rect 8654 4088 8758 4122
rect 8952 4088 9056 4122
rect 9250 4088 9354 4122
rect 9548 4088 9652 4122
rect 9846 4088 9950 4122
rect 10144 4088 10248 4122
rect 10442 4088 10546 4122
rect 10740 4088 10844 4122
rect 11038 4088 11142 4122
rect 11336 4088 11440 4122
rect 11634 4088 11738 4122
rect 13824 3760 14288 3794
rect 14842 3760 15306 3794
rect 15860 3760 16324 3794
rect 16878 3760 17342 3794
rect 17896 3760 18360 3794
rect 18914 3760 19378 3794
rect 19932 3760 20396 3794
rect 20950 3760 21414 3794
rect 21968 3760 22432 3794
rect 22986 3760 23450 3794
rect 24004 3760 24468 3794
rect 25022 3760 25486 3794
rect 26040 3760 26504 3794
rect 27058 3760 27522 3794
rect 28076 3760 28540 3794
rect 29094 3760 29558 3794
rect 30112 3760 30576 3794
rect 31130 3760 31594 3794
rect 32148 3760 32612 3794
rect 33166 3760 33630 3794
rect 1838 3684 2302 3718
rect 2856 3684 3320 3718
rect 3874 3684 4338 3718
rect 4892 3684 5356 3718
rect 5910 3684 6374 3718
rect 6928 3684 7392 3718
rect 8654 3686 8758 3720
rect 8952 3686 9056 3720
rect 9250 3686 9354 3720
rect 9548 3686 9652 3720
rect 9846 3686 9950 3720
rect 10144 3686 10248 3720
rect 10442 3686 10546 3720
rect 10740 3686 10844 3720
rect 11038 3686 11142 3720
rect 11336 3686 11440 3720
rect 11634 3686 11738 3720
rect 1544 3058 1578 3634
rect 2562 3058 2596 3634
rect 3580 3058 3614 3634
rect 4598 3058 4632 3634
rect 5616 3058 5650 3634
rect 6634 3058 6668 3634
rect 7652 3058 7686 3634
rect 8540 3060 8574 3636
rect 8838 3060 8872 3636
rect 9136 3060 9170 3636
rect 9434 3060 9468 3636
rect 9732 3060 9766 3636
rect 10030 3060 10064 3636
rect 10328 3060 10362 3636
rect 10626 3060 10660 3636
rect 10924 3060 10958 3636
rect 11222 3060 11256 3636
rect 11520 3060 11554 3636
rect 11818 3060 11852 3636
rect 13530 3134 13564 3710
rect 14548 3134 14582 3710
rect 15566 3134 15600 3710
rect 16584 3134 16618 3710
rect 17602 3134 17636 3710
rect 18620 3134 18654 3710
rect 19638 3134 19672 3710
rect 20656 3134 20690 3710
rect 21674 3134 21708 3710
rect 22692 3134 22726 3710
rect 23710 3134 23744 3710
rect 24728 3134 24762 3710
rect 25746 3134 25780 3710
rect 26764 3134 26798 3710
rect 27782 3134 27816 3710
rect 28800 3134 28834 3710
rect 29818 3134 29852 3710
rect 30836 3134 30870 3710
rect 31854 3134 31888 3710
rect 32872 3134 32906 3710
rect 33890 3134 33924 3710
rect 13824 3050 14288 3084
rect 14842 3050 15306 3084
rect 15860 3050 16324 3084
rect 16878 3050 17342 3084
rect 17896 3050 18360 3084
rect 18914 3050 19378 3084
rect 19932 3050 20396 3084
rect 20950 3050 21414 3084
rect 21968 3050 22432 3084
rect 22986 3050 23450 3084
rect 24004 3050 24468 3084
rect 25022 3050 25486 3084
rect 26040 3050 26504 3084
rect 27058 3050 27522 3084
rect 28076 3050 28540 3084
rect 29094 3050 29558 3084
rect 30112 3050 30576 3084
rect 31130 3050 31594 3084
rect 32148 3050 32612 3084
rect 33166 3050 33630 3084
rect 1838 2974 2302 3008
rect 2856 2974 3320 3008
rect 3874 2974 4338 3008
rect 4892 2974 5356 3008
rect 5910 2974 6374 3008
rect 6928 2974 7392 3008
rect 8654 2976 8758 3010
rect 8952 2976 9056 3010
rect 9250 2976 9354 3010
rect 9548 2976 9652 3010
rect 9846 2976 9950 3010
rect 10144 2976 10248 3010
rect 10442 2976 10546 3010
rect 10740 2976 10844 3010
rect 11038 2976 11142 3010
rect 11336 2976 11440 3010
rect 11634 2976 11738 3010
rect 1839 2573 2303 2607
rect 2857 2573 3321 2607
rect 3875 2573 4339 2607
rect 4893 2573 5357 2607
rect 5911 2573 6375 2607
rect 6929 2573 7393 2607
rect 8652 2574 8756 2608
rect 8950 2574 9054 2608
rect 9248 2574 9352 2608
rect 9546 2574 9650 2608
rect 9844 2574 9948 2608
rect 10142 2574 10246 2608
rect 10440 2574 10544 2608
rect 10738 2574 10842 2608
rect 11036 2574 11140 2608
rect 11334 2574 11438 2608
rect 11632 2574 11736 2608
rect 1545 1947 1579 2523
rect 2563 1947 2597 2523
rect 3581 1947 3615 2523
rect 4599 1947 4633 2523
rect 5617 1947 5651 2523
rect 6635 1947 6669 2523
rect 7653 1947 7687 2523
rect 8538 1948 8572 2524
rect 8836 1948 8870 2524
rect 9134 1948 9168 2524
rect 9432 1948 9466 2524
rect 9730 1948 9764 2524
rect 10028 1948 10062 2524
rect 10326 1948 10360 2524
rect 10624 1948 10658 2524
rect 10922 1948 10956 2524
rect 11220 1948 11254 2524
rect 11518 1948 11552 2524
rect 13824 2526 14288 2560
rect 14842 2526 15306 2560
rect 15860 2526 16324 2560
rect 16878 2526 17342 2560
rect 17896 2526 18360 2560
rect 18914 2526 19378 2560
rect 19932 2526 20396 2560
rect 20950 2526 21414 2560
rect 21968 2526 22432 2560
rect 22986 2526 23450 2560
rect 24004 2526 24468 2560
rect 25022 2526 25486 2560
rect 26040 2526 26504 2560
rect 27058 2526 27522 2560
rect 28076 2526 28540 2560
rect 29094 2526 29558 2560
rect 30112 2526 30576 2560
rect 31130 2526 31594 2560
rect 32148 2526 32612 2560
rect 33166 2526 33630 2560
rect 11816 1948 11850 2524
rect 13530 1900 13564 2476
rect 1839 1863 2303 1897
rect 2857 1863 3321 1897
rect 3875 1863 4339 1897
rect 4893 1863 5357 1897
rect 5911 1863 6375 1897
rect 6929 1863 7393 1897
rect 8652 1864 8756 1898
rect 8950 1864 9054 1898
rect 9248 1864 9352 1898
rect 9546 1864 9650 1898
rect 9844 1864 9948 1898
rect 10142 1864 10246 1898
rect 10440 1864 10544 1898
rect 10738 1864 10842 1898
rect 11036 1864 11140 1898
rect 11334 1864 11438 1898
rect 11632 1864 11736 1898
rect 14548 1900 14582 2476
rect 15566 1900 15600 2476
rect 16584 1900 16618 2476
rect 17602 1900 17636 2476
rect 18620 1900 18654 2476
rect 19638 1900 19672 2476
rect 20656 1900 20690 2476
rect 21674 1900 21708 2476
rect 22692 1900 22726 2476
rect 23710 1900 23744 2476
rect 24728 1900 24762 2476
rect 25746 1900 25780 2476
rect 26764 1900 26798 2476
rect 27782 1900 27816 2476
rect 28800 1900 28834 2476
rect 29818 1900 29852 2476
rect 30836 1900 30870 2476
rect 31854 1900 31888 2476
rect 32872 1900 32906 2476
rect 33890 1900 33924 2476
rect 13824 1816 14288 1850
rect 14842 1816 15306 1850
rect 15860 1816 16324 1850
rect 16878 1816 17342 1850
rect 17896 1816 18360 1850
rect 18914 1816 19378 1850
rect 19932 1816 20396 1850
rect 20950 1816 21414 1850
rect 21968 1816 22432 1850
rect 22986 1816 23450 1850
rect 24004 1816 24468 1850
rect 25022 1816 25486 1850
rect 26040 1816 26504 1850
rect 27058 1816 27522 1850
rect 28076 1816 28540 1850
rect 29094 1816 29558 1850
rect 30112 1816 30576 1850
rect 31130 1816 31594 1850
rect 32148 1816 32612 1850
rect 33166 1816 33630 1850
rect 1838 1460 2302 1494
rect 2856 1460 3320 1494
rect 3874 1460 4338 1494
rect 4892 1460 5356 1494
rect 5910 1460 6374 1494
rect 6928 1460 7392 1494
rect 8652 1464 8756 1498
rect 8950 1464 9054 1498
rect 9248 1464 9352 1498
rect 9546 1464 9650 1498
rect 9844 1464 9948 1498
rect 10142 1464 10246 1498
rect 10440 1464 10544 1498
rect 10738 1464 10842 1498
rect 11036 1464 11140 1498
rect 11334 1464 11438 1498
rect 11632 1464 11736 1498
rect 1544 834 1578 1410
rect 2562 834 2596 1410
rect 3580 834 3614 1410
rect 4598 834 4632 1410
rect 5616 834 5650 1410
rect 6634 834 6668 1410
rect 7652 834 7686 1410
rect 8538 838 8572 1414
rect 8836 838 8870 1414
rect 9134 838 9168 1414
rect 9432 838 9466 1414
rect 9730 838 9764 1414
rect 10028 838 10062 1414
rect 10326 838 10360 1414
rect 10624 838 10658 1414
rect 10922 838 10956 1414
rect 11220 838 11254 1414
rect 11518 838 11552 1414
rect 11816 838 11850 1414
rect 13824 1294 14288 1328
rect 14842 1294 15306 1328
rect 15860 1294 16324 1328
rect 16878 1294 17342 1328
rect 17896 1294 18360 1328
rect 18914 1294 19378 1328
rect 19932 1294 20396 1328
rect 20950 1294 21414 1328
rect 21968 1294 22432 1328
rect 22986 1294 23450 1328
rect 24004 1294 24468 1328
rect 25022 1294 25486 1328
rect 26040 1294 26504 1328
rect 27058 1294 27522 1328
rect 28076 1294 28540 1328
rect 29094 1294 29558 1328
rect 30112 1294 30576 1328
rect 31130 1294 31594 1328
rect 32148 1294 32612 1328
rect 33166 1294 33630 1328
rect 1838 750 2302 784
rect 2856 750 3320 784
rect 3874 750 4338 784
rect 4892 750 5356 784
rect 5910 750 6374 784
rect 6928 750 7392 784
rect 8652 754 8756 788
rect 8950 754 9054 788
rect 9248 754 9352 788
rect 9546 754 9650 788
rect 9844 754 9948 788
rect 10142 754 10246 788
rect 10440 754 10544 788
rect 10738 754 10842 788
rect 11036 754 11140 788
rect 11334 754 11438 788
rect 11632 754 11736 788
rect 13530 668 13564 1244
rect 14548 668 14582 1244
rect 15566 668 15600 1244
rect 16584 668 16618 1244
rect 17602 668 17636 1244
rect 18620 668 18654 1244
rect 19638 668 19672 1244
rect 20656 668 20690 1244
rect 21674 668 21708 1244
rect 22692 668 22726 1244
rect 23710 668 23744 1244
rect 24728 668 24762 1244
rect 25746 668 25780 1244
rect 26764 668 26798 1244
rect 27782 668 27816 1244
rect 28800 668 28834 1244
rect 29818 668 29852 1244
rect 30836 668 30870 1244
rect 31854 668 31888 1244
rect 32872 668 32906 1244
rect 33890 668 33924 1244
rect 13824 584 14288 618
rect 14842 584 15306 618
rect 15860 584 16324 618
rect 16878 584 17342 618
rect 17896 584 18360 618
rect 18914 584 19378 618
rect 19932 584 20396 618
rect 20950 584 21414 618
rect 21968 584 22432 618
rect 22986 584 23450 618
rect 24004 584 24468 618
rect 25022 584 25486 618
rect 26040 584 26504 618
rect 27058 584 27522 618
rect 28076 584 28540 618
rect 29094 584 29558 618
rect 30112 584 30576 618
rect 31130 584 31594 618
rect 32148 584 32612 618
rect 33166 584 33630 618
rect 35772 210 35872 14470
rect 52728 15262 52790 15362
rect 52790 15262 89710 15362
rect 89710 15262 89772 15362
rect 67826 14860 68290 14894
rect 68844 14860 69308 14894
rect 69862 14860 70326 14894
rect 70880 14860 71344 14894
rect 71898 14860 72362 14894
rect 72916 14860 73380 14894
rect 73934 14860 74398 14894
rect 74952 14860 75416 14894
rect 75970 14860 76434 14894
rect 76988 14860 77452 14894
rect 78006 14860 78470 14894
rect 79024 14860 79488 14894
rect 80042 14860 80506 14894
rect 81060 14860 81524 14894
rect 82078 14860 82542 14894
rect 83096 14860 83560 14894
rect 84114 14860 84578 14894
rect 85132 14860 85596 14894
rect 86150 14860 86614 14894
rect 87168 14860 87632 14894
rect 48736 8447 48956 8448
rect 50228 8447 50430 8448
rect 48736 8414 48786 8447
rect 48786 8414 48956 8447
rect 50228 8414 50404 8447
rect 50404 8414 50430 8447
rect 50464 8351 50500 8352
rect 48688 7778 48690 8350
rect 48690 7778 48724 8350
rect 48724 7778 48726 8350
rect 48908 8311 48992 8345
rect 49166 8311 49250 8345
rect 49424 8311 49508 8345
rect 49682 8311 49766 8345
rect 49940 8311 50024 8345
rect 50198 8311 50282 8345
rect 48804 7876 48838 8252
rect 49062 7876 49096 8252
rect 49320 7876 49354 8252
rect 49578 7876 49612 8252
rect 49836 7876 49870 8252
rect 50094 7876 50128 8252
rect 50352 7876 50386 8252
rect 48908 7783 48992 7817
rect 49166 7783 49250 7817
rect 49424 7783 49508 7817
rect 49682 7783 49766 7817
rect 49940 7783 50024 7817
rect 50198 7783 50282 7817
rect 50464 7777 50466 8351
rect 50466 7777 50500 8351
rect 50603 7911 50637 7945
rect 50695 7911 50729 7945
rect 50787 7911 50821 7945
rect 50464 7776 50500 7777
rect 50228 7715 50430 7716
rect 48736 7681 48786 7714
rect 48786 7681 48956 7714
rect 50228 7682 50404 7715
rect 50404 7682 50430 7715
rect 48736 7680 48956 7681
rect 50633 7574 50681 7622
rect 50737 7633 50783 7644
rect 50737 7604 50770 7633
rect 50770 7604 50783 7633
rect 48760 7514 48968 7516
rect 50232 7514 50430 7518
rect 48760 7480 48786 7514
rect 48786 7480 48968 7514
rect 50232 7480 50404 7514
rect 50404 7480 50430 7514
rect 48760 7478 48968 7480
rect 48688 7062 48690 7418
rect 48690 7062 48724 7418
rect 48908 7378 48992 7412
rect 49166 7378 49250 7412
rect 49424 7378 49508 7412
rect 49682 7378 49766 7412
rect 49940 7378 50024 7412
rect 50198 7378 50282 7412
rect 48804 7152 48838 7328
rect 49062 7152 49096 7328
rect 49320 7152 49354 7328
rect 49578 7152 49612 7328
rect 49836 7152 49870 7328
rect 50094 7152 50128 7328
rect 50352 7152 50386 7328
rect 48908 7068 48992 7102
rect 49166 7068 49250 7102
rect 49424 7068 49508 7102
rect 49682 7068 49766 7102
rect 49940 7068 50024 7102
rect 50198 7068 50282 7102
rect 50464 7062 50466 7418
rect 50466 7062 50500 7418
rect 50500 7062 50502 7418
rect 50603 7367 50637 7401
rect 50695 7367 50729 7401
rect 50787 7367 50821 7401
rect 48758 7000 48966 7002
rect 48758 6966 48786 7000
rect 48786 6966 48966 7000
rect 50230 6966 50404 7000
rect 50404 6966 50432 7000
rect 50230 6964 50432 6966
rect 48736 6483 48956 6484
rect 50228 6483 50430 6484
rect 48736 6450 48786 6483
rect 48786 6450 48956 6483
rect 50228 6450 50404 6483
rect 50404 6450 50430 6483
rect 50464 6387 50500 6388
rect 48688 5814 48690 6386
rect 48690 5814 48724 6386
rect 48724 5814 48726 6386
rect 48908 6347 48992 6381
rect 49166 6347 49250 6381
rect 49424 6347 49508 6381
rect 49682 6347 49766 6381
rect 49940 6347 50024 6381
rect 50198 6347 50282 6381
rect 48804 5912 48838 6288
rect 49062 5912 49096 6288
rect 49320 5912 49354 6288
rect 49578 5912 49612 6288
rect 49836 5912 49870 6288
rect 50094 5912 50128 6288
rect 50352 5912 50386 6288
rect 48908 5819 48992 5853
rect 49166 5819 49250 5853
rect 49424 5819 49508 5853
rect 49682 5819 49766 5853
rect 49940 5819 50024 5853
rect 50198 5819 50282 5853
rect 50464 5813 50466 6387
rect 50466 5813 50500 6387
rect 50603 5947 50637 5981
rect 50695 5947 50729 5981
rect 50787 5947 50821 5981
rect 50464 5812 50500 5813
rect 50228 5751 50430 5752
rect 48736 5717 48786 5750
rect 48786 5717 48956 5750
rect 50228 5718 50404 5751
rect 50404 5718 50430 5751
rect 48736 5716 48956 5717
rect 50633 5610 50681 5658
rect 50737 5669 50783 5680
rect 50737 5640 50770 5669
rect 50770 5640 50783 5669
rect 48760 5550 48968 5552
rect 50232 5550 50430 5554
rect 48760 5516 48786 5550
rect 48786 5516 48968 5550
rect 50232 5516 50404 5550
rect 50404 5516 50430 5550
rect 48760 5514 48968 5516
rect 48688 5098 48690 5454
rect 48690 5098 48724 5454
rect 48908 5414 48992 5448
rect 49166 5414 49250 5448
rect 49424 5414 49508 5448
rect 49682 5414 49766 5448
rect 49940 5414 50024 5448
rect 50198 5414 50282 5448
rect 48804 5188 48838 5364
rect 49062 5188 49096 5364
rect 49320 5188 49354 5364
rect 49578 5188 49612 5364
rect 49836 5188 49870 5364
rect 50094 5188 50128 5364
rect 50352 5188 50386 5364
rect 48908 5104 48992 5138
rect 49166 5104 49250 5138
rect 49424 5104 49508 5138
rect 49682 5104 49766 5138
rect 49940 5104 50024 5138
rect 50198 5104 50282 5138
rect 50464 5098 50466 5454
rect 50466 5098 50500 5454
rect 50500 5098 50502 5454
rect 50603 5403 50637 5437
rect 50695 5403 50729 5437
rect 50787 5403 50821 5437
rect 48758 5036 48966 5038
rect 48758 5002 48786 5036
rect 48786 5002 48966 5036
rect 50230 5002 50404 5036
rect 50404 5002 50432 5036
rect 50230 5000 50432 5002
rect 48736 4483 48956 4484
rect 50228 4483 50430 4484
rect 48736 4450 48786 4483
rect 48786 4450 48956 4483
rect 50228 4450 50404 4483
rect 50404 4450 50430 4483
rect 50464 4387 50500 4388
rect 48688 3814 48690 4386
rect 48690 3814 48724 4386
rect 48724 3814 48726 4386
rect 48908 4347 48992 4381
rect 49166 4347 49250 4381
rect 49424 4347 49508 4381
rect 49682 4347 49766 4381
rect 49940 4347 50024 4381
rect 50198 4347 50282 4381
rect 48804 3912 48838 4288
rect 49062 3912 49096 4288
rect 49320 3912 49354 4288
rect 49578 3912 49612 4288
rect 49836 3912 49870 4288
rect 50094 3912 50128 4288
rect 50352 3912 50386 4288
rect 48908 3819 48992 3853
rect 49166 3819 49250 3853
rect 49424 3819 49508 3853
rect 49682 3819 49766 3853
rect 49940 3819 50024 3853
rect 50198 3819 50282 3853
rect 50464 3813 50466 4387
rect 50466 3813 50500 4387
rect 50603 3947 50637 3981
rect 50695 3947 50729 3981
rect 50787 3947 50821 3981
rect 50464 3812 50500 3813
rect 50228 3751 50430 3752
rect 48736 3717 48786 3750
rect 48786 3717 48956 3750
rect 50228 3718 50404 3751
rect 50404 3718 50430 3751
rect 48736 3716 48956 3717
rect 50633 3610 50681 3658
rect 50737 3669 50783 3680
rect 50737 3640 50770 3669
rect 50770 3640 50783 3669
rect 48760 3550 48968 3552
rect 50232 3550 50430 3554
rect 48760 3516 48786 3550
rect 48786 3516 48968 3550
rect 50232 3516 50404 3550
rect 50404 3516 50430 3550
rect 48760 3514 48968 3516
rect 48688 3098 48690 3454
rect 48690 3098 48724 3454
rect 48908 3414 48992 3448
rect 49166 3414 49250 3448
rect 49424 3414 49508 3448
rect 49682 3414 49766 3448
rect 49940 3414 50024 3448
rect 50198 3414 50282 3448
rect 48804 3188 48838 3364
rect 49062 3188 49096 3364
rect 49320 3188 49354 3364
rect 49578 3188 49612 3364
rect 49836 3188 49870 3364
rect 50094 3188 50128 3364
rect 50352 3188 50386 3364
rect 48908 3104 48992 3138
rect 49166 3104 49250 3138
rect 49424 3104 49508 3138
rect 49682 3104 49766 3138
rect 49940 3104 50024 3138
rect 50198 3104 50282 3138
rect 50464 3098 50466 3454
rect 50466 3098 50500 3454
rect 50500 3098 50502 3454
rect 50603 3403 50637 3437
rect 50695 3403 50729 3437
rect 50787 3403 50821 3437
rect 48758 3036 48966 3038
rect 48758 3002 48786 3036
rect 48786 3002 48966 3036
rect 50230 3002 50404 3036
rect 50404 3002 50432 3036
rect 50230 3000 50432 3002
rect 48736 2393 48956 2394
rect 50228 2393 50430 2394
rect 48736 2360 48786 2393
rect 48786 2360 48956 2393
rect 50228 2360 50404 2393
rect 50404 2360 50430 2393
rect 50464 2297 50500 2298
rect 48688 1724 48690 2296
rect 48690 1724 48724 2296
rect 48724 1724 48726 2296
rect 48908 2257 48992 2291
rect 49166 2257 49250 2291
rect 49424 2257 49508 2291
rect 49682 2257 49766 2291
rect 49940 2257 50024 2291
rect 50198 2257 50282 2291
rect 48804 1822 48838 2198
rect 49062 1822 49096 2198
rect 49320 1822 49354 2198
rect 49578 1822 49612 2198
rect 49836 1822 49870 2198
rect 50094 1822 50128 2198
rect 50352 1822 50386 2198
rect 48908 1729 48992 1763
rect 49166 1729 49250 1763
rect 49424 1729 49508 1763
rect 49682 1729 49766 1763
rect 49940 1729 50024 1763
rect 50198 1729 50282 1763
rect 50464 1723 50466 2297
rect 50466 1723 50500 2297
rect 50603 1857 50637 1891
rect 50695 1857 50729 1891
rect 50787 1857 50821 1891
rect 50464 1722 50500 1723
rect 50228 1661 50430 1662
rect 48736 1627 48786 1660
rect 48786 1627 48956 1660
rect 50228 1628 50404 1661
rect 50404 1628 50430 1661
rect 48736 1626 48956 1627
rect 50633 1520 50681 1568
rect 50737 1579 50783 1590
rect 50737 1550 50770 1579
rect 50770 1550 50783 1579
rect 48760 1460 48968 1462
rect 50232 1460 50430 1464
rect 48760 1426 48786 1460
rect 48786 1426 48968 1460
rect 50232 1426 50404 1460
rect 50404 1426 50430 1460
rect 48760 1424 48968 1426
rect 48688 1008 48690 1364
rect 48690 1008 48724 1364
rect 48908 1324 48992 1358
rect 49166 1324 49250 1358
rect 49424 1324 49508 1358
rect 49682 1324 49766 1358
rect 49940 1324 50024 1358
rect 50198 1324 50282 1358
rect 48804 1098 48838 1274
rect 49062 1098 49096 1274
rect 49320 1098 49354 1274
rect 49578 1098 49612 1274
rect 49836 1098 49870 1274
rect 50094 1098 50128 1274
rect 50352 1098 50386 1274
rect 48908 1014 48992 1048
rect 49166 1014 49250 1048
rect 49424 1014 49508 1048
rect 49682 1014 49766 1048
rect 49940 1014 50024 1048
rect 50198 1014 50282 1048
rect 50464 1008 50466 1364
rect 50466 1008 50500 1364
rect 50500 1008 50502 1364
rect 50603 1313 50637 1347
rect 50695 1313 50729 1347
rect 50787 1313 50821 1347
rect 48758 946 48966 948
rect 48758 912 48786 946
rect 48786 912 48966 946
rect 50230 912 50404 946
rect 50404 912 50432 946
rect 50230 910 50432 912
rect -1272 -682 -1210 -582
rect -1210 -682 35710 -582
rect 35710 -682 35772 -582
rect 52628 210 52728 14470
rect 67532 14234 67566 14810
rect 68550 14234 68584 14810
rect 69568 14234 69602 14810
rect 70586 14234 70620 14810
rect 71604 14234 71638 14810
rect 72622 14234 72656 14810
rect 73640 14234 73674 14810
rect 74658 14234 74692 14810
rect 75676 14234 75710 14810
rect 76694 14234 76728 14810
rect 77712 14234 77746 14810
rect 78730 14234 78764 14810
rect 79748 14234 79782 14810
rect 80766 14234 80800 14810
rect 81784 14234 81818 14810
rect 82802 14234 82836 14810
rect 83820 14234 83854 14810
rect 84838 14234 84872 14810
rect 85856 14234 85890 14810
rect 86874 14234 86908 14810
rect 87892 14234 87926 14810
rect 67826 14150 68290 14184
rect 68844 14150 69308 14184
rect 69862 14150 70326 14184
rect 70880 14150 71344 14184
rect 71898 14150 72362 14184
rect 72916 14150 73380 14184
rect 73934 14150 74398 14184
rect 74952 14150 75416 14184
rect 75970 14150 76434 14184
rect 76988 14150 77452 14184
rect 78006 14150 78470 14184
rect 79024 14150 79488 14184
rect 80042 14150 80506 14184
rect 81060 14150 81524 14184
rect 82078 14150 82542 14184
rect 83096 14150 83560 14184
rect 84114 14150 84578 14184
rect 85132 14150 85596 14184
rect 86150 14150 86614 14184
rect 87168 14150 87632 14184
rect 56060 14066 56524 14100
rect 57078 14066 57542 14100
rect 58096 14066 58560 14100
rect 59114 14066 59578 14100
rect 60132 14066 60596 14100
rect 61150 14066 61614 14100
rect 62168 14066 62632 14100
rect 63186 14066 63650 14100
rect 64204 14066 64668 14100
rect 55766 13440 55800 14016
rect 56784 13440 56818 14016
rect 57802 13440 57836 14016
rect 58820 13440 58854 14016
rect 59838 13440 59872 14016
rect 60856 13440 60890 14016
rect 61874 13440 61908 14016
rect 62892 13440 62926 14016
rect 63910 13440 63944 14016
rect 64928 13440 64962 14016
rect 67826 13626 68290 13660
rect 68844 13626 69308 13660
rect 69862 13626 70326 13660
rect 70880 13626 71344 13660
rect 71898 13626 72362 13660
rect 72916 13626 73380 13660
rect 73934 13626 74398 13660
rect 74952 13626 75416 13660
rect 75970 13626 76434 13660
rect 76988 13626 77452 13660
rect 78006 13626 78470 13660
rect 79024 13626 79488 13660
rect 80042 13626 80506 13660
rect 81060 13626 81524 13660
rect 82078 13626 82542 13660
rect 83096 13626 83560 13660
rect 84114 13626 84578 13660
rect 85132 13626 85596 13660
rect 86150 13626 86614 13660
rect 87168 13626 87632 13660
rect 56060 13356 56524 13390
rect 57078 13356 57542 13390
rect 56060 13248 56524 13282
rect 58096 13356 58560 13390
rect 57078 13248 57542 13282
rect 59114 13356 59578 13390
rect 58096 13248 58560 13282
rect 60132 13356 60596 13390
rect 59114 13248 59578 13282
rect 61150 13356 61614 13390
rect 60132 13248 60596 13282
rect 62168 13356 62632 13390
rect 61150 13248 61614 13282
rect 63186 13356 63650 13390
rect 62168 13248 62632 13282
rect 64204 13356 64668 13390
rect 63186 13248 63650 13282
rect 64204 13248 64668 13282
rect 55766 12622 55800 13198
rect 56784 12622 56818 13198
rect 57802 12622 57836 13198
rect 58820 12622 58854 13198
rect 59838 12622 59872 13198
rect 60856 12622 60890 13198
rect 61874 12622 61908 13198
rect 62892 12622 62926 13198
rect 63910 12622 63944 13198
rect 64928 12622 64962 13198
rect 67532 13000 67566 13576
rect 68550 13000 68584 13576
rect 69568 13000 69602 13576
rect 70586 13000 70620 13576
rect 71604 13000 71638 13576
rect 72622 13000 72656 13576
rect 73640 13000 73674 13576
rect 74658 13000 74692 13576
rect 75676 13000 75710 13576
rect 76694 13000 76728 13576
rect 77712 13000 77746 13576
rect 78730 13000 78764 13576
rect 79748 13000 79782 13576
rect 80766 13000 80800 13576
rect 81784 13000 81818 13576
rect 82802 13000 82836 13576
rect 83820 13000 83854 13576
rect 84838 13000 84872 13576
rect 85856 13000 85890 13576
rect 86874 13000 86908 13576
rect 87892 13000 87926 13576
rect 67826 12916 68290 12950
rect 68844 12916 69308 12950
rect 69862 12916 70326 12950
rect 70880 12916 71344 12950
rect 71898 12916 72362 12950
rect 72916 12916 73380 12950
rect 73934 12916 74398 12950
rect 74952 12916 75416 12950
rect 75970 12916 76434 12950
rect 76988 12916 77452 12950
rect 78006 12916 78470 12950
rect 79024 12916 79488 12950
rect 80042 12916 80506 12950
rect 81060 12916 81524 12950
rect 82078 12916 82542 12950
rect 83096 12916 83560 12950
rect 84114 12916 84578 12950
rect 85132 12916 85596 12950
rect 86150 12916 86614 12950
rect 87168 12916 87632 12950
rect 56060 12538 56524 12572
rect 57078 12538 57542 12572
rect 56060 12430 56524 12464
rect 58096 12538 58560 12572
rect 57078 12430 57542 12464
rect 59114 12538 59578 12572
rect 58096 12430 58560 12464
rect 60132 12538 60596 12572
rect 59114 12430 59578 12464
rect 61150 12538 61614 12572
rect 60132 12430 60596 12464
rect 62168 12538 62632 12572
rect 61150 12430 61614 12464
rect 63186 12538 63650 12572
rect 62168 12430 62632 12464
rect 64204 12538 64668 12572
rect 63186 12430 63650 12464
rect 64204 12430 64668 12464
rect 55766 11804 55800 12380
rect 56784 11804 56818 12380
rect 57802 11804 57836 12380
rect 58820 11804 58854 12380
rect 59838 11804 59872 12380
rect 60856 11804 60890 12380
rect 61874 11804 61908 12380
rect 62892 11804 62926 12380
rect 63910 11804 63944 12380
rect 67826 12394 68290 12428
rect 68844 12394 69308 12428
rect 69862 12394 70326 12428
rect 70880 12394 71344 12428
rect 71898 12394 72362 12428
rect 72916 12394 73380 12428
rect 73934 12394 74398 12428
rect 74952 12394 75416 12428
rect 75970 12394 76434 12428
rect 76988 12394 77452 12428
rect 78006 12394 78470 12428
rect 79024 12394 79488 12428
rect 80042 12394 80506 12428
rect 81060 12394 81524 12428
rect 82078 12394 82542 12428
rect 83096 12394 83560 12428
rect 84114 12394 84578 12428
rect 85132 12394 85596 12428
rect 86150 12394 86614 12428
rect 87168 12394 87632 12428
rect 64928 11804 64962 12380
rect 67532 11768 67566 12344
rect 56060 11720 56524 11754
rect 57078 11720 57542 11754
rect 56060 11612 56524 11646
rect 58096 11720 58560 11754
rect 57078 11612 57542 11646
rect 59114 11720 59578 11754
rect 58096 11612 58560 11646
rect 60132 11720 60596 11754
rect 59114 11612 59578 11646
rect 61150 11720 61614 11754
rect 60132 11612 60596 11646
rect 62168 11720 62632 11754
rect 61150 11612 61614 11646
rect 63186 11720 63650 11754
rect 62168 11612 62632 11646
rect 64204 11720 64668 11754
rect 68550 11768 68584 12344
rect 69568 11768 69602 12344
rect 70586 11768 70620 12344
rect 71604 11768 71638 12344
rect 72622 11768 72656 12344
rect 73640 11768 73674 12344
rect 74658 11768 74692 12344
rect 75676 11768 75710 12344
rect 76694 11768 76728 12344
rect 77712 11768 77746 12344
rect 78730 11768 78764 12344
rect 79748 11768 79782 12344
rect 80766 11768 80800 12344
rect 81784 11768 81818 12344
rect 82802 11768 82836 12344
rect 83820 11768 83854 12344
rect 84838 11768 84872 12344
rect 85856 11768 85890 12344
rect 86874 11768 86908 12344
rect 87892 11768 87926 12344
rect 63186 11612 63650 11646
rect 67826 11684 68290 11718
rect 68844 11684 69308 11718
rect 69862 11684 70326 11718
rect 70880 11684 71344 11718
rect 71898 11684 72362 11718
rect 72916 11684 73380 11718
rect 73934 11684 74398 11718
rect 74952 11684 75416 11718
rect 75970 11684 76434 11718
rect 76988 11684 77452 11718
rect 78006 11684 78470 11718
rect 79024 11684 79488 11718
rect 80042 11684 80506 11718
rect 81060 11684 81524 11718
rect 82078 11684 82542 11718
rect 83096 11684 83560 11718
rect 84114 11684 84578 11718
rect 85132 11684 85596 11718
rect 86150 11684 86614 11718
rect 87168 11684 87632 11718
rect 64204 11612 64668 11646
rect 55766 10986 55800 11562
rect 56784 10986 56818 11562
rect 57802 10986 57836 11562
rect 58820 10986 58854 11562
rect 59838 10986 59872 11562
rect 60856 10986 60890 11562
rect 61874 10986 61908 11562
rect 62892 10986 62926 11562
rect 63910 10986 63944 11562
rect 64928 10986 64962 11562
rect 67824 11160 68288 11194
rect 68842 11160 69306 11194
rect 69860 11160 70324 11194
rect 70878 11160 71342 11194
rect 71896 11160 72360 11194
rect 72914 11160 73378 11194
rect 73932 11160 74396 11194
rect 74950 11160 75414 11194
rect 75968 11160 76432 11194
rect 76986 11160 77450 11194
rect 78004 11160 78468 11194
rect 79022 11160 79486 11194
rect 80040 11160 80504 11194
rect 81058 11160 81522 11194
rect 82076 11160 82540 11194
rect 83094 11160 83558 11194
rect 84112 11160 84576 11194
rect 85130 11160 85594 11194
rect 86148 11160 86612 11194
rect 87166 11160 87630 11194
rect 56060 10902 56524 10936
rect 57078 10902 57542 10936
rect 56060 10794 56524 10828
rect 58096 10902 58560 10936
rect 57078 10794 57542 10828
rect 59114 10902 59578 10936
rect 58096 10794 58560 10828
rect 60132 10902 60596 10936
rect 59114 10794 59578 10828
rect 61150 10902 61614 10936
rect 60132 10794 60596 10828
rect 62168 10902 62632 10936
rect 61150 10794 61614 10828
rect 63186 10902 63650 10936
rect 62168 10794 62632 10828
rect 64204 10902 64668 10936
rect 63186 10794 63650 10828
rect 64204 10794 64668 10828
rect 55766 10168 55800 10744
rect 56784 10168 56818 10744
rect 57802 10168 57836 10744
rect 58820 10168 58854 10744
rect 59838 10168 59872 10744
rect 60856 10168 60890 10744
rect 61874 10168 61908 10744
rect 62892 10168 62926 10744
rect 63910 10168 63944 10744
rect 64928 10168 64962 10744
rect 67530 10534 67564 11110
rect 68548 10534 68582 11110
rect 69566 10534 69600 11110
rect 70584 10534 70618 11110
rect 71602 10534 71636 11110
rect 72620 10534 72654 11110
rect 73638 10534 73672 11110
rect 74656 10534 74690 11110
rect 75674 10534 75708 11110
rect 76692 10534 76726 11110
rect 77710 10534 77744 11110
rect 78728 10534 78762 11110
rect 79746 10534 79780 11110
rect 80764 10534 80798 11110
rect 81782 10534 81816 11110
rect 82800 10534 82834 11110
rect 83818 10534 83852 11110
rect 84836 10534 84870 11110
rect 85854 10534 85888 11110
rect 86872 10534 86906 11110
rect 87890 10534 87924 11110
rect 67824 10450 68288 10484
rect 68842 10450 69306 10484
rect 69860 10450 70324 10484
rect 70878 10450 71342 10484
rect 71896 10450 72360 10484
rect 72914 10450 73378 10484
rect 73932 10450 74396 10484
rect 74950 10450 75414 10484
rect 75968 10450 76432 10484
rect 76986 10450 77450 10484
rect 78004 10450 78468 10484
rect 79022 10450 79486 10484
rect 80040 10450 80504 10484
rect 81058 10450 81522 10484
rect 82076 10450 82540 10484
rect 83094 10450 83558 10484
rect 84112 10450 84576 10484
rect 85130 10450 85594 10484
rect 86148 10450 86612 10484
rect 87166 10450 87630 10484
rect 56060 10084 56524 10118
rect 57078 10084 57542 10118
rect 56060 9976 56524 10010
rect 58096 10084 58560 10118
rect 57078 9976 57542 10010
rect 59114 10084 59578 10118
rect 58096 9976 58560 10010
rect 60132 10084 60596 10118
rect 59114 9976 59578 10010
rect 61150 10084 61614 10118
rect 60132 9976 60596 10010
rect 62168 10084 62632 10118
rect 61150 9976 61614 10010
rect 63186 10084 63650 10118
rect 62168 9976 62632 10010
rect 64204 10084 64668 10118
rect 63186 9976 63650 10010
rect 64204 9976 64668 10010
rect 55766 9350 55800 9926
rect 56784 9350 56818 9926
rect 57802 9350 57836 9926
rect 58820 9350 58854 9926
rect 59838 9350 59872 9926
rect 60856 9350 60890 9926
rect 61874 9350 61908 9926
rect 62892 9350 62926 9926
rect 63910 9350 63944 9926
rect 67824 9926 68288 9960
rect 68842 9926 69306 9960
rect 69860 9926 70324 9960
rect 70878 9926 71342 9960
rect 71896 9926 72360 9960
rect 72914 9926 73378 9960
rect 73932 9926 74396 9960
rect 74950 9926 75414 9960
rect 75968 9926 76432 9960
rect 76986 9926 77450 9960
rect 78004 9926 78468 9960
rect 79022 9926 79486 9960
rect 80040 9926 80504 9960
rect 81058 9926 81522 9960
rect 82076 9926 82540 9960
rect 83094 9926 83558 9960
rect 84112 9926 84576 9960
rect 85130 9926 85594 9960
rect 86148 9926 86612 9960
rect 87166 9926 87630 9960
rect 64928 9350 64962 9926
rect 67530 9300 67564 9876
rect 56060 9266 56524 9300
rect 57078 9266 57542 9300
rect 56060 9158 56524 9192
rect 58096 9266 58560 9300
rect 57078 9158 57542 9192
rect 59114 9266 59578 9300
rect 58096 9158 58560 9192
rect 60132 9266 60596 9300
rect 59114 9158 59578 9192
rect 61150 9266 61614 9300
rect 60132 9158 60596 9192
rect 62168 9266 62632 9300
rect 61150 9158 61614 9192
rect 63186 9266 63650 9300
rect 62168 9158 62632 9192
rect 64204 9266 64668 9300
rect 68548 9300 68582 9876
rect 69566 9300 69600 9876
rect 70584 9300 70618 9876
rect 71602 9300 71636 9876
rect 72620 9300 72654 9876
rect 73638 9300 73672 9876
rect 74656 9300 74690 9876
rect 75674 9300 75708 9876
rect 76692 9300 76726 9876
rect 77710 9300 77744 9876
rect 78728 9300 78762 9876
rect 79746 9300 79780 9876
rect 80764 9300 80798 9876
rect 81782 9300 81816 9876
rect 82800 9300 82834 9876
rect 83818 9300 83852 9876
rect 84836 9300 84870 9876
rect 85854 9300 85888 9876
rect 86872 9300 86906 9876
rect 87890 9300 87924 9876
rect 63186 9158 63650 9192
rect 67824 9216 68288 9250
rect 68842 9216 69306 9250
rect 69860 9216 70324 9250
rect 70878 9216 71342 9250
rect 71896 9216 72360 9250
rect 72914 9216 73378 9250
rect 73932 9216 74396 9250
rect 74950 9216 75414 9250
rect 75968 9216 76432 9250
rect 76986 9216 77450 9250
rect 78004 9216 78468 9250
rect 79022 9216 79486 9250
rect 80040 9216 80504 9250
rect 81058 9216 81522 9250
rect 82076 9216 82540 9250
rect 83094 9216 83558 9250
rect 84112 9216 84576 9250
rect 85130 9216 85594 9250
rect 86148 9216 86612 9250
rect 87166 9216 87630 9250
rect 64204 9158 64668 9192
rect 55766 8532 55800 9108
rect 56784 8532 56818 9108
rect 57802 8532 57836 9108
rect 58820 8532 58854 9108
rect 59838 8532 59872 9108
rect 60856 8532 60890 9108
rect 61874 8532 61908 9108
rect 62892 8532 62926 9108
rect 63910 8532 63944 9108
rect 64928 8532 64962 9108
rect 67824 8694 68288 8728
rect 68842 8694 69306 8728
rect 69860 8694 70324 8728
rect 70878 8694 71342 8728
rect 71896 8694 72360 8728
rect 72914 8694 73378 8728
rect 73932 8694 74396 8728
rect 74950 8694 75414 8728
rect 75968 8694 76432 8728
rect 76986 8694 77450 8728
rect 78004 8694 78468 8728
rect 79022 8694 79486 8728
rect 80040 8694 80504 8728
rect 81058 8694 81522 8728
rect 82076 8694 82540 8728
rect 83094 8694 83558 8728
rect 84112 8694 84576 8728
rect 85130 8694 85594 8728
rect 86148 8694 86612 8728
rect 87166 8694 87630 8728
rect 56060 8448 56524 8482
rect 57078 8448 57542 8482
rect 56060 8340 56524 8374
rect 58096 8448 58560 8482
rect 57078 8340 57542 8374
rect 59114 8448 59578 8482
rect 58096 8340 58560 8374
rect 60132 8448 60596 8482
rect 59114 8340 59578 8374
rect 61150 8448 61614 8482
rect 60132 8340 60596 8374
rect 62168 8448 62632 8482
rect 61150 8340 61614 8374
rect 63186 8448 63650 8482
rect 62168 8340 62632 8374
rect 64204 8448 64668 8482
rect 63186 8340 63650 8374
rect 64204 8340 64668 8374
rect 55766 7714 55800 8290
rect 56784 7714 56818 8290
rect 57802 7714 57836 8290
rect 58820 7714 58854 8290
rect 59838 7714 59872 8290
rect 60856 7714 60890 8290
rect 61874 7714 61908 8290
rect 62892 7714 62926 8290
rect 63910 7714 63944 8290
rect 64928 7714 64962 8290
rect 67530 8068 67564 8644
rect 68548 8068 68582 8644
rect 69566 8068 69600 8644
rect 70584 8068 70618 8644
rect 71602 8068 71636 8644
rect 72620 8068 72654 8644
rect 73638 8068 73672 8644
rect 74656 8068 74690 8644
rect 75674 8068 75708 8644
rect 76692 8068 76726 8644
rect 77710 8068 77744 8644
rect 78728 8068 78762 8644
rect 79746 8068 79780 8644
rect 80764 8068 80798 8644
rect 81782 8068 81816 8644
rect 82800 8068 82834 8644
rect 83818 8068 83852 8644
rect 84836 8068 84870 8644
rect 85854 8068 85888 8644
rect 86872 8068 86906 8644
rect 87890 8068 87924 8644
rect 67824 7984 68288 8018
rect 68842 7984 69306 8018
rect 69860 7984 70324 8018
rect 70878 7984 71342 8018
rect 71896 7984 72360 8018
rect 72914 7984 73378 8018
rect 73932 7984 74396 8018
rect 74950 7984 75414 8018
rect 75968 7984 76432 8018
rect 76986 7984 77450 8018
rect 78004 7984 78468 8018
rect 79022 7984 79486 8018
rect 80040 7984 80504 8018
rect 81058 7984 81522 8018
rect 82076 7984 82540 8018
rect 83094 7984 83558 8018
rect 84112 7984 84576 8018
rect 85130 7984 85594 8018
rect 86148 7984 86612 8018
rect 87166 7984 87630 8018
rect 56060 7630 56524 7664
rect 57078 7630 57542 7664
rect 58096 7630 58560 7664
rect 59114 7630 59578 7664
rect 60132 7630 60596 7664
rect 61150 7630 61614 7664
rect 62168 7630 62632 7664
rect 63186 7630 63650 7664
rect 64204 7630 64668 7664
rect 67824 7460 68288 7494
rect 68842 7460 69306 7494
rect 69860 7460 70324 7494
rect 70878 7460 71342 7494
rect 71896 7460 72360 7494
rect 72914 7460 73378 7494
rect 73932 7460 74396 7494
rect 74950 7460 75414 7494
rect 75968 7460 76432 7494
rect 76986 7460 77450 7494
rect 78004 7460 78468 7494
rect 79022 7460 79486 7494
rect 80040 7460 80504 7494
rect 81058 7460 81522 7494
rect 82076 7460 82540 7494
rect 83094 7460 83558 7494
rect 84112 7460 84576 7494
rect 85130 7460 85594 7494
rect 86148 7460 86612 7494
rect 87166 7460 87630 7494
rect 62720 6956 62784 6990
rect 62938 6956 63002 6990
rect 63156 6956 63220 6990
rect 63374 6956 63438 6990
rect 63592 6956 63656 6990
rect 63810 6956 63874 6990
rect 64028 6956 64092 6990
rect 64246 6956 64310 6990
rect 64464 6956 64528 6990
rect 64682 6956 64746 6990
rect 62626 6730 62660 6906
rect 62844 6730 62878 6906
rect 63062 6730 63096 6906
rect 63280 6730 63314 6906
rect 63498 6730 63532 6906
rect 63716 6730 63750 6906
rect 63934 6730 63968 6906
rect 64152 6730 64186 6906
rect 64370 6730 64404 6906
rect 64588 6730 64622 6906
rect 64806 6730 64840 6906
rect 67530 6834 67564 7410
rect 68548 6834 68582 7410
rect 69566 6834 69600 7410
rect 70584 6834 70618 7410
rect 71602 6834 71636 7410
rect 72620 6834 72654 7410
rect 73638 6834 73672 7410
rect 74656 6834 74690 7410
rect 75674 6834 75708 7410
rect 76692 6834 76726 7410
rect 77710 6834 77744 7410
rect 78728 6834 78762 7410
rect 79746 6834 79780 7410
rect 80764 6834 80798 7410
rect 81782 6834 81816 7410
rect 82800 6834 82834 7410
rect 83818 6834 83852 7410
rect 84836 6834 84870 7410
rect 85854 6834 85888 7410
rect 86872 6834 86906 7410
rect 87890 6834 87924 7410
rect 67824 6750 68288 6784
rect 68842 6750 69306 6784
rect 69860 6750 70324 6784
rect 70878 6750 71342 6784
rect 71896 6750 72360 6784
rect 72914 6750 73378 6784
rect 73932 6750 74396 6784
rect 74950 6750 75414 6784
rect 75968 6750 76432 6784
rect 76986 6750 77450 6784
rect 78004 6750 78468 6784
rect 79022 6750 79486 6784
rect 80040 6750 80504 6784
rect 81058 6750 81522 6784
rect 82076 6750 82540 6784
rect 83094 6750 83558 6784
rect 84112 6750 84576 6784
rect 85130 6750 85594 6784
rect 86148 6750 86612 6784
rect 87166 6750 87630 6784
rect 62720 6646 62784 6680
rect 62938 6646 63002 6680
rect 63156 6646 63220 6680
rect 63374 6646 63438 6680
rect 63592 6646 63656 6680
rect 63810 6646 63874 6680
rect 64028 6646 64092 6680
rect 64246 6646 64310 6680
rect 64464 6646 64528 6680
rect 64682 6646 64746 6680
rect 67824 6226 68288 6260
rect 68842 6226 69306 6260
rect 69860 6226 70324 6260
rect 70878 6226 71342 6260
rect 71896 6226 72360 6260
rect 72914 6226 73378 6260
rect 73932 6226 74396 6260
rect 74950 6226 75414 6260
rect 75968 6226 76432 6260
rect 76986 6226 77450 6260
rect 78004 6226 78468 6260
rect 79022 6226 79486 6260
rect 80040 6226 80504 6260
rect 81058 6226 81522 6260
rect 82076 6226 82540 6260
rect 83094 6226 83558 6260
rect 84112 6226 84576 6260
rect 85130 6226 85594 6260
rect 86148 6226 86612 6260
rect 87166 6226 87630 6260
rect 62720 6124 62784 6158
rect 62938 6124 63002 6158
rect 63156 6124 63220 6158
rect 63374 6124 63438 6158
rect 63592 6124 63656 6158
rect 63810 6124 63874 6158
rect 64028 6124 64092 6158
rect 64246 6124 64310 6158
rect 64464 6124 64528 6158
rect 64682 6124 64746 6158
rect 62626 5898 62660 6074
rect 62844 5898 62878 6074
rect 63062 5898 63096 6074
rect 63280 5898 63314 6074
rect 63498 5898 63532 6074
rect 63716 5898 63750 6074
rect 63934 5898 63968 6074
rect 64152 5898 64186 6074
rect 64370 5898 64404 6074
rect 64588 5898 64622 6074
rect 64806 5898 64840 6074
rect 62720 5814 62784 5848
rect 62938 5814 63002 5848
rect 63156 5814 63220 5848
rect 63374 5814 63438 5848
rect 63592 5814 63656 5848
rect 63810 5814 63874 5848
rect 64028 5814 64092 5848
rect 64246 5814 64310 5848
rect 64464 5814 64528 5848
rect 64682 5814 64746 5848
rect 67530 5600 67564 6176
rect 68548 5600 68582 6176
rect 69566 5600 69600 6176
rect 70584 5600 70618 6176
rect 71602 5600 71636 6176
rect 72620 5600 72654 6176
rect 73638 5600 73672 6176
rect 74656 5600 74690 6176
rect 75674 5600 75708 6176
rect 76692 5600 76726 6176
rect 77710 5600 77744 6176
rect 78728 5600 78762 6176
rect 79746 5600 79780 6176
rect 80764 5600 80798 6176
rect 81782 5600 81816 6176
rect 82800 5600 82834 6176
rect 83818 5600 83852 6176
rect 84836 5600 84870 6176
rect 85854 5600 85888 6176
rect 86872 5600 86906 6176
rect 87890 5600 87924 6176
rect 67824 5516 68288 5550
rect 68842 5516 69306 5550
rect 69860 5516 70324 5550
rect 70878 5516 71342 5550
rect 71896 5516 72360 5550
rect 72914 5516 73378 5550
rect 73932 5516 74396 5550
rect 74950 5516 75414 5550
rect 75968 5516 76432 5550
rect 76986 5516 77450 5550
rect 78004 5516 78468 5550
rect 79022 5516 79486 5550
rect 80040 5516 80504 5550
rect 81058 5516 81522 5550
rect 82076 5516 82540 5550
rect 83094 5516 83558 5550
rect 84112 5516 84576 5550
rect 85130 5516 85594 5550
rect 86148 5516 86612 5550
rect 87166 5516 87630 5550
rect 67824 4994 68288 5028
rect 68842 4994 69306 5028
rect 69860 4994 70324 5028
rect 70878 4994 71342 5028
rect 71896 4994 72360 5028
rect 72914 4994 73378 5028
rect 73932 4994 74396 5028
rect 74950 4994 75414 5028
rect 75968 4994 76432 5028
rect 76986 4994 77450 5028
rect 78004 4994 78468 5028
rect 79022 4994 79486 5028
rect 80040 4994 80504 5028
rect 81058 4994 81522 5028
rect 82076 4994 82540 5028
rect 83094 4994 83558 5028
rect 84112 4994 84576 5028
rect 85130 4994 85594 5028
rect 86148 4994 86612 5028
rect 87166 4994 87630 5028
rect 55839 4797 56303 4831
rect 56857 4797 57321 4831
rect 57875 4797 58339 4831
rect 58893 4797 59357 4831
rect 59911 4797 60375 4831
rect 60929 4797 61393 4831
rect 62654 4798 62758 4832
rect 62952 4798 63056 4832
rect 63250 4798 63354 4832
rect 63548 4798 63652 4832
rect 63846 4798 63950 4832
rect 64144 4798 64248 4832
rect 64442 4798 64546 4832
rect 64740 4798 64844 4832
rect 65038 4798 65142 4832
rect 65336 4798 65440 4832
rect 65634 4798 65738 4832
rect 55545 4171 55579 4747
rect 56563 4171 56597 4747
rect 57581 4171 57615 4747
rect 58599 4171 58633 4747
rect 59617 4171 59651 4747
rect 60635 4171 60669 4747
rect 61653 4171 61687 4747
rect 62540 4172 62574 4748
rect 62838 4172 62872 4748
rect 63136 4172 63170 4748
rect 63434 4172 63468 4748
rect 63732 4172 63766 4748
rect 64030 4172 64064 4748
rect 64328 4172 64362 4748
rect 64626 4172 64660 4748
rect 64924 4172 64958 4748
rect 65222 4172 65256 4748
rect 65520 4172 65554 4748
rect 65818 4172 65852 4748
rect 67530 4368 67564 4944
rect 68548 4368 68582 4944
rect 69566 4368 69600 4944
rect 70584 4368 70618 4944
rect 71602 4368 71636 4944
rect 72620 4368 72654 4944
rect 73638 4368 73672 4944
rect 74656 4368 74690 4944
rect 75674 4368 75708 4944
rect 76692 4368 76726 4944
rect 77710 4368 77744 4944
rect 78728 4368 78762 4944
rect 79746 4368 79780 4944
rect 80764 4368 80798 4944
rect 81782 4368 81816 4944
rect 82800 4368 82834 4944
rect 83818 4368 83852 4944
rect 84836 4368 84870 4944
rect 85854 4368 85888 4944
rect 86872 4368 86906 4944
rect 87890 4368 87924 4944
rect 67824 4284 68288 4318
rect 68842 4284 69306 4318
rect 69860 4284 70324 4318
rect 70878 4284 71342 4318
rect 71896 4284 72360 4318
rect 72914 4284 73378 4318
rect 73932 4284 74396 4318
rect 74950 4284 75414 4318
rect 75968 4284 76432 4318
rect 76986 4284 77450 4318
rect 78004 4284 78468 4318
rect 79022 4284 79486 4318
rect 80040 4284 80504 4318
rect 81058 4284 81522 4318
rect 82076 4284 82540 4318
rect 83094 4284 83558 4318
rect 84112 4284 84576 4318
rect 85130 4284 85594 4318
rect 86148 4284 86612 4318
rect 87166 4284 87630 4318
rect 55839 4087 56303 4121
rect 56857 4087 57321 4121
rect 57875 4087 58339 4121
rect 58893 4087 59357 4121
rect 59911 4087 60375 4121
rect 60929 4087 61393 4121
rect 62654 4088 62758 4122
rect 62952 4088 63056 4122
rect 63250 4088 63354 4122
rect 63548 4088 63652 4122
rect 63846 4088 63950 4122
rect 64144 4088 64248 4122
rect 64442 4088 64546 4122
rect 64740 4088 64844 4122
rect 65038 4088 65142 4122
rect 65336 4088 65440 4122
rect 65634 4088 65738 4122
rect 67824 3760 68288 3794
rect 68842 3760 69306 3794
rect 69860 3760 70324 3794
rect 70878 3760 71342 3794
rect 71896 3760 72360 3794
rect 72914 3760 73378 3794
rect 73932 3760 74396 3794
rect 74950 3760 75414 3794
rect 75968 3760 76432 3794
rect 76986 3760 77450 3794
rect 78004 3760 78468 3794
rect 79022 3760 79486 3794
rect 80040 3760 80504 3794
rect 81058 3760 81522 3794
rect 82076 3760 82540 3794
rect 83094 3760 83558 3794
rect 84112 3760 84576 3794
rect 85130 3760 85594 3794
rect 86148 3760 86612 3794
rect 87166 3760 87630 3794
rect 55838 3684 56302 3718
rect 56856 3684 57320 3718
rect 57874 3684 58338 3718
rect 58892 3684 59356 3718
rect 59910 3684 60374 3718
rect 60928 3684 61392 3718
rect 62654 3686 62758 3720
rect 62952 3686 63056 3720
rect 63250 3686 63354 3720
rect 63548 3686 63652 3720
rect 63846 3686 63950 3720
rect 64144 3686 64248 3720
rect 64442 3686 64546 3720
rect 64740 3686 64844 3720
rect 65038 3686 65142 3720
rect 65336 3686 65440 3720
rect 65634 3686 65738 3720
rect 55544 3058 55578 3634
rect 56562 3058 56596 3634
rect 57580 3058 57614 3634
rect 58598 3058 58632 3634
rect 59616 3058 59650 3634
rect 60634 3058 60668 3634
rect 61652 3058 61686 3634
rect 62540 3060 62574 3636
rect 62838 3060 62872 3636
rect 63136 3060 63170 3636
rect 63434 3060 63468 3636
rect 63732 3060 63766 3636
rect 64030 3060 64064 3636
rect 64328 3060 64362 3636
rect 64626 3060 64660 3636
rect 64924 3060 64958 3636
rect 65222 3060 65256 3636
rect 65520 3060 65554 3636
rect 65818 3060 65852 3636
rect 67530 3134 67564 3710
rect 68548 3134 68582 3710
rect 69566 3134 69600 3710
rect 70584 3134 70618 3710
rect 71602 3134 71636 3710
rect 72620 3134 72654 3710
rect 73638 3134 73672 3710
rect 74656 3134 74690 3710
rect 75674 3134 75708 3710
rect 76692 3134 76726 3710
rect 77710 3134 77744 3710
rect 78728 3134 78762 3710
rect 79746 3134 79780 3710
rect 80764 3134 80798 3710
rect 81782 3134 81816 3710
rect 82800 3134 82834 3710
rect 83818 3134 83852 3710
rect 84836 3134 84870 3710
rect 85854 3134 85888 3710
rect 86872 3134 86906 3710
rect 87890 3134 87924 3710
rect 67824 3050 68288 3084
rect 68842 3050 69306 3084
rect 69860 3050 70324 3084
rect 70878 3050 71342 3084
rect 71896 3050 72360 3084
rect 72914 3050 73378 3084
rect 73932 3050 74396 3084
rect 74950 3050 75414 3084
rect 75968 3050 76432 3084
rect 76986 3050 77450 3084
rect 78004 3050 78468 3084
rect 79022 3050 79486 3084
rect 80040 3050 80504 3084
rect 81058 3050 81522 3084
rect 82076 3050 82540 3084
rect 83094 3050 83558 3084
rect 84112 3050 84576 3084
rect 85130 3050 85594 3084
rect 86148 3050 86612 3084
rect 87166 3050 87630 3084
rect 55838 2974 56302 3008
rect 56856 2974 57320 3008
rect 57874 2974 58338 3008
rect 58892 2974 59356 3008
rect 59910 2974 60374 3008
rect 60928 2974 61392 3008
rect 62654 2976 62758 3010
rect 62952 2976 63056 3010
rect 63250 2976 63354 3010
rect 63548 2976 63652 3010
rect 63846 2976 63950 3010
rect 64144 2976 64248 3010
rect 64442 2976 64546 3010
rect 64740 2976 64844 3010
rect 65038 2976 65142 3010
rect 65336 2976 65440 3010
rect 65634 2976 65738 3010
rect 55839 2573 56303 2607
rect 56857 2573 57321 2607
rect 57875 2573 58339 2607
rect 58893 2573 59357 2607
rect 59911 2573 60375 2607
rect 60929 2573 61393 2607
rect 62652 2574 62756 2608
rect 62950 2574 63054 2608
rect 63248 2574 63352 2608
rect 63546 2574 63650 2608
rect 63844 2574 63948 2608
rect 64142 2574 64246 2608
rect 64440 2574 64544 2608
rect 64738 2574 64842 2608
rect 65036 2574 65140 2608
rect 65334 2574 65438 2608
rect 65632 2574 65736 2608
rect 55545 1947 55579 2523
rect 56563 1947 56597 2523
rect 57581 1947 57615 2523
rect 58599 1947 58633 2523
rect 59617 1947 59651 2523
rect 60635 1947 60669 2523
rect 61653 1947 61687 2523
rect 62538 1948 62572 2524
rect 62836 1948 62870 2524
rect 63134 1948 63168 2524
rect 63432 1948 63466 2524
rect 63730 1948 63764 2524
rect 64028 1948 64062 2524
rect 64326 1948 64360 2524
rect 64624 1948 64658 2524
rect 64922 1948 64956 2524
rect 65220 1948 65254 2524
rect 65518 1948 65552 2524
rect 67824 2526 68288 2560
rect 68842 2526 69306 2560
rect 69860 2526 70324 2560
rect 70878 2526 71342 2560
rect 71896 2526 72360 2560
rect 72914 2526 73378 2560
rect 73932 2526 74396 2560
rect 74950 2526 75414 2560
rect 75968 2526 76432 2560
rect 76986 2526 77450 2560
rect 78004 2526 78468 2560
rect 79022 2526 79486 2560
rect 80040 2526 80504 2560
rect 81058 2526 81522 2560
rect 82076 2526 82540 2560
rect 83094 2526 83558 2560
rect 84112 2526 84576 2560
rect 85130 2526 85594 2560
rect 86148 2526 86612 2560
rect 87166 2526 87630 2560
rect 65816 1948 65850 2524
rect 67530 1900 67564 2476
rect 55839 1863 56303 1897
rect 56857 1863 57321 1897
rect 57875 1863 58339 1897
rect 58893 1863 59357 1897
rect 59911 1863 60375 1897
rect 60929 1863 61393 1897
rect 62652 1864 62756 1898
rect 62950 1864 63054 1898
rect 63248 1864 63352 1898
rect 63546 1864 63650 1898
rect 63844 1864 63948 1898
rect 64142 1864 64246 1898
rect 64440 1864 64544 1898
rect 64738 1864 64842 1898
rect 65036 1864 65140 1898
rect 65334 1864 65438 1898
rect 65632 1864 65736 1898
rect 68548 1900 68582 2476
rect 69566 1900 69600 2476
rect 70584 1900 70618 2476
rect 71602 1900 71636 2476
rect 72620 1900 72654 2476
rect 73638 1900 73672 2476
rect 74656 1900 74690 2476
rect 75674 1900 75708 2476
rect 76692 1900 76726 2476
rect 77710 1900 77744 2476
rect 78728 1900 78762 2476
rect 79746 1900 79780 2476
rect 80764 1900 80798 2476
rect 81782 1900 81816 2476
rect 82800 1900 82834 2476
rect 83818 1900 83852 2476
rect 84836 1900 84870 2476
rect 85854 1900 85888 2476
rect 86872 1900 86906 2476
rect 87890 1900 87924 2476
rect 67824 1816 68288 1850
rect 68842 1816 69306 1850
rect 69860 1816 70324 1850
rect 70878 1816 71342 1850
rect 71896 1816 72360 1850
rect 72914 1816 73378 1850
rect 73932 1816 74396 1850
rect 74950 1816 75414 1850
rect 75968 1816 76432 1850
rect 76986 1816 77450 1850
rect 78004 1816 78468 1850
rect 79022 1816 79486 1850
rect 80040 1816 80504 1850
rect 81058 1816 81522 1850
rect 82076 1816 82540 1850
rect 83094 1816 83558 1850
rect 84112 1816 84576 1850
rect 85130 1816 85594 1850
rect 86148 1816 86612 1850
rect 87166 1816 87630 1850
rect 55838 1460 56302 1494
rect 56856 1460 57320 1494
rect 57874 1460 58338 1494
rect 58892 1460 59356 1494
rect 59910 1460 60374 1494
rect 60928 1460 61392 1494
rect 62652 1464 62756 1498
rect 62950 1464 63054 1498
rect 63248 1464 63352 1498
rect 63546 1464 63650 1498
rect 63844 1464 63948 1498
rect 64142 1464 64246 1498
rect 64440 1464 64544 1498
rect 64738 1464 64842 1498
rect 65036 1464 65140 1498
rect 65334 1464 65438 1498
rect 65632 1464 65736 1498
rect 55544 834 55578 1410
rect 56562 834 56596 1410
rect 57580 834 57614 1410
rect 58598 834 58632 1410
rect 59616 834 59650 1410
rect 60634 834 60668 1410
rect 61652 834 61686 1410
rect 62538 838 62572 1414
rect 62836 838 62870 1414
rect 63134 838 63168 1414
rect 63432 838 63466 1414
rect 63730 838 63764 1414
rect 64028 838 64062 1414
rect 64326 838 64360 1414
rect 64624 838 64658 1414
rect 64922 838 64956 1414
rect 65220 838 65254 1414
rect 65518 838 65552 1414
rect 65816 838 65850 1414
rect 67824 1294 68288 1328
rect 68842 1294 69306 1328
rect 69860 1294 70324 1328
rect 70878 1294 71342 1328
rect 71896 1294 72360 1328
rect 72914 1294 73378 1328
rect 73932 1294 74396 1328
rect 74950 1294 75414 1328
rect 75968 1294 76432 1328
rect 76986 1294 77450 1328
rect 78004 1294 78468 1328
rect 79022 1294 79486 1328
rect 80040 1294 80504 1328
rect 81058 1294 81522 1328
rect 82076 1294 82540 1328
rect 83094 1294 83558 1328
rect 84112 1294 84576 1328
rect 85130 1294 85594 1328
rect 86148 1294 86612 1328
rect 87166 1294 87630 1328
rect 55838 750 56302 784
rect 56856 750 57320 784
rect 57874 750 58338 784
rect 58892 750 59356 784
rect 59910 750 60374 784
rect 60928 750 61392 784
rect 62652 754 62756 788
rect 62950 754 63054 788
rect 63248 754 63352 788
rect 63546 754 63650 788
rect 63844 754 63948 788
rect 64142 754 64246 788
rect 64440 754 64544 788
rect 64738 754 64842 788
rect 65036 754 65140 788
rect 65334 754 65438 788
rect 65632 754 65736 788
rect 67530 668 67564 1244
rect 68548 668 68582 1244
rect 69566 668 69600 1244
rect 70584 668 70618 1244
rect 71602 668 71636 1244
rect 72620 668 72654 1244
rect 73638 668 73672 1244
rect 74656 668 74690 1244
rect 75674 668 75708 1244
rect 76692 668 76726 1244
rect 77710 668 77744 1244
rect 78728 668 78762 1244
rect 79746 668 79780 1244
rect 80764 668 80798 1244
rect 81782 668 81816 1244
rect 82800 668 82834 1244
rect 83818 668 83852 1244
rect 84836 668 84870 1244
rect 85854 668 85888 1244
rect 86872 668 86906 1244
rect 87890 668 87924 1244
rect 67824 584 68288 618
rect 68842 584 69306 618
rect 69860 584 70324 618
rect 70878 584 71342 618
rect 71896 584 72360 618
rect 72914 584 73378 618
rect 73932 584 74396 618
rect 74950 584 75414 618
rect 75968 584 76432 618
rect 76986 584 77450 618
rect 78004 584 78468 618
rect 79022 584 79486 618
rect 80040 584 80504 618
rect 81058 584 81522 618
rect 82076 584 82540 618
rect 83094 584 83558 618
rect 84112 584 84576 618
rect 85130 584 85594 618
rect 86148 584 86612 618
rect 87166 584 87630 618
rect 89772 210 89872 14470
rect 52728 -682 52790 -582
rect 52790 -682 89710 -582
rect 89710 -682 89772 -582
<< metal1 >>
rect 11322 28262 35778 28268
rect 11322 28162 11428 28262
rect 35672 28162 35778 28262
rect 11322 28156 35778 28162
rect -1414 27642 -1354 27648
rect -8742 16408 -8682 16414
rect -1414 16408 -1354 27582
rect 11322 27642 11434 28156
rect 12034 27856 12044 28156
rect 35056 27856 35066 28156
rect 11322 18278 11328 27642
rect 11428 18278 11434 27642
rect 14948 27774 31828 27806
rect 14948 27560 15011 27774
rect 31796 27560 31828 27774
rect 14948 27540 31828 27560
rect 35666 27642 35778 28156
rect 65322 28262 89778 28268
rect 65322 28162 65428 28262
rect 89672 28162 89778 28262
rect 65322 28156 89778 28162
rect 14948 27538 19302 27540
rect 14564 21978 14952 22038
rect 14564 21838 14624 21978
rect 14666 21937 14726 21978
rect 14658 21931 14746 21937
rect 14658 21897 14670 21931
rect 14734 21897 14746 21931
rect 14658 21891 14746 21897
rect 14564 21810 14576 21838
rect 14570 21462 14576 21810
rect 14610 21810 14624 21838
rect 14782 21838 14842 21978
rect 14892 21937 14952 21978
rect 14876 21931 14964 21937
rect 14876 21897 14888 21931
rect 14952 21897 14964 21931
rect 14876 21891 14964 21897
rect 14610 21462 14616 21810
rect 14782 21806 14794 21838
rect 14788 21492 14794 21806
rect 14570 21450 14616 21462
rect 14782 21462 14794 21492
rect 14828 21806 14842 21838
rect 14998 21838 15058 27538
rect 15100 21978 15106 22038
rect 15166 21978 15172 22038
rect 15212 21978 15218 22038
rect 15278 21978 15284 22038
rect 15322 21978 15328 22038
rect 15388 21978 15394 22038
rect 15106 21937 15166 21978
rect 15094 21931 15182 21937
rect 15094 21897 15106 21931
rect 15170 21897 15182 21931
rect 15094 21891 15182 21897
rect 14828 21492 14834 21806
rect 14828 21462 14842 21492
rect 14658 21403 14746 21409
rect 14658 21369 14670 21403
rect 14734 21369 14746 21403
rect 14658 21363 14746 21369
rect 14782 21326 14842 21462
rect 14998 21462 15012 21838
rect 15046 21462 15058 21838
rect 15218 21838 15278 21978
rect 15328 21937 15388 21978
rect 15312 21931 15400 21937
rect 15312 21897 15324 21931
rect 15388 21897 15400 21931
rect 15312 21891 15400 21897
rect 15218 21812 15230 21838
rect 14876 21403 14964 21409
rect 14876 21369 14888 21403
rect 14952 21369 14964 21403
rect 14876 21363 14964 21369
rect 14892 21326 14952 21363
rect 14436 21266 14442 21326
rect 14502 21266 14508 21326
rect 14776 21266 14782 21326
rect 14842 21266 14848 21326
rect 14886 21266 14892 21326
rect 14952 21266 14958 21326
rect 13054 20320 13060 20380
rect 13120 20320 13126 20380
rect 11322 17764 11434 18278
rect 13060 18148 13120 20320
rect 14442 19542 14502 21266
rect 14998 21220 15058 21462
rect 15224 21462 15230 21812
rect 15264 21812 15278 21838
rect 15434 21838 15494 27538
rect 15530 21931 15618 21937
rect 15530 21897 15542 21931
rect 15606 21897 15618 21931
rect 15530 21891 15618 21897
rect 15748 21931 15836 21937
rect 15748 21897 15760 21931
rect 15824 21897 15836 21931
rect 15748 21891 15836 21897
rect 15264 21462 15270 21812
rect 15224 21450 15270 21462
rect 15434 21462 15448 21838
rect 15482 21462 15494 21838
rect 15660 21838 15706 21850
rect 15660 21494 15666 21838
rect 15094 21403 15182 21409
rect 15094 21369 15106 21403
rect 15170 21369 15182 21403
rect 15094 21363 15182 21369
rect 15312 21403 15400 21409
rect 15312 21369 15324 21403
rect 15388 21369 15400 21403
rect 15312 21363 15400 21369
rect 15434 21220 15494 21462
rect 15654 21462 15666 21494
rect 15700 21494 15706 21838
rect 15872 21838 15932 27538
rect 15972 21978 15978 22038
rect 16038 21978 16044 22038
rect 16082 21978 16088 22038
rect 16148 21978 16154 22038
rect 16190 21978 16196 22038
rect 16256 21978 16262 22038
rect 15978 21937 16038 21978
rect 15966 21931 16054 21937
rect 15966 21897 15978 21931
rect 16042 21897 16054 21931
rect 15966 21891 16054 21897
rect 15700 21462 15714 21494
rect 15530 21403 15618 21409
rect 15530 21369 15542 21403
rect 15606 21369 15618 21403
rect 15530 21363 15618 21369
rect 15542 21326 15602 21363
rect 15654 21326 15714 21462
rect 15872 21462 15884 21838
rect 15918 21462 15932 21838
rect 16088 21838 16148 21978
rect 16196 21937 16256 21978
rect 16184 21931 16272 21937
rect 16184 21897 16196 21931
rect 16260 21897 16272 21931
rect 16184 21891 16272 21897
rect 16088 21810 16102 21838
rect 15748 21403 15836 21409
rect 15748 21369 15760 21403
rect 15824 21369 15836 21403
rect 15748 21363 15836 21369
rect 15762 21326 15822 21363
rect 15536 21266 15542 21326
rect 15602 21266 15608 21326
rect 15648 21266 15654 21326
rect 15714 21266 15720 21326
rect 15756 21266 15762 21326
rect 15822 21266 15828 21326
rect 15872 21220 15932 21462
rect 16096 21462 16102 21810
rect 16136 21810 16148 21838
rect 16306 21838 16366 27538
rect 18930 27364 18936 27424
rect 18996 27364 19002 27424
rect 17424 27148 18502 27208
rect 17424 26968 17484 27148
rect 17928 27067 17988 27148
rect 17720 27061 18208 27067
rect 17720 27027 17732 27061
rect 18196 27027 18208 27061
rect 17720 27021 18208 27027
rect 17424 26928 17438 26968
rect 17432 26392 17438 26928
rect 17472 26928 17484 26968
rect 18442 26968 18502 27148
rect 18936 27067 18996 27364
rect 19462 27178 19522 27540
rect 20012 27364 20018 27424
rect 20078 27364 20084 27424
rect 20970 27364 20976 27424
rect 21036 27364 21042 27424
rect 19456 27118 19462 27178
rect 19522 27118 19528 27178
rect 18738 27061 19226 27067
rect 18738 27027 18750 27061
rect 19214 27027 19226 27061
rect 18738 27021 19226 27027
rect 18442 26942 18456 26968
rect 17472 26392 17478 26928
rect 18450 26428 18456 26942
rect 17432 26380 17478 26392
rect 18444 26392 18456 26428
rect 18490 26942 18502 26968
rect 19462 26968 19522 27118
rect 20018 27067 20078 27364
rect 20976 27067 21036 27364
rect 21498 27178 21558 27540
rect 22006 27364 22012 27424
rect 22072 27364 22078 27424
rect 23012 27364 23018 27424
rect 23078 27364 23084 27424
rect 21492 27118 21498 27178
rect 21558 27118 21564 27178
rect 19756 27061 20244 27067
rect 19756 27027 19768 27061
rect 20232 27027 20244 27061
rect 19756 27021 20244 27027
rect 20774 27061 21262 27067
rect 20774 27027 20786 27061
rect 21250 27027 21262 27061
rect 20774 27021 21262 27027
rect 20976 27018 21036 27021
rect 19462 26944 19474 26968
rect 18490 26428 18496 26942
rect 19468 26432 19474 26944
rect 18490 26392 18504 26428
rect 17720 26333 18208 26339
rect 17720 26299 17732 26333
rect 18196 26299 18208 26333
rect 17720 26293 18208 26299
rect 18444 26246 18504 26392
rect 19464 26392 19474 26432
rect 19508 26944 19522 26968
rect 20486 26968 20532 26980
rect 19508 26432 19514 26944
rect 19508 26392 19524 26432
rect 20486 26420 20492 26968
rect 18948 26339 19008 26340
rect 18738 26333 19226 26339
rect 18738 26299 18750 26333
rect 19214 26299 19226 26333
rect 18738 26293 19226 26299
rect 17274 26186 17280 26246
rect 17340 26186 17346 26246
rect 18438 26186 18444 26246
rect 18504 26186 18510 26246
rect 17144 25982 17150 26042
rect 17210 25982 17216 26042
rect 17150 23114 17210 25982
rect 17280 23572 17340 26186
rect 18438 25982 18444 26042
rect 18504 25982 18510 26042
rect 17720 25925 18208 25931
rect 17720 25891 17732 25925
rect 18196 25891 18208 25925
rect 17720 25885 18208 25891
rect 17432 25832 17478 25844
rect 17432 25292 17438 25832
rect 17426 25256 17438 25292
rect 17472 25292 17478 25832
rect 18444 25832 18504 25982
rect 18948 25931 19008 26293
rect 18738 25925 19226 25931
rect 18738 25891 18750 25925
rect 19214 25891 19226 25925
rect 18738 25885 19226 25891
rect 18948 25882 19008 25885
rect 18444 25794 18456 25832
rect 17472 25256 17486 25292
rect 18450 25286 18456 25794
rect 17426 25106 17486 25256
rect 18444 25256 18456 25286
rect 18490 25794 18504 25832
rect 19464 25832 19524 26392
rect 20480 26392 20492 26420
rect 20526 26420 20532 26968
rect 21498 26968 21558 27118
rect 22012 27067 22072 27364
rect 22510 27230 22516 27290
rect 22576 27230 22582 27290
rect 21792 27061 22280 27067
rect 21792 27027 21804 27061
rect 22268 27027 22280 27061
rect 21792 27021 22280 27027
rect 22012 27018 22072 27021
rect 21498 26944 21510 26968
rect 21504 26450 21510 26944
rect 20526 26392 20540 26420
rect 19970 26339 20030 26346
rect 19756 26333 20244 26339
rect 19756 26299 19768 26333
rect 20232 26299 20244 26333
rect 19756 26293 20244 26299
rect 19970 25931 20030 26293
rect 20480 26142 20540 26392
rect 21488 26392 21510 26450
rect 21544 26944 21558 26968
rect 22516 26968 22576 27230
rect 23018 27067 23078 27364
rect 23536 27180 23596 27540
rect 24034 27364 24040 27424
rect 24100 27364 24106 27424
rect 25052 27364 25058 27424
rect 25118 27364 25124 27424
rect 23530 27120 23536 27180
rect 23596 27120 23602 27180
rect 22810 27061 23298 27067
rect 22810 27027 22822 27061
rect 23286 27027 23298 27061
rect 22810 27021 23298 27027
rect 21544 26450 21550 26944
rect 22516 26940 22528 26968
rect 21544 26392 21552 26450
rect 21000 26339 21060 26346
rect 20774 26333 21262 26339
rect 20774 26299 20786 26333
rect 21250 26299 21262 26333
rect 20774 26293 21262 26299
rect 20474 26082 20480 26142
rect 20540 26082 20546 26142
rect 21000 25931 21060 26293
rect 19756 25925 20244 25931
rect 19756 25891 19768 25925
rect 20232 25891 20244 25925
rect 19756 25885 20244 25891
rect 20774 25925 21262 25931
rect 20774 25891 20786 25925
rect 21250 25891 21262 25925
rect 20774 25885 21262 25891
rect 18490 25286 18496 25794
rect 19464 25792 19474 25832
rect 18490 25256 18504 25286
rect 19468 25282 19474 25792
rect 17720 25197 18208 25203
rect 17720 25163 17732 25197
rect 18196 25163 18208 25197
rect 17720 25157 18208 25163
rect 17938 25106 17998 25157
rect 18444 25106 18504 25256
rect 19460 25256 19474 25282
rect 19508 25792 19524 25832
rect 20486 25832 20532 25844
rect 19508 25282 19514 25792
rect 19508 25256 19520 25282
rect 20486 25276 20492 25832
rect 18930 25203 18990 25210
rect 18738 25197 19226 25203
rect 18738 25163 18750 25197
rect 19214 25163 19226 25197
rect 18738 25157 19226 25163
rect 17426 25046 18504 25106
rect 18438 24898 18498 24904
rect 17428 24838 18498 24898
rect 17428 24696 17488 24838
rect 17938 24795 17998 24838
rect 17720 24789 18208 24795
rect 17720 24755 17732 24789
rect 18196 24755 18208 24789
rect 17720 24749 18208 24755
rect 17428 24664 17438 24696
rect 17432 24120 17438 24664
rect 17472 24664 17488 24696
rect 18438 24696 18498 24838
rect 18930 24795 18990 25157
rect 19460 25108 19520 25256
rect 20478 25256 20492 25276
rect 20526 25276 20532 25832
rect 21488 25832 21552 26392
rect 22522 26392 22528 26940
rect 22562 26940 22576 26968
rect 23536 26968 23596 27120
rect 24040 27067 24100 27364
rect 25058 27067 25118 27364
rect 25568 27180 25628 27540
rect 26076 27364 26082 27424
rect 26142 27364 26148 27424
rect 27088 27364 27094 27424
rect 27154 27364 27160 27424
rect 25560 27120 25566 27180
rect 25626 27120 25632 27180
rect 23828 27061 24316 27067
rect 23828 27027 23840 27061
rect 24304 27027 24316 27061
rect 23828 27021 24316 27027
rect 24846 27061 25334 27067
rect 24846 27027 24858 27061
rect 25322 27027 25334 27061
rect 24846 27021 25334 27027
rect 22562 26392 22568 26940
rect 23536 26928 23546 26968
rect 23540 26446 23546 26928
rect 22522 26380 22568 26392
rect 23524 26392 23546 26446
rect 23580 26928 23596 26968
rect 24558 26968 24604 26980
rect 23580 26446 23586 26928
rect 23580 26392 23588 26446
rect 24558 26432 24564 26968
rect 22000 26339 22060 26352
rect 23018 26339 23078 26346
rect 21792 26333 22280 26339
rect 21792 26299 21804 26333
rect 22268 26299 22280 26333
rect 21792 26293 22280 26299
rect 22810 26333 23298 26339
rect 22810 26299 22822 26333
rect 23286 26299 23298 26333
rect 22810 26293 23298 26299
rect 22000 25931 22060 26293
rect 22510 26082 22516 26142
rect 22576 26082 22582 26142
rect 21792 25925 22280 25931
rect 21792 25891 21804 25925
rect 22268 25891 22280 25925
rect 21792 25885 22280 25891
rect 21488 25802 21510 25832
rect 21504 25284 21510 25802
rect 20526 25256 20538 25276
rect 19976 25203 20036 25210
rect 19756 25197 20244 25203
rect 19756 25163 19768 25197
rect 20232 25163 20244 25197
rect 19756 25157 20244 25163
rect 19454 25048 19460 25108
rect 19520 25048 19526 25108
rect 18738 24789 19226 24795
rect 18738 24755 18750 24789
rect 19214 24755 19226 24789
rect 18738 24749 19226 24755
rect 18438 24664 18456 24696
rect 17472 24120 17478 24664
rect 18450 24162 18456 24664
rect 17432 24108 17478 24120
rect 18438 24120 18456 24162
rect 18490 24664 18498 24696
rect 19460 24696 19520 25048
rect 19976 24795 20036 25157
rect 20478 25012 20538 25256
rect 21496 25256 21510 25284
rect 21544 25802 21552 25832
rect 22516 25832 22576 26082
rect 23018 25931 23078 26293
rect 22810 25925 23298 25931
rect 22810 25891 22822 25925
rect 23286 25891 23298 25925
rect 22810 25885 23298 25891
rect 21544 25284 21550 25802
rect 22516 25794 22528 25832
rect 22522 25292 22528 25794
rect 21544 25282 21556 25284
rect 21544 25256 21560 25282
rect 20774 25197 21262 25203
rect 20774 25163 20786 25197
rect 21250 25163 21262 25197
rect 20774 25157 21262 25163
rect 21496 25108 21560 25256
rect 22514 25256 22528 25292
rect 22562 25794 22576 25832
rect 23524 25832 23588 26392
rect 24554 26392 24564 26432
rect 24598 26432 24604 26968
rect 25568 26968 25628 27120
rect 26082 27067 26142 27364
rect 27094 27067 27154 27364
rect 27608 27182 27668 27540
rect 28106 27364 28112 27424
rect 28172 27364 28178 27424
rect 29118 27364 29124 27424
rect 29184 27364 29190 27424
rect 27602 27122 27608 27182
rect 27668 27122 27674 27182
rect 25864 27061 26352 27067
rect 25864 27027 25876 27061
rect 26340 27027 26352 27061
rect 25864 27021 26352 27027
rect 26882 27061 27370 27067
rect 26882 27027 26894 27061
rect 27358 27027 27370 27061
rect 26882 27021 27370 27027
rect 25568 26928 25582 26968
rect 25576 26448 25582 26928
rect 24598 26392 24614 26432
rect 24042 26339 24102 26342
rect 23828 26333 24316 26339
rect 23828 26299 23840 26333
rect 24304 26299 24316 26333
rect 23828 26293 24316 26299
rect 24042 25931 24102 26293
rect 24554 26246 24614 26392
rect 25566 26392 25582 26448
rect 25616 26928 25628 26968
rect 26594 26968 26640 26980
rect 25616 26448 25622 26928
rect 25616 26392 25630 26448
rect 26594 26430 26600 26968
rect 25060 26339 25120 26348
rect 24846 26333 25334 26339
rect 24846 26299 24858 26333
rect 25322 26299 25334 26333
rect 24846 26293 25334 26299
rect 24548 26186 24554 26246
rect 24614 26186 24620 26246
rect 24544 25982 24550 26042
rect 24610 25982 24616 26042
rect 23828 25925 24316 25931
rect 23828 25891 23840 25925
rect 24304 25891 24316 25925
rect 23828 25885 24316 25891
rect 24042 25884 24102 25885
rect 23524 25798 23546 25832
rect 22562 25292 22568 25794
rect 23540 25292 23546 25798
rect 22562 25256 22578 25292
rect 22024 25203 22084 25216
rect 21792 25197 22280 25203
rect 21792 25163 21804 25197
rect 22268 25163 22280 25197
rect 21792 25157 22280 25163
rect 21490 25048 21496 25108
rect 21556 25048 21562 25108
rect 20472 24952 20478 25012
rect 20538 24952 20544 25012
rect 21176 24946 21182 25010
rect 21246 24946 21252 25010
rect 21182 24916 21246 24946
rect 20480 24852 21246 24916
rect 19756 24789 20244 24795
rect 19756 24755 19768 24789
rect 20232 24755 20244 24789
rect 19756 24749 20244 24755
rect 18490 24162 18496 24664
rect 19460 24644 19474 24696
rect 18490 24120 18502 24162
rect 19468 24156 19474 24644
rect 17720 24061 18208 24067
rect 17720 24027 17732 24061
rect 18196 24027 18208 24061
rect 17720 24021 18208 24027
rect 18438 23722 18502 24120
rect 19460 24120 19474 24156
rect 19508 24644 19520 24696
rect 20480 24696 20544 24852
rect 20774 24789 21262 24795
rect 20774 24755 20786 24789
rect 21250 24755 21262 24789
rect 20774 24749 21262 24755
rect 20480 24650 20492 24696
rect 19508 24156 19514 24644
rect 19508 24120 19520 24156
rect 20486 24144 20492 24650
rect 18738 24061 19226 24067
rect 18738 24027 18750 24061
rect 19214 24027 19226 24061
rect 18738 24021 19226 24027
rect 19460 23970 19520 24120
rect 20476 24120 20492 24144
rect 20526 24650 20544 24696
rect 21496 24696 21560 25048
rect 22024 24795 22084 25157
rect 22514 25010 22578 25256
rect 23530 25256 23546 25292
rect 23580 25798 23588 25832
rect 24550 25832 24610 25982
rect 25060 25931 25120 26293
rect 24846 25925 25334 25931
rect 24846 25891 24858 25925
rect 25322 25891 25334 25925
rect 24846 25885 25334 25891
rect 24550 25806 24564 25832
rect 23580 25292 23586 25798
rect 23580 25290 23590 25292
rect 23580 25256 23594 25290
rect 23042 25203 23102 25206
rect 22810 25197 23298 25203
rect 22810 25163 22822 25197
rect 23286 25163 23298 25197
rect 22810 25157 23298 25163
rect 22348 24946 22354 25010
rect 22418 24946 22578 25010
rect 22510 24842 22516 24902
rect 22576 24842 22582 24902
rect 21792 24789 22280 24795
rect 21792 24755 21804 24789
rect 22268 24755 22280 24789
rect 21792 24749 22280 24755
rect 20526 24144 20532 24650
rect 21496 24648 21510 24696
rect 21504 24146 21510 24648
rect 20526 24120 20540 24144
rect 19756 24061 20244 24067
rect 19756 24027 19768 24061
rect 20232 24027 20244 24061
rect 19756 24021 20244 24027
rect 19454 23910 19460 23970
rect 19520 23910 19526 23970
rect 20476 23860 20540 24120
rect 21496 24120 21510 24146
rect 21544 24648 21560 24696
rect 22516 24696 22576 24842
rect 23042 24795 23102 25157
rect 23530 25108 23594 25256
rect 24558 25256 24564 25806
rect 24598 25806 24610 25832
rect 25566 25832 25630 26392
rect 26588 26392 26600 26430
rect 26634 26430 26640 26968
rect 27608 26968 27668 27122
rect 28112 27067 28172 27364
rect 28614 27230 28620 27290
rect 28680 27230 28686 27290
rect 27900 27061 28388 27067
rect 27900 27027 27912 27061
rect 28376 27027 28388 27061
rect 27900 27021 28388 27027
rect 27608 26930 27618 26968
rect 27612 26432 27618 26930
rect 26634 26392 26648 26430
rect 26076 26339 26136 26345
rect 25864 26333 26352 26339
rect 25864 26299 25876 26333
rect 26340 26299 26352 26333
rect 25864 26293 26352 26299
rect 26076 25931 26136 26293
rect 26588 26246 26648 26392
rect 27604 26392 27618 26432
rect 27652 26930 27668 26968
rect 28620 26968 28680 27230
rect 29124 27067 29184 27364
rect 29640 27182 29700 27540
rect 30146 27364 30152 27424
rect 30212 27364 30218 27424
rect 31158 27364 31164 27424
rect 31224 27364 31230 27424
rect 29634 27122 29640 27182
rect 29700 27122 29706 27182
rect 28918 27061 29406 27067
rect 28918 27027 28930 27061
rect 29394 27027 29406 27061
rect 28918 27021 29406 27027
rect 27652 26432 27658 26930
rect 28620 26926 28636 26968
rect 27652 26392 27668 26432
rect 28630 26424 28636 26926
rect 27088 26339 27148 26345
rect 26882 26333 27370 26339
rect 26882 26299 26894 26333
rect 27358 26299 27370 26333
rect 26882 26293 27370 26299
rect 26582 26186 26588 26246
rect 26648 26186 26654 26246
rect 26580 25982 26586 26042
rect 26646 25982 26652 26042
rect 25864 25925 26352 25931
rect 25864 25891 25876 25925
rect 26340 25891 26352 25925
rect 25864 25885 26352 25891
rect 26076 25882 26136 25885
rect 24598 25256 24604 25806
rect 25566 25800 25582 25832
rect 25576 25304 25582 25800
rect 24558 25244 24604 25256
rect 25568 25256 25582 25304
rect 25616 25800 25630 25832
rect 26586 25832 26646 25982
rect 27088 25931 27148 26293
rect 26882 25925 27370 25931
rect 26882 25891 26894 25925
rect 27358 25891 27370 25925
rect 26882 25885 27370 25891
rect 27088 25882 27148 25885
rect 26586 25800 26600 25832
rect 25616 25304 25622 25800
rect 25616 25302 25628 25304
rect 25616 25256 25632 25302
rect 26594 25286 26600 25800
rect 24042 25203 24102 25210
rect 23828 25197 24316 25203
rect 23828 25163 23840 25197
rect 24304 25163 24316 25197
rect 23828 25157 24316 25163
rect 24846 25197 25334 25203
rect 24846 25163 24858 25197
rect 25322 25163 25334 25197
rect 24846 25157 25334 25163
rect 23524 25048 23530 25108
rect 23590 25048 23596 25108
rect 22810 24789 23298 24795
rect 22810 24755 22822 24789
rect 23286 24755 23298 24789
rect 22810 24749 23298 24755
rect 23042 24748 23102 24749
rect 22516 24660 22528 24696
rect 21544 24146 21550 24648
rect 22522 24168 22528 24660
rect 21544 24144 21556 24146
rect 21544 24120 21560 24144
rect 20774 24061 21262 24067
rect 20774 24027 20786 24061
rect 21250 24027 21262 24061
rect 20774 24021 21262 24027
rect 20470 23796 20476 23860
rect 20540 23796 20546 23860
rect 18432 23658 18438 23722
rect 18502 23658 18508 23722
rect 18262 23572 18322 23578
rect 17274 23512 17280 23572
rect 17340 23512 17346 23572
rect 17866 23236 17926 23242
rect 17150 23054 17812 23114
rect 16526 21970 16806 22030
rect 16992 21978 16998 22038
rect 17058 21978 17064 22038
rect 16402 21931 16490 21937
rect 16402 21897 16414 21931
rect 16478 21897 16490 21931
rect 16402 21891 16490 21897
rect 16136 21462 16142 21810
rect 16096 21450 16142 21462
rect 16306 21462 16320 21838
rect 16354 21462 16366 21838
rect 16526 21838 16586 21970
rect 16634 21937 16694 21970
rect 16620 21931 16708 21937
rect 16620 21897 16632 21931
rect 16696 21897 16708 21931
rect 16620 21891 16708 21897
rect 16526 21814 16538 21838
rect 16532 21508 16538 21814
rect 15966 21403 16054 21409
rect 15966 21369 15978 21403
rect 16042 21369 16054 21403
rect 15966 21363 16054 21369
rect 16184 21403 16272 21409
rect 16184 21369 16196 21403
rect 16260 21369 16272 21403
rect 16184 21363 16272 21369
rect 16306 21220 16366 21462
rect 16524 21462 16538 21508
rect 16572 21814 16586 21838
rect 16746 21838 16806 21970
rect 16572 21508 16578 21814
rect 16746 21806 16756 21838
rect 16572 21462 16584 21508
rect 16402 21403 16490 21409
rect 16402 21369 16414 21403
rect 16478 21369 16490 21403
rect 16402 21363 16490 21369
rect 16414 21326 16474 21363
rect 16524 21326 16584 21462
rect 16750 21462 16756 21806
rect 16790 21806 16806 21838
rect 16790 21462 16796 21806
rect 16750 21450 16796 21462
rect 16620 21403 16708 21409
rect 16620 21369 16632 21403
rect 16696 21369 16708 21403
rect 16620 21363 16708 21369
rect 16408 21266 16414 21326
rect 16474 21266 16480 21326
rect 16518 21266 16524 21326
rect 16584 21266 16590 21326
rect 14992 21160 14998 21220
rect 15058 21160 15064 21220
rect 15428 21160 15434 21220
rect 15494 21160 15500 21220
rect 15866 21160 15872 21220
rect 15932 21160 15938 21220
rect 16300 21160 16306 21220
rect 16366 21160 16372 21220
rect 14566 21042 14842 21102
rect 14566 20900 14626 21042
rect 14670 20999 14730 21042
rect 14658 20993 14746 20999
rect 14658 20959 14670 20993
rect 14734 20959 14746 20993
rect 14658 20953 14746 20959
rect 14566 20866 14576 20900
rect 14570 20524 14576 20866
rect 14610 20866 14626 20900
rect 14782 20900 14842 21042
rect 14876 20993 14964 20999
rect 14876 20959 14888 20993
rect 14952 20959 14964 20993
rect 14876 20953 14964 20959
rect 14782 20870 14794 20900
rect 14610 20524 14616 20866
rect 14788 20558 14794 20870
rect 14570 20512 14616 20524
rect 14782 20524 14794 20558
rect 14828 20870 14842 20900
rect 14998 20900 15058 21160
rect 15212 21044 15218 21104
rect 15278 21044 15284 21104
rect 15094 20993 15182 20999
rect 15094 20959 15106 20993
rect 15170 20959 15182 20993
rect 15094 20953 15182 20959
rect 14998 20872 15012 20900
rect 14828 20558 14834 20870
rect 15006 20566 15012 20872
rect 14828 20524 14842 20558
rect 14658 20465 14746 20471
rect 14658 20431 14670 20465
rect 14734 20431 14746 20465
rect 14658 20425 14746 20431
rect 14782 20380 14842 20524
rect 14998 20524 15012 20566
rect 15046 20872 15058 20900
rect 15218 20900 15278 21044
rect 15312 20993 15400 20999
rect 15312 20959 15324 20993
rect 15388 20959 15400 20993
rect 15312 20953 15400 20959
rect 15218 20874 15230 20900
rect 15046 20566 15052 20872
rect 15046 20524 15058 20566
rect 14876 20465 14964 20471
rect 14876 20431 14888 20465
rect 14952 20431 14964 20465
rect 14876 20425 14964 20431
rect 14776 20320 14782 20380
rect 14842 20320 14848 20380
rect 14892 20182 14952 20425
rect 14998 20276 15058 20524
rect 15224 20524 15230 20874
rect 15264 20874 15278 20900
rect 15434 20900 15494 21160
rect 15530 20993 15618 20999
rect 15530 20959 15542 20993
rect 15606 20959 15618 20993
rect 15530 20953 15618 20959
rect 15748 20993 15836 20999
rect 15748 20959 15760 20993
rect 15824 20959 15836 20993
rect 15748 20953 15836 20959
rect 15264 20524 15270 20874
rect 15434 20870 15448 20900
rect 15442 20556 15448 20870
rect 15224 20512 15270 20524
rect 15434 20524 15448 20556
rect 15482 20870 15494 20900
rect 15660 20900 15706 20912
rect 15482 20556 15488 20870
rect 15660 20560 15666 20900
rect 15482 20524 15494 20556
rect 15094 20465 15182 20471
rect 15094 20431 15106 20465
rect 15170 20431 15182 20465
rect 15094 20425 15182 20431
rect 15312 20465 15400 20471
rect 15312 20431 15324 20465
rect 15388 20431 15400 20465
rect 15312 20425 15400 20431
rect 14992 20216 14998 20276
rect 15058 20216 15064 20276
rect 14564 20178 14952 20182
rect 14564 20122 14892 20178
rect 14564 19962 14624 20122
rect 14670 20061 14730 20122
rect 14658 20055 14746 20061
rect 14658 20021 14670 20055
rect 14734 20021 14746 20055
rect 14658 20015 14746 20021
rect 14564 19936 14576 19962
rect 14570 19586 14576 19936
rect 14610 19936 14624 19962
rect 14784 19962 14844 20122
rect 14886 20118 14892 20122
rect 14952 20118 14958 20178
rect 14892 20061 14952 20118
rect 14876 20055 14964 20061
rect 14876 20021 14888 20055
rect 14952 20021 14964 20055
rect 14876 20015 14964 20021
rect 14610 19586 14616 19936
rect 14784 19924 14794 19962
rect 14788 19612 14794 19924
rect 14570 19574 14616 19586
rect 14782 19586 14794 19612
rect 14828 19924 14844 19962
rect 14998 19962 15058 20216
rect 15106 20178 15166 20425
rect 15210 20320 15216 20380
rect 15276 20320 15282 20380
rect 15100 20118 15106 20178
rect 15166 20118 15172 20178
rect 15106 20061 15166 20118
rect 15094 20055 15182 20061
rect 15094 20021 15106 20055
rect 15170 20021 15182 20055
rect 15094 20015 15182 20021
rect 14998 19928 15012 19962
rect 14828 19612 14834 19924
rect 14828 19586 14842 19612
rect 15006 19610 15012 19928
rect 14658 19527 14746 19533
rect 14658 19493 14670 19527
rect 14734 19493 14746 19527
rect 14658 19487 14746 19493
rect 14442 19226 14502 19482
rect 14782 19442 14842 19586
rect 14998 19586 15012 19610
rect 15046 19928 15058 19962
rect 15216 19962 15276 20320
rect 15326 20178 15386 20425
rect 15434 20276 15494 20524
rect 15652 20524 15666 20560
rect 15700 20560 15706 20900
rect 15872 20900 15932 21160
rect 16082 21044 16088 21104
rect 16148 21044 16154 21104
rect 15966 20993 16054 20999
rect 15966 20959 15978 20993
rect 16042 20959 16054 20993
rect 15966 20953 16054 20959
rect 15872 20866 15884 20900
rect 15700 20524 15712 20560
rect 15878 20552 15884 20866
rect 15530 20465 15618 20471
rect 15530 20431 15542 20465
rect 15606 20431 15618 20465
rect 15530 20425 15618 20431
rect 15428 20216 15434 20276
rect 15494 20216 15500 20276
rect 15320 20118 15326 20178
rect 15386 20118 15392 20178
rect 15326 20061 15386 20118
rect 15312 20055 15400 20061
rect 15312 20021 15324 20055
rect 15388 20021 15400 20055
rect 15312 20015 15400 20021
rect 15216 19928 15230 19962
rect 15046 19610 15052 19928
rect 15046 19586 15058 19610
rect 14876 19527 14964 19533
rect 14876 19493 14888 19527
rect 14952 19493 14964 19527
rect 14876 19487 14964 19493
rect 14776 19382 14782 19442
rect 14842 19382 14848 19442
rect 14998 19344 15058 19586
rect 15224 19586 15230 19928
rect 15264 19928 15276 19962
rect 15434 19962 15494 20216
rect 15544 20178 15604 20425
rect 15652 20380 15712 20524
rect 15872 20524 15884 20552
rect 15918 20866 15932 20900
rect 16088 20900 16148 21044
rect 16184 20993 16272 20999
rect 16184 20959 16196 20993
rect 16260 20959 16272 20993
rect 16184 20953 16272 20959
rect 16088 20868 16102 20900
rect 15918 20552 15924 20866
rect 15918 20524 15932 20552
rect 15748 20465 15836 20471
rect 15748 20431 15760 20465
rect 15824 20431 15836 20465
rect 15748 20425 15836 20431
rect 15646 20320 15652 20380
rect 15712 20320 15718 20380
rect 15760 20178 15820 20425
rect 15872 20276 15932 20524
rect 16096 20524 16102 20868
rect 16136 20868 16148 20900
rect 16306 20900 16366 21160
rect 16526 21060 16806 21120
rect 16402 20993 16490 20999
rect 16402 20959 16414 20993
rect 16478 20959 16490 20993
rect 16402 20953 16490 20959
rect 16306 20878 16320 20900
rect 16136 20524 16142 20868
rect 16314 20554 16320 20878
rect 16096 20512 16142 20524
rect 16306 20524 16320 20554
rect 16354 20878 16366 20900
rect 16526 20900 16586 21060
rect 16636 20999 16696 21060
rect 16620 20993 16708 20999
rect 16620 20959 16632 20993
rect 16696 20959 16708 20993
rect 16620 20953 16708 20959
rect 16354 20554 16360 20878
rect 16526 20876 16538 20900
rect 16532 20560 16538 20876
rect 16354 20524 16366 20554
rect 15966 20465 16054 20471
rect 15966 20431 15978 20465
rect 16042 20431 16054 20465
rect 15966 20425 16054 20431
rect 16184 20465 16272 20471
rect 16184 20431 16196 20465
rect 16260 20431 16272 20465
rect 16184 20425 16272 20431
rect 15866 20216 15872 20276
rect 15932 20216 15938 20276
rect 15538 20118 15544 20178
rect 15604 20118 15610 20178
rect 15648 20118 15654 20178
rect 15714 20118 15720 20178
rect 15754 20118 15760 20178
rect 15820 20118 15826 20178
rect 15544 20061 15604 20118
rect 15530 20055 15618 20061
rect 15530 20021 15542 20055
rect 15606 20021 15618 20055
rect 15530 20015 15618 20021
rect 15264 19586 15270 19928
rect 15434 19926 15448 19962
rect 15442 19624 15448 19926
rect 15224 19574 15270 19586
rect 15434 19586 15448 19624
rect 15482 19926 15494 19962
rect 15654 19962 15714 20118
rect 15760 20061 15820 20118
rect 15748 20055 15836 20061
rect 15748 20021 15760 20055
rect 15824 20021 15836 20055
rect 15748 20015 15836 20021
rect 15654 19934 15666 19962
rect 15482 19624 15488 19926
rect 15482 19586 15494 19624
rect 15660 19616 15666 19934
rect 15094 19527 15182 19533
rect 15094 19493 15106 19527
rect 15170 19493 15182 19527
rect 15094 19487 15182 19493
rect 15312 19527 15400 19533
rect 15312 19493 15324 19527
rect 15388 19493 15400 19527
rect 15312 19487 15400 19493
rect 15434 19344 15494 19586
rect 15652 19586 15666 19616
rect 15700 19934 15714 19962
rect 15872 19962 15932 20216
rect 15978 20178 16038 20425
rect 16082 20320 16088 20380
rect 16148 20320 16154 20380
rect 15972 20118 15978 20178
rect 16038 20118 16044 20178
rect 15978 20061 16038 20118
rect 15966 20055 16054 20061
rect 15966 20021 15978 20055
rect 16042 20021 16054 20055
rect 15966 20015 16054 20021
rect 15700 19616 15706 19934
rect 15872 19922 15884 19962
rect 15878 19620 15884 19922
rect 15700 19586 15712 19616
rect 15530 19527 15618 19533
rect 15530 19493 15542 19527
rect 15606 19493 15618 19527
rect 15530 19487 15618 19493
rect 15652 19442 15712 19586
rect 15872 19586 15884 19620
rect 15918 19922 15932 19962
rect 16088 19962 16148 20320
rect 16196 20178 16256 20425
rect 16306 20276 16366 20524
rect 16526 20524 16538 20560
rect 16572 20876 16586 20900
rect 16746 20900 16806 21060
rect 16876 21044 16882 21104
rect 16942 21044 16948 21104
rect 16572 20560 16578 20876
rect 16746 20864 16756 20900
rect 16572 20524 16586 20560
rect 16402 20465 16490 20471
rect 16402 20431 16414 20465
rect 16478 20431 16490 20465
rect 16402 20425 16490 20431
rect 16300 20216 16306 20276
rect 16366 20216 16372 20276
rect 16190 20118 16196 20178
rect 16256 20118 16262 20178
rect 16196 20061 16256 20118
rect 16184 20055 16272 20061
rect 16184 20021 16196 20055
rect 16260 20021 16272 20055
rect 16184 20015 16272 20021
rect 16088 19936 16102 19962
rect 15918 19620 15924 19922
rect 15918 19586 15932 19620
rect 15748 19527 15836 19533
rect 15748 19493 15760 19527
rect 15824 19493 15836 19527
rect 15748 19487 15836 19493
rect 15646 19382 15652 19442
rect 15712 19382 15718 19442
rect 15872 19344 15932 19586
rect 16096 19586 16102 19936
rect 16136 19936 16148 19962
rect 16306 19962 16366 20216
rect 16412 20178 16472 20425
rect 16526 20380 16586 20524
rect 16750 20524 16756 20864
rect 16790 20864 16806 20900
rect 16790 20524 16796 20864
rect 16750 20512 16796 20524
rect 16620 20465 16708 20471
rect 16620 20431 16632 20465
rect 16696 20431 16708 20465
rect 16620 20425 16708 20431
rect 16520 20320 16526 20380
rect 16586 20320 16592 20380
rect 16406 20118 16412 20178
rect 16472 20118 16806 20178
rect 16412 20061 16472 20118
rect 16402 20055 16490 20061
rect 16402 20021 16414 20055
rect 16478 20021 16490 20055
rect 16402 20015 16490 20021
rect 16136 19586 16142 19936
rect 16306 19934 16320 19962
rect 16314 19620 16320 19934
rect 16096 19574 16142 19586
rect 16306 19586 16320 19620
rect 16354 19934 16366 19962
rect 16524 19962 16584 20118
rect 16632 20061 16692 20118
rect 16620 20055 16708 20061
rect 16620 20021 16632 20055
rect 16696 20021 16708 20055
rect 16620 20015 16708 20021
rect 16524 19944 16538 19962
rect 16354 19620 16360 19934
rect 16532 19620 16538 19944
rect 16354 19586 16366 19620
rect 15966 19527 16054 19533
rect 15966 19493 15978 19527
rect 16042 19493 16054 19527
rect 15966 19487 16054 19493
rect 16184 19527 16272 19533
rect 16184 19493 16196 19527
rect 16260 19493 16272 19527
rect 16184 19487 16272 19493
rect 16306 19344 16366 19586
rect 16526 19586 16538 19620
rect 16572 19944 16584 19962
rect 16746 19962 16806 20118
rect 16572 19620 16578 19944
rect 16746 19940 16756 19962
rect 16572 19586 16586 19620
rect 16402 19527 16490 19533
rect 16402 19493 16414 19527
rect 16478 19493 16490 19527
rect 16402 19487 16490 19493
rect 16526 19442 16586 19586
rect 16750 19586 16756 19940
rect 16790 19940 16806 19962
rect 16790 19586 16796 19940
rect 16750 19574 16796 19586
rect 16620 19527 16708 19533
rect 16620 19493 16632 19527
rect 16696 19493 16708 19527
rect 16620 19487 16708 19493
rect 16882 19442 16942 21044
rect 16520 19382 16526 19442
rect 16586 19382 16592 19442
rect 16876 19382 16882 19442
rect 16942 19382 16948 19442
rect 14992 19284 14998 19344
rect 15058 19284 15064 19344
rect 15428 19284 15434 19344
rect 15494 19284 15500 19344
rect 15866 19284 15872 19344
rect 15932 19284 15938 19344
rect 16300 19284 16306 19344
rect 16366 19284 16372 19344
rect 14436 19166 14442 19226
rect 14502 19166 14508 19226
rect 14566 19164 14952 19224
rect 14566 19024 14626 19164
rect 14672 19123 14732 19164
rect 14658 19117 14746 19123
rect 14658 19083 14670 19117
rect 14734 19083 14746 19117
rect 14658 19077 14746 19083
rect 14566 18994 14576 19024
rect 14570 18648 14576 18994
rect 14610 18994 14626 19024
rect 14782 19024 14842 19164
rect 14892 19123 14952 19164
rect 14876 19117 14964 19123
rect 14876 19083 14888 19117
rect 14952 19083 14964 19117
rect 14876 19077 14964 19083
rect 14782 19000 14794 19024
rect 14610 18648 14616 18994
rect 14788 18676 14794 19000
rect 14570 18636 14616 18648
rect 14782 18648 14794 18676
rect 14828 19000 14842 19024
rect 14998 19024 15058 19284
rect 15102 19166 15108 19226
rect 15168 19166 15174 19226
rect 15210 19166 15216 19226
rect 15276 19166 15282 19226
rect 15318 19166 15324 19226
rect 15384 19166 15390 19226
rect 15108 19123 15168 19166
rect 15094 19117 15182 19123
rect 15094 19083 15106 19117
rect 15170 19083 15182 19117
rect 15094 19077 15182 19083
rect 14828 18676 14834 19000
rect 14998 18996 15012 19024
rect 14828 18648 14842 18676
rect 14658 18589 14746 18595
rect 14658 18555 14670 18589
rect 14734 18555 14746 18589
rect 14658 18549 14746 18555
rect 14782 18506 14842 18648
rect 15006 18648 15012 18996
rect 15046 18996 15058 19024
rect 15216 19024 15276 19166
rect 15324 19123 15384 19166
rect 15312 19117 15400 19123
rect 15312 19083 15324 19117
rect 15388 19083 15400 19117
rect 15312 19077 15400 19083
rect 15216 19000 15230 19024
rect 15046 18648 15052 18996
rect 15006 18636 15052 18648
rect 15224 18648 15230 19000
rect 15264 19000 15276 19024
rect 15434 19024 15494 19284
rect 15530 19117 15618 19123
rect 15530 19083 15542 19117
rect 15606 19083 15618 19117
rect 15530 19077 15618 19083
rect 15748 19117 15836 19123
rect 15748 19083 15760 19117
rect 15824 19083 15836 19117
rect 15748 19077 15836 19083
rect 15264 18648 15270 19000
rect 15434 18994 15448 19024
rect 15224 18636 15270 18648
rect 15442 18648 15448 18994
rect 15482 18994 15494 19024
rect 15660 19024 15706 19036
rect 15482 18648 15488 18994
rect 15660 18678 15666 19024
rect 15442 18636 15488 18648
rect 15652 18648 15666 18678
rect 15700 18678 15706 19024
rect 15872 19024 15932 19284
rect 15964 19166 15970 19226
rect 16030 19166 16036 19226
rect 16082 19166 16088 19226
rect 16148 19166 16154 19226
rect 16191 19166 16197 19224
rect 16255 19166 16261 19224
rect 15970 19123 16030 19166
rect 15966 19117 16054 19123
rect 15966 19083 15978 19117
rect 16042 19083 16054 19117
rect 15966 19077 16054 19083
rect 15872 18990 15884 19024
rect 15700 18648 15712 18678
rect 14876 18589 14964 18595
rect 14876 18555 14888 18589
rect 14952 18555 14964 18589
rect 14876 18549 14964 18555
rect 15094 18589 15182 18595
rect 15094 18555 15106 18589
rect 15170 18555 15182 18589
rect 15094 18549 15182 18555
rect 15312 18589 15400 18595
rect 15312 18555 15324 18589
rect 15388 18555 15400 18589
rect 15312 18549 15400 18555
rect 15530 18589 15618 18595
rect 15530 18555 15542 18589
rect 15606 18555 15618 18589
rect 15530 18549 15618 18555
rect 14892 18506 14952 18549
rect 15546 18506 15606 18549
rect 15652 18506 15712 18648
rect 15878 18648 15884 18990
rect 15918 18990 15932 19024
rect 16088 19024 16148 19166
rect 16197 19123 16255 19166
rect 16184 19117 16272 19123
rect 16184 19083 16196 19117
rect 16260 19083 16272 19117
rect 16184 19077 16272 19083
rect 15918 18648 15924 18990
rect 16088 18984 16102 19024
rect 15878 18636 15924 18648
rect 16096 18648 16102 18984
rect 16136 18984 16148 19024
rect 16306 19024 16366 19284
rect 16526 19174 16806 19234
rect 16402 19117 16490 19123
rect 16402 19083 16414 19117
rect 16478 19083 16490 19117
rect 16402 19077 16490 19083
rect 16306 19002 16320 19024
rect 16136 18648 16142 18984
rect 16096 18636 16142 18648
rect 16314 18648 16320 19002
rect 16354 19002 16366 19024
rect 16526 19024 16586 19174
rect 16632 19123 16692 19174
rect 16620 19117 16708 19123
rect 16620 19083 16632 19117
rect 16696 19083 16708 19117
rect 16620 19077 16708 19083
rect 16354 18648 16360 19002
rect 16526 19000 16538 19024
rect 16532 18682 16538 19000
rect 16314 18636 16360 18648
rect 16526 18648 16538 18682
rect 16572 19000 16586 19024
rect 16746 19024 16806 19174
rect 16572 18682 16578 19000
rect 16746 18996 16756 19024
rect 16572 18648 16586 18682
rect 15748 18589 15836 18595
rect 15748 18555 15760 18589
rect 15824 18555 15836 18589
rect 15748 18549 15836 18555
rect 15966 18589 16054 18595
rect 15966 18555 15978 18589
rect 16042 18555 16054 18589
rect 15966 18549 16054 18555
rect 16184 18589 16272 18595
rect 16184 18555 16196 18589
rect 16260 18555 16272 18589
rect 16184 18549 16272 18555
rect 16402 18589 16490 18595
rect 16402 18555 16414 18589
rect 16478 18555 16490 18589
rect 16402 18549 16490 18555
rect 15762 18506 15822 18549
rect 16414 18506 16474 18549
rect 16526 18506 16586 18648
rect 16750 18648 16756 18996
rect 16790 18996 16806 19024
rect 16790 18648 16796 18996
rect 16750 18636 16796 18648
rect 16620 18589 16708 18595
rect 16620 18555 16632 18589
rect 16696 18555 16708 18589
rect 16620 18549 16708 18555
rect 16998 18506 17058 21978
rect 17752 20932 17812 23054
rect 17746 20872 17752 20932
rect 17812 20872 17818 20932
rect 17866 20828 17926 23176
rect 18262 23136 18322 23512
rect 20476 23426 20540 23796
rect 20982 23788 21042 24021
rect 21496 23970 21560 24120
rect 22514 24120 22528 24168
rect 22562 24660 22576 24696
rect 23530 24696 23594 25048
rect 24042 24795 24102 25157
rect 25070 24795 25130 25157
rect 25568 25106 25632 25256
rect 26588 25256 26600 25286
rect 26634 25800 26646 25832
rect 27604 25832 27668 26392
rect 28622 26392 28636 26424
rect 28670 26926 28680 26968
rect 29640 26968 29700 27122
rect 30152 27067 30212 27364
rect 31164 27067 31224 27364
rect 31676 27182 31736 27540
rect 32176 27364 32182 27424
rect 32242 27364 32248 27424
rect 31670 27122 31676 27182
rect 31736 27122 31742 27182
rect 29936 27061 30424 27067
rect 29936 27027 29948 27061
rect 30412 27027 30424 27061
rect 29936 27021 30424 27027
rect 30954 27061 31442 27067
rect 30954 27027 30966 27061
rect 31430 27027 31442 27061
rect 30954 27021 31442 27027
rect 29640 26940 29654 26968
rect 28670 26424 28676 26926
rect 29648 26440 29654 26940
rect 28670 26392 28682 26424
rect 28094 26339 28154 26345
rect 27900 26333 28388 26339
rect 27900 26299 27912 26333
rect 28376 26299 28388 26333
rect 27900 26293 28388 26299
rect 28094 25931 28154 26293
rect 28622 26240 28682 26392
rect 29640 26392 29654 26440
rect 29688 26940 29700 26968
rect 30666 26968 30712 26980
rect 29688 26440 29694 26940
rect 29688 26392 29700 26440
rect 30666 26424 30672 26968
rect 29112 26339 29172 26345
rect 28918 26333 29406 26339
rect 28918 26299 28930 26333
rect 29394 26299 29406 26333
rect 28918 26293 29406 26299
rect 28622 26180 28824 26240
rect 28616 26082 28622 26142
rect 28682 26082 28688 26142
rect 27900 25925 28388 25931
rect 27900 25891 27912 25925
rect 28376 25891 28388 25925
rect 27900 25885 28388 25891
rect 28094 25882 28154 25885
rect 26634 25286 26640 25800
rect 27604 25784 27618 25832
rect 27612 25300 27618 25784
rect 26634 25256 26648 25286
rect 26088 25203 26148 25215
rect 25864 25197 26352 25203
rect 25864 25163 25876 25197
rect 26340 25163 26352 25197
rect 25864 25157 26352 25163
rect 25562 25046 25568 25106
rect 25628 25046 25634 25106
rect 23828 24789 24316 24795
rect 23828 24755 23840 24789
rect 24304 24755 24316 24789
rect 23828 24749 24316 24755
rect 24846 24789 25334 24795
rect 24846 24755 24858 24789
rect 25322 24755 25334 24789
rect 24846 24749 25334 24755
rect 25070 24742 25130 24749
rect 22562 24168 22568 24660
rect 23530 24636 23546 24696
rect 22562 24120 22574 24168
rect 23540 24154 23546 24636
rect 21792 24061 22280 24067
rect 21792 24027 21804 24061
rect 22268 24027 22280 24061
rect 21792 24021 22280 24027
rect 21490 23910 21496 23970
rect 21556 23910 21562 23970
rect 22024 23788 22084 24021
rect 20982 23728 22084 23788
rect 20470 23362 20476 23426
rect 20540 23362 20546 23426
rect 20982 23324 21042 23728
rect 20444 23264 21042 23324
rect 18256 23076 18262 23136
rect 18322 23076 18328 23136
rect 19422 23076 19428 23136
rect 19488 23076 19494 23136
rect 17988 22030 17994 22090
rect 18054 22030 18060 22090
rect 17860 20768 17866 20828
rect 17926 20768 17932 20828
rect 14776 18446 14782 18506
rect 14842 18446 14848 18506
rect 14886 18446 14892 18506
rect 14952 18446 14958 18506
rect 15540 18446 15546 18506
rect 15606 18446 15612 18506
rect 15646 18446 15652 18506
rect 15712 18446 15718 18506
rect 15756 18446 15762 18506
rect 15822 18446 15828 18506
rect 16408 18446 16414 18506
rect 16474 18446 16480 18506
rect 16520 18446 16526 18506
rect 16586 18446 16592 18506
rect 16992 18446 16998 18506
rect 17058 18446 17064 18506
rect 17994 18418 18054 22030
rect 18124 21932 18130 21992
rect 18190 21932 18196 21992
rect 17988 18358 17994 18418
rect 18054 18358 18060 18418
rect 18130 18288 18190 21932
rect 18262 19468 18322 23076
rect 18706 23015 19194 23021
rect 18706 22981 18718 23015
rect 19182 22981 19194 23015
rect 18706 22975 19194 22981
rect 18418 22922 18464 22934
rect 18418 22382 18424 22922
rect 18410 22346 18424 22382
rect 18458 22382 18464 22922
rect 19428 22922 19488 23076
rect 19724 23015 20212 23021
rect 19724 22981 19736 23015
rect 20200 22981 20212 23015
rect 19724 22975 20212 22981
rect 19428 22896 19442 22922
rect 18458 22346 18470 22382
rect 19436 22370 19442 22896
rect 18410 22188 18470 22346
rect 19426 22346 19442 22370
rect 19476 22896 19488 22922
rect 20444 22922 20504 23264
rect 22514 23236 22574 24120
rect 23530 24120 23546 24154
rect 23580 24636 23594 24696
rect 24558 24696 24604 24708
rect 23580 24154 23586 24636
rect 23580 24152 23590 24154
rect 24558 24152 24564 24696
rect 23580 24120 23594 24152
rect 22810 24061 23298 24067
rect 22810 24027 22822 24061
rect 23286 24027 23298 24061
rect 22810 24021 23298 24027
rect 23530 23974 23594 24120
rect 24548 24120 24564 24152
rect 24598 24152 24604 24696
rect 25568 24696 25632 25046
rect 26088 24795 26148 25157
rect 26588 25008 26648 25256
rect 27604 25256 27618 25300
rect 27652 25784 27668 25832
rect 28622 25832 28682 26082
rect 28764 26038 28824 26180
rect 28758 25978 28764 26038
rect 28824 25978 28830 26038
rect 29112 25931 29172 26293
rect 28918 25925 29406 25931
rect 28918 25891 28930 25925
rect 29394 25891 29406 25925
rect 28918 25885 29406 25891
rect 29112 25882 29172 25885
rect 28622 25808 28636 25832
rect 27652 25300 27658 25784
rect 27652 25298 27664 25300
rect 27652 25256 27668 25298
rect 27088 25203 27148 25211
rect 26882 25197 27370 25203
rect 26882 25163 26894 25197
rect 27358 25163 27370 25197
rect 26882 25157 27370 25163
rect 26582 24948 26588 25008
rect 26648 24948 26654 25008
rect 27088 24795 27148 25157
rect 27604 25106 27668 25256
rect 28630 25256 28636 25808
rect 28670 25808 28682 25832
rect 29640 25832 29700 26392
rect 30656 26392 30672 26424
rect 30706 26424 30712 26968
rect 31676 26968 31736 27122
rect 32182 27067 32242 27364
rect 32696 27130 33776 27190
rect 31972 27061 32460 27067
rect 31972 27027 31984 27061
rect 32448 27027 32460 27061
rect 31972 27021 32460 27027
rect 31676 26936 31690 26968
rect 31684 26430 31690 26936
rect 30706 26392 30716 26424
rect 30130 26339 30190 26345
rect 29936 26333 30424 26339
rect 29936 26299 29948 26333
rect 30412 26299 30424 26333
rect 29936 26293 30424 26299
rect 30130 25931 30190 26293
rect 30656 26142 30716 26392
rect 31680 26392 31690 26430
rect 31724 26936 31736 26968
rect 32696 26968 32756 27130
rect 33198 27067 33258 27130
rect 32990 27061 33478 27067
rect 32990 27027 33002 27061
rect 33466 27027 33478 27061
rect 32990 27021 33478 27027
rect 32696 26938 32708 26968
rect 31724 26430 31730 26936
rect 32702 26432 32708 26938
rect 31724 26392 31740 26430
rect 31130 26339 31190 26345
rect 30954 26333 31442 26339
rect 30954 26299 30966 26333
rect 31430 26299 31442 26333
rect 30954 26293 31442 26299
rect 30650 26082 30656 26142
rect 30716 26082 30722 26142
rect 30652 25978 30658 26038
rect 30718 25978 30724 26038
rect 29936 25925 30424 25931
rect 29936 25891 29948 25925
rect 30412 25891 30424 25925
rect 29936 25885 30424 25891
rect 30130 25882 30190 25885
rect 28670 25256 28676 25808
rect 29640 25788 29654 25832
rect 29648 25292 29654 25788
rect 28630 25244 28676 25256
rect 29640 25256 29654 25292
rect 29688 25788 29700 25832
rect 30658 25832 30718 25978
rect 31130 25931 31190 26293
rect 30954 25925 31442 25931
rect 30954 25891 30966 25925
rect 31430 25891 31442 25925
rect 30954 25885 31442 25891
rect 31130 25882 31190 25885
rect 30658 25804 30672 25832
rect 29688 25292 29694 25788
rect 30666 25292 30672 25804
rect 29688 25256 29700 25292
rect 28094 25203 28154 25211
rect 29136 25203 29196 25211
rect 27900 25197 28388 25203
rect 27900 25163 27912 25197
rect 28376 25163 28388 25197
rect 27900 25157 28388 25163
rect 28918 25197 29406 25203
rect 28918 25163 28930 25197
rect 29394 25163 29406 25197
rect 28918 25157 29406 25163
rect 27598 25046 27604 25106
rect 27664 25046 27670 25106
rect 25864 24789 26352 24795
rect 25864 24755 25876 24789
rect 26340 24755 26352 24789
rect 25864 24749 26352 24755
rect 26882 24789 27370 24795
rect 26882 24755 26894 24789
rect 27358 24755 27370 24789
rect 26882 24749 27370 24755
rect 27088 24748 27148 24749
rect 25568 24656 25582 24696
rect 25576 24166 25582 24656
rect 24598 24120 24612 24152
rect 23828 24061 24316 24067
rect 23828 24027 23840 24061
rect 24304 24027 24316 24061
rect 23828 24021 24316 24027
rect 22990 23966 23050 23972
rect 22508 23176 22514 23236
rect 22574 23176 22580 23236
rect 21458 23076 21464 23136
rect 21524 23076 21530 23136
rect 20742 23015 21230 23021
rect 20742 22981 20754 23015
rect 21218 22981 21230 23015
rect 20742 22975 21230 22981
rect 19476 22370 19482 22896
rect 20444 22876 20460 22922
rect 20454 22370 20460 22876
rect 19476 22346 19486 22370
rect 18706 22287 19194 22293
rect 18706 22253 18718 22287
rect 19182 22253 19194 22287
rect 18706 22247 19194 22253
rect 18924 22188 18984 22247
rect 19426 22188 19486 22346
rect 20446 22346 20460 22370
rect 20494 22876 20504 22922
rect 21464 22922 21524 23076
rect 22990 23021 23050 23906
rect 23498 23970 23594 23974
rect 23498 23968 23530 23970
rect 23590 23910 23596 23970
rect 23984 23910 23990 23970
rect 24050 23910 24056 23970
rect 21760 23015 22248 23021
rect 21760 22981 21772 23015
rect 22236 22981 22248 23015
rect 21760 22975 22248 22981
rect 22778 23015 23266 23021
rect 22778 22981 22790 23015
rect 23254 22981 23266 23015
rect 22778 22975 23266 22981
rect 21464 22898 21478 22922
rect 20494 22370 20500 22876
rect 20494 22346 20506 22370
rect 19724 22287 20212 22293
rect 19724 22253 19736 22287
rect 20200 22253 20212 22287
rect 19724 22247 20212 22253
rect 18410 22128 19486 22188
rect 19426 21822 19432 21882
rect 19492 21822 19498 21882
rect 18706 21759 19194 21765
rect 18706 21725 18718 21759
rect 19182 21725 19194 21759
rect 18706 21719 19194 21725
rect 18418 21666 18464 21678
rect 18418 21126 18424 21666
rect 18414 21090 18424 21126
rect 18458 21126 18464 21666
rect 19432 21666 19492 21822
rect 19916 21765 19976 22247
rect 20446 22188 20506 22346
rect 21472 22346 21478 22898
rect 21512 22898 21524 22922
rect 22490 22922 22536 22934
rect 21512 22346 21518 22898
rect 22490 22374 22496 22922
rect 21472 22334 21518 22346
rect 22482 22346 22496 22374
rect 22530 22374 22536 22922
rect 23498 22922 23558 23908
rect 23990 23021 24050 23910
rect 24548 23722 24612 24120
rect 25568 24120 25582 24166
rect 25616 24656 25632 24696
rect 26594 24696 26640 24708
rect 25616 24166 25622 24656
rect 25616 24164 25628 24166
rect 25616 24120 25632 24164
rect 26594 24156 26600 24696
rect 24846 24061 25334 24067
rect 24846 24027 24858 24061
rect 25322 24027 25334 24061
rect 24846 24021 25334 24027
rect 25568 23978 25632 24120
rect 26584 24120 26600 24156
rect 26634 24156 26640 24696
rect 27604 24696 27668 25046
rect 28094 24795 28154 25157
rect 28616 24842 28622 24902
rect 28682 24842 28688 24902
rect 27900 24789 28388 24795
rect 27900 24755 27912 24789
rect 28376 24755 28388 24789
rect 27900 24749 28388 24755
rect 28094 24748 28154 24749
rect 27604 24644 27618 24696
rect 27612 24162 27618 24644
rect 26634 24120 26648 24156
rect 25864 24061 26352 24067
rect 25864 24027 25876 24061
rect 26340 24027 26352 24061
rect 25864 24021 26352 24027
rect 25034 23972 25094 23978
rect 24542 23658 24548 23722
rect 24612 23658 24618 23722
rect 24548 23438 24612 23658
rect 24548 23368 24612 23374
rect 25034 23021 25094 23912
rect 25536 23972 25632 23978
rect 25596 23968 25632 23972
rect 26050 23972 26110 23978
rect 25536 23908 25568 23912
rect 25628 23908 25634 23968
rect 23796 23015 24284 23021
rect 23796 22981 23808 23015
rect 24272 22981 24284 23015
rect 23796 22975 24284 22981
rect 24814 23015 25302 23021
rect 24814 22981 24826 23015
rect 25290 22981 25302 23015
rect 24814 22975 25302 22981
rect 25034 22968 25094 22975
rect 22530 22346 22542 22374
rect 20742 22287 21230 22293
rect 20742 22253 20754 22287
rect 21218 22253 21230 22287
rect 20742 22247 21230 22253
rect 21760 22287 22248 22293
rect 21760 22253 21772 22287
rect 22236 22253 22248 22287
rect 21760 22247 22248 22253
rect 20440 22128 20446 22188
rect 20506 22128 20512 22188
rect 20446 21992 20506 22128
rect 20440 21932 20446 21992
rect 20506 21932 20512 21992
rect 20954 21765 21014 22247
rect 21460 21934 21466 21994
rect 21526 21934 21532 21994
rect 21466 21882 21526 21934
rect 21460 21822 21466 21882
rect 21526 21822 21532 21882
rect 19724 21759 20212 21765
rect 19724 21725 19736 21759
rect 20200 21725 20212 21759
rect 19724 21719 20212 21725
rect 20742 21759 21230 21765
rect 20742 21725 20754 21759
rect 21218 21725 21230 21759
rect 20742 21719 21230 21725
rect 19432 21640 19442 21666
rect 18458 21090 18474 21126
rect 19436 21114 19442 21640
rect 18414 20932 18474 21090
rect 19430 21090 19442 21114
rect 19476 21640 19492 21666
rect 20454 21666 20500 21678
rect 19476 21114 19482 21640
rect 20454 21116 20460 21666
rect 19476 21090 19490 21114
rect 18706 21031 19194 21037
rect 18706 20997 18718 21031
rect 19182 20997 19194 21031
rect 18706 20991 19194 20997
rect 18928 20932 18988 20991
rect 19430 20932 19490 21090
rect 20448 21090 20460 21116
rect 20494 21116 20500 21666
rect 21466 21666 21526 21822
rect 21960 21765 22020 22247
rect 22482 22188 22542 22346
rect 23498 22346 23514 22922
rect 23548 22346 23558 22922
rect 24526 22922 24572 22934
rect 24526 22370 24532 22922
rect 22778 22287 23266 22293
rect 22778 22253 22790 22287
rect 23254 22253 23266 22287
rect 22778 22247 23266 22253
rect 22992 22192 23052 22247
rect 23498 22192 23558 22346
rect 24518 22346 24532 22370
rect 24566 22370 24572 22922
rect 25536 22922 25596 23908
rect 26050 23021 26110 23912
rect 26584 23722 26648 24120
rect 27604 24120 27618 24162
rect 27652 24644 27668 24696
rect 28622 24696 28682 24842
rect 29136 24795 29196 25157
rect 29640 25106 29700 25256
rect 30658 25256 30672 25292
rect 30706 25804 30718 25832
rect 31680 25832 31740 26392
rect 32696 26392 32708 26432
rect 32742 26938 32756 26968
rect 33716 26968 33776 27130
rect 32742 26432 32748 26938
rect 33716 26922 33726 26968
rect 32742 26392 32756 26432
rect 32160 26339 32220 26351
rect 31972 26333 32460 26339
rect 31972 26299 31984 26333
rect 32448 26299 32460 26333
rect 31972 26293 32460 26299
rect 32160 25931 32220 26293
rect 32696 26246 32756 26392
rect 33720 26392 33726 26922
rect 33760 26922 33776 26968
rect 33760 26392 33766 26922
rect 33720 26380 33766 26392
rect 32990 26333 33478 26339
rect 32990 26299 33002 26333
rect 33466 26299 33478 26333
rect 32990 26293 33478 26299
rect 32690 26186 32696 26246
rect 32756 26186 32762 26246
rect 33828 26186 33834 26246
rect 33894 26186 33900 26246
rect 32700 25970 33770 26030
rect 31972 25925 32460 25931
rect 31972 25891 31984 25925
rect 32448 25891 32460 25925
rect 31972 25885 32460 25891
rect 30706 25292 30712 25804
rect 31680 25796 31690 25832
rect 30706 25256 30718 25292
rect 31684 25288 31690 25796
rect 30136 25203 30196 25215
rect 29936 25197 30424 25203
rect 29936 25163 29948 25197
rect 30412 25163 30424 25197
rect 29936 25157 30424 25163
rect 29634 25046 29640 25106
rect 29700 25046 29706 25106
rect 28918 24789 29406 24795
rect 28918 24755 28930 24789
rect 29394 24755 29406 24789
rect 28918 24749 29406 24755
rect 29136 24748 29196 24749
rect 28622 24660 28636 24696
rect 27652 24162 27658 24644
rect 27652 24160 27664 24162
rect 27652 24120 27668 24160
rect 26882 24061 27370 24067
rect 26882 24027 26894 24061
rect 27358 24027 27370 24061
rect 26882 24021 27370 24027
rect 27078 23972 27138 23978
rect 27604 23972 27668 24120
rect 28630 24120 28636 24660
rect 28670 24660 28682 24696
rect 29640 24696 29700 25046
rect 30136 24795 30196 25157
rect 30658 24902 30718 25256
rect 31674 25256 31690 25288
rect 31724 25796 31740 25832
rect 32700 25832 32760 25970
rect 33206 25931 33266 25970
rect 32990 25925 33478 25931
rect 32990 25891 33002 25925
rect 33466 25891 33478 25925
rect 32990 25885 33478 25891
rect 32700 25804 32708 25832
rect 31724 25288 31730 25796
rect 31724 25286 31734 25288
rect 32702 25286 32708 25804
rect 31724 25256 31738 25286
rect 31162 25203 31222 25211
rect 30954 25197 31442 25203
rect 30954 25163 30966 25197
rect 31430 25163 31442 25197
rect 30954 25157 31442 25163
rect 30652 24842 30658 24902
rect 30718 24842 30724 24902
rect 31162 24795 31222 25157
rect 31674 25104 31738 25256
rect 32696 25256 32708 25286
rect 32742 25804 32760 25832
rect 33710 25832 33770 25970
rect 32742 25286 32748 25804
rect 33710 25798 33726 25832
rect 32742 25256 32756 25286
rect 32160 25203 32220 25209
rect 31972 25197 32460 25203
rect 31972 25163 31984 25197
rect 32448 25163 32460 25197
rect 31972 25157 32460 25163
rect 31668 25044 31674 25104
rect 31734 25044 31740 25104
rect 29936 24789 30424 24795
rect 29936 24755 29948 24789
rect 30412 24755 30424 24789
rect 29936 24749 30424 24755
rect 30954 24789 31442 24795
rect 30954 24755 30966 24789
rect 31430 24755 31442 24789
rect 30954 24749 31442 24755
rect 31162 24748 31222 24749
rect 28670 24120 28676 24660
rect 29640 24642 29654 24696
rect 29648 24150 29654 24642
rect 28630 24108 28676 24120
rect 29640 24120 29654 24150
rect 29688 24642 29700 24696
rect 30666 24696 30712 24708
rect 29688 24150 29694 24642
rect 30666 24154 30672 24696
rect 29688 24148 29700 24150
rect 29688 24120 29704 24148
rect 27900 24061 28388 24067
rect 27900 24027 27912 24061
rect 28376 24027 28388 24061
rect 27900 24021 28388 24027
rect 28918 24061 29406 24067
rect 28918 24027 28930 24061
rect 29394 24027 29406 24061
rect 28918 24021 29406 24027
rect 26578 23658 26584 23722
rect 26648 23658 26654 23722
rect 27078 23021 27138 23912
rect 27572 23968 27668 23972
rect 27572 23966 27604 23968
rect 27664 23908 27670 23968
rect 28100 23962 28160 23968
rect 25832 23015 26320 23021
rect 25832 22981 25844 23015
rect 26308 22981 26320 23015
rect 25832 22975 26320 22981
rect 26850 23015 27338 23021
rect 26850 22981 26862 23015
rect 27326 22981 27338 23015
rect 26850 22975 27338 22981
rect 24566 22346 24578 22370
rect 23796 22287 24284 22293
rect 23796 22253 23808 22287
rect 24272 22253 24284 22287
rect 23796 22247 24284 22253
rect 24012 22192 24072 22247
rect 24518 22192 24578 22346
rect 25536 22346 25550 22922
rect 25584 22346 25596 22922
rect 26562 22922 26608 22934
rect 26562 22372 26568 22922
rect 24814 22287 25302 22293
rect 24814 22253 24826 22287
rect 25290 22253 25302 22287
rect 24814 22247 25302 22253
rect 25022 22192 25082 22247
rect 25536 22192 25596 22346
rect 26552 22346 26568 22372
rect 26602 22372 26608 22922
rect 27572 22922 27632 23906
rect 28100 23021 28160 23902
rect 28588 23966 28648 23972
rect 27868 23015 28356 23021
rect 27868 22981 27880 23015
rect 28344 22981 28356 23015
rect 27868 22975 28356 22981
rect 28100 22974 28160 22975
rect 26602 22346 26612 22372
rect 25832 22287 26320 22293
rect 25832 22253 25844 22287
rect 26308 22253 26320 22287
rect 25832 22247 26320 22253
rect 26044 22192 26104 22247
rect 26552 22192 26612 22346
rect 27572 22346 27586 22922
rect 27620 22346 27632 22922
rect 26850 22287 27338 22293
rect 26850 22253 26862 22287
rect 27326 22253 27338 22287
rect 26850 22247 27338 22253
rect 27066 22192 27126 22247
rect 27572 22192 27632 22346
rect 28588 22922 28648 23906
rect 29100 23962 29160 23968
rect 29640 23966 29704 24120
rect 30656 24120 30672 24154
rect 30706 24154 30712 24696
rect 31674 24696 31738 25044
rect 32160 24795 32220 25157
rect 32696 25008 32756 25256
rect 33720 25256 33726 25798
rect 33760 25798 33770 25832
rect 33760 25256 33766 25798
rect 33720 25244 33766 25256
rect 32990 25197 33478 25203
rect 32990 25163 33002 25197
rect 33466 25163 33478 25197
rect 32990 25157 33478 25163
rect 32690 24948 32696 25008
rect 32756 24948 32762 25008
rect 32698 24894 32758 24896
rect 32698 24834 33770 24894
rect 31972 24789 32460 24795
rect 31972 24755 31984 24789
rect 32448 24755 32460 24789
rect 31972 24749 32460 24755
rect 32160 24746 32220 24749
rect 31674 24650 31690 24696
rect 30706 24120 30720 24154
rect 31684 24150 31690 24650
rect 29936 24061 30424 24067
rect 29936 24027 29948 24061
rect 30412 24027 30424 24061
rect 29936 24021 30424 24027
rect 29634 23906 29640 23966
rect 29700 23906 29706 23966
rect 29100 23021 29160 23902
rect 30656 23860 30720 24120
rect 31674 24120 31690 24150
rect 31724 24650 31738 24696
rect 32698 24696 32758 24834
rect 33202 24795 33262 24834
rect 32990 24789 33478 24795
rect 32990 24755 33002 24789
rect 33466 24755 33478 24789
rect 32990 24749 33478 24755
rect 32698 24670 32708 24696
rect 31724 24150 31730 24650
rect 32702 24150 32708 24670
rect 31724 24148 31734 24150
rect 31724 24120 31738 24148
rect 30954 24061 31442 24067
rect 30954 24027 30966 24061
rect 31430 24027 31442 24061
rect 30954 24021 31442 24027
rect 31674 23966 31738 24120
rect 32692 24120 32708 24150
rect 32742 24670 32758 24696
rect 33710 24696 33770 24834
rect 32742 24150 32748 24670
rect 33710 24646 33726 24696
rect 32742 24120 32756 24150
rect 31972 24061 32460 24067
rect 31972 24027 31984 24061
rect 32448 24027 32460 24061
rect 31972 24021 32460 24027
rect 31668 23906 31674 23966
rect 31734 23906 31740 23966
rect 30650 23796 30656 23860
rect 30720 23796 30726 23860
rect 32692 23722 32756 24120
rect 33720 24120 33726 24646
rect 33760 24646 33770 24696
rect 33760 24120 33766 24646
rect 33720 24108 33766 24120
rect 32990 24061 33478 24067
rect 32990 24027 33002 24061
rect 33466 24027 33478 24061
rect 32990 24021 33478 24027
rect 32686 23658 32692 23722
rect 32756 23658 32762 23722
rect 32664 23442 32724 23448
rect 32664 23140 32724 23382
rect 33834 23436 33894 26186
rect 33834 23370 33894 23376
rect 29604 23076 29610 23136
rect 29670 23076 29676 23136
rect 31638 23076 31644 23136
rect 31704 23076 31710 23136
rect 32664 23080 33740 23140
rect 28886 23015 29374 23021
rect 28886 22981 28898 23015
rect 29362 22981 29374 23015
rect 28886 22975 29374 22981
rect 29100 22968 29160 22975
rect 28588 22346 28604 22922
rect 28638 22346 28648 22922
rect 29610 22922 29670 23076
rect 29904 23015 30392 23021
rect 29904 22981 29916 23015
rect 30380 22981 30392 23015
rect 29904 22975 30392 22981
rect 30922 23015 31410 23021
rect 30922 22981 30934 23015
rect 31398 22981 31410 23015
rect 30922 22975 31410 22981
rect 29610 22894 29622 22922
rect 27868 22287 28356 22293
rect 27868 22253 27880 22287
rect 28344 22253 28356 22287
rect 27868 22247 28356 22253
rect 28092 22192 28152 22247
rect 28588 22192 28648 22346
rect 29616 22346 29622 22894
rect 29656 22894 29670 22922
rect 30634 22922 30680 22934
rect 29656 22346 29662 22894
rect 30634 22370 30640 22922
rect 29616 22334 29662 22346
rect 30626 22346 30640 22370
rect 30674 22370 30680 22922
rect 31644 22922 31704 23076
rect 31940 23015 32428 23021
rect 31940 22981 31952 23015
rect 32416 22981 32428 23015
rect 31940 22975 32428 22981
rect 31644 22898 31658 22922
rect 30674 22346 30686 22370
rect 28886 22287 29374 22293
rect 28886 22253 28898 22287
rect 29362 22253 29374 22287
rect 28886 22247 29374 22253
rect 29904 22287 30392 22293
rect 29904 22253 29916 22287
rect 30380 22253 30392 22287
rect 29904 22247 30392 22253
rect 29104 22192 29164 22247
rect 22476 22128 22482 22188
rect 22542 22128 22548 22188
rect 22992 22132 29164 22192
rect 23498 22032 23558 22132
rect 28588 22032 28648 22132
rect 23498 21972 28648 22032
rect 21760 21759 22248 21765
rect 21760 21725 21772 21759
rect 22236 21725 22248 21759
rect 21760 21719 22248 21725
rect 22778 21759 23266 21765
rect 22778 21725 22790 21759
rect 23254 21725 23266 21759
rect 22778 21719 23266 21725
rect 21466 21644 21478 21666
rect 20494 21090 20508 21116
rect 19910 21037 19970 21038
rect 19724 21031 20212 21037
rect 19724 20997 19736 21031
rect 20200 20997 20212 21031
rect 19724 20991 20212 20997
rect 18414 20872 19490 20932
rect 18412 20570 19488 20630
rect 18412 20410 18472 20570
rect 18926 20509 18986 20570
rect 18706 20503 19194 20509
rect 18706 20469 18718 20503
rect 19182 20469 19194 20503
rect 18706 20463 19194 20469
rect 18412 20376 18424 20410
rect 18418 19834 18424 20376
rect 18458 20376 18472 20410
rect 19428 20410 19488 20570
rect 19910 20509 19970 20991
rect 20448 20828 20508 21090
rect 21472 21090 21478 21644
rect 21512 21644 21526 21666
rect 22490 21666 22536 21678
rect 21512 21090 21518 21644
rect 22490 21120 22496 21666
rect 21472 21078 21518 21090
rect 22484 21090 22496 21120
rect 22530 21120 22536 21666
rect 23498 21666 23558 21972
rect 24516 21820 24522 21880
rect 24582 21820 24588 21880
rect 25026 21834 26084 21894
rect 23796 21759 24284 21765
rect 23796 21725 23808 21759
rect 24272 21725 24284 21759
rect 23796 21719 24284 21725
rect 23498 21622 23514 21666
rect 23508 21120 23514 21622
rect 22530 21090 22544 21120
rect 20948 21037 21008 21038
rect 21954 21037 22014 21038
rect 20742 21031 21230 21037
rect 20742 20997 20754 21031
rect 21218 20997 21230 21031
rect 20742 20991 21230 20997
rect 21760 21031 22248 21037
rect 21760 20997 21772 21031
rect 22236 20997 22248 21031
rect 21760 20991 22248 20997
rect 20448 20762 20508 20768
rect 20442 20564 20448 20624
rect 20508 20564 20514 20624
rect 19724 20503 20212 20509
rect 19724 20469 19736 20503
rect 20200 20469 20212 20503
rect 19724 20463 20212 20469
rect 19428 20388 19442 20410
rect 18458 19834 18464 20376
rect 19436 19862 19442 20388
rect 18418 19822 18464 19834
rect 19430 19834 19442 19862
rect 19476 20388 19488 20410
rect 20448 20410 20508 20564
rect 20948 20509 21008 20991
rect 21954 20509 22014 20991
rect 22484 20828 22544 21090
rect 23500 21090 23514 21120
rect 23548 21622 23558 21666
rect 24522 21666 24582 21820
rect 25026 21765 25086 21834
rect 26026 21796 26084 21834
rect 26550 21820 26556 21880
rect 26616 21820 26622 21880
rect 26026 21765 26086 21796
rect 24814 21759 25302 21765
rect 24814 21725 24826 21759
rect 25290 21725 25302 21759
rect 24814 21719 25302 21725
rect 25832 21759 26320 21765
rect 25832 21725 25844 21759
rect 26308 21725 26320 21759
rect 25832 21719 26320 21725
rect 24522 21638 24532 21666
rect 23548 21120 23554 21622
rect 23548 21090 23560 21120
rect 22778 21031 23266 21037
rect 22778 20997 22790 21031
rect 23254 20997 23266 21031
rect 22778 20991 23266 20997
rect 23004 20936 23064 20991
rect 23500 20936 23560 21090
rect 24526 21090 24532 21638
rect 24566 21638 24582 21666
rect 25544 21666 25590 21678
rect 24566 21090 24572 21638
rect 25544 21114 25550 21666
rect 24526 21078 24572 21090
rect 25538 21090 25550 21114
rect 25584 21114 25590 21666
rect 26556 21666 26616 21820
rect 26850 21759 27338 21765
rect 26850 21725 26862 21759
rect 27326 21725 27338 21759
rect 26850 21719 27338 21725
rect 27868 21759 28356 21765
rect 27868 21725 27880 21759
rect 28344 21725 28356 21759
rect 27868 21719 28356 21725
rect 26556 21636 26568 21666
rect 26562 21118 26568 21636
rect 25584 21090 25598 21114
rect 23796 21031 24284 21037
rect 23796 20997 23808 21031
rect 24272 20997 24284 21031
rect 23796 20991 24284 20997
rect 24814 21031 25302 21037
rect 24814 20997 24826 21031
rect 25290 20997 25302 21031
rect 24814 20991 25302 20997
rect 24016 20936 24076 20991
rect 23004 20876 24076 20936
rect 22478 20768 22484 20828
rect 22544 20768 22550 20828
rect 22476 20666 22482 20726
rect 22542 20666 22548 20726
rect 22482 20624 22542 20666
rect 22476 20564 22482 20624
rect 22542 20564 22548 20624
rect 20742 20503 21230 20509
rect 20742 20469 20754 20503
rect 21218 20469 21230 20503
rect 20742 20463 21230 20469
rect 21760 20503 22248 20509
rect 21760 20469 21772 20503
rect 22236 20469 22248 20503
rect 21760 20463 22248 20469
rect 19476 19862 19482 20388
rect 20448 20386 20460 20410
rect 19476 19834 19490 19862
rect 18706 19775 19194 19781
rect 18706 19741 18718 19775
rect 19182 19741 19194 19775
rect 18706 19735 19194 19741
rect 19430 19676 19490 19834
rect 20454 19834 20460 20386
rect 20494 20386 20508 20410
rect 21472 20410 21518 20422
rect 20494 19834 20500 20386
rect 21472 19858 21478 20410
rect 20454 19822 20500 19834
rect 21466 19834 21478 19858
rect 21512 19858 21518 20410
rect 22482 20410 22542 20564
rect 22778 20503 23266 20509
rect 22778 20469 22790 20503
rect 23254 20469 23266 20503
rect 22778 20463 23266 20469
rect 22482 20382 22496 20410
rect 21512 19834 21526 19858
rect 19922 19781 19982 19788
rect 20960 19781 21020 19788
rect 19724 19775 20212 19781
rect 19724 19741 19736 19775
rect 20200 19741 20212 19775
rect 19724 19735 20212 19741
rect 20742 19775 21230 19781
rect 20742 19741 20754 19775
rect 21218 19741 21230 19775
rect 20742 19735 21230 19741
rect 19424 19616 19430 19676
rect 19490 19616 19496 19676
rect 18256 19408 18262 19468
rect 18322 19408 18328 19468
rect 18412 19310 19488 19370
rect 18412 19154 18472 19310
rect 18926 19253 18986 19310
rect 18706 19247 19194 19253
rect 18706 19213 18718 19247
rect 19182 19213 19194 19247
rect 18706 19207 19194 19213
rect 18412 19116 18424 19154
rect 18418 18578 18424 19116
rect 18458 19116 18472 19154
rect 19428 19154 19488 19310
rect 19922 19253 19982 19735
rect 20438 19306 20444 19366
rect 20504 19306 20510 19366
rect 19724 19247 20212 19253
rect 19724 19213 19736 19247
rect 20200 19213 20212 19247
rect 19724 19207 20212 19213
rect 19428 19128 19442 19154
rect 18458 18578 18464 19116
rect 19436 18604 19442 19128
rect 18418 18566 18464 18578
rect 19426 18578 19442 18604
rect 19476 19128 19488 19154
rect 20444 19154 20504 19306
rect 20960 19253 21020 19735
rect 21466 19676 21526 19834
rect 22490 19834 22496 20382
rect 22530 20382 22542 20410
rect 23500 20410 23560 20876
rect 24512 20872 24518 20932
rect 24578 20872 24584 20932
rect 23796 20503 24284 20509
rect 23796 20469 23808 20503
rect 24272 20469 24284 20503
rect 23796 20463 24284 20469
rect 22530 19834 22536 20382
rect 23500 20372 23514 20410
rect 23508 19868 23514 20372
rect 22490 19822 22536 19834
rect 23498 19834 23514 19868
rect 23548 20372 23560 20410
rect 24518 20410 24578 20872
rect 25020 20509 25080 20991
rect 25538 20932 25598 21090
rect 26556 21090 26568 21118
rect 26602 21636 26616 21666
rect 27580 21666 27626 21678
rect 26602 21118 26608 21636
rect 27580 21118 27586 21666
rect 26602 21090 26616 21118
rect 26050 21037 26110 21044
rect 25832 21031 26320 21037
rect 25832 20997 25844 21031
rect 26308 20997 26320 21031
rect 25832 20991 26320 20997
rect 25532 20872 25538 20932
rect 25598 20872 25604 20932
rect 25532 20566 25538 20626
rect 25598 20566 25604 20626
rect 24814 20503 25302 20509
rect 24814 20469 24826 20503
rect 25290 20469 25302 20503
rect 24814 20463 25302 20469
rect 25020 20458 25080 20463
rect 24518 20386 24532 20410
rect 23548 19868 23554 20372
rect 23548 19834 23558 19868
rect 24526 19864 24532 20386
rect 21966 19781 22026 19788
rect 21760 19775 22248 19781
rect 21760 19741 21772 19775
rect 22236 19741 22248 19775
rect 21760 19735 22248 19741
rect 22778 19775 23266 19781
rect 22778 19741 22790 19775
rect 23254 19741 23266 19775
rect 22778 19735 23266 19741
rect 21460 19616 21466 19676
rect 21526 19616 21532 19676
rect 21466 19568 21526 19616
rect 21460 19508 21466 19568
rect 21526 19508 21532 19568
rect 21966 19518 22026 19735
rect 23002 19684 23062 19735
rect 23498 19684 23558 19834
rect 24520 19834 24532 19864
rect 24566 20386 24578 20410
rect 25538 20410 25598 20566
rect 26050 20509 26110 20991
rect 26556 20626 26616 21090
rect 27574 21090 27586 21118
rect 27620 21118 27626 21666
rect 28588 21666 28648 21972
rect 29606 21820 29612 21880
rect 29672 21820 29678 21880
rect 28886 21759 29374 21765
rect 28886 21725 28898 21759
rect 29362 21725 29374 21759
rect 28886 21719 29374 21725
rect 28588 21646 28604 21666
rect 28598 21118 28604 21646
rect 27620 21090 27634 21118
rect 27062 21037 27122 21044
rect 26850 21031 27338 21037
rect 26850 20997 26862 21031
rect 27326 20997 27338 21031
rect 26850 20991 27338 20997
rect 26550 20566 26556 20626
rect 26616 20566 26622 20626
rect 27062 20509 27122 20991
rect 27574 20932 27634 21090
rect 28588 21090 28604 21118
rect 28638 21646 28648 21666
rect 29612 21666 29672 21820
rect 30112 21765 30172 22247
rect 30626 22188 30686 22346
rect 31652 22346 31658 22898
rect 31692 22898 31704 22922
rect 32664 22922 32724 23080
rect 33178 23021 33238 23080
rect 32958 23015 33446 23021
rect 32958 22981 32970 23015
rect 33434 22981 33446 23015
rect 32958 22975 33446 22981
rect 31692 22346 31698 22898
rect 32664 22886 32676 22922
rect 32670 22374 32676 22886
rect 31652 22334 31698 22346
rect 32662 22346 32676 22374
rect 32710 22886 32724 22922
rect 33680 22922 33740 23080
rect 34082 23076 34088 23136
rect 34148 23076 34154 23136
rect 33680 22898 33694 22922
rect 32710 22374 32716 22886
rect 32710 22346 32722 22374
rect 32142 22293 32202 22299
rect 30922 22287 31410 22293
rect 30922 22253 30934 22287
rect 31398 22253 31410 22287
rect 30922 22247 31410 22253
rect 31940 22287 32428 22293
rect 31940 22253 31952 22287
rect 32416 22253 32428 22287
rect 31940 22247 32428 22253
rect 30620 22128 30626 22188
rect 30686 22128 30692 22188
rect 31136 21765 31196 22247
rect 31640 21820 31646 21880
rect 31706 21820 31712 21880
rect 29904 21759 30392 21765
rect 29904 21725 29916 21759
rect 30380 21725 30392 21759
rect 29904 21719 30392 21725
rect 30922 21759 31410 21765
rect 30922 21725 30934 21759
rect 31398 21725 31410 21759
rect 30922 21719 31410 21725
rect 28638 21118 28644 21646
rect 29612 21638 29622 21666
rect 28638 21090 28648 21118
rect 27868 21031 28356 21037
rect 27868 20997 27880 21031
rect 28344 20997 28356 21031
rect 27868 20991 28356 20997
rect 28092 20934 28152 20991
rect 28588 20934 28648 21090
rect 29616 21090 29622 21638
rect 29656 21638 29672 21666
rect 30634 21666 30680 21678
rect 29656 21090 29662 21638
rect 30634 21126 30640 21666
rect 29616 21078 29662 21090
rect 30624 21090 30640 21126
rect 30674 21126 30680 21666
rect 31646 21666 31706 21820
rect 32142 21765 32202 22247
rect 32662 22188 32722 22346
rect 33688 22346 33694 22898
rect 33728 22898 33740 22922
rect 33728 22346 33734 22898
rect 33688 22334 33734 22346
rect 32958 22287 33446 22293
rect 32958 22253 32970 22287
rect 33434 22253 33446 22287
rect 32958 22247 33446 22253
rect 32656 22128 32662 22188
rect 32722 22128 32728 22188
rect 33922 21934 33928 21994
rect 33988 21934 33994 21994
rect 32664 21826 33740 21886
rect 31940 21759 32428 21765
rect 31940 21725 31952 21759
rect 32416 21725 32428 21759
rect 31940 21719 32428 21725
rect 31646 21642 31658 21666
rect 30674 21090 30684 21126
rect 31652 21118 31658 21642
rect 30106 21037 30166 21038
rect 28886 21031 29374 21037
rect 28886 20997 28898 21031
rect 29362 20997 29374 21031
rect 28886 20991 29374 20997
rect 29904 21031 30392 21037
rect 29904 20997 29916 21031
rect 30380 20997 30392 21031
rect 29904 20991 30392 20997
rect 29104 20934 29164 20991
rect 27568 20872 27574 20932
rect 27634 20872 27640 20932
rect 28092 20874 29164 20934
rect 27566 20566 27572 20626
rect 27632 20566 27638 20626
rect 25832 20503 26320 20509
rect 25832 20469 25844 20503
rect 26308 20469 26320 20503
rect 25832 20463 26320 20469
rect 26850 20503 27338 20509
rect 26850 20469 26862 20503
rect 27326 20469 27338 20503
rect 26850 20463 27338 20469
rect 25538 20388 25550 20410
rect 24566 19864 24572 20386
rect 24566 19834 24580 19864
rect 23796 19775 24284 19781
rect 23796 19741 23808 19775
rect 24272 19741 24284 19775
rect 23796 19735 24284 19741
rect 24014 19684 24074 19735
rect 23002 19624 24074 19684
rect 24520 19678 24580 19834
rect 25544 19834 25550 20388
rect 25584 20388 25598 20410
rect 26562 20410 26608 20422
rect 25584 19834 25590 20388
rect 26562 19860 26568 20410
rect 25544 19822 25590 19834
rect 26556 19834 26568 19860
rect 26602 19860 26608 20410
rect 27572 20410 27632 20566
rect 27868 20503 28356 20509
rect 27868 20469 27880 20503
rect 28344 20469 28356 20503
rect 27868 20463 28356 20469
rect 27572 20384 27586 20410
rect 26602 19834 26616 19860
rect 26046 19781 26106 19784
rect 24814 19775 25302 19781
rect 24814 19741 24826 19775
rect 25290 19741 25302 19775
rect 24814 19735 25302 19741
rect 25832 19775 26320 19781
rect 25832 19741 25844 19775
rect 26308 19741 26320 19775
rect 25832 19735 26320 19741
rect 21966 19458 22742 19518
rect 21966 19253 22026 19458
rect 22682 19372 22742 19458
rect 22472 19306 22478 19366
rect 22538 19306 22544 19366
rect 22676 19312 22682 19372
rect 22742 19312 22748 19372
rect 20742 19247 21230 19253
rect 20742 19213 20754 19247
rect 21218 19213 21230 19247
rect 20742 19207 21230 19213
rect 21760 19247 22248 19253
rect 21760 19213 21772 19247
rect 22236 19213 22248 19247
rect 21760 19207 22248 19213
rect 20444 19128 20460 19154
rect 19476 18604 19482 19128
rect 19476 18578 19486 18604
rect 18706 18519 19194 18525
rect 18706 18485 18718 18519
rect 19182 18485 19194 18519
rect 18706 18479 19194 18485
rect 19426 18418 19486 18578
rect 20454 18578 20460 19128
rect 20494 19128 20504 19154
rect 21472 19154 21518 19166
rect 20494 18578 20500 19128
rect 21472 18600 21478 19154
rect 20454 18566 20500 18578
rect 21462 18578 21478 18600
rect 21512 18600 21518 19154
rect 22478 19154 22538 19306
rect 22778 19247 23266 19253
rect 22778 19213 22790 19247
rect 23254 19213 23266 19247
rect 22778 19207 23266 19213
rect 22478 19124 22496 19154
rect 22490 18614 22496 19124
rect 21512 18578 21522 18600
rect 19724 18519 20212 18525
rect 19724 18485 19736 18519
rect 20200 18485 20212 18519
rect 19724 18479 20212 18485
rect 20742 18519 21230 18525
rect 20742 18485 20754 18519
rect 21218 18485 21230 18519
rect 20742 18479 21230 18485
rect 19420 18358 19426 18418
rect 19486 18358 19492 18418
rect 19934 18304 19994 18479
rect 20958 18304 21018 18479
rect 21462 18418 21522 18578
rect 22484 18578 22496 18614
rect 22530 19124 22538 19154
rect 23498 19154 23558 19624
rect 24514 19618 24520 19678
rect 24580 19618 24586 19678
rect 25030 19546 25090 19735
rect 26046 19546 26106 19735
rect 26556 19678 26616 19834
rect 27580 19834 27586 20384
rect 27620 20384 27632 20410
rect 28588 20410 28648 20874
rect 29602 20768 29608 20828
rect 29668 20768 29674 20828
rect 28886 20503 29374 20509
rect 28886 20469 28898 20503
rect 29362 20469 29374 20503
rect 28886 20463 29374 20469
rect 27620 19834 27626 20384
rect 28588 20380 28604 20410
rect 28598 19866 28604 20380
rect 27580 19822 27626 19834
rect 28586 19834 28604 19866
rect 28638 20380 28648 20410
rect 29608 20410 29668 20768
rect 30106 20509 30166 20991
rect 30470 20886 30476 20946
rect 30536 20886 30542 20946
rect 30476 20626 30536 20886
rect 30624 20836 30684 21090
rect 31644 21090 31658 21118
rect 31692 21642 31706 21666
rect 32664 21666 32724 21826
rect 33178 21765 33238 21826
rect 32958 21759 33446 21765
rect 32958 21725 32970 21759
rect 33434 21725 33446 21759
rect 32958 21719 33446 21725
rect 31692 21118 31698 21642
rect 32664 21632 32676 21666
rect 32670 21130 32676 21632
rect 31692 21090 31704 21118
rect 31130 21037 31190 21038
rect 30922 21031 31410 21037
rect 30922 20997 30934 21031
rect 31398 20997 31410 21031
rect 30922 20991 31410 20997
rect 30618 20776 30624 20836
rect 30684 20776 30690 20836
rect 30470 20566 30476 20626
rect 30536 20566 30542 20626
rect 30622 20568 30628 20628
rect 30688 20568 30694 20628
rect 29904 20503 30392 20509
rect 29904 20469 29916 20503
rect 30380 20469 30392 20503
rect 29904 20463 30392 20469
rect 28638 19866 28644 20380
rect 29608 20378 29622 20410
rect 29616 19866 29622 20378
rect 28638 19834 28646 19866
rect 26850 19775 27338 19781
rect 26850 19741 26862 19775
rect 27326 19741 27338 19775
rect 26850 19735 27338 19741
rect 27868 19775 28356 19781
rect 27868 19741 27880 19775
rect 28344 19741 28356 19775
rect 27868 19735 28356 19741
rect 26550 19618 26556 19678
rect 26616 19618 26622 19678
rect 27060 19546 27120 19735
rect 28090 19682 28150 19735
rect 28586 19682 28646 19834
rect 29610 19834 29622 19866
rect 29656 20378 29668 20410
rect 30628 20410 30688 20568
rect 31130 20509 31190 20991
rect 31644 20726 31704 21090
rect 32664 21090 32676 21130
rect 32710 21632 32724 21666
rect 33680 21666 33740 21826
rect 33680 21644 33694 21666
rect 32710 21130 32716 21632
rect 32710 21090 32724 21130
rect 32136 21037 32196 21044
rect 31940 21031 32428 21037
rect 31940 20997 31952 21031
rect 32416 20997 32428 21031
rect 31940 20991 32428 20997
rect 31638 20666 31644 20726
rect 31704 20666 31710 20726
rect 32136 20509 32196 20991
rect 32664 20836 32724 21090
rect 33688 21090 33694 21644
rect 33728 21644 33740 21666
rect 33728 21090 33734 21644
rect 33688 21078 33734 21090
rect 32958 21031 33446 21037
rect 32958 20997 32970 21031
rect 33434 20997 33446 21031
rect 32958 20991 33446 20997
rect 32658 20776 32664 20836
rect 32724 20776 32730 20836
rect 33790 20776 33796 20836
rect 33856 20776 33862 20836
rect 32656 20568 32662 20628
rect 32722 20568 32728 20628
rect 30922 20503 31410 20509
rect 30922 20469 30934 20503
rect 31398 20469 31410 20503
rect 30922 20463 31410 20469
rect 31940 20503 32428 20509
rect 31940 20469 31952 20503
rect 32416 20469 32428 20503
rect 31940 20463 32428 20469
rect 30628 20390 30640 20410
rect 29656 19866 29662 20378
rect 29656 19834 29670 19866
rect 28886 19775 29374 19781
rect 28886 19741 28898 19775
rect 29362 19741 29374 19775
rect 28886 19735 29374 19741
rect 29102 19682 29162 19735
rect 28090 19622 29162 19682
rect 29610 19680 29670 19834
rect 30634 19834 30640 20390
rect 30674 20390 30688 20410
rect 31652 20410 31698 20422
rect 30674 19834 30680 20390
rect 31652 19862 31658 20410
rect 30634 19822 30680 19834
rect 31646 19834 31658 19862
rect 31692 19862 31698 20410
rect 32662 20410 32722 20568
rect 32958 20503 33446 20509
rect 32958 20469 32970 20503
rect 33434 20469 33446 20503
rect 32958 20463 33446 20469
rect 32662 20386 32676 20410
rect 32670 19870 32676 20386
rect 31692 19834 31706 19862
rect 30118 19781 30178 19788
rect 31142 19781 31202 19788
rect 29904 19775 30392 19781
rect 29904 19741 29916 19775
rect 30380 19741 30392 19775
rect 29904 19735 30392 19741
rect 30922 19775 31410 19781
rect 30922 19741 30934 19775
rect 31398 19741 31410 19775
rect 30922 19735 31410 19741
rect 25030 19486 27844 19546
rect 24516 19372 24576 19378
rect 25030 19372 25090 19486
rect 24576 19312 25090 19372
rect 24516 19306 24576 19312
rect 25530 19308 25536 19368
rect 25596 19308 25602 19368
rect 27564 19308 27570 19368
rect 27630 19308 27636 19368
rect 27784 19364 27844 19486
rect 23796 19247 24284 19253
rect 23796 19213 23808 19247
rect 24272 19213 24284 19247
rect 23796 19207 24284 19213
rect 24814 19247 25302 19253
rect 24814 19213 24826 19247
rect 25290 19213 25302 19247
rect 24814 19207 25302 19213
rect 22530 18614 22536 19124
rect 23498 19096 23514 19154
rect 22530 18578 22544 18614
rect 23508 18610 23514 19096
rect 21760 18519 22248 18525
rect 21760 18485 21772 18519
rect 22236 18485 22248 18519
rect 21760 18479 22248 18485
rect 21456 18358 21462 18418
rect 21522 18358 21528 18418
rect 21964 18304 22024 18479
rect 18124 18228 18130 18288
rect 18190 18228 18196 18288
rect 19934 18244 22024 18304
rect 13054 18088 13060 18148
rect 13120 18088 13126 18148
rect 12904 18042 12964 18048
rect 18130 18042 18190 18228
rect 12964 17982 18190 18042
rect 12904 17976 12964 17982
rect 12134 17924 12194 17930
rect 19934 17924 19994 18244
rect 21964 17994 22024 18244
rect 22484 18148 22544 18578
rect 23498 18578 23514 18610
rect 23548 19096 23558 19154
rect 24526 19154 24572 19166
rect 23548 18610 23554 19096
rect 24526 18622 24532 19154
rect 23548 18578 23558 18610
rect 22778 18519 23266 18525
rect 22778 18485 22790 18519
rect 23254 18485 23266 18519
rect 22778 18479 23266 18485
rect 23002 18424 23062 18479
rect 23498 18424 23558 18578
rect 24520 18578 24532 18622
rect 24566 18622 24572 19154
rect 25536 19154 25596 19308
rect 25832 19247 26320 19253
rect 25832 19213 25844 19247
rect 26308 19213 26320 19247
rect 25832 19207 26320 19213
rect 26850 19247 27338 19253
rect 26850 19213 26862 19247
rect 27326 19213 27338 19247
rect 26850 19207 27338 19213
rect 25536 19130 25550 19154
rect 24566 18578 24580 18622
rect 25544 18602 25550 19130
rect 23796 18519 24284 18525
rect 23796 18485 23808 18519
rect 24272 18485 24284 18519
rect 23796 18479 24284 18485
rect 24014 18424 24074 18479
rect 24520 18424 24580 18578
rect 25536 18578 25550 18602
rect 25584 19130 25596 19154
rect 26562 19154 26608 19166
rect 25584 18602 25590 19130
rect 26562 18616 26568 19154
rect 25584 18578 25596 18602
rect 24814 18519 25302 18525
rect 24814 18485 24826 18519
rect 25290 18485 25302 18519
rect 24814 18479 25302 18485
rect 25030 18424 25090 18479
rect 25536 18424 25596 18578
rect 26554 18578 26568 18616
rect 26602 18616 26608 19154
rect 27570 19154 27630 19308
rect 27778 19304 27784 19364
rect 27844 19304 27850 19364
rect 27868 19247 28356 19253
rect 27868 19213 27880 19247
rect 28344 19213 28356 19247
rect 27868 19207 28356 19213
rect 27570 19126 27586 19154
rect 26602 18578 26614 18616
rect 27580 18606 27586 19126
rect 25832 18519 26320 18525
rect 25832 18485 25844 18519
rect 26308 18485 26320 18519
rect 25832 18479 26320 18485
rect 26046 18424 26106 18479
rect 26554 18424 26614 18578
rect 27572 18578 27586 18606
rect 27620 19126 27630 19154
rect 28586 19154 28646 19622
rect 29604 19620 29610 19680
rect 29670 19620 29676 19680
rect 30118 19370 30178 19735
rect 30118 19364 30180 19370
rect 30118 19304 30120 19364
rect 30626 19306 30632 19366
rect 30692 19306 30698 19366
rect 30118 19298 30180 19304
rect 30118 19253 30178 19298
rect 28886 19247 29374 19253
rect 28886 19213 28898 19247
rect 29362 19213 29374 19247
rect 28886 19207 29374 19213
rect 29904 19247 30392 19253
rect 29904 19213 29916 19247
rect 30380 19213 30392 19247
rect 29904 19207 30392 19213
rect 27620 18606 27626 19126
rect 28586 19116 28604 19154
rect 28598 18608 28604 19116
rect 27620 18578 27632 18606
rect 26850 18519 27338 18525
rect 26850 18485 26862 18519
rect 27326 18485 27338 18519
rect 26850 18479 27338 18485
rect 27056 18424 27116 18479
rect 27572 18424 27632 18578
rect 28586 18578 28604 18608
rect 28638 19116 28646 19154
rect 29616 19154 29662 19166
rect 28638 18608 28644 19116
rect 28638 18578 28646 18608
rect 29616 18604 29622 19154
rect 27868 18519 28356 18525
rect 27868 18485 27880 18519
rect 28344 18485 28356 18519
rect 27868 18479 28356 18485
rect 28090 18424 28150 18479
rect 28586 18424 28646 18578
rect 29614 18578 29622 18604
rect 29656 18604 29662 19154
rect 30632 19154 30692 19306
rect 31142 19253 31202 19735
rect 31646 19680 31706 19834
rect 32662 19834 32676 19870
rect 32710 20386 32722 20410
rect 33688 20410 33734 20422
rect 32710 19870 32716 20386
rect 32710 19834 32722 19870
rect 33688 19858 33694 20410
rect 32148 19781 32208 19794
rect 31940 19775 32428 19781
rect 31940 19741 31952 19775
rect 32416 19741 32428 19775
rect 31940 19735 32428 19741
rect 31640 19620 31646 19680
rect 31706 19620 31712 19680
rect 32148 19253 32208 19735
rect 32662 19676 32722 19834
rect 33678 19834 33694 19858
rect 33728 19858 33734 20410
rect 33728 19834 33738 19858
rect 32958 19775 33446 19781
rect 32958 19741 32970 19775
rect 33434 19741 33446 19775
rect 32958 19735 33446 19741
rect 33176 19676 33236 19735
rect 33678 19676 33738 19834
rect 32662 19616 33738 19676
rect 33796 19568 33856 20776
rect 33928 20628 33988 21934
rect 33922 20568 33928 20628
rect 33988 20568 33994 20628
rect 33790 19508 33796 19568
rect 33856 19508 33862 19568
rect 32660 19306 32666 19366
rect 32726 19306 32732 19366
rect 30922 19247 31410 19253
rect 30922 19213 30934 19247
rect 31398 19213 31410 19247
rect 30922 19207 31410 19213
rect 31940 19247 32428 19253
rect 31940 19213 31952 19247
rect 32416 19213 32428 19247
rect 31940 19207 32428 19213
rect 30632 19128 30640 19154
rect 29656 18578 29674 18604
rect 28886 18519 29374 18525
rect 28886 18485 28898 18519
rect 29362 18485 29374 18519
rect 28886 18479 29374 18485
rect 29102 18424 29162 18479
rect 23002 18364 29162 18424
rect 29614 18418 29674 18578
rect 30634 18578 30640 19128
rect 30674 19128 30692 19154
rect 31652 19154 31698 19166
rect 30674 18578 30680 19128
rect 31652 18600 31658 19154
rect 30634 18566 30680 18578
rect 31650 18578 31658 18600
rect 31692 18600 31698 19154
rect 32666 19154 32726 19306
rect 32958 19247 33446 19253
rect 32958 19213 32970 19247
rect 33434 19213 33446 19247
rect 32958 19207 33446 19213
rect 32666 19124 32676 19154
rect 32670 18616 32676 19124
rect 31692 18578 31710 18600
rect 30122 18525 30182 18532
rect 29904 18519 30392 18525
rect 29904 18485 29916 18519
rect 30380 18485 30392 18519
rect 29904 18479 30392 18485
rect 30922 18519 31410 18525
rect 30922 18485 30934 18519
rect 31398 18485 31410 18519
rect 30922 18479 31410 18485
rect 29608 18358 29614 18418
rect 29674 18358 29680 18418
rect 30122 18306 30182 18479
rect 31142 18306 31202 18479
rect 31650 18418 31710 18578
rect 32664 18578 32676 18616
rect 32710 19124 32726 19154
rect 33688 19154 33734 19166
rect 32710 18616 32716 19124
rect 32710 18578 32724 18616
rect 33688 18604 33694 19154
rect 31940 18519 32428 18525
rect 31940 18485 31952 18519
rect 32416 18485 32428 18519
rect 31940 18479 32428 18485
rect 31644 18358 31650 18418
rect 31710 18358 31716 18418
rect 32144 18306 32204 18479
rect 32664 18422 32724 18578
rect 33680 18578 33694 18604
rect 33728 18604 33734 19154
rect 33728 18578 33740 18604
rect 32958 18519 33446 18525
rect 32958 18485 32970 18519
rect 33434 18485 33446 18519
rect 32958 18479 33446 18485
rect 33178 18422 33238 18479
rect 33680 18422 33740 18578
rect 32664 18362 33740 18422
rect 30122 18246 32204 18306
rect 22478 18088 22484 18148
rect 22544 18088 22550 18148
rect 30122 17994 30182 18246
rect 34088 18148 34148 23076
rect 35666 18278 35672 27642
rect 35772 18278 35778 27642
rect 47792 27680 48000 27710
rect 47792 27564 47824 27680
rect 47792 25538 48000 27564
rect 48306 27680 48488 27710
rect 48462 27564 48488 27680
rect 48306 25538 48488 27564
rect 65322 27642 65434 28156
rect 66034 27856 66044 28156
rect 89056 27856 89066 28156
rect 47022 25478 49087 25538
rect 47022 23538 47082 25478
rect 47251 25412 47556 25478
rect 47251 25378 47310 25412
rect 47530 25378 47556 25412
rect 47251 25364 47556 25378
rect 47251 25314 47312 25364
rect 47251 25284 47262 25314
rect 47252 25056 47262 25284
rect 47251 24996 47262 25056
rect 47252 24742 47262 24996
rect 47300 25056 47312 25314
rect 47362 25216 47422 25364
rect 47496 25315 47556 25364
rect 47752 25430 47812 25431
rect 48528 25430 48588 25436
rect 47752 25370 48528 25430
rect 47752 25315 47812 25370
rect 48010 25315 48070 25370
rect 48268 25315 48328 25370
rect 48528 25315 48588 25370
rect 48784 25412 49087 25478
rect 48784 25378 48802 25412
rect 49004 25378 49087 25412
rect 48784 25364 49087 25378
rect 48784 25315 48844 25364
rect 47470 25309 47578 25315
rect 47470 25275 47482 25309
rect 47566 25275 47578 25309
rect 47470 25269 47578 25275
rect 47728 25309 47836 25315
rect 47728 25275 47740 25309
rect 47824 25275 47836 25309
rect 47728 25269 47836 25275
rect 47986 25309 48094 25315
rect 47986 25275 47998 25309
rect 48082 25275 48094 25309
rect 47986 25269 48094 25275
rect 48244 25309 48352 25315
rect 48244 25275 48256 25309
rect 48340 25275 48352 25309
rect 48244 25269 48352 25275
rect 48502 25309 48610 25315
rect 48502 25275 48514 25309
rect 48598 25275 48610 25309
rect 48502 25269 48610 25275
rect 48760 25309 48868 25315
rect 48760 25275 48772 25309
rect 48856 25275 48868 25309
rect 48760 25269 48868 25275
rect 47362 25056 47378 25216
rect 47300 24996 47378 25056
rect 47300 24742 47312 24996
rect 47372 24874 47378 24996
rect 47252 24692 47312 24742
rect 47364 24840 47378 24874
rect 47412 24996 47422 25216
rect 47630 25216 47676 25228
rect 47412 24874 47418 24996
rect 47630 24885 47636 25216
rect 47412 24840 47424 24874
rect 47364 24692 47424 24840
rect 47622 24840 47636 24885
rect 47670 24885 47676 25216
rect 47888 25216 47934 25228
rect 47670 24840 47682 24885
rect 47888 24860 47894 25216
rect 47470 24781 47578 24787
rect 47470 24747 47482 24781
rect 47566 24747 47578 24781
rect 47470 24741 47578 24747
rect 47492 24692 47552 24741
rect 47251 24678 47552 24692
rect 47251 24644 47310 24678
rect 47530 24644 47552 24678
rect 47251 24632 47552 24644
rect 47622 24515 47682 24840
rect 47880 24840 47894 24860
rect 47928 24860 47934 25216
rect 48146 25216 48192 25228
rect 48146 24883 48152 25216
rect 47928 24840 47940 24860
rect 47728 24781 47836 24787
rect 47728 24747 47740 24781
rect 47824 24747 47836 24781
rect 47728 24741 47836 24747
rect 47880 24664 47940 24840
rect 48138 24840 48152 24883
rect 48186 24883 48192 25216
rect 48404 25216 48450 25228
rect 48186 24840 48198 24883
rect 48404 24878 48410 25216
rect 47986 24781 48094 24787
rect 47986 24747 47998 24781
rect 48082 24747 48094 24781
rect 47986 24741 48094 24747
rect 47874 24604 47880 24664
rect 47940 24604 47946 24664
rect 47250 24480 47554 24490
rect 47250 24442 47334 24480
rect 47542 24442 47554 24480
rect 47616 24455 47622 24515
rect 47682 24455 47688 24515
rect 47250 24430 47554 24442
rect 47250 24382 47310 24430
rect 47250 24026 47262 24382
rect 47298 24026 47310 24382
rect 47364 24292 47424 24430
rect 47494 24382 47554 24430
rect 47470 24376 47578 24382
rect 47470 24342 47482 24376
rect 47566 24342 47578 24376
rect 47470 24336 47578 24342
rect 47364 24242 47378 24292
rect 47372 24155 47378 24242
rect 47250 23977 47310 24026
rect 47366 24116 47378 24155
rect 47412 24242 47424 24292
rect 47622 24292 47682 24455
rect 47728 24376 47836 24382
rect 47728 24342 47740 24376
rect 47824 24342 47836 24376
rect 47728 24336 47836 24342
rect 47622 24255 47636 24292
rect 47412 24155 47418 24242
rect 47412 24116 47426 24155
rect 47366 23977 47426 24116
rect 47630 24116 47636 24255
rect 47670 24255 47682 24292
rect 47880 24322 47940 24604
rect 48138 24515 48198 24840
rect 48398 24840 48410 24878
rect 48444 24878 48450 25216
rect 48662 25216 48708 25228
rect 48662 24883 48668 25216
rect 48444 24840 48458 24878
rect 48244 24781 48352 24787
rect 48244 24747 48256 24781
rect 48340 24747 48352 24781
rect 48244 24741 48352 24747
rect 48398 24664 48458 24840
rect 48656 24840 48668 24883
rect 48702 24883 48708 25216
rect 48912 25216 48972 25364
rect 48912 24998 48926 25216
rect 48702 24840 48716 24883
rect 48920 24870 48926 24998
rect 48502 24781 48610 24787
rect 48502 24747 48514 24781
rect 48598 24747 48610 24781
rect 48502 24741 48610 24747
rect 48392 24604 48398 24664
rect 48458 24604 48464 24664
rect 48132 24455 48138 24515
rect 48198 24455 48204 24515
rect 47986 24376 48094 24382
rect 47986 24342 47998 24376
rect 48082 24342 48094 24376
rect 47986 24336 48094 24342
rect 47880 24292 47942 24322
rect 47880 24256 47894 24292
rect 47670 24116 47676 24255
rect 47630 24104 47676 24116
rect 47882 24116 47894 24256
rect 47928 24116 47942 24292
rect 48138 24292 48198 24455
rect 48244 24376 48352 24382
rect 48244 24342 48256 24376
rect 48340 24342 48352 24376
rect 48244 24336 48352 24342
rect 48138 24136 48152 24292
rect 47882 24076 47942 24116
rect 48146 24116 48152 24136
rect 48186 24136 48198 24292
rect 48398 24292 48458 24604
rect 48656 24515 48716 24840
rect 48914 24840 48926 24870
rect 48960 25058 48972 25216
rect 49026 25316 49087 25364
rect 49026 25058 49038 25316
rect 48960 24998 49038 25058
rect 48960 24870 48966 24998
rect 48960 24840 48974 24870
rect 48760 24781 48868 24787
rect 48760 24747 48772 24781
rect 48856 24747 48868 24781
rect 48760 24741 48868 24747
rect 48780 24692 48840 24741
rect 48914 24692 48974 24840
rect 49026 24740 49038 24998
rect 49074 25300 49087 25316
rect 49074 24940 49086 25300
rect 49074 24909 49424 24940
rect 49074 24875 49177 24909
rect 49211 24875 49269 24909
rect 49303 24875 49361 24909
rect 49395 24875 49424 24909
rect 49074 24844 49424 24875
rect 49074 24740 49086 24844
rect 49026 24692 49086 24740
rect 48780 24680 49086 24692
rect 48780 24646 48802 24680
rect 49004 24646 49086 24680
rect 48780 24632 49086 24646
rect 49519 24614 49579 24620
rect 49299 24608 49519 24614
rect 49201 24592 49261 24598
rect 49195 24532 49201 24592
rect 49261 24532 49267 24592
rect 49299 24568 49311 24608
rect 49357 24568 49519 24608
rect 49299 24554 49519 24568
rect 49519 24548 49579 24554
rect 49201 24526 49261 24532
rect 48502 24376 48610 24382
rect 48502 24342 48514 24376
rect 48598 24342 48610 24376
rect 48502 24336 48610 24342
rect 48186 24116 48192 24136
rect 48146 24104 48192 24116
rect 48398 24116 48410 24292
rect 48444 24116 48458 24292
rect 48656 24292 48716 24455
rect 48786 24482 49088 24492
rect 48786 24444 48806 24482
rect 49004 24444 49088 24482
rect 48786 24432 49088 24444
rect 48786 24382 48846 24432
rect 48760 24376 48868 24382
rect 48760 24342 48772 24376
rect 48856 24342 48868 24376
rect 48760 24336 48868 24342
rect 48656 24253 48668 24292
rect 48398 24076 48458 24116
rect 48662 24116 48668 24253
rect 48702 24253 48716 24292
rect 48914 24292 48974 24432
rect 48702 24116 48708 24253
rect 48914 24246 48926 24292
rect 48920 24149 48926 24246
rect 48662 24104 48708 24116
rect 48912 24116 48926 24149
rect 48960 24246 48974 24292
rect 49028 24396 49088 24432
rect 49028 24382 49424 24396
rect 48960 24149 48966 24246
rect 48960 24116 48972 24149
rect 47470 24066 47578 24072
rect 47470 24032 47482 24066
rect 47566 24032 47578 24066
rect 47470 24026 47578 24032
rect 47728 24066 47836 24072
rect 47728 24032 47740 24066
rect 47824 24032 47836 24066
rect 47728 24026 47836 24032
rect 47986 24066 48094 24072
rect 47986 24032 47998 24066
rect 48082 24032 48094 24066
rect 47986 24026 48094 24032
rect 48244 24066 48352 24072
rect 48244 24032 48256 24066
rect 48340 24032 48352 24066
rect 48244 24026 48352 24032
rect 48502 24066 48610 24072
rect 48502 24032 48514 24066
rect 48598 24032 48610 24066
rect 48502 24026 48610 24032
rect 48760 24066 48868 24072
rect 48760 24032 48772 24066
rect 48856 24032 48868 24066
rect 48760 24026 48868 24032
rect 47494 23977 47554 24026
rect 47250 23966 47554 23977
rect 47250 23934 47332 23966
rect 47244 23874 47250 23934
rect 47310 23930 47332 23934
rect 47540 23930 47554 23966
rect 47310 23874 47554 23930
rect 47752 23967 47812 24026
rect 48012 23967 48072 24026
rect 48270 23967 48330 24026
rect 48526 23967 48586 24026
rect 48784 23977 48844 24026
rect 48912 23977 48972 24116
rect 49028 24026 49038 24382
rect 49076 24365 49424 24382
rect 49076 24331 49177 24365
rect 49211 24331 49269 24365
rect 49303 24331 49361 24365
rect 49395 24331 49424 24365
rect 49076 24300 49424 24331
rect 49076 24026 49088 24300
rect 49028 23977 49088 24026
rect 47752 23907 48526 23967
rect 48586 23907 48592 23967
rect 48784 23964 49088 23977
rect 48784 23928 48804 23964
rect 49006 23928 49088 23964
rect 47250 23860 47554 23874
rect 47251 23842 47554 23860
rect 48784 23842 49088 23928
rect 47251 23782 49089 23842
rect 47022 23478 50478 23538
rect 47251 23412 47556 23478
rect 47251 23378 47310 23412
rect 47530 23378 47556 23412
rect 47251 23364 47556 23378
rect 47251 23314 47312 23364
rect 47251 23284 47262 23314
rect 47252 23056 47262 23284
rect 47251 22996 47262 23056
rect 47252 22742 47262 22996
rect 47300 23056 47312 23314
rect 47362 23216 47422 23364
rect 47496 23315 47556 23364
rect 47752 23430 47812 23431
rect 48528 23430 48588 23436
rect 47752 23370 48528 23430
rect 47752 23315 47812 23370
rect 48010 23315 48070 23370
rect 48268 23315 48328 23370
rect 48528 23315 48588 23370
rect 48784 23412 49087 23478
rect 48784 23378 48802 23412
rect 49004 23378 49087 23412
rect 48784 23364 49087 23378
rect 48784 23315 48844 23364
rect 47470 23309 47578 23315
rect 47470 23275 47482 23309
rect 47566 23275 47578 23309
rect 47470 23269 47578 23275
rect 47728 23309 47836 23315
rect 47728 23275 47740 23309
rect 47824 23275 47836 23309
rect 47728 23269 47836 23275
rect 47986 23309 48094 23315
rect 47986 23275 47998 23309
rect 48082 23275 48094 23309
rect 47986 23269 48094 23275
rect 48244 23309 48352 23315
rect 48244 23275 48256 23309
rect 48340 23275 48352 23309
rect 48244 23269 48352 23275
rect 48502 23309 48610 23315
rect 48502 23275 48514 23309
rect 48598 23275 48610 23309
rect 48502 23269 48610 23275
rect 48760 23309 48868 23315
rect 48760 23275 48772 23309
rect 48856 23275 48868 23309
rect 48760 23269 48868 23275
rect 47362 23056 47378 23216
rect 47300 22996 47378 23056
rect 47300 22742 47312 22996
rect 47372 22874 47378 22996
rect 47252 22692 47312 22742
rect 47364 22840 47378 22874
rect 47412 22996 47422 23216
rect 47630 23216 47676 23228
rect 47412 22874 47418 22996
rect 47630 22885 47636 23216
rect 47412 22840 47424 22874
rect 47364 22692 47424 22840
rect 47622 22840 47636 22885
rect 47670 22885 47676 23216
rect 47888 23216 47934 23228
rect 47670 22840 47682 22885
rect 47888 22860 47894 23216
rect 47470 22781 47578 22787
rect 47470 22747 47482 22781
rect 47566 22747 47578 22781
rect 47470 22741 47578 22747
rect 47492 22692 47552 22741
rect 47251 22678 47552 22692
rect 47251 22644 47310 22678
rect 47530 22644 47552 22678
rect 47251 22632 47552 22644
rect 47622 22515 47682 22840
rect 47880 22840 47894 22860
rect 47928 22860 47934 23216
rect 48146 23216 48192 23228
rect 48146 22883 48152 23216
rect 47928 22840 47940 22860
rect 47728 22781 47836 22787
rect 47728 22747 47740 22781
rect 47824 22747 47836 22781
rect 47728 22741 47836 22747
rect 47880 22664 47940 22840
rect 48138 22840 48152 22883
rect 48186 22883 48192 23216
rect 48404 23216 48450 23228
rect 48186 22840 48198 22883
rect 48404 22878 48410 23216
rect 47986 22781 48094 22787
rect 47986 22747 47998 22781
rect 48082 22747 48094 22781
rect 47986 22741 48094 22747
rect 47874 22604 47880 22664
rect 47940 22604 47946 22664
rect 47250 22480 47554 22490
rect 47250 22442 47334 22480
rect 47542 22442 47554 22480
rect 47616 22455 47622 22515
rect 47682 22455 47688 22515
rect 47250 22430 47554 22442
rect 47250 22382 47310 22430
rect 47250 22026 47262 22382
rect 47298 22026 47310 22382
rect 47364 22292 47424 22430
rect 47494 22382 47554 22430
rect 47470 22376 47578 22382
rect 47470 22342 47482 22376
rect 47566 22342 47578 22376
rect 47470 22336 47578 22342
rect 47364 22242 47378 22292
rect 47372 22155 47378 22242
rect 47250 21977 47310 22026
rect 47366 22116 47378 22155
rect 47412 22242 47424 22292
rect 47622 22292 47682 22455
rect 47728 22376 47836 22382
rect 47728 22342 47740 22376
rect 47824 22342 47836 22376
rect 47728 22336 47836 22342
rect 47622 22255 47636 22292
rect 47412 22155 47418 22242
rect 47412 22116 47426 22155
rect 47366 21977 47426 22116
rect 47630 22116 47636 22255
rect 47670 22255 47682 22292
rect 47880 22322 47940 22604
rect 48138 22515 48198 22840
rect 48398 22840 48410 22878
rect 48444 22878 48450 23216
rect 48662 23216 48708 23228
rect 48662 22883 48668 23216
rect 48444 22840 48458 22878
rect 48244 22781 48352 22787
rect 48244 22747 48256 22781
rect 48340 22747 48352 22781
rect 48244 22741 48352 22747
rect 48398 22664 48458 22840
rect 48656 22840 48668 22883
rect 48702 22883 48708 23216
rect 48912 23216 48972 23364
rect 48912 22998 48926 23216
rect 48702 22840 48716 22883
rect 48920 22870 48926 22998
rect 48502 22781 48610 22787
rect 48502 22747 48514 22781
rect 48598 22747 48610 22781
rect 48502 22741 48610 22747
rect 48392 22604 48398 22664
rect 48458 22604 48464 22664
rect 48132 22455 48138 22515
rect 48198 22455 48204 22515
rect 47986 22376 48094 22382
rect 47986 22342 47998 22376
rect 48082 22342 48094 22376
rect 47986 22336 48094 22342
rect 47880 22292 47942 22322
rect 47880 22256 47894 22292
rect 47670 22116 47676 22255
rect 47630 22104 47676 22116
rect 47882 22116 47894 22256
rect 47928 22116 47942 22292
rect 48138 22292 48198 22455
rect 48244 22376 48352 22382
rect 48244 22342 48256 22376
rect 48340 22342 48352 22376
rect 48244 22336 48352 22342
rect 48138 22136 48152 22292
rect 47882 22076 47942 22116
rect 48146 22116 48152 22136
rect 48186 22136 48198 22292
rect 48398 22292 48458 22604
rect 48656 22515 48716 22840
rect 48914 22840 48926 22870
rect 48960 23058 48972 23216
rect 49026 23316 49087 23364
rect 49026 23058 49038 23316
rect 48960 22998 49038 23058
rect 48960 22870 48966 22998
rect 48960 22840 48974 22870
rect 48760 22781 48868 22787
rect 48760 22747 48772 22781
rect 48856 22747 48868 22781
rect 48760 22741 48868 22747
rect 48780 22692 48840 22741
rect 48914 22692 48974 22840
rect 49026 22740 49038 22998
rect 49074 23300 49087 23316
rect 49074 22940 49086 23300
rect 49074 22909 49424 22940
rect 49074 22875 49177 22909
rect 49211 22875 49269 22909
rect 49303 22875 49361 22909
rect 49395 22875 49424 22909
rect 49074 22844 49424 22875
rect 49074 22740 49086 22844
rect 49026 22692 49086 22740
rect 48780 22680 49086 22692
rect 48780 22646 48802 22680
rect 49004 22646 49086 22680
rect 48780 22632 49086 22646
rect 49519 22614 49579 22620
rect 49299 22608 49519 22614
rect 49201 22592 49261 22598
rect 49195 22532 49201 22592
rect 49261 22532 49267 22592
rect 49299 22568 49311 22608
rect 49357 22568 49519 22608
rect 49299 22554 49519 22568
rect 49519 22548 49579 22554
rect 49201 22526 49261 22532
rect 48502 22376 48610 22382
rect 48502 22342 48514 22376
rect 48598 22342 48610 22376
rect 48502 22336 48610 22342
rect 48186 22116 48192 22136
rect 48146 22104 48192 22116
rect 48398 22116 48410 22292
rect 48444 22116 48458 22292
rect 48656 22292 48716 22455
rect 48786 22482 49088 22492
rect 48786 22444 48806 22482
rect 49004 22444 49088 22482
rect 48786 22432 49088 22444
rect 48786 22382 48846 22432
rect 48760 22376 48868 22382
rect 48760 22342 48772 22376
rect 48856 22342 48868 22376
rect 48760 22336 48868 22342
rect 48656 22253 48668 22292
rect 48398 22076 48458 22116
rect 48662 22116 48668 22253
rect 48702 22253 48716 22292
rect 48914 22292 48974 22432
rect 48702 22116 48708 22253
rect 48914 22246 48926 22292
rect 48920 22149 48926 22246
rect 48662 22104 48708 22116
rect 48912 22116 48926 22149
rect 48960 22246 48974 22292
rect 49028 22396 49088 22432
rect 49028 22382 49424 22396
rect 48960 22149 48966 22246
rect 48960 22116 48972 22149
rect 47470 22066 47578 22072
rect 47470 22032 47482 22066
rect 47566 22032 47578 22066
rect 47470 22026 47578 22032
rect 47728 22066 47836 22072
rect 47728 22032 47740 22066
rect 47824 22032 47836 22066
rect 47728 22026 47836 22032
rect 47986 22066 48094 22072
rect 47986 22032 47998 22066
rect 48082 22032 48094 22066
rect 47986 22026 48094 22032
rect 48244 22066 48352 22072
rect 48244 22032 48256 22066
rect 48340 22032 48352 22066
rect 48244 22026 48352 22032
rect 48502 22066 48610 22072
rect 48502 22032 48514 22066
rect 48598 22032 48610 22066
rect 48502 22026 48610 22032
rect 48760 22066 48868 22072
rect 48760 22032 48772 22066
rect 48856 22032 48868 22066
rect 48760 22026 48868 22032
rect 47494 21977 47554 22026
rect 47250 21966 47554 21977
rect 47250 21930 47332 21966
rect 47540 21930 47554 21966
rect 47250 21920 47554 21930
rect 46972 21860 46978 21920
rect 47038 21860 47554 21920
rect 47752 21967 47812 22026
rect 48012 21967 48072 22026
rect 48270 21967 48330 22026
rect 48526 21967 48586 22026
rect 48784 21977 48844 22026
rect 48912 21977 48972 22116
rect 49028 22026 49038 22382
rect 49076 22365 49424 22382
rect 49076 22331 49177 22365
rect 49211 22331 49269 22365
rect 49303 22331 49361 22365
rect 49395 22331 49424 22365
rect 49076 22300 49424 22331
rect 49076 22026 49088 22300
rect 49028 21977 49088 22026
rect 47752 21907 48526 21967
rect 48586 21907 48592 21967
rect 48784 21964 49088 21977
rect 48784 21928 48804 21964
rect 49006 21928 49088 21964
rect 47251 21842 47554 21860
rect 48784 21842 49088 21928
rect 47251 21782 49089 21842
rect 34082 18088 34088 18148
rect 34148 18088 34154 18148
rect 21964 17934 30182 17994
rect 12194 17864 19994 17924
rect 12134 17858 12194 17864
rect 35666 17764 35778 18278
rect 11322 17758 35778 17764
rect 11322 17658 11428 17758
rect 35672 17658 35778 17758
rect 11322 17652 35778 17658
rect -13107 16348 -8742 16408
rect -8682 16348 -8671 16408
rect -1420 16348 -1414 16408
rect -1354 16348 -1348 16408
rect -13107 16282 -12802 16348
rect -13107 16248 -13048 16282
rect -12828 16248 -12802 16282
rect -13107 16234 -12802 16248
rect -13107 16184 -13046 16234
rect -13107 16154 -13096 16184
rect -13106 15926 -13096 16154
rect -13107 15866 -13096 15926
rect -13106 15612 -13096 15866
rect -13058 15926 -13046 16184
rect -12996 16086 -12936 16234
rect -12862 16185 -12802 16234
rect -12606 16300 -12546 16301
rect -11830 16300 -11770 16306
rect -12606 16240 -11830 16300
rect -12606 16185 -12546 16240
rect -12348 16185 -12288 16240
rect -12090 16185 -12030 16240
rect -11830 16185 -11770 16240
rect -11574 16282 -11271 16348
rect -11574 16248 -11556 16282
rect -11354 16248 -11271 16282
rect -11574 16234 -11271 16248
rect -11574 16185 -11514 16234
rect -12888 16179 -12780 16185
rect -12888 16145 -12876 16179
rect -12792 16145 -12780 16179
rect -12888 16139 -12780 16145
rect -12630 16179 -12522 16185
rect -12630 16145 -12618 16179
rect -12534 16145 -12522 16179
rect -12630 16139 -12522 16145
rect -12372 16179 -12264 16185
rect -12372 16145 -12360 16179
rect -12276 16145 -12264 16179
rect -12372 16139 -12264 16145
rect -12114 16179 -12006 16185
rect -12114 16145 -12102 16179
rect -12018 16145 -12006 16179
rect -12114 16139 -12006 16145
rect -11856 16179 -11748 16185
rect -11856 16145 -11844 16179
rect -11760 16145 -11748 16179
rect -11856 16139 -11748 16145
rect -11598 16179 -11490 16185
rect -11598 16145 -11586 16179
rect -11502 16145 -11490 16179
rect -11598 16139 -11490 16145
rect -12996 15926 -12980 16086
rect -13058 15866 -12980 15926
rect -13058 15612 -13046 15866
rect -12986 15744 -12980 15866
rect -13106 15562 -13046 15612
rect -12994 15710 -12980 15744
rect -12946 15866 -12936 16086
rect -12728 16086 -12682 16098
rect -12946 15744 -12940 15866
rect -12728 15755 -12722 16086
rect -12946 15710 -12934 15744
rect -12994 15562 -12934 15710
rect -12736 15710 -12722 15755
rect -12688 15755 -12682 16086
rect -12470 16086 -12424 16098
rect -12688 15710 -12676 15755
rect -12470 15730 -12464 16086
rect -12888 15651 -12780 15657
rect -12888 15617 -12876 15651
rect -12792 15617 -12780 15651
rect -12888 15611 -12780 15617
rect -12866 15562 -12806 15611
rect -13107 15548 -12806 15562
rect -13107 15514 -13048 15548
rect -12828 15514 -12806 15548
rect -13107 15502 -12806 15514
rect -12736 15385 -12676 15710
rect -12478 15710 -12464 15730
rect -12430 15730 -12424 16086
rect -12212 16086 -12166 16098
rect -12212 15753 -12206 16086
rect -12430 15710 -12418 15730
rect -12630 15651 -12522 15657
rect -12630 15617 -12618 15651
rect -12534 15617 -12522 15651
rect -12630 15611 -12522 15617
rect -12478 15534 -12418 15710
rect -12220 15710 -12206 15753
rect -12172 15753 -12166 16086
rect -11954 16086 -11908 16098
rect -12172 15710 -12160 15753
rect -11954 15748 -11948 16086
rect -12372 15651 -12264 15657
rect -12372 15617 -12360 15651
rect -12276 15617 -12264 15651
rect -12372 15611 -12264 15617
rect -12484 15474 -12478 15534
rect -12418 15474 -12412 15534
rect -13108 15350 -12804 15360
rect -13108 15312 -13024 15350
rect -12816 15312 -12804 15350
rect -12742 15325 -12736 15385
rect -12676 15325 -12670 15385
rect -13108 15300 -12804 15312
rect -13108 15252 -13048 15300
rect -13108 14896 -13096 15252
rect -13060 14896 -13048 15252
rect -12994 15162 -12934 15300
rect -12864 15252 -12804 15300
rect -12888 15246 -12780 15252
rect -12888 15212 -12876 15246
rect -12792 15212 -12780 15246
rect -12888 15206 -12780 15212
rect -12994 15112 -12980 15162
rect -12986 15025 -12980 15112
rect -13108 14847 -13048 14896
rect -12992 14986 -12980 15025
rect -12946 15112 -12934 15162
rect -12736 15162 -12676 15325
rect -12630 15246 -12522 15252
rect -12630 15212 -12618 15246
rect -12534 15212 -12522 15246
rect -12630 15206 -12522 15212
rect -12736 15125 -12722 15162
rect -12946 15025 -12940 15112
rect -12946 14986 -12932 15025
rect -12992 14847 -12932 14986
rect -12728 14986 -12722 15125
rect -12688 15125 -12676 15162
rect -12478 15192 -12418 15474
rect -12220 15385 -12160 15710
rect -11960 15710 -11948 15748
rect -11914 15748 -11908 16086
rect -11696 16086 -11650 16098
rect -11696 15753 -11690 16086
rect -11914 15710 -11900 15748
rect -12114 15651 -12006 15657
rect -12114 15617 -12102 15651
rect -12018 15617 -12006 15651
rect -12114 15611 -12006 15617
rect -11960 15534 -11900 15710
rect -11702 15710 -11690 15753
rect -11656 15753 -11650 16086
rect -11446 16086 -11386 16234
rect -11446 15868 -11432 16086
rect -11656 15710 -11642 15753
rect -11438 15740 -11432 15868
rect -11856 15651 -11748 15657
rect -11856 15617 -11844 15651
rect -11760 15617 -11748 15651
rect -11856 15611 -11748 15617
rect -11966 15474 -11960 15534
rect -11900 15474 -11894 15534
rect -12226 15325 -12220 15385
rect -12160 15325 -12154 15385
rect -12372 15246 -12264 15252
rect -12372 15212 -12360 15246
rect -12276 15212 -12264 15246
rect -12372 15206 -12264 15212
rect -12478 15162 -12416 15192
rect -12478 15126 -12464 15162
rect -12688 14986 -12682 15125
rect -12476 15054 -12464 15126
rect -12728 14974 -12682 14986
rect -12478 14986 -12464 15054
rect -12430 14986 -12416 15162
rect -12220 15162 -12160 15325
rect -12114 15246 -12006 15252
rect -12114 15212 -12102 15246
rect -12018 15212 -12006 15246
rect -12114 15206 -12006 15212
rect -12220 15006 -12206 15162
rect -12478 14956 -12416 14986
rect -12212 14986 -12206 15006
rect -12172 15006 -12160 15162
rect -11960 15162 -11900 15474
rect -11702 15385 -11642 15710
rect -11444 15710 -11432 15740
rect -11398 15928 -11386 16086
rect -11332 16186 -11271 16234
rect -11332 15928 -11320 16186
rect -11398 15868 -11320 15928
rect -11398 15740 -11392 15868
rect -11398 15710 -11384 15740
rect -11598 15651 -11490 15657
rect -11598 15617 -11586 15651
rect -11502 15617 -11490 15651
rect -11598 15611 -11490 15617
rect -11578 15562 -11518 15611
rect -11444 15562 -11384 15710
rect -11332 15610 -11320 15868
rect -11284 16170 -11271 16186
rect -10507 16282 -10202 16348
rect -10507 16248 -10448 16282
rect -10228 16248 -10202 16282
rect -10507 16234 -10202 16248
rect -10507 16184 -10446 16234
rect -11284 15810 -11272 16170
rect -10507 16154 -10496 16184
rect -10506 15926 -10496 16154
rect -10507 15866 -10496 15926
rect -11284 15779 -10934 15810
rect -11284 15745 -11181 15779
rect -11147 15745 -11089 15779
rect -11055 15745 -10997 15779
rect -10963 15745 -10934 15779
rect -11284 15714 -10934 15745
rect -11284 15610 -11272 15714
rect -11332 15562 -11272 15610
rect -10506 15612 -10496 15866
rect -10458 15926 -10446 16184
rect -10396 16086 -10336 16234
rect -10262 16185 -10202 16234
rect -10006 16300 -9946 16301
rect -9230 16300 -9170 16306
rect -10006 16240 -9230 16300
rect -10006 16185 -9946 16240
rect -9748 16185 -9688 16240
rect -9490 16185 -9430 16240
rect -9230 16185 -9170 16240
rect -8974 16282 -8671 16348
rect -8974 16248 -8956 16282
rect -8754 16248 -8671 16282
rect -8974 16234 -8671 16248
rect -8974 16185 -8914 16234
rect -10288 16179 -10180 16185
rect -10288 16145 -10276 16179
rect -10192 16145 -10180 16179
rect -10288 16139 -10180 16145
rect -10030 16179 -9922 16185
rect -10030 16145 -10018 16179
rect -9934 16145 -9922 16179
rect -10030 16139 -9922 16145
rect -9772 16179 -9664 16185
rect -9772 16145 -9760 16179
rect -9676 16145 -9664 16179
rect -9772 16139 -9664 16145
rect -9514 16179 -9406 16185
rect -9514 16145 -9502 16179
rect -9418 16145 -9406 16179
rect -9514 16139 -9406 16145
rect -9256 16179 -9148 16185
rect -9256 16145 -9244 16179
rect -9160 16145 -9148 16179
rect -9256 16139 -9148 16145
rect -8998 16179 -8890 16185
rect -8998 16145 -8986 16179
rect -8902 16145 -8890 16179
rect -8998 16139 -8890 16145
rect -10396 15926 -10380 16086
rect -10458 15866 -10380 15926
rect -10458 15612 -10446 15866
rect -10386 15744 -10380 15866
rect -10506 15562 -10446 15612
rect -10394 15710 -10380 15744
rect -10346 15866 -10336 16086
rect -10128 16086 -10082 16098
rect -10346 15744 -10340 15866
rect -10128 15755 -10122 16086
rect -10346 15710 -10334 15744
rect -10394 15562 -10334 15710
rect -10136 15710 -10122 15755
rect -10088 15755 -10082 16086
rect -9870 16086 -9824 16098
rect -10088 15710 -10076 15755
rect -9870 15730 -9864 16086
rect -10288 15651 -10180 15657
rect -10288 15617 -10276 15651
rect -10192 15617 -10180 15651
rect -10288 15611 -10180 15617
rect -10266 15562 -10206 15611
rect -11578 15550 -11272 15562
rect -11578 15516 -11556 15550
rect -11354 15516 -11272 15550
rect -11578 15502 -11272 15516
rect -10507 15548 -10206 15562
rect -10507 15514 -10448 15548
rect -10228 15514 -10206 15548
rect -10507 15502 -10206 15514
rect -10839 15484 -10779 15490
rect -11059 15478 -10839 15484
rect -11157 15462 -11097 15468
rect -11163 15402 -11157 15462
rect -11097 15402 -11091 15462
rect -11059 15438 -11047 15478
rect -11001 15438 -10839 15478
rect -11059 15424 -10839 15438
rect -10839 15418 -10779 15424
rect -11157 15396 -11097 15402
rect -10136 15385 -10076 15710
rect -9878 15710 -9864 15730
rect -9830 15730 -9824 16086
rect -9612 16086 -9566 16098
rect -9612 15753 -9606 16086
rect -9830 15710 -9818 15730
rect -10030 15651 -9922 15657
rect -10030 15617 -10018 15651
rect -9934 15617 -9922 15651
rect -10030 15611 -9922 15617
rect -9878 15534 -9818 15710
rect -9620 15710 -9606 15753
rect -9572 15753 -9566 16086
rect -9354 16086 -9308 16098
rect -9572 15710 -9560 15753
rect -9354 15748 -9348 16086
rect -9772 15651 -9664 15657
rect -9772 15617 -9760 15651
rect -9676 15617 -9664 15651
rect -9772 15611 -9664 15617
rect -9884 15474 -9878 15534
rect -9818 15474 -9812 15534
rect -11856 15246 -11748 15252
rect -11856 15212 -11844 15246
rect -11760 15212 -11748 15246
rect -11856 15206 -11748 15212
rect -12172 14986 -12166 15006
rect -12212 14974 -12166 14986
rect -11960 14986 -11948 15162
rect -11914 14986 -11900 15162
rect -11702 15162 -11642 15325
rect -11572 15352 -11270 15362
rect -11572 15314 -11552 15352
rect -11354 15314 -11270 15352
rect -11572 15302 -11270 15314
rect -11572 15252 -11512 15302
rect -11598 15246 -11490 15252
rect -11598 15212 -11586 15246
rect -11502 15212 -11490 15246
rect -11598 15206 -11490 15212
rect -11702 15123 -11690 15162
rect -12888 14936 -12780 14942
rect -12888 14902 -12876 14936
rect -12792 14902 -12780 14936
rect -12888 14896 -12780 14902
rect -12630 14936 -12522 14942
rect -12630 14902 -12618 14936
rect -12534 14902 -12522 14936
rect -12630 14896 -12522 14902
rect -12484 14896 -12478 14956
rect -12418 14896 -12412 14956
rect -11960 14946 -11900 14986
rect -11696 14986 -11690 15123
rect -11656 15123 -11642 15162
rect -11444 15162 -11384 15302
rect -11656 14986 -11650 15123
rect -11444 15116 -11432 15162
rect -11438 15019 -11432 15116
rect -11696 14974 -11650 14986
rect -11446 14986 -11432 15019
rect -11398 15116 -11384 15162
rect -11330 15266 -11270 15302
rect -10508 15350 -10204 15360
rect -10508 15312 -10424 15350
rect -10216 15312 -10204 15350
rect -10142 15325 -10136 15385
rect -10076 15325 -10070 15385
rect -10508 15300 -10204 15312
rect -11330 15252 -10934 15266
rect -11398 15019 -11392 15116
rect -11398 14986 -11386 15019
rect -12372 14936 -12264 14942
rect -12372 14902 -12360 14936
rect -12276 14902 -12264 14936
rect -12372 14896 -12264 14902
rect -12114 14936 -12006 14942
rect -12114 14902 -12102 14936
rect -12018 14902 -12006 14936
rect -12114 14896 -12006 14902
rect -11856 14936 -11748 14942
rect -11856 14902 -11844 14936
rect -11760 14902 -11748 14936
rect -11856 14896 -11748 14902
rect -11598 14936 -11490 14942
rect -11598 14902 -11586 14936
rect -11502 14902 -11490 14936
rect -11598 14896 -11490 14902
rect -12864 14847 -12804 14896
rect -13108 14836 -12804 14847
rect -13108 14800 -13026 14836
rect -12818 14800 -12804 14836
rect -13108 14730 -12804 14800
rect -12606 14837 -12546 14896
rect -12346 14837 -12286 14896
rect -12088 14837 -12028 14896
rect -11832 14837 -11772 14896
rect -11574 14847 -11514 14896
rect -11446 14847 -11386 14986
rect -11330 14896 -11320 15252
rect -11282 15235 -10934 15252
rect -11282 15201 -11181 15235
rect -11147 15201 -11089 15235
rect -11055 15201 -10997 15235
rect -10963 15201 -10934 15235
rect -11282 15170 -10934 15201
rect -10508 15252 -10448 15300
rect -11282 14896 -11270 15170
rect -11330 14847 -11270 14896
rect -12606 14777 -11832 14837
rect -11772 14777 -11766 14837
rect -11574 14834 -11270 14847
rect -11574 14798 -11554 14834
rect -11352 14798 -11270 14834
rect -13107 14712 -12804 14730
rect -11574 14712 -11270 14798
rect -10508 14896 -10496 15252
rect -10460 14896 -10448 15252
rect -10394 15162 -10334 15300
rect -10264 15252 -10204 15300
rect -10288 15246 -10180 15252
rect -10288 15212 -10276 15246
rect -10192 15212 -10180 15246
rect -10288 15206 -10180 15212
rect -10394 15112 -10380 15162
rect -10386 15025 -10380 15112
rect -10508 14847 -10448 14896
rect -10392 14986 -10380 15025
rect -10346 15112 -10334 15162
rect -10136 15162 -10076 15325
rect -10030 15246 -9922 15252
rect -10030 15212 -10018 15246
rect -9934 15212 -9922 15246
rect -10030 15206 -9922 15212
rect -10136 15125 -10122 15162
rect -10346 15025 -10340 15112
rect -10346 14986 -10332 15025
rect -10392 14847 -10332 14986
rect -10128 14986 -10122 15125
rect -10088 15125 -10076 15162
rect -9878 15192 -9818 15474
rect -9620 15385 -9560 15710
rect -9360 15710 -9348 15748
rect -9314 15748 -9308 16086
rect -9096 16086 -9050 16098
rect -9096 15753 -9090 16086
rect -9314 15710 -9300 15748
rect -9514 15651 -9406 15657
rect -9514 15617 -9502 15651
rect -9418 15617 -9406 15651
rect -9514 15611 -9406 15617
rect -9360 15534 -9300 15710
rect -9102 15710 -9090 15753
rect -9056 15753 -9050 16086
rect -8846 16086 -8786 16234
rect -8846 15868 -8832 16086
rect -9056 15710 -9042 15753
rect -8838 15740 -8832 15868
rect -9256 15651 -9148 15657
rect -9256 15617 -9244 15651
rect -9160 15617 -9148 15651
rect -9256 15611 -9148 15617
rect -9366 15474 -9360 15534
rect -9300 15474 -9294 15534
rect -9626 15325 -9620 15385
rect -9560 15325 -9554 15385
rect -9772 15246 -9664 15252
rect -9772 15212 -9760 15246
rect -9676 15212 -9664 15246
rect -9772 15206 -9664 15212
rect -9878 15162 -9816 15192
rect -9878 15126 -9864 15162
rect -10088 14986 -10082 15125
rect -9876 15078 -9864 15126
rect -10128 14974 -10082 14986
rect -9878 14986 -9864 15078
rect -9830 14986 -9816 15162
rect -9620 15162 -9560 15325
rect -9514 15246 -9406 15252
rect -9514 15212 -9502 15246
rect -9418 15212 -9406 15246
rect -9514 15206 -9406 15212
rect -9620 15006 -9606 15162
rect -9878 14952 -9816 14986
rect -9612 14986 -9606 15006
rect -9572 15006 -9560 15162
rect -9360 15162 -9300 15474
rect -9102 15385 -9042 15710
rect -8844 15710 -8832 15740
rect -8798 15928 -8786 16086
rect -8732 16186 -8671 16234
rect -8732 15928 -8720 16186
rect -8798 15868 -8720 15928
rect -8798 15740 -8792 15868
rect -8798 15710 -8784 15740
rect -8998 15651 -8890 15657
rect -8998 15617 -8986 15651
rect -8902 15617 -8890 15651
rect -8998 15611 -8890 15617
rect -8978 15562 -8918 15611
rect -8844 15562 -8784 15710
rect -8732 15610 -8720 15868
rect -8684 16170 -8671 16186
rect -8684 15810 -8672 16170
rect -8684 15779 -7834 15810
rect -8684 15745 -8581 15779
rect -8547 15745 -8489 15779
rect -8455 15745 -8397 15779
rect -8363 15745 -8081 15779
rect -8047 15745 -7989 15779
rect -7955 15745 -7897 15779
rect -7863 15745 -7834 15779
rect -8684 15714 -7834 15745
rect -8684 15610 -8672 15714
rect -8732 15562 -8672 15610
rect -8978 15550 -8672 15562
rect -8978 15516 -8956 15550
rect -8754 15516 -8672 15550
rect -8978 15502 -8672 15516
rect -8239 15484 -8179 15490
rect -8459 15478 -8239 15484
rect -8557 15462 -8497 15468
rect -8563 15402 -8557 15462
rect -8497 15402 -8491 15462
rect -8459 15438 -8447 15478
rect -8401 15438 -8239 15478
rect -8459 15424 -8239 15438
rect -8179 15478 -7992 15484
rect -8179 15430 -8052 15478
rect -8004 15430 -7992 15478
rect -8179 15424 -7992 15430
rect -7962 15482 -7734 15488
rect -7962 15434 -7950 15482
rect -7902 15434 -7734 15482
rect -7962 15428 -7734 15434
rect -8239 15418 -8179 15424
rect -8557 15396 -8497 15402
rect 10305 15368 10427 15373
rect -1378 15364 35878 15368
rect -1378 15362 5912 15364
rect 6012 15362 8512 15364
rect 8612 15362 10316 15364
rect 10416 15362 35878 15364
rect -9256 15246 -9148 15252
rect -9256 15212 -9244 15246
rect -9160 15212 -9148 15246
rect -9256 15206 -9148 15212
rect -9572 14986 -9566 15006
rect -9612 14974 -9566 14986
rect -9360 14986 -9348 15162
rect -9314 14986 -9300 15162
rect -9102 15162 -9042 15325
rect -8972 15352 -8670 15362
rect -8972 15314 -8952 15352
rect -8754 15314 -8670 15352
rect -8972 15302 -8670 15314
rect -8972 15252 -8912 15302
rect -8998 15246 -8890 15252
rect -8998 15212 -8986 15246
rect -8902 15212 -8890 15246
rect -8998 15206 -8890 15212
rect -9102 15123 -9090 15162
rect -10288 14936 -10180 14942
rect -10288 14902 -10276 14936
rect -10192 14902 -10180 14936
rect -10288 14896 -10180 14902
rect -10030 14936 -9922 14942
rect -10030 14902 -10018 14936
rect -9934 14902 -9922 14936
rect -10030 14896 -9922 14902
rect -10264 14847 -10204 14896
rect -10508 14836 -10204 14847
rect -10508 14800 -10426 14836
rect -10218 14800 -10204 14836
rect -10508 14712 -10204 14800
rect -10006 14837 -9946 14896
rect -9884 14892 -9878 14952
rect -9818 14892 -9812 14952
rect -9360 14946 -9300 14986
rect -9096 14986 -9090 15123
rect -9056 15123 -9042 15162
rect -8844 15162 -8784 15302
rect -9056 14986 -9050 15123
rect -8844 15116 -8832 15162
rect -8838 15019 -8832 15116
rect -9096 14974 -9050 14986
rect -8846 14986 -8832 15019
rect -8798 15116 -8784 15162
rect -8730 15266 -8670 15302
rect -8730 15252 -7834 15266
rect -8798 15019 -8792 15116
rect -8798 14986 -8786 15019
rect -9772 14936 -9664 14942
rect -9772 14902 -9760 14936
rect -9676 14902 -9664 14936
rect -9772 14896 -9664 14902
rect -9514 14936 -9406 14942
rect -9514 14902 -9502 14936
rect -9418 14902 -9406 14936
rect -9514 14896 -9406 14902
rect -9256 14936 -9148 14942
rect -9256 14902 -9244 14936
rect -9160 14902 -9148 14936
rect -9256 14896 -9148 14902
rect -8998 14936 -8890 14942
rect -8998 14902 -8986 14936
rect -8902 14902 -8890 14936
rect -8998 14896 -8890 14902
rect -9746 14837 -9686 14896
rect -9488 14837 -9428 14896
rect -9232 14837 -9172 14896
rect -8974 14847 -8914 14896
rect -8846 14847 -8786 14986
rect -8730 14896 -8720 15252
rect -8682 15235 -7834 15252
rect -8682 15201 -8581 15235
rect -8547 15201 -8489 15235
rect -8455 15201 -8397 15235
rect -8363 15201 -8081 15235
rect -8047 15201 -7989 15235
rect -7955 15201 -7897 15235
rect -7863 15201 -7834 15235
rect -8682 15170 -7834 15201
rect -1378 15262 -1272 15362
rect 35772 15262 35878 15362
rect -1378 15256 35878 15262
rect -8682 14896 -8670 15170
rect -8730 14847 -8670 14896
rect -9946 14777 -9232 14837
rect -9172 14777 -9166 14837
rect -8974 14834 -8670 14847
rect -8974 14798 -8954 14834
rect -8752 14798 -8670 14834
rect -10006 14771 -9946 14777
rect -8974 14712 -8670 14798
rect -1792 14712 -1732 14718
rect -1378 14712 -1266 15256
rect 12898 15132 12904 15192
rect 12964 15132 12970 15192
rect 13054 15132 13060 15192
rect 13120 15132 13126 15192
rect 13286 15184 13346 15190
rect -13107 14652 -8750 14712
rect -8690 14652 -8669 14712
rect -1732 14652 -1266 14712
rect -8750 14646 -8690 14652
rect -1792 14646 -1732 14652
rect -1378 14470 -1266 14652
rect -1378 210 -1372 14470
rect -1272 210 -1266 14470
rect 12904 14354 12964 15132
rect 8878 14294 12964 14354
rect 8878 14216 8938 14294
rect 1754 14156 8938 14216
rect 1754 14016 1814 14156
rect 2264 14106 2324 14156
rect 2048 14100 2536 14106
rect 2048 14066 2060 14100
rect 2524 14066 2536 14100
rect 2048 14060 2536 14066
rect 1754 13986 1766 14016
rect 1760 13458 1766 13986
rect 1750 13440 1766 13458
rect 1800 13986 1814 14016
rect 2770 14016 2830 14156
rect 3272 14106 3332 14156
rect 4300 14106 4360 14156
rect 3066 14100 3554 14106
rect 3066 14066 3078 14100
rect 3542 14066 3554 14100
rect 3066 14060 3554 14066
rect 4084 14100 4572 14106
rect 4084 14066 4096 14100
rect 4560 14066 4572 14100
rect 4084 14060 4572 14066
rect 2770 13992 2784 14016
rect 1800 13458 1806 13986
rect 2778 13462 2784 13992
rect 1800 13440 1810 13458
rect 1750 13198 1810 13440
rect 2770 13440 2784 13462
rect 2818 13992 2830 14016
rect 3796 14016 3842 14028
rect 2818 13462 2824 13992
rect 3796 13464 3802 14016
rect 2818 13440 2830 13462
rect 2048 13390 2536 13396
rect 2048 13356 2060 13390
rect 2524 13356 2536 13390
rect 2048 13350 2536 13356
rect 2264 13288 2324 13350
rect 2048 13282 2536 13288
rect 2048 13248 2060 13282
rect 2524 13248 2536 13282
rect 2048 13242 2536 13248
rect 1750 13168 1766 13198
rect 1760 12644 1766 13168
rect 1752 12622 1766 12644
rect 1800 13168 1810 13198
rect 2770 13198 2830 13440
rect 3790 13440 3802 13464
rect 3836 13464 3842 14016
rect 4808 14016 4868 14156
rect 5314 14106 5374 14156
rect 6328 14106 6388 14156
rect 5102 14100 5590 14106
rect 5102 14066 5114 14100
rect 5578 14066 5590 14100
rect 5102 14060 5590 14066
rect 6120 14100 6608 14106
rect 6120 14066 6132 14100
rect 6596 14066 6608 14100
rect 6120 14060 6608 14066
rect 4808 13978 4820 14016
rect 3836 13440 3850 13464
rect 4814 13460 4820 13978
rect 3066 13390 3554 13396
rect 3066 13356 3078 13390
rect 3542 13356 3554 13390
rect 3066 13350 3554 13356
rect 3268 13288 3328 13350
rect 3066 13282 3554 13288
rect 3066 13248 3078 13282
rect 3542 13248 3554 13282
rect 3066 13242 3554 13248
rect 2770 13172 2784 13198
rect 1800 12644 1806 13168
rect 2778 12648 2784 13172
rect 1800 12622 1812 12644
rect 1752 12380 1812 12622
rect 2772 12622 2784 12648
rect 2818 13172 2830 13198
rect 3790 13198 3850 13440
rect 4808 13440 4820 13460
rect 4854 13978 4868 14016
rect 5832 14016 5878 14028
rect 6844 14016 6904 14156
rect 7360 14106 7420 14156
rect 8366 14106 8426 14156
rect 7138 14100 7626 14106
rect 7138 14066 7150 14100
rect 7614 14066 7626 14100
rect 7138 14060 7626 14066
rect 8156 14100 8644 14106
rect 8156 14066 8168 14100
rect 8632 14066 8644 14100
rect 8156 14060 8644 14066
rect 4854 13460 4860 13978
rect 5832 13468 5838 14016
rect 4854 13440 4868 13460
rect 4084 13390 4572 13396
rect 4084 13356 4096 13390
rect 4560 13356 4572 13390
rect 4084 13350 4572 13356
rect 4298 13288 4358 13350
rect 4084 13282 4572 13288
rect 4084 13248 4096 13282
rect 4560 13248 4572 13282
rect 4084 13242 4572 13248
rect 3790 13174 3802 13198
rect 2818 12648 2824 13172
rect 3796 12650 3802 13174
rect 2818 12622 2832 12648
rect 2048 12572 2536 12578
rect 2048 12538 2060 12572
rect 2524 12538 2536 12572
rect 2048 12532 2536 12538
rect 2264 12470 2324 12532
rect 2048 12464 2536 12470
rect 2048 12430 2060 12464
rect 2524 12430 2536 12464
rect 2048 12424 2536 12430
rect 1752 12354 1766 12380
rect 1760 11816 1766 12354
rect 1752 11804 1766 11816
rect 1800 12354 1812 12380
rect 2772 12380 2832 12622
rect 3792 12622 3802 12650
rect 3836 13174 3850 13198
rect 4808 13198 4868 13440
rect 5828 13440 5838 13468
rect 5872 13468 5878 14016
rect 6842 13982 6856 14016
rect 6844 13970 6856 13982
rect 5872 13440 5888 13468
rect 6850 13460 6856 13970
rect 5102 13390 5590 13396
rect 5102 13356 5114 13390
rect 5578 13356 5590 13390
rect 5102 13350 5590 13356
rect 5300 13288 5360 13350
rect 5102 13282 5590 13288
rect 5102 13248 5114 13282
rect 5578 13248 5590 13282
rect 5102 13242 5590 13248
rect 3836 12650 3842 13174
rect 4808 13170 4820 13198
rect 3836 12622 3852 12650
rect 4814 12646 4820 13170
rect 3066 12572 3554 12578
rect 3066 12538 3078 12572
rect 3542 12538 3554 12572
rect 3066 12532 3554 12538
rect 3280 12470 3340 12532
rect 3066 12464 3554 12470
rect 3066 12430 3078 12464
rect 3542 12430 3554 12464
rect 3066 12424 3554 12430
rect 2772 12358 2784 12380
rect 1800 11816 1806 12354
rect 2778 11820 2784 12358
rect 1800 11804 1812 11816
rect 1752 11562 1812 11804
rect 2772 11804 2784 11820
rect 2818 12358 2832 12380
rect 3792 12380 3852 12622
rect 4810 12622 4820 12646
rect 4854 13170 4868 13198
rect 5828 13198 5888 13440
rect 6840 13440 6856 13460
rect 6890 13970 6904 14016
rect 7868 14016 7914 14028
rect 6890 13460 6896 13970
rect 7868 13460 7874 14016
rect 6890 13440 6900 13460
rect 6120 13390 6608 13396
rect 6120 13356 6132 13390
rect 6596 13356 6608 13390
rect 6120 13350 6608 13356
rect 6330 13288 6390 13350
rect 6120 13282 6608 13288
rect 6120 13248 6132 13282
rect 6596 13248 6608 13282
rect 6120 13242 6608 13248
rect 5828 13178 5838 13198
rect 4854 12646 4860 13170
rect 5832 12654 5838 13178
rect 4854 12622 4870 12646
rect 4084 12572 4572 12578
rect 4084 12538 4096 12572
rect 4560 12538 4572 12572
rect 4084 12532 4572 12538
rect 4298 12470 4358 12532
rect 4084 12464 4572 12470
rect 4084 12430 4096 12464
rect 4560 12430 4572 12464
rect 4084 12424 4572 12430
rect 3792 12360 3802 12380
rect 2818 11820 2824 12358
rect 3796 11822 3802 12360
rect 2818 11804 2832 11820
rect 2048 11754 2536 11760
rect 2048 11720 2060 11754
rect 2524 11720 2536 11754
rect 2048 11714 2536 11720
rect 2258 11652 2318 11714
rect 2048 11646 2536 11652
rect 2048 11612 2060 11646
rect 2524 11612 2536 11646
rect 2048 11606 2536 11612
rect 1752 11526 1766 11562
rect 1760 11004 1766 11526
rect 1752 10986 1766 11004
rect 1800 11526 1812 11562
rect 2772 11562 2832 11804
rect 3792 11804 3802 11822
rect 3836 12360 3852 12380
rect 4810 12380 4870 12622
rect 5830 12622 5838 12654
rect 5872 13178 5888 13198
rect 6840 13198 6900 13440
rect 7862 13440 7874 13460
rect 7908 13460 7914 14016
rect 8878 14016 8938 14156
rect 9388 14106 9448 14294
rect 12134 14206 12194 14212
rect 10918 14146 12134 14206
rect 9174 14100 9662 14106
rect 9174 14066 9186 14100
rect 9650 14066 9662 14100
rect 9174 14060 9662 14066
rect 10192 14100 10680 14106
rect 10192 14066 10204 14100
rect 10668 14066 10680 14100
rect 10192 14060 10680 14066
rect 8878 13980 8892 14016
rect 8886 13460 8892 13980
rect 7908 13440 7922 13460
rect 7138 13390 7626 13396
rect 7138 13356 7150 13390
rect 7614 13356 7626 13390
rect 7138 13350 7626 13356
rect 7346 13288 7406 13350
rect 7138 13282 7626 13288
rect 7138 13248 7150 13282
rect 7614 13248 7626 13282
rect 7138 13242 7626 13248
rect 5872 12654 5878 13178
rect 6840 13170 6856 13198
rect 5872 12622 5890 12654
rect 6850 12646 6856 13170
rect 5102 12572 5590 12578
rect 5102 12538 5114 12572
rect 5578 12538 5590 12572
rect 5102 12532 5590 12538
rect 5300 12470 5360 12532
rect 5102 12464 5590 12470
rect 5102 12430 5114 12464
rect 5578 12430 5590 12464
rect 5102 12424 5590 12430
rect 3836 11822 3842 12360
rect 4810 12356 4820 12380
rect 3836 11804 3852 11822
rect 4814 11818 4820 12356
rect 3066 11754 3554 11760
rect 3066 11720 3078 11754
rect 3542 11720 3554 11754
rect 3066 11714 3554 11720
rect 3280 11652 3340 11714
rect 3066 11646 3554 11652
rect 3066 11612 3078 11646
rect 3542 11612 3554 11646
rect 3066 11606 3554 11612
rect 2772 11530 2784 11562
rect 1800 11004 1806 11526
rect 2778 11008 2784 11530
rect 1800 10986 1812 11004
rect 1752 10744 1812 10986
rect 2772 10986 2784 11008
rect 2818 11530 2832 11562
rect 3792 11562 3852 11804
rect 4810 11804 4820 11818
rect 4854 12356 4870 12380
rect 5830 12380 5890 12622
rect 6842 12622 6856 12646
rect 6890 13170 6900 13198
rect 7862 13198 7922 13440
rect 8882 13440 8892 13460
rect 8926 13980 8938 14016
rect 9904 14016 9950 14028
rect 8926 13460 8932 13980
rect 9904 13464 9910 14016
rect 8926 13440 8942 13460
rect 8156 13390 8644 13396
rect 8156 13356 8168 13390
rect 8632 13356 8644 13390
rect 8156 13350 8644 13356
rect 8368 13288 8428 13350
rect 8156 13282 8644 13288
rect 8156 13248 8168 13282
rect 8632 13248 8644 13282
rect 8156 13242 8644 13248
rect 7862 13170 7874 13198
rect 6890 12646 6896 13170
rect 7868 12646 7874 13170
rect 6890 12622 6902 12646
rect 6120 12572 6608 12578
rect 6120 12538 6132 12572
rect 6596 12538 6608 12572
rect 6120 12532 6608 12538
rect 6330 12470 6390 12532
rect 6120 12464 6608 12470
rect 6120 12430 6132 12464
rect 6596 12430 6608 12464
rect 6120 12424 6608 12430
rect 5830 12364 5838 12380
rect 4854 11818 4860 12356
rect 5832 11826 5838 12364
rect 4854 11804 4870 11818
rect 4084 11754 4572 11760
rect 4084 11720 4096 11754
rect 4560 11720 4572 11754
rect 4084 11714 4572 11720
rect 4292 11652 4352 11714
rect 4084 11646 4572 11652
rect 4084 11612 4096 11646
rect 4560 11612 4572 11646
rect 4084 11606 4572 11612
rect 3792 11532 3802 11562
rect 2818 11008 2824 11530
rect 3796 11010 3802 11532
rect 2818 10986 2832 11008
rect 2048 10936 2536 10942
rect 2048 10902 2060 10936
rect 2524 10902 2536 10936
rect 2048 10896 2536 10902
rect 2256 10834 2316 10896
rect 2048 10828 2536 10834
rect 2048 10794 2060 10828
rect 2524 10794 2536 10828
rect 2048 10788 2536 10794
rect 1752 10714 1766 10744
rect 1760 10184 1766 10714
rect 1752 10168 1766 10184
rect 1800 10714 1812 10744
rect 2772 10744 2832 10986
rect 3792 10986 3802 11010
rect 3836 11532 3852 11562
rect 4810 11562 4870 11804
rect 5830 11804 5838 11826
rect 5872 12364 5890 12380
rect 6842 12380 6902 12622
rect 7864 12622 7874 12646
rect 7908 13170 7922 13198
rect 8882 13198 8942 13440
rect 9898 13440 9910 13464
rect 9944 13464 9950 14016
rect 10918 14016 10978 14146
rect 12134 14140 12194 14146
rect 12794 14032 12800 14092
rect 12860 14032 12866 14092
rect 10918 13964 10928 14016
rect 9944 13440 9958 13464
rect 10922 13460 10928 13964
rect 9174 13390 9662 13396
rect 9174 13356 9186 13390
rect 9650 13356 9662 13390
rect 9174 13350 9662 13356
rect 9380 13288 9440 13350
rect 9174 13282 9662 13288
rect 9174 13248 9186 13282
rect 9650 13248 9662 13282
rect 9174 13242 9662 13248
rect 8882 13170 8892 13198
rect 7908 12646 7914 13170
rect 8886 12646 8892 13170
rect 7908 12622 7924 12646
rect 7138 12572 7626 12578
rect 7138 12538 7150 12572
rect 7614 12538 7626 12572
rect 7138 12532 7626 12538
rect 7346 12470 7406 12532
rect 7138 12464 7626 12470
rect 7138 12430 7150 12464
rect 7614 12430 7626 12464
rect 7138 12424 7626 12430
rect 5872 11826 5878 12364
rect 6842 12356 6856 12380
rect 5872 11804 5890 11826
rect 6850 11818 6856 12356
rect 5102 11754 5590 11760
rect 5102 11720 5114 11754
rect 5578 11720 5590 11754
rect 5102 11714 5590 11720
rect 5294 11652 5354 11714
rect 5102 11646 5590 11652
rect 5102 11612 5114 11646
rect 5578 11612 5590 11646
rect 5102 11606 5590 11612
rect 3836 11010 3842 11532
rect 4810 11528 4820 11562
rect 3836 10986 3852 11010
rect 4814 11006 4820 11528
rect 3066 10936 3554 10942
rect 3066 10902 3078 10936
rect 3542 10902 3554 10936
rect 3066 10896 3554 10902
rect 3274 10834 3334 10896
rect 3066 10828 3554 10834
rect 3066 10794 3078 10828
rect 3542 10794 3554 10828
rect 3066 10788 3554 10794
rect 2772 10718 2784 10744
rect 1800 10184 1806 10714
rect 2778 10188 2784 10718
rect 1800 10168 1812 10184
rect 1752 9926 1812 10168
rect 2772 10168 2784 10188
rect 2818 10718 2832 10744
rect 3792 10744 3852 10986
rect 4810 10986 4820 11006
rect 4854 11528 4870 11562
rect 5830 11562 5890 11804
rect 6842 11804 6856 11818
rect 6890 12356 6902 12380
rect 7864 12380 7924 12622
rect 8884 12622 8892 12646
rect 8926 13170 8942 13198
rect 9898 13198 9958 13440
rect 10920 13440 10928 13460
rect 10962 13964 10978 14016
rect 10962 13460 10968 13964
rect 10962 13440 10980 13460
rect 10192 13390 10680 13396
rect 10192 13356 10204 13390
rect 10668 13356 10680 13390
rect 10192 13350 10680 13356
rect 10400 13288 10460 13350
rect 10192 13282 10680 13288
rect 10192 13248 10204 13282
rect 10668 13248 10680 13282
rect 10192 13242 10680 13248
rect 9898 13174 9910 13198
rect 8926 12646 8932 13170
rect 9904 12650 9910 13174
rect 8926 12622 8944 12646
rect 8156 12572 8644 12578
rect 8156 12538 8168 12572
rect 8632 12538 8644 12572
rect 8156 12532 8644 12538
rect 8368 12470 8428 12532
rect 8156 12464 8644 12470
rect 8156 12430 8168 12464
rect 8632 12430 8644 12464
rect 8156 12424 8644 12430
rect 7864 12356 7874 12380
rect 6890 11818 6896 12356
rect 7868 11818 7874 12356
rect 6890 11804 6902 11818
rect 6120 11754 6608 11760
rect 6120 11720 6132 11754
rect 6596 11720 6608 11754
rect 6120 11714 6608 11720
rect 6324 11652 6384 11714
rect 6120 11646 6608 11652
rect 6120 11612 6132 11646
rect 6596 11612 6608 11646
rect 6120 11606 6608 11612
rect 5830 11536 5838 11562
rect 4854 11006 4860 11528
rect 5832 11014 5838 11536
rect 4854 10986 4870 11006
rect 4084 10936 4572 10942
rect 4084 10902 4096 10936
rect 4560 10902 4572 10936
rect 4084 10896 4572 10902
rect 4290 10834 4350 10896
rect 4084 10828 4572 10834
rect 4084 10794 4096 10828
rect 4560 10794 4572 10828
rect 4084 10788 4572 10794
rect 3792 10720 3802 10744
rect 2818 10188 2824 10718
rect 3796 10190 3802 10720
rect 2818 10168 2832 10188
rect 2048 10118 2536 10124
rect 2048 10084 2060 10118
rect 2524 10084 2536 10118
rect 2048 10078 2536 10084
rect 2258 10016 2318 10078
rect 2048 10010 2536 10016
rect 2048 9976 2060 10010
rect 2524 9976 2536 10010
rect 2048 9970 2536 9976
rect 1752 9894 1766 9926
rect 1760 9372 1766 9894
rect 1752 9350 1766 9372
rect 1800 9894 1812 9926
rect 2772 9926 2832 10168
rect 3792 10168 3802 10190
rect 3836 10720 3852 10744
rect 4810 10744 4870 10986
rect 5830 10986 5838 11014
rect 5872 11536 5890 11562
rect 6842 11562 6902 11804
rect 7864 11804 7874 11818
rect 7908 12356 7924 12380
rect 8884 12380 8944 12622
rect 9900 12622 9910 12650
rect 9944 13174 9958 13198
rect 10920 13198 10980 13440
rect 9944 12650 9950 13174
rect 10920 13170 10928 13198
rect 9944 12622 9960 12650
rect 9174 12572 9662 12578
rect 9174 12538 9186 12572
rect 9650 12538 9662 12572
rect 9174 12532 9662 12538
rect 9380 12470 9440 12532
rect 9174 12464 9662 12470
rect 9174 12430 9186 12464
rect 9650 12430 9662 12464
rect 9174 12424 9662 12430
rect 8884 12356 8892 12380
rect 7908 11818 7914 12356
rect 8886 11818 8892 12356
rect 7908 11804 7924 11818
rect 7138 11754 7626 11760
rect 7138 11720 7150 11754
rect 7614 11720 7626 11754
rect 7138 11714 7626 11720
rect 7340 11652 7400 11714
rect 7138 11646 7626 11652
rect 7138 11612 7150 11646
rect 7614 11612 7626 11646
rect 7138 11606 7626 11612
rect 5872 11014 5878 11536
rect 6842 11528 6856 11562
rect 5872 10986 5890 11014
rect 6850 11006 6856 11528
rect 5102 10936 5590 10942
rect 5102 10902 5114 10936
rect 5578 10902 5590 10936
rect 5102 10896 5590 10902
rect 5292 10834 5352 10896
rect 5102 10828 5590 10834
rect 5102 10794 5114 10828
rect 5578 10794 5590 10828
rect 5102 10788 5590 10794
rect 3836 10190 3842 10720
rect 4810 10716 4820 10744
rect 3836 10168 3852 10190
rect 4814 10186 4820 10716
rect 3066 10118 3554 10124
rect 3066 10084 3078 10118
rect 3542 10084 3554 10118
rect 3066 10078 3554 10084
rect 3272 10016 3332 10078
rect 3066 10010 3554 10016
rect 3066 9976 3078 10010
rect 3542 9976 3554 10010
rect 3066 9970 3554 9976
rect 2772 9898 2784 9926
rect 1800 9372 1806 9894
rect 2778 9376 2784 9898
rect 1800 9350 1812 9372
rect 1752 9108 1812 9350
rect 2772 9350 2784 9376
rect 2818 9898 2832 9926
rect 3792 9926 3852 10168
rect 4810 10168 4820 10186
rect 4854 10716 4870 10744
rect 5830 10744 5890 10986
rect 6842 10986 6856 11006
rect 6890 11528 6902 11562
rect 7864 11562 7924 11804
rect 8884 11804 8892 11818
rect 8926 12356 8944 12380
rect 9900 12380 9960 12622
rect 10922 12622 10928 13170
rect 10962 13170 10980 13198
rect 10962 12646 10968 13170
rect 10962 12622 10982 12646
rect 10192 12572 10680 12578
rect 10192 12538 10204 12572
rect 10668 12538 10680 12572
rect 10192 12532 10680 12538
rect 10400 12470 10460 12532
rect 10192 12464 10680 12470
rect 10192 12430 10204 12464
rect 10668 12430 10680 12464
rect 10192 12424 10680 12430
rect 9900 12360 9910 12380
rect 8926 11818 8932 12356
rect 9904 11822 9910 12360
rect 8926 11804 8944 11818
rect 8156 11754 8644 11760
rect 8156 11720 8168 11754
rect 8632 11720 8644 11754
rect 8156 11714 8644 11720
rect 8362 11652 8422 11714
rect 8156 11646 8644 11652
rect 8156 11612 8168 11646
rect 8632 11612 8644 11646
rect 8156 11606 8644 11612
rect 7864 11528 7874 11562
rect 6890 11006 6896 11528
rect 7868 11006 7874 11528
rect 6890 10986 6902 11006
rect 6120 10936 6608 10942
rect 6120 10902 6132 10936
rect 6596 10902 6608 10936
rect 6120 10896 6608 10902
rect 6322 10834 6382 10896
rect 6120 10828 6608 10834
rect 6120 10794 6132 10828
rect 6596 10794 6608 10828
rect 6120 10788 6608 10794
rect 5830 10724 5838 10744
rect 4854 10186 4860 10716
rect 5832 10194 5838 10724
rect 4854 10168 4870 10186
rect 4084 10118 4572 10124
rect 4084 10084 4096 10118
rect 4560 10084 4572 10118
rect 4084 10078 4572 10084
rect 4292 10016 4352 10078
rect 4084 10010 4572 10016
rect 4084 9976 4096 10010
rect 4560 9976 4572 10010
rect 4084 9970 4572 9976
rect 3792 9900 3802 9926
rect 2818 9376 2824 9898
rect 3796 9378 3802 9900
rect 2818 9350 2832 9376
rect 2048 9300 2536 9306
rect 2048 9266 2060 9300
rect 2524 9266 2536 9300
rect 2048 9260 2536 9266
rect 2260 9198 2320 9260
rect 2048 9192 2536 9198
rect 2048 9158 2060 9192
rect 2524 9158 2536 9192
rect 2048 9152 2536 9158
rect 1752 9082 1766 9108
rect 1760 8554 1766 9082
rect 1752 8532 1766 8554
rect 1800 9082 1812 9108
rect 2772 9108 2832 9350
rect 3792 9350 3802 9378
rect 3836 9900 3852 9926
rect 4810 9926 4870 10168
rect 5830 10168 5838 10194
rect 5872 10724 5890 10744
rect 6842 10744 6902 10986
rect 7864 10986 7874 11006
rect 7908 11528 7924 11562
rect 8884 11562 8944 11804
rect 9900 11804 9910 11822
rect 9944 12360 9960 12380
rect 10922 12380 10982 12622
rect 9944 11822 9950 12360
rect 9944 11804 9960 11822
rect 9174 11754 9662 11760
rect 9174 11720 9186 11754
rect 9650 11720 9662 11754
rect 9174 11714 9662 11720
rect 9374 11652 9434 11714
rect 9174 11646 9662 11652
rect 9174 11612 9186 11646
rect 9650 11612 9662 11646
rect 9174 11606 9662 11612
rect 8884 11528 8892 11562
rect 7908 11006 7914 11528
rect 8886 11006 8892 11528
rect 7908 10986 7924 11006
rect 7138 10936 7626 10942
rect 7138 10902 7150 10936
rect 7614 10902 7626 10936
rect 7138 10896 7626 10902
rect 7338 10834 7398 10896
rect 7138 10828 7626 10834
rect 7138 10794 7150 10828
rect 7614 10794 7626 10828
rect 7138 10788 7626 10794
rect 5872 10194 5878 10724
rect 6842 10716 6856 10744
rect 5872 10168 5890 10194
rect 6850 10186 6856 10716
rect 5102 10118 5590 10124
rect 5102 10084 5114 10118
rect 5578 10084 5590 10118
rect 5102 10078 5590 10084
rect 5294 10016 5354 10078
rect 5102 10010 5590 10016
rect 5102 9976 5114 10010
rect 5578 9976 5590 10010
rect 5102 9970 5590 9976
rect 3836 9378 3842 9900
rect 4810 9896 4820 9926
rect 3836 9350 3852 9378
rect 4814 9374 4820 9896
rect 3066 9300 3554 9306
rect 3066 9266 3078 9300
rect 3542 9266 3554 9300
rect 3066 9260 3554 9266
rect 3274 9198 3334 9260
rect 3066 9192 3554 9198
rect 3066 9158 3078 9192
rect 3542 9158 3554 9192
rect 3066 9152 3554 9158
rect 2772 9086 2784 9108
rect 1800 8554 1806 9082
rect 2778 8558 2784 9086
rect 1800 8532 1812 8554
rect 1752 8290 1812 8532
rect 2772 8532 2784 8558
rect 2818 9086 2832 9108
rect 3792 9108 3852 9350
rect 4810 9350 4820 9374
rect 4854 9896 4870 9926
rect 5830 9926 5890 10168
rect 6842 10168 6856 10186
rect 6890 10716 6902 10744
rect 7864 10744 7924 10986
rect 8884 10986 8892 11006
rect 8926 11528 8944 11562
rect 9900 11562 9960 11804
rect 10922 11804 10928 12380
rect 10962 12356 10982 12380
rect 10962 11818 10968 12356
rect 10962 11804 10982 11818
rect 10192 11754 10680 11760
rect 10192 11720 10204 11754
rect 10668 11720 10680 11754
rect 10192 11714 10680 11720
rect 10394 11652 10454 11714
rect 10192 11646 10680 11652
rect 10192 11612 10204 11646
rect 10668 11612 10680 11646
rect 10192 11606 10680 11612
rect 9900 11532 9910 11562
rect 8926 11006 8932 11528
rect 9904 11010 9910 11532
rect 8926 10986 8944 11006
rect 8156 10936 8644 10942
rect 8156 10902 8168 10936
rect 8632 10902 8644 10936
rect 8156 10896 8644 10902
rect 8360 10834 8420 10896
rect 8156 10828 8644 10834
rect 8156 10794 8168 10828
rect 8632 10794 8644 10828
rect 8156 10788 8644 10794
rect 7864 10716 7874 10744
rect 6890 10186 6896 10716
rect 7868 10186 7874 10716
rect 6890 10168 6902 10186
rect 6120 10118 6608 10124
rect 6120 10084 6132 10118
rect 6596 10084 6608 10118
rect 6120 10078 6608 10084
rect 6324 10016 6384 10078
rect 6120 10010 6608 10016
rect 6120 9976 6132 10010
rect 6596 9976 6608 10010
rect 6120 9970 6608 9976
rect 5830 9904 5838 9926
rect 4854 9374 4860 9896
rect 5832 9382 5838 9904
rect 4854 9350 4870 9374
rect 4084 9300 4572 9306
rect 4084 9266 4096 9300
rect 4560 9266 4572 9300
rect 4084 9260 4572 9266
rect 4294 9198 4354 9260
rect 4084 9192 4572 9198
rect 4084 9158 4096 9192
rect 4560 9158 4572 9192
rect 4084 9152 4572 9158
rect 3792 9088 3802 9108
rect 2818 8558 2824 9086
rect 3796 8560 3802 9088
rect 2818 8532 2832 8558
rect 2048 8482 2536 8488
rect 2048 8448 2060 8482
rect 2524 8448 2536 8482
rect 2048 8442 2536 8448
rect 2262 8380 2322 8442
rect 2048 8374 2536 8380
rect 2048 8340 2060 8374
rect 2524 8340 2536 8374
rect 2048 8334 2536 8340
rect 1752 8264 1766 8290
rect 1760 7714 1766 8264
rect 1800 8264 1812 8290
rect 2772 8290 2832 8532
rect 3792 8532 3802 8560
rect 3836 9088 3852 9108
rect 4810 9108 4870 9350
rect 5830 9350 5838 9382
rect 5872 9904 5890 9926
rect 6842 9926 6902 10168
rect 7864 10168 7874 10186
rect 7908 10716 7924 10744
rect 8884 10744 8944 10986
rect 9900 10986 9910 11010
rect 9944 11532 9960 11562
rect 10922 11562 10982 11804
rect 12800 11638 12860 14032
rect 13060 12758 13120 15132
rect 13060 12752 13122 12758
rect 13060 12692 13062 12752
rect 13060 12686 13122 12692
rect 12920 12480 12926 12540
rect 12986 12480 12992 12540
rect 12794 11578 12800 11638
rect 12860 11578 12866 11638
rect 9944 11010 9950 11532
rect 9944 10986 9960 11010
rect 9174 10936 9662 10942
rect 9174 10902 9186 10936
rect 9650 10902 9662 10936
rect 9174 10896 9662 10902
rect 9372 10834 9432 10896
rect 9174 10828 9662 10834
rect 9174 10794 9186 10828
rect 9650 10794 9662 10828
rect 9174 10788 9662 10794
rect 8884 10716 8892 10744
rect 7908 10186 7914 10716
rect 8886 10186 8892 10716
rect 7908 10168 7924 10186
rect 7138 10118 7626 10124
rect 7138 10084 7150 10118
rect 7614 10084 7626 10118
rect 7138 10078 7626 10084
rect 7340 10016 7400 10078
rect 7138 10010 7626 10016
rect 7138 9976 7150 10010
rect 7614 9976 7626 10010
rect 7138 9970 7626 9976
rect 5872 9382 5878 9904
rect 6842 9896 6856 9926
rect 5872 9350 5890 9382
rect 6850 9374 6856 9896
rect 5102 9300 5590 9306
rect 5102 9266 5114 9300
rect 5578 9266 5590 9300
rect 5102 9260 5590 9266
rect 5296 9198 5356 9260
rect 5102 9192 5590 9198
rect 5102 9158 5114 9192
rect 5578 9158 5590 9192
rect 5102 9152 5590 9158
rect 3836 8560 3842 9088
rect 4810 9084 4820 9108
rect 3836 8532 3852 8560
rect 4814 8556 4820 9084
rect 3066 8482 3554 8488
rect 3066 8448 3078 8482
rect 3542 8448 3554 8482
rect 3066 8442 3554 8448
rect 3276 8380 3336 8442
rect 3066 8374 3554 8380
rect 3066 8340 3078 8374
rect 3542 8340 3554 8374
rect 3066 8334 3554 8340
rect 2772 8268 2784 8290
rect 1800 7714 1806 8264
rect 1760 7702 1806 7714
rect 2778 7714 2784 8268
rect 2818 8268 2832 8290
rect 3792 8290 3852 8532
rect 4810 8532 4820 8556
rect 4854 9084 4870 9108
rect 5830 9108 5890 9350
rect 6842 9350 6856 9374
rect 6890 9896 6902 9926
rect 7864 9926 7924 10168
rect 8884 10168 8892 10186
rect 8926 10716 8944 10744
rect 9900 10744 9960 10986
rect 10922 10986 10928 11562
rect 10962 11528 10982 11562
rect 10962 11006 10968 11528
rect 10962 10986 10982 11006
rect 10192 10936 10680 10942
rect 10192 10902 10204 10936
rect 10668 10902 10680 10936
rect 10192 10896 10680 10902
rect 10392 10834 10452 10896
rect 10192 10828 10680 10834
rect 10192 10794 10204 10828
rect 10668 10794 10680 10828
rect 10192 10788 10680 10794
rect 9900 10720 9910 10744
rect 8926 10186 8932 10716
rect 9904 10190 9910 10720
rect 8926 10168 8944 10186
rect 8156 10118 8644 10124
rect 8156 10084 8168 10118
rect 8632 10084 8644 10118
rect 8156 10078 8644 10084
rect 8362 10016 8422 10078
rect 8156 10010 8644 10016
rect 8156 9976 8168 10010
rect 8632 9976 8644 10010
rect 8156 9970 8644 9976
rect 7864 9896 7874 9926
rect 6890 9374 6896 9896
rect 7868 9374 7874 9896
rect 6890 9350 6902 9374
rect 6120 9300 6608 9306
rect 6120 9266 6132 9300
rect 6596 9266 6608 9300
rect 6120 9260 6608 9266
rect 6326 9198 6386 9260
rect 6120 9192 6608 9198
rect 6120 9158 6132 9192
rect 6596 9158 6608 9192
rect 6120 9152 6608 9158
rect 5830 9092 5838 9108
rect 4854 8556 4860 9084
rect 5832 8564 5838 9092
rect 4854 8532 4870 8556
rect 4084 8482 4572 8488
rect 4084 8448 4096 8482
rect 4560 8448 4572 8482
rect 4084 8442 4572 8448
rect 4296 8380 4356 8442
rect 4084 8374 4572 8380
rect 4084 8340 4096 8374
rect 4560 8340 4572 8374
rect 4084 8334 4572 8340
rect 3792 8270 3802 8290
rect 2818 7714 2824 8268
rect 3796 7760 3802 8270
rect 2778 7702 2824 7714
rect 3786 7714 3802 7760
rect 3836 8270 3852 8290
rect 4810 8290 4870 8532
rect 5830 8532 5838 8564
rect 5872 9092 5890 9108
rect 6842 9108 6902 9350
rect 7864 9350 7874 9374
rect 7908 9896 7924 9926
rect 8884 9926 8944 10168
rect 9900 10168 9910 10190
rect 9944 10720 9960 10744
rect 10922 10744 10982 10986
rect 9944 10190 9950 10720
rect 9944 10168 9960 10190
rect 9174 10118 9662 10124
rect 9174 10084 9186 10118
rect 9650 10084 9662 10118
rect 9174 10078 9662 10084
rect 9374 10016 9434 10078
rect 9174 10010 9662 10016
rect 9174 9976 9186 10010
rect 9650 9976 9662 10010
rect 9174 9970 9662 9976
rect 8884 9896 8892 9926
rect 7908 9374 7914 9896
rect 8886 9374 8892 9896
rect 7908 9350 7924 9374
rect 7138 9300 7626 9306
rect 7138 9266 7150 9300
rect 7614 9266 7626 9300
rect 7138 9260 7626 9266
rect 7342 9198 7402 9260
rect 7138 9192 7626 9198
rect 7138 9158 7150 9192
rect 7614 9158 7626 9192
rect 7138 9152 7626 9158
rect 5872 8564 5878 9092
rect 6842 9084 6856 9108
rect 5872 8532 5890 8564
rect 6850 8556 6856 9084
rect 5102 8482 5590 8488
rect 5102 8448 5114 8482
rect 5578 8448 5590 8482
rect 5102 8442 5590 8448
rect 5298 8380 5358 8442
rect 5102 8374 5590 8380
rect 5102 8340 5114 8374
rect 5578 8340 5590 8374
rect 5102 8334 5590 8340
rect 3836 7760 3842 8270
rect 4810 8266 4820 8290
rect 3836 7714 3846 7760
rect 2048 7664 2536 7670
rect 2048 7630 2060 7664
rect 2524 7630 2536 7664
rect 2048 7624 2536 7630
rect 3066 7664 3554 7670
rect 3066 7630 3078 7664
rect 3542 7630 3554 7664
rect 3066 7624 3554 7630
rect 3786 7540 3846 7714
rect 4814 7714 4820 8266
rect 4854 8266 4870 8290
rect 5830 8290 5890 8532
rect 6842 8532 6856 8556
rect 6890 9084 6902 9108
rect 7864 9108 7924 9350
rect 8884 9350 8892 9374
rect 8926 9896 8944 9926
rect 9900 9926 9960 10168
rect 10922 10168 10928 10744
rect 10962 10716 10982 10744
rect 10962 10186 10968 10716
rect 10962 10168 10982 10186
rect 10192 10118 10680 10124
rect 10192 10084 10204 10118
rect 10668 10084 10680 10118
rect 10192 10078 10680 10084
rect 10394 10016 10454 10078
rect 10192 10010 10680 10016
rect 10192 9976 10204 10010
rect 10668 9976 10680 10010
rect 10192 9970 10680 9976
rect 9900 9900 9910 9926
rect 8926 9374 8932 9896
rect 9904 9378 9910 9900
rect 8926 9350 8944 9374
rect 8156 9300 8644 9306
rect 8156 9266 8168 9300
rect 8632 9266 8644 9300
rect 8156 9260 8644 9266
rect 8364 9198 8424 9260
rect 8156 9192 8644 9198
rect 8156 9158 8168 9192
rect 8632 9158 8644 9192
rect 8156 9152 8644 9158
rect 7864 9084 7874 9108
rect 6890 8556 6896 9084
rect 7868 8556 7874 9084
rect 6890 8532 6902 8556
rect 6120 8482 6608 8488
rect 6120 8448 6132 8482
rect 6596 8448 6608 8482
rect 6120 8442 6608 8448
rect 6328 8380 6388 8442
rect 6120 8374 6608 8380
rect 6120 8340 6132 8374
rect 6596 8340 6608 8374
rect 6120 8334 6608 8340
rect 5830 8274 5838 8290
rect 4854 7714 4860 8266
rect 5832 7762 5838 8274
rect 4814 7702 4860 7714
rect 5824 7714 5838 7762
rect 5872 8274 5890 8290
rect 6842 8290 6902 8532
rect 7864 8532 7874 8556
rect 7908 9084 7924 9108
rect 8884 9108 8944 9350
rect 9900 9350 9910 9378
rect 9944 9900 9960 9926
rect 10922 9926 10982 10168
rect 9944 9378 9950 9900
rect 9944 9350 9960 9378
rect 9174 9300 9662 9306
rect 9174 9266 9186 9300
rect 9650 9266 9662 9300
rect 9174 9260 9662 9266
rect 9376 9198 9436 9260
rect 9174 9192 9662 9198
rect 9174 9158 9186 9192
rect 9650 9158 9662 9192
rect 9174 9152 9662 9158
rect 8884 9084 8892 9108
rect 7908 8556 7914 9084
rect 8886 8556 8892 9084
rect 7908 8532 7924 8556
rect 7138 8482 7626 8488
rect 7138 8448 7150 8482
rect 7614 8448 7626 8482
rect 7138 8442 7626 8448
rect 7344 8380 7404 8442
rect 7138 8374 7626 8380
rect 7138 8340 7150 8374
rect 7614 8340 7626 8374
rect 7138 8334 7626 8340
rect 5872 7762 5878 8274
rect 6842 8266 6856 8290
rect 5872 7714 5884 7762
rect 4084 7664 4572 7670
rect 4084 7630 4096 7664
rect 4560 7630 4572 7664
rect 4084 7624 4572 7630
rect 5102 7664 5590 7670
rect 5102 7630 5114 7664
rect 5578 7630 5590 7664
rect 5102 7624 5590 7630
rect 5824 7540 5884 7714
rect 6850 7714 6856 8266
rect 6890 8266 6902 8290
rect 7864 8290 7924 8532
rect 8884 8532 8892 8556
rect 8926 9084 8944 9108
rect 9900 9108 9960 9350
rect 10922 9350 10928 9926
rect 10962 9896 10982 9926
rect 10962 9374 10968 9896
rect 10962 9350 10982 9374
rect 10192 9300 10680 9306
rect 10192 9266 10204 9300
rect 10668 9266 10680 9300
rect 10192 9260 10680 9266
rect 10396 9198 10456 9260
rect 10192 9192 10680 9198
rect 10192 9158 10204 9192
rect 10668 9158 10680 9192
rect 10192 9152 10680 9158
rect 9900 9088 9910 9108
rect 8926 8556 8932 9084
rect 9904 8560 9910 9088
rect 8926 8532 8944 8556
rect 8156 8482 8644 8488
rect 8156 8448 8168 8482
rect 8632 8448 8644 8482
rect 8156 8442 8644 8448
rect 8366 8380 8426 8442
rect 8156 8374 8644 8380
rect 8156 8340 8168 8374
rect 8632 8340 8644 8374
rect 8156 8334 8644 8340
rect 7864 8266 7874 8290
rect 6890 7714 6896 8266
rect 7868 7758 7874 8266
rect 6850 7702 6896 7714
rect 7860 7714 7874 7758
rect 7908 8266 7924 8290
rect 8884 8290 8944 8532
rect 9900 8532 9910 8560
rect 9944 9088 9960 9108
rect 10922 9108 10982 9350
rect 9944 8560 9950 9088
rect 9944 8532 9960 8560
rect 9174 8482 9662 8488
rect 9174 8448 9186 8482
rect 9650 8448 9662 8482
rect 9174 8442 9662 8448
rect 9378 8380 9438 8442
rect 9174 8374 9662 8380
rect 9174 8340 9186 8374
rect 9650 8340 9662 8374
rect 9174 8334 9662 8340
rect 8884 8266 8892 8290
rect 7908 7758 7914 8266
rect 7908 7714 7920 7758
rect 6120 7664 6608 7670
rect 6120 7630 6132 7664
rect 6596 7630 6608 7664
rect 6120 7624 6608 7630
rect 7138 7664 7626 7670
rect 7138 7630 7150 7664
rect 7614 7630 7626 7664
rect 7138 7624 7626 7630
rect 7860 7540 7920 7714
rect 8886 7714 8892 8266
rect 8926 8266 8944 8290
rect 9900 8290 9960 8532
rect 10922 8532 10928 9108
rect 10962 9084 10982 9108
rect 10962 8556 10968 9084
rect 10962 8532 10982 8556
rect 10192 8482 10680 8488
rect 10192 8448 10204 8482
rect 10668 8448 10680 8482
rect 10192 8442 10680 8448
rect 10398 8380 10458 8442
rect 10192 8374 10680 8380
rect 10192 8340 10204 8374
rect 10668 8340 10680 8374
rect 10192 8334 10680 8340
rect 9900 8270 9910 8290
rect 8926 7714 8932 8266
rect 9904 7756 9910 8270
rect 8886 7702 8932 7714
rect 9896 7714 9910 7756
rect 9944 8270 9960 8290
rect 10922 8290 10982 8532
rect 9944 7756 9950 8270
rect 10922 7768 10928 8290
rect 9944 7714 9956 7756
rect 8156 7664 8644 7670
rect 8156 7630 8168 7664
rect 8632 7630 8644 7664
rect 8156 7624 8644 7630
rect 9174 7664 9662 7670
rect 9174 7630 9186 7664
rect 9650 7630 9662 7664
rect 9174 7624 9662 7630
rect 9896 7540 9956 7714
rect 10916 7714 10928 7768
rect 10962 8266 10982 8290
rect 10962 7768 10968 8266
rect 10962 7714 10976 7768
rect 10192 7664 10680 7670
rect 10192 7630 10204 7664
rect 10668 7630 10680 7664
rect 10192 7624 10680 7630
rect 10410 7540 10470 7624
rect 10916 7540 10976 7714
rect 11902 7682 11962 7688
rect 3786 7480 10976 7540
rect 11640 7652 11700 7674
rect 7968 6320 7974 6380
rect 8034 6320 8040 6380
rect 1534 4926 2612 4986
rect 1534 4747 1594 4926
rect 2048 4837 2108 4926
rect 1827 4831 2315 4837
rect 1827 4797 1839 4831
rect 2303 4797 2315 4831
rect 1827 4791 2315 4797
rect 1534 4702 1545 4747
rect 1539 4171 1545 4702
rect 1579 4702 1594 4747
rect 2552 4747 2612 4926
rect 3558 4880 3564 4940
rect 3624 4880 3630 4940
rect 3944 4926 5154 4986
rect 7974 4984 8034 6320
rect 2845 4831 3333 4837
rect 2845 4797 2857 4831
rect 3321 4797 3333 4831
rect 2845 4791 3333 4797
rect 1579 4171 1585 4702
rect 2552 4698 2563 4747
rect 2557 4216 2563 4698
rect 1539 4159 1585 4171
rect 2550 4171 2563 4216
rect 2597 4698 2612 4747
rect 3564 4747 3624 4880
rect 4072 4837 4132 4926
rect 3863 4831 4351 4837
rect 3863 4797 3875 4831
rect 4339 4797 4351 4831
rect 3863 4791 4351 4797
rect 2597 4216 2603 4698
rect 2597 4171 2610 4216
rect 1827 4121 2315 4127
rect 1827 4087 1839 4121
rect 2303 4087 2315 4121
rect 1827 4081 2315 4087
rect 2550 4036 2610 4171
rect 3564 4171 3581 4747
rect 3615 4171 3624 4747
rect 4588 4747 4648 4926
rect 5094 4837 5154 4926
rect 5598 4880 5604 4940
rect 5664 4880 5670 4940
rect 6624 4924 8034 4984
rect 4881 4831 5369 4837
rect 4881 4797 4893 4831
rect 5357 4797 5369 4831
rect 4881 4791 5369 4797
rect 4588 4690 4599 4747
rect 4593 4212 4599 4690
rect 2845 4121 3333 4127
rect 2845 4087 2857 4121
rect 3321 4087 3333 4121
rect 2845 4081 3333 4087
rect 1406 3976 1412 4036
rect 1472 3976 1478 4036
rect 2544 3976 2550 4036
rect 2610 3976 2616 4036
rect 1412 1614 1472 3976
rect 1532 3760 2608 3820
rect 1532 3634 1592 3760
rect 2042 3724 2102 3760
rect 1826 3718 2314 3724
rect 1826 3684 1838 3718
rect 2302 3684 2314 3718
rect 1826 3678 2314 3684
rect 1532 3574 1544 3634
rect 1538 3058 1544 3574
rect 1578 3574 1592 3634
rect 2548 3634 2608 3760
rect 3060 3724 3120 4081
rect 3564 3940 3624 4171
rect 4586 4171 4599 4212
rect 4633 4690 4648 4747
rect 5604 4747 5664 4880
rect 5899 4831 6387 4837
rect 5899 4797 5911 4831
rect 6375 4797 6387 4831
rect 5899 4791 6387 4797
rect 5604 4702 5617 4747
rect 4633 4212 4639 4690
rect 4633 4171 4646 4212
rect 5611 4210 5617 4702
rect 3863 4121 4351 4127
rect 3863 4087 3875 4121
rect 4339 4087 4351 4121
rect 3863 4081 4351 4087
rect 3558 3880 3564 3940
rect 3624 3880 3630 3940
rect 2844 3718 3332 3724
rect 2844 3684 2856 3718
rect 3320 3684 3332 3718
rect 2844 3678 3332 3684
rect 2548 3588 2562 3634
rect 1578 3058 1584 3574
rect 2556 3104 2562 3588
rect 1538 3046 1584 3058
rect 2548 3058 2562 3104
rect 2596 3588 2608 3634
rect 3564 3634 3624 3880
rect 4080 3724 4140 4081
rect 4586 3824 4646 4171
rect 5604 4171 5617 4210
rect 5651 4702 5664 4747
rect 6624 4747 6684 4924
rect 7132 4837 7192 4924
rect 6917 4831 7405 4837
rect 6917 4797 6929 4831
rect 7393 4797 7405 4831
rect 6917 4791 7405 4797
rect 5651 4210 5657 4702
rect 6624 4694 6635 4747
rect 6629 4216 6635 4694
rect 5651 4171 5664 4210
rect 4881 4121 5369 4127
rect 4881 4087 4893 4121
rect 5357 4087 5369 4121
rect 4881 4081 5369 4087
rect 4580 3764 4586 3824
rect 4646 3764 4652 3824
rect 5088 3724 5148 4081
rect 5604 3940 5664 4171
rect 6624 4171 6635 4216
rect 6669 4694 6684 4747
rect 7640 4747 7700 4924
rect 7640 4700 7653 4747
rect 6669 4216 6675 4694
rect 6669 4171 6684 4216
rect 5899 4121 6387 4127
rect 5899 4087 5911 4121
rect 6375 4087 6387 4121
rect 5899 4081 6387 4087
rect 5598 3880 5604 3940
rect 5664 3880 5670 3940
rect 3862 3718 4350 3724
rect 3862 3684 3874 3718
rect 4338 3684 4350 3718
rect 3862 3678 4350 3684
rect 4880 3718 5368 3724
rect 4880 3684 4892 3718
rect 5356 3684 5368 3718
rect 4880 3678 5368 3684
rect 3564 3588 3580 3634
rect 2596 3104 2602 3588
rect 2596 3058 2608 3104
rect 3574 3100 3580 3588
rect 1826 3008 2314 3014
rect 1826 2974 1838 3008
rect 2302 2974 2314 3008
rect 1826 2968 2314 2974
rect 2548 2816 2608 3058
rect 3566 3058 3580 3100
rect 3614 3588 3624 3634
rect 4592 3634 4638 3646
rect 3614 3100 3620 3588
rect 4592 3110 4598 3634
rect 3614 3058 3626 3100
rect 2844 3008 3332 3014
rect 2844 2974 2856 3008
rect 3320 2974 3332 3008
rect 2844 2968 3332 2974
rect 2690 2864 2696 2924
rect 2756 2864 2762 2924
rect 2542 2756 2548 2816
rect 2608 2756 2614 2816
rect 2696 2714 2756 2864
rect 1532 2654 2756 2714
rect 1532 2523 1592 2654
rect 2048 2613 2108 2654
rect 1827 2607 2315 2613
rect 1827 2573 1839 2607
rect 2303 2573 2315 2607
rect 1827 2567 2315 2573
rect 1532 2482 1545 2523
rect 1539 1947 1545 2482
rect 1579 2482 1592 2523
rect 2550 2523 2610 2654
rect 3066 2613 3126 2968
rect 3566 2704 3626 3058
rect 4582 3058 4598 3110
rect 4632 3110 4638 3634
rect 5604 3634 5664 3880
rect 6110 3724 6170 4081
rect 6624 4036 6684 4171
rect 7647 4171 7653 4700
rect 7687 4700 7700 4747
rect 7687 4171 7693 4700
rect 7647 4159 7693 4171
rect 6917 4121 7405 4127
rect 6917 4087 6929 4121
rect 7393 4087 7405 4121
rect 6917 4081 7405 4087
rect 6618 3976 6624 4036
rect 6684 3976 6690 4036
rect 8104 3930 8164 7480
rect 10130 7356 10136 7416
rect 10196 7356 10202 7416
rect 11042 7356 11048 7416
rect 11108 7356 11114 7416
rect 9260 7246 9266 7306
rect 9326 7246 9332 7306
rect 8346 7138 8352 7198
rect 8412 7138 8418 7198
rect 8352 5644 8412 7138
rect 8476 7030 8482 7090
rect 8542 7030 8548 7090
rect 8482 5766 8542 7030
rect 8708 6990 8796 6996
rect 8708 6956 8720 6990
rect 8784 6956 8796 6990
rect 8708 6950 8796 6956
rect 8926 6990 9014 6996
rect 8926 6956 8938 6990
rect 9002 6956 9014 6990
rect 8926 6950 9014 6956
rect 9144 6990 9232 6996
rect 9144 6956 9156 6990
rect 9220 6956 9232 6990
rect 9144 6950 9232 6956
rect 8620 6906 8666 6918
rect 8620 6760 8626 6906
rect 8612 6730 8626 6760
rect 8660 6760 8666 6906
rect 8838 6906 8884 6918
rect 8660 6730 8672 6760
rect 8838 6752 8844 6906
rect 8612 6580 8672 6730
rect 8832 6730 8844 6752
rect 8878 6752 8884 6906
rect 9056 6906 9102 6918
rect 8878 6730 8892 6752
rect 9056 6742 9062 6906
rect 8708 6680 8796 6686
rect 8708 6646 8720 6680
rect 8784 6646 8796 6680
rect 8708 6640 8796 6646
rect 8720 6580 8780 6640
rect 8832 6580 8892 6730
rect 9048 6730 9062 6742
rect 9096 6742 9102 6906
rect 9266 6906 9326 7246
rect 10024 7138 10030 7198
rect 10090 7138 10096 7198
rect 9806 7030 9812 7090
rect 9872 7030 9878 7090
rect 9812 6996 9872 7030
rect 10030 6996 10090 7138
rect 9362 6990 9450 6996
rect 9362 6956 9374 6990
rect 9438 6956 9450 6990
rect 9362 6950 9450 6956
rect 9580 6990 9668 6996
rect 9580 6956 9592 6990
rect 9656 6956 9668 6990
rect 9580 6950 9668 6956
rect 9798 6990 9886 6996
rect 9798 6956 9810 6990
rect 9874 6956 9886 6990
rect 9798 6950 9886 6956
rect 10016 6990 10104 6996
rect 10016 6956 10028 6990
rect 10092 6956 10104 6990
rect 10016 6950 10104 6956
rect 9266 6890 9280 6906
rect 9096 6730 9108 6742
rect 8926 6680 9014 6686
rect 8926 6646 8938 6680
rect 9002 6646 9014 6680
rect 8926 6640 9014 6646
rect 8940 6590 9000 6640
rect 8612 6520 8892 6580
rect 8934 6530 8940 6590
rect 9000 6530 9006 6590
rect 8832 6262 8892 6520
rect 9048 6490 9108 6730
rect 9274 6730 9280 6890
rect 9314 6890 9326 6906
rect 9492 6906 9538 6918
rect 9314 6730 9320 6890
rect 9492 6756 9498 6906
rect 9274 6718 9320 6730
rect 9486 6730 9498 6756
rect 9532 6756 9538 6906
rect 9710 6906 9756 6918
rect 9710 6766 9716 6906
rect 9532 6730 9546 6756
rect 9144 6680 9232 6686
rect 9144 6646 9156 6680
rect 9220 6646 9232 6680
rect 9144 6640 9232 6646
rect 9362 6680 9450 6686
rect 9362 6646 9374 6680
rect 9438 6646 9450 6680
rect 9362 6640 9450 6646
rect 9042 6430 9048 6490
rect 9108 6430 9114 6490
rect 9044 6320 9050 6380
rect 9110 6320 9116 6380
rect 8614 6202 8892 6262
rect 8614 6074 8674 6202
rect 8724 6164 8784 6202
rect 8708 6158 8796 6164
rect 8708 6124 8720 6158
rect 8784 6124 8796 6158
rect 8708 6118 8796 6124
rect 8614 6048 8626 6074
rect 8620 5898 8626 6048
rect 8660 6048 8674 6074
rect 8832 6074 8892 6202
rect 8926 6158 9014 6164
rect 8926 6124 8938 6158
rect 9002 6124 9014 6158
rect 8926 6118 9014 6124
rect 8660 5898 8666 6048
rect 8620 5886 8666 5898
rect 8832 5898 8844 6074
rect 8878 5898 8892 6074
rect 9050 6074 9110 6320
rect 9158 6270 9218 6640
rect 9378 6270 9438 6640
rect 9486 6490 9546 6730
rect 9702 6730 9716 6766
rect 9750 6766 9756 6906
rect 9928 6906 9974 6918
rect 9750 6730 9762 6766
rect 9928 6764 9934 6906
rect 9580 6680 9668 6686
rect 9580 6646 9592 6680
rect 9656 6646 9668 6680
rect 9580 6640 9668 6646
rect 9596 6590 9656 6640
rect 9590 6530 9596 6590
rect 9656 6530 9662 6590
rect 9480 6430 9486 6490
rect 9546 6430 9552 6490
rect 9478 6320 9484 6380
rect 9544 6320 9550 6380
rect 9152 6210 9158 6270
rect 9218 6210 9224 6270
rect 9372 6210 9378 6270
rect 9438 6210 9444 6270
rect 9158 6164 9218 6210
rect 9378 6164 9438 6210
rect 9144 6158 9232 6164
rect 9144 6124 9156 6158
rect 9220 6124 9232 6158
rect 9144 6118 9232 6124
rect 9362 6158 9450 6164
rect 9362 6124 9374 6158
rect 9438 6124 9450 6158
rect 9362 6118 9450 6124
rect 9050 6038 9062 6074
rect 8708 5848 8796 5854
rect 8708 5814 8720 5848
rect 8784 5814 8796 5848
rect 8708 5808 8796 5814
rect 8476 5706 8482 5766
rect 8542 5706 8548 5766
rect 8346 5584 8352 5644
rect 8412 5584 8418 5644
rect 8832 5520 8892 5898
rect 9056 5898 9062 6038
rect 9096 6038 9110 6074
rect 9274 6074 9320 6086
rect 9096 5898 9102 6038
rect 9274 5938 9280 6074
rect 9056 5886 9102 5898
rect 9270 5898 9280 5938
rect 9314 5938 9320 6074
rect 9484 6074 9544 6320
rect 9580 6158 9668 6164
rect 9580 6124 9592 6158
rect 9656 6124 9668 6158
rect 9580 6118 9668 6124
rect 9484 6044 9498 6074
rect 9314 5898 9330 5938
rect 8926 5848 9014 5854
rect 8926 5814 8938 5848
rect 9002 5814 9014 5848
rect 8926 5808 9014 5814
rect 9144 5848 9232 5854
rect 9144 5814 9156 5848
rect 9220 5814 9232 5848
rect 9144 5808 9232 5814
rect 8940 5766 9000 5808
rect 8934 5706 8940 5766
rect 9000 5706 9006 5766
rect 9158 5644 9218 5808
rect 9152 5584 9158 5644
rect 9218 5584 9224 5644
rect 8826 5460 8832 5520
rect 8892 5460 8898 5520
rect 9270 5394 9330 5898
rect 9492 5898 9498 6044
rect 9532 6044 9544 6074
rect 9702 6074 9762 6730
rect 9922 6730 9934 6764
rect 9968 6764 9974 6906
rect 10136 6906 10196 7356
rect 10922 7246 10928 7306
rect 10988 7246 10994 7306
rect 10242 7138 10248 7198
rect 10308 7138 10314 7198
rect 10248 6996 10308 7138
rect 10460 7030 10466 7090
rect 10526 7030 10532 7090
rect 10466 6996 10526 7030
rect 10234 6990 10322 6996
rect 10234 6956 10246 6990
rect 10310 6956 10322 6990
rect 10234 6950 10322 6956
rect 10452 6990 10540 6996
rect 10452 6956 10464 6990
rect 10528 6956 10540 6990
rect 10452 6950 10540 6956
rect 10670 6990 10758 6996
rect 10670 6956 10682 6990
rect 10746 6956 10758 6990
rect 10670 6950 10758 6956
rect 10136 6860 10152 6906
rect 9968 6730 9982 6764
rect 9798 6680 9886 6686
rect 9798 6646 9810 6680
rect 9874 6646 9886 6680
rect 9798 6640 9886 6646
rect 9922 6490 9982 6730
rect 10146 6730 10152 6860
rect 10186 6860 10196 6906
rect 10364 6906 10410 6918
rect 10186 6730 10192 6860
rect 10364 6756 10370 6906
rect 10146 6718 10192 6730
rect 10358 6730 10370 6756
rect 10404 6756 10410 6906
rect 10582 6906 10628 6918
rect 10404 6730 10418 6756
rect 10582 6748 10588 6906
rect 10016 6680 10104 6686
rect 10016 6646 10028 6680
rect 10092 6646 10104 6680
rect 10016 6640 10104 6646
rect 10234 6680 10322 6686
rect 10234 6646 10246 6680
rect 10310 6646 10322 6680
rect 10234 6640 10322 6646
rect 10358 6490 10418 6730
rect 10576 6730 10588 6748
rect 10622 6748 10628 6906
rect 10800 6906 10846 6918
rect 10800 6766 10806 6906
rect 10622 6730 10636 6748
rect 10452 6680 10540 6686
rect 10452 6646 10464 6680
rect 10528 6646 10540 6680
rect 10452 6640 10540 6646
rect 10460 6530 10466 6590
rect 10526 6530 10532 6590
rect 10576 6588 10636 6730
rect 10794 6730 10806 6766
rect 10840 6766 10846 6906
rect 10928 6816 10988 7246
rect 10840 6730 10854 6766
rect 10670 6680 10758 6686
rect 10670 6646 10682 6680
rect 10746 6646 10758 6680
rect 10670 6640 10758 6646
rect 10684 6588 10744 6640
rect 10794 6588 10854 6730
rect 9812 6430 10418 6490
rect 9812 6380 9872 6430
rect 9806 6320 9812 6380
rect 9872 6320 9878 6380
rect 9916 6320 9922 6380
rect 9982 6320 9988 6380
rect 10352 6320 10358 6380
rect 10418 6320 10424 6380
rect 9798 6158 9886 6164
rect 9798 6124 9810 6158
rect 9874 6124 9886 6158
rect 9798 6118 9886 6124
rect 9532 5898 9538 6044
rect 9492 5886 9538 5898
rect 9702 5898 9716 6074
rect 9750 5898 9762 6074
rect 9922 6074 9982 6320
rect 10026 6210 10032 6270
rect 10092 6210 10098 6270
rect 10242 6210 10248 6270
rect 10308 6210 10314 6270
rect 10032 6164 10092 6210
rect 10248 6164 10308 6210
rect 10016 6158 10104 6164
rect 10016 6124 10028 6158
rect 10092 6124 10104 6158
rect 10016 6118 10104 6124
rect 10234 6158 10322 6164
rect 10234 6124 10246 6158
rect 10310 6124 10322 6158
rect 10234 6118 10322 6124
rect 9922 6056 9934 6074
rect 9362 5848 9450 5854
rect 9362 5814 9374 5848
rect 9438 5814 9450 5848
rect 9362 5808 9450 5814
rect 9580 5848 9668 5854
rect 9580 5814 9592 5848
rect 9656 5814 9668 5848
rect 9580 5808 9668 5814
rect 9376 5644 9436 5808
rect 9596 5766 9656 5808
rect 9590 5706 9596 5766
rect 9656 5706 9662 5766
rect 9370 5584 9376 5644
rect 9436 5584 9442 5644
rect 9264 5334 9270 5394
rect 9330 5334 9336 5394
rect 9606 5280 9654 5706
rect 9702 5520 9762 5898
rect 9928 5898 9934 6056
rect 9968 6056 9982 6074
rect 10146 6074 10192 6086
rect 9968 5898 9974 6056
rect 10146 5920 10152 6074
rect 9928 5886 9974 5898
rect 10140 5898 10152 5920
rect 10186 5920 10192 6074
rect 10358 6074 10418 6320
rect 10466 6164 10526 6530
rect 10576 6528 10854 6588
rect 10576 6470 10636 6528
rect 10570 6410 10576 6470
rect 10636 6410 10642 6470
rect 10576 6272 10636 6410
rect 10576 6212 10854 6272
rect 10452 6158 10540 6164
rect 10452 6124 10464 6158
rect 10528 6124 10540 6158
rect 10452 6118 10540 6124
rect 10358 6042 10370 6074
rect 10186 5898 10200 5920
rect 9798 5848 9886 5854
rect 9798 5814 9810 5848
rect 9874 5814 9886 5848
rect 9798 5808 9886 5814
rect 10016 5848 10104 5854
rect 10016 5814 10028 5848
rect 10092 5814 10104 5848
rect 10016 5808 10104 5814
rect 9812 5646 9872 5808
rect 10140 5766 10200 5898
rect 10364 5898 10370 6042
rect 10404 6042 10418 6074
rect 10576 6074 10636 6212
rect 10684 6164 10744 6212
rect 10670 6158 10758 6164
rect 10670 6124 10682 6158
rect 10746 6124 10758 6158
rect 10670 6118 10758 6124
rect 10576 6056 10588 6074
rect 10404 5898 10410 6042
rect 10582 5928 10588 6056
rect 10364 5886 10410 5898
rect 10574 5898 10588 5928
rect 10622 6056 10636 6074
rect 10794 6074 10854 6212
rect 10622 5928 10628 6056
rect 10794 6054 10806 6074
rect 10622 5898 10634 5928
rect 10234 5848 10322 5854
rect 10234 5814 10246 5848
rect 10310 5814 10322 5848
rect 10234 5808 10322 5814
rect 10452 5848 10540 5854
rect 10452 5814 10464 5848
rect 10528 5814 10540 5848
rect 10452 5808 10540 5814
rect 10134 5706 10140 5766
rect 10200 5706 10206 5766
rect 10468 5646 10528 5808
rect 9806 5586 9812 5646
rect 9872 5586 9878 5646
rect 10462 5586 10468 5646
rect 10528 5586 10534 5646
rect 10574 5520 10634 5898
rect 10800 5898 10806 6054
rect 10840 6054 10854 6074
rect 10840 5898 10846 6054
rect 10800 5886 10846 5898
rect 10670 5848 10758 5854
rect 10670 5814 10682 5848
rect 10746 5814 10758 5848
rect 10670 5808 10758 5814
rect 10928 5766 10988 6756
rect 10922 5706 10928 5766
rect 10988 5706 10994 5766
rect 9696 5460 9702 5520
rect 9762 5460 9768 5520
rect 10568 5460 10574 5520
rect 10634 5460 10640 5520
rect 11048 5394 11108 7356
rect 11164 6530 11170 6590
rect 11230 6530 11236 6590
rect 11170 6344 11230 6530
rect 11170 6276 11230 6284
rect 11042 5334 11048 5394
rect 11108 5334 11114 5394
rect 9598 5228 9604 5280
rect 9656 5228 9662 5280
rect 8274 5144 8280 5204
rect 8340 5144 8346 5204
rect 11640 5200 11700 7592
rect 8280 4960 8340 5144
rect 8412 5140 11700 5200
rect 8274 4900 8280 4960
rect 8340 4900 8346 4960
rect 6622 3870 8164 3930
rect 5898 3718 6386 3724
rect 5898 3684 5910 3718
rect 6374 3684 6386 3718
rect 5898 3678 6386 3684
rect 5604 3600 5616 3634
rect 4632 3058 4642 3110
rect 5610 3092 5616 3600
rect 3862 3008 4350 3014
rect 3862 2974 3874 3008
rect 4338 2974 4350 3008
rect 3862 2968 4350 2974
rect 3560 2644 3566 2704
rect 3626 2644 3632 2704
rect 2845 2607 3333 2613
rect 2845 2573 2857 2607
rect 3321 2573 3333 2607
rect 2845 2567 3333 2573
rect 2550 2482 2563 2523
rect 1579 1947 1585 2482
rect 1539 1935 1585 1947
rect 2557 1947 2563 2482
rect 2597 2482 2610 2523
rect 3566 2523 3626 2644
rect 4080 2613 4140 2968
rect 4582 2924 4642 3058
rect 5606 3058 5616 3092
rect 5650 3600 5664 3634
rect 6622 3634 6682 3870
rect 7132 3724 7192 3870
rect 6916 3718 7404 3724
rect 6916 3684 6928 3718
rect 7392 3684 7404 3718
rect 6916 3678 7404 3684
rect 7638 3634 7698 3870
rect 7742 3764 7748 3824
rect 7808 3764 7814 3824
rect 5650 3092 5656 3600
rect 6622 3588 6634 3634
rect 6624 3586 6634 3588
rect 6628 3096 6634 3586
rect 5650 3058 5666 3092
rect 4880 3008 5368 3014
rect 4880 2974 4892 3008
rect 5356 2974 5368 3008
rect 4880 2968 5368 2974
rect 4576 2864 4582 2924
rect 4642 2864 4648 2924
rect 4578 2756 4584 2816
rect 4644 2756 4650 2816
rect 3863 2607 4351 2613
rect 3863 2573 3875 2607
rect 4339 2573 4351 2607
rect 3863 2567 4351 2573
rect 3566 2494 3581 2523
rect 2597 1947 2603 2482
rect 3575 1984 3581 2494
rect 2557 1935 2603 1947
rect 3568 1947 3581 1984
rect 3615 2494 3626 2523
rect 4584 2523 4644 2756
rect 5108 2613 5168 2968
rect 5606 2710 5666 3058
rect 6620 3058 6634 3096
rect 6668 3586 6684 3634
rect 7638 3604 7652 3634
rect 7640 3602 7652 3604
rect 6668 3096 6674 3586
rect 6668 3058 6680 3096
rect 5898 3008 6386 3014
rect 5898 2974 5910 3008
rect 6374 2974 6386 3008
rect 5898 2968 6386 2974
rect 5604 2704 5666 2710
rect 5664 2644 5666 2704
rect 5604 2638 5666 2644
rect 4881 2607 5369 2613
rect 4881 2573 4893 2607
rect 5357 2573 5369 2607
rect 4881 2567 5369 2573
rect 3615 1984 3621 2494
rect 4584 2480 4599 2523
rect 3615 1947 3628 1984
rect 1827 1897 2315 1903
rect 1827 1863 1839 1897
rect 2303 1863 2315 1897
rect 1827 1857 2315 1863
rect 2845 1897 3333 1903
rect 2845 1863 2857 1897
rect 3321 1863 3333 1897
rect 2845 1857 3333 1863
rect 2544 1660 2550 1720
rect 2610 1660 2616 1720
rect 1406 1554 1412 1614
rect 1472 1554 1478 1614
rect 1826 1494 2314 1500
rect 1826 1460 1838 1494
rect 2302 1460 2314 1494
rect 1826 1454 2314 1460
rect 1538 1410 1584 1422
rect 1538 874 1544 1410
rect 1532 834 1544 874
rect 1578 874 1584 1410
rect 2550 1410 2610 1660
rect 3074 1500 3134 1857
rect 3568 1822 3628 1947
rect 4593 1947 4599 2480
rect 4633 2480 4644 2523
rect 5606 2523 5666 2638
rect 6118 2613 6178 2968
rect 6446 2864 6452 2924
rect 6512 2864 6518 2924
rect 6452 2714 6512 2864
rect 6620 2816 6680 3058
rect 7646 3058 7652 3602
rect 7686 3602 7700 3634
rect 7686 3058 7692 3602
rect 7646 3046 7692 3058
rect 6916 3008 7404 3014
rect 6916 2974 6928 3008
rect 7392 2974 7404 3008
rect 6916 2968 7404 2974
rect 6614 2756 6620 2816
rect 6680 2756 6686 2816
rect 6452 2654 7696 2714
rect 5899 2607 6387 2613
rect 5899 2573 5911 2607
rect 6375 2573 6387 2607
rect 5899 2567 6387 2573
rect 5606 2486 5617 2523
rect 4633 1947 4639 2480
rect 5611 1980 5617 2486
rect 4593 1935 4639 1947
rect 5602 1947 5617 1980
rect 5651 2486 5666 2523
rect 6622 2523 6682 2654
rect 7140 2613 7200 2654
rect 6917 2607 7405 2613
rect 6917 2573 6929 2607
rect 7393 2573 7405 2607
rect 6917 2567 7405 2573
rect 5651 1980 5657 2486
rect 6622 2482 6635 2523
rect 5651 1947 5662 1980
rect 3863 1897 4351 1903
rect 3863 1863 3875 1897
rect 4339 1863 4351 1897
rect 3863 1857 4351 1863
rect 4881 1897 5369 1903
rect 4881 1863 4893 1897
rect 5357 1863 5369 1897
rect 4881 1857 5369 1863
rect 3562 1762 3568 1822
rect 3628 1762 3634 1822
rect 2844 1494 3332 1500
rect 2844 1460 2856 1494
rect 3320 1460 3332 1494
rect 2844 1454 3332 1460
rect 2550 1366 2562 1410
rect 1578 834 1592 874
rect 2556 868 2562 1366
rect 1532 670 1592 834
rect 2548 834 2562 868
rect 2596 1366 2610 1410
rect 3568 1410 3628 1762
rect 4074 1500 4134 1857
rect 4578 1554 4584 1614
rect 4644 1554 4650 1614
rect 3862 1494 4350 1500
rect 3862 1460 3874 1494
rect 4338 1460 4350 1494
rect 3862 1454 4350 1460
rect 2596 868 2602 1366
rect 2596 834 2608 868
rect 1826 784 2314 790
rect 1826 750 1838 784
rect 2302 750 2314 784
rect 1826 744 2314 750
rect 2040 670 2100 744
rect 2548 670 2608 834
rect 3568 834 3580 1410
rect 3614 834 3628 1410
rect 4584 1410 4644 1554
rect 5098 1500 5158 1857
rect 5602 1828 5662 1947
rect 6629 1947 6635 2482
rect 6669 2482 6682 2523
rect 7636 2523 7696 2654
rect 7636 2488 7653 2523
rect 6669 1947 6675 2482
rect 6629 1935 6675 1947
rect 7647 1947 7653 2488
rect 7687 2488 7696 2523
rect 7687 1947 7693 2488
rect 7647 1935 7693 1947
rect 5899 1897 6387 1903
rect 5899 1863 5911 1897
rect 6375 1863 6387 1897
rect 5899 1857 6387 1863
rect 6917 1897 7405 1903
rect 6917 1863 6929 1897
rect 7393 1863 7405 1897
rect 6917 1857 7405 1863
rect 5598 1822 5662 1828
rect 5658 1762 5662 1822
rect 5598 1756 5662 1762
rect 4880 1494 5368 1500
rect 4880 1460 4892 1494
rect 5356 1460 5368 1494
rect 4880 1454 5368 1460
rect 4584 1358 4598 1410
rect 2844 784 3332 790
rect 2844 750 2856 784
rect 3320 750 3332 784
rect 2844 744 3332 750
rect 3054 670 3114 744
rect 1532 610 3054 670
rect 3114 610 3120 670
rect -1378 -576 -1266 210
rect 3568 110 3628 834
rect 4592 834 4598 1358
rect 4632 1358 4644 1410
rect 5602 1410 5662 1756
rect 6114 1500 6174 1857
rect 7748 1720 7808 3764
rect 8280 2920 8340 4900
rect 8412 3926 8472 5140
rect 8828 5060 8888 5066
rect 11902 5060 11962 7622
rect 8826 5000 8828 5006
rect 10012 5000 10018 5060
rect 10078 5000 10084 5060
rect 11206 5000 11212 5060
rect 11272 5000 11278 5060
rect 11896 5000 11902 5060
rect 11962 5000 11968 5060
rect 8826 4965 8888 5000
rect 8523 4903 8888 4965
rect 8523 4748 8585 4903
rect 8675 4838 8737 4903
rect 8642 4832 8770 4838
rect 8642 4798 8654 4832
rect 8758 4798 8770 4832
rect 8642 4792 8770 4798
rect 8826 4748 8888 4903
rect 9266 4900 9272 4960
rect 9332 4900 9338 4960
rect 9564 4900 9570 4960
rect 9630 4900 9636 4960
rect 9272 4838 9332 4900
rect 9570 4838 9630 4900
rect 8940 4832 9068 4838
rect 8940 4798 8952 4832
rect 9056 4798 9068 4832
rect 8940 4792 9068 4798
rect 9238 4832 9366 4838
rect 9238 4798 9250 4832
rect 9354 4798 9366 4832
rect 9238 4792 9366 4798
rect 9536 4832 9664 4838
rect 9536 4798 9548 4832
rect 9652 4798 9664 4832
rect 9536 4792 9664 4798
rect 9834 4832 9962 4838
rect 9834 4798 9846 4832
rect 9950 4798 9962 4832
rect 9834 4792 9962 4798
rect 8523 4715 8540 4748
rect 8534 4172 8540 4715
rect 8574 4716 8588 4748
rect 8574 4715 8585 4716
rect 8574 4172 8580 4715
rect 8826 4708 8838 4748
rect 8828 4696 8838 4708
rect 8534 4160 8580 4172
rect 8832 4172 8838 4696
rect 8872 4696 8888 4748
rect 9130 4748 9176 4760
rect 8872 4172 8878 4696
rect 9130 4221 9136 4748
rect 8832 4160 8878 4172
rect 9121 4172 9136 4221
rect 9170 4221 9176 4748
rect 9428 4748 9474 4760
rect 9428 4228 9434 4748
rect 9170 4172 9179 4221
rect 9420 4208 9434 4228
rect 8642 4122 8770 4128
rect 8642 4088 8654 4122
rect 8758 4088 8770 4122
rect 8642 4082 8770 4088
rect 8940 4122 9068 4128
rect 8940 4088 8952 4122
rect 9056 4088 9068 4122
rect 8940 4082 9068 4088
rect 8824 3926 8884 3932
rect 8402 3866 8408 3926
rect 8468 3866 8474 3926
rect 8884 3866 8886 3876
rect 8824 3836 8886 3866
rect 8528 3776 8886 3836
rect 8976 3818 9036 4082
rect 9121 4057 9179 4172
rect 9418 4172 9434 4208
rect 9468 4228 9474 4748
rect 9726 4748 9772 4760
rect 9468 4172 9480 4228
rect 9726 4186 9732 4748
rect 9720 4172 9732 4186
rect 9766 4186 9772 4748
rect 10018 4748 10078 5000
rect 10460 4900 10466 4960
rect 10526 4900 10532 4960
rect 10756 4900 10762 4960
rect 10822 4900 10828 4960
rect 10466 4838 10526 4900
rect 10762 4838 10822 4900
rect 10132 4832 10260 4838
rect 10132 4798 10144 4832
rect 10248 4798 10260 4832
rect 10132 4792 10260 4798
rect 10430 4832 10558 4838
rect 10430 4798 10442 4832
rect 10546 4798 10558 4832
rect 10430 4792 10558 4798
rect 10728 4832 10856 4838
rect 10728 4798 10740 4832
rect 10844 4798 10856 4832
rect 10728 4792 10856 4798
rect 11026 4832 11154 4838
rect 11026 4798 11038 4832
rect 11142 4798 11154 4832
rect 11026 4792 11154 4798
rect 10018 4688 10030 4748
rect 9766 4179 9780 4186
rect 9766 4172 9783 4179
rect 9238 4122 9366 4128
rect 9238 4088 9250 4122
rect 9354 4088 9366 4122
rect 9238 4082 9366 4088
rect 9115 3999 9121 4057
rect 9179 3999 9185 4057
rect 8528 3636 8588 3776
rect 8676 3726 8736 3776
rect 8642 3720 8770 3726
rect 8642 3686 8654 3720
rect 8758 3686 8770 3720
rect 8642 3680 8770 3686
rect 8528 3588 8540 3636
rect 8534 3060 8540 3588
rect 8574 3588 8588 3636
rect 8824 3636 8886 3776
rect 8970 3758 8976 3818
rect 9036 3758 9042 3818
rect 8940 3720 9068 3726
rect 8940 3686 8952 3720
rect 9056 3686 9068 3720
rect 8940 3680 9068 3686
rect 8824 3598 8838 3636
rect 8574 3060 8580 3588
rect 8826 3586 8838 3598
rect 8832 3100 8838 3586
rect 8534 3048 8580 3060
rect 8824 3060 8838 3100
rect 8872 3586 8886 3636
rect 9121 3636 9179 3999
rect 9418 3926 9478 4172
rect 9536 4122 9664 4128
rect 9536 4088 9548 4122
rect 9652 4088 9664 4122
rect 9536 4082 9664 4088
rect 9720 4057 9783 4172
rect 10024 4172 10030 4688
rect 10064 4688 10078 4748
rect 10322 4748 10368 4760
rect 10064 4172 10070 4688
rect 10322 4195 10328 4748
rect 10024 4160 10070 4172
rect 10316 4172 10328 4195
rect 10362 4195 10368 4748
rect 10620 4748 10666 4760
rect 10620 4230 10626 4748
rect 10612 4214 10626 4230
rect 10362 4172 10374 4195
rect 9834 4122 9962 4128
rect 9834 4088 9846 4122
rect 9950 4088 9962 4122
rect 9834 4082 9962 4088
rect 10132 4122 10260 4128
rect 10132 4088 10144 4122
rect 10248 4088 10260 4122
rect 10132 4082 10260 4088
rect 9719 3999 9725 4057
rect 9783 3999 9789 4057
rect 9412 3866 9418 3926
rect 9478 3866 9484 3926
rect 9268 3758 9274 3818
rect 9334 3758 9340 3818
rect 9568 3758 9574 3818
rect 9634 3758 9640 3818
rect 9274 3726 9334 3758
rect 9574 3726 9634 3758
rect 9238 3720 9366 3726
rect 9238 3686 9250 3720
rect 9354 3686 9366 3720
rect 9238 3680 9366 3686
rect 9536 3720 9664 3726
rect 9536 3686 9548 3720
rect 9652 3686 9664 3720
rect 9536 3680 9664 3686
rect 9121 3605 9136 3636
rect 8872 3100 8878 3586
rect 9130 3100 9136 3605
rect 8872 3060 8884 3100
rect 8642 3010 8770 3016
rect 8642 2976 8654 3010
rect 8758 2976 8770 3010
rect 8642 2970 8770 2976
rect 8274 2860 8280 2920
rect 8340 2860 8346 2920
rect 6612 1660 6618 1720
rect 6678 1660 6684 1720
rect 7742 1660 7748 1720
rect 7808 1660 7814 1720
rect 5898 1494 6386 1500
rect 5898 1460 5910 1494
rect 6374 1460 6386 1494
rect 5898 1454 6386 1460
rect 4632 834 4638 1358
rect 4592 822 4638 834
rect 5602 834 5616 1410
rect 5650 834 5662 1410
rect 6618 1410 6678 1660
rect 6916 1494 7404 1500
rect 6916 1460 6928 1494
rect 7392 1460 7404 1494
rect 6916 1454 7404 1460
rect 6618 1370 6634 1410
rect 6628 890 6634 1370
rect 3862 784 4350 790
rect 3862 750 3874 784
rect 4338 750 4350 784
rect 3862 744 4350 750
rect 4880 784 5368 790
rect 4880 750 4892 784
rect 5356 750 5368 784
rect 4880 744 5368 750
rect 4080 670 4140 744
rect 5104 670 5164 744
rect 4074 610 4080 670
rect 4140 610 4146 670
rect 5098 610 5104 670
rect 5164 610 5170 670
rect 5602 110 5662 834
rect 6622 834 6634 890
rect 6668 1370 6678 1410
rect 7646 1410 7692 1422
rect 6668 890 6674 1370
rect 6668 834 6682 890
rect 7646 874 7652 1410
rect 5898 784 6386 790
rect 5898 750 5910 784
rect 6374 750 6386 784
rect 5898 744 6386 750
rect 6004 670 6064 676
rect 6106 670 6166 744
rect 6622 670 6682 834
rect 7638 834 7652 874
rect 7686 874 7692 1410
rect 7686 834 7698 874
rect 6916 784 7404 790
rect 6916 750 6928 784
rect 7392 750 7404 784
rect 6916 744 7404 750
rect 7130 670 7190 744
rect 7638 670 7698 834
rect 8280 700 8340 2860
rect 8640 2608 8768 2614
rect 8640 2574 8652 2608
rect 8756 2574 8768 2608
rect 8640 2568 8768 2574
rect 8532 2524 8578 2536
rect 8532 1996 8538 2524
rect 8526 1948 8538 1996
rect 8572 1996 8578 2524
rect 8824 2524 8884 3060
rect 9122 3060 9136 3100
rect 9170 3605 9179 3636
rect 9428 3636 9474 3648
rect 9170 3100 9176 3605
rect 9428 3100 9434 3636
rect 9170 3060 9182 3100
rect 8978 3016 9026 3018
rect 8940 3010 9068 3016
rect 8940 2976 8952 3010
rect 9056 2976 9068 3010
rect 8940 2970 9068 2976
rect 8974 2920 9034 2970
rect 8968 2860 8974 2920
rect 9034 2860 9040 2920
rect 8974 2614 9034 2860
rect 8938 2608 9066 2614
rect 8938 2574 8950 2608
rect 9054 2574 9066 2608
rect 8938 2568 9066 2574
rect 8824 2486 8836 2524
rect 8572 1948 8586 1996
rect 8830 1994 8836 2486
rect 8526 1800 8586 1948
rect 8822 1948 8836 1994
rect 8870 2486 8884 2524
rect 9122 2524 9182 3060
rect 9420 3060 9434 3100
rect 9468 3100 9474 3636
rect 9720 3636 9783 3999
rect 9868 3818 9928 4082
rect 10010 3866 10016 3926
rect 10076 3866 10082 3926
rect 9862 3758 9868 3818
rect 9928 3758 9934 3818
rect 9834 3720 9962 3726
rect 9834 3686 9846 3720
rect 9950 3686 9962 3720
rect 9834 3680 9962 3686
rect 9720 3623 9732 3636
rect 9468 3060 9480 3100
rect 9726 3060 9732 3623
rect 9766 3623 9783 3636
rect 10016 3636 10076 3866
rect 10164 3818 10224 4082
rect 10316 4057 10374 4172
rect 10610 4172 10626 4214
rect 10660 4230 10666 4748
rect 10918 4748 10964 4760
rect 10660 4172 10672 4230
rect 10918 4223 10924 4748
rect 10913 4202 10924 4223
rect 10912 4172 10924 4202
rect 10958 4223 10964 4748
rect 11212 4748 11272 5000
rect 11324 4832 11452 4838
rect 11324 4798 11336 4832
rect 11440 4798 11452 4832
rect 11324 4792 11452 4798
rect 11622 4832 11750 4838
rect 11622 4798 11634 4832
rect 11738 4798 11750 4832
rect 11622 4792 11750 4798
rect 11212 4692 11222 4748
rect 10958 4202 10971 4223
rect 10958 4172 10972 4202
rect 10430 4122 10558 4128
rect 10430 4088 10442 4122
rect 10546 4088 10558 4122
rect 10430 4082 10558 4088
rect 10310 3999 10316 4057
rect 10374 3999 10380 4057
rect 10158 3758 10164 3818
rect 10224 3758 10230 3818
rect 10132 3720 10260 3726
rect 10132 3686 10144 3720
rect 10248 3686 10260 3720
rect 10132 3680 10260 3686
rect 9766 3060 9772 3623
rect 10016 3586 10030 3636
rect 10024 3060 10030 3586
rect 10064 3586 10076 3636
rect 10316 3636 10374 3999
rect 10610 3926 10670 4172
rect 10728 4122 10856 4128
rect 10728 4088 10740 4122
rect 10844 4088 10856 4122
rect 10728 4082 10856 4088
rect 10912 4057 10972 4172
rect 11216 4172 11222 4692
rect 11256 4692 11272 4748
rect 11514 4748 11560 4760
rect 11256 4172 11262 4692
rect 11514 4217 11520 4748
rect 11509 4210 11520 4217
rect 11216 4160 11262 4172
rect 11506 4172 11520 4210
rect 11554 4217 11560 4748
rect 11812 4748 11858 4760
rect 11554 4172 11567 4217
rect 11812 4212 11818 4748
rect 11026 4122 11154 4128
rect 11026 4088 11038 4122
rect 11142 4088 11154 4122
rect 11026 4082 11154 4088
rect 11324 4122 11452 4128
rect 11324 4088 11336 4122
rect 11440 4088 11452 4122
rect 11324 4082 11452 4088
rect 10912 3999 10913 4057
rect 10971 3999 10972 4057
rect 10604 3866 10610 3926
rect 10670 3866 10676 3926
rect 10458 3758 10464 3818
rect 10524 3758 10530 3818
rect 10760 3758 10766 3818
rect 10826 3758 10832 3818
rect 10464 3726 10524 3758
rect 10766 3726 10826 3758
rect 10430 3720 10558 3726
rect 10430 3686 10442 3720
rect 10546 3686 10558 3720
rect 10430 3680 10558 3686
rect 10728 3720 10856 3726
rect 10728 3686 10740 3720
rect 10844 3686 10856 3720
rect 10728 3680 10856 3686
rect 10620 3636 10666 3648
rect 10316 3607 10328 3636
rect 10064 3060 10070 3586
rect 10322 3066 10328 3607
rect 9238 3010 9366 3016
rect 9238 2976 9250 3010
rect 9354 2976 9366 3010
rect 9238 2970 9366 2976
rect 9420 2812 9480 3060
rect 9536 3010 9664 3016
rect 9536 2976 9548 3010
rect 9652 2976 9664 3010
rect 9536 2970 9664 2976
rect 9414 2752 9420 2812
rect 9480 2752 9486 2812
rect 9236 2608 9364 2614
rect 9236 2574 9248 2608
rect 9352 2574 9364 2608
rect 9236 2568 9364 2574
rect 9122 2486 9134 2524
rect 8870 1998 8876 2486
rect 9128 2002 9134 2486
rect 8870 1948 8890 1998
rect 9122 1948 9134 2002
rect 9168 2486 9182 2524
rect 9420 2524 9480 2752
rect 9534 2608 9662 2614
rect 9534 2574 9546 2608
rect 9650 2574 9662 2608
rect 9534 2568 9662 2574
rect 9720 2524 9780 3060
rect 10024 3048 10070 3060
rect 10314 3060 10328 3066
rect 10362 3608 10378 3636
rect 10362 3607 10374 3608
rect 10362 3066 10368 3607
rect 10620 3116 10626 3636
rect 10614 3102 10626 3116
rect 10362 3060 10374 3066
rect 10612 3060 10626 3102
rect 10660 3116 10666 3636
rect 10912 3636 10972 3999
rect 11056 3818 11116 4082
rect 11202 3866 11208 3926
rect 11268 3866 11274 3926
rect 11050 3758 11056 3818
rect 11116 3758 11122 3818
rect 11026 3720 11154 3726
rect 11026 3686 11038 3720
rect 11142 3686 11154 3720
rect 11026 3680 11154 3686
rect 10912 3616 10924 3636
rect 10660 3060 10674 3116
rect 10918 3060 10924 3616
rect 10958 3616 10972 3636
rect 11208 3636 11268 3866
rect 11360 3818 11420 4082
rect 11506 4057 11567 4172
rect 11804 4172 11818 4212
rect 11852 4212 11858 4748
rect 11852 4172 11864 4212
rect 11622 4122 11750 4128
rect 11622 4088 11634 4122
rect 11738 4088 11750 4122
rect 11622 4082 11750 4088
rect 11506 4048 11509 4057
rect 11508 3999 11509 4048
rect 11660 4054 11720 4082
rect 11804 4054 11864 4172
rect 11567 3999 11864 4054
rect 11508 3994 11864 3999
rect 11508 3842 11568 3994
rect 11354 3758 11360 3818
rect 11420 3758 11426 3818
rect 11508 3782 11866 3842
rect 11324 3720 11452 3726
rect 11324 3686 11336 3720
rect 11440 3686 11452 3720
rect 11324 3680 11452 3686
rect 10958 3060 10964 3616
rect 11208 3586 11222 3636
rect 11216 3060 11222 3586
rect 11256 3586 11268 3636
rect 11508 3636 11568 3782
rect 11656 3726 11716 3782
rect 11622 3720 11750 3726
rect 11622 3686 11634 3720
rect 11738 3686 11750 3720
rect 11622 3680 11750 3686
rect 11508 3604 11520 3636
rect 11256 3060 11262 3586
rect 11514 3104 11520 3604
rect 9834 3010 9962 3016
rect 9834 2976 9846 3010
rect 9950 2976 9962 3010
rect 9834 2970 9962 2976
rect 10132 3010 10260 3016
rect 10132 2976 10144 3010
rect 10248 2976 10260 3010
rect 10132 2970 10260 2976
rect 9870 2920 9930 2970
rect 10164 2920 10224 2970
rect 9864 2860 9870 2920
rect 9930 2860 9936 2920
rect 10158 2860 10164 2920
rect 10224 2860 10230 2920
rect 9874 2614 9930 2860
rect 10164 2614 10220 2860
rect 9832 2608 9960 2614
rect 9832 2574 9844 2608
rect 9948 2574 9960 2608
rect 9832 2568 9960 2574
rect 10130 2608 10258 2614
rect 10130 2574 10142 2608
rect 10246 2574 10258 2608
rect 10130 2568 10258 2574
rect 10022 2524 10068 2536
rect 10314 2530 10374 3060
rect 10430 3010 10558 3016
rect 10430 2976 10442 3010
rect 10546 2976 10558 3010
rect 10430 2970 10558 2976
rect 10614 2812 10674 3060
rect 10728 3010 10856 3016
rect 10728 2976 10740 3010
rect 10844 2976 10856 3010
rect 10728 2970 10856 2976
rect 10608 2752 10614 2812
rect 10674 2752 10680 2812
rect 10428 2608 10556 2614
rect 10428 2574 10440 2608
rect 10544 2574 10556 2608
rect 10428 2568 10556 2574
rect 9420 2486 9432 2524
rect 9168 2002 9174 2486
rect 9168 1948 9182 2002
rect 8640 1898 8768 1904
rect 8640 1864 8652 1898
rect 8756 1864 8768 1898
rect 8640 1858 8768 1864
rect 8672 1800 8732 1858
rect 8822 1800 8882 1948
rect 8938 1898 9066 1904
rect 8938 1864 8950 1898
rect 9054 1864 9066 1898
rect 8938 1858 9066 1864
rect 9122 1828 9182 1948
rect 9426 1948 9432 2486
rect 9466 2486 9480 2524
rect 9466 1948 9472 2486
rect 9724 2008 9730 2524
rect 9426 1936 9472 1948
rect 9716 1948 9730 2008
rect 9764 2008 9770 2524
rect 9764 1948 9776 2008
rect 10022 1996 10028 2524
rect 9236 1898 9364 1904
rect 9236 1864 9248 1898
rect 9352 1864 9364 1898
rect 9236 1858 9364 1864
rect 9534 1898 9662 1904
rect 9534 1864 9546 1898
rect 9650 1864 9662 1898
rect 9534 1858 9662 1864
rect 8526 1740 8882 1800
rect 9116 1768 9122 1828
rect 9182 1768 9188 1828
rect 8524 1734 8586 1740
rect 8584 1680 8586 1734
rect 8524 1668 8584 1674
rect 8966 1566 8972 1626
rect 9032 1566 9038 1626
rect 8972 1504 9032 1566
rect 8640 1498 8768 1504
rect 8640 1464 8652 1498
rect 8756 1464 8768 1498
rect 8640 1458 8768 1464
rect 8938 1498 9066 1504
rect 8938 1464 8950 1498
rect 9054 1464 9066 1498
rect 8938 1458 9066 1464
rect 8532 1414 8578 1426
rect 8532 890 8538 1414
rect 8524 838 8538 890
rect 8572 890 8578 1414
rect 8830 1414 8876 1426
rect 8572 838 8584 890
rect 8830 886 8836 1414
rect 8524 700 8584 838
rect 8824 838 8836 886
rect 8870 886 8876 1414
rect 9122 1414 9182 1768
rect 9270 1626 9330 1858
rect 9410 1674 9416 1734
rect 9476 1674 9482 1734
rect 9264 1566 9270 1626
rect 9330 1566 9336 1626
rect 9236 1498 9364 1504
rect 9236 1464 9248 1498
rect 9352 1464 9364 1498
rect 9236 1458 9364 1464
rect 9122 1370 9134 1414
rect 8870 838 8884 886
rect 8640 788 8768 794
rect 8640 754 8652 788
rect 8756 754 8768 788
rect 8640 748 8768 754
rect 8672 700 8732 748
rect 8824 700 8884 838
rect 9128 838 9134 1370
rect 9168 1370 9182 1414
rect 9416 1414 9476 1674
rect 9566 1626 9626 1858
rect 9716 1828 9776 1948
rect 10014 1948 10028 1996
rect 10062 1996 10068 2524
rect 10320 2524 10366 2530
rect 10614 2524 10674 2752
rect 10726 2608 10854 2614
rect 10726 2574 10738 2608
rect 10842 2574 10854 2608
rect 10726 2568 10854 2574
rect 10062 1990 10074 1996
rect 10062 1948 10080 1990
rect 10320 1978 10326 2524
rect 10316 1948 10326 1978
rect 10360 1978 10366 2524
rect 10612 2486 10624 2524
rect 10360 1948 10376 1978
rect 9832 1898 9960 1904
rect 9832 1864 9844 1898
rect 9948 1864 9960 1898
rect 9832 1858 9960 1864
rect 9710 1768 9716 1828
rect 9776 1768 9782 1828
rect 9560 1566 9566 1626
rect 9626 1566 9632 1626
rect 9534 1498 9662 1504
rect 9534 1464 9546 1498
rect 9650 1464 9662 1498
rect 9534 1458 9662 1464
rect 9716 1414 9776 1768
rect 10014 1734 10074 1948
rect 10130 1898 10258 1904
rect 10130 1864 10142 1898
rect 10246 1864 10258 1898
rect 10130 1858 10258 1864
rect 10316 1828 10376 1948
rect 10618 1948 10624 2486
rect 10658 2486 10674 2524
rect 10908 2524 10968 3060
rect 11216 3048 11262 3060
rect 11504 3060 11520 3104
rect 11554 3604 11568 3636
rect 11806 3636 11866 3782
rect 11554 3104 11560 3604
rect 11806 3600 11818 3636
rect 11554 3060 11564 3104
rect 11812 3100 11818 3600
rect 11806 3060 11818 3100
rect 11852 3600 11866 3636
rect 11852 3100 11858 3600
rect 11852 3060 11866 3100
rect 11026 3010 11154 3016
rect 11026 2976 11038 3010
rect 11142 2976 11154 3010
rect 11026 2970 11154 2976
rect 11324 3010 11452 3016
rect 11324 2976 11336 3010
rect 11440 2976 11452 3010
rect 11324 2970 11452 2976
rect 11058 2920 11118 2970
rect 11360 2920 11420 2970
rect 11052 2860 11058 2920
rect 11118 2860 11124 2920
rect 11354 2860 11360 2920
rect 11420 2860 11426 2920
rect 11062 2614 11118 2860
rect 11364 2614 11420 2860
rect 11024 2608 11152 2614
rect 11024 2574 11036 2608
rect 11140 2574 11152 2608
rect 11024 2568 11152 2574
rect 11322 2608 11450 2614
rect 11322 2574 11334 2608
rect 11438 2574 11450 2608
rect 11322 2568 11450 2574
rect 10908 2496 10922 2524
rect 10658 1948 10664 2486
rect 10916 2002 10922 2496
rect 10618 1936 10664 1948
rect 10910 1948 10922 2002
rect 10956 2496 10968 2524
rect 11214 2524 11260 2536
rect 10956 2002 10962 2496
rect 10956 1948 10970 2002
rect 11214 1998 11220 2524
rect 10428 1898 10556 1904
rect 10428 1864 10440 1898
rect 10544 1864 10556 1898
rect 10428 1858 10556 1864
rect 10726 1898 10854 1904
rect 10726 1864 10738 1898
rect 10842 1864 10854 1898
rect 10726 1858 10854 1864
rect 10310 1768 10316 1828
rect 10376 1768 10382 1828
rect 10008 1674 10014 1734
rect 10074 1674 10080 1734
rect 9864 1566 9870 1626
rect 9930 1566 9936 1626
rect 10160 1566 10166 1626
rect 10226 1566 10232 1626
rect 9870 1504 9930 1566
rect 10166 1504 10226 1566
rect 9832 1498 9960 1504
rect 9832 1464 9844 1498
rect 9948 1464 9960 1498
rect 9832 1458 9960 1464
rect 10130 1498 10258 1504
rect 10130 1464 10142 1498
rect 10246 1464 10258 1498
rect 10130 1458 10258 1464
rect 9416 1380 9432 1414
rect 9168 838 9174 1370
rect 9424 1356 9432 1380
rect 9128 826 9174 838
rect 9426 838 9432 1356
rect 9466 1356 9484 1414
rect 9716 1380 9730 1414
rect 9466 838 9472 1356
rect 9426 826 9472 838
rect 9724 838 9730 1380
rect 9764 1380 9776 1414
rect 10022 1414 10068 1426
rect 9764 838 9770 1380
rect 10022 878 10028 1414
rect 10014 876 10028 878
rect 9724 826 9770 838
rect 10012 838 10028 876
rect 10062 878 10068 1414
rect 10316 1414 10376 1768
rect 10464 1626 10524 1858
rect 10606 1674 10612 1734
rect 10672 1674 10678 1734
rect 10458 1566 10464 1626
rect 10524 1566 10530 1626
rect 10428 1498 10556 1504
rect 10428 1464 10440 1498
rect 10544 1464 10556 1498
rect 10428 1458 10556 1464
rect 10316 1382 10326 1414
rect 10062 838 10074 878
rect 10320 838 10326 1382
rect 10360 1382 10376 1414
rect 10612 1414 10672 1674
rect 10760 1626 10820 1858
rect 10910 1828 10970 1948
rect 11212 1948 11220 1998
rect 11254 1998 11260 2524
rect 11504 2524 11564 3060
rect 11812 3048 11858 3060
rect 11622 3010 11750 3016
rect 11622 2976 11634 3010
rect 11738 2976 11750 3010
rect 11622 2970 11750 2976
rect 11902 2812 11962 5000
rect 11620 2608 11748 2614
rect 11620 2574 11632 2608
rect 11736 2574 11748 2608
rect 11620 2568 11748 2574
rect 11810 2524 11856 2536
rect 11254 1948 11272 1998
rect 11024 1898 11152 1904
rect 11024 1864 11036 1898
rect 11140 1864 11152 1898
rect 11024 1858 11152 1864
rect 10904 1768 10910 1828
rect 10970 1768 10976 1828
rect 10754 1566 10760 1626
rect 10820 1566 10826 1626
rect 10726 1498 10854 1504
rect 10726 1464 10738 1498
rect 10842 1464 10854 1498
rect 10726 1458 10854 1464
rect 10910 1414 10970 1768
rect 11212 1734 11272 1948
rect 11504 1948 11518 2524
rect 11552 2488 11568 2524
rect 11802 2492 11816 2524
rect 11552 1948 11564 2488
rect 11810 2000 11816 2492
rect 11802 1978 11816 2000
rect 11800 1948 11816 1978
rect 11850 2492 11862 2524
rect 11850 2000 11856 2492
rect 11850 1948 11862 2000
rect 11322 1898 11450 1904
rect 11322 1864 11334 1898
rect 11438 1864 11450 1898
rect 11322 1858 11450 1864
rect 11504 1828 11564 1948
rect 11620 1898 11748 1904
rect 11620 1864 11632 1898
rect 11736 1864 11748 1898
rect 11620 1858 11748 1864
rect 11498 1768 11504 1828
rect 11564 1824 11570 1828
rect 11652 1824 11712 1858
rect 11802 1824 11862 1948
rect 11564 1768 11862 1824
rect 11504 1764 11862 1768
rect 11206 1674 11212 1734
rect 11272 1674 11278 1734
rect 11050 1566 11056 1626
rect 11116 1566 11122 1626
rect 11354 1566 11360 1626
rect 11420 1566 11426 1626
rect 11504 1602 11564 1764
rect 11056 1504 11116 1566
rect 11360 1504 11420 1566
rect 11504 1542 11864 1602
rect 11024 1498 11152 1504
rect 11024 1464 11036 1498
rect 11140 1464 11152 1498
rect 11024 1458 11152 1464
rect 11322 1498 11450 1504
rect 11322 1464 11334 1498
rect 11438 1464 11450 1498
rect 11322 1458 11450 1464
rect 10360 838 10366 1382
rect 10612 1376 10624 1414
rect 10616 1354 10624 1376
rect 8938 788 9066 794
rect 8938 754 8950 788
rect 9054 754 9066 788
rect 8938 748 9066 754
rect 9236 788 9364 794
rect 9236 754 9248 788
rect 9352 754 9364 788
rect 9236 748 9364 754
rect 9534 788 9662 794
rect 9534 754 9546 788
rect 9650 754 9662 788
rect 9534 748 9662 754
rect 9832 788 9960 794
rect 9832 754 9844 788
rect 9948 754 9960 788
rect 9832 748 9960 754
rect 9270 700 9330 748
rect 9568 700 9628 748
rect 6064 610 7698 670
rect 8274 640 8280 700
rect 8340 640 8346 700
rect 8524 640 8884 700
rect 9264 640 9270 700
rect 9330 640 9336 700
rect 9562 640 9568 700
rect 9628 640 9634 700
rect 6004 604 6064 610
rect 8824 600 8884 640
rect 10012 600 10072 838
rect 10320 826 10366 838
rect 10618 838 10624 1354
rect 10658 1354 10676 1414
rect 10910 1388 10922 1414
rect 10658 838 10664 1354
rect 10618 826 10664 838
rect 10916 838 10922 1388
rect 10956 1388 10970 1414
rect 11214 1414 11260 1426
rect 10956 838 10962 1388
rect 11214 886 11220 1414
rect 11206 838 11220 886
rect 11254 886 11260 1414
rect 11504 1414 11564 1542
rect 11654 1504 11714 1542
rect 11620 1498 11748 1504
rect 11620 1464 11632 1498
rect 11736 1464 11748 1498
rect 11620 1458 11748 1464
rect 11504 1358 11518 1414
rect 11254 874 11266 886
rect 11254 838 11268 874
rect 10916 826 10962 838
rect 10130 788 10258 794
rect 10130 754 10142 788
rect 10246 754 10258 788
rect 10130 748 10258 754
rect 10428 788 10556 794
rect 10428 754 10440 788
rect 10544 754 10556 788
rect 10428 748 10556 754
rect 10726 788 10854 794
rect 10726 754 10738 788
rect 10842 754 10854 788
rect 10726 748 10854 754
rect 11024 788 11152 794
rect 11024 754 11036 788
rect 11140 754 11152 788
rect 11024 748 11152 754
rect 10464 700 10524 748
rect 10766 700 10826 748
rect 10458 640 10464 700
rect 10524 640 10530 700
rect 10760 640 10766 700
rect 10826 640 10832 700
rect 11208 600 11268 838
rect 11512 838 11518 1358
rect 11552 1358 11564 1414
rect 11804 1414 11864 1542
rect 11804 1388 11816 1414
rect 11552 838 11558 1358
rect 11512 826 11558 838
rect 11810 838 11816 1388
rect 11850 1388 11864 1414
rect 11850 838 11856 1388
rect 11810 826 11856 838
rect 11322 788 11450 794
rect 11322 754 11334 788
rect 11438 754 11450 788
rect 11322 748 11450 754
rect 11620 788 11748 794
rect 11620 754 11632 788
rect 11736 754 11748 788
rect 11620 748 11748 754
rect 11902 600 11962 2752
rect 12026 3818 12086 3824
rect 12026 1626 12086 3758
rect 12926 2996 12986 12480
rect 12920 2936 12926 2996
rect 12986 2936 12992 2996
rect 13060 2778 13120 12686
rect 13286 11424 13346 15124
rect 14020 14946 33432 15006
rect 14020 14900 14080 14946
rect 13814 14894 14302 14900
rect 13814 14860 13826 14894
rect 14290 14860 14302 14894
rect 13814 14854 14302 14860
rect 13526 14810 13572 14822
rect 13526 14268 13532 14810
rect 13518 14234 13532 14268
rect 13566 14268 13572 14810
rect 14536 14810 14596 14946
rect 15048 14900 15108 14946
rect 16056 14900 16116 14946
rect 14832 14894 15320 14900
rect 14832 14860 14844 14894
rect 15308 14860 15320 14894
rect 14832 14854 15320 14860
rect 15850 14894 16338 14900
rect 15850 14860 15862 14894
rect 16326 14860 16338 14894
rect 15850 14854 16338 14860
rect 13566 14234 13578 14268
rect 13518 14092 13578 14234
rect 14536 14234 14550 14810
rect 14584 14234 14596 14810
rect 15562 14810 15608 14822
rect 15562 14272 15568 14810
rect 13814 14184 14302 14190
rect 13814 14150 13826 14184
rect 14290 14150 14302 14184
rect 13814 14144 14302 14150
rect 13512 14032 13518 14092
rect 13578 14032 13584 14092
rect 13518 13576 13578 14032
rect 14026 13666 14086 14144
rect 14536 13994 14596 14234
rect 15554 14234 15568 14272
rect 15602 14272 15608 14810
rect 16574 14810 16634 14946
rect 17066 14900 17126 14946
rect 18078 14900 18138 14946
rect 16868 14894 17356 14900
rect 16868 14860 16880 14894
rect 17344 14860 17356 14894
rect 16868 14854 17356 14860
rect 17886 14894 18374 14900
rect 17886 14860 17898 14894
rect 18362 14860 18374 14894
rect 17886 14854 18374 14860
rect 15602 14234 15614 14272
rect 14832 14184 15320 14190
rect 14832 14150 14844 14184
rect 15308 14150 15320 14184
rect 14832 14144 15320 14150
rect 14530 13934 14536 13994
rect 14596 13934 14602 13994
rect 13814 13660 14302 13666
rect 13814 13626 13826 13660
rect 14290 13626 14302 13660
rect 13814 13620 14302 13626
rect 13518 13542 13532 13576
rect 13526 13000 13532 13542
rect 13566 13542 13578 13576
rect 14536 13576 14596 13934
rect 15028 13666 15088 14144
rect 15554 14092 15614 14234
rect 16574 14234 16586 14810
rect 16620 14234 16634 14810
rect 17598 14810 17644 14822
rect 17598 14264 17604 14810
rect 16050 14190 16110 14192
rect 15850 14184 16338 14190
rect 15850 14150 15862 14184
rect 16326 14150 16338 14184
rect 15850 14144 16338 14150
rect 15548 14032 15554 14092
rect 15614 14032 15620 14092
rect 14832 13660 15320 13666
rect 14832 13626 14844 13660
rect 15308 13626 15320 13660
rect 14832 13620 15320 13626
rect 13566 13000 13572 13542
rect 14536 13528 14550 13576
rect 13526 12988 13572 13000
rect 14544 13000 14550 13528
rect 14584 13528 14596 13576
rect 15554 13576 15614 14032
rect 16050 13666 16110 14144
rect 16574 13994 16634 14234
rect 17588 14234 17604 14264
rect 17638 14264 17644 14810
rect 18608 14810 18668 14946
rect 19126 14900 19186 14946
rect 20114 14900 20174 14946
rect 18904 14894 19392 14900
rect 18904 14860 18916 14894
rect 19380 14860 19392 14894
rect 18904 14854 19392 14860
rect 19922 14894 20410 14900
rect 19922 14860 19934 14894
rect 20398 14860 20410 14894
rect 19922 14854 20410 14860
rect 17638 14234 17648 14264
rect 16868 14184 17356 14190
rect 16868 14150 16880 14184
rect 17344 14150 17356 14184
rect 16868 14144 17356 14150
rect 17588 14092 17648 14234
rect 18608 14234 18622 14810
rect 18656 14234 18668 14810
rect 19634 14810 19680 14822
rect 19634 14278 19640 14810
rect 17886 14184 18374 14190
rect 17886 14150 17898 14184
rect 18362 14150 18374 14184
rect 17886 14144 18374 14150
rect 17582 14032 17588 14092
rect 17648 14032 17654 14092
rect 18608 13994 18668 14234
rect 19628 14234 19640 14278
rect 19674 14278 19680 14810
rect 20642 14810 20702 14946
rect 21158 14900 21218 14946
rect 22160 14900 22220 14946
rect 20940 14894 21428 14900
rect 20940 14860 20952 14894
rect 21416 14860 21428 14894
rect 20940 14854 21428 14860
rect 21958 14894 22446 14900
rect 21958 14860 21970 14894
rect 22434 14860 22446 14894
rect 21958 14854 22446 14860
rect 19674 14234 19688 14278
rect 18904 14184 19392 14190
rect 18904 14150 18916 14184
rect 19380 14150 19392 14184
rect 18904 14144 19392 14150
rect 19628 14092 19688 14234
rect 20642 14234 20658 14810
rect 20692 14234 20702 14810
rect 21670 14810 21716 14822
rect 21670 14274 21676 14810
rect 19922 14184 20410 14190
rect 19922 14150 19934 14184
rect 20398 14150 20410 14184
rect 19922 14144 20410 14150
rect 19622 14032 19628 14092
rect 19688 14032 19694 14092
rect 20642 13994 20702 14234
rect 21664 14234 21676 14274
rect 21710 14274 21716 14810
rect 22682 14810 22742 14946
rect 23188 14900 23248 14946
rect 24206 14900 24266 14946
rect 22976 14894 23464 14900
rect 22976 14860 22988 14894
rect 23452 14860 23464 14894
rect 22976 14854 23464 14860
rect 23994 14894 24482 14900
rect 23994 14860 24006 14894
rect 24470 14860 24482 14894
rect 23994 14854 24482 14860
rect 23188 14852 23248 14854
rect 21710 14234 21724 14274
rect 20940 14184 21428 14190
rect 20940 14150 20952 14184
rect 21416 14150 21428 14184
rect 20940 14144 21428 14150
rect 21664 14092 21724 14234
rect 22682 14234 22694 14810
rect 22728 14234 22742 14810
rect 23706 14810 23752 14822
rect 23706 14274 23712 14810
rect 21958 14184 22446 14190
rect 21958 14150 21970 14184
rect 22434 14150 22446 14184
rect 21958 14144 22446 14150
rect 21658 14032 21664 14092
rect 21724 14032 21730 14092
rect 22682 13994 22742 14234
rect 23698 14234 23712 14274
rect 23746 14274 23752 14810
rect 24716 14810 24776 14946
rect 25224 14900 25284 14946
rect 26244 14900 26304 14946
rect 25012 14894 25500 14900
rect 25012 14860 25024 14894
rect 25488 14860 25500 14894
rect 25012 14854 25500 14860
rect 26030 14894 26518 14900
rect 26030 14860 26042 14894
rect 26506 14860 26518 14894
rect 26030 14854 26518 14860
rect 23746 14234 23758 14274
rect 22976 14184 23464 14190
rect 22976 14150 22988 14184
rect 23452 14150 23464 14184
rect 22976 14144 23464 14150
rect 23698 14092 23758 14234
rect 24716 14234 24730 14810
rect 24764 14234 24776 14810
rect 25742 14810 25788 14822
rect 25742 14280 25748 14810
rect 23994 14184 24482 14190
rect 23994 14150 24006 14184
rect 24470 14150 24482 14184
rect 23994 14144 24482 14150
rect 23692 14032 23698 14092
rect 23758 14032 23764 14092
rect 24716 13994 24776 14234
rect 25734 14234 25748 14280
rect 25782 14280 25788 14810
rect 26754 14810 26814 14946
rect 27252 14900 27312 14946
rect 28280 14900 28340 14946
rect 27048 14894 27536 14900
rect 27048 14860 27060 14894
rect 27524 14860 27536 14894
rect 27048 14854 27536 14860
rect 28066 14894 28554 14900
rect 28066 14860 28078 14894
rect 28542 14860 28554 14894
rect 28066 14854 28554 14860
rect 25782 14234 25794 14280
rect 25012 14184 25500 14190
rect 25012 14150 25024 14184
rect 25488 14150 25500 14184
rect 25012 14144 25500 14150
rect 25734 14092 25794 14234
rect 26754 14234 26766 14810
rect 26800 14234 26814 14810
rect 27778 14810 27824 14822
rect 27778 14282 27784 14810
rect 26030 14184 26518 14190
rect 26030 14150 26042 14184
rect 26506 14150 26518 14184
rect 26030 14144 26518 14150
rect 25728 14032 25734 14092
rect 25794 14032 25800 14092
rect 26754 13994 26814 14234
rect 27770 14234 27784 14282
rect 27818 14282 27824 14810
rect 28786 14810 28846 14946
rect 29282 14900 29342 14946
rect 30312 14900 30372 14946
rect 29084 14894 29572 14900
rect 29084 14860 29096 14894
rect 29560 14860 29572 14894
rect 29084 14854 29572 14860
rect 30102 14894 30590 14900
rect 30102 14860 30114 14894
rect 30578 14860 30590 14894
rect 30102 14854 30590 14860
rect 27818 14234 27830 14282
rect 27048 14184 27536 14190
rect 27048 14150 27060 14184
rect 27524 14150 27536 14184
rect 27048 14144 27536 14150
rect 27770 14092 27830 14234
rect 28786 14234 28802 14810
rect 28836 14234 28846 14810
rect 29814 14810 29860 14822
rect 29814 14288 29820 14810
rect 28066 14184 28554 14190
rect 28066 14150 28078 14184
rect 28542 14150 28554 14184
rect 28066 14144 28554 14150
rect 27764 14032 27770 14092
rect 27830 14032 27836 14092
rect 28786 13994 28846 14234
rect 29806 14234 29820 14288
rect 29854 14288 29860 14810
rect 30824 14810 30884 14946
rect 31360 14900 31420 14946
rect 32334 14900 32394 14946
rect 31120 14894 31608 14900
rect 31120 14860 31132 14894
rect 31596 14860 31608 14894
rect 31120 14854 31608 14860
rect 32138 14894 32626 14900
rect 32138 14860 32150 14894
rect 32614 14860 32626 14894
rect 32138 14854 32626 14860
rect 29854 14234 29866 14288
rect 29084 14184 29572 14190
rect 29084 14150 29096 14184
rect 29560 14150 29572 14184
rect 29084 14144 29572 14150
rect 29806 14092 29866 14234
rect 30824 14234 30838 14810
rect 30872 14234 30884 14810
rect 31850 14810 31896 14822
rect 31850 14280 31856 14810
rect 30102 14184 30590 14190
rect 30102 14150 30114 14184
rect 30578 14150 30590 14184
rect 30102 14144 30590 14150
rect 29800 14032 29806 14092
rect 29866 14032 29872 14092
rect 30824 13994 30884 14234
rect 31844 14234 31856 14280
rect 31890 14280 31896 14810
rect 32862 14810 32922 14946
rect 33372 14900 33432 14946
rect 33156 14894 33644 14900
rect 33156 14860 33168 14894
rect 33632 14860 33644 14894
rect 33156 14854 33644 14860
rect 31890 14234 31904 14280
rect 31120 14184 31608 14190
rect 31120 14150 31132 14184
rect 31596 14150 31608 14184
rect 31120 14144 31608 14150
rect 16568 13934 16574 13994
rect 16634 13934 16640 13994
rect 18602 13934 18608 13994
rect 18668 13934 18674 13994
rect 20636 13934 20642 13994
rect 20702 13934 20708 13994
rect 22676 13934 22682 13994
rect 22742 13934 22748 13994
rect 24710 13934 24716 13994
rect 24776 13934 24782 13994
rect 26748 13934 26754 13994
rect 26814 13934 26820 13994
rect 28780 13934 28786 13994
rect 28846 13934 28852 13994
rect 30818 13934 30824 13994
rect 30884 13934 30890 13994
rect 23168 13880 23228 13888
rect 23168 13820 25276 13880
rect 20140 13702 21210 13762
rect 22676 13722 22682 13782
rect 22742 13722 22748 13782
rect 20140 13666 20200 13702
rect 15850 13660 16338 13666
rect 15850 13626 15862 13660
rect 16326 13626 16338 13660
rect 15850 13620 16338 13626
rect 16868 13660 17356 13666
rect 16868 13626 16880 13660
rect 17344 13626 17356 13660
rect 16868 13620 17356 13626
rect 17886 13660 18374 13666
rect 17886 13626 17898 13660
rect 18362 13626 18374 13660
rect 17886 13620 18374 13626
rect 18904 13660 19392 13666
rect 18904 13626 18916 13660
rect 19380 13626 19392 13660
rect 18904 13620 19392 13626
rect 19922 13660 20410 13666
rect 19922 13626 19934 13660
rect 20398 13626 20410 13660
rect 19922 13620 20410 13626
rect 15554 13544 15568 13576
rect 14584 13000 14590 13528
rect 14544 12988 14590 13000
rect 15562 13000 15568 13544
rect 15602 13544 15614 13576
rect 16580 13576 16626 13588
rect 15602 13000 15608 13544
rect 16580 13028 16586 13576
rect 15562 12988 15608 13000
rect 16574 13000 16586 13028
rect 16620 13028 16626 13576
rect 17598 13576 17644 13588
rect 18616 13576 18662 13588
rect 19634 13576 19680 13588
rect 17598 13048 17604 13576
rect 16620 13000 16634 13028
rect 13814 12950 14302 12956
rect 13814 12916 13826 12950
rect 14290 12916 14302 12950
rect 13814 12910 14302 12916
rect 14832 12950 15320 12956
rect 14832 12916 14844 12950
rect 15308 12916 15320 12950
rect 14832 12910 15320 12916
rect 15850 12950 16338 12956
rect 15850 12916 15862 12950
rect 16326 12916 16338 12950
rect 15850 12910 16338 12916
rect 16574 12858 16634 13000
rect 17592 13000 17604 13048
rect 17638 13048 17644 13576
rect 18606 13542 18622 13576
rect 18616 13076 18622 13542
rect 17638 13000 17652 13048
rect 16868 12950 17356 12956
rect 16868 12916 16880 12950
rect 17344 12916 17356 12950
rect 16868 12910 17356 12916
rect 17222 12862 17282 12910
rect 17592 12862 17652 13000
rect 18606 13000 18622 13076
rect 18656 13542 18666 13576
rect 18656 13076 18662 13542
rect 18656 13060 18666 13076
rect 18656 13000 18670 13060
rect 19634 13056 19640 13576
rect 19626 13000 19640 13056
rect 19674 13056 19680 13576
rect 20646 13576 20706 13702
rect 21150 13666 21210 13702
rect 20940 13660 21428 13666
rect 20940 13626 20952 13660
rect 21416 13626 21428 13660
rect 20940 13620 21428 13626
rect 21958 13660 22446 13666
rect 21958 13626 21970 13660
rect 22434 13626 22446 13660
rect 21958 13620 22446 13626
rect 20646 13526 20658 13576
rect 19674 13000 19686 13056
rect 20652 13050 20658 13526
rect 20646 13036 20658 13050
rect 17886 12950 18374 12956
rect 17886 12916 17898 12950
rect 18362 12916 18374 12950
rect 17886 12910 18374 12916
rect 18094 12862 18154 12910
rect 18606 12862 18666 13000
rect 18904 12950 19392 12956
rect 18904 12916 18916 12950
rect 19380 12916 19392 12950
rect 18904 12910 19392 12916
rect 19134 12862 19194 12910
rect 19626 12862 19686 13000
rect 20644 13000 20658 13036
rect 20692 13526 20706 13576
rect 21670 13576 21716 13588
rect 20692 13050 20698 13526
rect 21670 13076 21676 13576
rect 20692 13000 20706 13050
rect 21658 13000 21676 13076
rect 21710 13076 21716 13576
rect 22682 13576 22742 13722
rect 23168 13666 23228 13820
rect 24202 13666 24262 13820
rect 24708 13722 24714 13782
rect 24774 13722 24780 13782
rect 22976 13660 23464 13666
rect 22976 13626 22988 13660
rect 23452 13626 23464 13660
rect 22976 13620 23464 13626
rect 23994 13660 24482 13666
rect 23994 13626 24006 13660
rect 24470 13626 24482 13660
rect 23994 13620 24482 13626
rect 22682 13542 22694 13576
rect 21710 13000 21718 13076
rect 22688 13062 22694 13542
rect 22682 13058 22694 13062
rect 19922 12950 20410 12956
rect 19922 12916 19934 12950
rect 20398 12916 20410 12950
rect 19922 12910 20410 12916
rect 16574 12798 17146 12858
rect 17216 12802 17222 12862
rect 17282 12802 17288 12862
rect 17586 12802 17592 12862
rect 17652 12802 17658 12862
rect 18088 12802 18094 12862
rect 18154 12802 18160 12862
rect 18600 12802 18606 12862
rect 18666 12802 18672 12862
rect 19128 12802 19134 12862
rect 19194 12802 19200 12862
rect 19620 12802 19626 12862
rect 19686 12802 19692 12862
rect 15040 12692 15046 12752
rect 15106 12692 15112 12752
rect 16062 12692 16068 12752
rect 16128 12692 16134 12752
rect 13516 12480 13522 12540
rect 13582 12480 13588 12540
rect 14014 12480 14020 12540
rect 14080 12480 14086 12540
rect 14526 12480 14532 12540
rect 14592 12480 14598 12540
rect 13522 12344 13582 12480
rect 14020 12434 14080 12480
rect 13814 12428 14302 12434
rect 13814 12394 13826 12428
rect 14290 12394 14302 12428
rect 13814 12388 14302 12394
rect 13522 12304 13532 12344
rect 13526 11768 13532 12304
rect 13566 12304 13582 12344
rect 14532 12344 14592 12480
rect 15046 12434 15106 12692
rect 16068 12434 16128 12692
rect 17086 12654 17146 12798
rect 17086 12648 17148 12654
rect 17086 12588 17088 12648
rect 17086 12582 17148 12588
rect 16568 12480 16574 12540
rect 16634 12480 16640 12540
rect 14832 12428 15320 12434
rect 14832 12394 14844 12428
rect 15308 12394 15320 12428
rect 14832 12388 15320 12394
rect 15850 12428 16338 12434
rect 15850 12394 15862 12428
rect 16326 12394 16338 12428
rect 15850 12388 16338 12394
rect 13566 11768 13572 12304
rect 14532 12298 14550 12344
rect 13526 11756 13572 11768
rect 14544 11768 14550 12298
rect 14584 12298 14592 12344
rect 15562 12344 15608 12356
rect 14584 11768 14590 12298
rect 15562 11826 15568 12344
rect 14544 11756 14590 11768
rect 15548 11768 15568 11826
rect 15602 11768 15608 12344
rect 16574 12344 16634 12480
rect 17086 12434 17146 12582
rect 16868 12428 17356 12434
rect 16868 12394 16880 12428
rect 17344 12394 17356 12428
rect 16868 12388 17356 12394
rect 16574 12292 16586 12344
rect 13814 11718 14302 11724
rect 13814 11684 13826 11718
rect 14290 11684 14302 11718
rect 13814 11678 14302 11684
rect 14832 11718 15320 11724
rect 14832 11684 14844 11718
rect 15308 11684 15320 11718
rect 14832 11678 15320 11684
rect 15030 11578 15036 11638
rect 15096 11578 15102 11638
rect 13280 11364 13286 11424
rect 13346 11364 13352 11424
rect 13286 10182 13346 11364
rect 13518 11268 14596 11328
rect 13518 11110 13578 11268
rect 14026 11200 14086 11268
rect 13812 11194 14300 11200
rect 13812 11160 13824 11194
rect 14288 11160 14300 11194
rect 13812 11154 14300 11160
rect 13518 11084 13530 11110
rect 13524 10534 13530 11084
rect 13564 11084 13578 11110
rect 14536 11110 14596 11268
rect 15036 11200 15096 11578
rect 15548 11546 15608 11768
rect 16580 11768 16586 12292
rect 16620 12292 16634 12344
rect 17592 12344 17652 12802
rect 18082 12588 18088 12648
rect 18148 12588 18154 12648
rect 19102 12588 19108 12648
rect 19168 12588 19174 12648
rect 18088 12434 18148 12588
rect 18602 12480 18608 12540
rect 18668 12480 18674 12540
rect 17886 12428 18374 12434
rect 17886 12394 17898 12428
rect 18362 12394 18374 12428
rect 17886 12388 18374 12394
rect 16620 11768 16626 12292
rect 17592 12280 17604 12344
rect 17598 11832 17604 12280
rect 16580 11756 16626 11768
rect 17584 11768 17604 11832
rect 17638 12280 17652 12344
rect 18608 12344 18668 12480
rect 19108 12434 19168 12588
rect 18904 12428 19392 12434
rect 18904 12394 18916 12428
rect 19380 12394 19392 12428
rect 18904 12388 19392 12394
rect 18608 12310 18622 12344
rect 17638 11768 17644 12280
rect 15850 11718 16338 11724
rect 15850 11684 15862 11718
rect 16326 11684 16338 11718
rect 15850 11678 16338 11684
rect 16868 11718 17356 11724
rect 16868 11684 16880 11718
rect 17344 11684 17356 11718
rect 16868 11678 17356 11684
rect 17072 11650 17132 11678
rect 16046 11590 16052 11650
rect 16112 11590 16118 11650
rect 17066 11590 17072 11650
rect 17132 11590 17138 11650
rect 15542 11486 15548 11546
rect 15608 11486 15614 11546
rect 15548 11252 15554 11312
rect 15614 11252 15620 11312
rect 14830 11194 15318 11200
rect 14830 11160 14842 11194
rect 15306 11160 15318 11194
rect 14830 11154 15318 11160
rect 13564 10534 13570 11084
rect 14536 11078 14548 11110
rect 14542 10578 14548 11078
rect 13524 10522 13570 10534
rect 14536 10534 14548 10578
rect 14582 11078 14596 11110
rect 15554 11110 15614 11252
rect 16052 11200 16112 11590
rect 16566 11486 16572 11546
rect 16632 11486 16638 11546
rect 15848 11194 16336 11200
rect 15848 11160 15860 11194
rect 16324 11160 16336 11194
rect 15848 11154 16336 11160
rect 15554 11084 15566 11110
rect 14582 10578 14588 11078
rect 14582 10534 14596 10578
rect 13812 10484 14300 10490
rect 13812 10450 13824 10484
rect 14288 10450 14300 10484
rect 13812 10444 14300 10450
rect 14536 10382 14596 10534
rect 15560 10534 15566 11084
rect 15600 11084 15614 11110
rect 16572 11110 16632 11486
rect 17072 11200 17132 11590
rect 17584 11546 17644 11768
rect 18616 11768 18622 12310
rect 18656 12310 18668 12344
rect 19626 12344 19686 12802
rect 20140 12752 20200 12910
rect 20644 12752 20704 13000
rect 20940 12950 21428 12956
rect 20940 12916 20952 12950
rect 21416 12916 21428 12950
rect 20940 12910 21428 12916
rect 21160 12752 21220 12910
rect 21658 12862 21718 13000
rect 22680 13000 22694 13058
rect 22728 13542 22742 13576
rect 23706 13576 23752 13588
rect 22728 13062 22734 13542
rect 23706 13066 23712 13576
rect 22728 13000 22742 13062
rect 23694 13000 23712 13066
rect 23746 13066 23752 13576
rect 24714 13576 24774 13722
rect 25216 13666 25276 13820
rect 26240 13732 27322 13792
rect 26240 13666 26300 13732
rect 25012 13660 25500 13666
rect 25012 13626 25024 13660
rect 25488 13626 25500 13660
rect 25012 13620 25500 13626
rect 26030 13660 26518 13666
rect 26030 13626 26042 13660
rect 26506 13626 26518 13660
rect 26030 13620 26518 13626
rect 24714 13542 24730 13576
rect 23746 13000 23754 13066
rect 24724 13026 24730 13542
rect 21958 12950 22446 12956
rect 21958 12916 21970 12950
rect 22434 12916 22446 12950
rect 21958 12910 22446 12916
rect 21652 12802 21658 12862
rect 21718 12802 21724 12862
rect 20134 12692 20140 12752
rect 20200 12692 20206 12752
rect 20638 12692 20644 12752
rect 20704 12692 20710 12752
rect 21154 12692 21160 12752
rect 21220 12692 21226 12752
rect 20140 12434 20200 12692
rect 20636 12480 20642 12540
rect 20702 12480 20708 12540
rect 19922 12428 20410 12434
rect 19922 12394 19934 12428
rect 20398 12394 20410 12428
rect 19922 12388 20410 12394
rect 18656 11768 18662 12310
rect 19626 12302 19640 12344
rect 19634 11810 19640 12302
rect 18616 11756 18662 11768
rect 19626 11768 19640 11810
rect 19674 12302 19686 12344
rect 20642 12344 20702 12480
rect 21160 12434 21220 12692
rect 20940 12428 21428 12434
rect 20940 12394 20952 12428
rect 21416 12394 21428 12428
rect 20940 12388 21428 12394
rect 19674 11810 19680 12302
rect 20642 12282 20658 12344
rect 19674 11768 19686 11810
rect 17886 11718 18374 11724
rect 17886 11684 17898 11718
rect 18362 11684 18374 11718
rect 17886 11678 18374 11684
rect 18904 11718 19392 11724
rect 18904 11684 18916 11718
rect 19380 11684 19392 11718
rect 18904 11678 19392 11684
rect 18084 11650 18144 11678
rect 19110 11650 19170 11678
rect 18078 11590 18084 11650
rect 18144 11590 18150 11650
rect 19104 11590 19110 11650
rect 19170 11590 19176 11650
rect 17578 11486 17584 11546
rect 17644 11486 17650 11546
rect 17584 11252 17590 11312
rect 17650 11252 17656 11312
rect 16866 11194 17354 11200
rect 16866 11160 16878 11194
rect 17342 11160 17354 11194
rect 16866 11154 17354 11160
rect 15600 10534 15606 11084
rect 16572 11078 16584 11110
rect 16578 10574 16584 11078
rect 15560 10522 15606 10534
rect 16570 10534 16584 10574
rect 16618 11078 16632 11110
rect 17590 11110 17650 11252
rect 18084 11200 18144 11590
rect 18598 11486 18604 11546
rect 18664 11486 18670 11546
rect 17884 11194 18372 11200
rect 17884 11160 17896 11194
rect 18360 11160 18372 11194
rect 17884 11154 18372 11160
rect 17590 11080 17602 11110
rect 16618 10574 16624 11078
rect 16618 10534 16630 10574
rect 14830 10484 15318 10490
rect 14830 10450 14842 10484
rect 15306 10450 15318 10484
rect 14830 10444 15318 10450
rect 15848 10484 16336 10490
rect 15848 10450 15860 10484
rect 16324 10450 16336 10484
rect 15848 10444 16336 10450
rect 13392 10322 13398 10382
rect 13458 10322 13464 10382
rect 14530 10322 14536 10382
rect 14596 10322 14602 10382
rect 13280 10122 13286 10182
rect 13346 10122 13352 10182
rect 13174 10020 13180 10080
rect 13240 10020 13246 10080
rect 13180 6590 13240 10020
rect 13286 8946 13346 10122
rect 13280 8886 13286 8946
rect 13346 8886 13352 8946
rect 13174 6530 13180 6590
rect 13240 6530 13246 6590
rect 13180 5286 13240 6530
rect 13286 6344 13346 8886
rect 13398 7608 13458 10322
rect 14528 10122 14534 10182
rect 14594 10122 14600 10182
rect 14534 10078 14594 10122
rect 13518 10018 14594 10078
rect 13518 10016 14082 10018
rect 13518 9876 13578 10016
rect 14022 9966 14082 10016
rect 13812 9960 14300 9966
rect 13812 9926 13824 9960
rect 14288 9926 14300 9960
rect 13812 9920 14300 9926
rect 13518 9844 13530 9876
rect 13524 9300 13530 9844
rect 13564 9844 13578 9876
rect 14534 9876 14594 10018
rect 15038 9966 15098 10444
rect 15546 10242 15552 10302
rect 15612 10242 15618 10302
rect 14830 9960 15318 9966
rect 14830 9926 14842 9960
rect 15306 9926 15318 9960
rect 14830 9920 15318 9926
rect 13564 9300 13570 9844
rect 14534 9840 14548 9876
rect 13524 9288 13570 9300
rect 14542 9300 14548 9840
rect 14582 9840 14594 9876
rect 15552 9876 15612 10242
rect 16066 10188 16126 10444
rect 16570 10406 16630 10534
rect 17596 10534 17602 11080
rect 17636 11080 17650 11110
rect 18604 11110 18664 11486
rect 19110 11200 19170 11590
rect 19626 11546 19686 11768
rect 20652 11768 20658 12282
rect 20692 12282 20702 12344
rect 21658 12344 21718 12802
rect 22180 12752 22240 12910
rect 22680 12864 22740 13000
rect 22976 12950 23464 12956
rect 22976 12916 22988 12950
rect 23452 12916 23464 12950
rect 22976 12910 23464 12916
rect 22680 12804 22858 12864
rect 22174 12692 22180 12752
rect 22240 12692 22246 12752
rect 22676 12692 22682 12752
rect 22742 12692 22748 12752
rect 22180 12434 22240 12692
rect 21958 12428 22446 12434
rect 21958 12394 21970 12428
rect 22434 12394 22446 12428
rect 21958 12388 22446 12394
rect 22682 12344 22742 12692
rect 22798 12540 22858 12804
rect 23176 12692 23182 12752
rect 23242 12692 23248 12752
rect 22798 12474 22858 12480
rect 23182 12434 23242 12692
rect 23322 12648 23382 12910
rect 23694 12862 23754 13000
rect 24716 13000 24730 13026
rect 24764 13542 24774 13576
rect 25742 13576 25788 13588
rect 24764 13026 24770 13542
rect 25742 13060 25748 13576
rect 24764 13000 24776 13026
rect 23994 12950 24482 12956
rect 23994 12916 24006 12950
rect 24470 12916 24482 12950
rect 23994 12910 24482 12916
rect 23688 12802 23694 12862
rect 23754 12802 23760 12862
rect 23316 12588 23322 12648
rect 23382 12588 23388 12648
rect 22976 12428 23464 12434
rect 22976 12394 22988 12428
rect 23452 12394 23464 12428
rect 22976 12388 23464 12394
rect 21658 12288 21676 12344
rect 20692 11768 20698 12282
rect 21670 11810 21676 12288
rect 20652 11756 20698 11768
rect 21662 11768 21676 11810
rect 21710 12288 21718 12344
rect 22678 12292 22694 12344
rect 21710 11810 21716 12288
rect 22688 11816 22694 12292
rect 21710 11768 21722 11810
rect 19922 11718 20410 11724
rect 19922 11684 19934 11718
rect 20398 11684 20410 11718
rect 19922 11678 20410 11684
rect 20940 11718 21428 11724
rect 20940 11684 20952 11718
rect 21416 11684 21428 11718
rect 20940 11678 21428 11684
rect 21662 11546 21722 11768
rect 22680 11768 22694 11816
rect 22728 12300 22742 12344
rect 23694 12344 23754 12802
rect 24202 12692 24208 12752
rect 24268 12692 24274 12752
rect 24208 12434 24268 12692
rect 24330 12648 24390 12910
rect 24716 12864 24776 13000
rect 25730 13000 25748 13060
rect 25782 13060 25788 13576
rect 26752 13576 26812 13732
rect 27262 13666 27322 13732
rect 28278 13732 28850 13792
rect 28278 13666 28338 13732
rect 27048 13660 27536 13666
rect 27048 13626 27060 13660
rect 27524 13626 27536 13660
rect 27048 13620 27536 13626
rect 28066 13660 28554 13666
rect 28066 13626 28078 13660
rect 28542 13626 28554 13660
rect 28066 13620 28554 13626
rect 26752 13536 26766 13576
rect 26760 13066 26766 13536
rect 25782 13000 25790 13060
rect 25012 12950 25500 12956
rect 25012 12916 25024 12950
rect 25488 12916 25500 12950
rect 25012 12910 25500 12916
rect 24522 12804 24776 12864
rect 24324 12588 24330 12648
rect 24390 12588 24396 12648
rect 24522 12538 24582 12804
rect 24712 12692 24718 12752
rect 24778 12692 24784 12752
rect 25220 12692 25226 12752
rect 25286 12692 25292 12752
rect 24522 12472 24582 12478
rect 23994 12428 24482 12434
rect 23994 12394 24006 12428
rect 24470 12394 24482 12428
rect 23994 12388 24482 12394
rect 24718 12344 24778 12692
rect 25226 12434 25286 12692
rect 25372 12648 25432 12910
rect 25730 12862 25790 13000
rect 26756 13000 26766 13066
rect 26800 13536 26812 13576
rect 27778 13576 27824 13588
rect 26800 13066 26806 13536
rect 26800 13000 26816 13066
rect 27778 13050 27784 13576
rect 26030 12950 26518 12956
rect 26030 12916 26042 12950
rect 26506 12916 26518 12950
rect 26030 12910 26518 12916
rect 25724 12802 25730 12862
rect 25790 12802 25796 12862
rect 25366 12588 25372 12648
rect 25432 12588 25438 12648
rect 25012 12428 25500 12434
rect 25012 12394 25024 12428
rect 25488 12394 25500 12428
rect 25012 12388 25500 12394
rect 25730 12344 25790 12802
rect 26234 12752 26294 12910
rect 26756 12752 26816 13000
rect 27768 13000 27784 13050
rect 27818 13050 27824 13576
rect 28790 13576 28850 13732
rect 29084 13660 29572 13666
rect 29084 13626 29096 13660
rect 29560 13626 29572 13660
rect 29084 13620 29572 13626
rect 30102 13660 30590 13666
rect 30102 13626 30114 13660
rect 30578 13626 30590 13660
rect 30102 13620 30590 13626
rect 28790 13550 28802 13576
rect 28796 13056 28802 13550
rect 27818 13000 27828 13050
rect 28788 13000 28802 13056
rect 28836 13550 28850 13576
rect 29814 13576 29860 13588
rect 28836 13056 28842 13550
rect 28836 13054 28848 13056
rect 28836 13000 28850 13054
rect 29814 13036 29820 13576
rect 27246 12956 27306 12958
rect 27048 12950 27536 12956
rect 27048 12916 27060 12950
rect 27524 12916 27536 12950
rect 27048 12910 27536 12916
rect 27246 12752 27306 12910
rect 27768 12862 27828 13000
rect 28278 12956 28338 12958
rect 28066 12950 28554 12956
rect 28066 12916 28078 12950
rect 28542 12916 28554 12950
rect 28066 12910 28554 12916
rect 27762 12802 27768 12862
rect 27828 12802 27834 12862
rect 26228 12692 26234 12752
rect 26294 12692 26300 12752
rect 26750 12692 26756 12752
rect 26816 12692 26822 12752
rect 27240 12692 27246 12752
rect 27306 12692 27312 12752
rect 26234 12434 26294 12692
rect 26750 12480 26756 12540
rect 26816 12480 26822 12540
rect 26030 12428 26518 12434
rect 26030 12394 26042 12428
rect 26506 12394 26518 12428
rect 26030 12388 26518 12394
rect 22728 12292 22738 12300
rect 23694 12296 23712 12344
rect 22728 11816 22734 12292
rect 23706 11816 23712 12296
rect 22728 11768 22740 11816
rect 21958 11718 22446 11724
rect 21958 11684 21970 11718
rect 22434 11684 22446 11718
rect 21958 11678 22446 11684
rect 22162 11618 22222 11678
rect 22680 11618 22740 11768
rect 23700 11768 23712 11816
rect 23746 12296 23754 12344
rect 24714 12304 24730 12344
rect 23746 11816 23752 12296
rect 23746 11768 23760 11816
rect 24724 11786 24730 12304
rect 22976 11718 23464 11724
rect 22976 11684 22988 11718
rect 23452 11684 23464 11718
rect 22976 11678 23464 11684
rect 23182 11618 23242 11678
rect 22162 11558 23242 11618
rect 23700 11546 23760 11768
rect 24718 11768 24730 11786
rect 24764 12306 24780 12344
rect 24764 12304 24778 12306
rect 24764 11786 24770 12304
rect 25730 12298 25748 12344
rect 25742 11822 25748 12298
rect 24764 11768 24778 11786
rect 23994 11718 24482 11724
rect 23994 11684 24006 11718
rect 24470 11684 24482 11718
rect 23994 11678 24482 11684
rect 24206 11622 24266 11678
rect 24718 11622 24778 11768
rect 25730 11768 25748 11822
rect 25782 12298 25790 12344
rect 26756 12344 26816 12480
rect 27246 12434 27306 12692
rect 27048 12428 27536 12434
rect 27048 12394 27060 12428
rect 27524 12394 27536 12428
rect 27048 12388 27536 12394
rect 26756 12302 26766 12344
rect 25782 11822 25788 12298
rect 25782 11768 25790 11822
rect 25012 11718 25500 11724
rect 25012 11684 25024 11718
rect 25488 11684 25500 11718
rect 25012 11678 25500 11684
rect 25208 11622 25268 11678
rect 24206 11562 25268 11622
rect 25730 11546 25790 11768
rect 26760 11768 26766 12302
rect 26800 12302 26816 12344
rect 27768 12344 27828 12802
rect 28278 12752 28338 12910
rect 28790 12752 28850 13000
rect 29806 13000 29820 13036
rect 29854 13036 29860 13576
rect 30824 13576 30884 13934
rect 31328 13666 31388 14144
rect 31844 14092 31904 14234
rect 32862 14234 32874 14810
rect 32908 14234 32922 14810
rect 33886 14810 33932 14822
rect 33886 14288 33892 14810
rect 32138 14184 32626 14190
rect 32138 14150 32150 14184
rect 32614 14150 32626 14184
rect 32138 14144 32626 14150
rect 31838 14032 31844 14092
rect 31904 14032 31910 14092
rect 31120 13660 31608 13666
rect 31120 13626 31132 13660
rect 31596 13626 31608 13660
rect 31120 13620 31608 13626
rect 30824 13536 30838 13576
rect 29854 13000 29866 13036
rect 29084 12950 29572 12956
rect 29084 12916 29096 12950
rect 29560 12916 29572 12950
rect 29084 12910 29572 12916
rect 29292 12862 29352 12910
rect 29806 12862 29866 13000
rect 30832 13000 30838 13536
rect 30872 13536 30884 13576
rect 31844 13576 31904 14032
rect 32354 13666 32414 14144
rect 32862 13994 32922 14234
rect 33874 14234 33892 14288
rect 33926 14288 33932 14810
rect 35766 14470 35878 15256
rect 33926 14234 33934 14288
rect 33156 14184 33644 14190
rect 33156 14150 33168 14184
rect 33632 14150 33644 14184
rect 33156 14144 33644 14150
rect 32856 13934 32862 13994
rect 32922 13934 32928 13994
rect 32138 13660 32626 13666
rect 32138 13626 32150 13660
rect 32614 13626 32626 13660
rect 32138 13620 32626 13626
rect 31844 13544 31856 13576
rect 30872 13000 30878 13536
rect 30832 12988 30878 13000
rect 31850 13000 31856 13544
rect 31890 13544 31904 13576
rect 32862 13576 32922 13934
rect 33376 13666 33436 14144
rect 33874 14092 33934 14234
rect 33868 14032 33874 14092
rect 33934 14032 33940 14092
rect 33156 13660 33644 13666
rect 33156 13626 33168 13660
rect 33632 13626 33644 13660
rect 33156 13620 33644 13626
rect 32862 13548 32874 13576
rect 31890 13000 31896 13544
rect 31850 12988 31896 13000
rect 32868 13000 32874 13548
rect 32908 13548 32922 13576
rect 33874 13576 33934 14032
rect 34592 13934 34598 13994
rect 34658 13934 34664 13994
rect 33874 13550 33892 13576
rect 32908 13000 32914 13548
rect 32868 12988 32914 13000
rect 33886 13000 33892 13550
rect 33926 13550 33934 13576
rect 33926 13000 33932 13550
rect 33886 12988 33932 13000
rect 30102 12950 30590 12956
rect 30102 12916 30114 12950
rect 30578 12916 30590 12950
rect 30102 12910 30590 12916
rect 31120 12950 31608 12956
rect 31120 12916 31132 12950
rect 31596 12916 31608 12950
rect 31120 12910 31608 12916
rect 32138 12950 32626 12956
rect 32138 12916 32150 12950
rect 32614 12916 32626 12950
rect 32138 12910 32626 12916
rect 33156 12950 33644 12956
rect 33156 12916 33168 12950
rect 33632 12916 33644 12950
rect 33156 12910 33644 12916
rect 30314 12862 30374 12910
rect 29800 12802 29806 12862
rect 29866 12802 29872 12862
rect 30308 12802 30314 12862
rect 30374 12802 30380 12862
rect 29292 12796 29352 12802
rect 28272 12692 28278 12752
rect 28338 12692 28344 12752
rect 28784 12692 28790 12752
rect 28850 12692 28856 12752
rect 28258 12588 28264 12648
rect 28324 12588 28330 12648
rect 29296 12588 29302 12648
rect 29362 12588 29368 12648
rect 28264 12434 28324 12588
rect 28782 12480 28788 12540
rect 28848 12480 28854 12540
rect 28066 12428 28554 12434
rect 28066 12394 28078 12428
rect 28542 12394 28554 12428
rect 28066 12388 28554 12394
rect 26800 11768 26806 12302
rect 26760 11756 26806 11768
rect 27768 11768 27784 12344
rect 27818 11768 27828 12344
rect 28788 12344 28848 12480
rect 29302 12434 29362 12588
rect 29084 12428 29572 12434
rect 29084 12394 29096 12428
rect 29560 12394 29572 12428
rect 29084 12388 29572 12394
rect 28788 12302 28802 12344
rect 26030 11718 26518 11724
rect 26030 11684 26042 11718
rect 26506 11684 26518 11718
rect 26030 11678 26518 11684
rect 27048 11718 27536 11724
rect 27048 11684 27060 11718
rect 27524 11684 27536 11718
rect 27048 11678 27536 11684
rect 26254 11576 27316 11636
rect 19620 11486 19626 11546
rect 19686 11486 19692 11546
rect 21656 11486 21662 11546
rect 21722 11486 21728 11546
rect 23694 11486 23700 11546
rect 23760 11486 23766 11546
rect 25724 11486 25730 11546
rect 25790 11486 25796 11546
rect 20640 11364 20646 11424
rect 20706 11364 20712 11424
rect 22674 11364 22680 11424
rect 22740 11364 22746 11424
rect 24704 11364 24710 11424
rect 24770 11364 24776 11424
rect 18902 11194 19390 11200
rect 18902 11160 18914 11194
rect 19378 11160 19390 11194
rect 18902 11154 19390 11160
rect 19920 11194 20408 11200
rect 19920 11160 19932 11194
rect 20396 11160 20408 11194
rect 19920 11154 20408 11160
rect 17636 10534 17642 11080
rect 18604 11066 18620 11110
rect 18614 10584 18620 11066
rect 17596 10522 17642 10534
rect 18606 10534 18620 10584
rect 18654 11066 18664 11110
rect 19632 11110 19678 11122
rect 18654 10584 18660 11066
rect 18654 10534 18666 10584
rect 19632 10570 19638 11110
rect 16866 10484 17354 10490
rect 16866 10450 16878 10484
rect 17342 10450 17354 10484
rect 16866 10444 17354 10450
rect 17884 10484 18372 10490
rect 17884 10450 17896 10484
rect 18360 10450 18372 10484
rect 17884 10444 18372 10450
rect 16564 10346 16570 10406
rect 16630 10346 16636 10406
rect 16060 10128 16066 10188
rect 16126 10128 16132 10188
rect 16066 9966 16126 10128
rect 15848 9960 16336 9966
rect 15848 9926 15860 9960
rect 16324 9926 16336 9960
rect 15848 9920 16336 9926
rect 14582 9300 14588 9840
rect 15552 9834 15566 9876
rect 15560 9358 15566 9834
rect 14542 9288 14588 9300
rect 15554 9300 15566 9358
rect 15600 9834 15612 9876
rect 16570 9876 16630 10346
rect 17068 10194 17128 10444
rect 17586 10242 17592 10302
rect 17652 10242 17658 10302
rect 17068 10188 17130 10194
rect 17068 10128 17070 10188
rect 17068 10122 17130 10128
rect 17068 9966 17128 10122
rect 16866 9960 17354 9966
rect 16866 9926 16878 9960
rect 17342 9926 17354 9960
rect 16866 9920 17354 9926
rect 15600 9358 15606 9834
rect 16570 9832 16584 9876
rect 15600 9300 15614 9358
rect 16578 9348 16584 9832
rect 13812 9250 14300 9256
rect 13812 9216 13824 9250
rect 14288 9216 14300 9250
rect 13812 9210 14300 9216
rect 14830 9250 15318 9256
rect 14830 9216 14842 9250
rect 15306 9216 15318 9250
rect 14830 9210 15318 9216
rect 14528 9090 14534 9150
rect 14594 9090 14600 9150
rect 13812 8728 14300 8734
rect 13812 8694 13824 8728
rect 14288 8694 14300 8728
rect 13812 8688 14300 8694
rect 13524 8644 13570 8656
rect 13524 8114 13530 8644
rect 13514 8068 13530 8114
rect 13564 8114 13570 8644
rect 14534 8644 14594 9090
rect 15040 9048 15100 9210
rect 15034 8988 15040 9048
rect 15100 8988 15106 9048
rect 15554 8846 15614 9300
rect 16572 9300 16584 9348
rect 16618 9832 16630 9876
rect 17592 9876 17652 10242
rect 18084 10194 18144 10444
rect 18606 10406 18666 10534
rect 19624 10534 19638 10570
rect 19672 10570 19678 11110
rect 20646 11110 20706 11364
rect 20938 11194 21426 11200
rect 20938 11160 20950 11194
rect 21414 11160 21426 11194
rect 20938 11154 21426 11160
rect 21956 11194 22444 11200
rect 21956 11160 21968 11194
rect 22432 11160 22444 11194
rect 21956 11154 22444 11160
rect 20646 11054 20656 11110
rect 19672 10534 19684 10570
rect 18902 10484 19390 10490
rect 18902 10450 18914 10484
rect 19378 10450 19390 10484
rect 18902 10444 19390 10450
rect 18600 10346 18606 10406
rect 18666 10346 18672 10406
rect 18082 10188 18144 10194
rect 18142 10128 18144 10188
rect 18082 10122 18144 10128
rect 18084 9966 18144 10122
rect 17884 9960 18372 9966
rect 17884 9926 17896 9960
rect 18360 9926 18372 9960
rect 17884 9920 18372 9926
rect 17592 9834 17602 9876
rect 16618 9348 16624 9832
rect 16618 9300 16632 9348
rect 15848 9250 16336 9256
rect 15848 9216 15860 9250
rect 16324 9216 16336 9250
rect 15848 9210 16336 9216
rect 16572 9150 16632 9300
rect 17596 9300 17602 9834
rect 17636 9834 17652 9876
rect 18606 9876 18666 10346
rect 19102 10188 19162 10444
rect 19624 10302 19684 10534
rect 20650 10534 20656 11054
rect 20690 11054 20706 11110
rect 21668 11110 21714 11122
rect 20690 10534 20696 11054
rect 21668 10564 21674 11110
rect 20650 10522 20696 10534
rect 21658 10534 21674 10564
rect 21708 10564 21714 11110
rect 22680 11110 22740 11364
rect 22974 11194 23462 11200
rect 22974 11160 22986 11194
rect 23450 11160 23462 11194
rect 22974 11154 23462 11160
rect 23992 11194 24480 11200
rect 23992 11160 24004 11194
rect 24468 11160 24480 11194
rect 23992 11154 24480 11160
rect 22680 11060 22692 11110
rect 21708 10534 21718 10564
rect 19920 10484 20408 10490
rect 19920 10450 19932 10484
rect 20396 10450 20408 10484
rect 19920 10444 20408 10450
rect 20938 10484 21426 10490
rect 20938 10450 20950 10484
rect 21414 10450 21426 10484
rect 20938 10444 21426 10450
rect 19618 10242 19624 10302
rect 19684 10242 19690 10302
rect 20114 10246 20174 10444
rect 21156 10246 21216 10444
rect 21658 10302 21718 10534
rect 22686 10534 22692 11060
rect 22726 11060 22740 11110
rect 23704 11110 23750 11122
rect 22726 10534 22732 11060
rect 23704 10576 23710 11110
rect 22686 10522 22732 10534
rect 23698 10534 23710 10576
rect 23744 10576 23750 11110
rect 24710 11110 24770 11364
rect 26254 11200 26314 11576
rect 26744 11486 26750 11546
rect 26810 11486 26816 11546
rect 25010 11194 25498 11200
rect 25010 11160 25022 11194
rect 25486 11160 25498 11194
rect 25010 11154 25498 11160
rect 26028 11194 26516 11200
rect 26028 11160 26040 11194
rect 26504 11160 26516 11194
rect 26028 11154 26516 11160
rect 24710 11066 24728 11110
rect 23744 10534 23758 10576
rect 21956 10484 22444 10490
rect 21956 10450 21968 10484
rect 22432 10450 22444 10484
rect 21956 10444 22444 10450
rect 22974 10484 23462 10490
rect 22974 10450 22986 10484
rect 23450 10450 23462 10484
rect 22974 10444 23462 10450
rect 19618 10130 19624 10190
rect 19684 10130 19690 10190
rect 20114 10186 21216 10246
rect 21652 10242 21658 10302
rect 21718 10242 21724 10302
rect 19102 9966 19162 10128
rect 18902 9960 19390 9966
rect 18902 9926 18914 9960
rect 19378 9926 19390 9960
rect 18902 9920 19390 9926
rect 17636 9300 17642 9834
rect 18606 9828 18620 9876
rect 18614 9350 18620 9828
rect 17596 9288 17642 9300
rect 18608 9300 18620 9350
rect 18654 9828 18666 9876
rect 19624 9876 19684 10130
rect 20114 9966 20174 10186
rect 20636 10020 20642 10080
rect 20702 10020 20708 10080
rect 19920 9960 20408 9966
rect 19920 9926 19932 9960
rect 20396 9926 20408 9960
rect 19920 9920 20408 9926
rect 18654 9350 18660 9828
rect 19624 9818 19638 9876
rect 18654 9300 18668 9350
rect 16866 9250 17354 9256
rect 16866 9216 16878 9250
rect 17342 9216 17354 9250
rect 16866 9210 17354 9216
rect 17884 9250 18372 9256
rect 17884 9216 17896 9250
rect 18360 9216 18372 9250
rect 17884 9210 18372 9216
rect 16566 9090 16572 9150
rect 16632 9090 16638 9150
rect 16564 8886 16570 8946
rect 16630 8886 16636 8946
rect 17078 8940 17138 9210
rect 18100 8940 18160 9210
rect 18608 9150 18668 9300
rect 19632 9300 19638 9818
rect 19672 9818 19684 9876
rect 20642 9876 20702 10020
rect 21156 9966 21216 10186
rect 21654 10130 21660 10190
rect 21720 10130 21726 10190
rect 20938 9960 21426 9966
rect 20938 9926 20950 9960
rect 21414 9926 21426 9960
rect 20938 9920 21426 9926
rect 20642 9830 20656 9876
rect 19672 9300 19678 9818
rect 19632 9288 19678 9300
rect 20650 9300 20656 9830
rect 20690 9830 20702 9876
rect 21660 9876 21720 10130
rect 22156 9966 22216 10444
rect 22670 10020 22676 10080
rect 22736 10020 22742 10080
rect 21956 9960 22444 9966
rect 21956 9926 21968 9960
rect 22432 9926 22444 9960
rect 21956 9920 22444 9926
rect 20690 9300 20696 9830
rect 21660 9808 21674 9876
rect 20650 9288 20696 9300
rect 21668 9300 21674 9808
rect 21708 9808 21720 9876
rect 22676 9876 22736 10020
rect 23190 9966 23250 10444
rect 23698 10302 23758 10534
rect 24722 10534 24728 11066
rect 24762 11066 24770 11110
rect 25740 11110 25786 11122
rect 24762 10534 24768 11066
rect 25740 10586 25746 11110
rect 24722 10522 24768 10534
rect 25732 10534 25746 10586
rect 25780 10586 25786 11110
rect 26750 11110 26810 11486
rect 27256 11370 27316 11576
rect 27768 11546 27828 11768
rect 28796 11768 28802 12302
rect 28836 12302 28848 12344
rect 29806 12344 29866 12802
rect 31328 12692 31334 12752
rect 31394 12692 31400 12752
rect 32348 12692 32354 12752
rect 32414 12692 32420 12752
rect 30296 12588 30302 12648
rect 30362 12588 30368 12648
rect 30302 12434 30362 12588
rect 30814 12480 30820 12540
rect 30880 12480 30886 12540
rect 30102 12428 30590 12434
rect 30102 12394 30114 12428
rect 30578 12394 30590 12428
rect 30102 12388 30590 12394
rect 30302 12376 30362 12388
rect 28836 11768 28842 12302
rect 29806 12286 29820 12344
rect 29814 11816 29820 12286
rect 28796 11756 28842 11768
rect 29804 11768 29820 11816
rect 29854 12286 29866 12344
rect 30820 12344 30880 12480
rect 31334 12434 31394 12692
rect 32354 12434 32414 12692
rect 32856 12480 32862 12540
rect 32922 12480 32928 12540
rect 33360 12480 33366 12540
rect 33426 12480 33432 12540
rect 33870 12480 33876 12540
rect 33936 12480 33942 12540
rect 31120 12428 31608 12434
rect 31120 12394 31132 12428
rect 31596 12394 31608 12428
rect 31120 12388 31608 12394
rect 32138 12428 32626 12434
rect 32138 12394 32150 12428
rect 32614 12394 32626 12428
rect 32138 12388 32626 12394
rect 30820 12298 30838 12344
rect 29854 11816 29860 12286
rect 29854 11768 29864 11816
rect 28066 11718 28554 11724
rect 28066 11684 28078 11718
rect 28542 11684 28554 11718
rect 28066 11678 28554 11684
rect 29084 11718 29572 11724
rect 29084 11684 29096 11718
rect 29560 11684 29572 11718
rect 29084 11678 29572 11684
rect 28268 11650 28328 11678
rect 29302 11650 29362 11678
rect 28260 11590 28266 11650
rect 28326 11590 28332 11650
rect 29296 11590 29302 11650
rect 29362 11590 29368 11650
rect 27762 11486 27768 11546
rect 27828 11486 27834 11546
rect 28268 11370 28328 11590
rect 28782 11486 28788 11546
rect 28848 11486 28854 11546
rect 27256 11310 28328 11370
rect 27256 11200 27316 11310
rect 28268 11200 28328 11310
rect 27046 11194 27534 11200
rect 27046 11160 27058 11194
rect 27522 11160 27534 11194
rect 27046 11154 27534 11160
rect 28064 11194 28552 11200
rect 28064 11160 28076 11194
rect 28540 11160 28552 11194
rect 28064 11154 28552 11160
rect 26750 11062 26764 11110
rect 25780 10534 25792 10586
rect 26758 10566 26764 11062
rect 23992 10484 24480 10490
rect 23992 10450 24004 10484
rect 24468 10450 24480 10484
rect 23992 10444 24480 10450
rect 25010 10484 25498 10490
rect 25010 10450 25022 10484
rect 25486 10450 25498 10484
rect 25010 10444 25498 10450
rect 23692 10242 23698 10302
rect 23758 10242 23764 10302
rect 24212 10246 24272 10444
rect 25220 10246 25280 10444
rect 25732 10302 25792 10534
rect 26750 10534 26764 10566
rect 26798 11062 26810 11110
rect 27776 11110 27822 11122
rect 26798 10566 26804 11062
rect 27776 10570 27782 11110
rect 26798 10534 26810 10566
rect 26028 10484 26516 10490
rect 26028 10450 26040 10484
rect 26504 10450 26516 10484
rect 26028 10444 26516 10450
rect 23690 10130 23696 10190
rect 23756 10130 23762 10190
rect 24212 10186 25280 10246
rect 25726 10242 25732 10302
rect 25792 10242 25798 10302
rect 25922 10238 25928 10298
rect 25988 10238 25994 10298
rect 22974 9960 23462 9966
rect 22974 9926 22986 9960
rect 23450 9926 23462 9960
rect 22974 9920 23462 9926
rect 22676 9828 22692 9876
rect 21708 9300 21714 9808
rect 21668 9288 21714 9300
rect 22686 9300 22692 9828
rect 22726 9828 22736 9876
rect 23696 9876 23756 10130
rect 24212 9966 24272 10186
rect 24710 10020 24716 10080
rect 24776 10020 24782 10080
rect 23992 9960 24480 9966
rect 23992 9926 24004 9960
rect 24468 9926 24480 9960
rect 23992 9920 24480 9926
rect 22726 9300 22732 9828
rect 23696 9826 23710 9876
rect 22686 9288 22732 9300
rect 23704 9300 23710 9826
rect 23744 9826 23756 9876
rect 24716 9876 24776 10020
rect 25220 9966 25280 10186
rect 25726 10130 25732 10190
rect 25792 10130 25798 10190
rect 25010 9960 25498 9966
rect 25010 9926 25022 9960
rect 25486 9926 25498 9960
rect 25010 9920 25498 9926
rect 24716 9838 24728 9876
rect 23744 9300 23750 9826
rect 24722 9346 24728 9838
rect 23704 9288 23750 9300
rect 24716 9300 24728 9346
rect 24762 9838 24776 9876
rect 25732 9876 25792 10130
rect 25928 10080 25988 10238
rect 26222 10082 26282 10444
rect 26750 10406 26810 10534
rect 27766 10534 27782 10570
rect 27816 10570 27822 11110
rect 28788 11110 28848 11486
rect 29302 11362 29362 11590
rect 29804 11546 29864 11768
rect 30832 11768 30838 12298
rect 30872 12298 30880 12344
rect 31850 12344 31896 12356
rect 30872 11768 30878 12298
rect 31850 11826 31856 12344
rect 30832 11756 30878 11768
rect 31840 11768 31856 11826
rect 31890 11826 31896 12344
rect 32862 12344 32922 12480
rect 33366 12434 33426 12480
rect 33156 12428 33644 12434
rect 33156 12394 33168 12428
rect 33632 12394 33644 12428
rect 33156 12388 33644 12394
rect 32862 12288 32874 12344
rect 31890 11768 31900 11826
rect 30102 11718 30590 11724
rect 30102 11684 30114 11718
rect 30578 11684 30590 11718
rect 30102 11678 30590 11684
rect 31120 11718 31608 11724
rect 31120 11684 31132 11718
rect 31596 11684 31608 11718
rect 31120 11678 31608 11684
rect 30318 11650 30378 11678
rect 30312 11590 30318 11650
rect 30378 11590 30384 11650
rect 31840 11546 31900 11768
rect 32868 11768 32874 12288
rect 32908 12288 32922 12344
rect 33876 12344 33936 12480
rect 33876 12308 33892 12344
rect 32908 11768 32914 12288
rect 32868 11756 32914 11768
rect 33886 11768 33892 12308
rect 33926 12308 33936 12344
rect 33926 11768 33932 12308
rect 33886 11756 33932 11768
rect 32138 11718 32626 11724
rect 32138 11684 32150 11718
rect 32614 11684 32626 11718
rect 32138 11678 32626 11684
rect 33156 11718 33644 11724
rect 33156 11684 33168 11718
rect 33632 11684 33644 11718
rect 33156 11678 33644 11684
rect 29798 11486 29804 11546
rect 29864 11486 29870 11546
rect 31834 11486 31840 11546
rect 31900 11486 31906 11546
rect 29302 11302 32390 11362
rect 29302 11200 29362 11302
rect 32330 11200 32390 11302
rect 33368 11276 33936 11336
rect 33368 11200 33428 11276
rect 29082 11194 29570 11200
rect 29082 11160 29094 11194
rect 29558 11160 29570 11194
rect 29082 11154 29570 11160
rect 30100 11194 30588 11200
rect 30100 11160 30112 11194
rect 30576 11160 30588 11194
rect 30100 11154 30588 11160
rect 31118 11194 31606 11200
rect 31118 11160 31130 11194
rect 31594 11160 31606 11194
rect 31118 11154 31606 11160
rect 32136 11194 32624 11200
rect 32136 11160 32148 11194
rect 32612 11160 32624 11194
rect 32136 11154 32624 11160
rect 33154 11194 33642 11200
rect 33154 11160 33166 11194
rect 33630 11160 33642 11194
rect 33154 11154 33642 11160
rect 28788 11052 28800 11110
rect 28794 10580 28800 11052
rect 27816 10534 27826 10570
rect 27046 10484 27534 10490
rect 27046 10450 27058 10484
rect 27522 10450 27534 10484
rect 27046 10444 27534 10450
rect 26744 10346 26750 10406
rect 26810 10346 26816 10406
rect 25922 10020 25928 10080
rect 25988 10020 25994 10080
rect 26216 10022 26222 10082
rect 26282 10022 26288 10082
rect 26222 9966 26282 10022
rect 26028 9960 26516 9966
rect 26028 9926 26040 9960
rect 26504 9926 26516 9960
rect 26028 9920 26516 9926
rect 24762 9346 24768 9838
rect 25732 9832 25746 9876
rect 24762 9300 24776 9346
rect 18902 9250 19390 9256
rect 18902 9216 18914 9250
rect 19378 9216 19390 9250
rect 18902 9210 19390 9216
rect 19920 9250 20408 9256
rect 19920 9216 19932 9250
rect 20396 9216 20408 9250
rect 19920 9210 20408 9216
rect 20938 9250 21426 9256
rect 20938 9216 20950 9250
rect 21414 9216 21426 9250
rect 20938 9210 21426 9216
rect 21956 9250 22444 9256
rect 21956 9216 21968 9250
rect 22432 9216 22444 9250
rect 21956 9210 22444 9216
rect 22974 9250 23462 9256
rect 22974 9216 22986 9250
rect 23450 9216 23462 9250
rect 22974 9210 23462 9216
rect 23992 9250 24480 9256
rect 23992 9216 24004 9250
rect 24468 9216 24480 9250
rect 23992 9210 24480 9216
rect 18602 9090 18608 9150
rect 18668 9090 18674 9150
rect 15548 8786 15554 8846
rect 15614 8786 15620 8846
rect 14830 8728 15318 8734
rect 14830 8694 14842 8728
rect 15306 8694 15318 8728
rect 14830 8688 15318 8694
rect 14534 8606 14548 8644
rect 13564 8068 13574 8114
rect 14542 8110 14548 8606
rect 13514 7906 13574 8068
rect 14532 8068 14548 8110
rect 14582 8606 14594 8644
rect 15554 8644 15614 8786
rect 15848 8728 16336 8734
rect 15848 8694 15860 8728
rect 16324 8694 16336 8728
rect 15848 8688 16336 8694
rect 14582 8110 14588 8606
rect 15554 8604 15566 8644
rect 14582 8068 14592 8110
rect 13812 8018 14300 8024
rect 13812 7984 13824 8018
rect 14288 7984 14300 8018
rect 13812 7978 14300 7984
rect 14026 7906 14086 7978
rect 14532 7906 14592 8068
rect 15560 8068 15566 8604
rect 15600 8604 15614 8644
rect 16570 8644 16630 8886
rect 17072 8880 17078 8940
rect 17138 8880 17144 8940
rect 18094 8880 18100 8940
rect 18160 8880 18166 8940
rect 17582 8786 17588 8846
rect 17648 8786 17654 8846
rect 16866 8728 17354 8734
rect 16866 8694 16878 8728
rect 17342 8694 17354 8728
rect 16866 8688 17354 8694
rect 15600 8068 15606 8604
rect 16570 8592 16584 8644
rect 15560 8056 15606 8068
rect 16578 8068 16584 8592
rect 16618 8592 16630 8644
rect 17588 8644 17648 8786
rect 18100 8734 18160 8880
rect 17884 8728 18372 8734
rect 17884 8694 17896 8728
rect 18360 8694 18372 8728
rect 17884 8688 18372 8694
rect 17588 8600 17602 8644
rect 16618 8068 16624 8592
rect 17596 8104 17602 8600
rect 16578 8056 16624 8068
rect 17588 8068 17602 8104
rect 17636 8600 17648 8644
rect 18608 8644 18668 9090
rect 19114 8940 19174 9210
rect 20132 9048 20192 9210
rect 21152 9160 21212 9210
rect 22152 9160 22212 9210
rect 23190 9160 23250 9210
rect 24218 9160 24278 9210
rect 20634 9090 20640 9150
rect 20700 9090 20706 9150
rect 21152 9100 24278 9160
rect 20126 8988 20132 9048
rect 20192 8988 20198 9048
rect 19108 8880 19114 8940
rect 19174 8880 19180 8940
rect 20126 8880 20132 8940
rect 20192 8880 20198 8940
rect 19114 8734 19174 8880
rect 19618 8786 19624 8846
rect 19684 8786 19690 8846
rect 18902 8728 19390 8734
rect 18902 8694 18914 8728
rect 19378 8694 19390 8728
rect 18902 8688 19390 8694
rect 17636 8104 17642 8600
rect 17636 8068 17648 8104
rect 14830 8018 15318 8024
rect 14830 7984 14842 8018
rect 15306 7984 15318 8018
rect 14830 7978 15318 7984
rect 15848 8018 16336 8024
rect 15848 7984 15860 8018
rect 16324 7984 16336 8018
rect 15848 7978 16336 7984
rect 16866 8018 17354 8024
rect 16866 7984 16878 8018
rect 17342 7984 17354 8018
rect 16866 7978 17354 7984
rect 15036 7922 15096 7978
rect 13514 7846 14592 7906
rect 15030 7862 15036 7922
rect 15096 7862 15102 7922
rect 15940 7862 15946 7922
rect 16006 7862 16012 7922
rect 15030 7646 15036 7706
rect 15096 7646 15102 7706
rect 15036 7640 15098 7646
rect 13398 7602 13460 7608
rect 13398 7542 13400 7602
rect 13398 7536 13460 7542
rect 13280 6284 13286 6344
rect 13346 6284 13352 6344
rect 13180 5280 13244 5286
rect 13180 5228 13192 5280
rect 13180 5222 13244 5228
rect 13180 4100 13240 5222
rect 13286 4226 13346 6284
rect 13398 5358 13458 7536
rect 15038 7500 15098 7640
rect 15946 7500 16006 7862
rect 16074 7706 16134 7978
rect 16942 7862 16948 7922
rect 17008 7862 17014 7922
rect 16074 7640 16134 7646
rect 16948 7500 17008 7862
rect 17088 7706 17148 7978
rect 17588 7820 17648 8068
rect 18608 8068 18620 8644
rect 18654 8068 18668 8644
rect 19624 8644 19684 8786
rect 20132 8734 20192 8880
rect 19920 8728 20408 8734
rect 19920 8694 19932 8728
rect 20396 8694 20408 8728
rect 19920 8688 20408 8694
rect 19624 8608 19638 8644
rect 17884 8018 18372 8024
rect 17884 7984 17896 8018
rect 18360 7984 18372 8018
rect 17884 7978 18372 7984
rect 18100 7922 18160 7978
rect 18094 7862 18100 7922
rect 18160 7862 18166 7922
rect 17582 7760 17588 7820
rect 17648 7760 17654 7820
rect 17082 7646 17088 7706
rect 17148 7646 17154 7706
rect 18100 7500 18160 7862
rect 13812 7494 14300 7500
rect 13812 7460 13824 7494
rect 14288 7460 14300 7494
rect 13812 7454 14300 7460
rect 14830 7494 15318 7500
rect 14830 7460 14842 7494
rect 15306 7460 15318 7494
rect 14830 7454 15318 7460
rect 15848 7494 16336 7500
rect 15848 7460 15860 7494
rect 16324 7460 16336 7494
rect 15848 7454 16336 7460
rect 16866 7494 17354 7500
rect 16866 7460 16878 7494
rect 17342 7460 17354 7494
rect 16866 7454 17354 7460
rect 17884 7494 18372 7500
rect 17884 7460 17896 7494
rect 18360 7460 18372 7494
rect 17884 7454 18372 7460
rect 13524 7410 13570 7422
rect 13524 6872 13530 7410
rect 13518 6834 13530 6872
rect 13564 6872 13570 7410
rect 14542 7410 14588 7422
rect 14542 6872 14548 7410
rect 13564 6834 13578 6872
rect 13518 6704 13578 6834
rect 14536 6834 14548 6872
rect 14582 6872 14588 7410
rect 15560 7410 15606 7422
rect 15560 6884 15566 7410
rect 14582 6834 14596 6872
rect 13812 6784 14300 6790
rect 13812 6750 13824 6784
rect 14288 6750 14300 6784
rect 13812 6744 14300 6750
rect 14016 6704 14076 6744
rect 14536 6704 14596 6834
rect 15552 6834 15566 6884
rect 15600 6884 15606 7410
rect 16578 7410 16624 7422
rect 16578 6892 16584 7410
rect 15600 6834 15612 6884
rect 14830 6784 15318 6790
rect 14830 6750 14842 6784
rect 15306 6750 15318 6784
rect 14830 6744 15318 6750
rect 13518 6644 14596 6704
rect 14536 6590 14596 6644
rect 15028 6634 15034 6694
rect 15094 6634 15100 6694
rect 14530 6530 14536 6590
rect 14596 6530 14602 6590
rect 14526 6320 14532 6380
rect 14592 6320 14598 6380
rect 13812 6260 14300 6266
rect 13812 6226 13824 6260
rect 14288 6226 14300 6260
rect 13812 6220 14300 6226
rect 13524 6176 13570 6188
rect 13524 5634 13530 6176
rect 13514 5600 13530 5634
rect 13564 5634 13570 6176
rect 14532 6176 14592 6320
rect 15034 6266 15094 6634
rect 15552 6478 15612 6834
rect 16570 6834 16584 6892
rect 16618 6892 16624 7410
rect 17596 7410 17642 7422
rect 16618 6834 16630 6892
rect 17596 6880 17602 7410
rect 15848 6784 16336 6790
rect 15848 6750 15860 6784
rect 16324 6750 16336 6784
rect 15848 6744 16336 6750
rect 16042 6694 16102 6744
rect 16036 6634 16042 6694
rect 16102 6634 16108 6694
rect 15546 6418 15552 6478
rect 15612 6418 15618 6478
rect 16570 6380 16630 6834
rect 17590 6834 17602 6880
rect 17636 6880 17642 7410
rect 18608 7410 18668 8068
rect 19632 8068 19638 8608
rect 19672 8608 19684 8644
rect 20640 8644 20700 9090
rect 21146 8880 21152 8940
rect 21212 8880 21218 8940
rect 24218 8924 24278 9100
rect 24716 9034 24776 9300
rect 25740 9300 25746 9832
rect 25780 9832 25792 9876
rect 26750 9876 26810 10346
rect 27252 10088 27312 10444
rect 27766 10190 27826 10534
rect 28786 10534 28800 10580
rect 28834 11052 28848 11110
rect 29812 11110 29858 11122
rect 28834 10580 28840 11052
rect 29812 10590 29818 11110
rect 28834 10534 28846 10580
rect 28064 10484 28552 10490
rect 28064 10450 28076 10484
rect 28540 10450 28552 10484
rect 28064 10444 28552 10450
rect 27760 10130 27766 10190
rect 27826 10130 27832 10190
rect 27250 10082 27312 10088
rect 27310 10022 27312 10082
rect 27250 10016 27312 10022
rect 27762 10016 27768 10076
rect 27828 10016 27834 10076
rect 27252 9966 27312 10016
rect 27046 9960 27534 9966
rect 27046 9926 27058 9960
rect 27522 9926 27534 9960
rect 27046 9920 27534 9926
rect 26750 9832 26764 9876
rect 25780 9300 25786 9832
rect 25740 9288 25786 9300
rect 26758 9300 26764 9832
rect 26798 9832 26810 9876
rect 27768 9876 27828 10016
rect 28276 9966 28336 10444
rect 28786 10406 28846 10534
rect 29804 10534 29818 10590
rect 29852 10590 29858 11110
rect 30830 11110 30876 11122
rect 29852 10534 29864 10590
rect 30830 10578 30836 11110
rect 29082 10484 29570 10490
rect 29082 10450 29094 10484
rect 29558 10450 29570 10484
rect 29082 10444 29570 10450
rect 28780 10346 28786 10406
rect 28846 10346 28852 10406
rect 28064 9960 28552 9966
rect 28064 9926 28076 9960
rect 28540 9926 28552 9960
rect 28064 9920 28552 9926
rect 27768 9846 27782 9876
rect 26798 9300 26804 9832
rect 27776 9340 27782 9846
rect 26758 9288 26804 9300
rect 27768 9300 27782 9340
rect 27816 9846 27828 9876
rect 28786 9876 28846 10346
rect 29302 9966 29362 10444
rect 29804 10190 29864 10534
rect 30820 10534 30836 10578
rect 30870 10578 30876 11110
rect 31848 11110 31894 11122
rect 31848 10578 31854 11110
rect 30870 10534 30880 10578
rect 30100 10484 30588 10490
rect 30100 10450 30112 10484
rect 30576 10450 30588 10484
rect 30100 10444 30588 10450
rect 29798 10130 29804 10190
rect 29864 10130 29870 10190
rect 30310 10140 30370 10444
rect 30820 10298 30880 10534
rect 31844 10534 31854 10578
rect 31888 10578 31894 11110
rect 32866 11110 32912 11122
rect 32866 10584 32872 11110
rect 31888 10534 31904 10578
rect 31118 10484 31606 10490
rect 31118 10450 31130 10484
rect 31594 10450 31606 10484
rect 31118 10444 31606 10450
rect 31326 10300 31386 10444
rect 30814 10238 30820 10298
rect 30880 10238 30886 10298
rect 31324 10294 31386 10300
rect 31384 10234 31386 10294
rect 31324 10228 31386 10234
rect 31326 10140 31386 10228
rect 31844 10190 31904 10534
rect 32860 10534 32872 10584
rect 32906 10584 32912 11110
rect 33876 11110 33936 11276
rect 33978 11252 33984 11312
rect 34044 11252 34050 11312
rect 33876 11082 33890 11110
rect 33884 10592 33890 11082
rect 32906 10534 32920 10584
rect 32136 10484 32624 10490
rect 32136 10450 32148 10484
rect 32612 10450 32624 10484
rect 32136 10444 32624 10450
rect 30310 10080 31386 10140
rect 31838 10130 31844 10190
rect 31904 10130 31910 10190
rect 29798 10016 29804 10076
rect 29864 10016 29870 10076
rect 29082 9960 29570 9966
rect 29082 9926 29094 9960
rect 29558 9926 29570 9960
rect 29082 9920 29570 9926
rect 27816 9340 27822 9846
rect 28786 9836 28800 9876
rect 27816 9300 27828 9340
rect 28794 9334 28800 9836
rect 25010 9250 25498 9256
rect 25010 9216 25022 9250
rect 25486 9216 25498 9250
rect 25010 9210 25498 9216
rect 26028 9250 26516 9256
rect 26028 9216 26040 9250
rect 26504 9216 26516 9250
rect 26028 9210 26516 9216
rect 27046 9250 27534 9256
rect 27046 9216 27058 9250
rect 27522 9216 27534 9250
rect 27046 9210 27534 9216
rect 25222 9162 25282 9210
rect 24710 8974 24716 9034
rect 24776 8974 24782 9034
rect 25222 8924 25282 9102
rect 21152 8734 21212 8880
rect 24218 8864 25282 8924
rect 26746 8776 26752 8836
rect 26812 8776 26818 8836
rect 20938 8728 21426 8734
rect 20938 8694 20950 8728
rect 21414 8694 21426 8728
rect 20938 8688 21426 8694
rect 21956 8728 22444 8734
rect 21956 8694 21968 8728
rect 22432 8694 22444 8728
rect 21956 8688 22444 8694
rect 22974 8728 23462 8734
rect 22974 8694 22986 8728
rect 23450 8694 23462 8728
rect 22974 8688 23462 8694
rect 23992 8728 24480 8734
rect 23992 8694 24004 8728
rect 24468 8694 24480 8728
rect 23992 8688 24480 8694
rect 25010 8728 25498 8734
rect 25010 8694 25022 8728
rect 25486 8694 25498 8728
rect 25010 8688 25498 8694
rect 26028 8728 26516 8734
rect 26028 8694 26040 8728
rect 26504 8694 26516 8728
rect 26028 8688 26516 8694
rect 19672 8068 19678 8608
rect 20640 8606 20656 8644
rect 19632 8056 19678 8068
rect 20650 8068 20656 8606
rect 20690 8606 20700 8644
rect 21668 8644 21714 8656
rect 20690 8068 20696 8606
rect 21668 8110 21674 8644
rect 20650 8056 20696 8068
rect 21660 8068 21674 8110
rect 21708 8110 21714 8644
rect 22686 8644 22732 8656
rect 21708 8068 21720 8110
rect 22686 8106 22692 8644
rect 18902 8018 19390 8024
rect 18902 7984 18914 8018
rect 19378 7984 19390 8018
rect 18902 7978 19390 7984
rect 19920 8018 20408 8024
rect 19920 7984 19932 8018
rect 20396 7984 20408 8018
rect 19920 7978 20408 7984
rect 20938 8018 21426 8024
rect 20938 7984 20950 8018
rect 21414 7984 21426 8018
rect 20938 7978 21426 7984
rect 19110 7922 19170 7978
rect 20116 7922 20176 7978
rect 21160 7922 21220 7978
rect 21660 7928 21720 8068
rect 22680 8068 22692 8106
rect 22726 8106 22732 8644
rect 23704 8644 23750 8656
rect 22726 8068 22740 8106
rect 23704 8100 23710 8644
rect 21956 8018 22444 8024
rect 21956 7984 21968 8018
rect 22432 7984 22444 8018
rect 21956 7978 22444 7984
rect 19104 7862 19110 7922
rect 19170 7862 19176 7922
rect 20110 7862 20116 7922
rect 20176 7862 20182 7922
rect 21154 7862 21160 7922
rect 21220 7862 21226 7922
rect 21654 7868 21660 7928
rect 21720 7868 21726 7928
rect 19110 7500 19170 7862
rect 20108 7646 20114 7706
rect 20174 7646 20180 7706
rect 21148 7646 21154 7706
rect 21214 7646 21220 7706
rect 20114 7500 20174 7646
rect 20632 7542 20638 7602
rect 20698 7542 20704 7602
rect 18902 7494 19390 7500
rect 18902 7460 18914 7494
rect 19378 7460 19390 7494
rect 18902 7454 19390 7460
rect 19920 7494 20408 7500
rect 19920 7460 19932 7494
rect 20396 7460 20408 7494
rect 19920 7454 20408 7460
rect 18608 7328 18620 7410
rect 18614 6880 18620 7328
rect 17636 6834 17650 6880
rect 16866 6784 17354 6790
rect 16866 6750 16878 6784
rect 17342 6750 17354 6784
rect 16866 6744 17354 6750
rect 17056 6694 17116 6744
rect 17050 6634 17056 6694
rect 17116 6634 17122 6694
rect 17590 6478 17650 6834
rect 18610 6834 18620 6880
rect 18654 7328 18668 7410
rect 19632 7410 19678 7422
rect 18654 6880 18660 7328
rect 18654 6834 18670 6880
rect 19632 6878 19638 7410
rect 17884 6784 18372 6790
rect 17884 6750 17896 6784
rect 18360 6750 18372 6784
rect 17884 6744 18372 6750
rect 18094 6694 18154 6744
rect 18088 6634 18094 6694
rect 18154 6634 18160 6694
rect 17584 6418 17590 6478
rect 17650 6418 17656 6478
rect 16564 6320 16570 6380
rect 16630 6320 16636 6380
rect 18094 6266 18154 6634
rect 18610 6380 18670 6834
rect 19628 6834 19638 6878
rect 19672 6878 19678 7410
rect 20638 7410 20698 7542
rect 21154 7500 21214 7646
rect 20938 7494 21426 7500
rect 20938 7460 20950 7494
rect 21414 7460 21426 7494
rect 20938 7454 21426 7460
rect 20638 7346 20656 7410
rect 19672 6834 19688 6878
rect 18902 6784 19390 6790
rect 18902 6750 18914 6784
rect 19378 6750 19390 6784
rect 18902 6744 19390 6750
rect 19112 6694 19172 6744
rect 19628 6700 19688 6834
rect 20650 6834 20656 7346
rect 20690 7346 20698 7410
rect 21660 7410 21720 7868
rect 22168 7706 22228 7978
rect 22162 7646 22168 7706
rect 22228 7646 22234 7706
rect 22168 7500 22228 7646
rect 22680 7602 22740 8068
rect 23696 8068 23710 8100
rect 23744 8100 23750 8644
rect 24722 8644 24768 8656
rect 24722 8102 24728 8644
rect 23744 8068 23756 8100
rect 22974 8018 23462 8024
rect 22974 7984 22986 8018
rect 23450 7984 23462 8018
rect 22974 7978 23462 7984
rect 23176 7706 23236 7978
rect 23696 7928 23756 8068
rect 24718 8068 24728 8102
rect 24762 8102 24768 8644
rect 25740 8644 25786 8656
rect 24762 8068 24778 8102
rect 25740 8100 25746 8644
rect 23992 8018 24480 8024
rect 23992 7984 24004 8018
rect 24468 7984 24480 8018
rect 23992 7978 24480 7984
rect 23690 7868 23696 7928
rect 23756 7868 23762 7928
rect 24220 7706 24280 7978
rect 23170 7646 23176 7706
rect 23236 7646 23242 7706
rect 24214 7646 24220 7706
rect 24280 7646 24286 7706
rect 22674 7542 22680 7602
rect 22740 7542 22746 7602
rect 21956 7494 22444 7500
rect 21956 7460 21968 7494
rect 22432 7460 22444 7494
rect 21956 7454 22444 7460
rect 21660 7374 21674 7410
rect 20690 6834 20696 7346
rect 21668 6892 21674 7374
rect 20650 6822 20696 6834
rect 21664 6834 21674 6892
rect 21708 7374 21720 7410
rect 22680 7410 22740 7542
rect 23176 7500 23236 7646
rect 24220 7500 24280 7646
rect 24718 7602 24778 8068
rect 25732 8068 25746 8100
rect 25780 8100 25786 8644
rect 26752 8644 26812 8776
rect 27046 8728 27534 8734
rect 27046 8694 27058 8728
rect 27522 8694 27534 8728
rect 27046 8688 27534 8694
rect 25780 8068 25792 8100
rect 25010 8018 25498 8024
rect 25010 7984 25022 8018
rect 25486 7984 25498 8018
rect 25010 7978 25498 7984
rect 25210 7706 25270 7978
rect 25732 7928 25792 8068
rect 26752 8068 26764 8644
rect 26798 8068 26812 8644
rect 27768 8644 27828 9300
rect 28788 9300 28800 9334
rect 28834 9836 28846 9876
rect 29804 9876 29864 10016
rect 30310 9966 30370 10080
rect 31326 9966 31386 10080
rect 31836 10016 31842 10076
rect 31902 10016 31908 10076
rect 30100 9960 30588 9966
rect 30100 9926 30112 9960
rect 30576 9926 30588 9960
rect 30100 9920 30588 9926
rect 31118 9960 31606 9966
rect 31118 9926 31130 9960
rect 31594 9926 31606 9960
rect 31118 9920 31606 9926
rect 28834 9334 28840 9836
rect 29804 9834 29818 9876
rect 28834 9300 28848 9334
rect 28064 9250 28552 9256
rect 28064 9216 28076 9250
rect 28540 9216 28552 9250
rect 28064 9210 28552 9216
rect 28264 8940 28324 9210
rect 28258 8880 28264 8940
rect 28324 8880 28330 8940
rect 28264 8734 28324 8880
rect 28064 8728 28552 8734
rect 28064 8694 28076 8728
rect 28540 8694 28552 8728
rect 28064 8688 28552 8694
rect 27768 8604 27782 8644
rect 27776 8100 27782 8604
rect 26028 8018 26516 8024
rect 26028 7984 26040 8018
rect 26504 7984 26516 8018
rect 26028 7978 26516 7984
rect 25726 7868 25732 7928
rect 25792 7868 25798 7928
rect 26228 7706 26288 7978
rect 25204 7646 25210 7706
rect 25270 7646 25276 7706
rect 26222 7646 26228 7706
rect 26288 7646 26294 7706
rect 24712 7542 24718 7602
rect 24778 7542 24784 7602
rect 22974 7494 23462 7500
rect 22974 7460 22986 7494
rect 23450 7460 23462 7494
rect 22974 7454 23462 7460
rect 23992 7494 24480 7500
rect 23992 7460 24004 7494
rect 24468 7460 24480 7494
rect 23992 7454 24480 7460
rect 21708 6892 21714 7374
rect 22680 7372 22692 7410
rect 21708 6834 21724 6892
rect 19920 6784 20408 6790
rect 19920 6750 19932 6784
rect 20396 6750 20408 6784
rect 19920 6744 20408 6750
rect 20938 6784 21426 6790
rect 20938 6750 20950 6784
rect 21414 6750 21426 6784
rect 20938 6744 21426 6750
rect 21664 6700 21724 6834
rect 22686 6834 22692 7372
rect 22726 7372 22740 7410
rect 23704 7410 23750 7422
rect 22726 6834 22732 7372
rect 23704 6884 23710 7410
rect 22686 6822 22732 6834
rect 23696 6834 23710 6884
rect 23744 6884 23750 7410
rect 24718 7410 24778 7542
rect 25210 7500 25270 7646
rect 26752 7602 26812 8068
rect 27770 8068 27782 8100
rect 27816 8604 27828 8644
rect 28788 8644 28848 9300
rect 29812 9300 29818 9834
rect 29852 9834 29864 9876
rect 30830 9876 30876 9888
rect 29852 9300 29858 9834
rect 30830 9358 30836 9876
rect 29812 9288 29858 9300
rect 30822 9300 30836 9358
rect 30870 9358 30876 9876
rect 31842 9876 31902 10016
rect 32344 9966 32404 10444
rect 32860 10406 32920 10534
rect 33878 10534 33890 10592
rect 33924 11082 33936 11110
rect 33924 10592 33930 11082
rect 33924 10534 33938 10592
rect 33154 10484 33642 10490
rect 33154 10450 33166 10484
rect 33630 10450 33642 10484
rect 33154 10444 33642 10450
rect 33878 10424 33938 10534
rect 32854 10346 32860 10406
rect 32920 10346 32926 10406
rect 33872 10364 33878 10424
rect 33938 10364 33944 10424
rect 32860 10128 32920 10346
rect 32860 10068 33934 10128
rect 33984 10076 34044 11252
rect 34472 10234 34478 10294
rect 34538 10234 34544 10294
rect 34222 10130 34228 10190
rect 34288 10130 34294 10190
rect 32136 9960 32624 9966
rect 32136 9926 32148 9960
rect 32612 9926 32624 9960
rect 32136 9920 32624 9926
rect 31842 9834 31854 9876
rect 30870 9300 30882 9358
rect 29294 9256 29354 9258
rect 29082 9250 29570 9256
rect 29082 9216 29094 9250
rect 29558 9216 29570 9250
rect 29082 9210 29570 9216
rect 30100 9250 30588 9256
rect 30100 9216 30112 9250
rect 30576 9216 30588 9250
rect 30100 9210 30588 9216
rect 29294 8940 29354 9210
rect 30316 9162 30376 9210
rect 30310 9102 30316 9162
rect 30376 9102 30382 9162
rect 30448 9106 30454 9166
rect 30514 9106 30520 9166
rect 30454 8940 30514 9106
rect 30822 8940 30882 9300
rect 31848 9300 31854 9834
rect 31888 9834 31902 9876
rect 32860 9876 32920 10068
rect 33364 9966 33424 10068
rect 33154 9960 33642 9966
rect 33154 9926 33166 9960
rect 33630 9926 33642 9960
rect 33154 9920 33642 9926
rect 32860 9842 32872 9876
rect 31888 9300 31894 9834
rect 32866 9340 32872 9842
rect 31848 9288 31894 9300
rect 32860 9300 32872 9340
rect 32906 9842 32920 9876
rect 33874 9876 33934 10068
rect 33978 10016 33984 10076
rect 34044 10016 34050 10076
rect 33874 9852 33890 9876
rect 32906 9340 32912 9842
rect 32906 9300 32920 9340
rect 31118 9250 31606 9256
rect 31118 9216 31130 9250
rect 31594 9216 31606 9250
rect 31118 9210 31606 9216
rect 32136 9250 32624 9256
rect 32136 9216 32148 9250
rect 32612 9216 32624 9250
rect 32136 9210 32624 9216
rect 32342 9166 32402 9210
rect 31330 9106 31336 9166
rect 31396 9106 31402 9166
rect 32336 9106 32342 9166
rect 32402 9106 32408 9166
rect 32860 9162 32920 9300
rect 33884 9300 33890 9852
rect 33924 9852 33934 9876
rect 33924 9300 33930 9852
rect 33884 9288 33930 9300
rect 33154 9250 33642 9256
rect 33154 9216 33166 9250
rect 33630 9216 33642 9250
rect 33154 9210 33642 9216
rect 29288 8880 29294 8940
rect 29354 8880 29360 8940
rect 30448 8880 30454 8940
rect 30514 8880 30520 8940
rect 30816 8880 30822 8940
rect 30882 8880 30888 8940
rect 29294 8734 29354 8880
rect 30454 8734 30514 8880
rect 30822 8836 30882 8880
rect 30816 8776 30822 8836
rect 30882 8776 30888 8836
rect 31336 8734 31396 9106
rect 32854 9102 32860 9162
rect 32920 9102 32926 9162
rect 32854 8974 32860 9034
rect 32920 8974 32926 9034
rect 31832 8778 31838 8838
rect 31898 8778 31904 8838
rect 29082 8728 29570 8734
rect 29082 8694 29094 8728
rect 29558 8694 29570 8728
rect 29082 8688 29570 8694
rect 30100 8728 30588 8734
rect 30100 8694 30112 8728
rect 30576 8694 30588 8728
rect 30100 8688 30588 8694
rect 31118 8728 31606 8734
rect 31118 8694 31130 8728
rect 31594 8694 31606 8728
rect 31118 8688 31606 8694
rect 31336 8686 31396 8688
rect 27816 8100 27822 8604
rect 28788 8598 28800 8644
rect 28794 8112 28800 8598
rect 27816 8068 27830 8100
rect 27046 8018 27534 8024
rect 27046 7984 27058 8018
rect 27522 7984 27534 8018
rect 27046 7978 27534 7984
rect 27262 7706 27322 7978
rect 27770 7928 27830 8068
rect 28786 8068 28800 8112
rect 28834 8598 28848 8644
rect 29812 8644 29858 8656
rect 28834 8112 28840 8598
rect 28834 8068 28846 8112
rect 29812 8108 29818 8644
rect 28064 8018 28552 8024
rect 28064 7984 28076 8018
rect 28540 7984 28552 8018
rect 28064 7978 28552 7984
rect 27764 7868 27770 7928
rect 27830 7868 27836 7928
rect 27756 7760 27762 7820
rect 27822 7760 27828 7820
rect 27256 7646 27262 7706
rect 27322 7646 27328 7706
rect 26746 7542 26752 7602
rect 26812 7542 26818 7602
rect 27258 7538 27264 7598
rect 27324 7538 27330 7598
rect 27264 7500 27324 7538
rect 25010 7494 25498 7500
rect 25010 7460 25022 7494
rect 25486 7460 25498 7494
rect 25010 7454 25498 7460
rect 26028 7494 26516 7500
rect 26028 7460 26040 7494
rect 26504 7460 26516 7494
rect 26028 7454 26516 7460
rect 27046 7494 27534 7500
rect 27046 7460 27058 7494
rect 27522 7460 27534 7494
rect 27046 7454 27534 7460
rect 24718 7374 24728 7410
rect 23744 6834 23756 6884
rect 21956 6784 22444 6790
rect 21956 6750 21968 6784
rect 22432 6750 22444 6784
rect 21956 6744 22444 6750
rect 22974 6784 23462 6790
rect 22974 6750 22986 6784
rect 23450 6750 23462 6784
rect 22974 6744 23462 6750
rect 23696 6700 23756 6834
rect 24722 6834 24728 7374
rect 24762 7374 24778 7410
rect 25740 7410 25786 7422
rect 24762 6834 24768 7374
rect 25740 6896 25746 7410
rect 24722 6822 24768 6834
rect 25730 6834 25746 6896
rect 25780 6896 25786 7410
rect 26758 7410 26804 7422
rect 25780 6834 25790 6896
rect 26758 6876 26764 7410
rect 23992 6784 24480 6790
rect 23992 6750 24004 6784
rect 24468 6750 24480 6784
rect 23992 6744 24480 6750
rect 25010 6784 25498 6790
rect 25010 6750 25022 6784
rect 25486 6750 25498 6784
rect 25010 6744 25498 6750
rect 25730 6700 25790 6834
rect 26752 6834 26764 6876
rect 26798 6876 26804 7410
rect 27762 7410 27822 7760
rect 28286 7598 28346 7978
rect 28786 7604 28846 8068
rect 29806 8068 29818 8108
rect 29852 8108 29858 8644
rect 30830 8644 30876 8656
rect 30830 8112 30836 8644
rect 29852 8068 29866 8108
rect 29082 8018 29570 8024
rect 29082 7984 29094 8018
rect 29558 7984 29570 8018
rect 29082 7978 29570 7984
rect 28280 7538 28286 7598
rect 28346 7538 28352 7598
rect 28780 7544 28786 7604
rect 28846 7544 28852 7604
rect 28286 7500 28346 7538
rect 28064 7494 28552 7500
rect 28064 7460 28076 7494
rect 28540 7460 28552 7494
rect 28064 7454 28552 7460
rect 27762 7374 27782 7410
rect 26798 6834 26812 6876
rect 26028 6784 26516 6790
rect 26028 6750 26040 6784
rect 26504 6750 26516 6784
rect 26028 6744 26516 6750
rect 19106 6634 19112 6694
rect 19172 6634 19178 6694
rect 19622 6640 19628 6700
rect 19688 6640 19694 6700
rect 23690 6640 23696 6700
rect 23756 6640 23762 6700
rect 25724 6640 25730 6700
rect 25790 6640 25796 6700
rect 18604 6320 18610 6380
rect 18670 6320 18676 6380
rect 14830 6260 15318 6266
rect 14830 6226 14842 6260
rect 15306 6226 15318 6260
rect 14830 6220 15318 6226
rect 15848 6260 16336 6266
rect 15848 6226 15860 6260
rect 16324 6226 16336 6260
rect 15848 6220 16336 6226
rect 16866 6260 17354 6266
rect 16866 6226 16878 6260
rect 17342 6226 17354 6260
rect 16866 6220 17354 6226
rect 17884 6260 18372 6266
rect 17884 6226 17896 6260
rect 18360 6226 18372 6260
rect 17884 6220 18372 6226
rect 14532 6122 14548 6176
rect 13564 5600 13574 5634
rect 14542 5630 14548 6122
rect 13514 5468 13574 5600
rect 14538 5600 14548 5630
rect 14582 6122 14592 6176
rect 15560 6176 15606 6188
rect 14582 5630 14588 6122
rect 15560 5646 15566 6176
rect 14582 5600 14598 5630
rect 13812 5550 14300 5556
rect 13812 5516 13824 5550
rect 14288 5516 14300 5550
rect 13812 5510 14300 5516
rect 14034 5468 14094 5510
rect 14538 5468 14598 5600
rect 15552 5600 15566 5646
rect 15600 5646 15606 6176
rect 16578 6176 16624 6188
rect 15600 5600 15612 5646
rect 16578 5630 16584 6176
rect 14830 5550 15318 5556
rect 14830 5516 14842 5550
rect 15306 5516 15318 5550
rect 14830 5510 15318 5516
rect 13514 5408 14598 5468
rect 13392 5298 13398 5358
rect 13458 5298 13464 5358
rect 14538 5262 14598 5408
rect 13514 5202 14598 5262
rect 13514 4944 13574 5202
rect 14026 5034 14086 5202
rect 14538 5142 14598 5202
rect 14532 5082 14538 5142
rect 14598 5082 14604 5142
rect 13812 5028 14300 5034
rect 13812 4994 13824 5028
rect 14288 4994 14300 5028
rect 13812 4988 14300 4994
rect 13514 4908 13530 4944
rect 13524 4368 13530 4908
rect 13564 4908 13574 4944
rect 14538 4944 14598 5082
rect 15030 5034 15090 5510
rect 15552 5456 15612 5600
rect 16570 5600 16584 5630
rect 16618 5630 16624 6176
rect 17596 6176 17642 6188
rect 17596 5642 17602 6176
rect 16618 5600 16630 5630
rect 15848 5550 16336 5556
rect 15848 5516 15860 5550
rect 16324 5516 16336 5550
rect 15848 5510 16336 5516
rect 15546 5396 15552 5456
rect 15612 5396 15618 5456
rect 15550 5202 15556 5262
rect 15616 5202 15622 5262
rect 14830 5028 15318 5034
rect 14830 4994 14842 5028
rect 15306 4994 15318 5028
rect 14830 4988 15318 4994
rect 13564 4368 13570 4908
rect 14538 4904 14548 4944
rect 13524 4356 13570 4368
rect 14542 4368 14548 4904
rect 14582 4904 14598 4944
rect 15556 4944 15616 5202
rect 16050 5198 16110 5510
rect 16570 5358 16630 5600
rect 17588 5600 17602 5642
rect 17636 5642 17642 6176
rect 18610 6176 18670 6320
rect 19112 6266 19172 6634
rect 18902 6260 19390 6266
rect 18902 6226 18914 6260
rect 19378 6226 19390 6260
rect 18902 6220 19390 6226
rect 18610 6146 18620 6176
rect 18614 5664 18620 6146
rect 17636 5600 17648 5642
rect 16866 5550 17354 5556
rect 16866 5516 16878 5550
rect 17342 5516 17354 5550
rect 16866 5510 17354 5516
rect 16564 5298 16570 5358
rect 16630 5298 16636 5358
rect 17084 5198 17144 5510
rect 17588 5456 17648 5600
rect 18606 5600 18620 5664
rect 18654 6146 18670 6176
rect 19628 6176 19688 6640
rect 21664 6634 21724 6640
rect 22674 6530 22680 6590
rect 22740 6530 22746 6590
rect 24710 6530 24716 6590
rect 24776 6530 24782 6590
rect 21656 6418 21662 6478
rect 21722 6418 21728 6478
rect 20640 6320 20646 6380
rect 20706 6320 20712 6380
rect 19920 6260 20408 6266
rect 19920 6226 19932 6260
rect 20396 6226 20408 6260
rect 19920 6220 20408 6226
rect 18654 5664 18660 6146
rect 19628 6134 19638 6176
rect 18654 5600 18666 5664
rect 19632 5640 19638 6134
rect 17884 5550 18372 5556
rect 17884 5516 17896 5550
rect 18360 5516 18372 5550
rect 17884 5510 18372 5516
rect 17582 5396 17588 5456
rect 17648 5396 17654 5456
rect 18094 5358 18154 5510
rect 18088 5298 18094 5358
rect 18154 5298 18160 5358
rect 17586 5202 17592 5262
rect 17652 5202 17658 5262
rect 16050 5138 17144 5198
rect 16050 5034 16110 5138
rect 17084 5034 17144 5138
rect 15848 5028 16336 5034
rect 15848 4994 15860 5028
rect 16324 4994 16336 5028
rect 15848 4988 16336 4994
rect 16866 5028 17354 5034
rect 16866 4994 16878 5028
rect 17342 4994 17354 5028
rect 16866 4988 17354 4994
rect 14582 4368 14588 4904
rect 15556 4900 15566 4944
rect 14542 4356 14588 4368
rect 15560 4368 15566 4900
rect 15600 4900 15616 4944
rect 16578 4944 16624 4956
rect 15600 4368 15606 4900
rect 16578 4410 16584 4944
rect 15560 4356 15606 4368
rect 16570 4368 16584 4410
rect 16618 4410 16624 4944
rect 17592 4944 17652 5202
rect 18094 5034 18154 5298
rect 18606 5142 18666 5600
rect 19626 5600 19638 5640
rect 19672 6134 19688 6176
rect 20646 6176 20706 6320
rect 20938 6260 21426 6266
rect 20938 6226 20950 6260
rect 21414 6226 21426 6260
rect 20938 6220 21426 6226
rect 20646 6140 20656 6176
rect 19672 5640 19678 6134
rect 19672 5600 19686 5640
rect 20650 5634 20656 6140
rect 18902 5550 19390 5556
rect 18902 5516 18914 5550
rect 19378 5516 19390 5550
rect 18902 5510 19390 5516
rect 19116 5358 19176 5510
rect 19626 5456 19686 5600
rect 20640 5600 20656 5634
rect 20690 6140 20706 6176
rect 21662 6176 21722 6418
rect 21956 6260 22444 6266
rect 21956 6226 21968 6260
rect 22432 6226 22444 6260
rect 21956 6220 22444 6226
rect 21662 6150 21674 6176
rect 20690 5634 20696 6140
rect 21668 5656 21674 6150
rect 20690 5600 20700 5634
rect 19920 5550 20408 5556
rect 19920 5516 19932 5550
rect 20396 5516 20408 5550
rect 19920 5510 20408 5516
rect 19620 5396 19626 5456
rect 19686 5396 19692 5456
rect 20140 5364 20200 5510
rect 18600 5082 18606 5142
rect 18666 5082 18672 5142
rect 17884 5028 18372 5034
rect 17884 4994 17896 5028
rect 18360 4994 18372 5028
rect 17884 4988 18372 4994
rect 17592 4892 17602 4944
rect 16618 4368 16630 4410
rect 13812 4318 14300 4324
rect 13812 4284 13824 4318
rect 14288 4284 14300 4318
rect 13812 4278 14300 4284
rect 14830 4318 15318 4324
rect 14830 4284 14842 4318
rect 15306 4284 15318 4318
rect 14830 4278 15318 4284
rect 15848 4318 16336 4324
rect 15848 4284 15860 4318
rect 16324 4284 16336 4318
rect 15848 4278 16336 4284
rect 13280 4166 13286 4226
rect 13346 4166 13352 4226
rect 16570 4100 16630 4368
rect 17596 4368 17602 4892
rect 17636 4892 17652 4944
rect 18606 4944 18666 5082
rect 19116 5034 19176 5298
rect 20138 5358 20200 5364
rect 20198 5298 20200 5358
rect 20138 5292 20200 5298
rect 19614 5202 19620 5262
rect 19680 5202 19686 5262
rect 18902 5028 19390 5034
rect 18902 4994 18914 5028
rect 19378 4994 19390 5028
rect 18902 4988 19390 4994
rect 18606 4904 18620 4944
rect 17636 4368 17642 4892
rect 18614 4422 18620 4904
rect 17596 4356 17642 4368
rect 18608 4368 18620 4422
rect 18654 4904 18666 4944
rect 19620 4944 19680 5202
rect 20140 5034 20200 5292
rect 20640 5142 20700 5600
rect 21658 5600 21674 5656
rect 21708 6150 21722 6176
rect 22680 6176 22740 6530
rect 22974 6260 23462 6266
rect 22974 6226 22986 6260
rect 23450 6226 23462 6260
rect 22974 6220 23462 6226
rect 23992 6260 24480 6266
rect 23992 6226 24004 6260
rect 24468 6226 24480 6260
rect 23992 6220 24480 6226
rect 21708 5656 21714 6150
rect 22680 6144 22692 6176
rect 21708 5600 21718 5656
rect 20938 5550 21426 5556
rect 20938 5516 20950 5550
rect 21414 5516 21426 5550
rect 20938 5510 21426 5516
rect 21142 5358 21202 5510
rect 21488 5476 21548 5482
rect 21658 5476 21718 5600
rect 22686 5600 22692 6144
rect 22726 6144 22740 6176
rect 23704 6176 23750 6188
rect 22726 5600 22732 6144
rect 23704 5670 23710 6176
rect 22686 5588 22732 5600
rect 23700 5600 23710 5670
rect 23744 5670 23750 6176
rect 24716 6176 24776 6530
rect 26258 6492 26318 6744
rect 26752 6702 26812 6834
rect 27776 6834 27782 7374
rect 27816 6834 27822 7410
rect 28786 7410 28846 7544
rect 29264 7500 29324 7978
rect 29806 7928 29866 8068
rect 30820 8068 30836 8112
rect 30870 8112 30876 8644
rect 31838 8644 31898 8778
rect 32136 8728 32624 8734
rect 32136 8694 32148 8728
rect 32612 8694 32624 8728
rect 32136 8688 32624 8694
rect 31838 8594 31854 8644
rect 30870 8068 30880 8112
rect 31848 8096 31854 8594
rect 30100 8018 30588 8024
rect 30100 7984 30112 8018
rect 30576 7984 30588 8018
rect 30100 7978 30588 7984
rect 29800 7868 29806 7928
rect 29866 7868 29872 7928
rect 29796 7760 29802 7820
rect 29862 7760 29868 7820
rect 29082 7494 29570 7500
rect 29082 7460 29094 7494
rect 29558 7460 29570 7494
rect 29082 7454 29570 7460
rect 28786 7316 28800 7410
rect 28794 6876 28800 7316
rect 27776 6822 27822 6834
rect 28786 6834 28800 6876
rect 28834 7316 28846 7410
rect 29802 7410 29862 7760
rect 30288 7646 30294 7706
rect 30354 7646 30360 7706
rect 30294 7500 30354 7646
rect 30820 7604 30880 8068
rect 31844 8068 31854 8096
rect 31888 8594 31898 8644
rect 32860 8644 32920 8974
rect 33154 8728 33642 8734
rect 33154 8694 33166 8728
rect 33630 8694 33642 8728
rect 33154 8688 33642 8694
rect 31888 8096 31894 8594
rect 32860 8592 32872 8644
rect 32866 8096 32872 8592
rect 31888 8068 31904 8096
rect 31118 8018 31606 8024
rect 31118 7984 31130 8018
rect 31594 7984 31606 8018
rect 31118 7978 31606 7984
rect 31844 7928 31904 8068
rect 32860 8068 32872 8096
rect 32906 8592 32920 8644
rect 33884 8644 33930 8656
rect 32906 8096 32912 8592
rect 33884 8102 33890 8644
rect 32906 8068 32920 8096
rect 32136 8018 32624 8024
rect 32136 7984 32148 8018
rect 32612 7984 32624 8018
rect 32136 7978 32624 7984
rect 31838 7868 31844 7928
rect 31904 7868 31910 7928
rect 31834 7760 31840 7820
rect 31900 7760 31906 7820
rect 31326 7646 31332 7706
rect 31392 7646 31398 7706
rect 30814 7544 30820 7604
rect 30880 7544 30886 7604
rect 31332 7500 31392 7646
rect 30100 7494 30588 7500
rect 30100 7460 30112 7494
rect 30576 7460 30588 7494
rect 30100 7454 30588 7460
rect 31118 7494 31606 7500
rect 31118 7460 31130 7494
rect 31594 7460 31606 7494
rect 31118 7454 31606 7460
rect 29802 7344 29818 7410
rect 28834 6876 28840 7316
rect 28834 6834 28846 6876
rect 27046 6784 27534 6790
rect 27046 6750 27058 6784
rect 27522 6750 27534 6784
rect 27046 6744 27534 6750
rect 28064 6784 28552 6790
rect 28064 6750 28076 6784
rect 28540 6750 28552 6784
rect 28064 6744 28552 6750
rect 26746 6642 26752 6702
rect 26812 6642 26818 6702
rect 27100 6642 27106 6702
rect 27166 6642 27172 6702
rect 26742 6530 26748 6590
rect 26808 6530 26814 6590
rect 26252 6432 26258 6492
rect 26318 6432 26324 6492
rect 25010 6260 25498 6266
rect 25010 6226 25022 6260
rect 25486 6226 25498 6260
rect 25010 6220 25498 6226
rect 26028 6260 26516 6266
rect 26028 6226 26040 6260
rect 26504 6226 26516 6260
rect 26028 6220 26516 6226
rect 24716 6138 24728 6176
rect 23744 5600 23760 5670
rect 21956 5550 22444 5556
rect 21956 5516 21968 5550
rect 22432 5516 22444 5550
rect 21956 5510 22444 5516
rect 22974 5550 23462 5556
rect 22974 5516 22986 5550
rect 23450 5516 23462 5550
rect 22974 5510 23462 5516
rect 21652 5416 21658 5476
rect 21718 5416 21724 5476
rect 21136 5298 21142 5358
rect 21202 5298 21208 5358
rect 20634 5082 20640 5142
rect 20700 5082 20706 5142
rect 19920 5028 20408 5034
rect 19920 4994 19932 5028
rect 20396 4994 20408 5028
rect 19920 4988 20408 4994
rect 18654 4422 18660 4904
rect 19620 4884 19638 4944
rect 18654 4368 18668 4422
rect 16866 4318 17354 4324
rect 16866 4284 16878 4318
rect 17342 4284 17354 4318
rect 16866 4278 17354 4284
rect 17884 4318 18372 4324
rect 17884 4284 17896 4318
rect 18360 4284 18372 4318
rect 17884 4278 18372 4284
rect 17090 4112 17150 4278
rect 13174 4040 13180 4100
rect 13240 4040 13246 4100
rect 16564 4040 16570 4100
rect 16630 4040 16636 4100
rect 17084 4052 17090 4112
rect 17150 4052 17156 4112
rect 15546 3930 15552 3990
rect 15612 3930 15618 3990
rect 17582 3930 17588 3990
rect 17648 3930 17654 3990
rect 13812 3794 14300 3800
rect 13812 3760 13824 3794
rect 14288 3760 14300 3794
rect 13812 3754 14300 3760
rect 14830 3794 15318 3800
rect 14830 3760 14842 3794
rect 15306 3760 15318 3794
rect 14830 3754 15318 3760
rect 13524 3710 13570 3722
rect 13524 3160 13530 3710
rect 13518 3134 13530 3160
rect 13564 3160 13570 3710
rect 14542 3710 14588 3722
rect 14542 3188 14548 3710
rect 13564 3134 13578 3160
rect 13518 2996 13578 3134
rect 14530 3134 14548 3188
rect 14582 3188 14588 3710
rect 15552 3710 15612 3930
rect 17200 3836 17206 3896
rect 17266 3836 17272 3896
rect 17206 3800 17266 3836
rect 15848 3794 16336 3800
rect 15848 3760 15860 3794
rect 16324 3760 16336 3794
rect 15848 3754 16336 3760
rect 16866 3794 17354 3800
rect 16866 3760 16878 3794
rect 17342 3760 17354 3794
rect 16866 3754 17354 3760
rect 15552 3650 15566 3710
rect 14582 3134 14590 3188
rect 13812 3084 14300 3090
rect 13812 3050 13824 3084
rect 14288 3050 14300 3084
rect 13812 3044 14300 3050
rect 14032 2996 14092 3044
rect 14530 2996 14590 3134
rect 15560 3134 15566 3650
rect 15600 3650 15612 3710
rect 16578 3710 16624 3722
rect 15600 3134 15606 3650
rect 16578 3178 16584 3710
rect 15560 3122 15606 3134
rect 16572 3134 16584 3178
rect 16618 3178 16624 3710
rect 17588 3710 17648 3930
rect 18090 3896 18150 4278
rect 18608 3990 18668 4368
rect 19632 4368 19638 4884
rect 19672 4884 19680 4944
rect 20640 4944 20700 5082
rect 21142 5034 21202 5298
rect 21488 5262 21548 5416
rect 21482 5202 21488 5262
rect 21548 5202 21554 5262
rect 21658 5208 21664 5268
rect 21724 5208 21730 5268
rect 20938 5028 21426 5034
rect 20938 4994 20950 5028
rect 21414 4994 21426 5028
rect 20938 4988 21426 4994
rect 20640 4904 20656 4944
rect 19672 4368 19678 4884
rect 20650 4434 20656 4904
rect 19632 4356 19678 4368
rect 20644 4368 20656 4434
rect 20690 4904 20700 4944
rect 21664 4944 21724 5208
rect 22180 5206 22240 5510
rect 23194 5370 23254 5510
rect 23700 5476 23760 5600
rect 24722 5600 24728 6138
rect 24762 6138 24776 6176
rect 25740 6176 25786 6188
rect 24762 5600 24768 6138
rect 25740 5670 25746 6176
rect 24722 5588 24768 5600
rect 25732 5600 25746 5670
rect 25780 5670 25786 6176
rect 26748 6176 26808 6530
rect 27106 6384 27166 6642
rect 27296 6492 27356 6744
rect 28272 6492 28332 6744
rect 27290 6432 27296 6492
rect 27356 6432 27362 6492
rect 28266 6432 28272 6492
rect 28332 6432 28338 6492
rect 28786 6380 28846 6834
rect 29812 6834 29818 7344
rect 29852 7344 29862 7410
rect 30830 7410 30876 7422
rect 29852 6834 29858 7344
rect 30830 6878 30836 7410
rect 29812 6822 29858 6834
rect 30824 6834 30836 6878
rect 30870 6878 30876 7410
rect 31840 7410 31900 7760
rect 32358 7706 32418 7978
rect 32860 7886 32920 8068
rect 33874 8068 33890 8102
rect 33924 8102 33930 8644
rect 33924 8068 33934 8102
rect 33154 8018 33642 8024
rect 33154 7984 33166 8018
rect 33630 7984 33642 8018
rect 33154 7978 33642 7984
rect 33368 7886 33428 7978
rect 33874 7886 33934 8068
rect 32860 7826 33934 7886
rect 32352 7646 32358 7706
rect 32418 7646 32424 7706
rect 32856 7544 32862 7604
rect 32922 7544 32928 7604
rect 32136 7494 32624 7500
rect 32136 7460 32148 7494
rect 32612 7460 32624 7494
rect 32136 7454 32624 7460
rect 31840 7358 31854 7410
rect 31848 6884 31854 7358
rect 30870 6834 30884 6878
rect 29082 6784 29570 6790
rect 29082 6750 29094 6784
rect 29558 6750 29570 6784
rect 29082 6744 29570 6750
rect 30100 6784 30588 6790
rect 30100 6750 30112 6784
rect 30576 6750 30588 6784
rect 30100 6744 30588 6750
rect 29288 6492 29348 6744
rect 30824 6702 30884 6834
rect 31842 6834 31854 6884
rect 31888 7358 31900 7410
rect 32862 7410 32922 7544
rect 33154 7494 33642 7500
rect 33154 7460 33166 7494
rect 33630 7460 33642 7494
rect 33154 7454 33642 7460
rect 32862 7376 32872 7410
rect 31888 6884 31894 7358
rect 31888 6834 31902 6884
rect 32866 6878 32872 7376
rect 31118 6784 31606 6790
rect 31118 6750 31130 6784
rect 31594 6750 31606 6784
rect 31118 6744 31606 6750
rect 30818 6642 30824 6702
rect 30884 6642 30890 6702
rect 29282 6432 29288 6492
rect 29348 6432 29354 6492
rect 31308 6432 31314 6492
rect 31374 6432 31380 6492
rect 27106 6318 27166 6324
rect 28780 6320 28786 6380
rect 28846 6320 28852 6380
rect 30816 6320 30822 6380
rect 30882 6320 30888 6380
rect 27046 6260 27534 6266
rect 27046 6226 27058 6260
rect 27522 6226 27534 6260
rect 27046 6220 27534 6226
rect 28064 6260 28552 6266
rect 28064 6226 28076 6260
rect 28540 6226 28552 6260
rect 28064 6220 28552 6226
rect 26748 6134 26764 6176
rect 25780 5600 25792 5670
rect 23992 5550 24480 5556
rect 23992 5516 24004 5550
rect 24468 5516 24480 5550
rect 23992 5510 24480 5516
rect 25010 5550 25498 5556
rect 25010 5516 25022 5550
rect 25486 5516 25498 5550
rect 25010 5510 25498 5516
rect 23694 5416 23700 5476
rect 23760 5416 23766 5476
rect 24216 5370 24276 5510
rect 25230 5370 25290 5510
rect 25732 5476 25792 5600
rect 26758 5600 26764 6134
rect 26798 6134 26808 6176
rect 27776 6176 27822 6188
rect 26798 5600 26804 6134
rect 27776 5636 27782 6176
rect 26758 5588 26804 5600
rect 27772 5600 27782 5636
rect 27816 5636 27822 6176
rect 28786 6176 28846 6320
rect 29082 6260 29570 6266
rect 29082 6226 29094 6260
rect 29558 6226 29570 6260
rect 29082 6220 29570 6226
rect 30100 6260 30588 6266
rect 30100 6226 30112 6260
rect 30576 6226 30588 6260
rect 30100 6220 30588 6226
rect 28786 6138 28800 6176
rect 28794 5652 28800 6138
rect 27816 5600 27832 5636
rect 26028 5550 26516 5556
rect 26028 5516 26040 5550
rect 26504 5516 26516 5550
rect 26028 5510 26516 5516
rect 27046 5550 27534 5556
rect 27046 5516 27058 5550
rect 27522 5516 27534 5550
rect 27046 5510 27534 5516
rect 25726 5416 25732 5476
rect 25792 5416 25798 5476
rect 26232 5470 26292 5510
rect 27258 5470 27318 5510
rect 27772 5476 27832 5600
rect 28790 5600 28800 5652
rect 28834 6138 28846 6176
rect 29812 6176 29858 6188
rect 28834 5652 28840 6138
rect 28834 5600 28850 5652
rect 29812 5644 29818 6176
rect 28064 5550 28552 5556
rect 28064 5516 28076 5550
rect 28540 5516 28552 5550
rect 28064 5510 28552 5516
rect 26232 5410 27318 5470
rect 27766 5416 27772 5476
rect 27832 5416 27838 5476
rect 26232 5370 26292 5410
rect 23194 5310 26292 5370
rect 26744 5318 26750 5378
rect 26810 5318 26816 5378
rect 23194 5206 23254 5310
rect 23686 5208 23692 5268
rect 23752 5208 23758 5268
rect 22180 5146 23254 5206
rect 22180 5034 22240 5146
rect 23194 5034 23254 5146
rect 21956 5028 22444 5034
rect 21956 4994 21968 5028
rect 22432 4994 22444 5028
rect 21956 4988 22444 4994
rect 22974 5028 23462 5034
rect 22974 4994 22986 5028
rect 23450 4994 23462 5028
rect 22974 4988 23462 4994
rect 20690 4434 20696 4904
rect 21664 4900 21674 4944
rect 20690 4368 20704 4434
rect 18902 4318 19390 4324
rect 18902 4284 18914 4318
rect 19378 4284 19390 4318
rect 18902 4278 19390 4284
rect 19920 4318 20408 4324
rect 19920 4284 19932 4318
rect 20396 4284 20408 4318
rect 19920 4278 20408 4284
rect 18602 3930 18608 3990
rect 18668 3930 18674 3990
rect 19112 3896 19172 4278
rect 20644 3990 20704 4368
rect 21668 4368 21674 4900
rect 21708 4900 21724 4944
rect 22686 4944 22732 4956
rect 21708 4368 21714 4900
rect 22686 4420 22692 4944
rect 21668 4356 21714 4368
rect 22674 4368 22692 4420
rect 22726 4420 22732 4944
rect 23692 4944 23752 5208
rect 24216 5034 24276 5310
rect 25230 5034 25290 5310
rect 25730 5208 25736 5268
rect 25796 5208 25802 5268
rect 23992 5028 24480 5034
rect 23992 4994 24004 5028
rect 24468 4994 24480 5028
rect 23992 4988 24480 4994
rect 25010 5028 25498 5034
rect 25010 4994 25022 5028
rect 25486 4994 25498 5028
rect 25010 4988 25498 4994
rect 23692 4900 23710 4944
rect 22726 4368 22734 4420
rect 20938 4318 21426 4324
rect 20938 4284 20950 4318
rect 21414 4284 21426 4318
rect 20938 4278 21426 4284
rect 21956 4318 22444 4324
rect 21956 4284 21968 4318
rect 22432 4284 22444 4318
rect 21956 4278 22444 4284
rect 19618 3930 19624 3990
rect 19684 3930 19690 3990
rect 20638 3930 20644 3990
rect 20704 3930 20710 3990
rect 18084 3836 18090 3896
rect 18150 3836 18156 3896
rect 19106 3836 19112 3896
rect 19172 3836 19178 3896
rect 18090 3800 18150 3836
rect 19112 3800 19172 3836
rect 17884 3794 18372 3800
rect 17884 3760 17896 3794
rect 18360 3760 18372 3794
rect 17884 3754 18372 3760
rect 18902 3794 19390 3800
rect 18902 3760 18914 3794
rect 19378 3760 19390 3794
rect 18902 3754 19390 3760
rect 17588 3660 17602 3710
rect 17596 3196 17602 3660
rect 16618 3134 16632 3178
rect 14830 3084 15318 3090
rect 14830 3050 14842 3084
rect 15306 3050 15318 3084
rect 14830 3044 15318 3050
rect 15848 3084 16336 3090
rect 15848 3050 15860 3084
rect 16324 3050 16336 3084
rect 15848 3044 16336 3050
rect 13512 2936 13518 2996
rect 13578 2936 13584 2996
rect 14026 2936 14032 2996
rect 14092 2936 14098 2996
rect 14524 2936 14530 2996
rect 14590 2936 14596 2996
rect 15046 2778 15106 3044
rect 16068 2778 16128 3044
rect 16572 2996 16632 3134
rect 17586 3134 17602 3196
rect 17636 3660 17648 3710
rect 18614 3710 18660 3722
rect 17636 3196 17642 3660
rect 17636 3134 17646 3196
rect 18614 3174 18620 3710
rect 16866 3084 17354 3090
rect 16866 3050 16878 3084
rect 17342 3050 17354 3084
rect 16866 3044 17354 3050
rect 16566 2936 16572 2996
rect 16632 2936 16638 2996
rect 17080 2884 17140 3044
rect 17074 2824 17080 2884
rect 17140 2824 17146 2884
rect 13054 2718 13060 2778
rect 13120 2718 13126 2778
rect 15040 2718 15046 2778
rect 15106 2718 15112 2778
rect 16062 2718 16068 2778
rect 16128 2718 16134 2778
rect 17586 2674 17646 3134
rect 18604 3134 18620 3174
rect 18654 3174 18660 3710
rect 19624 3710 19684 3930
rect 21154 3896 21214 4278
rect 22170 4112 22230 4278
rect 22674 4226 22734 4368
rect 23704 4368 23710 4900
rect 23744 4900 23752 4944
rect 24722 4944 24768 4956
rect 23744 4368 23750 4900
rect 24722 4420 24728 4944
rect 23704 4356 23750 4368
rect 24716 4368 24728 4420
rect 24762 4420 24768 4944
rect 25736 4944 25796 5208
rect 26232 5034 26292 5310
rect 26028 5028 26516 5034
rect 26028 4994 26040 5028
rect 26504 4994 26516 5028
rect 26028 4988 26516 4994
rect 25736 4896 25746 4944
rect 24762 4368 24776 4420
rect 22974 4318 23462 4324
rect 22974 4284 22986 4318
rect 23450 4284 23462 4318
rect 22974 4278 23462 4284
rect 23992 4318 24480 4324
rect 23992 4284 24004 4318
rect 24468 4284 24480 4318
rect 23992 4278 24480 4284
rect 24716 4226 24776 4368
rect 25740 4368 25746 4896
rect 25780 4896 25796 4944
rect 26750 4944 26810 5318
rect 27258 5034 27318 5410
rect 27758 5208 27764 5268
rect 27824 5208 27830 5268
rect 27046 5028 27534 5034
rect 27046 4994 27058 5028
rect 27522 4994 27534 5028
rect 27046 4988 27534 4994
rect 26750 4908 26764 4944
rect 25780 4368 25786 4896
rect 26758 4412 26764 4908
rect 25740 4356 25786 4368
rect 26752 4368 26764 4412
rect 26798 4908 26810 4944
rect 27764 4944 27824 5208
rect 28278 5034 28338 5510
rect 28790 5142 28850 5600
rect 29802 5600 29818 5644
rect 29852 5644 29858 6176
rect 30822 6176 30882 6320
rect 31314 6266 31374 6432
rect 31118 6260 31606 6266
rect 31118 6226 31130 6260
rect 31594 6226 31606 6260
rect 31118 6220 31606 6226
rect 30822 6118 30836 6176
rect 29852 5600 29862 5644
rect 30830 5640 30836 6118
rect 29082 5550 29570 5556
rect 29082 5516 29094 5550
rect 29558 5516 29570 5550
rect 29082 5510 29570 5516
rect 28784 5082 28790 5142
rect 28850 5082 28856 5142
rect 28064 5028 28552 5034
rect 28064 4994 28076 5028
rect 28540 4994 28552 5028
rect 28064 4988 28552 4994
rect 26798 4412 26804 4908
rect 27764 4896 27782 4944
rect 26798 4368 26812 4412
rect 25010 4318 25498 4324
rect 25010 4284 25022 4318
rect 25486 4284 25498 4318
rect 25010 4278 25498 4284
rect 26028 4318 26516 4324
rect 26028 4284 26040 4318
rect 26504 4284 26516 4318
rect 26028 4278 26516 4284
rect 26752 4226 26812 4368
rect 27776 4368 27782 4896
rect 27816 4896 27824 4944
rect 28790 4944 28850 5082
rect 29294 5034 29354 5510
rect 29802 5268 29862 5600
rect 30820 5600 30836 5640
rect 30870 6118 30882 6176
rect 31842 6176 31902 6834
rect 32858 6834 32872 6878
rect 32906 7376 32922 7410
rect 33884 7410 33930 7422
rect 32906 6878 32912 7376
rect 32906 6834 32918 6878
rect 33884 6864 33890 7410
rect 32136 6784 32624 6790
rect 32136 6750 32148 6784
rect 32612 6750 32624 6784
rect 32136 6744 32624 6750
rect 32344 6492 32404 6744
rect 32858 6652 32918 6834
rect 33874 6834 33890 6864
rect 33924 6864 33930 7410
rect 33924 6834 33934 6864
rect 33154 6784 33642 6790
rect 33154 6750 33166 6784
rect 33630 6750 33642 6784
rect 33154 6744 33642 6750
rect 33364 6652 33424 6744
rect 33874 6652 33934 6834
rect 32858 6592 33934 6652
rect 32338 6432 32344 6492
rect 32404 6432 32410 6492
rect 32858 6380 32918 6592
rect 32852 6320 32858 6380
rect 32918 6320 32924 6380
rect 32136 6260 32624 6266
rect 32136 6226 32148 6260
rect 32612 6226 32624 6260
rect 32136 6220 32624 6226
rect 33154 6260 33642 6266
rect 33154 6226 33166 6260
rect 33630 6226 33642 6260
rect 33154 6220 33642 6226
rect 31842 6134 31854 6176
rect 30870 5640 30876 6118
rect 31848 5654 31854 6134
rect 30870 5600 30880 5640
rect 30100 5550 30588 5556
rect 30100 5516 30112 5550
rect 30576 5516 30588 5550
rect 30100 5510 30588 5516
rect 29796 5208 29802 5268
rect 29862 5208 29868 5268
rect 30328 5034 30388 5510
rect 30820 5142 30880 5600
rect 31842 5600 31854 5654
rect 31888 6134 31902 6176
rect 32866 6176 32912 6188
rect 31888 5654 31894 6134
rect 31888 5600 31902 5654
rect 32866 5646 32872 6176
rect 31118 5550 31606 5556
rect 31118 5516 31130 5550
rect 31594 5516 31606 5550
rect 31118 5510 31606 5516
rect 31346 5144 31406 5510
rect 31842 5268 31902 5600
rect 32856 5600 32872 5646
rect 32906 5646 32912 6176
rect 33884 6176 33930 6188
rect 32906 5600 32916 5646
rect 33884 5628 33890 6176
rect 32136 5550 32624 5556
rect 32136 5516 32148 5550
rect 32612 5516 32624 5550
rect 32136 5510 32624 5516
rect 32360 5272 32420 5510
rect 32856 5474 32916 5600
rect 33876 5600 33890 5628
rect 33924 5628 33930 6176
rect 33924 5600 33936 5628
rect 33154 5550 33642 5556
rect 33154 5516 33166 5550
rect 33630 5516 33642 5550
rect 33154 5510 33642 5516
rect 33362 5476 33422 5510
rect 33876 5476 33936 5600
rect 33362 5474 33936 5476
rect 32856 5414 33936 5474
rect 32856 5378 32916 5414
rect 32850 5318 32856 5378
rect 32916 5318 32922 5378
rect 31836 5208 31842 5268
rect 31902 5208 31908 5268
rect 32354 5212 32360 5272
rect 32420 5212 32426 5272
rect 30814 5082 30820 5142
rect 30880 5082 30886 5142
rect 29082 5028 29570 5034
rect 29082 4994 29094 5028
rect 29558 4994 29570 5028
rect 29082 4988 29570 4994
rect 30100 5028 30588 5034
rect 30100 4994 30112 5028
rect 30576 4994 30588 5028
rect 30100 4988 30588 4994
rect 28790 4898 28800 4944
rect 27816 4368 27822 4896
rect 28794 4428 28800 4898
rect 27776 4356 27822 4368
rect 28788 4368 28800 4428
rect 28834 4898 28850 4944
rect 29812 4944 29858 4956
rect 28834 4428 28840 4898
rect 28834 4368 28848 4428
rect 29812 4412 29818 4944
rect 27046 4318 27534 4324
rect 27046 4284 27058 4318
rect 27522 4284 27534 4318
rect 27046 4278 27534 4284
rect 28064 4318 28552 4324
rect 28064 4284 28076 4318
rect 28540 4284 28552 4318
rect 28064 4278 28552 4284
rect 22668 4166 22674 4226
rect 22734 4166 22740 4226
rect 24710 4166 24716 4226
rect 24776 4166 24782 4226
rect 26746 4166 26752 4226
rect 26812 4166 26818 4226
rect 27258 4116 27318 4278
rect 22164 4052 22170 4112
rect 22230 4052 22236 4112
rect 27252 4056 27258 4116
rect 27318 4056 27324 4116
rect 21656 3930 21662 3990
rect 21722 3930 21728 3990
rect 23686 3930 23692 3990
rect 23752 3930 23758 3990
rect 25724 3930 25730 3990
rect 25790 3930 25796 3990
rect 27760 3930 27766 3990
rect 27826 3930 27832 3990
rect 21148 3836 21154 3896
rect 21214 3836 21220 3896
rect 19920 3794 20408 3800
rect 19920 3760 19932 3794
rect 20396 3760 20408 3794
rect 19920 3754 20408 3760
rect 20938 3794 21426 3800
rect 20938 3760 20950 3794
rect 21414 3760 21426 3794
rect 20938 3754 21426 3760
rect 18654 3134 18664 3174
rect 17884 3084 18372 3090
rect 17884 3050 17896 3084
rect 18360 3050 18372 3084
rect 17884 3044 18372 3050
rect 18092 2884 18152 3044
rect 18604 2996 18664 3134
rect 19624 3134 19638 3710
rect 19672 3134 19684 3710
rect 20650 3710 20696 3722
rect 20650 3174 20656 3710
rect 18902 3084 19390 3090
rect 18902 3050 18914 3084
rect 19378 3050 19390 3084
rect 18902 3044 19390 3050
rect 18598 2936 18604 2996
rect 18664 2936 18670 2996
rect 19106 2884 19166 3044
rect 18086 2824 18092 2884
rect 18152 2824 18158 2884
rect 19100 2824 19106 2884
rect 19166 2824 19172 2884
rect 18600 2718 18606 2778
rect 18666 2718 18672 2778
rect 19112 2718 19118 2778
rect 19178 2718 19184 2778
rect 12648 2614 12654 2674
rect 12714 2614 12720 2674
rect 17076 2614 17082 2674
rect 17142 2614 17148 2674
rect 17580 2614 17586 2674
rect 17646 2614 17652 2674
rect 18096 2614 18102 2674
rect 18162 2614 18168 2674
rect 12020 1566 12026 1626
rect 12086 1566 12092 1626
rect 8818 540 8824 600
rect 8884 540 8890 600
rect 10006 540 10012 600
rect 10072 540 10078 600
rect 11202 540 11208 600
rect 11268 540 11274 600
rect 11896 540 11902 600
rect 11962 540 11968 600
rect 12654 110 12714 2614
rect 17082 2566 17142 2614
rect 13812 2560 14300 2566
rect 13812 2526 13824 2560
rect 14288 2526 14300 2560
rect 13812 2520 14300 2526
rect 14830 2560 15318 2566
rect 14830 2526 14842 2560
rect 15306 2526 15318 2560
rect 14830 2520 15318 2526
rect 15848 2560 16336 2566
rect 15848 2526 15860 2560
rect 16324 2526 16336 2560
rect 15848 2520 16336 2526
rect 16866 2560 17354 2566
rect 16866 2526 16878 2560
rect 17342 2526 17354 2560
rect 16866 2520 17354 2526
rect 13524 2476 13570 2488
rect 13524 1926 13530 2476
rect 13518 1900 13530 1926
rect 13564 1926 13570 2476
rect 14542 2476 14588 2488
rect 14542 1928 14548 2476
rect 13564 1900 13578 1926
rect 13518 1444 13578 1900
rect 14530 1900 14548 1928
rect 14582 1928 14588 2476
rect 15560 2476 15606 2488
rect 15560 1932 15566 2476
rect 14582 1900 14590 1928
rect 13812 1850 14300 1856
rect 13812 1816 13824 1850
rect 14288 1816 14300 1850
rect 13812 1810 14300 1816
rect 13512 1384 13518 1444
rect 13578 1384 13584 1444
rect 13518 1244 13578 1384
rect 14016 1334 14076 1810
rect 14530 1542 14590 1900
rect 15548 1900 15566 1932
rect 15600 1932 15606 2476
rect 16578 2476 16624 2488
rect 16578 1940 16584 2476
rect 15600 1900 15608 1932
rect 14830 1850 15318 1856
rect 14830 1816 14842 1850
rect 15306 1816 15318 1850
rect 14830 1810 15318 1816
rect 14524 1482 14530 1542
rect 14590 1482 14596 1542
rect 13812 1328 14300 1334
rect 13812 1294 13824 1328
rect 14288 1294 14300 1328
rect 13812 1288 14300 1294
rect 13518 1188 13530 1244
rect 13524 668 13530 1188
rect 13564 1188 13578 1244
rect 14530 1244 14590 1482
rect 15038 1334 15098 1810
rect 15548 1444 15608 1900
rect 16568 1900 16584 1940
rect 16618 1940 16624 2476
rect 17586 2476 17646 2614
rect 18102 2566 18162 2614
rect 17884 2560 18372 2566
rect 17884 2526 17896 2560
rect 18360 2526 18372 2560
rect 17884 2520 18372 2526
rect 18606 2476 18666 2718
rect 19118 2566 19178 2718
rect 19624 2674 19684 3134
rect 20636 3134 20656 3174
rect 20690 3134 20696 3710
rect 21662 3710 21722 3930
rect 22168 3854 23238 3914
rect 22168 3800 22228 3854
rect 21956 3794 22444 3800
rect 21956 3760 21968 3794
rect 22432 3760 22444 3794
rect 21956 3754 22444 3760
rect 21662 3654 21674 3710
rect 21668 3186 21674 3654
rect 19920 3084 20408 3090
rect 19920 3050 19932 3084
rect 20396 3050 20408 3084
rect 19920 3044 20408 3050
rect 20136 2778 20196 3044
rect 20636 2996 20696 3134
rect 21662 3134 21674 3186
rect 21708 3654 21722 3710
rect 22680 3710 22740 3854
rect 23178 3800 23238 3854
rect 22974 3794 23462 3800
rect 22974 3760 22986 3794
rect 23450 3760 23462 3794
rect 22974 3754 23462 3760
rect 22680 3674 22692 3710
rect 21708 3186 21714 3654
rect 21708 3134 21722 3186
rect 22686 3178 22692 3674
rect 22678 3170 22692 3178
rect 22672 3134 22692 3170
rect 22726 3674 22740 3710
rect 23692 3710 23752 3930
rect 24192 3858 25280 3918
rect 24192 3800 24252 3858
rect 23992 3794 24480 3800
rect 23992 3760 24004 3794
rect 24468 3760 24480 3794
rect 23992 3754 24480 3760
rect 22726 3178 22732 3674
rect 23692 3660 23710 3710
rect 23704 3184 23710 3660
rect 22726 3134 22738 3178
rect 20938 3084 21426 3090
rect 20938 3050 20950 3084
rect 21414 3050 21426 3084
rect 20938 3044 21426 3050
rect 20630 2936 20636 2996
rect 20696 2936 20702 2996
rect 21148 2778 21208 3044
rect 20130 2718 20136 2778
rect 20196 2718 20202 2778
rect 20636 2718 20642 2778
rect 20702 2718 20708 2778
rect 21142 2718 21148 2778
rect 21208 2718 21214 2778
rect 19618 2614 19624 2674
rect 19684 2614 19690 2674
rect 18902 2560 19390 2566
rect 18902 2526 18914 2560
rect 19378 2526 19390 2560
rect 18902 2520 19390 2526
rect 17586 2424 17602 2476
rect 16618 1900 16628 1940
rect 15848 1850 16336 1856
rect 15848 1816 15860 1850
rect 16324 1816 16336 1850
rect 15848 1810 16336 1816
rect 15542 1384 15548 1444
rect 15608 1384 15614 1444
rect 14830 1328 15318 1334
rect 14830 1294 14842 1328
rect 15306 1294 15318 1328
rect 14830 1288 15318 1294
rect 14530 1206 14548 1244
rect 13564 668 13570 1188
rect 14542 718 14548 1206
rect 13524 656 13570 668
rect 14532 668 14548 718
rect 14582 1206 14590 1244
rect 15548 1244 15608 1384
rect 16064 1334 16124 1810
rect 16568 1542 16628 1900
rect 17596 1900 17602 2424
rect 17636 2424 17646 2476
rect 17636 1900 17642 2424
rect 18604 2420 18620 2476
rect 18614 1942 18620 2420
rect 17596 1888 17642 1900
rect 18604 1900 18620 1942
rect 18654 2424 18666 2476
rect 19624 2476 19684 2614
rect 20136 2566 20196 2718
rect 19920 2560 20408 2566
rect 19920 2526 19932 2560
rect 20396 2526 20408 2560
rect 19920 2520 20408 2526
rect 20642 2476 20702 2718
rect 21148 2566 21208 2718
rect 21662 2674 21722 3134
rect 21956 3084 22444 3090
rect 21956 3050 21968 3084
rect 22432 3050 22444 3084
rect 21956 3044 22444 3050
rect 22012 2824 22018 2884
rect 22078 2824 22084 2884
rect 21656 2614 21662 2674
rect 21722 2614 21728 2674
rect 20938 2560 21426 2566
rect 20938 2526 20950 2560
rect 21414 2526 21426 2560
rect 20938 2520 21426 2526
rect 19624 2426 19638 2476
rect 18654 2420 18664 2424
rect 18654 1942 18660 2420
rect 18654 1900 18664 1942
rect 16866 1850 17354 1856
rect 16866 1816 16878 1850
rect 17342 1816 17354 1850
rect 16866 1810 17354 1816
rect 17884 1850 18372 1856
rect 17884 1816 17896 1850
rect 18360 1816 18372 1850
rect 17884 1810 18372 1816
rect 18604 1756 18664 1900
rect 19632 1900 19638 2426
rect 19672 2426 19684 2476
rect 19672 1900 19678 2426
rect 20636 2410 20656 2476
rect 20650 1934 20656 2410
rect 19632 1888 19678 1900
rect 20642 1900 20656 1934
rect 20690 2436 20702 2476
rect 21662 2476 21722 2614
rect 22018 2566 22078 2824
rect 22160 2778 22220 3044
rect 22540 2996 22600 3002
rect 22154 2718 22160 2778
rect 22220 2718 22226 2778
rect 22540 2766 22600 2936
rect 22678 2886 22738 3134
rect 23698 3134 23710 3184
rect 23744 3660 23752 3710
rect 24716 3710 24776 3858
rect 25220 3800 25280 3858
rect 25010 3794 25498 3800
rect 25010 3760 25022 3794
rect 25486 3760 25498 3794
rect 25010 3754 25498 3760
rect 24716 3678 24728 3710
rect 23744 3184 23750 3660
rect 24722 3188 24728 3678
rect 23744 3134 23758 3184
rect 22974 3084 23462 3090
rect 22974 3050 22986 3084
rect 23450 3050 23462 3084
rect 22974 3044 23462 3050
rect 22672 2826 22678 2886
rect 22738 2826 22744 2886
rect 23180 2778 23240 3044
rect 23300 2822 23306 2882
rect 23366 2822 23372 2882
rect 22540 2706 22740 2766
rect 23174 2718 23180 2778
rect 23240 2718 23246 2778
rect 21956 2560 22444 2566
rect 21956 2526 21968 2560
rect 22432 2526 22444 2560
rect 21956 2520 22444 2526
rect 20690 1934 20696 2436
rect 21662 2416 21674 2476
rect 20690 1900 20702 1934
rect 18902 1850 19390 1856
rect 18902 1816 18914 1850
rect 19378 1816 19390 1850
rect 18902 1810 19390 1816
rect 19920 1850 20408 1856
rect 19920 1816 19932 1850
rect 20396 1816 20408 1850
rect 19920 1810 20408 1816
rect 19108 1756 19168 1810
rect 18604 1696 19168 1756
rect 20124 1748 20184 1810
rect 20642 1748 20702 1900
rect 21668 1900 21674 2416
rect 21708 2416 21722 2476
rect 22680 2476 22740 2706
rect 23306 2566 23366 2822
rect 23698 2674 23758 3134
rect 24714 3134 24728 3188
rect 24762 3678 24776 3710
rect 25730 3710 25790 3930
rect 26028 3794 26516 3800
rect 26028 3760 26040 3794
rect 26504 3760 26516 3794
rect 26028 3754 26516 3760
rect 27046 3794 27534 3800
rect 27046 3760 27058 3794
rect 27522 3760 27534 3794
rect 27046 3754 27534 3760
rect 24762 3188 24768 3678
rect 25730 3666 25746 3710
rect 24762 3134 24774 3188
rect 25740 3172 25746 3666
rect 23992 3084 24480 3090
rect 23992 3050 24004 3084
rect 24468 3050 24480 3084
rect 23992 3044 24480 3050
rect 24202 2778 24262 3044
rect 24346 2822 24352 2882
rect 24412 2822 24418 2882
rect 24196 2718 24202 2778
rect 24262 2718 24268 2778
rect 23692 2614 23698 2674
rect 23758 2614 23764 2674
rect 22974 2560 23462 2566
rect 22974 2526 22986 2560
rect 23450 2526 23462 2560
rect 22974 2520 23462 2526
rect 22680 2448 22692 2476
rect 21708 1900 21714 2416
rect 22686 1924 22692 2448
rect 21668 1888 21714 1900
rect 22680 1900 22692 1924
rect 22726 2448 22740 2476
rect 23698 2476 23758 2614
rect 24352 2566 24412 2822
rect 24714 2778 24774 3134
rect 25734 3134 25746 3172
rect 25780 3666 25790 3710
rect 26758 3710 26804 3722
rect 25780 3172 25786 3666
rect 26758 3194 26764 3710
rect 25780 3134 25794 3172
rect 25010 3084 25498 3090
rect 25010 3050 25022 3084
rect 25486 3050 25498 3084
rect 25010 3044 25498 3050
rect 24900 2998 24960 3004
rect 24708 2718 24714 2778
rect 24774 2718 24780 2778
rect 24900 2670 24960 2938
rect 25220 2778 25280 3044
rect 25214 2718 25220 2778
rect 25280 2718 25286 2778
rect 24716 2610 24960 2670
rect 23992 2560 24480 2566
rect 23992 2526 24004 2560
rect 24468 2526 24480 2560
rect 23992 2520 24480 2526
rect 22726 1924 22732 2448
rect 23698 2410 23710 2476
rect 22726 1900 22740 1924
rect 20938 1850 21426 1856
rect 20938 1816 20950 1850
rect 21414 1816 21426 1850
rect 20938 1810 21426 1816
rect 21956 1850 22444 1856
rect 21956 1816 21968 1850
rect 22432 1816 22444 1850
rect 21956 1810 22444 1816
rect 21150 1748 21210 1810
rect 20124 1688 21210 1748
rect 22170 1638 22230 1810
rect 22680 1742 22740 1900
rect 23704 1900 23710 2410
rect 23744 2410 23758 2476
rect 24716 2476 24776 2610
rect 25220 2566 25280 2718
rect 25734 2674 25794 3134
rect 26750 3134 26764 3194
rect 26798 3194 26804 3710
rect 27766 3710 27826 3930
rect 28276 3896 28336 4278
rect 28788 3990 28848 4368
rect 29806 4368 29818 4412
rect 29852 4412 29858 4944
rect 30820 4944 30880 5082
rect 31346 5034 31406 5084
rect 32360 5034 32420 5212
rect 32858 5144 33936 5202
rect 32852 5084 32858 5144
rect 32918 5142 33936 5144
rect 32918 5084 32924 5142
rect 31118 5028 31606 5034
rect 31118 4994 31130 5028
rect 31594 4994 31606 5028
rect 31118 4988 31606 4994
rect 32136 5028 32624 5034
rect 32136 4994 32148 5028
rect 32612 4994 32624 5028
rect 32136 4988 32624 4994
rect 30820 4898 30836 4944
rect 30830 4416 30836 4898
rect 29852 4368 29866 4412
rect 29082 4318 29570 4324
rect 29082 4284 29094 4318
rect 29558 4284 29570 4318
rect 29082 4278 29570 4284
rect 28782 3930 28788 3990
rect 28848 3930 28854 3990
rect 29296 3896 29356 4278
rect 29806 4226 29866 4368
rect 30822 4368 30836 4416
rect 30870 4898 30880 4944
rect 31848 4944 31894 4956
rect 30870 4416 30876 4898
rect 30870 4368 30882 4416
rect 31848 4412 31854 4944
rect 30100 4318 30588 4324
rect 30100 4284 30112 4318
rect 30576 4284 30588 4318
rect 30100 4278 30588 4284
rect 29800 4166 29806 4226
rect 29866 4166 29872 4226
rect 29802 3930 29808 3990
rect 29868 3930 29874 3990
rect 28270 3836 28276 3896
rect 28336 3836 28342 3896
rect 29290 3836 29296 3896
rect 29356 3836 29362 3896
rect 28276 3800 28336 3836
rect 29296 3800 29356 3836
rect 28064 3794 28552 3800
rect 28064 3760 28076 3794
rect 28540 3760 28552 3794
rect 28064 3754 28552 3760
rect 29082 3794 29570 3800
rect 29082 3760 29094 3794
rect 29558 3760 29570 3794
rect 29082 3754 29570 3760
rect 27766 3666 27782 3710
rect 26798 3134 26810 3194
rect 27776 3188 27782 3666
rect 26028 3084 26516 3090
rect 26028 3050 26040 3084
rect 26504 3050 26516 3084
rect 26028 3044 26516 3050
rect 26238 2778 26298 3044
rect 26750 2996 26810 3134
rect 27766 3134 27782 3188
rect 27816 3666 27826 3710
rect 28794 3710 28840 3722
rect 27816 3188 27822 3666
rect 27816 3134 27826 3188
rect 28794 3166 28800 3710
rect 27046 3084 27534 3090
rect 27046 3050 27058 3084
rect 27522 3050 27534 3084
rect 27046 3044 27534 3050
rect 26744 2936 26750 2996
rect 26810 2936 26816 2996
rect 27258 2778 27318 3044
rect 26232 2718 26238 2778
rect 26298 2718 26304 2778
rect 26744 2718 26750 2778
rect 26810 2718 26816 2778
rect 27252 2718 27258 2778
rect 27318 2718 27324 2778
rect 25728 2614 25734 2674
rect 25794 2614 25800 2674
rect 25010 2560 25498 2566
rect 25010 2526 25022 2560
rect 25486 2526 25498 2560
rect 25010 2520 25498 2526
rect 24716 2442 24728 2476
rect 23744 1900 23750 2410
rect 24722 1966 24728 2442
rect 23704 1888 23750 1900
rect 24716 1900 24728 1966
rect 24762 2442 24776 2476
rect 25734 2476 25794 2614
rect 26238 2566 26298 2718
rect 26028 2560 26516 2566
rect 26028 2526 26040 2560
rect 26504 2526 26516 2560
rect 26028 2520 26516 2526
rect 26750 2476 26810 2718
rect 27258 2566 27318 2718
rect 27766 2674 27826 3134
rect 28784 3134 28800 3166
rect 28834 3166 28840 3710
rect 29808 3710 29868 3930
rect 30310 3896 30370 4278
rect 30822 3990 30882 4368
rect 31838 4368 31854 4412
rect 31888 4412 31894 4944
rect 32858 4944 32918 5084
rect 33360 5034 33420 5142
rect 33154 5028 33642 5034
rect 33154 4994 33166 5028
rect 33630 4994 33642 5028
rect 33154 4988 33642 4994
rect 32858 4910 32872 4944
rect 31888 4368 31898 4412
rect 31118 4318 31606 4324
rect 31118 4284 31130 4318
rect 31594 4284 31606 4318
rect 31118 4278 31606 4284
rect 30816 3930 30822 3990
rect 30882 3930 30888 3990
rect 31346 3896 31406 4278
rect 31838 4226 31898 4368
rect 32866 4368 32872 4910
rect 32906 4910 32918 4944
rect 33876 4944 33936 5142
rect 32906 4368 32912 4910
rect 33876 4906 33890 4944
rect 32866 4356 32912 4368
rect 33884 4368 33890 4906
rect 33924 4906 33936 4944
rect 33924 4368 33930 4906
rect 33884 4356 33930 4368
rect 32136 4318 32624 4324
rect 32136 4284 32148 4318
rect 32612 4284 32624 4318
rect 32136 4278 32624 4284
rect 33154 4318 33642 4324
rect 33154 4284 33166 4318
rect 33630 4284 33642 4318
rect 33154 4278 33642 4284
rect 31832 4166 31838 4226
rect 31898 4166 31904 4226
rect 32358 4116 32418 4278
rect 33984 4226 34044 10016
rect 34106 9102 34112 9162
rect 34172 9102 34178 9162
rect 34112 7604 34172 9102
rect 34228 8838 34288 10130
rect 34344 8880 34350 8940
rect 34410 8880 34416 8940
rect 34222 8778 34228 8838
rect 34288 8778 34294 8838
rect 34106 7544 34112 7604
rect 34172 7544 34178 7604
rect 34102 6642 34108 6702
rect 34168 6642 34174 6702
rect 34108 5378 34168 6642
rect 34228 5476 34288 8778
rect 34222 5416 34228 5476
rect 34288 5416 34294 5476
rect 34102 5318 34108 5378
rect 34168 5318 34174 5378
rect 34350 5144 34410 8880
rect 34478 7712 34538 10234
rect 34476 7706 34538 7712
rect 34536 7646 34538 7706
rect 34476 7640 34538 7646
rect 34478 5272 34538 7640
rect 34472 5212 34478 5272
rect 34538 5212 34544 5272
rect 34344 5084 34350 5144
rect 34410 5084 34416 5144
rect 33978 4166 33984 4226
rect 34044 4166 34050 4226
rect 32352 4056 32358 4116
rect 32418 4056 32424 4116
rect 32358 3992 32418 4056
rect 31838 3930 31844 3990
rect 31904 3930 31910 3990
rect 32358 3932 34104 3992
rect 30304 3836 30310 3896
rect 30370 3836 30376 3896
rect 31340 3836 31346 3896
rect 31406 3836 31412 3896
rect 30310 3800 30370 3836
rect 30100 3794 30588 3800
rect 30100 3760 30112 3794
rect 30576 3760 30588 3794
rect 30100 3754 30588 3760
rect 31118 3794 31606 3800
rect 31118 3760 31130 3794
rect 31594 3760 31606 3794
rect 31118 3754 31606 3760
rect 30318 3750 30378 3754
rect 29808 3644 29818 3710
rect 29812 3182 29818 3644
rect 28834 3134 28844 3166
rect 28064 3084 28552 3090
rect 28064 3050 28076 3084
rect 28540 3050 28552 3084
rect 28064 3044 28552 3050
rect 28280 2882 28340 3044
rect 28784 2996 28844 3134
rect 29804 3134 29818 3182
rect 29852 3644 29868 3710
rect 30830 3710 30876 3722
rect 29852 3182 29858 3644
rect 30830 3184 30836 3710
rect 29852 3134 29864 3182
rect 29082 3084 29570 3090
rect 29082 3050 29094 3084
rect 29558 3050 29570 3084
rect 29082 3044 29570 3050
rect 28778 2936 28784 2996
rect 28844 2936 28850 2996
rect 29298 2882 29358 3044
rect 28274 2822 28280 2882
rect 28340 2822 28346 2882
rect 29292 2822 29298 2882
rect 29358 2822 29364 2882
rect 29804 2674 29864 3134
rect 30818 3134 30836 3184
rect 30870 3184 30876 3710
rect 31844 3710 31904 3930
rect 32136 3794 32624 3800
rect 32136 3760 32148 3794
rect 32612 3760 32624 3794
rect 32136 3754 32624 3760
rect 33154 3794 33642 3800
rect 33154 3760 33166 3794
rect 33630 3760 33642 3794
rect 33154 3754 33642 3760
rect 31844 3650 31854 3710
rect 30870 3134 30878 3184
rect 30100 3084 30588 3090
rect 30100 3050 30112 3084
rect 30576 3050 30588 3084
rect 30100 3044 30588 3050
rect 30306 2888 30366 3044
rect 30818 2996 30878 3134
rect 31848 3134 31854 3650
rect 31888 3650 31904 3710
rect 32866 3710 32912 3722
rect 31888 3134 31894 3650
rect 32866 3178 32872 3710
rect 31848 3122 31894 3134
rect 32860 3134 32872 3178
rect 32906 3178 32912 3710
rect 33884 3710 33930 3722
rect 32906 3134 32920 3178
rect 33884 3176 33890 3710
rect 31118 3084 31606 3090
rect 31118 3050 31130 3084
rect 31594 3050 31606 3084
rect 31118 3044 31606 3050
rect 32136 3084 32624 3090
rect 32136 3050 32148 3084
rect 32612 3050 32624 3084
rect 32136 3044 32624 3050
rect 30812 2936 30818 2996
rect 30878 2936 30884 2996
rect 30306 2882 30368 2888
rect 30306 2822 30308 2882
rect 30306 2816 30368 2822
rect 27760 2614 27766 2674
rect 27826 2614 27832 2674
rect 28282 2614 28288 2674
rect 28348 2614 28354 2674
rect 28782 2614 28788 2674
rect 28848 2614 28854 2674
rect 29290 2614 29296 2674
rect 29356 2614 29362 2674
rect 29798 2614 29804 2674
rect 29864 2614 29870 2674
rect 30148 2614 30154 2674
rect 30214 2614 30220 2674
rect 30306 2672 30366 2816
rect 31330 2778 31390 3044
rect 32332 2778 32392 3044
rect 32860 2996 32920 3134
rect 33878 3134 33890 3176
rect 33924 3176 33930 3710
rect 33924 3134 33938 3176
rect 33154 3084 33642 3090
rect 33154 3050 33166 3084
rect 33630 3050 33642 3084
rect 33154 3044 33642 3050
rect 33372 2996 33432 3044
rect 33878 2996 33938 3134
rect 32854 2936 32860 2996
rect 32920 2936 32926 2996
rect 33366 2936 33372 2996
rect 33432 2936 33438 2996
rect 33872 2936 33878 2996
rect 33938 2936 33944 2996
rect 31324 2718 31330 2778
rect 31390 2718 31396 2778
rect 32326 2718 32332 2778
rect 32392 2718 32398 2778
rect 27046 2560 27534 2566
rect 27046 2526 27058 2560
rect 27522 2526 27534 2560
rect 27046 2520 27534 2526
rect 24762 1966 24768 2442
rect 25734 2400 25746 2476
rect 24762 1900 24776 1966
rect 22974 1850 23462 1856
rect 22974 1816 22986 1850
rect 23450 1816 23462 1850
rect 22974 1810 23462 1816
rect 23992 1850 24480 1856
rect 23992 1816 24004 1850
rect 24468 1816 24480 1850
rect 23992 1810 24480 1816
rect 22674 1682 22680 1742
rect 22740 1682 22746 1742
rect 23182 1638 23242 1810
rect 24208 1638 24268 1810
rect 24716 1742 24776 1900
rect 25740 1900 25746 2400
rect 25780 2400 25794 2476
rect 26746 2426 26764 2476
rect 25780 1900 25786 2400
rect 26758 1932 26764 2426
rect 25740 1888 25786 1900
rect 26748 1900 26764 1932
rect 26798 2428 26810 2476
rect 27766 2476 27826 2614
rect 28288 2566 28348 2614
rect 28064 2560 28552 2566
rect 28064 2526 28076 2560
rect 28540 2526 28552 2560
rect 28064 2520 28552 2526
rect 28288 2514 28348 2520
rect 28788 2476 28848 2614
rect 29296 2566 29356 2614
rect 29082 2560 29570 2566
rect 29082 2526 29094 2560
rect 29558 2526 29570 2560
rect 29082 2520 29570 2526
rect 26798 2426 26806 2428
rect 26798 1932 26804 2426
rect 27766 2420 27782 2476
rect 26798 1900 26808 1932
rect 25010 1850 25498 1856
rect 25010 1816 25022 1850
rect 25486 1816 25498 1850
rect 25010 1810 25498 1816
rect 26028 1850 26516 1856
rect 26028 1816 26040 1850
rect 26504 1816 26516 1850
rect 26028 1810 26516 1816
rect 26236 1750 26296 1810
rect 26748 1750 26808 1900
rect 27776 1900 27782 2420
rect 27816 2420 27826 2476
rect 27816 1900 27822 2420
rect 28782 2416 28800 2476
rect 28794 1938 28800 2416
rect 28784 1900 28800 1938
rect 28834 2416 28848 2476
rect 29804 2476 29864 2614
rect 30154 2566 30214 2614
rect 30306 2612 30884 2672
rect 30100 2560 30588 2566
rect 30100 2526 30112 2560
rect 30576 2526 30588 2560
rect 30100 2520 30588 2526
rect 29804 2442 29818 2476
rect 28834 1938 28840 2416
rect 28834 1900 28844 1938
rect 29812 1900 29818 2442
rect 29852 2442 29864 2476
rect 30824 2476 30884 2612
rect 34044 2610 34104 3932
rect 31118 2560 31606 2566
rect 31118 2526 31130 2560
rect 31594 2526 31606 2560
rect 31118 2520 31606 2526
rect 32136 2560 32624 2566
rect 32136 2526 32148 2560
rect 32612 2526 32624 2560
rect 32136 2520 32624 2526
rect 33154 2560 33642 2566
rect 33154 2526 33166 2560
rect 33630 2526 33642 2560
rect 33154 2520 33642 2526
rect 33884 2550 34104 2610
rect 29852 1900 29858 2442
rect 30824 2438 30836 2476
rect 27776 1888 27822 1900
rect 28794 1888 28840 1900
rect 29812 1888 29858 1900
rect 30830 1900 30836 2438
rect 30870 2438 30884 2476
rect 31848 2476 31894 2488
rect 30870 1900 30876 2438
rect 31848 1932 31854 2476
rect 30830 1888 30876 1900
rect 31838 1900 31854 1932
rect 31888 1932 31894 2476
rect 32866 2476 32912 2488
rect 32866 1948 32872 2476
rect 31888 1900 31898 1932
rect 27046 1850 27534 1856
rect 27046 1816 27058 1850
rect 27522 1816 27534 1850
rect 27046 1810 27534 1816
rect 28064 1850 28552 1856
rect 28064 1816 28076 1850
rect 28540 1816 28552 1850
rect 28064 1810 28552 1816
rect 29082 1850 29570 1856
rect 29082 1816 29094 1850
rect 29558 1816 29570 1850
rect 29082 1810 29570 1816
rect 30100 1850 30588 1856
rect 30100 1816 30112 1850
rect 30576 1816 30588 1850
rect 30100 1810 30588 1816
rect 31118 1850 31606 1856
rect 31118 1816 31130 1850
rect 31594 1816 31606 1850
rect 31118 1810 31606 1816
rect 27254 1750 27314 1810
rect 24710 1682 24716 1742
rect 24776 1682 24782 1742
rect 26236 1690 27314 1750
rect 22170 1578 24268 1638
rect 16562 1482 16568 1542
rect 16628 1482 16634 1542
rect 18600 1482 18606 1542
rect 18666 1482 18672 1542
rect 20632 1482 20638 1542
rect 20698 1482 20704 1542
rect 22670 1482 22676 1542
rect 22736 1482 22742 1542
rect 24704 1482 24710 1542
rect 24770 1482 24776 1542
rect 26744 1482 26750 1542
rect 26810 1482 26816 1542
rect 28778 1482 28784 1542
rect 28844 1482 28850 1542
rect 30812 1482 30818 1542
rect 30878 1482 30884 1542
rect 15848 1328 16336 1334
rect 15848 1294 15860 1328
rect 16324 1294 16336 1328
rect 15848 1288 16336 1294
rect 14582 718 14588 1206
rect 15548 1196 15566 1244
rect 14582 668 14592 718
rect 13812 618 14300 624
rect 13812 584 13824 618
rect 14288 584 14300 618
rect 13812 578 14300 584
rect 14016 512 14076 578
rect 14532 512 14592 668
rect 15560 668 15566 1196
rect 15600 1196 15608 1244
rect 16568 1244 16628 1482
rect 17580 1384 17586 1444
rect 17646 1384 17652 1444
rect 16866 1328 17354 1334
rect 16866 1294 16878 1328
rect 17342 1294 17354 1328
rect 16866 1288 17354 1294
rect 16568 1212 16584 1244
rect 15600 668 15606 1196
rect 16578 696 16584 1212
rect 15560 656 15606 668
rect 16570 668 16584 696
rect 16618 1212 16628 1244
rect 17586 1244 17646 1384
rect 17884 1328 18372 1334
rect 17884 1294 17896 1328
rect 18360 1294 18372 1328
rect 17884 1288 18372 1294
rect 16618 696 16624 1212
rect 17586 1188 17602 1244
rect 16618 668 16630 696
rect 14830 618 15318 624
rect 14830 584 14842 618
rect 15306 584 15318 618
rect 14830 578 15318 584
rect 15848 618 16336 624
rect 15848 584 15860 618
rect 16324 584 16336 618
rect 15848 578 16336 584
rect 15064 512 15124 578
rect 16054 512 16114 578
rect 16570 512 16630 668
rect 17596 668 17602 1188
rect 17636 1188 17646 1244
rect 18606 1244 18666 1482
rect 19616 1384 19622 1444
rect 19682 1384 19688 1444
rect 18902 1328 19390 1334
rect 18902 1294 18914 1328
rect 19378 1294 19390 1328
rect 18902 1288 19390 1294
rect 18606 1198 18620 1244
rect 17636 668 17642 1188
rect 18614 696 18620 1198
rect 17596 656 17642 668
rect 18606 668 18620 696
rect 18654 1198 18666 1244
rect 19622 1244 19682 1384
rect 19920 1328 20408 1334
rect 19920 1294 19932 1328
rect 20396 1294 20408 1328
rect 19920 1288 20408 1294
rect 18654 696 18660 1198
rect 19622 1194 19638 1244
rect 18654 668 18666 696
rect 16866 618 17354 624
rect 16866 584 16878 618
rect 17342 584 17354 618
rect 16866 578 17354 584
rect 17884 618 18372 624
rect 17884 584 17896 618
rect 18360 584 18372 618
rect 17884 578 18372 584
rect 17076 512 17136 578
rect 18098 512 18158 578
rect 18606 512 18666 668
rect 19632 668 19638 1194
rect 19672 1194 19682 1244
rect 20638 1244 20698 1482
rect 21652 1384 21658 1444
rect 21718 1384 21724 1444
rect 20938 1328 21426 1334
rect 20938 1294 20950 1328
rect 21414 1294 21426 1328
rect 20938 1288 21426 1294
rect 19672 668 19678 1194
rect 20638 1188 20656 1244
rect 20650 702 20656 1188
rect 19632 656 19678 668
rect 20640 668 20656 702
rect 20690 1188 20698 1244
rect 21658 1244 21718 1384
rect 21956 1328 22444 1334
rect 21956 1294 21968 1328
rect 22432 1294 22444 1328
rect 21956 1288 22444 1294
rect 21658 1196 21674 1244
rect 20690 702 20696 1188
rect 20690 668 20700 702
rect 18902 618 19390 624
rect 18902 584 18914 618
rect 19378 584 19390 618
rect 18902 578 19390 584
rect 19920 618 20408 624
rect 19920 584 19932 618
rect 20396 584 20408 618
rect 19920 578 20408 584
rect 19120 512 19180 578
rect 20130 512 20190 578
rect 20640 512 20700 668
rect 21668 668 21674 1196
rect 21708 1196 21718 1244
rect 22676 1244 22736 1482
rect 23688 1384 23694 1444
rect 23754 1384 23760 1444
rect 22974 1328 23462 1334
rect 22974 1294 22986 1328
rect 23450 1294 23462 1328
rect 22974 1288 23462 1294
rect 22676 1200 22692 1244
rect 21708 668 21714 1196
rect 22686 726 22692 1200
rect 21668 656 21714 668
rect 22680 668 22692 726
rect 22726 1200 22736 1244
rect 23694 1244 23754 1384
rect 23992 1328 24480 1334
rect 23992 1294 24004 1328
rect 24468 1294 24480 1328
rect 23992 1288 24480 1294
rect 23694 1202 23710 1244
rect 22726 726 22732 1200
rect 22726 668 22740 726
rect 20938 618 21426 624
rect 20938 584 20950 618
rect 21414 584 21426 618
rect 20938 578 21426 584
rect 21956 618 22444 624
rect 21956 584 21968 618
rect 22432 584 22444 618
rect 21956 578 22444 584
rect 21158 512 21218 578
rect 22176 512 22236 578
rect 22680 512 22740 668
rect 23704 668 23710 1202
rect 23744 1202 23754 1244
rect 24710 1244 24770 1482
rect 25722 1384 25728 1444
rect 25788 1384 25794 1444
rect 25010 1328 25498 1334
rect 25010 1294 25022 1328
rect 25486 1294 25498 1328
rect 25010 1288 25498 1294
rect 23744 668 23750 1202
rect 24710 1188 24728 1244
rect 24722 698 24728 1188
rect 23704 656 23750 668
rect 24718 668 24728 698
rect 24762 1188 24770 1244
rect 25728 1244 25788 1384
rect 26028 1328 26516 1334
rect 26028 1294 26040 1328
rect 26504 1294 26516 1328
rect 26028 1288 26516 1294
rect 25728 1202 25746 1244
rect 24762 698 24768 1188
rect 24762 668 24778 698
rect 22974 618 23462 624
rect 22974 584 22986 618
rect 23450 584 23462 618
rect 22974 578 23462 584
rect 23992 618 24480 624
rect 23992 584 24004 618
rect 24468 584 24480 618
rect 23992 578 24480 584
rect 23192 512 23252 578
rect 24214 512 24274 578
rect 24718 512 24778 668
rect 25740 668 25746 1202
rect 25780 1202 25788 1244
rect 26750 1244 26810 1482
rect 27758 1384 27764 1444
rect 27824 1384 27830 1444
rect 27046 1328 27534 1334
rect 27046 1294 27058 1328
rect 27522 1294 27534 1328
rect 27046 1288 27534 1294
rect 25780 668 25786 1202
rect 26750 1198 26764 1244
rect 26758 712 26764 1198
rect 25740 656 25786 668
rect 26752 668 26764 712
rect 26798 1198 26810 1244
rect 27764 1244 27824 1384
rect 28064 1328 28552 1334
rect 28064 1294 28076 1328
rect 28540 1294 28552 1328
rect 28064 1288 28552 1294
rect 27764 1198 27782 1244
rect 26798 712 26804 1198
rect 26798 668 26812 712
rect 25010 618 25498 624
rect 25010 584 25022 618
rect 25486 584 25498 618
rect 25010 578 25498 584
rect 26028 618 26516 624
rect 26028 584 26040 618
rect 26504 584 26516 618
rect 26028 578 26516 584
rect 25236 512 25296 578
rect 26244 512 26304 578
rect 26752 512 26812 668
rect 27776 668 27782 1198
rect 27816 1198 27824 1244
rect 28784 1244 28844 1482
rect 29798 1384 29804 1444
rect 29864 1384 29870 1444
rect 29082 1328 29570 1334
rect 29082 1294 29094 1328
rect 29558 1294 29570 1328
rect 29082 1288 29570 1294
rect 27816 668 27822 1198
rect 28784 1186 28800 1244
rect 28794 708 28800 1186
rect 27776 656 27822 668
rect 28788 668 28800 708
rect 28834 1186 28844 1244
rect 29804 1244 29864 1384
rect 30100 1328 30588 1334
rect 30100 1294 30112 1328
rect 30576 1294 30588 1328
rect 30100 1288 30588 1294
rect 29804 1212 29818 1244
rect 28834 708 28840 1186
rect 28834 668 28848 708
rect 27248 624 27308 626
rect 27046 618 27534 624
rect 27046 584 27058 618
rect 27522 584 27534 618
rect 27046 578 27534 584
rect 28064 618 28552 624
rect 28064 584 28076 618
rect 28540 584 28552 618
rect 28064 578 28552 584
rect 27248 512 27308 578
rect 28294 512 28354 578
rect 28788 512 28848 668
rect 29812 668 29818 1212
rect 29852 1212 29864 1244
rect 30818 1244 30878 1482
rect 31316 1334 31376 1810
rect 31838 1444 31898 1900
rect 32856 1900 32872 1948
rect 32906 1948 32912 2476
rect 33884 2476 33944 2550
rect 32906 1900 32916 1948
rect 33884 1934 33890 2476
rect 32136 1850 32624 1856
rect 32136 1816 32148 1850
rect 32612 1816 32624 1850
rect 32136 1810 32624 1816
rect 31832 1384 31838 1444
rect 31898 1384 31904 1444
rect 31118 1328 31606 1334
rect 31118 1294 31130 1328
rect 31594 1294 31606 1328
rect 31118 1288 31606 1294
rect 29852 668 29858 1212
rect 30818 1202 30836 1244
rect 30830 702 30836 1202
rect 29812 656 29858 668
rect 30826 668 30836 702
rect 30870 1202 30878 1244
rect 31838 1244 31898 1384
rect 32344 1334 32404 1810
rect 32856 1542 32916 1900
rect 33874 1900 33890 1934
rect 33924 2400 33944 2476
rect 33924 1934 33930 2400
rect 33924 1900 33934 1934
rect 33154 1850 33642 1856
rect 33154 1816 33166 1850
rect 33630 1816 33642 1850
rect 33154 1810 33642 1816
rect 32850 1482 32856 1542
rect 32916 1482 32922 1542
rect 32136 1328 32624 1334
rect 32136 1294 32148 1328
rect 32612 1294 32624 1328
rect 32136 1288 32624 1294
rect 31838 1204 31854 1244
rect 30870 702 30876 1202
rect 30870 668 30886 702
rect 29082 618 29570 624
rect 29082 584 29094 618
rect 29558 584 29570 618
rect 29082 578 29570 584
rect 30100 618 30588 624
rect 30100 584 30112 618
rect 30576 584 30588 618
rect 30100 578 30588 584
rect 29292 512 29352 578
rect 30304 512 30364 578
rect 30826 512 30886 668
rect 31848 668 31854 1204
rect 31888 1204 31898 1244
rect 32856 1244 32916 1482
rect 33336 1334 33396 1810
rect 33874 1444 33934 1900
rect 34598 1542 34658 13934
rect 34750 2614 34756 2674
rect 34816 2614 34822 2674
rect 34592 1482 34598 1542
rect 34658 1482 34664 1542
rect 33868 1384 33874 1444
rect 33934 1384 33940 1444
rect 33154 1328 33642 1334
rect 33154 1294 33166 1328
rect 33630 1294 33642 1328
rect 33154 1288 33642 1294
rect 33336 1286 33396 1288
rect 32856 1214 32872 1244
rect 31888 668 31894 1204
rect 32866 696 32872 1214
rect 31848 656 31894 668
rect 32854 668 32872 696
rect 32906 1214 32916 1244
rect 33874 1244 33934 1384
rect 32906 696 32912 1214
rect 33874 1208 33890 1244
rect 32906 668 32914 696
rect 31118 618 31606 624
rect 31118 584 31130 618
rect 31594 584 31606 618
rect 31118 578 31606 584
rect 32136 618 32624 624
rect 32136 584 32148 618
rect 32612 584 32624 618
rect 32136 578 32624 584
rect 31326 512 31386 578
rect 32392 512 32452 578
rect 32854 512 32914 668
rect 33884 668 33890 1208
rect 33924 1208 33934 1244
rect 33924 668 33930 1208
rect 33884 656 33930 668
rect 33154 618 33642 624
rect 33154 584 33166 618
rect 33630 584 33642 618
rect 33154 578 33642 584
rect 33354 512 33414 578
rect 14016 452 33414 512
rect 34756 110 34816 2614
rect 35766 210 35772 14470
rect 35872 210 35878 14470
rect 48494 8574 48554 8578
rect 50076 8574 50476 23478
rect 65322 18278 65328 27642
rect 65428 18278 65434 27642
rect 68948 27774 85828 27806
rect 68948 27560 69011 27774
rect 85796 27560 85828 27774
rect 68948 27540 85828 27560
rect 89666 27642 89778 28156
rect 68948 27538 73302 27540
rect 68564 21978 68952 22038
rect 68564 21838 68624 21978
rect 68666 21937 68726 21978
rect 68658 21931 68746 21937
rect 68658 21897 68670 21931
rect 68734 21897 68746 21931
rect 68658 21891 68746 21897
rect 68564 21810 68576 21838
rect 68570 21462 68576 21810
rect 68610 21810 68624 21838
rect 68782 21838 68842 21978
rect 68892 21937 68952 21978
rect 68876 21931 68964 21937
rect 68876 21897 68888 21931
rect 68952 21897 68964 21931
rect 68876 21891 68964 21897
rect 68610 21462 68616 21810
rect 68782 21806 68794 21838
rect 68788 21492 68794 21806
rect 68570 21450 68616 21462
rect 68782 21462 68794 21492
rect 68828 21806 68842 21838
rect 68998 21838 69058 27538
rect 69100 21978 69106 22038
rect 69166 21978 69172 22038
rect 69212 21978 69218 22038
rect 69278 21978 69284 22038
rect 69322 21978 69328 22038
rect 69388 21978 69394 22038
rect 69106 21937 69166 21978
rect 69094 21931 69182 21937
rect 69094 21897 69106 21931
rect 69170 21897 69182 21931
rect 69094 21891 69182 21897
rect 68828 21492 68834 21806
rect 68828 21462 68842 21492
rect 68658 21403 68746 21409
rect 68658 21369 68670 21403
rect 68734 21369 68746 21403
rect 68658 21363 68746 21369
rect 68782 21326 68842 21462
rect 68998 21462 69012 21838
rect 69046 21462 69058 21838
rect 69218 21838 69278 21978
rect 69328 21937 69388 21978
rect 69312 21931 69400 21937
rect 69312 21897 69324 21931
rect 69388 21897 69400 21931
rect 69312 21891 69400 21897
rect 69218 21812 69230 21838
rect 68876 21403 68964 21409
rect 68876 21369 68888 21403
rect 68952 21369 68964 21403
rect 68876 21363 68964 21369
rect 68892 21326 68952 21363
rect 68436 21266 68442 21326
rect 68502 21266 68508 21326
rect 68776 21266 68782 21326
rect 68842 21266 68848 21326
rect 68886 21266 68892 21326
rect 68952 21266 68958 21326
rect 67054 20320 67060 20380
rect 67120 20320 67126 20380
rect 65322 17764 65434 18278
rect 67060 18148 67120 20320
rect 68442 19542 68502 21266
rect 68998 21220 69058 21462
rect 69224 21462 69230 21812
rect 69264 21812 69278 21838
rect 69434 21838 69494 27538
rect 69530 21931 69618 21937
rect 69530 21897 69542 21931
rect 69606 21897 69618 21931
rect 69530 21891 69618 21897
rect 69748 21931 69836 21937
rect 69748 21897 69760 21931
rect 69824 21897 69836 21931
rect 69748 21891 69836 21897
rect 69264 21462 69270 21812
rect 69224 21450 69270 21462
rect 69434 21462 69448 21838
rect 69482 21462 69494 21838
rect 69660 21838 69706 21850
rect 69660 21494 69666 21838
rect 69094 21403 69182 21409
rect 69094 21369 69106 21403
rect 69170 21369 69182 21403
rect 69094 21363 69182 21369
rect 69312 21403 69400 21409
rect 69312 21369 69324 21403
rect 69388 21369 69400 21403
rect 69312 21363 69400 21369
rect 69434 21220 69494 21462
rect 69654 21462 69666 21494
rect 69700 21494 69706 21838
rect 69872 21838 69932 27538
rect 69972 21978 69978 22038
rect 70038 21978 70044 22038
rect 70082 21978 70088 22038
rect 70148 21978 70154 22038
rect 70190 21978 70196 22038
rect 70256 21978 70262 22038
rect 69978 21937 70038 21978
rect 69966 21931 70054 21937
rect 69966 21897 69978 21931
rect 70042 21897 70054 21931
rect 69966 21891 70054 21897
rect 69700 21462 69714 21494
rect 69530 21403 69618 21409
rect 69530 21369 69542 21403
rect 69606 21369 69618 21403
rect 69530 21363 69618 21369
rect 69542 21326 69602 21363
rect 69654 21326 69714 21462
rect 69872 21462 69884 21838
rect 69918 21462 69932 21838
rect 70088 21838 70148 21978
rect 70196 21937 70256 21978
rect 70184 21931 70272 21937
rect 70184 21897 70196 21931
rect 70260 21897 70272 21931
rect 70184 21891 70272 21897
rect 70088 21810 70102 21838
rect 69748 21403 69836 21409
rect 69748 21369 69760 21403
rect 69824 21369 69836 21403
rect 69748 21363 69836 21369
rect 69762 21326 69822 21363
rect 69536 21266 69542 21326
rect 69602 21266 69608 21326
rect 69648 21266 69654 21326
rect 69714 21266 69720 21326
rect 69756 21266 69762 21326
rect 69822 21266 69828 21326
rect 69872 21220 69932 21462
rect 70096 21462 70102 21810
rect 70136 21810 70148 21838
rect 70306 21838 70366 27538
rect 72930 27364 72936 27424
rect 72996 27364 73002 27424
rect 71424 27148 72502 27208
rect 71424 26968 71484 27148
rect 71928 27067 71988 27148
rect 71720 27061 72208 27067
rect 71720 27027 71732 27061
rect 72196 27027 72208 27061
rect 71720 27021 72208 27027
rect 71424 26928 71438 26968
rect 71432 26392 71438 26928
rect 71472 26928 71484 26968
rect 72442 26968 72502 27148
rect 72936 27067 72996 27364
rect 73462 27178 73522 27540
rect 74012 27364 74018 27424
rect 74078 27364 74084 27424
rect 74970 27364 74976 27424
rect 75036 27364 75042 27424
rect 73456 27118 73462 27178
rect 73522 27118 73528 27178
rect 72738 27061 73226 27067
rect 72738 27027 72750 27061
rect 73214 27027 73226 27061
rect 72738 27021 73226 27027
rect 72442 26942 72456 26968
rect 71472 26392 71478 26928
rect 72450 26428 72456 26942
rect 71432 26380 71478 26392
rect 72444 26392 72456 26428
rect 72490 26942 72502 26968
rect 73462 26968 73522 27118
rect 74018 27067 74078 27364
rect 74976 27067 75036 27364
rect 75498 27178 75558 27540
rect 76006 27364 76012 27424
rect 76072 27364 76078 27424
rect 77012 27364 77018 27424
rect 77078 27364 77084 27424
rect 75492 27118 75498 27178
rect 75558 27118 75564 27178
rect 73756 27061 74244 27067
rect 73756 27027 73768 27061
rect 74232 27027 74244 27061
rect 73756 27021 74244 27027
rect 74774 27061 75262 27067
rect 74774 27027 74786 27061
rect 75250 27027 75262 27061
rect 74774 27021 75262 27027
rect 74976 27018 75036 27021
rect 73462 26944 73474 26968
rect 72490 26428 72496 26942
rect 73468 26432 73474 26944
rect 72490 26392 72504 26428
rect 71720 26333 72208 26339
rect 71720 26299 71732 26333
rect 72196 26299 72208 26333
rect 71720 26293 72208 26299
rect 72444 26246 72504 26392
rect 73464 26392 73474 26432
rect 73508 26944 73522 26968
rect 74486 26968 74532 26980
rect 73508 26432 73514 26944
rect 73508 26392 73524 26432
rect 74486 26420 74492 26968
rect 72948 26339 73008 26340
rect 72738 26333 73226 26339
rect 72738 26299 72750 26333
rect 73214 26299 73226 26333
rect 72738 26293 73226 26299
rect 71274 26186 71280 26246
rect 71340 26186 71346 26246
rect 72438 26186 72444 26246
rect 72504 26186 72510 26246
rect 71144 25982 71150 26042
rect 71210 25982 71216 26042
rect 71150 23114 71210 25982
rect 71280 23572 71340 26186
rect 72438 25982 72444 26042
rect 72504 25982 72510 26042
rect 71720 25925 72208 25931
rect 71720 25891 71732 25925
rect 72196 25891 72208 25925
rect 71720 25885 72208 25891
rect 71432 25832 71478 25844
rect 71432 25292 71438 25832
rect 71426 25256 71438 25292
rect 71472 25292 71478 25832
rect 72444 25832 72504 25982
rect 72948 25931 73008 26293
rect 72738 25925 73226 25931
rect 72738 25891 72750 25925
rect 73214 25891 73226 25925
rect 72738 25885 73226 25891
rect 72948 25882 73008 25885
rect 72444 25794 72456 25832
rect 71472 25256 71486 25292
rect 72450 25286 72456 25794
rect 71426 25106 71486 25256
rect 72444 25256 72456 25286
rect 72490 25794 72504 25832
rect 73464 25832 73524 26392
rect 74480 26392 74492 26420
rect 74526 26420 74532 26968
rect 75498 26968 75558 27118
rect 76012 27067 76072 27364
rect 76510 27230 76516 27290
rect 76576 27230 76582 27290
rect 75792 27061 76280 27067
rect 75792 27027 75804 27061
rect 76268 27027 76280 27061
rect 75792 27021 76280 27027
rect 76012 27018 76072 27021
rect 75498 26944 75510 26968
rect 75504 26450 75510 26944
rect 74526 26392 74540 26420
rect 73970 26339 74030 26346
rect 73756 26333 74244 26339
rect 73756 26299 73768 26333
rect 74232 26299 74244 26333
rect 73756 26293 74244 26299
rect 73970 25931 74030 26293
rect 74480 26142 74540 26392
rect 75488 26392 75510 26450
rect 75544 26944 75558 26968
rect 76516 26968 76576 27230
rect 77018 27067 77078 27364
rect 77536 27180 77596 27540
rect 78034 27364 78040 27424
rect 78100 27364 78106 27424
rect 79052 27364 79058 27424
rect 79118 27364 79124 27424
rect 77530 27120 77536 27180
rect 77596 27120 77602 27180
rect 76810 27061 77298 27067
rect 76810 27027 76822 27061
rect 77286 27027 77298 27061
rect 76810 27021 77298 27027
rect 75544 26450 75550 26944
rect 76516 26940 76528 26968
rect 75544 26392 75552 26450
rect 75000 26339 75060 26346
rect 74774 26333 75262 26339
rect 74774 26299 74786 26333
rect 75250 26299 75262 26333
rect 74774 26293 75262 26299
rect 74474 26082 74480 26142
rect 74540 26082 74546 26142
rect 75000 25931 75060 26293
rect 73756 25925 74244 25931
rect 73756 25891 73768 25925
rect 74232 25891 74244 25925
rect 73756 25885 74244 25891
rect 74774 25925 75262 25931
rect 74774 25891 74786 25925
rect 75250 25891 75262 25925
rect 74774 25885 75262 25891
rect 72490 25286 72496 25794
rect 73464 25792 73474 25832
rect 72490 25256 72504 25286
rect 73468 25282 73474 25792
rect 71720 25197 72208 25203
rect 71720 25163 71732 25197
rect 72196 25163 72208 25197
rect 71720 25157 72208 25163
rect 71938 25106 71998 25157
rect 72444 25106 72504 25256
rect 73460 25256 73474 25282
rect 73508 25792 73524 25832
rect 74486 25832 74532 25844
rect 73508 25282 73514 25792
rect 73508 25256 73520 25282
rect 74486 25276 74492 25832
rect 72930 25203 72990 25210
rect 72738 25197 73226 25203
rect 72738 25163 72750 25197
rect 73214 25163 73226 25197
rect 72738 25157 73226 25163
rect 71426 25046 72504 25106
rect 72438 24898 72498 24904
rect 71428 24838 72498 24898
rect 71428 24696 71488 24838
rect 71938 24795 71998 24838
rect 71720 24789 72208 24795
rect 71720 24755 71732 24789
rect 72196 24755 72208 24789
rect 71720 24749 72208 24755
rect 71428 24664 71438 24696
rect 71432 24120 71438 24664
rect 71472 24664 71488 24696
rect 72438 24696 72498 24838
rect 72930 24795 72990 25157
rect 73460 25108 73520 25256
rect 74478 25256 74492 25276
rect 74526 25276 74532 25832
rect 75488 25832 75552 26392
rect 76522 26392 76528 26940
rect 76562 26940 76576 26968
rect 77536 26968 77596 27120
rect 78040 27067 78100 27364
rect 79058 27067 79118 27364
rect 79568 27180 79628 27540
rect 80076 27364 80082 27424
rect 80142 27364 80148 27424
rect 81088 27364 81094 27424
rect 81154 27364 81160 27424
rect 79560 27120 79566 27180
rect 79626 27120 79632 27180
rect 77828 27061 78316 27067
rect 77828 27027 77840 27061
rect 78304 27027 78316 27061
rect 77828 27021 78316 27027
rect 78846 27061 79334 27067
rect 78846 27027 78858 27061
rect 79322 27027 79334 27061
rect 78846 27021 79334 27027
rect 76562 26392 76568 26940
rect 77536 26928 77546 26968
rect 77540 26446 77546 26928
rect 76522 26380 76568 26392
rect 77524 26392 77546 26446
rect 77580 26928 77596 26968
rect 78558 26968 78604 26980
rect 77580 26446 77586 26928
rect 77580 26392 77588 26446
rect 78558 26432 78564 26968
rect 76000 26339 76060 26352
rect 77018 26339 77078 26346
rect 75792 26333 76280 26339
rect 75792 26299 75804 26333
rect 76268 26299 76280 26333
rect 75792 26293 76280 26299
rect 76810 26333 77298 26339
rect 76810 26299 76822 26333
rect 77286 26299 77298 26333
rect 76810 26293 77298 26299
rect 76000 25931 76060 26293
rect 76510 26082 76516 26142
rect 76576 26082 76582 26142
rect 75792 25925 76280 25931
rect 75792 25891 75804 25925
rect 76268 25891 76280 25925
rect 75792 25885 76280 25891
rect 75488 25802 75510 25832
rect 75504 25284 75510 25802
rect 74526 25256 74538 25276
rect 73976 25203 74036 25210
rect 73756 25197 74244 25203
rect 73756 25163 73768 25197
rect 74232 25163 74244 25197
rect 73756 25157 74244 25163
rect 73454 25048 73460 25108
rect 73520 25048 73526 25108
rect 72738 24789 73226 24795
rect 72738 24755 72750 24789
rect 73214 24755 73226 24789
rect 72738 24749 73226 24755
rect 72438 24664 72456 24696
rect 71472 24120 71478 24664
rect 72450 24162 72456 24664
rect 71432 24108 71478 24120
rect 72438 24120 72456 24162
rect 72490 24664 72498 24696
rect 73460 24696 73520 25048
rect 73976 24795 74036 25157
rect 74478 25012 74538 25256
rect 75496 25256 75510 25284
rect 75544 25802 75552 25832
rect 76516 25832 76576 26082
rect 77018 25931 77078 26293
rect 76810 25925 77298 25931
rect 76810 25891 76822 25925
rect 77286 25891 77298 25925
rect 76810 25885 77298 25891
rect 75544 25284 75550 25802
rect 76516 25794 76528 25832
rect 76522 25292 76528 25794
rect 75544 25282 75556 25284
rect 75544 25256 75560 25282
rect 74774 25197 75262 25203
rect 74774 25163 74786 25197
rect 75250 25163 75262 25197
rect 74774 25157 75262 25163
rect 75496 25108 75560 25256
rect 76514 25256 76528 25292
rect 76562 25794 76576 25832
rect 77524 25832 77588 26392
rect 78554 26392 78564 26432
rect 78598 26432 78604 26968
rect 79568 26968 79628 27120
rect 80082 27067 80142 27364
rect 81094 27067 81154 27364
rect 81608 27182 81668 27540
rect 82106 27364 82112 27424
rect 82172 27364 82178 27424
rect 83118 27364 83124 27424
rect 83184 27364 83190 27424
rect 81602 27122 81608 27182
rect 81668 27122 81674 27182
rect 79864 27061 80352 27067
rect 79864 27027 79876 27061
rect 80340 27027 80352 27061
rect 79864 27021 80352 27027
rect 80882 27061 81370 27067
rect 80882 27027 80894 27061
rect 81358 27027 81370 27061
rect 80882 27021 81370 27027
rect 79568 26928 79582 26968
rect 79576 26448 79582 26928
rect 78598 26392 78614 26432
rect 78042 26339 78102 26342
rect 77828 26333 78316 26339
rect 77828 26299 77840 26333
rect 78304 26299 78316 26333
rect 77828 26293 78316 26299
rect 78042 25931 78102 26293
rect 78554 26246 78614 26392
rect 79566 26392 79582 26448
rect 79616 26928 79628 26968
rect 80594 26968 80640 26980
rect 79616 26448 79622 26928
rect 79616 26392 79630 26448
rect 80594 26430 80600 26968
rect 79060 26339 79120 26348
rect 78846 26333 79334 26339
rect 78846 26299 78858 26333
rect 79322 26299 79334 26333
rect 78846 26293 79334 26299
rect 78548 26186 78554 26246
rect 78614 26186 78620 26246
rect 78544 25982 78550 26042
rect 78610 25982 78616 26042
rect 77828 25925 78316 25931
rect 77828 25891 77840 25925
rect 78304 25891 78316 25925
rect 77828 25885 78316 25891
rect 78042 25884 78102 25885
rect 77524 25798 77546 25832
rect 76562 25292 76568 25794
rect 77540 25292 77546 25798
rect 76562 25256 76578 25292
rect 76024 25203 76084 25216
rect 75792 25197 76280 25203
rect 75792 25163 75804 25197
rect 76268 25163 76280 25197
rect 75792 25157 76280 25163
rect 75490 25048 75496 25108
rect 75556 25048 75562 25108
rect 74472 24952 74478 25012
rect 74538 24952 74544 25012
rect 75176 24946 75182 25010
rect 75246 24946 75252 25010
rect 75182 24916 75246 24946
rect 74480 24852 75246 24916
rect 73756 24789 74244 24795
rect 73756 24755 73768 24789
rect 74232 24755 74244 24789
rect 73756 24749 74244 24755
rect 72490 24162 72496 24664
rect 73460 24644 73474 24696
rect 72490 24120 72502 24162
rect 73468 24156 73474 24644
rect 71720 24061 72208 24067
rect 71720 24027 71732 24061
rect 72196 24027 72208 24061
rect 71720 24021 72208 24027
rect 72438 23722 72502 24120
rect 73460 24120 73474 24156
rect 73508 24644 73520 24696
rect 74480 24696 74544 24852
rect 74774 24789 75262 24795
rect 74774 24755 74786 24789
rect 75250 24755 75262 24789
rect 74774 24749 75262 24755
rect 74480 24650 74492 24696
rect 73508 24156 73514 24644
rect 73508 24120 73520 24156
rect 74486 24144 74492 24650
rect 72738 24061 73226 24067
rect 72738 24027 72750 24061
rect 73214 24027 73226 24061
rect 72738 24021 73226 24027
rect 73460 23970 73520 24120
rect 74476 24120 74492 24144
rect 74526 24650 74544 24696
rect 75496 24696 75560 25048
rect 76024 24795 76084 25157
rect 76514 25010 76578 25256
rect 77530 25256 77546 25292
rect 77580 25798 77588 25832
rect 78550 25832 78610 25982
rect 79060 25931 79120 26293
rect 78846 25925 79334 25931
rect 78846 25891 78858 25925
rect 79322 25891 79334 25925
rect 78846 25885 79334 25891
rect 78550 25806 78564 25832
rect 77580 25292 77586 25798
rect 77580 25290 77590 25292
rect 77580 25256 77594 25290
rect 77042 25203 77102 25206
rect 76810 25197 77298 25203
rect 76810 25163 76822 25197
rect 77286 25163 77298 25197
rect 76810 25157 77298 25163
rect 76348 24946 76354 25010
rect 76418 24946 76578 25010
rect 76510 24842 76516 24902
rect 76576 24842 76582 24902
rect 75792 24789 76280 24795
rect 75792 24755 75804 24789
rect 76268 24755 76280 24789
rect 75792 24749 76280 24755
rect 74526 24144 74532 24650
rect 75496 24648 75510 24696
rect 75504 24146 75510 24648
rect 74526 24120 74540 24144
rect 73756 24061 74244 24067
rect 73756 24027 73768 24061
rect 74232 24027 74244 24061
rect 73756 24021 74244 24027
rect 73454 23910 73460 23970
rect 73520 23910 73526 23970
rect 74476 23860 74540 24120
rect 75496 24120 75510 24146
rect 75544 24648 75560 24696
rect 76516 24696 76576 24842
rect 77042 24795 77102 25157
rect 77530 25108 77594 25256
rect 78558 25256 78564 25806
rect 78598 25806 78610 25832
rect 79566 25832 79630 26392
rect 80588 26392 80600 26430
rect 80634 26430 80640 26968
rect 81608 26968 81668 27122
rect 82112 27067 82172 27364
rect 82614 27230 82620 27290
rect 82680 27230 82686 27290
rect 81900 27061 82388 27067
rect 81900 27027 81912 27061
rect 82376 27027 82388 27061
rect 81900 27021 82388 27027
rect 81608 26930 81618 26968
rect 81612 26432 81618 26930
rect 80634 26392 80648 26430
rect 80076 26339 80136 26345
rect 79864 26333 80352 26339
rect 79864 26299 79876 26333
rect 80340 26299 80352 26333
rect 79864 26293 80352 26299
rect 80076 25931 80136 26293
rect 80588 26246 80648 26392
rect 81604 26392 81618 26432
rect 81652 26930 81668 26968
rect 82620 26968 82680 27230
rect 83124 27067 83184 27364
rect 83640 27182 83700 27540
rect 84146 27364 84152 27424
rect 84212 27364 84218 27424
rect 85158 27364 85164 27424
rect 85224 27364 85230 27424
rect 83634 27122 83640 27182
rect 83700 27122 83706 27182
rect 82918 27061 83406 27067
rect 82918 27027 82930 27061
rect 83394 27027 83406 27061
rect 82918 27021 83406 27027
rect 81652 26432 81658 26930
rect 82620 26926 82636 26968
rect 81652 26392 81668 26432
rect 82630 26424 82636 26926
rect 81088 26339 81148 26345
rect 80882 26333 81370 26339
rect 80882 26299 80894 26333
rect 81358 26299 81370 26333
rect 80882 26293 81370 26299
rect 80582 26186 80588 26246
rect 80648 26186 80654 26246
rect 80580 25982 80586 26042
rect 80646 25982 80652 26042
rect 79864 25925 80352 25931
rect 79864 25891 79876 25925
rect 80340 25891 80352 25925
rect 79864 25885 80352 25891
rect 80076 25882 80136 25885
rect 78598 25256 78604 25806
rect 79566 25800 79582 25832
rect 79576 25304 79582 25800
rect 78558 25244 78604 25256
rect 79568 25256 79582 25304
rect 79616 25800 79630 25832
rect 80586 25832 80646 25982
rect 81088 25931 81148 26293
rect 80882 25925 81370 25931
rect 80882 25891 80894 25925
rect 81358 25891 81370 25925
rect 80882 25885 81370 25891
rect 81088 25882 81148 25885
rect 80586 25800 80600 25832
rect 79616 25304 79622 25800
rect 79616 25302 79628 25304
rect 79616 25256 79632 25302
rect 80594 25286 80600 25800
rect 78042 25203 78102 25210
rect 77828 25197 78316 25203
rect 77828 25163 77840 25197
rect 78304 25163 78316 25197
rect 77828 25157 78316 25163
rect 78846 25197 79334 25203
rect 78846 25163 78858 25197
rect 79322 25163 79334 25197
rect 78846 25157 79334 25163
rect 77524 25048 77530 25108
rect 77590 25048 77596 25108
rect 76810 24789 77298 24795
rect 76810 24755 76822 24789
rect 77286 24755 77298 24789
rect 76810 24749 77298 24755
rect 77042 24748 77102 24749
rect 76516 24660 76528 24696
rect 75544 24146 75550 24648
rect 76522 24168 76528 24660
rect 75544 24144 75556 24146
rect 75544 24120 75560 24144
rect 74774 24061 75262 24067
rect 74774 24027 74786 24061
rect 75250 24027 75262 24061
rect 74774 24021 75262 24027
rect 74470 23796 74476 23860
rect 74540 23796 74546 23860
rect 72432 23658 72438 23722
rect 72502 23658 72508 23722
rect 72262 23572 72322 23578
rect 71274 23512 71280 23572
rect 71340 23512 71346 23572
rect 71866 23236 71926 23242
rect 71150 23054 71812 23114
rect 70526 21970 70806 22030
rect 70992 21978 70998 22038
rect 71058 21978 71064 22038
rect 70402 21931 70490 21937
rect 70402 21897 70414 21931
rect 70478 21897 70490 21931
rect 70402 21891 70490 21897
rect 70136 21462 70142 21810
rect 70096 21450 70142 21462
rect 70306 21462 70320 21838
rect 70354 21462 70366 21838
rect 70526 21838 70586 21970
rect 70634 21937 70694 21970
rect 70620 21931 70708 21937
rect 70620 21897 70632 21931
rect 70696 21897 70708 21931
rect 70620 21891 70708 21897
rect 70526 21814 70538 21838
rect 70532 21508 70538 21814
rect 69966 21403 70054 21409
rect 69966 21369 69978 21403
rect 70042 21369 70054 21403
rect 69966 21363 70054 21369
rect 70184 21403 70272 21409
rect 70184 21369 70196 21403
rect 70260 21369 70272 21403
rect 70184 21363 70272 21369
rect 70306 21220 70366 21462
rect 70524 21462 70538 21508
rect 70572 21814 70586 21838
rect 70746 21838 70806 21970
rect 70572 21508 70578 21814
rect 70746 21806 70756 21838
rect 70572 21462 70584 21508
rect 70402 21403 70490 21409
rect 70402 21369 70414 21403
rect 70478 21369 70490 21403
rect 70402 21363 70490 21369
rect 70414 21326 70474 21363
rect 70524 21326 70584 21462
rect 70750 21462 70756 21806
rect 70790 21806 70806 21838
rect 70790 21462 70796 21806
rect 70750 21450 70796 21462
rect 70620 21403 70708 21409
rect 70620 21369 70632 21403
rect 70696 21369 70708 21403
rect 70620 21363 70708 21369
rect 70408 21266 70414 21326
rect 70474 21266 70480 21326
rect 70518 21266 70524 21326
rect 70584 21266 70590 21326
rect 68992 21160 68998 21220
rect 69058 21160 69064 21220
rect 69428 21160 69434 21220
rect 69494 21160 69500 21220
rect 69866 21160 69872 21220
rect 69932 21160 69938 21220
rect 70300 21160 70306 21220
rect 70366 21160 70372 21220
rect 68566 21042 68842 21102
rect 68566 20900 68626 21042
rect 68670 20999 68730 21042
rect 68658 20993 68746 20999
rect 68658 20959 68670 20993
rect 68734 20959 68746 20993
rect 68658 20953 68746 20959
rect 68566 20866 68576 20900
rect 68570 20524 68576 20866
rect 68610 20866 68626 20900
rect 68782 20900 68842 21042
rect 68876 20993 68964 20999
rect 68876 20959 68888 20993
rect 68952 20959 68964 20993
rect 68876 20953 68964 20959
rect 68782 20870 68794 20900
rect 68610 20524 68616 20866
rect 68788 20558 68794 20870
rect 68570 20512 68616 20524
rect 68782 20524 68794 20558
rect 68828 20870 68842 20900
rect 68998 20900 69058 21160
rect 69212 21044 69218 21104
rect 69278 21044 69284 21104
rect 69094 20993 69182 20999
rect 69094 20959 69106 20993
rect 69170 20959 69182 20993
rect 69094 20953 69182 20959
rect 68998 20872 69012 20900
rect 68828 20558 68834 20870
rect 69006 20566 69012 20872
rect 68828 20524 68842 20558
rect 68658 20465 68746 20471
rect 68658 20431 68670 20465
rect 68734 20431 68746 20465
rect 68658 20425 68746 20431
rect 68782 20380 68842 20524
rect 68998 20524 69012 20566
rect 69046 20872 69058 20900
rect 69218 20900 69278 21044
rect 69312 20993 69400 20999
rect 69312 20959 69324 20993
rect 69388 20959 69400 20993
rect 69312 20953 69400 20959
rect 69218 20874 69230 20900
rect 69046 20566 69052 20872
rect 69046 20524 69058 20566
rect 68876 20465 68964 20471
rect 68876 20431 68888 20465
rect 68952 20431 68964 20465
rect 68876 20425 68964 20431
rect 68776 20320 68782 20380
rect 68842 20320 68848 20380
rect 68892 20182 68952 20425
rect 68998 20276 69058 20524
rect 69224 20524 69230 20874
rect 69264 20874 69278 20900
rect 69434 20900 69494 21160
rect 69530 20993 69618 20999
rect 69530 20959 69542 20993
rect 69606 20959 69618 20993
rect 69530 20953 69618 20959
rect 69748 20993 69836 20999
rect 69748 20959 69760 20993
rect 69824 20959 69836 20993
rect 69748 20953 69836 20959
rect 69264 20524 69270 20874
rect 69434 20870 69448 20900
rect 69442 20556 69448 20870
rect 69224 20512 69270 20524
rect 69434 20524 69448 20556
rect 69482 20870 69494 20900
rect 69660 20900 69706 20912
rect 69482 20556 69488 20870
rect 69660 20560 69666 20900
rect 69482 20524 69494 20556
rect 69094 20465 69182 20471
rect 69094 20431 69106 20465
rect 69170 20431 69182 20465
rect 69094 20425 69182 20431
rect 69312 20465 69400 20471
rect 69312 20431 69324 20465
rect 69388 20431 69400 20465
rect 69312 20425 69400 20431
rect 68992 20216 68998 20276
rect 69058 20216 69064 20276
rect 68564 20178 68952 20182
rect 68564 20122 68892 20178
rect 68564 19962 68624 20122
rect 68670 20061 68730 20122
rect 68658 20055 68746 20061
rect 68658 20021 68670 20055
rect 68734 20021 68746 20055
rect 68658 20015 68746 20021
rect 68564 19936 68576 19962
rect 68570 19586 68576 19936
rect 68610 19936 68624 19962
rect 68784 19962 68844 20122
rect 68886 20118 68892 20122
rect 68952 20118 68958 20178
rect 68892 20061 68952 20118
rect 68876 20055 68964 20061
rect 68876 20021 68888 20055
rect 68952 20021 68964 20055
rect 68876 20015 68964 20021
rect 68610 19586 68616 19936
rect 68784 19924 68794 19962
rect 68788 19612 68794 19924
rect 68570 19574 68616 19586
rect 68782 19586 68794 19612
rect 68828 19924 68844 19962
rect 68998 19962 69058 20216
rect 69106 20178 69166 20425
rect 69210 20320 69216 20380
rect 69276 20320 69282 20380
rect 69100 20118 69106 20178
rect 69166 20118 69172 20178
rect 69106 20061 69166 20118
rect 69094 20055 69182 20061
rect 69094 20021 69106 20055
rect 69170 20021 69182 20055
rect 69094 20015 69182 20021
rect 68998 19928 69012 19962
rect 68828 19612 68834 19924
rect 68828 19586 68842 19612
rect 69006 19610 69012 19928
rect 68658 19527 68746 19533
rect 68658 19493 68670 19527
rect 68734 19493 68746 19527
rect 68658 19487 68746 19493
rect 68442 19226 68502 19482
rect 68782 19442 68842 19586
rect 68998 19586 69012 19610
rect 69046 19928 69058 19962
rect 69216 19962 69276 20320
rect 69326 20178 69386 20425
rect 69434 20276 69494 20524
rect 69652 20524 69666 20560
rect 69700 20560 69706 20900
rect 69872 20900 69932 21160
rect 70082 21044 70088 21104
rect 70148 21044 70154 21104
rect 69966 20993 70054 20999
rect 69966 20959 69978 20993
rect 70042 20959 70054 20993
rect 69966 20953 70054 20959
rect 69872 20866 69884 20900
rect 69700 20524 69712 20560
rect 69878 20552 69884 20866
rect 69530 20465 69618 20471
rect 69530 20431 69542 20465
rect 69606 20431 69618 20465
rect 69530 20425 69618 20431
rect 69428 20216 69434 20276
rect 69494 20216 69500 20276
rect 69320 20118 69326 20178
rect 69386 20118 69392 20178
rect 69326 20061 69386 20118
rect 69312 20055 69400 20061
rect 69312 20021 69324 20055
rect 69388 20021 69400 20055
rect 69312 20015 69400 20021
rect 69216 19928 69230 19962
rect 69046 19610 69052 19928
rect 69046 19586 69058 19610
rect 68876 19527 68964 19533
rect 68876 19493 68888 19527
rect 68952 19493 68964 19527
rect 68876 19487 68964 19493
rect 68776 19382 68782 19442
rect 68842 19382 68848 19442
rect 68998 19344 69058 19586
rect 69224 19586 69230 19928
rect 69264 19928 69276 19962
rect 69434 19962 69494 20216
rect 69544 20178 69604 20425
rect 69652 20380 69712 20524
rect 69872 20524 69884 20552
rect 69918 20866 69932 20900
rect 70088 20900 70148 21044
rect 70184 20993 70272 20999
rect 70184 20959 70196 20993
rect 70260 20959 70272 20993
rect 70184 20953 70272 20959
rect 70088 20868 70102 20900
rect 69918 20552 69924 20866
rect 69918 20524 69932 20552
rect 69748 20465 69836 20471
rect 69748 20431 69760 20465
rect 69824 20431 69836 20465
rect 69748 20425 69836 20431
rect 69646 20320 69652 20380
rect 69712 20320 69718 20380
rect 69760 20178 69820 20425
rect 69872 20276 69932 20524
rect 70096 20524 70102 20868
rect 70136 20868 70148 20900
rect 70306 20900 70366 21160
rect 70526 21060 70806 21120
rect 70402 20993 70490 20999
rect 70402 20959 70414 20993
rect 70478 20959 70490 20993
rect 70402 20953 70490 20959
rect 70306 20878 70320 20900
rect 70136 20524 70142 20868
rect 70314 20554 70320 20878
rect 70096 20512 70142 20524
rect 70306 20524 70320 20554
rect 70354 20878 70366 20900
rect 70526 20900 70586 21060
rect 70636 20999 70696 21060
rect 70620 20993 70708 20999
rect 70620 20959 70632 20993
rect 70696 20959 70708 20993
rect 70620 20953 70708 20959
rect 70354 20554 70360 20878
rect 70526 20876 70538 20900
rect 70532 20560 70538 20876
rect 70354 20524 70366 20554
rect 69966 20465 70054 20471
rect 69966 20431 69978 20465
rect 70042 20431 70054 20465
rect 69966 20425 70054 20431
rect 70184 20465 70272 20471
rect 70184 20431 70196 20465
rect 70260 20431 70272 20465
rect 70184 20425 70272 20431
rect 69866 20216 69872 20276
rect 69932 20216 69938 20276
rect 69538 20118 69544 20178
rect 69604 20118 69610 20178
rect 69648 20118 69654 20178
rect 69714 20118 69720 20178
rect 69754 20118 69760 20178
rect 69820 20118 69826 20178
rect 69544 20061 69604 20118
rect 69530 20055 69618 20061
rect 69530 20021 69542 20055
rect 69606 20021 69618 20055
rect 69530 20015 69618 20021
rect 69264 19586 69270 19928
rect 69434 19926 69448 19962
rect 69442 19624 69448 19926
rect 69224 19574 69270 19586
rect 69434 19586 69448 19624
rect 69482 19926 69494 19962
rect 69654 19962 69714 20118
rect 69760 20061 69820 20118
rect 69748 20055 69836 20061
rect 69748 20021 69760 20055
rect 69824 20021 69836 20055
rect 69748 20015 69836 20021
rect 69654 19934 69666 19962
rect 69482 19624 69488 19926
rect 69482 19586 69494 19624
rect 69660 19616 69666 19934
rect 69094 19527 69182 19533
rect 69094 19493 69106 19527
rect 69170 19493 69182 19527
rect 69094 19487 69182 19493
rect 69312 19527 69400 19533
rect 69312 19493 69324 19527
rect 69388 19493 69400 19527
rect 69312 19487 69400 19493
rect 69434 19344 69494 19586
rect 69652 19586 69666 19616
rect 69700 19934 69714 19962
rect 69872 19962 69932 20216
rect 69978 20178 70038 20425
rect 70082 20320 70088 20380
rect 70148 20320 70154 20380
rect 69972 20118 69978 20178
rect 70038 20118 70044 20178
rect 69978 20061 70038 20118
rect 69966 20055 70054 20061
rect 69966 20021 69978 20055
rect 70042 20021 70054 20055
rect 69966 20015 70054 20021
rect 69700 19616 69706 19934
rect 69872 19922 69884 19962
rect 69878 19620 69884 19922
rect 69700 19586 69712 19616
rect 69530 19527 69618 19533
rect 69530 19493 69542 19527
rect 69606 19493 69618 19527
rect 69530 19487 69618 19493
rect 69652 19442 69712 19586
rect 69872 19586 69884 19620
rect 69918 19922 69932 19962
rect 70088 19962 70148 20320
rect 70196 20178 70256 20425
rect 70306 20276 70366 20524
rect 70526 20524 70538 20560
rect 70572 20876 70586 20900
rect 70746 20900 70806 21060
rect 70876 21044 70882 21104
rect 70942 21044 70948 21104
rect 70572 20560 70578 20876
rect 70746 20864 70756 20900
rect 70572 20524 70586 20560
rect 70402 20465 70490 20471
rect 70402 20431 70414 20465
rect 70478 20431 70490 20465
rect 70402 20425 70490 20431
rect 70300 20216 70306 20276
rect 70366 20216 70372 20276
rect 70190 20118 70196 20178
rect 70256 20118 70262 20178
rect 70196 20061 70256 20118
rect 70184 20055 70272 20061
rect 70184 20021 70196 20055
rect 70260 20021 70272 20055
rect 70184 20015 70272 20021
rect 70088 19936 70102 19962
rect 69918 19620 69924 19922
rect 69918 19586 69932 19620
rect 69748 19527 69836 19533
rect 69748 19493 69760 19527
rect 69824 19493 69836 19527
rect 69748 19487 69836 19493
rect 69646 19382 69652 19442
rect 69712 19382 69718 19442
rect 69872 19344 69932 19586
rect 70096 19586 70102 19936
rect 70136 19936 70148 19962
rect 70306 19962 70366 20216
rect 70412 20178 70472 20425
rect 70526 20380 70586 20524
rect 70750 20524 70756 20864
rect 70790 20864 70806 20900
rect 70790 20524 70796 20864
rect 70750 20512 70796 20524
rect 70620 20465 70708 20471
rect 70620 20431 70632 20465
rect 70696 20431 70708 20465
rect 70620 20425 70708 20431
rect 70520 20320 70526 20380
rect 70586 20320 70592 20380
rect 70406 20118 70412 20178
rect 70472 20118 70806 20178
rect 70412 20061 70472 20118
rect 70402 20055 70490 20061
rect 70402 20021 70414 20055
rect 70478 20021 70490 20055
rect 70402 20015 70490 20021
rect 70136 19586 70142 19936
rect 70306 19934 70320 19962
rect 70314 19620 70320 19934
rect 70096 19574 70142 19586
rect 70306 19586 70320 19620
rect 70354 19934 70366 19962
rect 70524 19962 70584 20118
rect 70632 20061 70692 20118
rect 70620 20055 70708 20061
rect 70620 20021 70632 20055
rect 70696 20021 70708 20055
rect 70620 20015 70708 20021
rect 70524 19944 70538 19962
rect 70354 19620 70360 19934
rect 70532 19620 70538 19944
rect 70354 19586 70366 19620
rect 69966 19527 70054 19533
rect 69966 19493 69978 19527
rect 70042 19493 70054 19527
rect 69966 19487 70054 19493
rect 70184 19527 70272 19533
rect 70184 19493 70196 19527
rect 70260 19493 70272 19527
rect 70184 19487 70272 19493
rect 70306 19344 70366 19586
rect 70526 19586 70538 19620
rect 70572 19944 70584 19962
rect 70746 19962 70806 20118
rect 70572 19620 70578 19944
rect 70746 19940 70756 19962
rect 70572 19586 70586 19620
rect 70402 19527 70490 19533
rect 70402 19493 70414 19527
rect 70478 19493 70490 19527
rect 70402 19487 70490 19493
rect 70526 19442 70586 19586
rect 70750 19586 70756 19940
rect 70790 19940 70806 19962
rect 70790 19586 70796 19940
rect 70750 19574 70796 19586
rect 70620 19527 70708 19533
rect 70620 19493 70632 19527
rect 70696 19493 70708 19527
rect 70620 19487 70708 19493
rect 70882 19442 70942 21044
rect 70520 19382 70526 19442
rect 70586 19382 70592 19442
rect 70876 19382 70882 19442
rect 70942 19382 70948 19442
rect 68992 19284 68998 19344
rect 69058 19284 69064 19344
rect 69428 19284 69434 19344
rect 69494 19284 69500 19344
rect 69866 19284 69872 19344
rect 69932 19284 69938 19344
rect 70300 19284 70306 19344
rect 70366 19284 70372 19344
rect 68436 19166 68442 19226
rect 68502 19166 68508 19226
rect 68566 19164 68952 19224
rect 68566 19024 68626 19164
rect 68672 19123 68732 19164
rect 68658 19117 68746 19123
rect 68658 19083 68670 19117
rect 68734 19083 68746 19117
rect 68658 19077 68746 19083
rect 68566 18994 68576 19024
rect 68570 18648 68576 18994
rect 68610 18994 68626 19024
rect 68782 19024 68842 19164
rect 68892 19123 68952 19164
rect 68876 19117 68964 19123
rect 68876 19083 68888 19117
rect 68952 19083 68964 19117
rect 68876 19077 68964 19083
rect 68782 19000 68794 19024
rect 68610 18648 68616 18994
rect 68788 18676 68794 19000
rect 68570 18636 68616 18648
rect 68782 18648 68794 18676
rect 68828 19000 68842 19024
rect 68998 19024 69058 19284
rect 69102 19166 69108 19226
rect 69168 19166 69174 19226
rect 69210 19166 69216 19226
rect 69276 19166 69282 19226
rect 69318 19166 69324 19226
rect 69384 19166 69390 19226
rect 69108 19123 69168 19166
rect 69094 19117 69182 19123
rect 69094 19083 69106 19117
rect 69170 19083 69182 19117
rect 69094 19077 69182 19083
rect 68828 18676 68834 19000
rect 68998 18996 69012 19024
rect 68828 18648 68842 18676
rect 68658 18589 68746 18595
rect 68658 18555 68670 18589
rect 68734 18555 68746 18589
rect 68658 18549 68746 18555
rect 68782 18506 68842 18648
rect 69006 18648 69012 18996
rect 69046 18996 69058 19024
rect 69216 19024 69276 19166
rect 69324 19123 69384 19166
rect 69312 19117 69400 19123
rect 69312 19083 69324 19117
rect 69388 19083 69400 19117
rect 69312 19077 69400 19083
rect 69216 19000 69230 19024
rect 69046 18648 69052 18996
rect 69006 18636 69052 18648
rect 69224 18648 69230 19000
rect 69264 19000 69276 19024
rect 69434 19024 69494 19284
rect 69530 19117 69618 19123
rect 69530 19083 69542 19117
rect 69606 19083 69618 19117
rect 69530 19077 69618 19083
rect 69748 19117 69836 19123
rect 69748 19083 69760 19117
rect 69824 19083 69836 19117
rect 69748 19077 69836 19083
rect 69264 18648 69270 19000
rect 69434 18994 69448 19024
rect 69224 18636 69270 18648
rect 69442 18648 69448 18994
rect 69482 18994 69494 19024
rect 69660 19024 69706 19036
rect 69482 18648 69488 18994
rect 69660 18678 69666 19024
rect 69442 18636 69488 18648
rect 69652 18648 69666 18678
rect 69700 18678 69706 19024
rect 69872 19024 69932 19284
rect 69964 19166 69970 19226
rect 70030 19166 70036 19226
rect 70082 19166 70088 19226
rect 70148 19166 70154 19226
rect 70191 19166 70197 19224
rect 70255 19166 70261 19224
rect 69970 19123 70030 19166
rect 69966 19117 70054 19123
rect 69966 19083 69978 19117
rect 70042 19083 70054 19117
rect 69966 19077 70054 19083
rect 69872 18990 69884 19024
rect 69700 18648 69712 18678
rect 68876 18589 68964 18595
rect 68876 18555 68888 18589
rect 68952 18555 68964 18589
rect 68876 18549 68964 18555
rect 69094 18589 69182 18595
rect 69094 18555 69106 18589
rect 69170 18555 69182 18589
rect 69094 18549 69182 18555
rect 69312 18589 69400 18595
rect 69312 18555 69324 18589
rect 69388 18555 69400 18589
rect 69312 18549 69400 18555
rect 69530 18589 69618 18595
rect 69530 18555 69542 18589
rect 69606 18555 69618 18589
rect 69530 18549 69618 18555
rect 68892 18506 68952 18549
rect 69546 18506 69606 18549
rect 69652 18506 69712 18648
rect 69878 18648 69884 18990
rect 69918 18990 69932 19024
rect 70088 19024 70148 19166
rect 70197 19123 70255 19166
rect 70184 19117 70272 19123
rect 70184 19083 70196 19117
rect 70260 19083 70272 19117
rect 70184 19077 70272 19083
rect 69918 18648 69924 18990
rect 70088 18984 70102 19024
rect 69878 18636 69924 18648
rect 70096 18648 70102 18984
rect 70136 18984 70148 19024
rect 70306 19024 70366 19284
rect 70526 19174 70806 19234
rect 70402 19117 70490 19123
rect 70402 19083 70414 19117
rect 70478 19083 70490 19117
rect 70402 19077 70490 19083
rect 70306 19002 70320 19024
rect 70136 18648 70142 18984
rect 70096 18636 70142 18648
rect 70314 18648 70320 19002
rect 70354 19002 70366 19024
rect 70526 19024 70586 19174
rect 70632 19123 70692 19174
rect 70620 19117 70708 19123
rect 70620 19083 70632 19117
rect 70696 19083 70708 19117
rect 70620 19077 70708 19083
rect 70354 18648 70360 19002
rect 70526 19000 70538 19024
rect 70532 18682 70538 19000
rect 70314 18636 70360 18648
rect 70526 18648 70538 18682
rect 70572 19000 70586 19024
rect 70746 19024 70806 19174
rect 70572 18682 70578 19000
rect 70746 18996 70756 19024
rect 70572 18648 70586 18682
rect 69748 18589 69836 18595
rect 69748 18555 69760 18589
rect 69824 18555 69836 18589
rect 69748 18549 69836 18555
rect 69966 18589 70054 18595
rect 69966 18555 69978 18589
rect 70042 18555 70054 18589
rect 69966 18549 70054 18555
rect 70184 18589 70272 18595
rect 70184 18555 70196 18589
rect 70260 18555 70272 18589
rect 70184 18549 70272 18555
rect 70402 18589 70490 18595
rect 70402 18555 70414 18589
rect 70478 18555 70490 18589
rect 70402 18549 70490 18555
rect 69762 18506 69822 18549
rect 70414 18506 70474 18549
rect 70526 18506 70586 18648
rect 70750 18648 70756 18996
rect 70790 18996 70806 19024
rect 70790 18648 70796 18996
rect 70750 18636 70796 18648
rect 70620 18589 70708 18595
rect 70620 18555 70632 18589
rect 70696 18555 70708 18589
rect 70620 18549 70708 18555
rect 70998 18506 71058 21978
rect 71752 20932 71812 23054
rect 71746 20872 71752 20932
rect 71812 20872 71818 20932
rect 71866 20828 71926 23176
rect 72262 23136 72322 23512
rect 74476 23426 74540 23796
rect 74982 23788 75042 24021
rect 75496 23970 75560 24120
rect 76514 24120 76528 24168
rect 76562 24660 76576 24696
rect 77530 24696 77594 25048
rect 78042 24795 78102 25157
rect 79070 24795 79130 25157
rect 79568 25106 79632 25256
rect 80588 25256 80600 25286
rect 80634 25800 80646 25832
rect 81604 25832 81668 26392
rect 82622 26392 82636 26424
rect 82670 26926 82680 26968
rect 83640 26968 83700 27122
rect 84152 27067 84212 27364
rect 85164 27067 85224 27364
rect 85676 27182 85736 27540
rect 86176 27364 86182 27424
rect 86242 27364 86248 27424
rect 85670 27122 85676 27182
rect 85736 27122 85742 27182
rect 83936 27061 84424 27067
rect 83936 27027 83948 27061
rect 84412 27027 84424 27061
rect 83936 27021 84424 27027
rect 84954 27061 85442 27067
rect 84954 27027 84966 27061
rect 85430 27027 85442 27061
rect 84954 27021 85442 27027
rect 83640 26940 83654 26968
rect 82670 26424 82676 26926
rect 83648 26440 83654 26940
rect 82670 26392 82682 26424
rect 82094 26339 82154 26345
rect 81900 26333 82388 26339
rect 81900 26299 81912 26333
rect 82376 26299 82388 26333
rect 81900 26293 82388 26299
rect 82094 25931 82154 26293
rect 82622 26240 82682 26392
rect 83640 26392 83654 26440
rect 83688 26940 83700 26968
rect 84666 26968 84712 26980
rect 83688 26440 83694 26940
rect 83688 26392 83700 26440
rect 84666 26424 84672 26968
rect 83112 26339 83172 26345
rect 82918 26333 83406 26339
rect 82918 26299 82930 26333
rect 83394 26299 83406 26333
rect 82918 26293 83406 26299
rect 82622 26180 82824 26240
rect 82616 26082 82622 26142
rect 82682 26082 82688 26142
rect 81900 25925 82388 25931
rect 81900 25891 81912 25925
rect 82376 25891 82388 25925
rect 81900 25885 82388 25891
rect 82094 25882 82154 25885
rect 80634 25286 80640 25800
rect 81604 25784 81618 25832
rect 81612 25300 81618 25784
rect 80634 25256 80648 25286
rect 80088 25203 80148 25215
rect 79864 25197 80352 25203
rect 79864 25163 79876 25197
rect 80340 25163 80352 25197
rect 79864 25157 80352 25163
rect 79562 25046 79568 25106
rect 79628 25046 79634 25106
rect 77828 24789 78316 24795
rect 77828 24755 77840 24789
rect 78304 24755 78316 24789
rect 77828 24749 78316 24755
rect 78846 24789 79334 24795
rect 78846 24755 78858 24789
rect 79322 24755 79334 24789
rect 78846 24749 79334 24755
rect 79070 24742 79130 24749
rect 76562 24168 76568 24660
rect 77530 24636 77546 24696
rect 76562 24120 76574 24168
rect 77540 24154 77546 24636
rect 75792 24061 76280 24067
rect 75792 24027 75804 24061
rect 76268 24027 76280 24061
rect 75792 24021 76280 24027
rect 75490 23910 75496 23970
rect 75556 23910 75562 23970
rect 76024 23788 76084 24021
rect 74982 23728 76084 23788
rect 74470 23362 74476 23426
rect 74540 23362 74546 23426
rect 74982 23324 75042 23728
rect 74444 23264 75042 23324
rect 72256 23076 72262 23136
rect 72322 23076 72328 23136
rect 73422 23076 73428 23136
rect 73488 23076 73494 23136
rect 71988 22030 71994 22090
rect 72054 22030 72060 22090
rect 71860 20768 71866 20828
rect 71926 20768 71932 20828
rect 68776 18446 68782 18506
rect 68842 18446 68848 18506
rect 68886 18446 68892 18506
rect 68952 18446 68958 18506
rect 69540 18446 69546 18506
rect 69606 18446 69612 18506
rect 69646 18446 69652 18506
rect 69712 18446 69718 18506
rect 69756 18446 69762 18506
rect 69822 18446 69828 18506
rect 70408 18446 70414 18506
rect 70474 18446 70480 18506
rect 70520 18446 70526 18506
rect 70586 18446 70592 18506
rect 70992 18446 70998 18506
rect 71058 18446 71064 18506
rect 71994 18418 72054 22030
rect 72124 21932 72130 21992
rect 72190 21932 72196 21992
rect 71988 18358 71994 18418
rect 72054 18358 72060 18418
rect 72130 18288 72190 21932
rect 72262 19468 72322 23076
rect 72706 23015 73194 23021
rect 72706 22981 72718 23015
rect 73182 22981 73194 23015
rect 72706 22975 73194 22981
rect 72418 22922 72464 22934
rect 72418 22382 72424 22922
rect 72410 22346 72424 22382
rect 72458 22382 72464 22922
rect 73428 22922 73488 23076
rect 73724 23015 74212 23021
rect 73724 22981 73736 23015
rect 74200 22981 74212 23015
rect 73724 22975 74212 22981
rect 73428 22896 73442 22922
rect 72458 22346 72470 22382
rect 73436 22370 73442 22896
rect 72410 22188 72470 22346
rect 73426 22346 73442 22370
rect 73476 22896 73488 22922
rect 74444 22922 74504 23264
rect 76514 23236 76574 24120
rect 77530 24120 77546 24154
rect 77580 24636 77594 24696
rect 78558 24696 78604 24708
rect 77580 24154 77586 24636
rect 77580 24152 77590 24154
rect 78558 24152 78564 24696
rect 77580 24120 77594 24152
rect 76810 24061 77298 24067
rect 76810 24027 76822 24061
rect 77286 24027 77298 24061
rect 76810 24021 77298 24027
rect 77530 23974 77594 24120
rect 78548 24120 78564 24152
rect 78598 24152 78604 24696
rect 79568 24696 79632 25046
rect 80088 24795 80148 25157
rect 80588 25008 80648 25256
rect 81604 25256 81618 25300
rect 81652 25784 81668 25832
rect 82622 25832 82682 26082
rect 82764 26038 82824 26180
rect 82758 25978 82764 26038
rect 82824 25978 82830 26038
rect 83112 25931 83172 26293
rect 82918 25925 83406 25931
rect 82918 25891 82930 25925
rect 83394 25891 83406 25925
rect 82918 25885 83406 25891
rect 83112 25882 83172 25885
rect 82622 25808 82636 25832
rect 81652 25300 81658 25784
rect 81652 25298 81664 25300
rect 81652 25256 81668 25298
rect 81088 25203 81148 25211
rect 80882 25197 81370 25203
rect 80882 25163 80894 25197
rect 81358 25163 81370 25197
rect 80882 25157 81370 25163
rect 80582 24948 80588 25008
rect 80648 24948 80654 25008
rect 81088 24795 81148 25157
rect 81604 25106 81668 25256
rect 82630 25256 82636 25808
rect 82670 25808 82682 25832
rect 83640 25832 83700 26392
rect 84656 26392 84672 26424
rect 84706 26424 84712 26968
rect 85676 26968 85736 27122
rect 86182 27067 86242 27364
rect 86696 27130 87776 27190
rect 85972 27061 86460 27067
rect 85972 27027 85984 27061
rect 86448 27027 86460 27061
rect 85972 27021 86460 27027
rect 85676 26936 85690 26968
rect 85684 26430 85690 26936
rect 84706 26392 84716 26424
rect 84130 26339 84190 26345
rect 83936 26333 84424 26339
rect 83936 26299 83948 26333
rect 84412 26299 84424 26333
rect 83936 26293 84424 26299
rect 84130 25931 84190 26293
rect 84656 26142 84716 26392
rect 85680 26392 85690 26430
rect 85724 26936 85736 26968
rect 86696 26968 86756 27130
rect 87198 27067 87258 27130
rect 86990 27061 87478 27067
rect 86990 27027 87002 27061
rect 87466 27027 87478 27061
rect 86990 27021 87478 27027
rect 86696 26938 86708 26968
rect 85724 26430 85730 26936
rect 86702 26432 86708 26938
rect 85724 26392 85740 26430
rect 85130 26339 85190 26345
rect 84954 26333 85442 26339
rect 84954 26299 84966 26333
rect 85430 26299 85442 26333
rect 84954 26293 85442 26299
rect 84650 26082 84656 26142
rect 84716 26082 84722 26142
rect 84652 25978 84658 26038
rect 84718 25978 84724 26038
rect 83936 25925 84424 25931
rect 83936 25891 83948 25925
rect 84412 25891 84424 25925
rect 83936 25885 84424 25891
rect 84130 25882 84190 25885
rect 82670 25256 82676 25808
rect 83640 25788 83654 25832
rect 83648 25292 83654 25788
rect 82630 25244 82676 25256
rect 83640 25256 83654 25292
rect 83688 25788 83700 25832
rect 84658 25832 84718 25978
rect 85130 25931 85190 26293
rect 84954 25925 85442 25931
rect 84954 25891 84966 25925
rect 85430 25891 85442 25925
rect 84954 25885 85442 25891
rect 85130 25882 85190 25885
rect 84658 25804 84672 25832
rect 83688 25292 83694 25788
rect 84666 25292 84672 25804
rect 83688 25256 83700 25292
rect 82094 25203 82154 25211
rect 83136 25203 83196 25211
rect 81900 25197 82388 25203
rect 81900 25163 81912 25197
rect 82376 25163 82388 25197
rect 81900 25157 82388 25163
rect 82918 25197 83406 25203
rect 82918 25163 82930 25197
rect 83394 25163 83406 25197
rect 82918 25157 83406 25163
rect 81598 25046 81604 25106
rect 81664 25046 81670 25106
rect 79864 24789 80352 24795
rect 79864 24755 79876 24789
rect 80340 24755 80352 24789
rect 79864 24749 80352 24755
rect 80882 24789 81370 24795
rect 80882 24755 80894 24789
rect 81358 24755 81370 24789
rect 80882 24749 81370 24755
rect 81088 24748 81148 24749
rect 79568 24656 79582 24696
rect 79576 24166 79582 24656
rect 78598 24120 78612 24152
rect 77828 24061 78316 24067
rect 77828 24027 77840 24061
rect 78304 24027 78316 24061
rect 77828 24021 78316 24027
rect 76990 23966 77050 23972
rect 76508 23176 76514 23236
rect 76574 23176 76580 23236
rect 75458 23076 75464 23136
rect 75524 23076 75530 23136
rect 74742 23015 75230 23021
rect 74742 22981 74754 23015
rect 75218 22981 75230 23015
rect 74742 22975 75230 22981
rect 73476 22370 73482 22896
rect 74444 22876 74460 22922
rect 74454 22370 74460 22876
rect 73476 22346 73486 22370
rect 72706 22287 73194 22293
rect 72706 22253 72718 22287
rect 73182 22253 73194 22287
rect 72706 22247 73194 22253
rect 72924 22188 72984 22247
rect 73426 22188 73486 22346
rect 74446 22346 74460 22370
rect 74494 22876 74504 22922
rect 75464 22922 75524 23076
rect 76990 23021 77050 23906
rect 77498 23970 77594 23974
rect 77498 23968 77530 23970
rect 77590 23910 77596 23970
rect 77984 23910 77990 23970
rect 78050 23910 78056 23970
rect 75760 23015 76248 23021
rect 75760 22981 75772 23015
rect 76236 22981 76248 23015
rect 75760 22975 76248 22981
rect 76778 23015 77266 23021
rect 76778 22981 76790 23015
rect 77254 22981 77266 23015
rect 76778 22975 77266 22981
rect 75464 22898 75478 22922
rect 74494 22370 74500 22876
rect 74494 22346 74506 22370
rect 73724 22287 74212 22293
rect 73724 22253 73736 22287
rect 74200 22253 74212 22287
rect 73724 22247 74212 22253
rect 72410 22128 73486 22188
rect 73426 21822 73432 21882
rect 73492 21822 73498 21882
rect 72706 21759 73194 21765
rect 72706 21725 72718 21759
rect 73182 21725 73194 21759
rect 72706 21719 73194 21725
rect 72418 21666 72464 21678
rect 72418 21126 72424 21666
rect 72414 21090 72424 21126
rect 72458 21126 72464 21666
rect 73432 21666 73492 21822
rect 73916 21765 73976 22247
rect 74446 22188 74506 22346
rect 75472 22346 75478 22898
rect 75512 22898 75524 22922
rect 76490 22922 76536 22934
rect 75512 22346 75518 22898
rect 76490 22374 76496 22922
rect 75472 22334 75518 22346
rect 76482 22346 76496 22374
rect 76530 22374 76536 22922
rect 77498 22922 77558 23908
rect 77990 23021 78050 23910
rect 78548 23722 78612 24120
rect 79568 24120 79582 24166
rect 79616 24656 79632 24696
rect 80594 24696 80640 24708
rect 79616 24166 79622 24656
rect 79616 24164 79628 24166
rect 79616 24120 79632 24164
rect 80594 24156 80600 24696
rect 78846 24061 79334 24067
rect 78846 24027 78858 24061
rect 79322 24027 79334 24061
rect 78846 24021 79334 24027
rect 79568 23978 79632 24120
rect 80584 24120 80600 24156
rect 80634 24156 80640 24696
rect 81604 24696 81668 25046
rect 82094 24795 82154 25157
rect 82616 24842 82622 24902
rect 82682 24842 82688 24902
rect 81900 24789 82388 24795
rect 81900 24755 81912 24789
rect 82376 24755 82388 24789
rect 81900 24749 82388 24755
rect 82094 24748 82154 24749
rect 81604 24644 81618 24696
rect 81612 24162 81618 24644
rect 80634 24120 80648 24156
rect 79864 24061 80352 24067
rect 79864 24027 79876 24061
rect 80340 24027 80352 24061
rect 79864 24021 80352 24027
rect 79034 23972 79094 23978
rect 78542 23658 78548 23722
rect 78612 23658 78618 23722
rect 78548 23438 78612 23658
rect 78548 23368 78612 23374
rect 79034 23021 79094 23912
rect 79536 23972 79632 23978
rect 79596 23968 79632 23972
rect 80050 23972 80110 23978
rect 79536 23908 79568 23912
rect 79628 23908 79634 23968
rect 77796 23015 78284 23021
rect 77796 22981 77808 23015
rect 78272 22981 78284 23015
rect 77796 22975 78284 22981
rect 78814 23015 79302 23021
rect 78814 22981 78826 23015
rect 79290 22981 79302 23015
rect 78814 22975 79302 22981
rect 79034 22968 79094 22975
rect 76530 22346 76542 22374
rect 74742 22287 75230 22293
rect 74742 22253 74754 22287
rect 75218 22253 75230 22287
rect 74742 22247 75230 22253
rect 75760 22287 76248 22293
rect 75760 22253 75772 22287
rect 76236 22253 76248 22287
rect 75760 22247 76248 22253
rect 74440 22128 74446 22188
rect 74506 22128 74512 22188
rect 74446 21992 74506 22128
rect 74440 21932 74446 21992
rect 74506 21932 74512 21992
rect 74954 21765 75014 22247
rect 75460 21934 75466 21994
rect 75526 21934 75532 21994
rect 75466 21882 75526 21934
rect 75460 21822 75466 21882
rect 75526 21822 75532 21882
rect 73724 21759 74212 21765
rect 73724 21725 73736 21759
rect 74200 21725 74212 21759
rect 73724 21719 74212 21725
rect 74742 21759 75230 21765
rect 74742 21725 74754 21759
rect 75218 21725 75230 21759
rect 74742 21719 75230 21725
rect 73432 21640 73442 21666
rect 72458 21090 72474 21126
rect 73436 21114 73442 21640
rect 72414 20932 72474 21090
rect 73430 21090 73442 21114
rect 73476 21640 73492 21666
rect 74454 21666 74500 21678
rect 73476 21114 73482 21640
rect 74454 21116 74460 21666
rect 73476 21090 73490 21114
rect 72706 21031 73194 21037
rect 72706 20997 72718 21031
rect 73182 20997 73194 21031
rect 72706 20991 73194 20997
rect 72928 20932 72988 20991
rect 73430 20932 73490 21090
rect 74448 21090 74460 21116
rect 74494 21116 74500 21666
rect 75466 21666 75526 21822
rect 75960 21765 76020 22247
rect 76482 22188 76542 22346
rect 77498 22346 77514 22922
rect 77548 22346 77558 22922
rect 78526 22922 78572 22934
rect 78526 22370 78532 22922
rect 76778 22287 77266 22293
rect 76778 22253 76790 22287
rect 77254 22253 77266 22287
rect 76778 22247 77266 22253
rect 76992 22192 77052 22247
rect 77498 22192 77558 22346
rect 78518 22346 78532 22370
rect 78566 22370 78572 22922
rect 79536 22922 79596 23908
rect 80050 23021 80110 23912
rect 80584 23722 80648 24120
rect 81604 24120 81618 24162
rect 81652 24644 81668 24696
rect 82622 24696 82682 24842
rect 83136 24795 83196 25157
rect 83640 25106 83700 25256
rect 84658 25256 84672 25292
rect 84706 25804 84718 25832
rect 85680 25832 85740 26392
rect 86696 26392 86708 26432
rect 86742 26938 86756 26968
rect 87716 26968 87776 27130
rect 86742 26432 86748 26938
rect 87716 26922 87726 26968
rect 86742 26392 86756 26432
rect 86160 26339 86220 26351
rect 85972 26333 86460 26339
rect 85972 26299 85984 26333
rect 86448 26299 86460 26333
rect 85972 26293 86460 26299
rect 86160 25931 86220 26293
rect 86696 26246 86756 26392
rect 87720 26392 87726 26922
rect 87760 26922 87776 26968
rect 87760 26392 87766 26922
rect 87720 26380 87766 26392
rect 86990 26333 87478 26339
rect 86990 26299 87002 26333
rect 87466 26299 87478 26333
rect 86990 26293 87478 26299
rect 86690 26186 86696 26246
rect 86756 26186 86762 26246
rect 87828 26186 87834 26246
rect 87894 26186 87900 26246
rect 86700 25970 87770 26030
rect 85972 25925 86460 25931
rect 85972 25891 85984 25925
rect 86448 25891 86460 25925
rect 85972 25885 86460 25891
rect 84706 25292 84712 25804
rect 85680 25796 85690 25832
rect 84706 25256 84718 25292
rect 85684 25288 85690 25796
rect 84136 25203 84196 25215
rect 83936 25197 84424 25203
rect 83936 25163 83948 25197
rect 84412 25163 84424 25197
rect 83936 25157 84424 25163
rect 83634 25046 83640 25106
rect 83700 25046 83706 25106
rect 82918 24789 83406 24795
rect 82918 24755 82930 24789
rect 83394 24755 83406 24789
rect 82918 24749 83406 24755
rect 83136 24748 83196 24749
rect 82622 24660 82636 24696
rect 81652 24162 81658 24644
rect 81652 24160 81664 24162
rect 81652 24120 81668 24160
rect 80882 24061 81370 24067
rect 80882 24027 80894 24061
rect 81358 24027 81370 24061
rect 80882 24021 81370 24027
rect 81078 23972 81138 23978
rect 81604 23972 81668 24120
rect 82630 24120 82636 24660
rect 82670 24660 82682 24696
rect 83640 24696 83700 25046
rect 84136 24795 84196 25157
rect 84658 24902 84718 25256
rect 85674 25256 85690 25288
rect 85724 25796 85740 25832
rect 86700 25832 86760 25970
rect 87206 25931 87266 25970
rect 86990 25925 87478 25931
rect 86990 25891 87002 25925
rect 87466 25891 87478 25925
rect 86990 25885 87478 25891
rect 86700 25804 86708 25832
rect 85724 25288 85730 25796
rect 85724 25286 85734 25288
rect 86702 25286 86708 25804
rect 85724 25256 85738 25286
rect 85162 25203 85222 25211
rect 84954 25197 85442 25203
rect 84954 25163 84966 25197
rect 85430 25163 85442 25197
rect 84954 25157 85442 25163
rect 84652 24842 84658 24902
rect 84718 24842 84724 24902
rect 85162 24795 85222 25157
rect 85674 25104 85738 25256
rect 86696 25256 86708 25286
rect 86742 25804 86760 25832
rect 87710 25832 87770 25970
rect 86742 25286 86748 25804
rect 87710 25798 87726 25832
rect 86742 25256 86756 25286
rect 86160 25203 86220 25209
rect 85972 25197 86460 25203
rect 85972 25163 85984 25197
rect 86448 25163 86460 25197
rect 85972 25157 86460 25163
rect 85668 25044 85674 25104
rect 85734 25044 85740 25104
rect 83936 24789 84424 24795
rect 83936 24755 83948 24789
rect 84412 24755 84424 24789
rect 83936 24749 84424 24755
rect 84954 24789 85442 24795
rect 84954 24755 84966 24789
rect 85430 24755 85442 24789
rect 84954 24749 85442 24755
rect 85162 24748 85222 24749
rect 82670 24120 82676 24660
rect 83640 24642 83654 24696
rect 83648 24150 83654 24642
rect 82630 24108 82676 24120
rect 83640 24120 83654 24150
rect 83688 24642 83700 24696
rect 84666 24696 84712 24708
rect 83688 24150 83694 24642
rect 84666 24154 84672 24696
rect 83688 24148 83700 24150
rect 83688 24120 83704 24148
rect 81900 24061 82388 24067
rect 81900 24027 81912 24061
rect 82376 24027 82388 24061
rect 81900 24021 82388 24027
rect 82918 24061 83406 24067
rect 82918 24027 82930 24061
rect 83394 24027 83406 24061
rect 82918 24021 83406 24027
rect 80578 23658 80584 23722
rect 80648 23658 80654 23722
rect 81078 23021 81138 23912
rect 81572 23968 81668 23972
rect 81572 23966 81604 23968
rect 81664 23908 81670 23968
rect 82100 23962 82160 23968
rect 79832 23015 80320 23021
rect 79832 22981 79844 23015
rect 80308 22981 80320 23015
rect 79832 22975 80320 22981
rect 80850 23015 81338 23021
rect 80850 22981 80862 23015
rect 81326 22981 81338 23015
rect 80850 22975 81338 22981
rect 78566 22346 78578 22370
rect 77796 22287 78284 22293
rect 77796 22253 77808 22287
rect 78272 22253 78284 22287
rect 77796 22247 78284 22253
rect 78012 22192 78072 22247
rect 78518 22192 78578 22346
rect 79536 22346 79550 22922
rect 79584 22346 79596 22922
rect 80562 22922 80608 22934
rect 80562 22372 80568 22922
rect 78814 22287 79302 22293
rect 78814 22253 78826 22287
rect 79290 22253 79302 22287
rect 78814 22247 79302 22253
rect 79022 22192 79082 22247
rect 79536 22192 79596 22346
rect 80552 22346 80568 22372
rect 80602 22372 80608 22922
rect 81572 22922 81632 23906
rect 82100 23021 82160 23902
rect 82588 23966 82648 23972
rect 81868 23015 82356 23021
rect 81868 22981 81880 23015
rect 82344 22981 82356 23015
rect 81868 22975 82356 22981
rect 82100 22974 82160 22975
rect 80602 22346 80612 22372
rect 79832 22287 80320 22293
rect 79832 22253 79844 22287
rect 80308 22253 80320 22287
rect 79832 22247 80320 22253
rect 80044 22192 80104 22247
rect 80552 22192 80612 22346
rect 81572 22346 81586 22922
rect 81620 22346 81632 22922
rect 80850 22287 81338 22293
rect 80850 22253 80862 22287
rect 81326 22253 81338 22287
rect 80850 22247 81338 22253
rect 81066 22192 81126 22247
rect 81572 22192 81632 22346
rect 82588 22922 82648 23906
rect 83100 23962 83160 23968
rect 83640 23966 83704 24120
rect 84656 24120 84672 24154
rect 84706 24154 84712 24696
rect 85674 24696 85738 25044
rect 86160 24795 86220 25157
rect 86696 25008 86756 25256
rect 87720 25256 87726 25798
rect 87760 25798 87770 25832
rect 87760 25256 87766 25798
rect 87720 25244 87766 25256
rect 86990 25197 87478 25203
rect 86990 25163 87002 25197
rect 87466 25163 87478 25197
rect 86990 25157 87478 25163
rect 86690 24948 86696 25008
rect 86756 24948 86762 25008
rect 86698 24894 86758 24896
rect 86698 24834 87770 24894
rect 85972 24789 86460 24795
rect 85972 24755 85984 24789
rect 86448 24755 86460 24789
rect 85972 24749 86460 24755
rect 86160 24746 86220 24749
rect 85674 24650 85690 24696
rect 84706 24120 84720 24154
rect 85684 24150 85690 24650
rect 83936 24061 84424 24067
rect 83936 24027 83948 24061
rect 84412 24027 84424 24061
rect 83936 24021 84424 24027
rect 83634 23906 83640 23966
rect 83700 23906 83706 23966
rect 83100 23021 83160 23902
rect 84656 23860 84720 24120
rect 85674 24120 85690 24150
rect 85724 24650 85738 24696
rect 86698 24696 86758 24834
rect 87202 24795 87262 24834
rect 86990 24789 87478 24795
rect 86990 24755 87002 24789
rect 87466 24755 87478 24789
rect 86990 24749 87478 24755
rect 86698 24670 86708 24696
rect 85724 24150 85730 24650
rect 86702 24150 86708 24670
rect 85724 24148 85734 24150
rect 85724 24120 85738 24148
rect 84954 24061 85442 24067
rect 84954 24027 84966 24061
rect 85430 24027 85442 24061
rect 84954 24021 85442 24027
rect 85674 23966 85738 24120
rect 86692 24120 86708 24150
rect 86742 24670 86758 24696
rect 87710 24696 87770 24834
rect 86742 24150 86748 24670
rect 87710 24646 87726 24696
rect 86742 24120 86756 24150
rect 85972 24061 86460 24067
rect 85972 24027 85984 24061
rect 86448 24027 86460 24061
rect 85972 24021 86460 24027
rect 85668 23906 85674 23966
rect 85734 23906 85740 23966
rect 84650 23796 84656 23860
rect 84720 23796 84726 23860
rect 86692 23722 86756 24120
rect 87720 24120 87726 24646
rect 87760 24646 87770 24696
rect 87760 24120 87766 24646
rect 87720 24108 87766 24120
rect 86990 24061 87478 24067
rect 86990 24027 87002 24061
rect 87466 24027 87478 24061
rect 86990 24021 87478 24027
rect 86686 23658 86692 23722
rect 86756 23658 86762 23722
rect 86664 23442 86724 23448
rect 86664 23140 86724 23382
rect 87834 23436 87894 26186
rect 87834 23370 87894 23376
rect 83604 23076 83610 23136
rect 83670 23076 83676 23136
rect 85638 23076 85644 23136
rect 85704 23076 85710 23136
rect 86664 23080 87740 23140
rect 82886 23015 83374 23021
rect 82886 22981 82898 23015
rect 83362 22981 83374 23015
rect 82886 22975 83374 22981
rect 83100 22968 83160 22975
rect 82588 22346 82604 22922
rect 82638 22346 82648 22922
rect 83610 22922 83670 23076
rect 83904 23015 84392 23021
rect 83904 22981 83916 23015
rect 84380 22981 84392 23015
rect 83904 22975 84392 22981
rect 84922 23015 85410 23021
rect 84922 22981 84934 23015
rect 85398 22981 85410 23015
rect 84922 22975 85410 22981
rect 83610 22894 83622 22922
rect 81868 22287 82356 22293
rect 81868 22253 81880 22287
rect 82344 22253 82356 22287
rect 81868 22247 82356 22253
rect 82092 22192 82152 22247
rect 82588 22192 82648 22346
rect 83616 22346 83622 22894
rect 83656 22894 83670 22922
rect 84634 22922 84680 22934
rect 83656 22346 83662 22894
rect 84634 22370 84640 22922
rect 83616 22334 83662 22346
rect 84626 22346 84640 22370
rect 84674 22370 84680 22922
rect 85644 22922 85704 23076
rect 85940 23015 86428 23021
rect 85940 22981 85952 23015
rect 86416 22981 86428 23015
rect 85940 22975 86428 22981
rect 85644 22898 85658 22922
rect 84674 22346 84686 22370
rect 82886 22287 83374 22293
rect 82886 22253 82898 22287
rect 83362 22253 83374 22287
rect 82886 22247 83374 22253
rect 83904 22287 84392 22293
rect 83904 22253 83916 22287
rect 84380 22253 84392 22287
rect 83904 22247 84392 22253
rect 83104 22192 83164 22247
rect 76476 22128 76482 22188
rect 76542 22128 76548 22188
rect 76992 22132 83164 22192
rect 77498 22032 77558 22132
rect 82588 22032 82648 22132
rect 77498 21972 82648 22032
rect 75760 21759 76248 21765
rect 75760 21725 75772 21759
rect 76236 21725 76248 21759
rect 75760 21719 76248 21725
rect 76778 21759 77266 21765
rect 76778 21725 76790 21759
rect 77254 21725 77266 21759
rect 76778 21719 77266 21725
rect 75466 21644 75478 21666
rect 74494 21090 74508 21116
rect 73910 21037 73970 21038
rect 73724 21031 74212 21037
rect 73724 20997 73736 21031
rect 74200 20997 74212 21031
rect 73724 20991 74212 20997
rect 72414 20872 73490 20932
rect 72412 20570 73488 20630
rect 72412 20410 72472 20570
rect 72926 20509 72986 20570
rect 72706 20503 73194 20509
rect 72706 20469 72718 20503
rect 73182 20469 73194 20503
rect 72706 20463 73194 20469
rect 72412 20376 72424 20410
rect 72418 19834 72424 20376
rect 72458 20376 72472 20410
rect 73428 20410 73488 20570
rect 73910 20509 73970 20991
rect 74448 20828 74508 21090
rect 75472 21090 75478 21644
rect 75512 21644 75526 21666
rect 76490 21666 76536 21678
rect 75512 21090 75518 21644
rect 76490 21120 76496 21666
rect 75472 21078 75518 21090
rect 76484 21090 76496 21120
rect 76530 21120 76536 21666
rect 77498 21666 77558 21972
rect 78516 21820 78522 21880
rect 78582 21820 78588 21880
rect 79026 21834 80084 21894
rect 77796 21759 78284 21765
rect 77796 21725 77808 21759
rect 78272 21725 78284 21759
rect 77796 21719 78284 21725
rect 77498 21622 77514 21666
rect 77508 21120 77514 21622
rect 76530 21090 76544 21120
rect 74948 21037 75008 21038
rect 75954 21037 76014 21038
rect 74742 21031 75230 21037
rect 74742 20997 74754 21031
rect 75218 20997 75230 21031
rect 74742 20991 75230 20997
rect 75760 21031 76248 21037
rect 75760 20997 75772 21031
rect 76236 20997 76248 21031
rect 75760 20991 76248 20997
rect 74448 20762 74508 20768
rect 74442 20564 74448 20624
rect 74508 20564 74514 20624
rect 73724 20503 74212 20509
rect 73724 20469 73736 20503
rect 74200 20469 74212 20503
rect 73724 20463 74212 20469
rect 73428 20388 73442 20410
rect 72458 19834 72464 20376
rect 73436 19862 73442 20388
rect 72418 19822 72464 19834
rect 73430 19834 73442 19862
rect 73476 20388 73488 20410
rect 74448 20410 74508 20564
rect 74948 20509 75008 20991
rect 75954 20509 76014 20991
rect 76484 20828 76544 21090
rect 77500 21090 77514 21120
rect 77548 21622 77558 21666
rect 78522 21666 78582 21820
rect 79026 21765 79086 21834
rect 80026 21796 80084 21834
rect 80550 21820 80556 21880
rect 80616 21820 80622 21880
rect 80026 21765 80086 21796
rect 78814 21759 79302 21765
rect 78814 21725 78826 21759
rect 79290 21725 79302 21759
rect 78814 21719 79302 21725
rect 79832 21759 80320 21765
rect 79832 21725 79844 21759
rect 80308 21725 80320 21759
rect 79832 21719 80320 21725
rect 78522 21638 78532 21666
rect 77548 21120 77554 21622
rect 77548 21090 77560 21120
rect 76778 21031 77266 21037
rect 76778 20997 76790 21031
rect 77254 20997 77266 21031
rect 76778 20991 77266 20997
rect 77004 20936 77064 20991
rect 77500 20936 77560 21090
rect 78526 21090 78532 21638
rect 78566 21638 78582 21666
rect 79544 21666 79590 21678
rect 78566 21090 78572 21638
rect 79544 21114 79550 21666
rect 78526 21078 78572 21090
rect 79538 21090 79550 21114
rect 79584 21114 79590 21666
rect 80556 21666 80616 21820
rect 80850 21759 81338 21765
rect 80850 21725 80862 21759
rect 81326 21725 81338 21759
rect 80850 21719 81338 21725
rect 81868 21759 82356 21765
rect 81868 21725 81880 21759
rect 82344 21725 82356 21759
rect 81868 21719 82356 21725
rect 80556 21636 80568 21666
rect 80562 21118 80568 21636
rect 79584 21090 79598 21114
rect 77796 21031 78284 21037
rect 77796 20997 77808 21031
rect 78272 20997 78284 21031
rect 77796 20991 78284 20997
rect 78814 21031 79302 21037
rect 78814 20997 78826 21031
rect 79290 20997 79302 21031
rect 78814 20991 79302 20997
rect 78016 20936 78076 20991
rect 77004 20876 78076 20936
rect 76478 20768 76484 20828
rect 76544 20768 76550 20828
rect 76476 20666 76482 20726
rect 76542 20666 76548 20726
rect 76482 20624 76542 20666
rect 76476 20564 76482 20624
rect 76542 20564 76548 20624
rect 74742 20503 75230 20509
rect 74742 20469 74754 20503
rect 75218 20469 75230 20503
rect 74742 20463 75230 20469
rect 75760 20503 76248 20509
rect 75760 20469 75772 20503
rect 76236 20469 76248 20503
rect 75760 20463 76248 20469
rect 73476 19862 73482 20388
rect 74448 20386 74460 20410
rect 73476 19834 73490 19862
rect 72706 19775 73194 19781
rect 72706 19741 72718 19775
rect 73182 19741 73194 19775
rect 72706 19735 73194 19741
rect 73430 19676 73490 19834
rect 74454 19834 74460 20386
rect 74494 20386 74508 20410
rect 75472 20410 75518 20422
rect 74494 19834 74500 20386
rect 75472 19858 75478 20410
rect 74454 19822 74500 19834
rect 75466 19834 75478 19858
rect 75512 19858 75518 20410
rect 76482 20410 76542 20564
rect 76778 20503 77266 20509
rect 76778 20469 76790 20503
rect 77254 20469 77266 20503
rect 76778 20463 77266 20469
rect 76482 20382 76496 20410
rect 75512 19834 75526 19858
rect 73922 19781 73982 19788
rect 74960 19781 75020 19788
rect 73724 19775 74212 19781
rect 73724 19741 73736 19775
rect 74200 19741 74212 19775
rect 73724 19735 74212 19741
rect 74742 19775 75230 19781
rect 74742 19741 74754 19775
rect 75218 19741 75230 19775
rect 74742 19735 75230 19741
rect 73424 19616 73430 19676
rect 73490 19616 73496 19676
rect 72256 19408 72262 19468
rect 72322 19408 72328 19468
rect 72412 19310 73488 19370
rect 72412 19154 72472 19310
rect 72926 19253 72986 19310
rect 72706 19247 73194 19253
rect 72706 19213 72718 19247
rect 73182 19213 73194 19247
rect 72706 19207 73194 19213
rect 72412 19116 72424 19154
rect 72418 18578 72424 19116
rect 72458 19116 72472 19154
rect 73428 19154 73488 19310
rect 73922 19253 73982 19735
rect 74438 19306 74444 19366
rect 74504 19306 74510 19366
rect 73724 19247 74212 19253
rect 73724 19213 73736 19247
rect 74200 19213 74212 19247
rect 73724 19207 74212 19213
rect 73428 19128 73442 19154
rect 72458 18578 72464 19116
rect 73436 18604 73442 19128
rect 72418 18566 72464 18578
rect 73426 18578 73442 18604
rect 73476 19128 73488 19154
rect 74444 19154 74504 19306
rect 74960 19253 75020 19735
rect 75466 19676 75526 19834
rect 76490 19834 76496 20382
rect 76530 20382 76542 20410
rect 77500 20410 77560 20876
rect 78512 20872 78518 20932
rect 78578 20872 78584 20932
rect 77796 20503 78284 20509
rect 77796 20469 77808 20503
rect 78272 20469 78284 20503
rect 77796 20463 78284 20469
rect 76530 19834 76536 20382
rect 77500 20372 77514 20410
rect 77508 19868 77514 20372
rect 76490 19822 76536 19834
rect 77498 19834 77514 19868
rect 77548 20372 77560 20410
rect 78518 20410 78578 20872
rect 79020 20509 79080 20991
rect 79538 20932 79598 21090
rect 80556 21090 80568 21118
rect 80602 21636 80616 21666
rect 81580 21666 81626 21678
rect 80602 21118 80608 21636
rect 81580 21118 81586 21666
rect 80602 21090 80616 21118
rect 80050 21037 80110 21044
rect 79832 21031 80320 21037
rect 79832 20997 79844 21031
rect 80308 20997 80320 21031
rect 79832 20991 80320 20997
rect 79532 20872 79538 20932
rect 79598 20872 79604 20932
rect 79532 20566 79538 20626
rect 79598 20566 79604 20626
rect 78814 20503 79302 20509
rect 78814 20469 78826 20503
rect 79290 20469 79302 20503
rect 78814 20463 79302 20469
rect 79020 20458 79080 20463
rect 78518 20386 78532 20410
rect 77548 19868 77554 20372
rect 77548 19834 77558 19868
rect 78526 19864 78532 20386
rect 75966 19781 76026 19788
rect 75760 19775 76248 19781
rect 75760 19741 75772 19775
rect 76236 19741 76248 19775
rect 75760 19735 76248 19741
rect 76778 19775 77266 19781
rect 76778 19741 76790 19775
rect 77254 19741 77266 19775
rect 76778 19735 77266 19741
rect 75460 19616 75466 19676
rect 75526 19616 75532 19676
rect 75466 19568 75526 19616
rect 75460 19508 75466 19568
rect 75526 19508 75532 19568
rect 75966 19518 76026 19735
rect 77002 19684 77062 19735
rect 77498 19684 77558 19834
rect 78520 19834 78532 19864
rect 78566 20386 78578 20410
rect 79538 20410 79598 20566
rect 80050 20509 80110 20991
rect 80556 20626 80616 21090
rect 81574 21090 81586 21118
rect 81620 21118 81626 21666
rect 82588 21666 82648 21972
rect 83606 21820 83612 21880
rect 83672 21820 83678 21880
rect 82886 21759 83374 21765
rect 82886 21725 82898 21759
rect 83362 21725 83374 21759
rect 82886 21719 83374 21725
rect 82588 21646 82604 21666
rect 82598 21118 82604 21646
rect 81620 21090 81634 21118
rect 81062 21037 81122 21044
rect 80850 21031 81338 21037
rect 80850 20997 80862 21031
rect 81326 20997 81338 21031
rect 80850 20991 81338 20997
rect 80550 20566 80556 20626
rect 80616 20566 80622 20626
rect 81062 20509 81122 20991
rect 81574 20932 81634 21090
rect 82588 21090 82604 21118
rect 82638 21646 82648 21666
rect 83612 21666 83672 21820
rect 84112 21765 84172 22247
rect 84626 22188 84686 22346
rect 85652 22346 85658 22898
rect 85692 22898 85704 22922
rect 86664 22922 86724 23080
rect 87178 23021 87238 23080
rect 86958 23015 87446 23021
rect 86958 22981 86970 23015
rect 87434 22981 87446 23015
rect 86958 22975 87446 22981
rect 85692 22346 85698 22898
rect 86664 22886 86676 22922
rect 86670 22374 86676 22886
rect 85652 22334 85698 22346
rect 86662 22346 86676 22374
rect 86710 22886 86724 22922
rect 87680 22922 87740 23080
rect 88082 23076 88088 23136
rect 88148 23076 88154 23136
rect 87680 22898 87694 22922
rect 86710 22374 86716 22886
rect 86710 22346 86722 22374
rect 86142 22293 86202 22299
rect 84922 22287 85410 22293
rect 84922 22253 84934 22287
rect 85398 22253 85410 22287
rect 84922 22247 85410 22253
rect 85940 22287 86428 22293
rect 85940 22253 85952 22287
rect 86416 22253 86428 22287
rect 85940 22247 86428 22253
rect 84620 22128 84626 22188
rect 84686 22128 84692 22188
rect 85136 21765 85196 22247
rect 85640 21820 85646 21880
rect 85706 21820 85712 21880
rect 83904 21759 84392 21765
rect 83904 21725 83916 21759
rect 84380 21725 84392 21759
rect 83904 21719 84392 21725
rect 84922 21759 85410 21765
rect 84922 21725 84934 21759
rect 85398 21725 85410 21759
rect 84922 21719 85410 21725
rect 82638 21118 82644 21646
rect 83612 21638 83622 21666
rect 82638 21090 82648 21118
rect 81868 21031 82356 21037
rect 81868 20997 81880 21031
rect 82344 20997 82356 21031
rect 81868 20991 82356 20997
rect 82092 20934 82152 20991
rect 82588 20934 82648 21090
rect 83616 21090 83622 21638
rect 83656 21638 83672 21666
rect 84634 21666 84680 21678
rect 83656 21090 83662 21638
rect 84634 21126 84640 21666
rect 83616 21078 83662 21090
rect 84624 21090 84640 21126
rect 84674 21126 84680 21666
rect 85646 21666 85706 21820
rect 86142 21765 86202 22247
rect 86662 22188 86722 22346
rect 87688 22346 87694 22898
rect 87728 22898 87740 22922
rect 87728 22346 87734 22898
rect 87688 22334 87734 22346
rect 86958 22287 87446 22293
rect 86958 22253 86970 22287
rect 87434 22253 87446 22287
rect 86958 22247 87446 22253
rect 86656 22128 86662 22188
rect 86722 22128 86728 22188
rect 87922 21934 87928 21994
rect 87988 21934 87994 21994
rect 86664 21826 87740 21886
rect 85940 21759 86428 21765
rect 85940 21725 85952 21759
rect 86416 21725 86428 21759
rect 85940 21719 86428 21725
rect 85646 21642 85658 21666
rect 84674 21090 84684 21126
rect 85652 21118 85658 21642
rect 84106 21037 84166 21038
rect 82886 21031 83374 21037
rect 82886 20997 82898 21031
rect 83362 20997 83374 21031
rect 82886 20991 83374 20997
rect 83904 21031 84392 21037
rect 83904 20997 83916 21031
rect 84380 20997 84392 21031
rect 83904 20991 84392 20997
rect 83104 20934 83164 20991
rect 81568 20872 81574 20932
rect 81634 20872 81640 20932
rect 82092 20874 83164 20934
rect 81566 20566 81572 20626
rect 81632 20566 81638 20626
rect 79832 20503 80320 20509
rect 79832 20469 79844 20503
rect 80308 20469 80320 20503
rect 79832 20463 80320 20469
rect 80850 20503 81338 20509
rect 80850 20469 80862 20503
rect 81326 20469 81338 20503
rect 80850 20463 81338 20469
rect 79538 20388 79550 20410
rect 78566 19864 78572 20386
rect 78566 19834 78580 19864
rect 77796 19775 78284 19781
rect 77796 19741 77808 19775
rect 78272 19741 78284 19775
rect 77796 19735 78284 19741
rect 78014 19684 78074 19735
rect 77002 19624 78074 19684
rect 78520 19678 78580 19834
rect 79544 19834 79550 20388
rect 79584 20388 79598 20410
rect 80562 20410 80608 20422
rect 79584 19834 79590 20388
rect 80562 19860 80568 20410
rect 79544 19822 79590 19834
rect 80556 19834 80568 19860
rect 80602 19860 80608 20410
rect 81572 20410 81632 20566
rect 81868 20503 82356 20509
rect 81868 20469 81880 20503
rect 82344 20469 82356 20503
rect 81868 20463 82356 20469
rect 81572 20384 81586 20410
rect 80602 19834 80616 19860
rect 80046 19781 80106 19784
rect 78814 19775 79302 19781
rect 78814 19741 78826 19775
rect 79290 19741 79302 19775
rect 78814 19735 79302 19741
rect 79832 19775 80320 19781
rect 79832 19741 79844 19775
rect 80308 19741 80320 19775
rect 79832 19735 80320 19741
rect 75966 19458 76742 19518
rect 75966 19253 76026 19458
rect 76682 19372 76742 19458
rect 76472 19306 76478 19366
rect 76538 19306 76544 19366
rect 76676 19312 76682 19372
rect 76742 19312 76748 19372
rect 74742 19247 75230 19253
rect 74742 19213 74754 19247
rect 75218 19213 75230 19247
rect 74742 19207 75230 19213
rect 75760 19247 76248 19253
rect 75760 19213 75772 19247
rect 76236 19213 76248 19247
rect 75760 19207 76248 19213
rect 74444 19128 74460 19154
rect 73476 18604 73482 19128
rect 73476 18578 73486 18604
rect 72706 18519 73194 18525
rect 72706 18485 72718 18519
rect 73182 18485 73194 18519
rect 72706 18479 73194 18485
rect 73426 18418 73486 18578
rect 74454 18578 74460 19128
rect 74494 19128 74504 19154
rect 75472 19154 75518 19166
rect 74494 18578 74500 19128
rect 75472 18600 75478 19154
rect 74454 18566 74500 18578
rect 75462 18578 75478 18600
rect 75512 18600 75518 19154
rect 76478 19154 76538 19306
rect 76778 19247 77266 19253
rect 76778 19213 76790 19247
rect 77254 19213 77266 19247
rect 76778 19207 77266 19213
rect 76478 19124 76496 19154
rect 76490 18614 76496 19124
rect 75512 18578 75522 18600
rect 73724 18519 74212 18525
rect 73724 18485 73736 18519
rect 74200 18485 74212 18519
rect 73724 18479 74212 18485
rect 74742 18519 75230 18525
rect 74742 18485 74754 18519
rect 75218 18485 75230 18519
rect 74742 18479 75230 18485
rect 73420 18358 73426 18418
rect 73486 18358 73492 18418
rect 73934 18304 73994 18479
rect 74958 18304 75018 18479
rect 75462 18418 75522 18578
rect 76484 18578 76496 18614
rect 76530 19124 76538 19154
rect 77498 19154 77558 19624
rect 78514 19618 78520 19678
rect 78580 19618 78586 19678
rect 79030 19546 79090 19735
rect 80046 19546 80106 19735
rect 80556 19678 80616 19834
rect 81580 19834 81586 20384
rect 81620 20384 81632 20410
rect 82588 20410 82648 20874
rect 83602 20768 83608 20828
rect 83668 20768 83674 20828
rect 82886 20503 83374 20509
rect 82886 20469 82898 20503
rect 83362 20469 83374 20503
rect 82886 20463 83374 20469
rect 81620 19834 81626 20384
rect 82588 20380 82604 20410
rect 82598 19866 82604 20380
rect 81580 19822 81626 19834
rect 82586 19834 82604 19866
rect 82638 20380 82648 20410
rect 83608 20410 83668 20768
rect 84106 20509 84166 20991
rect 84470 20886 84476 20946
rect 84536 20886 84542 20946
rect 84476 20626 84536 20886
rect 84624 20836 84684 21090
rect 85644 21090 85658 21118
rect 85692 21642 85706 21666
rect 86664 21666 86724 21826
rect 87178 21765 87238 21826
rect 86958 21759 87446 21765
rect 86958 21725 86970 21759
rect 87434 21725 87446 21759
rect 86958 21719 87446 21725
rect 85692 21118 85698 21642
rect 86664 21632 86676 21666
rect 86670 21130 86676 21632
rect 85692 21090 85704 21118
rect 85130 21037 85190 21038
rect 84922 21031 85410 21037
rect 84922 20997 84934 21031
rect 85398 20997 85410 21031
rect 84922 20991 85410 20997
rect 84618 20776 84624 20836
rect 84684 20776 84690 20836
rect 84470 20566 84476 20626
rect 84536 20566 84542 20626
rect 84622 20568 84628 20628
rect 84688 20568 84694 20628
rect 83904 20503 84392 20509
rect 83904 20469 83916 20503
rect 84380 20469 84392 20503
rect 83904 20463 84392 20469
rect 82638 19866 82644 20380
rect 83608 20378 83622 20410
rect 83616 19866 83622 20378
rect 82638 19834 82646 19866
rect 80850 19775 81338 19781
rect 80850 19741 80862 19775
rect 81326 19741 81338 19775
rect 80850 19735 81338 19741
rect 81868 19775 82356 19781
rect 81868 19741 81880 19775
rect 82344 19741 82356 19775
rect 81868 19735 82356 19741
rect 80550 19618 80556 19678
rect 80616 19618 80622 19678
rect 81060 19546 81120 19735
rect 82090 19682 82150 19735
rect 82586 19682 82646 19834
rect 83610 19834 83622 19866
rect 83656 20378 83668 20410
rect 84628 20410 84688 20568
rect 85130 20509 85190 20991
rect 85644 20726 85704 21090
rect 86664 21090 86676 21130
rect 86710 21632 86724 21666
rect 87680 21666 87740 21826
rect 87680 21644 87694 21666
rect 86710 21130 86716 21632
rect 86710 21090 86724 21130
rect 86136 21037 86196 21044
rect 85940 21031 86428 21037
rect 85940 20997 85952 21031
rect 86416 20997 86428 21031
rect 85940 20991 86428 20997
rect 85638 20666 85644 20726
rect 85704 20666 85710 20726
rect 86136 20509 86196 20991
rect 86664 20836 86724 21090
rect 87688 21090 87694 21644
rect 87728 21644 87740 21666
rect 87728 21090 87734 21644
rect 87688 21078 87734 21090
rect 86958 21031 87446 21037
rect 86958 20997 86970 21031
rect 87434 20997 87446 21031
rect 86958 20991 87446 20997
rect 86658 20776 86664 20836
rect 86724 20776 86730 20836
rect 87790 20776 87796 20836
rect 87856 20776 87862 20836
rect 86656 20568 86662 20628
rect 86722 20568 86728 20628
rect 84922 20503 85410 20509
rect 84922 20469 84934 20503
rect 85398 20469 85410 20503
rect 84922 20463 85410 20469
rect 85940 20503 86428 20509
rect 85940 20469 85952 20503
rect 86416 20469 86428 20503
rect 85940 20463 86428 20469
rect 84628 20390 84640 20410
rect 83656 19866 83662 20378
rect 83656 19834 83670 19866
rect 82886 19775 83374 19781
rect 82886 19741 82898 19775
rect 83362 19741 83374 19775
rect 82886 19735 83374 19741
rect 83102 19682 83162 19735
rect 82090 19622 83162 19682
rect 83610 19680 83670 19834
rect 84634 19834 84640 20390
rect 84674 20390 84688 20410
rect 85652 20410 85698 20422
rect 84674 19834 84680 20390
rect 85652 19862 85658 20410
rect 84634 19822 84680 19834
rect 85646 19834 85658 19862
rect 85692 19862 85698 20410
rect 86662 20410 86722 20568
rect 86958 20503 87446 20509
rect 86958 20469 86970 20503
rect 87434 20469 87446 20503
rect 86958 20463 87446 20469
rect 86662 20386 86676 20410
rect 86670 19870 86676 20386
rect 85692 19834 85706 19862
rect 84118 19781 84178 19788
rect 85142 19781 85202 19788
rect 83904 19775 84392 19781
rect 83904 19741 83916 19775
rect 84380 19741 84392 19775
rect 83904 19735 84392 19741
rect 84922 19775 85410 19781
rect 84922 19741 84934 19775
rect 85398 19741 85410 19775
rect 84922 19735 85410 19741
rect 79030 19486 81844 19546
rect 78516 19372 78576 19378
rect 79030 19372 79090 19486
rect 78576 19312 79090 19372
rect 78516 19306 78576 19312
rect 79530 19308 79536 19368
rect 79596 19308 79602 19368
rect 81564 19308 81570 19368
rect 81630 19308 81636 19368
rect 81784 19364 81844 19486
rect 77796 19247 78284 19253
rect 77796 19213 77808 19247
rect 78272 19213 78284 19247
rect 77796 19207 78284 19213
rect 78814 19247 79302 19253
rect 78814 19213 78826 19247
rect 79290 19213 79302 19247
rect 78814 19207 79302 19213
rect 76530 18614 76536 19124
rect 77498 19096 77514 19154
rect 76530 18578 76544 18614
rect 77508 18610 77514 19096
rect 75760 18519 76248 18525
rect 75760 18485 75772 18519
rect 76236 18485 76248 18519
rect 75760 18479 76248 18485
rect 75456 18358 75462 18418
rect 75522 18358 75528 18418
rect 75964 18304 76024 18479
rect 72124 18228 72130 18288
rect 72190 18228 72196 18288
rect 73934 18244 76024 18304
rect 67054 18088 67060 18148
rect 67120 18088 67126 18148
rect 66904 18042 66964 18048
rect 72130 18042 72190 18228
rect 66964 17982 72190 18042
rect 66904 17976 66964 17982
rect 66134 17924 66194 17930
rect 73934 17924 73994 18244
rect 75964 17994 76024 18244
rect 76484 18148 76544 18578
rect 77498 18578 77514 18610
rect 77548 19096 77558 19154
rect 78526 19154 78572 19166
rect 77548 18610 77554 19096
rect 78526 18622 78532 19154
rect 77548 18578 77558 18610
rect 76778 18519 77266 18525
rect 76778 18485 76790 18519
rect 77254 18485 77266 18519
rect 76778 18479 77266 18485
rect 77002 18424 77062 18479
rect 77498 18424 77558 18578
rect 78520 18578 78532 18622
rect 78566 18622 78572 19154
rect 79536 19154 79596 19308
rect 79832 19247 80320 19253
rect 79832 19213 79844 19247
rect 80308 19213 80320 19247
rect 79832 19207 80320 19213
rect 80850 19247 81338 19253
rect 80850 19213 80862 19247
rect 81326 19213 81338 19247
rect 80850 19207 81338 19213
rect 79536 19130 79550 19154
rect 78566 18578 78580 18622
rect 79544 18602 79550 19130
rect 77796 18519 78284 18525
rect 77796 18485 77808 18519
rect 78272 18485 78284 18519
rect 77796 18479 78284 18485
rect 78014 18424 78074 18479
rect 78520 18424 78580 18578
rect 79536 18578 79550 18602
rect 79584 19130 79596 19154
rect 80562 19154 80608 19166
rect 79584 18602 79590 19130
rect 80562 18616 80568 19154
rect 79584 18578 79596 18602
rect 78814 18519 79302 18525
rect 78814 18485 78826 18519
rect 79290 18485 79302 18519
rect 78814 18479 79302 18485
rect 79030 18424 79090 18479
rect 79536 18424 79596 18578
rect 80554 18578 80568 18616
rect 80602 18616 80608 19154
rect 81570 19154 81630 19308
rect 81778 19304 81784 19364
rect 81844 19304 81850 19364
rect 81868 19247 82356 19253
rect 81868 19213 81880 19247
rect 82344 19213 82356 19247
rect 81868 19207 82356 19213
rect 81570 19126 81586 19154
rect 80602 18578 80614 18616
rect 81580 18606 81586 19126
rect 79832 18519 80320 18525
rect 79832 18485 79844 18519
rect 80308 18485 80320 18519
rect 79832 18479 80320 18485
rect 80046 18424 80106 18479
rect 80554 18424 80614 18578
rect 81572 18578 81586 18606
rect 81620 19126 81630 19154
rect 82586 19154 82646 19622
rect 83604 19620 83610 19680
rect 83670 19620 83676 19680
rect 84118 19370 84178 19735
rect 84118 19364 84180 19370
rect 84118 19304 84120 19364
rect 84626 19306 84632 19366
rect 84692 19306 84698 19366
rect 84118 19298 84180 19304
rect 84118 19253 84178 19298
rect 82886 19247 83374 19253
rect 82886 19213 82898 19247
rect 83362 19213 83374 19247
rect 82886 19207 83374 19213
rect 83904 19247 84392 19253
rect 83904 19213 83916 19247
rect 84380 19213 84392 19247
rect 83904 19207 84392 19213
rect 81620 18606 81626 19126
rect 82586 19116 82604 19154
rect 82598 18608 82604 19116
rect 81620 18578 81632 18606
rect 80850 18519 81338 18525
rect 80850 18485 80862 18519
rect 81326 18485 81338 18519
rect 80850 18479 81338 18485
rect 81056 18424 81116 18479
rect 81572 18424 81632 18578
rect 82586 18578 82604 18608
rect 82638 19116 82646 19154
rect 83616 19154 83662 19166
rect 82638 18608 82644 19116
rect 82638 18578 82646 18608
rect 83616 18604 83622 19154
rect 81868 18519 82356 18525
rect 81868 18485 81880 18519
rect 82344 18485 82356 18519
rect 81868 18479 82356 18485
rect 82090 18424 82150 18479
rect 82586 18424 82646 18578
rect 83614 18578 83622 18604
rect 83656 18604 83662 19154
rect 84632 19154 84692 19306
rect 85142 19253 85202 19735
rect 85646 19680 85706 19834
rect 86662 19834 86676 19870
rect 86710 20386 86722 20410
rect 87688 20410 87734 20422
rect 86710 19870 86716 20386
rect 86710 19834 86722 19870
rect 87688 19858 87694 20410
rect 86148 19781 86208 19794
rect 85940 19775 86428 19781
rect 85940 19741 85952 19775
rect 86416 19741 86428 19775
rect 85940 19735 86428 19741
rect 85640 19620 85646 19680
rect 85706 19620 85712 19680
rect 86148 19253 86208 19735
rect 86662 19676 86722 19834
rect 87678 19834 87694 19858
rect 87728 19858 87734 20410
rect 87728 19834 87738 19858
rect 86958 19775 87446 19781
rect 86958 19741 86970 19775
rect 87434 19741 87446 19775
rect 86958 19735 87446 19741
rect 87176 19676 87236 19735
rect 87678 19676 87738 19834
rect 86662 19616 87738 19676
rect 87796 19568 87856 20776
rect 87928 20628 87988 21934
rect 87922 20568 87928 20628
rect 87988 20568 87994 20628
rect 87790 19508 87796 19568
rect 87856 19508 87862 19568
rect 86660 19306 86666 19366
rect 86726 19306 86732 19366
rect 84922 19247 85410 19253
rect 84922 19213 84934 19247
rect 85398 19213 85410 19247
rect 84922 19207 85410 19213
rect 85940 19247 86428 19253
rect 85940 19213 85952 19247
rect 86416 19213 86428 19247
rect 85940 19207 86428 19213
rect 84632 19128 84640 19154
rect 83656 18578 83674 18604
rect 82886 18519 83374 18525
rect 82886 18485 82898 18519
rect 83362 18485 83374 18519
rect 82886 18479 83374 18485
rect 83102 18424 83162 18479
rect 77002 18364 83162 18424
rect 83614 18418 83674 18578
rect 84634 18578 84640 19128
rect 84674 19128 84692 19154
rect 85652 19154 85698 19166
rect 84674 18578 84680 19128
rect 85652 18600 85658 19154
rect 84634 18566 84680 18578
rect 85650 18578 85658 18600
rect 85692 18600 85698 19154
rect 86666 19154 86726 19306
rect 86958 19247 87446 19253
rect 86958 19213 86970 19247
rect 87434 19213 87446 19247
rect 86958 19207 87446 19213
rect 86666 19124 86676 19154
rect 86670 18616 86676 19124
rect 85692 18578 85710 18600
rect 84122 18525 84182 18532
rect 83904 18519 84392 18525
rect 83904 18485 83916 18519
rect 84380 18485 84392 18519
rect 83904 18479 84392 18485
rect 84922 18519 85410 18525
rect 84922 18485 84934 18519
rect 85398 18485 85410 18519
rect 84922 18479 85410 18485
rect 83608 18358 83614 18418
rect 83674 18358 83680 18418
rect 84122 18306 84182 18479
rect 85142 18306 85202 18479
rect 85650 18418 85710 18578
rect 86664 18578 86676 18616
rect 86710 19124 86726 19154
rect 87688 19154 87734 19166
rect 86710 18616 86716 19124
rect 86710 18578 86724 18616
rect 87688 18604 87694 19154
rect 85940 18519 86428 18525
rect 85940 18485 85952 18519
rect 86416 18485 86428 18519
rect 85940 18479 86428 18485
rect 85644 18358 85650 18418
rect 85710 18358 85716 18418
rect 86144 18306 86204 18479
rect 86664 18422 86724 18578
rect 87680 18578 87694 18604
rect 87728 18604 87734 19154
rect 87728 18578 87740 18604
rect 86958 18519 87446 18525
rect 86958 18485 86970 18519
rect 87434 18485 87446 18519
rect 86958 18479 87446 18485
rect 87178 18422 87238 18479
rect 87680 18422 87740 18578
rect 86664 18362 87740 18422
rect 84122 18246 86204 18306
rect 76478 18088 76484 18148
rect 76544 18088 76550 18148
rect 84122 17994 84182 18246
rect 88088 18148 88148 23076
rect 89666 18278 89672 27642
rect 89772 18278 89778 27642
rect 88082 18088 88088 18148
rect 88148 18088 88154 18148
rect 75964 17934 84182 17994
rect 66194 17864 73994 17924
rect 66134 17858 66194 17864
rect 89666 17764 89778 18278
rect 65322 17758 89778 17764
rect 65322 17658 65428 17758
rect 89672 17658 89778 17758
rect 65322 17652 89778 17658
rect 64305 15368 64427 15373
rect 52622 15364 89878 15368
rect 52622 15362 59912 15364
rect 60012 15362 62512 15364
rect 62612 15362 64316 15364
rect 64416 15362 89878 15364
rect 52622 15262 52728 15362
rect 89772 15262 89878 15362
rect 52622 15256 89878 15262
rect 52622 14470 52734 15256
rect 66898 15132 66904 15192
rect 66964 15132 66970 15192
rect 67054 15132 67060 15192
rect 67120 15132 67126 15192
rect 67286 15184 67346 15190
rect 50938 9048 50944 9108
rect 51004 9048 51010 9108
rect 48494 8514 50513 8574
rect 48358 7491 48364 7551
rect 48424 7491 48430 7551
rect 48364 6176 48424 7491
rect 48494 6610 48554 8514
rect 48677 8448 48982 8514
rect 48677 8414 48736 8448
rect 48956 8414 48982 8448
rect 48677 8400 48982 8414
rect 48677 8350 48738 8400
rect 48677 8320 48688 8350
rect 48678 8092 48688 8320
rect 48677 8032 48688 8092
rect 48678 7778 48688 8032
rect 48726 8092 48738 8350
rect 48788 8252 48848 8400
rect 48922 8351 48982 8400
rect 49178 8466 49238 8467
rect 49954 8466 50014 8472
rect 49178 8406 49954 8466
rect 49178 8351 49238 8406
rect 49436 8351 49496 8406
rect 49694 8351 49754 8406
rect 49954 8351 50014 8406
rect 50210 8448 50513 8514
rect 50210 8414 50228 8448
rect 50430 8414 50513 8448
rect 50210 8400 50513 8414
rect 50210 8351 50270 8400
rect 48896 8345 49004 8351
rect 48896 8311 48908 8345
rect 48992 8311 49004 8345
rect 48896 8305 49004 8311
rect 49154 8345 49262 8351
rect 49154 8311 49166 8345
rect 49250 8311 49262 8345
rect 49154 8305 49262 8311
rect 49412 8345 49520 8351
rect 49412 8311 49424 8345
rect 49508 8311 49520 8345
rect 49412 8305 49520 8311
rect 49670 8345 49778 8351
rect 49670 8311 49682 8345
rect 49766 8311 49778 8345
rect 49670 8305 49778 8311
rect 49928 8345 50036 8351
rect 49928 8311 49940 8345
rect 50024 8311 50036 8345
rect 49928 8305 50036 8311
rect 50186 8345 50294 8351
rect 50186 8311 50198 8345
rect 50282 8311 50294 8345
rect 50186 8305 50294 8311
rect 48788 8092 48804 8252
rect 48726 8032 48804 8092
rect 48726 7778 48738 8032
rect 48798 7910 48804 8032
rect 48678 7728 48738 7778
rect 48790 7876 48804 7910
rect 48838 8032 48848 8252
rect 49056 8252 49102 8264
rect 48838 7910 48844 8032
rect 49056 7921 49062 8252
rect 48838 7876 48850 7910
rect 48790 7728 48850 7876
rect 49048 7876 49062 7921
rect 49096 7921 49102 8252
rect 49314 8252 49360 8264
rect 49096 7876 49108 7921
rect 49314 7896 49320 8252
rect 48896 7817 49004 7823
rect 48896 7783 48908 7817
rect 48992 7783 49004 7817
rect 48896 7777 49004 7783
rect 48918 7728 48978 7777
rect 48677 7714 48978 7728
rect 48677 7680 48736 7714
rect 48956 7680 48978 7714
rect 48677 7668 48978 7680
rect 49048 7551 49108 7876
rect 49306 7876 49320 7896
rect 49354 7896 49360 8252
rect 49572 8252 49618 8264
rect 49572 7919 49578 8252
rect 49354 7876 49366 7896
rect 49154 7817 49262 7823
rect 49154 7783 49166 7817
rect 49250 7783 49262 7817
rect 49154 7777 49262 7783
rect 49306 7700 49366 7876
rect 49564 7876 49578 7919
rect 49612 7919 49618 8252
rect 49830 8252 49876 8264
rect 49612 7876 49624 7919
rect 49830 7914 49836 8252
rect 49412 7817 49520 7823
rect 49412 7783 49424 7817
rect 49508 7783 49520 7817
rect 49412 7777 49520 7783
rect 49300 7640 49306 7700
rect 49366 7640 49372 7700
rect 48676 7516 48980 7526
rect 48676 7478 48760 7516
rect 48968 7478 48980 7516
rect 49042 7491 49048 7551
rect 49108 7491 49114 7551
rect 48676 7466 48980 7478
rect 48676 7418 48736 7466
rect 48676 7062 48688 7418
rect 48724 7062 48736 7418
rect 48790 7328 48850 7466
rect 48920 7418 48980 7466
rect 48896 7412 49004 7418
rect 48896 7378 48908 7412
rect 48992 7378 49004 7412
rect 48896 7372 49004 7378
rect 48790 7278 48804 7328
rect 48798 7191 48804 7278
rect 48676 7013 48736 7062
rect 48792 7152 48804 7191
rect 48838 7278 48850 7328
rect 49048 7328 49108 7491
rect 49154 7412 49262 7418
rect 49154 7378 49166 7412
rect 49250 7378 49262 7412
rect 49154 7372 49262 7378
rect 49048 7291 49062 7328
rect 48838 7191 48844 7278
rect 48838 7152 48852 7191
rect 48792 7013 48852 7152
rect 49056 7152 49062 7291
rect 49096 7291 49108 7328
rect 49306 7358 49366 7640
rect 49564 7551 49624 7876
rect 49824 7876 49836 7914
rect 49870 7914 49876 8252
rect 50088 8252 50134 8264
rect 50088 7919 50094 8252
rect 49870 7876 49884 7914
rect 49670 7817 49778 7823
rect 49670 7783 49682 7817
rect 49766 7783 49778 7817
rect 49670 7777 49778 7783
rect 49824 7700 49884 7876
rect 50082 7876 50094 7919
rect 50128 7919 50134 8252
rect 50338 8252 50398 8400
rect 50338 8034 50352 8252
rect 50128 7876 50142 7919
rect 50346 7906 50352 8034
rect 49928 7817 50036 7823
rect 49928 7783 49940 7817
rect 50024 7783 50036 7817
rect 49928 7777 50036 7783
rect 49818 7640 49824 7700
rect 49884 7640 49890 7700
rect 49558 7491 49564 7551
rect 49624 7491 49630 7551
rect 49412 7412 49520 7418
rect 49412 7378 49424 7412
rect 49508 7378 49520 7412
rect 49412 7372 49520 7378
rect 49306 7328 49368 7358
rect 49306 7292 49320 7328
rect 49096 7152 49102 7291
rect 49056 7140 49102 7152
rect 49308 7152 49320 7292
rect 49354 7152 49368 7328
rect 49564 7328 49624 7491
rect 49670 7412 49778 7418
rect 49670 7378 49682 7412
rect 49766 7378 49778 7412
rect 49670 7372 49778 7378
rect 49564 7172 49578 7328
rect 49308 7112 49368 7152
rect 49572 7152 49578 7172
rect 49612 7172 49624 7328
rect 49824 7328 49884 7640
rect 50082 7551 50142 7876
rect 50340 7876 50352 7906
rect 50386 8094 50398 8252
rect 50452 8352 50513 8400
rect 50452 8094 50464 8352
rect 50386 8034 50464 8094
rect 50386 7906 50392 8034
rect 50386 7876 50400 7906
rect 50186 7817 50294 7823
rect 50186 7783 50198 7817
rect 50282 7783 50294 7817
rect 50186 7777 50294 7783
rect 50206 7728 50266 7777
rect 50340 7728 50400 7876
rect 50452 7776 50464 8034
rect 50500 8336 50513 8352
rect 50500 7976 50512 8336
rect 50500 7945 50850 7976
rect 50500 7911 50603 7945
rect 50637 7911 50695 7945
rect 50729 7911 50787 7945
rect 50821 7911 50850 7945
rect 50500 7880 50850 7911
rect 50500 7776 50512 7880
rect 50452 7728 50512 7776
rect 50206 7716 50512 7728
rect 50206 7682 50228 7716
rect 50430 7682 50512 7716
rect 50206 7668 50512 7682
rect 50944 7656 51004 9048
rect 50944 7650 51005 7656
rect 50725 7644 50945 7650
rect 50627 7628 50687 7634
rect 50621 7568 50627 7628
rect 50687 7568 50693 7628
rect 50725 7604 50737 7644
rect 50783 7604 50945 7644
rect 50725 7590 50945 7604
rect 50945 7584 51005 7590
rect 50627 7562 50687 7568
rect 49928 7412 50036 7418
rect 49928 7378 49940 7412
rect 50024 7378 50036 7412
rect 49928 7372 50036 7378
rect 49612 7152 49618 7172
rect 49572 7140 49618 7152
rect 49824 7152 49836 7328
rect 49870 7152 49884 7328
rect 50082 7328 50142 7491
rect 50212 7518 50514 7528
rect 50212 7480 50232 7518
rect 50430 7480 50514 7518
rect 50212 7468 50514 7480
rect 50212 7418 50272 7468
rect 50186 7412 50294 7418
rect 50186 7378 50198 7412
rect 50282 7378 50294 7412
rect 50186 7372 50294 7378
rect 50082 7289 50094 7328
rect 49824 7112 49884 7152
rect 50088 7152 50094 7289
rect 50128 7289 50142 7328
rect 50340 7328 50400 7468
rect 50128 7152 50134 7289
rect 50340 7282 50352 7328
rect 50346 7185 50352 7282
rect 50088 7140 50134 7152
rect 50338 7152 50352 7185
rect 50386 7282 50400 7328
rect 50454 7432 50514 7468
rect 50454 7418 50850 7432
rect 50386 7185 50392 7282
rect 50386 7152 50398 7185
rect 48896 7102 49004 7108
rect 48896 7068 48908 7102
rect 48992 7068 49004 7102
rect 48896 7062 49004 7068
rect 49154 7102 49262 7108
rect 49154 7068 49166 7102
rect 49250 7068 49262 7102
rect 49154 7062 49262 7068
rect 49412 7102 49520 7108
rect 49412 7068 49424 7102
rect 49508 7068 49520 7102
rect 49412 7062 49520 7068
rect 49670 7102 49778 7108
rect 49670 7068 49682 7102
rect 49766 7068 49778 7102
rect 49670 7062 49778 7068
rect 49928 7102 50036 7108
rect 49928 7068 49940 7102
rect 50024 7068 50036 7102
rect 49928 7062 50036 7068
rect 50186 7102 50294 7108
rect 50186 7068 50198 7102
rect 50282 7068 50294 7102
rect 50186 7062 50294 7068
rect 48920 7013 48980 7062
rect 48676 7002 48980 7013
rect 48676 6966 48758 7002
rect 48966 6966 48980 7002
rect 48676 6896 48980 6966
rect 49178 7003 49238 7062
rect 49438 7003 49498 7062
rect 49696 7003 49756 7062
rect 49952 7003 50012 7062
rect 50210 7013 50270 7062
rect 50338 7013 50398 7152
rect 50454 7062 50464 7418
rect 50502 7401 50850 7418
rect 50502 7367 50603 7401
rect 50637 7367 50695 7401
rect 50729 7367 50787 7401
rect 50821 7367 50850 7401
rect 50502 7336 50850 7367
rect 50502 7062 50514 7336
rect 50454 7013 50514 7062
rect 49178 6943 49952 7003
rect 50012 6943 50018 7003
rect 50210 7000 50514 7013
rect 50210 6964 50230 7000
rect 50432 6964 50514 7000
rect 48677 6878 48980 6896
rect 50210 6878 50514 6964
rect 52622 6878 52628 14470
rect 48677 6818 52628 6878
rect 48494 6550 50513 6610
rect 48358 6116 48364 6176
rect 48424 6116 48430 6176
rect 48494 4610 48554 6550
rect 48677 6484 48982 6550
rect 48677 6450 48736 6484
rect 48956 6450 48982 6484
rect 48677 6436 48982 6450
rect 48677 6386 48738 6436
rect 48677 6356 48688 6386
rect 48678 6128 48688 6356
rect 48677 6068 48688 6128
rect 48678 5814 48688 6068
rect 48726 6128 48738 6386
rect 48788 6288 48848 6436
rect 48922 6387 48982 6436
rect 49178 6502 49238 6503
rect 49954 6502 50014 6508
rect 49178 6442 49954 6502
rect 49178 6387 49238 6442
rect 49436 6387 49496 6442
rect 49694 6387 49754 6442
rect 49954 6387 50014 6442
rect 50210 6484 50513 6550
rect 50210 6450 50228 6484
rect 50430 6450 50513 6484
rect 50210 6436 50513 6450
rect 50210 6387 50270 6436
rect 48896 6381 49004 6387
rect 48896 6347 48908 6381
rect 48992 6347 49004 6381
rect 48896 6341 49004 6347
rect 49154 6381 49262 6387
rect 49154 6347 49166 6381
rect 49250 6347 49262 6381
rect 49154 6341 49262 6347
rect 49412 6381 49520 6387
rect 49412 6347 49424 6381
rect 49508 6347 49520 6381
rect 49412 6341 49520 6347
rect 49670 6381 49778 6387
rect 49670 6347 49682 6381
rect 49766 6347 49778 6381
rect 49670 6341 49778 6347
rect 49928 6381 50036 6387
rect 49928 6347 49940 6381
rect 50024 6347 50036 6381
rect 49928 6341 50036 6347
rect 50186 6381 50294 6387
rect 50186 6347 50198 6381
rect 50282 6347 50294 6381
rect 50186 6341 50294 6347
rect 48788 6128 48804 6288
rect 48726 6068 48804 6128
rect 48726 5814 48738 6068
rect 48798 5946 48804 6068
rect 48678 5764 48738 5814
rect 48790 5912 48804 5946
rect 48838 6068 48848 6288
rect 49056 6288 49102 6300
rect 48838 5946 48844 6068
rect 49056 5957 49062 6288
rect 48838 5912 48850 5946
rect 48790 5764 48850 5912
rect 49048 5912 49062 5957
rect 49096 5957 49102 6288
rect 49314 6288 49360 6300
rect 49096 5912 49108 5957
rect 49314 5932 49320 6288
rect 48896 5853 49004 5859
rect 48896 5819 48908 5853
rect 48992 5819 49004 5853
rect 48896 5813 49004 5819
rect 48918 5764 48978 5813
rect 48677 5750 48978 5764
rect 48677 5716 48736 5750
rect 48956 5716 48978 5750
rect 48677 5704 48978 5716
rect 49048 5587 49108 5912
rect 49306 5912 49320 5932
rect 49354 5932 49360 6288
rect 49572 6288 49618 6300
rect 49572 5955 49578 6288
rect 49354 5912 49366 5932
rect 49154 5853 49262 5859
rect 49154 5819 49166 5853
rect 49250 5819 49262 5853
rect 49154 5813 49262 5819
rect 49306 5736 49366 5912
rect 49564 5912 49578 5955
rect 49612 5955 49618 6288
rect 49830 6288 49876 6300
rect 49612 5912 49624 5955
rect 49830 5950 49836 6288
rect 49412 5853 49520 5859
rect 49412 5819 49424 5853
rect 49508 5819 49520 5853
rect 49412 5813 49520 5819
rect 49300 5676 49306 5736
rect 49366 5676 49372 5736
rect 48676 5552 48980 5562
rect 48676 5514 48760 5552
rect 48968 5514 48980 5552
rect 49042 5527 49048 5587
rect 49108 5527 49114 5587
rect 48676 5502 48980 5514
rect 48676 5454 48736 5502
rect 48676 5098 48688 5454
rect 48724 5098 48736 5454
rect 48790 5364 48850 5502
rect 48920 5454 48980 5502
rect 48896 5448 49004 5454
rect 48896 5414 48908 5448
rect 48992 5414 49004 5448
rect 48896 5408 49004 5414
rect 48790 5314 48804 5364
rect 48798 5227 48804 5314
rect 48676 5049 48736 5098
rect 48792 5188 48804 5227
rect 48838 5314 48850 5364
rect 49048 5364 49108 5527
rect 49154 5448 49262 5454
rect 49154 5414 49166 5448
rect 49250 5414 49262 5448
rect 49154 5408 49262 5414
rect 49048 5327 49062 5364
rect 48838 5227 48844 5314
rect 48838 5188 48852 5227
rect 48792 5049 48852 5188
rect 49056 5188 49062 5327
rect 49096 5327 49108 5364
rect 49306 5394 49366 5676
rect 49564 5587 49624 5912
rect 49824 5912 49836 5950
rect 49870 5950 49876 6288
rect 50088 6288 50134 6300
rect 50088 5955 50094 6288
rect 49870 5912 49884 5950
rect 49670 5853 49778 5859
rect 49670 5819 49682 5853
rect 49766 5819 49778 5853
rect 49670 5813 49778 5819
rect 49824 5736 49884 5912
rect 50082 5912 50094 5955
rect 50128 5955 50134 6288
rect 50338 6288 50398 6436
rect 50338 6070 50352 6288
rect 50128 5912 50142 5955
rect 50346 5942 50352 6070
rect 49928 5853 50036 5859
rect 49928 5819 49940 5853
rect 50024 5819 50036 5853
rect 49928 5813 50036 5819
rect 49818 5676 49824 5736
rect 49884 5676 49890 5736
rect 49558 5527 49564 5587
rect 49624 5527 49630 5587
rect 49412 5448 49520 5454
rect 49412 5414 49424 5448
rect 49508 5414 49520 5448
rect 49412 5408 49520 5414
rect 49306 5364 49368 5394
rect 49306 5328 49320 5364
rect 49096 5188 49102 5327
rect 49056 5176 49102 5188
rect 49308 5188 49320 5328
rect 49354 5188 49368 5364
rect 49564 5364 49624 5527
rect 49670 5448 49778 5454
rect 49670 5414 49682 5448
rect 49766 5414 49778 5448
rect 49670 5408 49778 5414
rect 49564 5208 49578 5364
rect 49308 5148 49368 5188
rect 49572 5188 49578 5208
rect 49612 5208 49624 5364
rect 49824 5364 49884 5676
rect 50082 5587 50142 5912
rect 50340 5912 50352 5942
rect 50386 6130 50398 6288
rect 50452 6388 50513 6436
rect 50452 6130 50464 6388
rect 50386 6070 50464 6130
rect 50386 5942 50392 6070
rect 50386 5912 50400 5942
rect 50186 5853 50294 5859
rect 50186 5819 50198 5853
rect 50282 5819 50294 5853
rect 50186 5813 50294 5819
rect 50206 5764 50266 5813
rect 50340 5764 50400 5912
rect 50452 5812 50464 6070
rect 50500 6372 50513 6388
rect 50500 6012 50512 6372
rect 50500 5981 50850 6012
rect 50500 5947 50603 5981
rect 50637 5947 50695 5981
rect 50729 5947 50787 5981
rect 50821 5947 50850 5981
rect 50500 5916 50850 5947
rect 50500 5812 50512 5916
rect 50452 5764 50512 5812
rect 50206 5752 50512 5764
rect 50206 5718 50228 5752
rect 50430 5718 50512 5752
rect 50206 5704 50512 5718
rect 50945 5686 51005 5692
rect 50725 5680 50945 5686
rect 50627 5664 50687 5670
rect 50621 5604 50627 5664
rect 50687 5604 50693 5664
rect 50725 5640 50737 5680
rect 50783 5640 50945 5680
rect 50725 5626 50945 5640
rect 51005 5626 51006 5686
rect 50945 5620 51005 5626
rect 50627 5598 50687 5604
rect 49928 5448 50036 5454
rect 49928 5414 49940 5448
rect 50024 5414 50036 5448
rect 49928 5408 50036 5414
rect 49612 5188 49618 5208
rect 49572 5176 49618 5188
rect 49824 5188 49836 5364
rect 49870 5188 49884 5364
rect 50082 5364 50142 5527
rect 50212 5554 50514 5564
rect 50212 5516 50232 5554
rect 50430 5516 50514 5554
rect 50212 5504 50514 5516
rect 50212 5454 50272 5504
rect 50186 5448 50294 5454
rect 50186 5414 50198 5448
rect 50282 5414 50294 5448
rect 50186 5408 50294 5414
rect 50082 5325 50094 5364
rect 49824 5148 49884 5188
rect 50088 5188 50094 5325
rect 50128 5325 50142 5364
rect 50340 5364 50400 5504
rect 50128 5188 50134 5325
rect 50340 5318 50352 5364
rect 50346 5221 50352 5318
rect 50088 5176 50134 5188
rect 50338 5188 50352 5221
rect 50386 5318 50400 5364
rect 50454 5468 50514 5504
rect 50454 5454 50850 5468
rect 50386 5221 50392 5318
rect 50386 5188 50398 5221
rect 48896 5138 49004 5144
rect 48896 5104 48908 5138
rect 48992 5104 49004 5138
rect 48896 5098 49004 5104
rect 49154 5138 49262 5144
rect 49154 5104 49166 5138
rect 49250 5104 49262 5138
rect 49154 5098 49262 5104
rect 49412 5138 49520 5144
rect 49412 5104 49424 5138
rect 49508 5104 49520 5138
rect 49412 5098 49520 5104
rect 49670 5138 49778 5144
rect 49670 5104 49682 5138
rect 49766 5104 49778 5138
rect 49670 5098 49778 5104
rect 49928 5138 50036 5144
rect 49928 5104 49940 5138
rect 50024 5104 50036 5138
rect 49928 5098 50036 5104
rect 50186 5138 50294 5144
rect 50186 5104 50198 5138
rect 50282 5104 50294 5138
rect 50186 5098 50294 5104
rect 48920 5049 48980 5098
rect 48676 5038 48980 5049
rect 48676 5002 48758 5038
rect 48966 5002 48980 5038
rect 48676 4932 48980 5002
rect 49178 5039 49238 5098
rect 49438 5039 49498 5098
rect 49696 5039 49756 5098
rect 49952 5039 50012 5098
rect 50210 5049 50270 5098
rect 50338 5049 50398 5188
rect 50454 5098 50464 5454
rect 50502 5437 50850 5454
rect 50502 5403 50603 5437
rect 50637 5403 50695 5437
rect 50729 5403 50787 5437
rect 50821 5403 50850 5437
rect 50502 5372 50850 5403
rect 50502 5098 50514 5372
rect 50454 5049 50514 5098
rect 49178 4979 49952 5039
rect 50012 4979 50018 5039
rect 50210 5036 50514 5049
rect 50210 5000 50230 5036
rect 50432 5000 50514 5036
rect 48677 4914 48980 4932
rect 50210 4914 50514 5000
rect 52622 4914 52628 6818
rect 48677 4854 52628 4914
rect 48494 4550 50513 4610
rect 48494 2520 48554 4550
rect 48677 4484 48982 4550
rect 48677 4450 48736 4484
rect 48956 4450 48982 4484
rect 48677 4436 48982 4450
rect 48677 4386 48738 4436
rect 48677 4356 48688 4386
rect 48678 4128 48688 4356
rect 48677 4068 48688 4128
rect 48678 3814 48688 4068
rect 48726 4128 48738 4386
rect 48788 4288 48848 4436
rect 48922 4387 48982 4436
rect 49178 4502 49238 4503
rect 49954 4502 50014 4508
rect 49178 4442 49954 4502
rect 49178 4387 49238 4442
rect 49436 4387 49496 4442
rect 49694 4387 49754 4442
rect 49954 4387 50014 4442
rect 50210 4484 50513 4550
rect 50210 4450 50228 4484
rect 50430 4450 50513 4484
rect 50210 4436 50513 4450
rect 50210 4387 50270 4436
rect 48896 4381 49004 4387
rect 48896 4347 48908 4381
rect 48992 4347 49004 4381
rect 48896 4341 49004 4347
rect 49154 4381 49262 4387
rect 49154 4347 49166 4381
rect 49250 4347 49262 4381
rect 49154 4341 49262 4347
rect 49412 4381 49520 4387
rect 49412 4347 49424 4381
rect 49508 4347 49520 4381
rect 49412 4341 49520 4347
rect 49670 4381 49778 4387
rect 49670 4347 49682 4381
rect 49766 4347 49778 4381
rect 49670 4341 49778 4347
rect 49928 4381 50036 4387
rect 49928 4347 49940 4381
rect 50024 4347 50036 4381
rect 49928 4341 50036 4347
rect 50186 4381 50294 4387
rect 50186 4347 50198 4381
rect 50282 4347 50294 4381
rect 50186 4341 50294 4347
rect 48788 4128 48804 4288
rect 48726 4068 48804 4128
rect 48726 3814 48738 4068
rect 48798 3946 48804 4068
rect 48678 3764 48738 3814
rect 48790 3912 48804 3946
rect 48838 4068 48848 4288
rect 49056 4288 49102 4300
rect 48838 3946 48844 4068
rect 49056 3957 49062 4288
rect 48838 3912 48850 3946
rect 48790 3764 48850 3912
rect 49048 3912 49062 3957
rect 49096 3957 49102 4288
rect 49314 4288 49360 4300
rect 49096 3912 49108 3957
rect 49314 3932 49320 4288
rect 48896 3853 49004 3859
rect 48896 3819 48908 3853
rect 48992 3819 49004 3853
rect 48896 3813 49004 3819
rect 48918 3764 48978 3813
rect 48677 3750 48978 3764
rect 48677 3716 48736 3750
rect 48956 3716 48978 3750
rect 48677 3704 48978 3716
rect 49048 3587 49108 3912
rect 49306 3912 49320 3932
rect 49354 3932 49360 4288
rect 49572 4288 49618 4300
rect 49572 3955 49578 4288
rect 49354 3912 49366 3932
rect 49154 3853 49262 3859
rect 49154 3819 49166 3853
rect 49250 3819 49262 3853
rect 49154 3813 49262 3819
rect 49306 3736 49366 3912
rect 49564 3912 49578 3955
rect 49612 3955 49618 4288
rect 49830 4288 49876 4300
rect 49612 3912 49624 3955
rect 49830 3950 49836 4288
rect 49412 3853 49520 3859
rect 49412 3819 49424 3853
rect 49508 3819 49520 3853
rect 49412 3813 49520 3819
rect 49300 3676 49306 3736
rect 49366 3676 49372 3736
rect 48676 3552 48980 3562
rect 48676 3514 48760 3552
rect 48968 3514 48980 3552
rect 49042 3527 49048 3587
rect 49108 3527 49114 3587
rect 48676 3502 48980 3514
rect 48676 3454 48736 3502
rect 48676 3098 48688 3454
rect 48724 3098 48736 3454
rect 48790 3364 48850 3502
rect 48920 3454 48980 3502
rect 48896 3448 49004 3454
rect 48896 3414 48908 3448
rect 48992 3414 49004 3448
rect 48896 3408 49004 3414
rect 48790 3314 48804 3364
rect 48798 3227 48804 3314
rect 48676 3049 48736 3098
rect 48792 3188 48804 3227
rect 48838 3314 48850 3364
rect 49048 3364 49108 3527
rect 49154 3448 49262 3454
rect 49154 3414 49166 3448
rect 49250 3414 49262 3448
rect 49154 3408 49262 3414
rect 49048 3327 49062 3364
rect 48838 3227 48844 3314
rect 48838 3188 48852 3227
rect 48792 3049 48852 3188
rect 49056 3188 49062 3327
rect 49096 3327 49108 3364
rect 49306 3394 49366 3676
rect 49564 3587 49624 3912
rect 49824 3912 49836 3950
rect 49870 3950 49876 4288
rect 50088 4288 50134 4300
rect 50088 3955 50094 4288
rect 49870 3912 49884 3950
rect 49670 3853 49778 3859
rect 49670 3819 49682 3853
rect 49766 3819 49778 3853
rect 49670 3813 49778 3819
rect 49824 3736 49884 3912
rect 50082 3912 50094 3955
rect 50128 3955 50134 4288
rect 50338 4288 50398 4436
rect 50338 4070 50352 4288
rect 50128 3912 50142 3955
rect 50346 3942 50352 4070
rect 49928 3853 50036 3859
rect 49928 3819 49940 3853
rect 50024 3819 50036 3853
rect 49928 3813 50036 3819
rect 49818 3676 49824 3736
rect 49884 3676 49890 3736
rect 49558 3527 49564 3587
rect 49624 3527 49630 3587
rect 49412 3448 49520 3454
rect 49412 3414 49424 3448
rect 49508 3414 49520 3448
rect 49412 3408 49520 3414
rect 49306 3364 49368 3394
rect 49306 3328 49320 3364
rect 49096 3188 49102 3327
rect 49056 3176 49102 3188
rect 49308 3188 49320 3328
rect 49354 3188 49368 3364
rect 49564 3364 49624 3527
rect 49670 3448 49778 3454
rect 49670 3414 49682 3448
rect 49766 3414 49778 3448
rect 49670 3408 49778 3414
rect 49564 3208 49578 3364
rect 49308 3148 49368 3188
rect 49572 3188 49578 3208
rect 49612 3208 49624 3364
rect 49824 3364 49884 3676
rect 50082 3587 50142 3912
rect 50340 3912 50352 3942
rect 50386 4130 50398 4288
rect 50452 4388 50513 4436
rect 50452 4130 50464 4388
rect 50386 4070 50464 4130
rect 50386 3942 50392 4070
rect 50386 3912 50400 3942
rect 50186 3853 50294 3859
rect 50186 3819 50198 3853
rect 50282 3819 50294 3853
rect 50186 3813 50294 3819
rect 50206 3764 50266 3813
rect 50340 3764 50400 3912
rect 50452 3812 50464 4070
rect 50500 4372 50513 4388
rect 50500 4012 50512 4372
rect 50500 3981 50850 4012
rect 50500 3947 50603 3981
rect 50637 3947 50695 3981
rect 50729 3947 50787 3981
rect 50821 3947 50850 3981
rect 50500 3916 50850 3947
rect 50500 3812 50512 3916
rect 50452 3764 50512 3812
rect 50206 3752 50512 3764
rect 50206 3718 50228 3752
rect 50430 3718 50512 3752
rect 50206 3704 50512 3718
rect 50945 3686 51005 3692
rect 50725 3680 50945 3686
rect 50627 3664 50687 3670
rect 50621 3604 50627 3664
rect 50687 3604 50693 3664
rect 50725 3640 50737 3680
rect 50783 3640 50945 3680
rect 50725 3626 50945 3640
rect 50945 3620 51005 3626
rect 50627 3598 50687 3604
rect 49928 3448 50036 3454
rect 49928 3414 49940 3448
rect 50024 3414 50036 3448
rect 49928 3408 50036 3414
rect 49612 3188 49618 3208
rect 49572 3176 49618 3188
rect 49824 3188 49836 3364
rect 49870 3188 49884 3364
rect 50082 3364 50142 3527
rect 50212 3554 50514 3564
rect 50212 3516 50232 3554
rect 50430 3516 50514 3554
rect 50212 3504 50514 3516
rect 50212 3454 50272 3504
rect 50186 3448 50294 3454
rect 50186 3414 50198 3448
rect 50282 3414 50294 3448
rect 50186 3408 50294 3414
rect 50082 3325 50094 3364
rect 49824 3148 49884 3188
rect 50088 3188 50094 3325
rect 50128 3325 50142 3364
rect 50340 3364 50400 3504
rect 50128 3188 50134 3325
rect 50340 3318 50352 3364
rect 50346 3221 50352 3318
rect 50088 3176 50134 3188
rect 50338 3188 50352 3221
rect 50386 3318 50400 3364
rect 50454 3468 50514 3504
rect 50454 3454 50850 3468
rect 50386 3221 50392 3318
rect 50386 3188 50398 3221
rect 48896 3138 49004 3144
rect 48896 3104 48908 3138
rect 48992 3104 49004 3138
rect 48896 3098 49004 3104
rect 49154 3138 49262 3144
rect 49154 3104 49166 3138
rect 49250 3104 49262 3138
rect 49154 3098 49262 3104
rect 49412 3138 49520 3144
rect 49412 3104 49424 3138
rect 49508 3104 49520 3138
rect 49412 3098 49520 3104
rect 49670 3138 49778 3144
rect 49670 3104 49682 3138
rect 49766 3104 49778 3138
rect 49670 3098 49778 3104
rect 49928 3138 50036 3144
rect 49928 3104 49940 3138
rect 50024 3104 50036 3138
rect 49928 3098 50036 3104
rect 50186 3138 50294 3144
rect 50186 3104 50198 3138
rect 50282 3104 50294 3138
rect 50186 3098 50294 3104
rect 48920 3049 48980 3098
rect 48676 3038 48980 3049
rect 48676 3002 48758 3038
rect 48966 3002 48980 3038
rect 48676 2932 48980 3002
rect 49178 3039 49238 3098
rect 49438 3039 49498 3098
rect 49696 3039 49756 3098
rect 49952 3039 50012 3098
rect 50210 3049 50270 3098
rect 50338 3049 50398 3188
rect 50454 3098 50464 3454
rect 50502 3437 50850 3454
rect 50502 3403 50603 3437
rect 50637 3403 50695 3437
rect 50729 3403 50787 3437
rect 50821 3403 50850 3437
rect 50502 3372 50850 3403
rect 50502 3098 50514 3372
rect 50454 3049 50514 3098
rect 49178 2979 49952 3039
rect 50012 2979 50018 3039
rect 50210 3036 50514 3049
rect 50210 3000 50230 3036
rect 50432 3000 50514 3036
rect 48677 2914 48980 2932
rect 50210 2914 50514 3000
rect 52622 2914 52628 4854
rect 48677 2854 52628 2914
rect 48494 2462 50513 2520
rect 48498 2460 50513 2462
rect 48677 2394 48982 2460
rect 48677 2360 48736 2394
rect 48956 2360 48982 2394
rect 48677 2346 48982 2360
rect 48677 2296 48738 2346
rect 48677 2266 48688 2296
rect 48678 2038 48688 2266
rect 48677 1978 48688 2038
rect 48678 1724 48688 1978
rect 48726 2038 48738 2296
rect 48788 2198 48848 2346
rect 48922 2297 48982 2346
rect 49178 2412 49238 2413
rect 49954 2412 50014 2418
rect 49178 2352 49954 2412
rect 49178 2297 49238 2352
rect 49436 2297 49496 2352
rect 49694 2297 49754 2352
rect 49954 2297 50014 2352
rect 50210 2394 50513 2460
rect 50210 2360 50228 2394
rect 50430 2360 50513 2394
rect 50210 2346 50513 2360
rect 50210 2297 50270 2346
rect 48896 2291 49004 2297
rect 48896 2257 48908 2291
rect 48992 2257 49004 2291
rect 48896 2251 49004 2257
rect 49154 2291 49262 2297
rect 49154 2257 49166 2291
rect 49250 2257 49262 2291
rect 49154 2251 49262 2257
rect 49412 2291 49520 2297
rect 49412 2257 49424 2291
rect 49508 2257 49520 2291
rect 49412 2251 49520 2257
rect 49670 2291 49778 2297
rect 49670 2257 49682 2291
rect 49766 2257 49778 2291
rect 49670 2251 49778 2257
rect 49928 2291 50036 2297
rect 49928 2257 49940 2291
rect 50024 2257 50036 2291
rect 49928 2251 50036 2257
rect 50186 2291 50294 2297
rect 50186 2257 50198 2291
rect 50282 2257 50294 2291
rect 50186 2251 50294 2257
rect 48788 2038 48804 2198
rect 48726 1978 48804 2038
rect 48726 1724 48738 1978
rect 48798 1856 48804 1978
rect 48678 1674 48738 1724
rect 48790 1822 48804 1856
rect 48838 1978 48848 2198
rect 49056 2198 49102 2210
rect 48838 1856 48844 1978
rect 49056 1867 49062 2198
rect 48838 1822 48850 1856
rect 48790 1674 48850 1822
rect 49048 1822 49062 1867
rect 49096 1867 49102 2198
rect 49314 2198 49360 2210
rect 49096 1822 49108 1867
rect 49314 1842 49320 2198
rect 48896 1763 49004 1769
rect 48896 1729 48908 1763
rect 48992 1729 49004 1763
rect 48896 1723 49004 1729
rect 48918 1674 48978 1723
rect 48677 1660 48978 1674
rect 48677 1626 48736 1660
rect 48956 1626 48978 1660
rect 48677 1614 48978 1626
rect 49048 1497 49108 1822
rect 49306 1822 49320 1842
rect 49354 1842 49360 2198
rect 49572 2198 49618 2210
rect 49572 1865 49578 2198
rect 49354 1822 49366 1842
rect 49154 1763 49262 1769
rect 49154 1729 49166 1763
rect 49250 1729 49262 1763
rect 49154 1723 49262 1729
rect 49306 1646 49366 1822
rect 49564 1822 49578 1865
rect 49612 1865 49618 2198
rect 49830 2198 49876 2210
rect 49612 1822 49624 1865
rect 49830 1860 49836 2198
rect 49412 1763 49520 1769
rect 49412 1729 49424 1763
rect 49508 1729 49520 1763
rect 49412 1723 49520 1729
rect 49300 1586 49306 1646
rect 49366 1586 49372 1646
rect 48676 1462 48980 1472
rect 48676 1424 48760 1462
rect 48968 1424 48980 1462
rect 49042 1437 49048 1497
rect 49108 1437 49114 1497
rect 48676 1412 48980 1424
rect 48676 1364 48736 1412
rect 48676 1008 48688 1364
rect 48724 1008 48736 1364
rect 48790 1274 48850 1412
rect 48920 1364 48980 1412
rect 48896 1358 49004 1364
rect 48896 1324 48908 1358
rect 48992 1324 49004 1358
rect 48896 1318 49004 1324
rect 48790 1224 48804 1274
rect 48798 1137 48804 1224
rect 48676 959 48736 1008
rect 48792 1098 48804 1137
rect 48838 1224 48850 1274
rect 49048 1274 49108 1437
rect 49154 1358 49262 1364
rect 49154 1324 49166 1358
rect 49250 1324 49262 1358
rect 49154 1318 49262 1324
rect 49048 1237 49062 1274
rect 48838 1137 48844 1224
rect 48838 1098 48852 1137
rect 48792 959 48852 1098
rect 49056 1098 49062 1237
rect 49096 1237 49108 1274
rect 49306 1304 49366 1586
rect 49564 1497 49624 1822
rect 49824 1822 49836 1860
rect 49870 1860 49876 2198
rect 50088 2198 50134 2210
rect 50088 1865 50094 2198
rect 49870 1822 49884 1860
rect 49670 1763 49778 1769
rect 49670 1729 49682 1763
rect 49766 1729 49778 1763
rect 49670 1723 49778 1729
rect 49824 1646 49884 1822
rect 50082 1822 50094 1865
rect 50128 1865 50134 2198
rect 50338 2198 50398 2346
rect 50338 1980 50352 2198
rect 50128 1822 50142 1865
rect 50346 1852 50352 1980
rect 49928 1763 50036 1769
rect 49928 1729 49940 1763
rect 50024 1729 50036 1763
rect 49928 1723 50036 1729
rect 49818 1586 49824 1646
rect 49884 1586 49890 1646
rect 49558 1437 49564 1497
rect 49624 1437 49630 1497
rect 49412 1358 49520 1364
rect 49412 1324 49424 1358
rect 49508 1324 49520 1358
rect 49412 1318 49520 1324
rect 49306 1274 49368 1304
rect 49306 1238 49320 1274
rect 49096 1098 49102 1237
rect 49056 1086 49102 1098
rect 49308 1098 49320 1238
rect 49354 1098 49368 1274
rect 49564 1274 49624 1437
rect 49670 1358 49778 1364
rect 49670 1324 49682 1358
rect 49766 1324 49778 1358
rect 49670 1318 49778 1324
rect 49564 1118 49578 1274
rect 49308 1058 49368 1098
rect 49572 1098 49578 1118
rect 49612 1118 49624 1274
rect 49824 1274 49884 1586
rect 50082 1497 50142 1822
rect 50340 1822 50352 1852
rect 50386 2040 50398 2198
rect 50452 2298 50513 2346
rect 50452 2040 50464 2298
rect 50386 1980 50464 2040
rect 50386 1852 50392 1980
rect 50386 1822 50400 1852
rect 50186 1763 50294 1769
rect 50186 1729 50198 1763
rect 50282 1729 50294 1763
rect 50186 1723 50294 1729
rect 50206 1674 50266 1723
rect 50340 1674 50400 1822
rect 50452 1722 50464 1980
rect 50500 2282 50513 2298
rect 50500 1922 50512 2282
rect 50500 1891 50850 1922
rect 50500 1857 50603 1891
rect 50637 1857 50695 1891
rect 50729 1857 50787 1891
rect 50821 1857 50850 1891
rect 50500 1826 50850 1857
rect 50500 1722 50512 1826
rect 50452 1674 50512 1722
rect 50206 1662 50512 1674
rect 50206 1628 50228 1662
rect 50430 1628 50512 1662
rect 50206 1614 50512 1628
rect 50945 1596 51005 1602
rect 50725 1590 50945 1596
rect 50627 1574 50687 1580
rect 50621 1514 50627 1574
rect 50687 1514 50693 1574
rect 50725 1550 50737 1590
rect 50783 1550 50945 1590
rect 50725 1536 50945 1550
rect 50945 1530 51005 1536
rect 50627 1508 50687 1514
rect 49928 1358 50036 1364
rect 49928 1324 49940 1358
rect 50024 1324 50036 1358
rect 49928 1318 50036 1324
rect 49612 1098 49618 1118
rect 49572 1086 49618 1098
rect 49824 1098 49836 1274
rect 49870 1098 49884 1274
rect 50082 1274 50142 1437
rect 50212 1464 50514 1474
rect 50212 1426 50232 1464
rect 50430 1426 50514 1464
rect 50212 1414 50514 1426
rect 50212 1364 50272 1414
rect 50186 1358 50294 1364
rect 50186 1324 50198 1358
rect 50282 1324 50294 1358
rect 50186 1318 50294 1324
rect 50082 1235 50094 1274
rect 49824 1058 49884 1098
rect 50088 1098 50094 1235
rect 50128 1235 50142 1274
rect 50340 1274 50400 1414
rect 50128 1098 50134 1235
rect 50340 1228 50352 1274
rect 50346 1131 50352 1228
rect 50088 1086 50134 1098
rect 50338 1098 50352 1131
rect 50386 1228 50400 1274
rect 50454 1378 50514 1414
rect 50454 1364 50850 1378
rect 50386 1131 50392 1228
rect 50386 1098 50398 1131
rect 48896 1048 49004 1054
rect 48896 1014 48908 1048
rect 48992 1014 49004 1048
rect 48896 1008 49004 1014
rect 49154 1048 49262 1054
rect 49154 1014 49166 1048
rect 49250 1014 49262 1048
rect 49154 1008 49262 1014
rect 49412 1048 49520 1054
rect 49412 1014 49424 1048
rect 49508 1014 49520 1048
rect 49412 1008 49520 1014
rect 49670 1048 49778 1054
rect 49670 1014 49682 1048
rect 49766 1014 49778 1048
rect 49670 1008 49778 1014
rect 49928 1048 50036 1054
rect 49928 1014 49940 1048
rect 50024 1014 50036 1048
rect 49928 1008 50036 1014
rect 50186 1048 50294 1054
rect 50186 1014 50198 1048
rect 50282 1014 50294 1048
rect 50186 1008 50294 1014
rect 48920 959 48980 1008
rect 48676 948 48980 959
rect 48676 912 48758 948
rect 48966 912 48980 948
rect 48676 842 48980 912
rect 49178 949 49238 1008
rect 49438 949 49498 1008
rect 49696 949 49756 1008
rect 49952 949 50012 1008
rect 50210 959 50270 1008
rect 50338 959 50398 1098
rect 50454 1008 50464 1364
rect 50502 1347 50850 1364
rect 50502 1313 50603 1347
rect 50637 1313 50695 1347
rect 50729 1313 50787 1347
rect 50821 1313 50850 1347
rect 50502 1282 50850 1313
rect 50502 1008 50514 1282
rect 50454 959 50514 1008
rect 49178 889 49952 949
rect 50012 889 50018 949
rect 50210 946 50514 959
rect 50210 910 50230 946
rect 50432 910 50514 946
rect 48677 824 48980 842
rect 50210 824 50514 910
rect 52622 824 52628 2854
rect 48677 764 52628 824
rect 3432 64 34918 110
rect 3432 -90 3478 64
rect 34878 -90 34918 64
rect 3432 -136 34918 -90
rect -666 -576 -656 -276
rect 35156 -576 35166 -276
rect 35766 -576 35878 210
rect -1378 -582 35878 -576
rect -1378 -682 -1272 -582
rect 35772 -682 35878 -582
rect -1378 -688 35878 -682
rect 52622 210 52628 764
rect 52728 210 52734 14470
rect 66904 14354 66964 15132
rect 62878 14294 66964 14354
rect 62878 14216 62938 14294
rect 55754 14156 62938 14216
rect 55754 14016 55814 14156
rect 56264 14106 56324 14156
rect 56048 14100 56536 14106
rect 56048 14066 56060 14100
rect 56524 14066 56536 14100
rect 56048 14060 56536 14066
rect 55754 13986 55766 14016
rect 55760 13458 55766 13986
rect 55750 13440 55766 13458
rect 55800 13986 55814 14016
rect 56770 14016 56830 14156
rect 57272 14106 57332 14156
rect 58300 14106 58360 14156
rect 57066 14100 57554 14106
rect 57066 14066 57078 14100
rect 57542 14066 57554 14100
rect 57066 14060 57554 14066
rect 58084 14100 58572 14106
rect 58084 14066 58096 14100
rect 58560 14066 58572 14100
rect 58084 14060 58572 14066
rect 56770 13992 56784 14016
rect 55800 13458 55806 13986
rect 56778 13462 56784 13992
rect 55800 13440 55810 13458
rect 55750 13198 55810 13440
rect 56770 13440 56784 13462
rect 56818 13992 56830 14016
rect 57796 14016 57842 14028
rect 56818 13462 56824 13992
rect 57796 13464 57802 14016
rect 56818 13440 56830 13462
rect 56048 13390 56536 13396
rect 56048 13356 56060 13390
rect 56524 13356 56536 13390
rect 56048 13350 56536 13356
rect 56264 13288 56324 13350
rect 56048 13282 56536 13288
rect 56048 13248 56060 13282
rect 56524 13248 56536 13282
rect 56048 13242 56536 13248
rect 55750 13168 55766 13198
rect 55760 12644 55766 13168
rect 55752 12622 55766 12644
rect 55800 13168 55810 13198
rect 56770 13198 56830 13440
rect 57790 13440 57802 13464
rect 57836 13464 57842 14016
rect 58808 14016 58868 14156
rect 59314 14106 59374 14156
rect 60328 14106 60388 14156
rect 59102 14100 59590 14106
rect 59102 14066 59114 14100
rect 59578 14066 59590 14100
rect 59102 14060 59590 14066
rect 60120 14100 60608 14106
rect 60120 14066 60132 14100
rect 60596 14066 60608 14100
rect 60120 14060 60608 14066
rect 58808 13978 58820 14016
rect 57836 13440 57850 13464
rect 58814 13460 58820 13978
rect 57066 13390 57554 13396
rect 57066 13356 57078 13390
rect 57542 13356 57554 13390
rect 57066 13350 57554 13356
rect 57268 13288 57328 13350
rect 57066 13282 57554 13288
rect 57066 13248 57078 13282
rect 57542 13248 57554 13282
rect 57066 13242 57554 13248
rect 56770 13172 56784 13198
rect 55800 12644 55806 13168
rect 56778 12648 56784 13172
rect 55800 12622 55812 12644
rect 55752 12380 55812 12622
rect 56772 12622 56784 12648
rect 56818 13172 56830 13198
rect 57790 13198 57850 13440
rect 58808 13440 58820 13460
rect 58854 13978 58868 14016
rect 59832 14016 59878 14028
rect 60844 14016 60904 14156
rect 61360 14106 61420 14156
rect 62366 14106 62426 14156
rect 61138 14100 61626 14106
rect 61138 14066 61150 14100
rect 61614 14066 61626 14100
rect 61138 14060 61626 14066
rect 62156 14100 62644 14106
rect 62156 14066 62168 14100
rect 62632 14066 62644 14100
rect 62156 14060 62644 14066
rect 58854 13460 58860 13978
rect 59832 13468 59838 14016
rect 58854 13440 58868 13460
rect 58084 13390 58572 13396
rect 58084 13356 58096 13390
rect 58560 13356 58572 13390
rect 58084 13350 58572 13356
rect 58298 13288 58358 13350
rect 58084 13282 58572 13288
rect 58084 13248 58096 13282
rect 58560 13248 58572 13282
rect 58084 13242 58572 13248
rect 57790 13174 57802 13198
rect 56818 12648 56824 13172
rect 57796 12650 57802 13174
rect 56818 12622 56832 12648
rect 56048 12572 56536 12578
rect 56048 12538 56060 12572
rect 56524 12538 56536 12572
rect 56048 12532 56536 12538
rect 56264 12470 56324 12532
rect 56048 12464 56536 12470
rect 56048 12430 56060 12464
rect 56524 12430 56536 12464
rect 56048 12424 56536 12430
rect 55752 12354 55766 12380
rect 55760 11816 55766 12354
rect 55752 11804 55766 11816
rect 55800 12354 55812 12380
rect 56772 12380 56832 12622
rect 57792 12622 57802 12650
rect 57836 13174 57850 13198
rect 58808 13198 58868 13440
rect 59828 13440 59838 13468
rect 59872 13468 59878 14016
rect 60842 13982 60856 14016
rect 60844 13970 60856 13982
rect 59872 13440 59888 13468
rect 60850 13460 60856 13970
rect 59102 13390 59590 13396
rect 59102 13356 59114 13390
rect 59578 13356 59590 13390
rect 59102 13350 59590 13356
rect 59300 13288 59360 13350
rect 59102 13282 59590 13288
rect 59102 13248 59114 13282
rect 59578 13248 59590 13282
rect 59102 13242 59590 13248
rect 57836 12650 57842 13174
rect 58808 13170 58820 13198
rect 57836 12622 57852 12650
rect 58814 12646 58820 13170
rect 57066 12572 57554 12578
rect 57066 12538 57078 12572
rect 57542 12538 57554 12572
rect 57066 12532 57554 12538
rect 57280 12470 57340 12532
rect 57066 12464 57554 12470
rect 57066 12430 57078 12464
rect 57542 12430 57554 12464
rect 57066 12424 57554 12430
rect 56772 12358 56784 12380
rect 55800 11816 55806 12354
rect 56778 11820 56784 12358
rect 55800 11804 55812 11816
rect 55752 11562 55812 11804
rect 56772 11804 56784 11820
rect 56818 12358 56832 12380
rect 57792 12380 57852 12622
rect 58810 12622 58820 12646
rect 58854 13170 58868 13198
rect 59828 13198 59888 13440
rect 60840 13440 60856 13460
rect 60890 13970 60904 14016
rect 61868 14016 61914 14028
rect 60890 13460 60896 13970
rect 61868 13460 61874 14016
rect 60890 13440 60900 13460
rect 60120 13390 60608 13396
rect 60120 13356 60132 13390
rect 60596 13356 60608 13390
rect 60120 13350 60608 13356
rect 60330 13288 60390 13350
rect 60120 13282 60608 13288
rect 60120 13248 60132 13282
rect 60596 13248 60608 13282
rect 60120 13242 60608 13248
rect 59828 13178 59838 13198
rect 58854 12646 58860 13170
rect 59832 12654 59838 13178
rect 58854 12622 58870 12646
rect 58084 12572 58572 12578
rect 58084 12538 58096 12572
rect 58560 12538 58572 12572
rect 58084 12532 58572 12538
rect 58298 12470 58358 12532
rect 58084 12464 58572 12470
rect 58084 12430 58096 12464
rect 58560 12430 58572 12464
rect 58084 12424 58572 12430
rect 57792 12360 57802 12380
rect 56818 11820 56824 12358
rect 57796 11822 57802 12360
rect 56818 11804 56832 11820
rect 56048 11754 56536 11760
rect 56048 11720 56060 11754
rect 56524 11720 56536 11754
rect 56048 11714 56536 11720
rect 56258 11652 56318 11714
rect 56048 11646 56536 11652
rect 56048 11612 56060 11646
rect 56524 11612 56536 11646
rect 56048 11606 56536 11612
rect 55752 11526 55766 11562
rect 55760 11004 55766 11526
rect 55752 10986 55766 11004
rect 55800 11526 55812 11562
rect 56772 11562 56832 11804
rect 57792 11804 57802 11822
rect 57836 12360 57852 12380
rect 58810 12380 58870 12622
rect 59830 12622 59838 12654
rect 59872 13178 59888 13198
rect 60840 13198 60900 13440
rect 61862 13440 61874 13460
rect 61908 13460 61914 14016
rect 62878 14016 62938 14156
rect 63388 14106 63448 14294
rect 66134 14206 66194 14212
rect 64918 14146 66134 14206
rect 63174 14100 63662 14106
rect 63174 14066 63186 14100
rect 63650 14066 63662 14100
rect 63174 14060 63662 14066
rect 64192 14100 64680 14106
rect 64192 14066 64204 14100
rect 64668 14066 64680 14100
rect 64192 14060 64680 14066
rect 62878 13980 62892 14016
rect 62886 13460 62892 13980
rect 61908 13440 61922 13460
rect 61138 13390 61626 13396
rect 61138 13356 61150 13390
rect 61614 13356 61626 13390
rect 61138 13350 61626 13356
rect 61346 13288 61406 13350
rect 61138 13282 61626 13288
rect 61138 13248 61150 13282
rect 61614 13248 61626 13282
rect 61138 13242 61626 13248
rect 59872 12654 59878 13178
rect 60840 13170 60856 13198
rect 59872 12622 59890 12654
rect 60850 12646 60856 13170
rect 59102 12572 59590 12578
rect 59102 12538 59114 12572
rect 59578 12538 59590 12572
rect 59102 12532 59590 12538
rect 59300 12470 59360 12532
rect 59102 12464 59590 12470
rect 59102 12430 59114 12464
rect 59578 12430 59590 12464
rect 59102 12424 59590 12430
rect 57836 11822 57842 12360
rect 58810 12356 58820 12380
rect 57836 11804 57852 11822
rect 58814 11818 58820 12356
rect 57066 11754 57554 11760
rect 57066 11720 57078 11754
rect 57542 11720 57554 11754
rect 57066 11714 57554 11720
rect 57280 11652 57340 11714
rect 57066 11646 57554 11652
rect 57066 11612 57078 11646
rect 57542 11612 57554 11646
rect 57066 11606 57554 11612
rect 56772 11530 56784 11562
rect 55800 11004 55806 11526
rect 56778 11008 56784 11530
rect 55800 10986 55812 11004
rect 55752 10744 55812 10986
rect 56772 10986 56784 11008
rect 56818 11530 56832 11562
rect 57792 11562 57852 11804
rect 58810 11804 58820 11818
rect 58854 12356 58870 12380
rect 59830 12380 59890 12622
rect 60842 12622 60856 12646
rect 60890 13170 60900 13198
rect 61862 13198 61922 13440
rect 62882 13440 62892 13460
rect 62926 13980 62938 14016
rect 63904 14016 63950 14028
rect 62926 13460 62932 13980
rect 63904 13464 63910 14016
rect 62926 13440 62942 13460
rect 62156 13390 62644 13396
rect 62156 13356 62168 13390
rect 62632 13356 62644 13390
rect 62156 13350 62644 13356
rect 62368 13288 62428 13350
rect 62156 13282 62644 13288
rect 62156 13248 62168 13282
rect 62632 13248 62644 13282
rect 62156 13242 62644 13248
rect 61862 13170 61874 13198
rect 60890 12646 60896 13170
rect 61868 12646 61874 13170
rect 60890 12622 60902 12646
rect 60120 12572 60608 12578
rect 60120 12538 60132 12572
rect 60596 12538 60608 12572
rect 60120 12532 60608 12538
rect 60330 12470 60390 12532
rect 60120 12464 60608 12470
rect 60120 12430 60132 12464
rect 60596 12430 60608 12464
rect 60120 12424 60608 12430
rect 59830 12364 59838 12380
rect 58854 11818 58860 12356
rect 59832 11826 59838 12364
rect 58854 11804 58870 11818
rect 58084 11754 58572 11760
rect 58084 11720 58096 11754
rect 58560 11720 58572 11754
rect 58084 11714 58572 11720
rect 58292 11652 58352 11714
rect 58084 11646 58572 11652
rect 58084 11612 58096 11646
rect 58560 11612 58572 11646
rect 58084 11606 58572 11612
rect 57792 11532 57802 11562
rect 56818 11008 56824 11530
rect 57796 11010 57802 11532
rect 56818 10986 56832 11008
rect 56048 10936 56536 10942
rect 56048 10902 56060 10936
rect 56524 10902 56536 10936
rect 56048 10896 56536 10902
rect 56256 10834 56316 10896
rect 56048 10828 56536 10834
rect 56048 10794 56060 10828
rect 56524 10794 56536 10828
rect 56048 10788 56536 10794
rect 55752 10714 55766 10744
rect 55760 10184 55766 10714
rect 55752 10168 55766 10184
rect 55800 10714 55812 10744
rect 56772 10744 56832 10986
rect 57792 10986 57802 11010
rect 57836 11532 57852 11562
rect 58810 11562 58870 11804
rect 59830 11804 59838 11826
rect 59872 12364 59890 12380
rect 60842 12380 60902 12622
rect 61864 12622 61874 12646
rect 61908 13170 61922 13198
rect 62882 13198 62942 13440
rect 63898 13440 63910 13464
rect 63944 13464 63950 14016
rect 64918 14016 64978 14146
rect 66134 14140 66194 14146
rect 66794 14032 66800 14092
rect 66860 14032 66866 14092
rect 64918 13964 64928 14016
rect 63944 13440 63958 13464
rect 64922 13460 64928 13964
rect 63174 13390 63662 13396
rect 63174 13356 63186 13390
rect 63650 13356 63662 13390
rect 63174 13350 63662 13356
rect 63380 13288 63440 13350
rect 63174 13282 63662 13288
rect 63174 13248 63186 13282
rect 63650 13248 63662 13282
rect 63174 13242 63662 13248
rect 62882 13170 62892 13198
rect 61908 12646 61914 13170
rect 62886 12646 62892 13170
rect 61908 12622 61924 12646
rect 61138 12572 61626 12578
rect 61138 12538 61150 12572
rect 61614 12538 61626 12572
rect 61138 12532 61626 12538
rect 61346 12470 61406 12532
rect 61138 12464 61626 12470
rect 61138 12430 61150 12464
rect 61614 12430 61626 12464
rect 61138 12424 61626 12430
rect 59872 11826 59878 12364
rect 60842 12356 60856 12380
rect 59872 11804 59890 11826
rect 60850 11818 60856 12356
rect 59102 11754 59590 11760
rect 59102 11720 59114 11754
rect 59578 11720 59590 11754
rect 59102 11714 59590 11720
rect 59294 11652 59354 11714
rect 59102 11646 59590 11652
rect 59102 11612 59114 11646
rect 59578 11612 59590 11646
rect 59102 11606 59590 11612
rect 57836 11010 57842 11532
rect 58810 11528 58820 11562
rect 57836 10986 57852 11010
rect 58814 11006 58820 11528
rect 57066 10936 57554 10942
rect 57066 10902 57078 10936
rect 57542 10902 57554 10936
rect 57066 10896 57554 10902
rect 57274 10834 57334 10896
rect 57066 10828 57554 10834
rect 57066 10794 57078 10828
rect 57542 10794 57554 10828
rect 57066 10788 57554 10794
rect 56772 10718 56784 10744
rect 55800 10184 55806 10714
rect 56778 10188 56784 10718
rect 55800 10168 55812 10184
rect 55752 9926 55812 10168
rect 56772 10168 56784 10188
rect 56818 10718 56832 10744
rect 57792 10744 57852 10986
rect 58810 10986 58820 11006
rect 58854 11528 58870 11562
rect 59830 11562 59890 11804
rect 60842 11804 60856 11818
rect 60890 12356 60902 12380
rect 61864 12380 61924 12622
rect 62884 12622 62892 12646
rect 62926 13170 62942 13198
rect 63898 13198 63958 13440
rect 64920 13440 64928 13460
rect 64962 13964 64978 14016
rect 64962 13460 64968 13964
rect 64962 13440 64980 13460
rect 64192 13390 64680 13396
rect 64192 13356 64204 13390
rect 64668 13356 64680 13390
rect 64192 13350 64680 13356
rect 64400 13288 64460 13350
rect 64192 13282 64680 13288
rect 64192 13248 64204 13282
rect 64668 13248 64680 13282
rect 64192 13242 64680 13248
rect 63898 13174 63910 13198
rect 62926 12646 62932 13170
rect 63904 12650 63910 13174
rect 62926 12622 62944 12646
rect 62156 12572 62644 12578
rect 62156 12538 62168 12572
rect 62632 12538 62644 12572
rect 62156 12532 62644 12538
rect 62368 12470 62428 12532
rect 62156 12464 62644 12470
rect 62156 12430 62168 12464
rect 62632 12430 62644 12464
rect 62156 12424 62644 12430
rect 61864 12356 61874 12380
rect 60890 11818 60896 12356
rect 61868 11818 61874 12356
rect 60890 11804 60902 11818
rect 60120 11754 60608 11760
rect 60120 11720 60132 11754
rect 60596 11720 60608 11754
rect 60120 11714 60608 11720
rect 60324 11652 60384 11714
rect 60120 11646 60608 11652
rect 60120 11612 60132 11646
rect 60596 11612 60608 11646
rect 60120 11606 60608 11612
rect 59830 11536 59838 11562
rect 58854 11006 58860 11528
rect 59832 11014 59838 11536
rect 58854 10986 58870 11006
rect 58084 10936 58572 10942
rect 58084 10902 58096 10936
rect 58560 10902 58572 10936
rect 58084 10896 58572 10902
rect 58290 10834 58350 10896
rect 58084 10828 58572 10834
rect 58084 10794 58096 10828
rect 58560 10794 58572 10828
rect 58084 10788 58572 10794
rect 57792 10720 57802 10744
rect 56818 10188 56824 10718
rect 57796 10190 57802 10720
rect 56818 10168 56832 10188
rect 56048 10118 56536 10124
rect 56048 10084 56060 10118
rect 56524 10084 56536 10118
rect 56048 10078 56536 10084
rect 56258 10016 56318 10078
rect 56048 10010 56536 10016
rect 56048 9976 56060 10010
rect 56524 9976 56536 10010
rect 56048 9970 56536 9976
rect 55752 9894 55766 9926
rect 55760 9372 55766 9894
rect 55752 9350 55766 9372
rect 55800 9894 55812 9926
rect 56772 9926 56832 10168
rect 57792 10168 57802 10190
rect 57836 10720 57852 10744
rect 58810 10744 58870 10986
rect 59830 10986 59838 11014
rect 59872 11536 59890 11562
rect 60842 11562 60902 11804
rect 61864 11804 61874 11818
rect 61908 12356 61924 12380
rect 62884 12380 62944 12622
rect 63900 12622 63910 12650
rect 63944 13174 63958 13198
rect 64920 13198 64980 13440
rect 63944 12650 63950 13174
rect 64920 13170 64928 13198
rect 63944 12622 63960 12650
rect 63174 12572 63662 12578
rect 63174 12538 63186 12572
rect 63650 12538 63662 12572
rect 63174 12532 63662 12538
rect 63380 12470 63440 12532
rect 63174 12464 63662 12470
rect 63174 12430 63186 12464
rect 63650 12430 63662 12464
rect 63174 12424 63662 12430
rect 62884 12356 62892 12380
rect 61908 11818 61914 12356
rect 62886 11818 62892 12356
rect 61908 11804 61924 11818
rect 61138 11754 61626 11760
rect 61138 11720 61150 11754
rect 61614 11720 61626 11754
rect 61138 11714 61626 11720
rect 61340 11652 61400 11714
rect 61138 11646 61626 11652
rect 61138 11612 61150 11646
rect 61614 11612 61626 11646
rect 61138 11606 61626 11612
rect 59872 11014 59878 11536
rect 60842 11528 60856 11562
rect 59872 10986 59890 11014
rect 60850 11006 60856 11528
rect 59102 10936 59590 10942
rect 59102 10902 59114 10936
rect 59578 10902 59590 10936
rect 59102 10896 59590 10902
rect 59292 10834 59352 10896
rect 59102 10828 59590 10834
rect 59102 10794 59114 10828
rect 59578 10794 59590 10828
rect 59102 10788 59590 10794
rect 57836 10190 57842 10720
rect 58810 10716 58820 10744
rect 57836 10168 57852 10190
rect 58814 10186 58820 10716
rect 57066 10118 57554 10124
rect 57066 10084 57078 10118
rect 57542 10084 57554 10118
rect 57066 10078 57554 10084
rect 57272 10016 57332 10078
rect 57066 10010 57554 10016
rect 57066 9976 57078 10010
rect 57542 9976 57554 10010
rect 57066 9970 57554 9976
rect 56772 9898 56784 9926
rect 55800 9372 55806 9894
rect 56778 9376 56784 9898
rect 55800 9350 55812 9372
rect 55752 9108 55812 9350
rect 56772 9350 56784 9376
rect 56818 9898 56832 9926
rect 57792 9926 57852 10168
rect 58810 10168 58820 10186
rect 58854 10716 58870 10744
rect 59830 10744 59890 10986
rect 60842 10986 60856 11006
rect 60890 11528 60902 11562
rect 61864 11562 61924 11804
rect 62884 11804 62892 11818
rect 62926 12356 62944 12380
rect 63900 12380 63960 12622
rect 64922 12622 64928 13170
rect 64962 13170 64980 13198
rect 64962 12646 64968 13170
rect 64962 12622 64982 12646
rect 64192 12572 64680 12578
rect 64192 12538 64204 12572
rect 64668 12538 64680 12572
rect 64192 12532 64680 12538
rect 64400 12470 64460 12532
rect 64192 12464 64680 12470
rect 64192 12430 64204 12464
rect 64668 12430 64680 12464
rect 64192 12424 64680 12430
rect 63900 12360 63910 12380
rect 62926 11818 62932 12356
rect 63904 11822 63910 12360
rect 62926 11804 62944 11818
rect 62156 11754 62644 11760
rect 62156 11720 62168 11754
rect 62632 11720 62644 11754
rect 62156 11714 62644 11720
rect 62362 11652 62422 11714
rect 62156 11646 62644 11652
rect 62156 11612 62168 11646
rect 62632 11612 62644 11646
rect 62156 11606 62644 11612
rect 61864 11528 61874 11562
rect 60890 11006 60896 11528
rect 61868 11006 61874 11528
rect 60890 10986 60902 11006
rect 60120 10936 60608 10942
rect 60120 10902 60132 10936
rect 60596 10902 60608 10936
rect 60120 10896 60608 10902
rect 60322 10834 60382 10896
rect 60120 10828 60608 10834
rect 60120 10794 60132 10828
rect 60596 10794 60608 10828
rect 60120 10788 60608 10794
rect 59830 10724 59838 10744
rect 58854 10186 58860 10716
rect 59832 10194 59838 10724
rect 58854 10168 58870 10186
rect 58084 10118 58572 10124
rect 58084 10084 58096 10118
rect 58560 10084 58572 10118
rect 58084 10078 58572 10084
rect 58292 10016 58352 10078
rect 58084 10010 58572 10016
rect 58084 9976 58096 10010
rect 58560 9976 58572 10010
rect 58084 9970 58572 9976
rect 57792 9900 57802 9926
rect 56818 9376 56824 9898
rect 57796 9378 57802 9900
rect 56818 9350 56832 9376
rect 56048 9300 56536 9306
rect 56048 9266 56060 9300
rect 56524 9266 56536 9300
rect 56048 9260 56536 9266
rect 56260 9198 56320 9260
rect 56048 9192 56536 9198
rect 56048 9158 56060 9192
rect 56524 9158 56536 9192
rect 56048 9152 56536 9158
rect 55752 9082 55766 9108
rect 55760 8554 55766 9082
rect 55752 8532 55766 8554
rect 55800 9082 55812 9108
rect 56772 9108 56832 9350
rect 57792 9350 57802 9378
rect 57836 9900 57852 9926
rect 58810 9926 58870 10168
rect 59830 10168 59838 10194
rect 59872 10724 59890 10744
rect 60842 10744 60902 10986
rect 61864 10986 61874 11006
rect 61908 11528 61924 11562
rect 62884 11562 62944 11804
rect 63900 11804 63910 11822
rect 63944 12360 63960 12380
rect 64922 12380 64982 12622
rect 63944 11822 63950 12360
rect 63944 11804 63960 11822
rect 63174 11754 63662 11760
rect 63174 11720 63186 11754
rect 63650 11720 63662 11754
rect 63174 11714 63662 11720
rect 63374 11652 63434 11714
rect 63174 11646 63662 11652
rect 63174 11612 63186 11646
rect 63650 11612 63662 11646
rect 63174 11606 63662 11612
rect 62884 11528 62892 11562
rect 61908 11006 61914 11528
rect 62886 11006 62892 11528
rect 61908 10986 61924 11006
rect 61138 10936 61626 10942
rect 61138 10902 61150 10936
rect 61614 10902 61626 10936
rect 61138 10896 61626 10902
rect 61338 10834 61398 10896
rect 61138 10828 61626 10834
rect 61138 10794 61150 10828
rect 61614 10794 61626 10828
rect 61138 10788 61626 10794
rect 59872 10194 59878 10724
rect 60842 10716 60856 10744
rect 59872 10168 59890 10194
rect 60850 10186 60856 10716
rect 59102 10118 59590 10124
rect 59102 10084 59114 10118
rect 59578 10084 59590 10118
rect 59102 10078 59590 10084
rect 59294 10016 59354 10078
rect 59102 10010 59590 10016
rect 59102 9976 59114 10010
rect 59578 9976 59590 10010
rect 59102 9970 59590 9976
rect 57836 9378 57842 9900
rect 58810 9896 58820 9926
rect 57836 9350 57852 9378
rect 58814 9374 58820 9896
rect 57066 9300 57554 9306
rect 57066 9266 57078 9300
rect 57542 9266 57554 9300
rect 57066 9260 57554 9266
rect 57274 9198 57334 9260
rect 57066 9192 57554 9198
rect 57066 9158 57078 9192
rect 57542 9158 57554 9192
rect 57066 9152 57554 9158
rect 56772 9086 56784 9108
rect 55800 8554 55806 9082
rect 56778 8558 56784 9086
rect 55800 8532 55812 8554
rect 55752 8290 55812 8532
rect 56772 8532 56784 8558
rect 56818 9086 56832 9108
rect 57792 9108 57852 9350
rect 58810 9350 58820 9374
rect 58854 9896 58870 9926
rect 59830 9926 59890 10168
rect 60842 10168 60856 10186
rect 60890 10716 60902 10744
rect 61864 10744 61924 10986
rect 62884 10986 62892 11006
rect 62926 11528 62944 11562
rect 63900 11562 63960 11804
rect 64922 11804 64928 12380
rect 64962 12356 64982 12380
rect 64962 11818 64968 12356
rect 64962 11804 64982 11818
rect 64192 11754 64680 11760
rect 64192 11720 64204 11754
rect 64668 11720 64680 11754
rect 64192 11714 64680 11720
rect 64394 11652 64454 11714
rect 64192 11646 64680 11652
rect 64192 11612 64204 11646
rect 64668 11612 64680 11646
rect 64192 11606 64680 11612
rect 63900 11532 63910 11562
rect 62926 11006 62932 11528
rect 63904 11010 63910 11532
rect 62926 10986 62944 11006
rect 62156 10936 62644 10942
rect 62156 10902 62168 10936
rect 62632 10902 62644 10936
rect 62156 10896 62644 10902
rect 62360 10834 62420 10896
rect 62156 10828 62644 10834
rect 62156 10794 62168 10828
rect 62632 10794 62644 10828
rect 62156 10788 62644 10794
rect 61864 10716 61874 10744
rect 60890 10186 60896 10716
rect 61868 10186 61874 10716
rect 60890 10168 60902 10186
rect 60120 10118 60608 10124
rect 60120 10084 60132 10118
rect 60596 10084 60608 10118
rect 60120 10078 60608 10084
rect 60324 10016 60384 10078
rect 60120 10010 60608 10016
rect 60120 9976 60132 10010
rect 60596 9976 60608 10010
rect 60120 9970 60608 9976
rect 59830 9904 59838 9926
rect 58854 9374 58860 9896
rect 59832 9382 59838 9904
rect 58854 9350 58870 9374
rect 58084 9300 58572 9306
rect 58084 9266 58096 9300
rect 58560 9266 58572 9300
rect 58084 9260 58572 9266
rect 58294 9198 58354 9260
rect 58084 9192 58572 9198
rect 58084 9158 58096 9192
rect 58560 9158 58572 9192
rect 58084 9152 58572 9158
rect 57792 9088 57802 9108
rect 56818 8558 56824 9086
rect 57796 8560 57802 9088
rect 56818 8532 56832 8558
rect 56048 8482 56536 8488
rect 56048 8448 56060 8482
rect 56524 8448 56536 8482
rect 56048 8442 56536 8448
rect 56262 8380 56322 8442
rect 56048 8374 56536 8380
rect 56048 8340 56060 8374
rect 56524 8340 56536 8374
rect 56048 8334 56536 8340
rect 55752 8264 55766 8290
rect 55760 7714 55766 8264
rect 55800 8264 55812 8290
rect 56772 8290 56832 8532
rect 57792 8532 57802 8560
rect 57836 9088 57852 9108
rect 58810 9108 58870 9350
rect 59830 9350 59838 9382
rect 59872 9904 59890 9926
rect 60842 9926 60902 10168
rect 61864 10168 61874 10186
rect 61908 10716 61924 10744
rect 62884 10744 62944 10986
rect 63900 10986 63910 11010
rect 63944 11532 63960 11562
rect 64922 11562 64982 11804
rect 66800 11638 66860 14032
rect 67060 12758 67120 15132
rect 67060 12752 67122 12758
rect 67060 12692 67062 12752
rect 67060 12686 67122 12692
rect 66920 12480 66926 12540
rect 66986 12480 66992 12540
rect 66794 11578 66800 11638
rect 66860 11578 66866 11638
rect 63944 11010 63950 11532
rect 63944 10986 63960 11010
rect 63174 10936 63662 10942
rect 63174 10902 63186 10936
rect 63650 10902 63662 10936
rect 63174 10896 63662 10902
rect 63372 10834 63432 10896
rect 63174 10828 63662 10834
rect 63174 10794 63186 10828
rect 63650 10794 63662 10828
rect 63174 10788 63662 10794
rect 62884 10716 62892 10744
rect 61908 10186 61914 10716
rect 62886 10186 62892 10716
rect 61908 10168 61924 10186
rect 61138 10118 61626 10124
rect 61138 10084 61150 10118
rect 61614 10084 61626 10118
rect 61138 10078 61626 10084
rect 61340 10016 61400 10078
rect 61138 10010 61626 10016
rect 61138 9976 61150 10010
rect 61614 9976 61626 10010
rect 61138 9970 61626 9976
rect 59872 9382 59878 9904
rect 60842 9896 60856 9926
rect 59872 9350 59890 9382
rect 60850 9374 60856 9896
rect 59102 9300 59590 9306
rect 59102 9266 59114 9300
rect 59578 9266 59590 9300
rect 59102 9260 59590 9266
rect 59296 9198 59356 9260
rect 59102 9192 59590 9198
rect 59102 9158 59114 9192
rect 59578 9158 59590 9192
rect 59102 9152 59590 9158
rect 57836 8560 57842 9088
rect 58810 9084 58820 9108
rect 57836 8532 57852 8560
rect 58814 8556 58820 9084
rect 57066 8482 57554 8488
rect 57066 8448 57078 8482
rect 57542 8448 57554 8482
rect 57066 8442 57554 8448
rect 57276 8380 57336 8442
rect 57066 8374 57554 8380
rect 57066 8340 57078 8374
rect 57542 8340 57554 8374
rect 57066 8334 57554 8340
rect 56772 8268 56784 8290
rect 55800 7714 55806 8264
rect 55760 7702 55806 7714
rect 56778 7714 56784 8268
rect 56818 8268 56832 8290
rect 57792 8290 57852 8532
rect 58810 8532 58820 8556
rect 58854 9084 58870 9108
rect 59830 9108 59890 9350
rect 60842 9350 60856 9374
rect 60890 9896 60902 9926
rect 61864 9926 61924 10168
rect 62884 10168 62892 10186
rect 62926 10716 62944 10744
rect 63900 10744 63960 10986
rect 64922 10986 64928 11562
rect 64962 11528 64982 11562
rect 64962 11006 64968 11528
rect 64962 10986 64982 11006
rect 64192 10936 64680 10942
rect 64192 10902 64204 10936
rect 64668 10902 64680 10936
rect 64192 10896 64680 10902
rect 64392 10834 64452 10896
rect 64192 10828 64680 10834
rect 64192 10794 64204 10828
rect 64668 10794 64680 10828
rect 64192 10788 64680 10794
rect 63900 10720 63910 10744
rect 62926 10186 62932 10716
rect 63904 10190 63910 10720
rect 62926 10168 62944 10186
rect 62156 10118 62644 10124
rect 62156 10084 62168 10118
rect 62632 10084 62644 10118
rect 62156 10078 62644 10084
rect 62362 10016 62422 10078
rect 62156 10010 62644 10016
rect 62156 9976 62168 10010
rect 62632 9976 62644 10010
rect 62156 9970 62644 9976
rect 61864 9896 61874 9926
rect 60890 9374 60896 9896
rect 61868 9374 61874 9896
rect 60890 9350 60902 9374
rect 60120 9300 60608 9306
rect 60120 9266 60132 9300
rect 60596 9266 60608 9300
rect 60120 9260 60608 9266
rect 60326 9198 60386 9260
rect 60120 9192 60608 9198
rect 60120 9158 60132 9192
rect 60596 9158 60608 9192
rect 60120 9152 60608 9158
rect 59830 9092 59838 9108
rect 58854 8556 58860 9084
rect 59832 8564 59838 9092
rect 58854 8532 58870 8556
rect 58084 8482 58572 8488
rect 58084 8448 58096 8482
rect 58560 8448 58572 8482
rect 58084 8442 58572 8448
rect 58296 8380 58356 8442
rect 58084 8374 58572 8380
rect 58084 8340 58096 8374
rect 58560 8340 58572 8374
rect 58084 8334 58572 8340
rect 57792 8270 57802 8290
rect 56818 7714 56824 8268
rect 57796 7760 57802 8270
rect 56778 7702 56824 7714
rect 57786 7714 57802 7760
rect 57836 8270 57852 8290
rect 58810 8290 58870 8532
rect 59830 8532 59838 8564
rect 59872 9092 59890 9108
rect 60842 9108 60902 9350
rect 61864 9350 61874 9374
rect 61908 9896 61924 9926
rect 62884 9926 62944 10168
rect 63900 10168 63910 10190
rect 63944 10720 63960 10744
rect 64922 10744 64982 10986
rect 63944 10190 63950 10720
rect 63944 10168 63960 10190
rect 63174 10118 63662 10124
rect 63174 10084 63186 10118
rect 63650 10084 63662 10118
rect 63174 10078 63662 10084
rect 63374 10016 63434 10078
rect 63174 10010 63662 10016
rect 63174 9976 63186 10010
rect 63650 9976 63662 10010
rect 63174 9970 63662 9976
rect 62884 9896 62892 9926
rect 61908 9374 61914 9896
rect 62886 9374 62892 9896
rect 61908 9350 61924 9374
rect 61138 9300 61626 9306
rect 61138 9266 61150 9300
rect 61614 9266 61626 9300
rect 61138 9260 61626 9266
rect 61342 9198 61402 9260
rect 61138 9192 61626 9198
rect 61138 9158 61150 9192
rect 61614 9158 61626 9192
rect 61138 9152 61626 9158
rect 59872 8564 59878 9092
rect 60842 9084 60856 9108
rect 59872 8532 59890 8564
rect 60850 8556 60856 9084
rect 59102 8482 59590 8488
rect 59102 8448 59114 8482
rect 59578 8448 59590 8482
rect 59102 8442 59590 8448
rect 59298 8380 59358 8442
rect 59102 8374 59590 8380
rect 59102 8340 59114 8374
rect 59578 8340 59590 8374
rect 59102 8334 59590 8340
rect 57836 7760 57842 8270
rect 58810 8266 58820 8290
rect 57836 7714 57846 7760
rect 56048 7664 56536 7670
rect 56048 7630 56060 7664
rect 56524 7630 56536 7664
rect 56048 7624 56536 7630
rect 57066 7664 57554 7670
rect 57066 7630 57078 7664
rect 57542 7630 57554 7664
rect 57066 7624 57554 7630
rect 57786 7540 57846 7714
rect 58814 7714 58820 8266
rect 58854 8266 58870 8290
rect 59830 8290 59890 8532
rect 60842 8532 60856 8556
rect 60890 9084 60902 9108
rect 61864 9108 61924 9350
rect 62884 9350 62892 9374
rect 62926 9896 62944 9926
rect 63900 9926 63960 10168
rect 64922 10168 64928 10744
rect 64962 10716 64982 10744
rect 64962 10186 64968 10716
rect 64962 10168 64982 10186
rect 64192 10118 64680 10124
rect 64192 10084 64204 10118
rect 64668 10084 64680 10118
rect 64192 10078 64680 10084
rect 64394 10016 64454 10078
rect 64192 10010 64680 10016
rect 64192 9976 64204 10010
rect 64668 9976 64680 10010
rect 64192 9970 64680 9976
rect 63900 9900 63910 9926
rect 62926 9374 62932 9896
rect 63904 9378 63910 9900
rect 62926 9350 62944 9374
rect 62156 9300 62644 9306
rect 62156 9266 62168 9300
rect 62632 9266 62644 9300
rect 62156 9260 62644 9266
rect 62364 9198 62424 9260
rect 62156 9192 62644 9198
rect 62156 9158 62168 9192
rect 62632 9158 62644 9192
rect 62156 9152 62644 9158
rect 61864 9084 61874 9108
rect 60890 8556 60896 9084
rect 61868 8556 61874 9084
rect 60890 8532 60902 8556
rect 60120 8482 60608 8488
rect 60120 8448 60132 8482
rect 60596 8448 60608 8482
rect 60120 8442 60608 8448
rect 60328 8380 60388 8442
rect 60120 8374 60608 8380
rect 60120 8340 60132 8374
rect 60596 8340 60608 8374
rect 60120 8334 60608 8340
rect 59830 8274 59838 8290
rect 58854 7714 58860 8266
rect 59832 7762 59838 8274
rect 58814 7702 58860 7714
rect 59824 7714 59838 7762
rect 59872 8274 59890 8290
rect 60842 8290 60902 8532
rect 61864 8532 61874 8556
rect 61908 9084 61924 9108
rect 62884 9108 62944 9350
rect 63900 9350 63910 9378
rect 63944 9900 63960 9926
rect 64922 9926 64982 10168
rect 63944 9378 63950 9900
rect 63944 9350 63960 9378
rect 63174 9300 63662 9306
rect 63174 9266 63186 9300
rect 63650 9266 63662 9300
rect 63174 9260 63662 9266
rect 63376 9198 63436 9260
rect 63174 9192 63662 9198
rect 63174 9158 63186 9192
rect 63650 9158 63662 9192
rect 63174 9152 63662 9158
rect 62884 9084 62892 9108
rect 61908 8556 61914 9084
rect 62886 8556 62892 9084
rect 61908 8532 61924 8556
rect 61138 8482 61626 8488
rect 61138 8448 61150 8482
rect 61614 8448 61626 8482
rect 61138 8442 61626 8448
rect 61344 8380 61404 8442
rect 61138 8374 61626 8380
rect 61138 8340 61150 8374
rect 61614 8340 61626 8374
rect 61138 8334 61626 8340
rect 59872 7762 59878 8274
rect 60842 8266 60856 8290
rect 59872 7714 59884 7762
rect 58084 7664 58572 7670
rect 58084 7630 58096 7664
rect 58560 7630 58572 7664
rect 58084 7624 58572 7630
rect 59102 7664 59590 7670
rect 59102 7630 59114 7664
rect 59578 7630 59590 7664
rect 59102 7624 59590 7630
rect 59824 7540 59884 7714
rect 60850 7714 60856 8266
rect 60890 8266 60902 8290
rect 61864 8290 61924 8532
rect 62884 8532 62892 8556
rect 62926 9084 62944 9108
rect 63900 9108 63960 9350
rect 64922 9350 64928 9926
rect 64962 9896 64982 9926
rect 64962 9374 64968 9896
rect 64962 9350 64982 9374
rect 64192 9300 64680 9306
rect 64192 9266 64204 9300
rect 64668 9266 64680 9300
rect 64192 9260 64680 9266
rect 64396 9198 64456 9260
rect 64192 9192 64680 9198
rect 64192 9158 64204 9192
rect 64668 9158 64680 9192
rect 64192 9152 64680 9158
rect 63900 9088 63910 9108
rect 62926 8556 62932 9084
rect 63904 8560 63910 9088
rect 62926 8532 62944 8556
rect 62156 8482 62644 8488
rect 62156 8448 62168 8482
rect 62632 8448 62644 8482
rect 62156 8442 62644 8448
rect 62366 8380 62426 8442
rect 62156 8374 62644 8380
rect 62156 8340 62168 8374
rect 62632 8340 62644 8374
rect 62156 8334 62644 8340
rect 61864 8266 61874 8290
rect 60890 7714 60896 8266
rect 61868 7758 61874 8266
rect 60850 7702 60896 7714
rect 61860 7714 61874 7758
rect 61908 8266 61924 8290
rect 62884 8290 62944 8532
rect 63900 8532 63910 8560
rect 63944 9088 63960 9108
rect 64922 9108 64982 9350
rect 63944 8560 63950 9088
rect 63944 8532 63960 8560
rect 63174 8482 63662 8488
rect 63174 8448 63186 8482
rect 63650 8448 63662 8482
rect 63174 8442 63662 8448
rect 63378 8380 63438 8442
rect 63174 8374 63662 8380
rect 63174 8340 63186 8374
rect 63650 8340 63662 8374
rect 63174 8334 63662 8340
rect 62884 8266 62892 8290
rect 61908 7758 61914 8266
rect 61908 7714 61920 7758
rect 60120 7664 60608 7670
rect 60120 7630 60132 7664
rect 60596 7630 60608 7664
rect 60120 7624 60608 7630
rect 61138 7664 61626 7670
rect 61138 7630 61150 7664
rect 61614 7630 61626 7664
rect 61138 7624 61626 7630
rect 61860 7540 61920 7714
rect 62886 7714 62892 8266
rect 62926 8266 62944 8290
rect 63900 8290 63960 8532
rect 64922 8532 64928 9108
rect 64962 9084 64982 9108
rect 64962 8556 64968 9084
rect 64962 8532 64982 8556
rect 64192 8482 64680 8488
rect 64192 8448 64204 8482
rect 64668 8448 64680 8482
rect 64192 8442 64680 8448
rect 64398 8380 64458 8442
rect 64192 8374 64680 8380
rect 64192 8340 64204 8374
rect 64668 8340 64680 8374
rect 64192 8334 64680 8340
rect 63900 8270 63910 8290
rect 62926 7714 62932 8266
rect 63904 7756 63910 8270
rect 62886 7702 62932 7714
rect 63896 7714 63910 7756
rect 63944 8270 63960 8290
rect 64922 8290 64982 8532
rect 63944 7756 63950 8270
rect 64922 7768 64928 8290
rect 63944 7714 63956 7756
rect 62156 7664 62644 7670
rect 62156 7630 62168 7664
rect 62632 7630 62644 7664
rect 62156 7624 62644 7630
rect 63174 7664 63662 7670
rect 63174 7630 63186 7664
rect 63650 7630 63662 7664
rect 63174 7624 63662 7630
rect 63896 7540 63956 7714
rect 64916 7714 64928 7768
rect 64962 8266 64982 8290
rect 64962 7768 64968 8266
rect 64962 7714 64976 7768
rect 64192 7664 64680 7670
rect 64192 7630 64204 7664
rect 64668 7630 64680 7664
rect 64192 7624 64680 7630
rect 64410 7540 64470 7624
rect 64916 7540 64976 7714
rect 65902 7682 65962 7688
rect 57786 7480 64976 7540
rect 65640 7652 65700 7674
rect 61968 6320 61974 6380
rect 62034 6320 62040 6380
rect 55534 4926 56612 4986
rect 55534 4747 55594 4926
rect 56048 4837 56108 4926
rect 55827 4831 56315 4837
rect 55827 4797 55839 4831
rect 56303 4797 56315 4831
rect 55827 4791 56315 4797
rect 55534 4702 55545 4747
rect 55539 4171 55545 4702
rect 55579 4702 55594 4747
rect 56552 4747 56612 4926
rect 57558 4880 57564 4940
rect 57624 4880 57630 4940
rect 57932 4926 59154 4986
rect 61974 4984 62034 6320
rect 56845 4831 57333 4837
rect 56845 4797 56857 4831
rect 57321 4797 57333 4831
rect 56845 4791 57333 4797
rect 55579 4171 55585 4702
rect 56552 4698 56563 4747
rect 56557 4216 56563 4698
rect 55539 4159 55585 4171
rect 56550 4171 56563 4216
rect 56597 4698 56612 4747
rect 57564 4747 57624 4880
rect 58072 4837 58132 4926
rect 57863 4831 58351 4837
rect 57863 4797 57875 4831
rect 58339 4797 58351 4831
rect 57863 4791 58351 4797
rect 56597 4216 56603 4698
rect 56597 4171 56610 4216
rect 55827 4121 56315 4127
rect 55827 4087 55839 4121
rect 56303 4087 56315 4121
rect 55827 4081 56315 4087
rect 56550 4036 56610 4171
rect 57564 4171 57581 4747
rect 57615 4171 57624 4747
rect 58588 4747 58648 4926
rect 59094 4837 59154 4926
rect 59598 4880 59604 4940
rect 59664 4880 59670 4940
rect 60624 4924 62034 4984
rect 58881 4831 59369 4837
rect 58881 4797 58893 4831
rect 59357 4797 59369 4831
rect 58881 4791 59369 4797
rect 58588 4690 58599 4747
rect 58593 4212 58599 4690
rect 56845 4121 57333 4127
rect 56845 4087 56857 4121
rect 57321 4087 57333 4121
rect 56845 4081 57333 4087
rect 55406 3976 55412 4036
rect 55472 3976 55478 4036
rect 56544 3976 56550 4036
rect 56610 3976 56616 4036
rect 55412 1614 55472 3976
rect 55532 3760 56608 3820
rect 55532 3634 55592 3760
rect 56042 3724 56102 3760
rect 55826 3718 56314 3724
rect 55826 3684 55838 3718
rect 56302 3684 56314 3718
rect 55826 3678 56314 3684
rect 55532 3574 55544 3634
rect 55538 3058 55544 3574
rect 55578 3574 55592 3634
rect 56548 3634 56608 3760
rect 57060 3724 57120 4081
rect 57564 3940 57624 4171
rect 58586 4171 58599 4212
rect 58633 4690 58648 4747
rect 59604 4747 59664 4880
rect 59899 4831 60387 4837
rect 59899 4797 59911 4831
rect 60375 4797 60387 4831
rect 59899 4791 60387 4797
rect 59604 4702 59617 4747
rect 58633 4212 58639 4690
rect 58633 4171 58646 4212
rect 59611 4210 59617 4702
rect 57863 4121 58351 4127
rect 57863 4087 57875 4121
rect 58339 4087 58351 4121
rect 57863 4081 58351 4087
rect 57558 3880 57564 3940
rect 57624 3880 57630 3940
rect 56844 3718 57332 3724
rect 56844 3684 56856 3718
rect 57320 3684 57332 3718
rect 56844 3678 57332 3684
rect 56548 3588 56562 3634
rect 55578 3058 55584 3574
rect 56556 3104 56562 3588
rect 55538 3046 55584 3058
rect 56548 3058 56562 3104
rect 56596 3588 56608 3634
rect 57564 3634 57624 3880
rect 58080 3724 58140 4081
rect 58586 3824 58646 4171
rect 59604 4171 59617 4210
rect 59651 4702 59664 4747
rect 60624 4747 60684 4924
rect 61132 4837 61192 4924
rect 60917 4831 61405 4837
rect 60917 4797 60929 4831
rect 61393 4797 61405 4831
rect 60917 4791 61405 4797
rect 59651 4210 59657 4702
rect 60624 4694 60635 4747
rect 60629 4216 60635 4694
rect 59651 4171 59664 4210
rect 58881 4121 59369 4127
rect 58881 4087 58893 4121
rect 59357 4087 59369 4121
rect 58881 4081 59369 4087
rect 58580 3764 58586 3824
rect 58646 3764 58652 3824
rect 59088 3724 59148 4081
rect 59604 3940 59664 4171
rect 60624 4171 60635 4216
rect 60669 4694 60684 4747
rect 61640 4747 61700 4924
rect 61640 4700 61653 4747
rect 60669 4216 60675 4694
rect 60669 4171 60684 4216
rect 59899 4121 60387 4127
rect 59899 4087 59911 4121
rect 60375 4087 60387 4121
rect 59899 4081 60387 4087
rect 59598 3880 59604 3940
rect 59664 3880 59670 3940
rect 57862 3718 58350 3724
rect 57862 3684 57874 3718
rect 58338 3684 58350 3718
rect 57862 3678 58350 3684
rect 58880 3718 59368 3724
rect 58880 3684 58892 3718
rect 59356 3684 59368 3718
rect 58880 3678 59368 3684
rect 57564 3588 57580 3634
rect 56596 3104 56602 3588
rect 56596 3058 56608 3104
rect 57574 3100 57580 3588
rect 55826 3008 56314 3014
rect 55826 2974 55838 3008
rect 56302 2974 56314 3008
rect 55826 2968 56314 2974
rect 56548 2816 56608 3058
rect 57566 3058 57580 3100
rect 57614 3588 57624 3634
rect 58592 3634 58638 3646
rect 57614 3100 57620 3588
rect 58592 3110 58598 3634
rect 57614 3058 57626 3100
rect 56844 3008 57332 3014
rect 56844 2974 56856 3008
rect 57320 2974 57332 3008
rect 56844 2968 57332 2974
rect 56690 2864 56696 2924
rect 56756 2864 56762 2924
rect 56542 2756 56548 2816
rect 56608 2756 56614 2816
rect 56696 2714 56756 2864
rect 55532 2654 56756 2714
rect 55532 2523 55592 2654
rect 56048 2613 56108 2654
rect 55827 2607 56315 2613
rect 55827 2573 55839 2607
rect 56303 2573 56315 2607
rect 55827 2567 56315 2573
rect 55532 2482 55545 2523
rect 55539 1947 55545 2482
rect 55579 2482 55592 2523
rect 56550 2523 56610 2654
rect 57066 2613 57126 2968
rect 57566 2704 57626 3058
rect 58582 3058 58598 3110
rect 58632 3110 58638 3634
rect 59604 3634 59664 3880
rect 60110 3724 60170 4081
rect 60624 4036 60684 4171
rect 61647 4171 61653 4700
rect 61687 4700 61700 4747
rect 61687 4171 61693 4700
rect 61647 4159 61693 4171
rect 60917 4121 61405 4127
rect 60917 4087 60929 4121
rect 61393 4087 61405 4121
rect 60917 4081 61405 4087
rect 60618 3976 60624 4036
rect 60684 3976 60690 4036
rect 62104 3930 62164 7480
rect 64130 7356 64136 7416
rect 64196 7356 64202 7416
rect 65042 7356 65048 7416
rect 65108 7356 65114 7416
rect 63260 7246 63266 7306
rect 63326 7246 63332 7306
rect 62346 7138 62352 7198
rect 62412 7138 62418 7198
rect 62352 5644 62412 7138
rect 62476 7030 62482 7090
rect 62542 7030 62548 7090
rect 62482 5766 62542 7030
rect 62708 6990 62796 6996
rect 62708 6956 62720 6990
rect 62784 6956 62796 6990
rect 62708 6950 62796 6956
rect 62926 6990 63014 6996
rect 62926 6956 62938 6990
rect 63002 6956 63014 6990
rect 62926 6950 63014 6956
rect 63144 6990 63232 6996
rect 63144 6956 63156 6990
rect 63220 6956 63232 6990
rect 63144 6950 63232 6956
rect 62620 6906 62666 6918
rect 62620 6760 62626 6906
rect 62612 6730 62626 6760
rect 62660 6760 62666 6906
rect 62838 6906 62884 6918
rect 62660 6730 62672 6760
rect 62838 6752 62844 6906
rect 62612 6580 62672 6730
rect 62832 6730 62844 6752
rect 62878 6752 62884 6906
rect 63056 6906 63102 6918
rect 62878 6730 62892 6752
rect 63056 6742 63062 6906
rect 62708 6680 62796 6686
rect 62708 6646 62720 6680
rect 62784 6646 62796 6680
rect 62708 6640 62796 6646
rect 62720 6580 62780 6640
rect 62832 6580 62892 6730
rect 63048 6730 63062 6742
rect 63096 6742 63102 6906
rect 63266 6906 63326 7246
rect 64024 7138 64030 7198
rect 64090 7138 64096 7198
rect 63806 7030 63812 7090
rect 63872 7030 63878 7090
rect 63812 6996 63872 7030
rect 64030 6996 64090 7138
rect 63362 6990 63450 6996
rect 63362 6956 63374 6990
rect 63438 6956 63450 6990
rect 63362 6950 63450 6956
rect 63580 6990 63668 6996
rect 63580 6956 63592 6990
rect 63656 6956 63668 6990
rect 63580 6950 63668 6956
rect 63798 6990 63886 6996
rect 63798 6956 63810 6990
rect 63874 6956 63886 6990
rect 63798 6950 63886 6956
rect 64016 6990 64104 6996
rect 64016 6956 64028 6990
rect 64092 6956 64104 6990
rect 64016 6950 64104 6956
rect 63266 6890 63280 6906
rect 63096 6730 63108 6742
rect 62926 6680 63014 6686
rect 62926 6646 62938 6680
rect 63002 6646 63014 6680
rect 62926 6640 63014 6646
rect 62940 6590 63000 6640
rect 62612 6520 62892 6580
rect 62934 6530 62940 6590
rect 63000 6530 63006 6590
rect 62832 6262 62892 6520
rect 63048 6490 63108 6730
rect 63274 6730 63280 6890
rect 63314 6890 63326 6906
rect 63492 6906 63538 6918
rect 63314 6730 63320 6890
rect 63492 6756 63498 6906
rect 63274 6718 63320 6730
rect 63486 6730 63498 6756
rect 63532 6756 63538 6906
rect 63710 6906 63756 6918
rect 63710 6766 63716 6906
rect 63532 6730 63546 6756
rect 63144 6680 63232 6686
rect 63144 6646 63156 6680
rect 63220 6646 63232 6680
rect 63144 6640 63232 6646
rect 63362 6680 63450 6686
rect 63362 6646 63374 6680
rect 63438 6646 63450 6680
rect 63362 6640 63450 6646
rect 63042 6430 63048 6490
rect 63108 6430 63114 6490
rect 63044 6320 63050 6380
rect 63110 6320 63116 6380
rect 62614 6202 62892 6262
rect 62614 6074 62674 6202
rect 62724 6164 62784 6202
rect 62708 6158 62796 6164
rect 62708 6124 62720 6158
rect 62784 6124 62796 6158
rect 62708 6118 62796 6124
rect 62614 6048 62626 6074
rect 62620 5898 62626 6048
rect 62660 6048 62674 6074
rect 62832 6074 62892 6202
rect 62926 6158 63014 6164
rect 62926 6124 62938 6158
rect 63002 6124 63014 6158
rect 62926 6118 63014 6124
rect 62660 5898 62666 6048
rect 62620 5886 62666 5898
rect 62832 5898 62844 6074
rect 62878 5898 62892 6074
rect 63050 6074 63110 6320
rect 63158 6270 63218 6640
rect 63378 6270 63438 6640
rect 63486 6490 63546 6730
rect 63702 6730 63716 6766
rect 63750 6766 63756 6906
rect 63928 6906 63974 6918
rect 63750 6730 63762 6766
rect 63928 6764 63934 6906
rect 63580 6680 63668 6686
rect 63580 6646 63592 6680
rect 63656 6646 63668 6680
rect 63580 6640 63668 6646
rect 63596 6590 63656 6640
rect 63590 6530 63596 6590
rect 63656 6530 63662 6590
rect 63480 6430 63486 6490
rect 63546 6430 63552 6490
rect 63478 6320 63484 6380
rect 63544 6320 63550 6380
rect 63152 6210 63158 6270
rect 63218 6210 63224 6270
rect 63372 6210 63378 6270
rect 63438 6210 63444 6270
rect 63158 6164 63218 6210
rect 63378 6164 63438 6210
rect 63144 6158 63232 6164
rect 63144 6124 63156 6158
rect 63220 6124 63232 6158
rect 63144 6118 63232 6124
rect 63362 6158 63450 6164
rect 63362 6124 63374 6158
rect 63438 6124 63450 6158
rect 63362 6118 63450 6124
rect 63050 6038 63062 6074
rect 62708 5848 62796 5854
rect 62708 5814 62720 5848
rect 62784 5814 62796 5848
rect 62708 5808 62796 5814
rect 62476 5706 62482 5766
rect 62542 5706 62548 5766
rect 62346 5584 62352 5644
rect 62412 5584 62418 5644
rect 62832 5520 62892 5898
rect 63056 5898 63062 6038
rect 63096 6038 63110 6074
rect 63274 6074 63320 6086
rect 63096 5898 63102 6038
rect 63274 5938 63280 6074
rect 63056 5886 63102 5898
rect 63270 5898 63280 5938
rect 63314 5938 63320 6074
rect 63484 6074 63544 6320
rect 63580 6158 63668 6164
rect 63580 6124 63592 6158
rect 63656 6124 63668 6158
rect 63580 6118 63668 6124
rect 63484 6044 63498 6074
rect 63314 5898 63330 5938
rect 62926 5848 63014 5854
rect 62926 5814 62938 5848
rect 63002 5814 63014 5848
rect 62926 5808 63014 5814
rect 63144 5848 63232 5854
rect 63144 5814 63156 5848
rect 63220 5814 63232 5848
rect 63144 5808 63232 5814
rect 62940 5766 63000 5808
rect 62934 5706 62940 5766
rect 63000 5706 63006 5766
rect 63158 5644 63218 5808
rect 63152 5584 63158 5644
rect 63218 5584 63224 5644
rect 62826 5460 62832 5520
rect 62892 5460 62898 5520
rect 63270 5394 63330 5898
rect 63492 5898 63498 6044
rect 63532 6044 63544 6074
rect 63702 6074 63762 6730
rect 63922 6730 63934 6764
rect 63968 6764 63974 6906
rect 64136 6906 64196 7356
rect 64922 7246 64928 7306
rect 64988 7246 64994 7306
rect 64242 7138 64248 7198
rect 64308 7138 64314 7198
rect 64248 6996 64308 7138
rect 64460 7030 64466 7090
rect 64526 7030 64532 7090
rect 64466 6996 64526 7030
rect 64234 6990 64322 6996
rect 64234 6956 64246 6990
rect 64310 6956 64322 6990
rect 64234 6950 64322 6956
rect 64452 6990 64540 6996
rect 64452 6956 64464 6990
rect 64528 6956 64540 6990
rect 64452 6950 64540 6956
rect 64670 6990 64758 6996
rect 64670 6956 64682 6990
rect 64746 6956 64758 6990
rect 64670 6950 64758 6956
rect 64136 6860 64152 6906
rect 63968 6730 63982 6764
rect 63798 6680 63886 6686
rect 63798 6646 63810 6680
rect 63874 6646 63886 6680
rect 63798 6640 63886 6646
rect 63922 6490 63982 6730
rect 64146 6730 64152 6860
rect 64186 6860 64196 6906
rect 64364 6906 64410 6918
rect 64186 6730 64192 6860
rect 64364 6756 64370 6906
rect 64146 6718 64192 6730
rect 64358 6730 64370 6756
rect 64404 6756 64410 6906
rect 64582 6906 64628 6918
rect 64404 6730 64418 6756
rect 64582 6748 64588 6906
rect 64016 6680 64104 6686
rect 64016 6646 64028 6680
rect 64092 6646 64104 6680
rect 64016 6640 64104 6646
rect 64234 6680 64322 6686
rect 64234 6646 64246 6680
rect 64310 6646 64322 6680
rect 64234 6640 64322 6646
rect 64358 6490 64418 6730
rect 64576 6730 64588 6748
rect 64622 6748 64628 6906
rect 64800 6906 64846 6918
rect 64800 6766 64806 6906
rect 64622 6730 64636 6748
rect 64452 6680 64540 6686
rect 64452 6646 64464 6680
rect 64528 6646 64540 6680
rect 64452 6640 64540 6646
rect 64460 6530 64466 6590
rect 64526 6530 64532 6590
rect 64576 6588 64636 6730
rect 64794 6730 64806 6766
rect 64840 6766 64846 6906
rect 64928 6816 64988 7246
rect 64840 6730 64854 6766
rect 64670 6680 64758 6686
rect 64670 6646 64682 6680
rect 64746 6646 64758 6680
rect 64670 6640 64758 6646
rect 64684 6588 64744 6640
rect 64794 6588 64854 6730
rect 63812 6430 64418 6490
rect 63812 6380 63872 6430
rect 63806 6320 63812 6380
rect 63872 6320 63878 6380
rect 63916 6320 63922 6380
rect 63982 6320 63988 6380
rect 64352 6320 64358 6380
rect 64418 6320 64424 6380
rect 63798 6158 63886 6164
rect 63798 6124 63810 6158
rect 63874 6124 63886 6158
rect 63798 6118 63886 6124
rect 63532 5898 63538 6044
rect 63492 5886 63538 5898
rect 63702 5898 63716 6074
rect 63750 5898 63762 6074
rect 63922 6074 63982 6320
rect 64026 6210 64032 6270
rect 64092 6210 64098 6270
rect 64242 6210 64248 6270
rect 64308 6210 64314 6270
rect 64032 6164 64092 6210
rect 64248 6164 64308 6210
rect 64016 6158 64104 6164
rect 64016 6124 64028 6158
rect 64092 6124 64104 6158
rect 64016 6118 64104 6124
rect 64234 6158 64322 6164
rect 64234 6124 64246 6158
rect 64310 6124 64322 6158
rect 64234 6118 64322 6124
rect 63922 6056 63934 6074
rect 63362 5848 63450 5854
rect 63362 5814 63374 5848
rect 63438 5814 63450 5848
rect 63362 5808 63450 5814
rect 63580 5848 63668 5854
rect 63580 5814 63592 5848
rect 63656 5814 63668 5848
rect 63580 5808 63668 5814
rect 63376 5644 63436 5808
rect 63596 5766 63656 5808
rect 63590 5706 63596 5766
rect 63656 5706 63662 5766
rect 63370 5584 63376 5644
rect 63436 5584 63442 5644
rect 63264 5334 63270 5394
rect 63330 5334 63336 5394
rect 63606 5280 63654 5706
rect 63702 5520 63762 5898
rect 63928 5898 63934 6056
rect 63968 6056 63982 6074
rect 64146 6074 64192 6086
rect 63968 5898 63974 6056
rect 64146 5920 64152 6074
rect 63928 5886 63974 5898
rect 64140 5898 64152 5920
rect 64186 5920 64192 6074
rect 64358 6074 64418 6320
rect 64466 6164 64526 6530
rect 64576 6528 64854 6588
rect 64576 6470 64636 6528
rect 64570 6410 64576 6470
rect 64636 6410 64642 6470
rect 64576 6272 64636 6410
rect 64576 6212 64854 6272
rect 64452 6158 64540 6164
rect 64452 6124 64464 6158
rect 64528 6124 64540 6158
rect 64452 6118 64540 6124
rect 64358 6042 64370 6074
rect 64186 5898 64200 5920
rect 63798 5848 63886 5854
rect 63798 5814 63810 5848
rect 63874 5814 63886 5848
rect 63798 5808 63886 5814
rect 64016 5848 64104 5854
rect 64016 5814 64028 5848
rect 64092 5814 64104 5848
rect 64016 5808 64104 5814
rect 63812 5646 63872 5808
rect 64140 5766 64200 5898
rect 64364 5898 64370 6042
rect 64404 6042 64418 6074
rect 64576 6074 64636 6212
rect 64684 6164 64744 6212
rect 64670 6158 64758 6164
rect 64670 6124 64682 6158
rect 64746 6124 64758 6158
rect 64670 6118 64758 6124
rect 64576 6056 64588 6074
rect 64404 5898 64410 6042
rect 64582 5928 64588 6056
rect 64364 5886 64410 5898
rect 64574 5898 64588 5928
rect 64622 6056 64636 6074
rect 64794 6074 64854 6212
rect 64622 5928 64628 6056
rect 64794 6054 64806 6074
rect 64622 5898 64634 5928
rect 64234 5848 64322 5854
rect 64234 5814 64246 5848
rect 64310 5814 64322 5848
rect 64234 5808 64322 5814
rect 64452 5848 64540 5854
rect 64452 5814 64464 5848
rect 64528 5814 64540 5848
rect 64452 5808 64540 5814
rect 64134 5706 64140 5766
rect 64200 5706 64206 5766
rect 64468 5646 64528 5808
rect 63806 5586 63812 5646
rect 63872 5586 63878 5646
rect 64462 5586 64468 5646
rect 64528 5586 64534 5646
rect 64574 5520 64634 5898
rect 64800 5898 64806 6054
rect 64840 6054 64854 6074
rect 64840 5898 64846 6054
rect 64800 5886 64846 5898
rect 64670 5848 64758 5854
rect 64670 5814 64682 5848
rect 64746 5814 64758 5848
rect 64670 5808 64758 5814
rect 64928 5766 64988 6756
rect 64922 5706 64928 5766
rect 64988 5706 64994 5766
rect 63696 5460 63702 5520
rect 63762 5460 63768 5520
rect 64568 5460 64574 5520
rect 64634 5460 64640 5520
rect 65048 5394 65108 7356
rect 65164 6530 65170 6590
rect 65230 6530 65236 6590
rect 65170 6344 65230 6530
rect 65170 6276 65230 6284
rect 65042 5334 65048 5394
rect 65108 5334 65114 5394
rect 63598 5228 63604 5280
rect 63656 5228 63662 5280
rect 65640 5200 65700 7592
rect 62412 5140 65700 5200
rect 62274 4900 62280 4960
rect 62340 4900 62346 4960
rect 60622 3870 62164 3930
rect 59898 3718 60386 3724
rect 59898 3684 59910 3718
rect 60374 3684 60386 3718
rect 59898 3678 60386 3684
rect 59604 3600 59616 3634
rect 58632 3058 58642 3110
rect 59610 3092 59616 3600
rect 57862 3008 58350 3014
rect 57862 2974 57874 3008
rect 58338 2974 58350 3008
rect 57862 2968 58350 2974
rect 57560 2644 57566 2704
rect 57626 2644 57632 2704
rect 56845 2607 57333 2613
rect 56845 2573 56857 2607
rect 57321 2573 57333 2607
rect 56845 2567 57333 2573
rect 56550 2482 56563 2523
rect 55579 1947 55585 2482
rect 55539 1935 55585 1947
rect 56557 1947 56563 2482
rect 56597 2482 56610 2523
rect 57566 2523 57626 2644
rect 58080 2613 58140 2968
rect 58582 2924 58642 3058
rect 59606 3058 59616 3092
rect 59650 3600 59664 3634
rect 60622 3634 60682 3870
rect 61132 3724 61192 3870
rect 60916 3718 61404 3724
rect 60916 3684 60928 3718
rect 61392 3684 61404 3718
rect 60916 3678 61404 3684
rect 61638 3634 61698 3870
rect 61742 3764 61748 3824
rect 61808 3764 61814 3824
rect 59650 3092 59656 3600
rect 60622 3588 60634 3634
rect 60624 3586 60634 3588
rect 60628 3096 60634 3586
rect 59650 3058 59666 3092
rect 58880 3008 59368 3014
rect 58880 2974 58892 3008
rect 59356 2974 59368 3008
rect 58880 2968 59368 2974
rect 58576 2864 58582 2924
rect 58642 2864 58648 2924
rect 58578 2756 58584 2816
rect 58644 2756 58650 2816
rect 57863 2607 58351 2613
rect 57863 2573 57875 2607
rect 58339 2573 58351 2607
rect 57863 2567 58351 2573
rect 57566 2494 57581 2523
rect 56597 1947 56603 2482
rect 57575 1984 57581 2494
rect 56557 1935 56603 1947
rect 57568 1947 57581 1984
rect 57615 2494 57626 2523
rect 58584 2523 58644 2756
rect 59108 2613 59168 2968
rect 59606 2710 59666 3058
rect 60620 3058 60634 3096
rect 60668 3586 60684 3634
rect 61638 3604 61652 3634
rect 61640 3602 61652 3604
rect 60668 3096 60674 3586
rect 60668 3058 60680 3096
rect 59898 3008 60386 3014
rect 59898 2974 59910 3008
rect 60374 2974 60386 3008
rect 59898 2968 60386 2974
rect 59604 2704 59666 2710
rect 59664 2644 59666 2704
rect 59604 2638 59666 2644
rect 58881 2607 59369 2613
rect 58881 2573 58893 2607
rect 59357 2573 59369 2607
rect 58881 2567 59369 2573
rect 57615 1984 57621 2494
rect 58584 2480 58599 2523
rect 57615 1947 57628 1984
rect 55827 1897 56315 1903
rect 55827 1863 55839 1897
rect 56303 1863 56315 1897
rect 55827 1857 56315 1863
rect 56845 1897 57333 1903
rect 56845 1863 56857 1897
rect 57321 1863 57333 1897
rect 56845 1857 57333 1863
rect 56544 1660 56550 1720
rect 56610 1660 56616 1720
rect 55406 1554 55412 1614
rect 55472 1554 55478 1614
rect 55826 1494 56314 1500
rect 55826 1460 55838 1494
rect 56302 1460 56314 1494
rect 55826 1454 56314 1460
rect 55538 1410 55584 1422
rect 55538 874 55544 1410
rect 55532 834 55544 874
rect 55578 874 55584 1410
rect 56550 1410 56610 1660
rect 57074 1500 57134 1857
rect 57568 1822 57628 1947
rect 58593 1947 58599 2480
rect 58633 2480 58644 2523
rect 59606 2523 59666 2638
rect 60118 2613 60178 2968
rect 60446 2864 60452 2924
rect 60512 2864 60518 2924
rect 60452 2714 60512 2864
rect 60620 2816 60680 3058
rect 61646 3058 61652 3602
rect 61686 3602 61700 3634
rect 61686 3058 61692 3602
rect 61646 3046 61692 3058
rect 60916 3008 61404 3014
rect 60916 2974 60928 3008
rect 61392 2974 61404 3008
rect 60916 2968 61404 2974
rect 60614 2756 60620 2816
rect 60680 2756 60686 2816
rect 60452 2654 61696 2714
rect 59899 2607 60387 2613
rect 59899 2573 59911 2607
rect 60375 2573 60387 2607
rect 59899 2567 60387 2573
rect 59606 2486 59617 2523
rect 58633 1947 58639 2480
rect 59611 1980 59617 2486
rect 58593 1935 58639 1947
rect 59602 1947 59617 1980
rect 59651 2486 59666 2523
rect 60622 2523 60682 2654
rect 61140 2613 61200 2654
rect 60917 2607 61405 2613
rect 60917 2573 60929 2607
rect 61393 2573 61405 2607
rect 60917 2567 61405 2573
rect 59651 1980 59657 2486
rect 60622 2482 60635 2523
rect 59651 1947 59662 1980
rect 57863 1897 58351 1903
rect 57863 1863 57875 1897
rect 58339 1863 58351 1897
rect 57863 1857 58351 1863
rect 58881 1897 59369 1903
rect 58881 1863 58893 1897
rect 59357 1863 59369 1897
rect 58881 1857 59369 1863
rect 57562 1762 57568 1822
rect 57628 1762 57634 1822
rect 56844 1494 57332 1500
rect 56844 1460 56856 1494
rect 57320 1460 57332 1494
rect 56844 1454 57332 1460
rect 56550 1366 56562 1410
rect 55578 834 55592 874
rect 56556 868 56562 1366
rect 55532 670 55592 834
rect 56548 834 56562 868
rect 56596 1366 56610 1410
rect 57568 1410 57628 1762
rect 58074 1500 58134 1857
rect 58578 1554 58584 1614
rect 58644 1554 58650 1614
rect 57862 1494 58350 1500
rect 57862 1460 57874 1494
rect 58338 1460 58350 1494
rect 57862 1454 58350 1460
rect 56596 868 56602 1366
rect 56596 834 56608 868
rect 55826 784 56314 790
rect 55826 750 55838 784
rect 56302 750 56314 784
rect 55826 744 56314 750
rect 56040 670 56100 744
rect 56548 670 56608 834
rect 57568 834 57580 1410
rect 57614 834 57628 1410
rect 58584 1410 58644 1554
rect 59098 1500 59158 1857
rect 59602 1828 59662 1947
rect 60629 1947 60635 2482
rect 60669 2482 60682 2523
rect 61636 2523 61696 2654
rect 61636 2488 61653 2523
rect 60669 1947 60675 2482
rect 60629 1935 60675 1947
rect 61647 1947 61653 2488
rect 61687 2488 61696 2523
rect 61687 1947 61693 2488
rect 61647 1935 61693 1947
rect 59899 1897 60387 1903
rect 59899 1863 59911 1897
rect 60375 1863 60387 1897
rect 59899 1857 60387 1863
rect 60917 1897 61405 1903
rect 60917 1863 60929 1897
rect 61393 1863 61405 1897
rect 60917 1857 61405 1863
rect 59598 1822 59662 1828
rect 59658 1762 59662 1822
rect 59598 1756 59662 1762
rect 58880 1494 59368 1500
rect 58880 1460 58892 1494
rect 59356 1460 59368 1494
rect 58880 1454 59368 1460
rect 58584 1358 58598 1410
rect 56844 784 57332 790
rect 56844 750 56856 784
rect 57320 750 57332 784
rect 56844 744 57332 750
rect 57054 670 57114 744
rect 55532 610 57054 670
rect 57114 610 57120 670
rect 52622 -576 52734 210
rect 57568 110 57628 834
rect 58592 834 58598 1358
rect 58632 1358 58644 1410
rect 59602 1410 59662 1756
rect 60114 1500 60174 1857
rect 61748 1720 61808 3764
rect 62280 2920 62340 4900
rect 62412 3926 62472 5140
rect 62828 5060 62888 5066
rect 65902 5060 65962 7622
rect 62826 5000 62828 5006
rect 64012 5000 64018 5060
rect 64078 5000 64084 5060
rect 65206 5000 65212 5060
rect 65272 5000 65278 5060
rect 65896 5000 65902 5060
rect 65962 5000 65968 5060
rect 62826 4965 62888 5000
rect 62523 4903 62888 4965
rect 62523 4748 62585 4903
rect 62675 4838 62737 4903
rect 62642 4832 62770 4838
rect 62642 4798 62654 4832
rect 62758 4798 62770 4832
rect 62642 4792 62770 4798
rect 62826 4748 62888 4903
rect 63266 4900 63272 4960
rect 63332 4900 63338 4960
rect 63564 4900 63570 4960
rect 63630 4900 63636 4960
rect 63272 4838 63332 4900
rect 63570 4838 63630 4900
rect 62940 4832 63068 4838
rect 62940 4798 62952 4832
rect 63056 4798 63068 4832
rect 62940 4792 63068 4798
rect 63238 4832 63366 4838
rect 63238 4798 63250 4832
rect 63354 4798 63366 4832
rect 63238 4792 63366 4798
rect 63536 4832 63664 4838
rect 63536 4798 63548 4832
rect 63652 4798 63664 4832
rect 63536 4792 63664 4798
rect 63834 4832 63962 4838
rect 63834 4798 63846 4832
rect 63950 4798 63962 4832
rect 63834 4792 63962 4798
rect 62523 4715 62540 4748
rect 62534 4172 62540 4715
rect 62574 4716 62588 4748
rect 62574 4715 62585 4716
rect 62574 4172 62580 4715
rect 62826 4708 62838 4748
rect 62828 4696 62838 4708
rect 62534 4160 62580 4172
rect 62832 4172 62838 4696
rect 62872 4696 62888 4748
rect 63130 4748 63176 4760
rect 62872 4172 62878 4696
rect 63130 4221 63136 4748
rect 62832 4160 62878 4172
rect 63121 4172 63136 4221
rect 63170 4221 63176 4748
rect 63428 4748 63474 4760
rect 63428 4228 63434 4748
rect 63170 4172 63179 4221
rect 63420 4208 63434 4228
rect 62642 4122 62770 4128
rect 62642 4088 62654 4122
rect 62758 4088 62770 4122
rect 62642 4082 62770 4088
rect 62940 4122 63068 4128
rect 62940 4088 62952 4122
rect 63056 4088 63068 4122
rect 62940 4082 63068 4088
rect 62824 3926 62884 3932
rect 62402 3866 62408 3926
rect 62468 3866 62474 3926
rect 62884 3866 62886 3876
rect 62824 3836 62886 3866
rect 62528 3776 62886 3836
rect 62976 3818 63036 4082
rect 63121 4057 63179 4172
rect 63418 4172 63434 4208
rect 63468 4228 63474 4748
rect 63726 4748 63772 4760
rect 63468 4172 63480 4228
rect 63726 4186 63732 4748
rect 63720 4172 63732 4186
rect 63766 4186 63772 4748
rect 64018 4748 64078 5000
rect 64460 4900 64466 4960
rect 64526 4900 64532 4960
rect 64756 4900 64762 4960
rect 64822 4900 64828 4960
rect 64466 4838 64526 4900
rect 64762 4838 64822 4900
rect 64132 4832 64260 4838
rect 64132 4798 64144 4832
rect 64248 4798 64260 4832
rect 64132 4792 64260 4798
rect 64430 4832 64558 4838
rect 64430 4798 64442 4832
rect 64546 4798 64558 4832
rect 64430 4792 64558 4798
rect 64728 4832 64856 4838
rect 64728 4798 64740 4832
rect 64844 4798 64856 4832
rect 64728 4792 64856 4798
rect 65026 4832 65154 4838
rect 65026 4798 65038 4832
rect 65142 4798 65154 4832
rect 65026 4792 65154 4798
rect 64018 4688 64030 4748
rect 63766 4179 63780 4186
rect 63766 4172 63783 4179
rect 63238 4122 63366 4128
rect 63238 4088 63250 4122
rect 63354 4088 63366 4122
rect 63238 4082 63366 4088
rect 63115 3999 63121 4057
rect 63179 3999 63185 4057
rect 62528 3636 62588 3776
rect 62676 3726 62736 3776
rect 62642 3720 62770 3726
rect 62642 3686 62654 3720
rect 62758 3686 62770 3720
rect 62642 3680 62770 3686
rect 62528 3588 62540 3636
rect 62534 3060 62540 3588
rect 62574 3588 62588 3636
rect 62824 3636 62886 3776
rect 62970 3758 62976 3818
rect 63036 3758 63042 3818
rect 62940 3720 63068 3726
rect 62940 3686 62952 3720
rect 63056 3686 63068 3720
rect 62940 3680 63068 3686
rect 62824 3598 62838 3636
rect 62574 3060 62580 3588
rect 62826 3586 62838 3598
rect 62832 3100 62838 3586
rect 62534 3048 62580 3060
rect 62824 3060 62838 3100
rect 62872 3586 62886 3636
rect 63121 3636 63179 3999
rect 63418 3926 63478 4172
rect 63536 4122 63664 4128
rect 63536 4088 63548 4122
rect 63652 4088 63664 4122
rect 63536 4082 63664 4088
rect 63720 4057 63783 4172
rect 64024 4172 64030 4688
rect 64064 4688 64078 4748
rect 64322 4748 64368 4760
rect 64064 4172 64070 4688
rect 64322 4195 64328 4748
rect 64024 4160 64070 4172
rect 64316 4172 64328 4195
rect 64362 4195 64368 4748
rect 64620 4748 64666 4760
rect 64620 4230 64626 4748
rect 64612 4214 64626 4230
rect 64362 4172 64374 4195
rect 63834 4122 63962 4128
rect 63834 4088 63846 4122
rect 63950 4088 63962 4122
rect 63834 4082 63962 4088
rect 64132 4122 64260 4128
rect 64132 4088 64144 4122
rect 64248 4088 64260 4122
rect 64132 4082 64260 4088
rect 63719 3999 63725 4057
rect 63783 3999 63789 4057
rect 63412 3866 63418 3926
rect 63478 3866 63484 3926
rect 63268 3758 63274 3818
rect 63334 3758 63340 3818
rect 63568 3758 63574 3818
rect 63634 3758 63640 3818
rect 63274 3726 63334 3758
rect 63574 3726 63634 3758
rect 63238 3720 63366 3726
rect 63238 3686 63250 3720
rect 63354 3686 63366 3720
rect 63238 3680 63366 3686
rect 63536 3720 63664 3726
rect 63536 3686 63548 3720
rect 63652 3686 63664 3720
rect 63536 3680 63664 3686
rect 63121 3605 63136 3636
rect 62872 3100 62878 3586
rect 63130 3100 63136 3605
rect 62872 3060 62884 3100
rect 62642 3010 62770 3016
rect 62642 2976 62654 3010
rect 62758 2976 62770 3010
rect 62642 2970 62770 2976
rect 62274 2860 62280 2920
rect 62340 2860 62346 2920
rect 60612 1660 60618 1720
rect 60678 1660 60684 1720
rect 61742 1660 61748 1720
rect 61808 1660 61814 1720
rect 59898 1494 60386 1500
rect 59898 1460 59910 1494
rect 60374 1460 60386 1494
rect 59898 1454 60386 1460
rect 58632 834 58638 1358
rect 58592 822 58638 834
rect 59602 834 59616 1410
rect 59650 834 59662 1410
rect 60618 1410 60678 1660
rect 60916 1494 61404 1500
rect 60916 1460 60928 1494
rect 61392 1460 61404 1494
rect 60916 1454 61404 1460
rect 60618 1370 60634 1410
rect 60628 890 60634 1370
rect 57862 784 58350 790
rect 57862 750 57874 784
rect 58338 750 58350 784
rect 57862 744 58350 750
rect 58880 784 59368 790
rect 58880 750 58892 784
rect 59356 750 59368 784
rect 58880 744 59368 750
rect 58080 670 58140 744
rect 59104 670 59164 744
rect 58074 610 58080 670
rect 58140 610 58146 670
rect 59098 610 59104 670
rect 59164 610 59170 670
rect 59602 110 59662 834
rect 60622 834 60634 890
rect 60668 1370 60678 1410
rect 61646 1410 61692 1422
rect 60668 890 60674 1370
rect 60668 834 60682 890
rect 61646 874 61652 1410
rect 59898 784 60386 790
rect 59898 750 59910 784
rect 60374 750 60386 784
rect 59898 744 60386 750
rect 60004 670 60064 676
rect 60106 670 60166 744
rect 60622 670 60682 834
rect 61638 834 61652 874
rect 61686 874 61692 1410
rect 61686 834 61698 874
rect 60916 784 61404 790
rect 60916 750 60928 784
rect 61392 750 61404 784
rect 60916 744 61404 750
rect 61130 670 61190 744
rect 61638 670 61698 834
rect 62280 700 62340 2860
rect 62640 2608 62768 2614
rect 62640 2574 62652 2608
rect 62756 2574 62768 2608
rect 62640 2568 62768 2574
rect 62532 2524 62578 2536
rect 62532 1996 62538 2524
rect 62526 1948 62538 1996
rect 62572 1996 62578 2524
rect 62824 2524 62884 3060
rect 63122 3060 63136 3100
rect 63170 3605 63179 3636
rect 63428 3636 63474 3648
rect 63170 3100 63176 3605
rect 63428 3100 63434 3636
rect 63170 3060 63182 3100
rect 62978 3016 63026 3018
rect 62940 3010 63068 3016
rect 62940 2976 62952 3010
rect 63056 2976 63068 3010
rect 62940 2970 63068 2976
rect 62974 2920 63034 2970
rect 62968 2860 62974 2920
rect 63034 2860 63040 2920
rect 62974 2614 63034 2860
rect 62938 2608 63066 2614
rect 62938 2574 62950 2608
rect 63054 2574 63066 2608
rect 62938 2568 63066 2574
rect 62824 2486 62836 2524
rect 62572 1948 62586 1996
rect 62830 1994 62836 2486
rect 62526 1800 62586 1948
rect 62822 1948 62836 1994
rect 62870 2486 62884 2524
rect 63122 2524 63182 3060
rect 63420 3060 63434 3100
rect 63468 3100 63474 3636
rect 63720 3636 63783 3999
rect 63868 3818 63928 4082
rect 64010 3866 64016 3926
rect 64076 3866 64082 3926
rect 63862 3758 63868 3818
rect 63928 3758 63934 3818
rect 63834 3720 63962 3726
rect 63834 3686 63846 3720
rect 63950 3686 63962 3720
rect 63834 3680 63962 3686
rect 63720 3623 63732 3636
rect 63468 3060 63480 3100
rect 63726 3060 63732 3623
rect 63766 3623 63783 3636
rect 64016 3636 64076 3866
rect 64164 3818 64224 4082
rect 64316 4057 64374 4172
rect 64610 4172 64626 4214
rect 64660 4230 64666 4748
rect 64918 4748 64964 4760
rect 64660 4172 64672 4230
rect 64918 4223 64924 4748
rect 64913 4202 64924 4223
rect 64912 4172 64924 4202
rect 64958 4223 64964 4748
rect 65212 4748 65272 5000
rect 65324 4832 65452 4838
rect 65324 4798 65336 4832
rect 65440 4798 65452 4832
rect 65324 4792 65452 4798
rect 65622 4832 65750 4838
rect 65622 4798 65634 4832
rect 65738 4798 65750 4832
rect 65622 4792 65750 4798
rect 65212 4692 65222 4748
rect 64958 4202 64971 4223
rect 64958 4172 64972 4202
rect 64430 4122 64558 4128
rect 64430 4088 64442 4122
rect 64546 4088 64558 4122
rect 64430 4082 64558 4088
rect 64310 3999 64316 4057
rect 64374 3999 64380 4057
rect 64158 3758 64164 3818
rect 64224 3758 64230 3818
rect 64132 3720 64260 3726
rect 64132 3686 64144 3720
rect 64248 3686 64260 3720
rect 64132 3680 64260 3686
rect 63766 3060 63772 3623
rect 64016 3586 64030 3636
rect 64024 3060 64030 3586
rect 64064 3586 64076 3636
rect 64316 3636 64374 3999
rect 64610 3926 64670 4172
rect 64728 4122 64856 4128
rect 64728 4088 64740 4122
rect 64844 4088 64856 4122
rect 64728 4082 64856 4088
rect 64912 4057 64972 4172
rect 65216 4172 65222 4692
rect 65256 4692 65272 4748
rect 65514 4748 65560 4760
rect 65256 4172 65262 4692
rect 65514 4217 65520 4748
rect 65509 4210 65520 4217
rect 65216 4160 65262 4172
rect 65506 4172 65520 4210
rect 65554 4217 65560 4748
rect 65812 4748 65858 4760
rect 65554 4172 65567 4217
rect 65812 4212 65818 4748
rect 65026 4122 65154 4128
rect 65026 4088 65038 4122
rect 65142 4088 65154 4122
rect 65026 4082 65154 4088
rect 65324 4122 65452 4128
rect 65324 4088 65336 4122
rect 65440 4088 65452 4122
rect 65324 4082 65452 4088
rect 64912 3999 64913 4057
rect 64971 3999 64972 4057
rect 64604 3866 64610 3926
rect 64670 3866 64676 3926
rect 64458 3758 64464 3818
rect 64524 3758 64530 3818
rect 64760 3758 64766 3818
rect 64826 3758 64832 3818
rect 64464 3726 64524 3758
rect 64766 3726 64826 3758
rect 64430 3720 64558 3726
rect 64430 3686 64442 3720
rect 64546 3686 64558 3720
rect 64430 3680 64558 3686
rect 64728 3720 64856 3726
rect 64728 3686 64740 3720
rect 64844 3686 64856 3720
rect 64728 3680 64856 3686
rect 64620 3636 64666 3648
rect 64316 3607 64328 3636
rect 64064 3060 64070 3586
rect 64322 3066 64328 3607
rect 63238 3010 63366 3016
rect 63238 2976 63250 3010
rect 63354 2976 63366 3010
rect 63238 2970 63366 2976
rect 63420 2812 63480 3060
rect 63536 3010 63664 3016
rect 63536 2976 63548 3010
rect 63652 2976 63664 3010
rect 63536 2970 63664 2976
rect 63414 2752 63420 2812
rect 63480 2752 63486 2812
rect 63236 2608 63364 2614
rect 63236 2574 63248 2608
rect 63352 2574 63364 2608
rect 63236 2568 63364 2574
rect 63122 2486 63134 2524
rect 62870 1998 62876 2486
rect 63128 2002 63134 2486
rect 62870 1948 62890 1998
rect 63122 1948 63134 2002
rect 63168 2486 63182 2524
rect 63420 2524 63480 2752
rect 63534 2608 63662 2614
rect 63534 2574 63546 2608
rect 63650 2574 63662 2608
rect 63534 2568 63662 2574
rect 63720 2524 63780 3060
rect 64024 3048 64070 3060
rect 64314 3060 64328 3066
rect 64362 3608 64378 3636
rect 64362 3607 64374 3608
rect 64362 3066 64368 3607
rect 64620 3116 64626 3636
rect 64614 3102 64626 3116
rect 64362 3060 64374 3066
rect 64612 3060 64626 3102
rect 64660 3116 64666 3636
rect 64912 3636 64972 3999
rect 65056 3818 65116 4082
rect 65202 3866 65208 3926
rect 65268 3866 65274 3926
rect 65050 3758 65056 3818
rect 65116 3758 65122 3818
rect 65026 3720 65154 3726
rect 65026 3686 65038 3720
rect 65142 3686 65154 3720
rect 65026 3680 65154 3686
rect 64912 3616 64924 3636
rect 64660 3060 64674 3116
rect 64918 3060 64924 3616
rect 64958 3616 64972 3636
rect 65208 3636 65268 3866
rect 65360 3818 65420 4082
rect 65506 4057 65567 4172
rect 65804 4172 65818 4212
rect 65852 4212 65858 4748
rect 65852 4172 65864 4212
rect 65622 4122 65750 4128
rect 65622 4088 65634 4122
rect 65738 4088 65750 4122
rect 65622 4082 65750 4088
rect 65506 4048 65509 4057
rect 65508 3999 65509 4048
rect 65660 4054 65720 4082
rect 65804 4054 65864 4172
rect 65567 3999 65864 4054
rect 65508 3994 65864 3999
rect 65508 3842 65568 3994
rect 65354 3758 65360 3818
rect 65420 3758 65426 3818
rect 65508 3782 65866 3842
rect 65324 3720 65452 3726
rect 65324 3686 65336 3720
rect 65440 3686 65452 3720
rect 65324 3680 65452 3686
rect 64958 3060 64964 3616
rect 65208 3586 65222 3636
rect 65216 3060 65222 3586
rect 65256 3586 65268 3636
rect 65508 3636 65568 3782
rect 65656 3726 65716 3782
rect 65622 3720 65750 3726
rect 65622 3686 65634 3720
rect 65738 3686 65750 3720
rect 65622 3680 65750 3686
rect 65508 3604 65520 3636
rect 65256 3060 65262 3586
rect 65514 3104 65520 3604
rect 63834 3010 63962 3016
rect 63834 2976 63846 3010
rect 63950 2976 63962 3010
rect 63834 2970 63962 2976
rect 64132 3010 64260 3016
rect 64132 2976 64144 3010
rect 64248 2976 64260 3010
rect 64132 2970 64260 2976
rect 63870 2920 63930 2970
rect 64164 2920 64224 2970
rect 63864 2860 63870 2920
rect 63930 2860 63936 2920
rect 64158 2860 64164 2920
rect 64224 2860 64230 2920
rect 63874 2614 63930 2860
rect 64164 2614 64220 2860
rect 63832 2608 63960 2614
rect 63832 2574 63844 2608
rect 63948 2574 63960 2608
rect 63832 2568 63960 2574
rect 64130 2608 64258 2614
rect 64130 2574 64142 2608
rect 64246 2574 64258 2608
rect 64130 2568 64258 2574
rect 64022 2524 64068 2536
rect 64314 2530 64374 3060
rect 64430 3010 64558 3016
rect 64430 2976 64442 3010
rect 64546 2976 64558 3010
rect 64430 2970 64558 2976
rect 64614 2812 64674 3060
rect 64728 3010 64856 3016
rect 64728 2976 64740 3010
rect 64844 2976 64856 3010
rect 64728 2970 64856 2976
rect 64608 2752 64614 2812
rect 64674 2752 64680 2812
rect 64428 2608 64556 2614
rect 64428 2574 64440 2608
rect 64544 2574 64556 2608
rect 64428 2568 64556 2574
rect 63420 2486 63432 2524
rect 63168 2002 63174 2486
rect 63168 1948 63182 2002
rect 62640 1898 62768 1904
rect 62640 1864 62652 1898
rect 62756 1864 62768 1898
rect 62640 1858 62768 1864
rect 62672 1800 62732 1858
rect 62822 1800 62882 1948
rect 62938 1898 63066 1904
rect 62938 1864 62950 1898
rect 63054 1864 63066 1898
rect 62938 1858 63066 1864
rect 63122 1828 63182 1948
rect 63426 1948 63432 2486
rect 63466 2486 63480 2524
rect 63466 1948 63472 2486
rect 63724 2008 63730 2524
rect 63426 1936 63472 1948
rect 63716 1948 63730 2008
rect 63764 2008 63770 2524
rect 63764 1948 63776 2008
rect 64022 1996 64028 2524
rect 63236 1898 63364 1904
rect 63236 1864 63248 1898
rect 63352 1864 63364 1898
rect 63236 1858 63364 1864
rect 63534 1898 63662 1904
rect 63534 1864 63546 1898
rect 63650 1864 63662 1898
rect 63534 1858 63662 1864
rect 62526 1740 62882 1800
rect 63116 1768 63122 1828
rect 63182 1768 63188 1828
rect 62524 1734 62586 1740
rect 62584 1680 62586 1734
rect 62524 1668 62584 1674
rect 62966 1566 62972 1626
rect 63032 1566 63038 1626
rect 62972 1504 63032 1566
rect 62640 1498 62768 1504
rect 62640 1464 62652 1498
rect 62756 1464 62768 1498
rect 62640 1458 62768 1464
rect 62938 1498 63066 1504
rect 62938 1464 62950 1498
rect 63054 1464 63066 1498
rect 62938 1458 63066 1464
rect 62532 1414 62578 1426
rect 62532 890 62538 1414
rect 62524 838 62538 890
rect 62572 890 62578 1414
rect 62830 1414 62876 1426
rect 62572 838 62584 890
rect 62830 886 62836 1414
rect 62524 700 62584 838
rect 62824 838 62836 886
rect 62870 886 62876 1414
rect 63122 1414 63182 1768
rect 63270 1626 63330 1858
rect 63410 1674 63416 1734
rect 63476 1674 63482 1734
rect 63264 1566 63270 1626
rect 63330 1566 63336 1626
rect 63236 1498 63364 1504
rect 63236 1464 63248 1498
rect 63352 1464 63364 1498
rect 63236 1458 63364 1464
rect 63122 1370 63134 1414
rect 62870 838 62884 886
rect 62640 788 62768 794
rect 62640 754 62652 788
rect 62756 754 62768 788
rect 62640 748 62768 754
rect 62672 700 62732 748
rect 62824 700 62884 838
rect 63128 838 63134 1370
rect 63168 1370 63182 1414
rect 63416 1414 63476 1674
rect 63566 1626 63626 1858
rect 63716 1828 63776 1948
rect 64014 1948 64028 1996
rect 64062 1996 64068 2524
rect 64320 2524 64366 2530
rect 64614 2524 64674 2752
rect 64726 2608 64854 2614
rect 64726 2574 64738 2608
rect 64842 2574 64854 2608
rect 64726 2568 64854 2574
rect 64062 1990 64074 1996
rect 64062 1948 64080 1990
rect 64320 1978 64326 2524
rect 64316 1948 64326 1978
rect 64360 1978 64366 2524
rect 64612 2486 64624 2524
rect 64360 1948 64376 1978
rect 63832 1898 63960 1904
rect 63832 1864 63844 1898
rect 63948 1864 63960 1898
rect 63832 1858 63960 1864
rect 63710 1768 63716 1828
rect 63776 1768 63782 1828
rect 63560 1566 63566 1626
rect 63626 1566 63632 1626
rect 63534 1498 63662 1504
rect 63534 1464 63546 1498
rect 63650 1464 63662 1498
rect 63534 1458 63662 1464
rect 63716 1414 63776 1768
rect 64014 1734 64074 1948
rect 64130 1898 64258 1904
rect 64130 1864 64142 1898
rect 64246 1864 64258 1898
rect 64130 1858 64258 1864
rect 64316 1828 64376 1948
rect 64618 1948 64624 2486
rect 64658 2486 64674 2524
rect 64908 2524 64968 3060
rect 65216 3048 65262 3060
rect 65504 3060 65520 3104
rect 65554 3604 65568 3636
rect 65806 3636 65866 3782
rect 65554 3104 65560 3604
rect 65806 3600 65818 3636
rect 65554 3060 65564 3104
rect 65812 3100 65818 3600
rect 65806 3060 65818 3100
rect 65852 3600 65866 3636
rect 65852 3100 65858 3600
rect 65852 3060 65866 3100
rect 65026 3010 65154 3016
rect 65026 2976 65038 3010
rect 65142 2976 65154 3010
rect 65026 2970 65154 2976
rect 65324 3010 65452 3016
rect 65324 2976 65336 3010
rect 65440 2976 65452 3010
rect 65324 2970 65452 2976
rect 65058 2920 65118 2970
rect 65360 2920 65420 2970
rect 65052 2860 65058 2920
rect 65118 2860 65124 2920
rect 65354 2860 65360 2920
rect 65420 2860 65426 2920
rect 65062 2614 65118 2860
rect 65364 2614 65420 2860
rect 65024 2608 65152 2614
rect 65024 2574 65036 2608
rect 65140 2574 65152 2608
rect 65024 2568 65152 2574
rect 65322 2608 65450 2614
rect 65322 2574 65334 2608
rect 65438 2574 65450 2608
rect 65322 2568 65450 2574
rect 64908 2496 64922 2524
rect 64658 1948 64664 2486
rect 64916 2002 64922 2496
rect 64618 1936 64664 1948
rect 64910 1948 64922 2002
rect 64956 2496 64968 2524
rect 65214 2524 65260 2536
rect 64956 2002 64962 2496
rect 64956 1948 64970 2002
rect 65214 1998 65220 2524
rect 64428 1898 64556 1904
rect 64428 1864 64440 1898
rect 64544 1864 64556 1898
rect 64428 1858 64556 1864
rect 64726 1898 64854 1904
rect 64726 1864 64738 1898
rect 64842 1864 64854 1898
rect 64726 1858 64854 1864
rect 64310 1768 64316 1828
rect 64376 1768 64382 1828
rect 64008 1674 64014 1734
rect 64074 1674 64080 1734
rect 63864 1566 63870 1626
rect 63930 1566 63936 1626
rect 64160 1566 64166 1626
rect 64226 1566 64232 1626
rect 63870 1504 63930 1566
rect 64166 1504 64226 1566
rect 63832 1498 63960 1504
rect 63832 1464 63844 1498
rect 63948 1464 63960 1498
rect 63832 1458 63960 1464
rect 64130 1498 64258 1504
rect 64130 1464 64142 1498
rect 64246 1464 64258 1498
rect 64130 1458 64258 1464
rect 63416 1380 63432 1414
rect 63168 838 63174 1370
rect 63424 1356 63432 1380
rect 63128 826 63174 838
rect 63426 838 63432 1356
rect 63466 1356 63484 1414
rect 63716 1380 63730 1414
rect 63466 838 63472 1356
rect 63426 826 63472 838
rect 63724 838 63730 1380
rect 63764 1380 63776 1414
rect 64022 1414 64068 1426
rect 63764 838 63770 1380
rect 64022 878 64028 1414
rect 64014 876 64028 878
rect 63724 826 63770 838
rect 64012 838 64028 876
rect 64062 878 64068 1414
rect 64316 1414 64376 1768
rect 64464 1626 64524 1858
rect 64606 1674 64612 1734
rect 64672 1674 64678 1734
rect 64458 1566 64464 1626
rect 64524 1566 64530 1626
rect 64428 1498 64556 1504
rect 64428 1464 64440 1498
rect 64544 1464 64556 1498
rect 64428 1458 64556 1464
rect 64316 1382 64326 1414
rect 64062 838 64074 878
rect 64320 838 64326 1382
rect 64360 1382 64376 1414
rect 64612 1414 64672 1674
rect 64760 1626 64820 1858
rect 64910 1828 64970 1948
rect 65212 1948 65220 1998
rect 65254 1998 65260 2524
rect 65504 2524 65564 3060
rect 65812 3048 65858 3060
rect 65622 3010 65750 3016
rect 65622 2976 65634 3010
rect 65738 2976 65750 3010
rect 65622 2970 65750 2976
rect 65902 2812 65962 5000
rect 65620 2608 65748 2614
rect 65620 2574 65632 2608
rect 65736 2574 65748 2608
rect 65620 2568 65748 2574
rect 65810 2524 65856 2536
rect 65254 1948 65272 1998
rect 65024 1898 65152 1904
rect 65024 1864 65036 1898
rect 65140 1864 65152 1898
rect 65024 1858 65152 1864
rect 64904 1768 64910 1828
rect 64970 1768 64976 1828
rect 64754 1566 64760 1626
rect 64820 1566 64826 1626
rect 64726 1498 64854 1504
rect 64726 1464 64738 1498
rect 64842 1464 64854 1498
rect 64726 1458 64854 1464
rect 64910 1414 64970 1768
rect 65212 1734 65272 1948
rect 65504 1948 65518 2524
rect 65552 2488 65568 2524
rect 65802 2492 65816 2524
rect 65552 1948 65564 2488
rect 65810 2000 65816 2492
rect 65802 1978 65816 2000
rect 65800 1948 65816 1978
rect 65850 2492 65862 2524
rect 65850 2000 65856 2492
rect 65850 1948 65862 2000
rect 65322 1898 65450 1904
rect 65322 1864 65334 1898
rect 65438 1864 65450 1898
rect 65322 1858 65450 1864
rect 65504 1828 65564 1948
rect 65620 1898 65748 1904
rect 65620 1864 65632 1898
rect 65736 1864 65748 1898
rect 65620 1858 65748 1864
rect 65498 1768 65504 1828
rect 65564 1824 65570 1828
rect 65652 1824 65712 1858
rect 65802 1824 65862 1948
rect 65564 1768 65862 1824
rect 65504 1764 65862 1768
rect 65206 1674 65212 1734
rect 65272 1674 65278 1734
rect 65050 1566 65056 1626
rect 65116 1566 65122 1626
rect 65354 1566 65360 1626
rect 65420 1566 65426 1626
rect 65504 1602 65564 1764
rect 65056 1504 65116 1566
rect 65360 1504 65420 1566
rect 65504 1542 65864 1602
rect 65024 1498 65152 1504
rect 65024 1464 65036 1498
rect 65140 1464 65152 1498
rect 65024 1458 65152 1464
rect 65322 1498 65450 1504
rect 65322 1464 65334 1498
rect 65438 1464 65450 1498
rect 65322 1458 65450 1464
rect 64360 838 64366 1382
rect 64612 1376 64624 1414
rect 64616 1354 64624 1376
rect 62938 788 63066 794
rect 62938 754 62950 788
rect 63054 754 63066 788
rect 62938 748 63066 754
rect 63236 788 63364 794
rect 63236 754 63248 788
rect 63352 754 63364 788
rect 63236 748 63364 754
rect 63534 788 63662 794
rect 63534 754 63546 788
rect 63650 754 63662 788
rect 63534 748 63662 754
rect 63832 788 63960 794
rect 63832 754 63844 788
rect 63948 754 63960 788
rect 63832 748 63960 754
rect 63270 700 63330 748
rect 63568 700 63628 748
rect 60064 610 61698 670
rect 62274 640 62280 700
rect 62340 640 62346 700
rect 62524 640 62884 700
rect 63264 640 63270 700
rect 63330 640 63336 700
rect 63562 640 63568 700
rect 63628 640 63634 700
rect 60004 604 60064 610
rect 62824 600 62884 640
rect 64012 600 64072 838
rect 64320 826 64366 838
rect 64618 838 64624 1354
rect 64658 1354 64676 1414
rect 64910 1388 64922 1414
rect 64658 838 64664 1354
rect 64618 826 64664 838
rect 64916 838 64922 1388
rect 64956 1388 64970 1414
rect 65214 1414 65260 1426
rect 64956 838 64962 1388
rect 65214 886 65220 1414
rect 65206 838 65220 886
rect 65254 886 65260 1414
rect 65504 1414 65564 1542
rect 65654 1504 65714 1542
rect 65620 1498 65748 1504
rect 65620 1464 65632 1498
rect 65736 1464 65748 1498
rect 65620 1458 65748 1464
rect 65504 1358 65518 1414
rect 65254 874 65266 886
rect 65254 838 65268 874
rect 64916 826 64962 838
rect 64130 788 64258 794
rect 64130 754 64142 788
rect 64246 754 64258 788
rect 64130 748 64258 754
rect 64428 788 64556 794
rect 64428 754 64440 788
rect 64544 754 64556 788
rect 64428 748 64556 754
rect 64726 788 64854 794
rect 64726 754 64738 788
rect 64842 754 64854 788
rect 64726 748 64854 754
rect 65024 788 65152 794
rect 65024 754 65036 788
rect 65140 754 65152 788
rect 65024 748 65152 754
rect 64464 700 64524 748
rect 64766 700 64826 748
rect 64458 640 64464 700
rect 64524 640 64530 700
rect 64760 640 64766 700
rect 64826 640 64832 700
rect 65208 600 65268 838
rect 65512 838 65518 1358
rect 65552 1358 65564 1414
rect 65804 1414 65864 1542
rect 65804 1388 65816 1414
rect 65552 838 65558 1358
rect 65512 826 65558 838
rect 65810 838 65816 1388
rect 65850 1388 65864 1414
rect 65850 838 65856 1388
rect 65810 826 65856 838
rect 65322 788 65450 794
rect 65322 754 65334 788
rect 65438 754 65450 788
rect 65322 748 65450 754
rect 65620 788 65748 794
rect 65620 754 65632 788
rect 65736 754 65748 788
rect 65620 748 65748 754
rect 65902 600 65962 2752
rect 66026 3818 66086 3824
rect 66026 1626 66086 3758
rect 66926 2996 66986 12480
rect 66920 2936 66926 2996
rect 66986 2936 66992 2996
rect 67060 2778 67120 12686
rect 67286 11424 67346 15124
rect 68020 14946 87432 15006
rect 68020 14900 68080 14946
rect 67814 14894 68302 14900
rect 67814 14860 67826 14894
rect 68290 14860 68302 14894
rect 67814 14854 68302 14860
rect 67526 14810 67572 14822
rect 67526 14268 67532 14810
rect 67518 14234 67532 14268
rect 67566 14268 67572 14810
rect 68536 14810 68596 14946
rect 69048 14900 69108 14946
rect 70056 14900 70116 14946
rect 68832 14894 69320 14900
rect 68832 14860 68844 14894
rect 69308 14860 69320 14894
rect 68832 14854 69320 14860
rect 69850 14894 70338 14900
rect 69850 14860 69862 14894
rect 70326 14860 70338 14894
rect 69850 14854 70338 14860
rect 67566 14234 67578 14268
rect 67518 14092 67578 14234
rect 68536 14234 68550 14810
rect 68584 14234 68596 14810
rect 69562 14810 69608 14822
rect 69562 14272 69568 14810
rect 67814 14184 68302 14190
rect 67814 14150 67826 14184
rect 68290 14150 68302 14184
rect 67814 14144 68302 14150
rect 67512 14032 67518 14092
rect 67578 14032 67584 14092
rect 67518 13576 67578 14032
rect 68026 13666 68086 14144
rect 68536 13994 68596 14234
rect 69554 14234 69568 14272
rect 69602 14272 69608 14810
rect 70574 14810 70634 14946
rect 71066 14900 71126 14946
rect 72078 14900 72138 14946
rect 70868 14894 71356 14900
rect 70868 14860 70880 14894
rect 71344 14860 71356 14894
rect 70868 14854 71356 14860
rect 71886 14894 72374 14900
rect 71886 14860 71898 14894
rect 72362 14860 72374 14894
rect 71886 14854 72374 14860
rect 69602 14234 69614 14272
rect 68832 14184 69320 14190
rect 68832 14150 68844 14184
rect 69308 14150 69320 14184
rect 68832 14144 69320 14150
rect 68530 13934 68536 13994
rect 68596 13934 68602 13994
rect 67814 13660 68302 13666
rect 67814 13626 67826 13660
rect 68290 13626 68302 13660
rect 67814 13620 68302 13626
rect 67518 13542 67532 13576
rect 67526 13000 67532 13542
rect 67566 13542 67578 13576
rect 68536 13576 68596 13934
rect 69028 13666 69088 14144
rect 69554 14092 69614 14234
rect 70574 14234 70586 14810
rect 70620 14234 70634 14810
rect 71598 14810 71644 14822
rect 71598 14264 71604 14810
rect 70050 14190 70110 14192
rect 69850 14184 70338 14190
rect 69850 14150 69862 14184
rect 70326 14150 70338 14184
rect 69850 14144 70338 14150
rect 69548 14032 69554 14092
rect 69614 14032 69620 14092
rect 68832 13660 69320 13666
rect 68832 13626 68844 13660
rect 69308 13626 69320 13660
rect 68832 13620 69320 13626
rect 67566 13000 67572 13542
rect 68536 13528 68550 13576
rect 67526 12988 67572 13000
rect 68544 13000 68550 13528
rect 68584 13528 68596 13576
rect 69554 13576 69614 14032
rect 70050 13666 70110 14144
rect 70574 13994 70634 14234
rect 71588 14234 71604 14264
rect 71638 14264 71644 14810
rect 72608 14810 72668 14946
rect 73126 14900 73186 14946
rect 74114 14900 74174 14946
rect 72904 14894 73392 14900
rect 72904 14860 72916 14894
rect 73380 14860 73392 14894
rect 72904 14854 73392 14860
rect 73922 14894 74410 14900
rect 73922 14860 73934 14894
rect 74398 14860 74410 14894
rect 73922 14854 74410 14860
rect 71638 14234 71648 14264
rect 70868 14184 71356 14190
rect 70868 14150 70880 14184
rect 71344 14150 71356 14184
rect 70868 14144 71356 14150
rect 71588 14092 71648 14234
rect 72608 14234 72622 14810
rect 72656 14234 72668 14810
rect 73634 14810 73680 14822
rect 73634 14278 73640 14810
rect 71886 14184 72374 14190
rect 71886 14150 71898 14184
rect 72362 14150 72374 14184
rect 71886 14144 72374 14150
rect 71582 14032 71588 14092
rect 71648 14032 71654 14092
rect 72608 13994 72668 14234
rect 73628 14234 73640 14278
rect 73674 14278 73680 14810
rect 74642 14810 74702 14946
rect 75158 14900 75218 14946
rect 76160 14900 76220 14946
rect 74940 14894 75428 14900
rect 74940 14860 74952 14894
rect 75416 14860 75428 14894
rect 74940 14854 75428 14860
rect 75958 14894 76446 14900
rect 75958 14860 75970 14894
rect 76434 14860 76446 14894
rect 75958 14854 76446 14860
rect 73674 14234 73688 14278
rect 72904 14184 73392 14190
rect 72904 14150 72916 14184
rect 73380 14150 73392 14184
rect 72904 14144 73392 14150
rect 73628 14092 73688 14234
rect 74642 14234 74658 14810
rect 74692 14234 74702 14810
rect 75670 14810 75716 14822
rect 75670 14274 75676 14810
rect 73922 14184 74410 14190
rect 73922 14150 73934 14184
rect 74398 14150 74410 14184
rect 73922 14144 74410 14150
rect 73622 14032 73628 14092
rect 73688 14032 73694 14092
rect 74642 13994 74702 14234
rect 75664 14234 75676 14274
rect 75710 14274 75716 14810
rect 76682 14810 76742 14946
rect 77188 14900 77248 14946
rect 78206 14900 78266 14946
rect 76976 14894 77464 14900
rect 76976 14860 76988 14894
rect 77452 14860 77464 14894
rect 76976 14854 77464 14860
rect 77994 14894 78482 14900
rect 77994 14860 78006 14894
rect 78470 14860 78482 14894
rect 77994 14854 78482 14860
rect 77188 14852 77248 14854
rect 75710 14234 75724 14274
rect 74940 14184 75428 14190
rect 74940 14150 74952 14184
rect 75416 14150 75428 14184
rect 74940 14144 75428 14150
rect 75664 14092 75724 14234
rect 76682 14234 76694 14810
rect 76728 14234 76742 14810
rect 77706 14810 77752 14822
rect 77706 14274 77712 14810
rect 75958 14184 76446 14190
rect 75958 14150 75970 14184
rect 76434 14150 76446 14184
rect 75958 14144 76446 14150
rect 75658 14032 75664 14092
rect 75724 14032 75730 14092
rect 76682 13994 76742 14234
rect 77698 14234 77712 14274
rect 77746 14274 77752 14810
rect 78716 14810 78776 14946
rect 79224 14900 79284 14946
rect 80244 14900 80304 14946
rect 79012 14894 79500 14900
rect 79012 14860 79024 14894
rect 79488 14860 79500 14894
rect 79012 14854 79500 14860
rect 80030 14894 80518 14900
rect 80030 14860 80042 14894
rect 80506 14860 80518 14894
rect 80030 14854 80518 14860
rect 77746 14234 77758 14274
rect 76976 14184 77464 14190
rect 76976 14150 76988 14184
rect 77452 14150 77464 14184
rect 76976 14144 77464 14150
rect 77698 14092 77758 14234
rect 78716 14234 78730 14810
rect 78764 14234 78776 14810
rect 79742 14810 79788 14822
rect 79742 14280 79748 14810
rect 77994 14184 78482 14190
rect 77994 14150 78006 14184
rect 78470 14150 78482 14184
rect 77994 14144 78482 14150
rect 77692 14032 77698 14092
rect 77758 14032 77764 14092
rect 78716 13994 78776 14234
rect 79734 14234 79748 14280
rect 79782 14280 79788 14810
rect 80754 14810 80814 14946
rect 81252 14900 81312 14946
rect 82280 14900 82340 14946
rect 81048 14894 81536 14900
rect 81048 14860 81060 14894
rect 81524 14860 81536 14894
rect 81048 14854 81536 14860
rect 82066 14894 82554 14900
rect 82066 14860 82078 14894
rect 82542 14860 82554 14894
rect 82066 14854 82554 14860
rect 79782 14234 79794 14280
rect 79012 14184 79500 14190
rect 79012 14150 79024 14184
rect 79488 14150 79500 14184
rect 79012 14144 79500 14150
rect 79734 14092 79794 14234
rect 80754 14234 80766 14810
rect 80800 14234 80814 14810
rect 81778 14810 81824 14822
rect 81778 14282 81784 14810
rect 80030 14184 80518 14190
rect 80030 14150 80042 14184
rect 80506 14150 80518 14184
rect 80030 14144 80518 14150
rect 79728 14032 79734 14092
rect 79794 14032 79800 14092
rect 80754 13994 80814 14234
rect 81770 14234 81784 14282
rect 81818 14282 81824 14810
rect 82786 14810 82846 14946
rect 83282 14900 83342 14946
rect 84312 14900 84372 14946
rect 83084 14894 83572 14900
rect 83084 14860 83096 14894
rect 83560 14860 83572 14894
rect 83084 14854 83572 14860
rect 84102 14894 84590 14900
rect 84102 14860 84114 14894
rect 84578 14860 84590 14894
rect 84102 14854 84590 14860
rect 81818 14234 81830 14282
rect 81048 14184 81536 14190
rect 81048 14150 81060 14184
rect 81524 14150 81536 14184
rect 81048 14144 81536 14150
rect 81770 14092 81830 14234
rect 82786 14234 82802 14810
rect 82836 14234 82846 14810
rect 83814 14810 83860 14822
rect 83814 14288 83820 14810
rect 82066 14184 82554 14190
rect 82066 14150 82078 14184
rect 82542 14150 82554 14184
rect 82066 14144 82554 14150
rect 81764 14032 81770 14092
rect 81830 14032 81836 14092
rect 82786 13994 82846 14234
rect 83806 14234 83820 14288
rect 83854 14288 83860 14810
rect 84824 14810 84884 14946
rect 85360 14900 85420 14946
rect 86334 14900 86394 14946
rect 85120 14894 85608 14900
rect 85120 14860 85132 14894
rect 85596 14860 85608 14894
rect 85120 14854 85608 14860
rect 86138 14894 86626 14900
rect 86138 14860 86150 14894
rect 86614 14860 86626 14894
rect 86138 14854 86626 14860
rect 83854 14234 83866 14288
rect 83084 14184 83572 14190
rect 83084 14150 83096 14184
rect 83560 14150 83572 14184
rect 83084 14144 83572 14150
rect 83806 14092 83866 14234
rect 84824 14234 84838 14810
rect 84872 14234 84884 14810
rect 85850 14810 85896 14822
rect 85850 14280 85856 14810
rect 84102 14184 84590 14190
rect 84102 14150 84114 14184
rect 84578 14150 84590 14184
rect 84102 14144 84590 14150
rect 83800 14032 83806 14092
rect 83866 14032 83872 14092
rect 84824 13994 84884 14234
rect 85844 14234 85856 14280
rect 85890 14280 85896 14810
rect 86862 14810 86922 14946
rect 87372 14900 87432 14946
rect 87156 14894 87644 14900
rect 87156 14860 87168 14894
rect 87632 14860 87644 14894
rect 87156 14854 87644 14860
rect 85890 14234 85904 14280
rect 85120 14184 85608 14190
rect 85120 14150 85132 14184
rect 85596 14150 85608 14184
rect 85120 14144 85608 14150
rect 70568 13934 70574 13994
rect 70634 13934 70640 13994
rect 72602 13934 72608 13994
rect 72668 13934 72674 13994
rect 74636 13934 74642 13994
rect 74702 13934 74708 13994
rect 76676 13934 76682 13994
rect 76742 13934 76748 13994
rect 78710 13934 78716 13994
rect 78776 13934 78782 13994
rect 80748 13934 80754 13994
rect 80814 13934 80820 13994
rect 82780 13934 82786 13994
rect 82846 13934 82852 13994
rect 84818 13934 84824 13994
rect 84884 13934 84890 13994
rect 77168 13880 77228 13888
rect 77168 13820 79276 13880
rect 74140 13702 75210 13762
rect 76676 13722 76682 13782
rect 76742 13722 76748 13782
rect 74140 13666 74200 13702
rect 69850 13660 70338 13666
rect 69850 13626 69862 13660
rect 70326 13626 70338 13660
rect 69850 13620 70338 13626
rect 70868 13660 71356 13666
rect 70868 13626 70880 13660
rect 71344 13626 71356 13660
rect 70868 13620 71356 13626
rect 71886 13660 72374 13666
rect 71886 13626 71898 13660
rect 72362 13626 72374 13660
rect 71886 13620 72374 13626
rect 72904 13660 73392 13666
rect 72904 13626 72916 13660
rect 73380 13626 73392 13660
rect 72904 13620 73392 13626
rect 73922 13660 74410 13666
rect 73922 13626 73934 13660
rect 74398 13626 74410 13660
rect 73922 13620 74410 13626
rect 69554 13544 69568 13576
rect 68584 13000 68590 13528
rect 68544 12988 68590 13000
rect 69562 13000 69568 13544
rect 69602 13544 69614 13576
rect 70580 13576 70626 13588
rect 69602 13000 69608 13544
rect 70580 13028 70586 13576
rect 69562 12988 69608 13000
rect 70574 13000 70586 13028
rect 70620 13028 70626 13576
rect 71598 13576 71644 13588
rect 72616 13576 72662 13588
rect 73634 13576 73680 13588
rect 71598 13048 71604 13576
rect 70620 13000 70634 13028
rect 67814 12950 68302 12956
rect 67814 12916 67826 12950
rect 68290 12916 68302 12950
rect 67814 12910 68302 12916
rect 68832 12950 69320 12956
rect 68832 12916 68844 12950
rect 69308 12916 69320 12950
rect 68832 12910 69320 12916
rect 69850 12950 70338 12956
rect 69850 12916 69862 12950
rect 70326 12916 70338 12950
rect 69850 12910 70338 12916
rect 70574 12858 70634 13000
rect 71592 13000 71604 13048
rect 71638 13048 71644 13576
rect 72606 13542 72622 13576
rect 72616 13076 72622 13542
rect 71638 13000 71652 13048
rect 70868 12950 71356 12956
rect 70868 12916 70880 12950
rect 71344 12916 71356 12950
rect 70868 12910 71356 12916
rect 71222 12862 71282 12910
rect 71592 12862 71652 13000
rect 72606 13000 72622 13076
rect 72656 13542 72666 13576
rect 72656 13076 72662 13542
rect 72656 13060 72666 13076
rect 72656 13000 72670 13060
rect 73634 13056 73640 13576
rect 73626 13000 73640 13056
rect 73674 13056 73680 13576
rect 74646 13576 74706 13702
rect 75150 13666 75210 13702
rect 74940 13660 75428 13666
rect 74940 13626 74952 13660
rect 75416 13626 75428 13660
rect 74940 13620 75428 13626
rect 75958 13660 76446 13666
rect 75958 13626 75970 13660
rect 76434 13626 76446 13660
rect 75958 13620 76446 13626
rect 74646 13526 74658 13576
rect 73674 13000 73686 13056
rect 74652 13050 74658 13526
rect 74646 13036 74658 13050
rect 71886 12950 72374 12956
rect 71886 12916 71898 12950
rect 72362 12916 72374 12950
rect 71886 12910 72374 12916
rect 72094 12862 72154 12910
rect 72606 12862 72666 13000
rect 72904 12950 73392 12956
rect 72904 12916 72916 12950
rect 73380 12916 73392 12950
rect 72904 12910 73392 12916
rect 73134 12862 73194 12910
rect 73626 12862 73686 13000
rect 74644 13000 74658 13036
rect 74692 13526 74706 13576
rect 75670 13576 75716 13588
rect 74692 13050 74698 13526
rect 75670 13076 75676 13576
rect 74692 13000 74706 13050
rect 75658 13000 75676 13076
rect 75710 13076 75716 13576
rect 76682 13576 76742 13722
rect 77168 13666 77228 13820
rect 78202 13666 78262 13820
rect 78708 13722 78714 13782
rect 78774 13722 78780 13782
rect 76976 13660 77464 13666
rect 76976 13626 76988 13660
rect 77452 13626 77464 13660
rect 76976 13620 77464 13626
rect 77994 13660 78482 13666
rect 77994 13626 78006 13660
rect 78470 13626 78482 13660
rect 77994 13620 78482 13626
rect 76682 13542 76694 13576
rect 75710 13000 75718 13076
rect 76688 13062 76694 13542
rect 76682 13058 76694 13062
rect 73922 12950 74410 12956
rect 73922 12916 73934 12950
rect 74398 12916 74410 12950
rect 73922 12910 74410 12916
rect 70574 12798 71146 12858
rect 71216 12802 71222 12862
rect 71282 12802 71288 12862
rect 71586 12802 71592 12862
rect 71652 12802 71658 12862
rect 72088 12802 72094 12862
rect 72154 12802 72160 12862
rect 72600 12802 72606 12862
rect 72666 12802 72672 12862
rect 73128 12802 73134 12862
rect 73194 12802 73200 12862
rect 73620 12802 73626 12862
rect 73686 12802 73692 12862
rect 69040 12692 69046 12752
rect 69106 12692 69112 12752
rect 70062 12692 70068 12752
rect 70128 12692 70134 12752
rect 67516 12480 67522 12540
rect 67582 12480 67588 12540
rect 68014 12480 68020 12540
rect 68080 12480 68086 12540
rect 68526 12480 68532 12540
rect 68592 12480 68598 12540
rect 67522 12344 67582 12480
rect 68020 12434 68080 12480
rect 67814 12428 68302 12434
rect 67814 12394 67826 12428
rect 68290 12394 68302 12428
rect 67814 12388 68302 12394
rect 67522 12304 67532 12344
rect 67526 11768 67532 12304
rect 67566 12304 67582 12344
rect 68532 12344 68592 12480
rect 69046 12434 69106 12692
rect 70068 12434 70128 12692
rect 71086 12654 71146 12798
rect 71086 12648 71148 12654
rect 71086 12588 71088 12648
rect 71086 12582 71148 12588
rect 70568 12480 70574 12540
rect 70634 12480 70640 12540
rect 68832 12428 69320 12434
rect 68832 12394 68844 12428
rect 69308 12394 69320 12428
rect 68832 12388 69320 12394
rect 69850 12428 70338 12434
rect 69850 12394 69862 12428
rect 70326 12394 70338 12428
rect 69850 12388 70338 12394
rect 67566 11768 67572 12304
rect 68532 12298 68550 12344
rect 67526 11756 67572 11768
rect 68544 11768 68550 12298
rect 68584 12298 68592 12344
rect 69562 12344 69608 12356
rect 68584 11768 68590 12298
rect 69562 11826 69568 12344
rect 68544 11756 68590 11768
rect 69548 11768 69568 11826
rect 69602 11768 69608 12344
rect 70574 12344 70634 12480
rect 71086 12434 71146 12582
rect 70868 12428 71356 12434
rect 70868 12394 70880 12428
rect 71344 12394 71356 12428
rect 70868 12388 71356 12394
rect 70574 12292 70586 12344
rect 67814 11718 68302 11724
rect 67814 11684 67826 11718
rect 68290 11684 68302 11718
rect 67814 11678 68302 11684
rect 68832 11718 69320 11724
rect 68832 11684 68844 11718
rect 69308 11684 69320 11718
rect 68832 11678 69320 11684
rect 69030 11578 69036 11638
rect 69096 11578 69102 11638
rect 67280 11364 67286 11424
rect 67346 11364 67352 11424
rect 67286 10182 67346 11364
rect 67518 11268 68596 11328
rect 67518 11110 67578 11268
rect 68026 11200 68086 11268
rect 67812 11194 68300 11200
rect 67812 11160 67824 11194
rect 68288 11160 68300 11194
rect 67812 11154 68300 11160
rect 67518 11084 67530 11110
rect 67524 10534 67530 11084
rect 67564 11084 67578 11110
rect 68536 11110 68596 11268
rect 69036 11200 69096 11578
rect 69548 11546 69608 11768
rect 70580 11768 70586 12292
rect 70620 12292 70634 12344
rect 71592 12344 71652 12802
rect 72082 12588 72088 12648
rect 72148 12588 72154 12648
rect 73102 12588 73108 12648
rect 73168 12588 73174 12648
rect 72088 12434 72148 12588
rect 72602 12480 72608 12540
rect 72668 12480 72674 12540
rect 71886 12428 72374 12434
rect 71886 12394 71898 12428
rect 72362 12394 72374 12428
rect 71886 12388 72374 12394
rect 70620 11768 70626 12292
rect 71592 12280 71604 12344
rect 71598 11832 71604 12280
rect 70580 11756 70626 11768
rect 71584 11768 71604 11832
rect 71638 12280 71652 12344
rect 72608 12344 72668 12480
rect 73108 12434 73168 12588
rect 72904 12428 73392 12434
rect 72904 12394 72916 12428
rect 73380 12394 73392 12428
rect 72904 12388 73392 12394
rect 72608 12310 72622 12344
rect 71638 11768 71644 12280
rect 69850 11718 70338 11724
rect 69850 11684 69862 11718
rect 70326 11684 70338 11718
rect 69850 11678 70338 11684
rect 70868 11718 71356 11724
rect 70868 11684 70880 11718
rect 71344 11684 71356 11718
rect 70868 11678 71356 11684
rect 71072 11650 71132 11678
rect 70046 11590 70052 11650
rect 70112 11590 70118 11650
rect 71066 11590 71072 11650
rect 71132 11590 71138 11650
rect 69542 11486 69548 11546
rect 69608 11486 69614 11546
rect 69548 11252 69554 11312
rect 69614 11252 69620 11312
rect 68830 11194 69318 11200
rect 68830 11160 68842 11194
rect 69306 11160 69318 11194
rect 68830 11154 69318 11160
rect 67564 10534 67570 11084
rect 68536 11078 68548 11110
rect 68542 10578 68548 11078
rect 67524 10522 67570 10534
rect 68536 10534 68548 10578
rect 68582 11078 68596 11110
rect 69554 11110 69614 11252
rect 70052 11200 70112 11590
rect 70566 11486 70572 11546
rect 70632 11486 70638 11546
rect 69848 11194 70336 11200
rect 69848 11160 69860 11194
rect 70324 11160 70336 11194
rect 69848 11154 70336 11160
rect 69554 11084 69566 11110
rect 68582 10578 68588 11078
rect 68582 10534 68596 10578
rect 67812 10484 68300 10490
rect 67812 10450 67824 10484
rect 68288 10450 68300 10484
rect 67812 10444 68300 10450
rect 68536 10382 68596 10534
rect 69560 10534 69566 11084
rect 69600 11084 69614 11110
rect 70572 11110 70632 11486
rect 71072 11200 71132 11590
rect 71584 11546 71644 11768
rect 72616 11768 72622 12310
rect 72656 12310 72668 12344
rect 73626 12344 73686 12802
rect 74140 12752 74200 12910
rect 74644 12752 74704 13000
rect 74940 12950 75428 12956
rect 74940 12916 74952 12950
rect 75416 12916 75428 12950
rect 74940 12910 75428 12916
rect 75160 12752 75220 12910
rect 75658 12862 75718 13000
rect 76680 13000 76694 13058
rect 76728 13542 76742 13576
rect 77706 13576 77752 13588
rect 76728 13062 76734 13542
rect 77706 13066 77712 13576
rect 76728 13000 76742 13062
rect 77694 13000 77712 13066
rect 77746 13066 77752 13576
rect 78714 13576 78774 13722
rect 79216 13666 79276 13820
rect 80240 13732 81322 13792
rect 80240 13666 80300 13732
rect 79012 13660 79500 13666
rect 79012 13626 79024 13660
rect 79488 13626 79500 13660
rect 79012 13620 79500 13626
rect 80030 13660 80518 13666
rect 80030 13626 80042 13660
rect 80506 13626 80518 13660
rect 80030 13620 80518 13626
rect 78714 13542 78730 13576
rect 77746 13000 77754 13066
rect 78724 13026 78730 13542
rect 75958 12950 76446 12956
rect 75958 12916 75970 12950
rect 76434 12916 76446 12950
rect 75958 12910 76446 12916
rect 75652 12802 75658 12862
rect 75718 12802 75724 12862
rect 74134 12692 74140 12752
rect 74200 12692 74206 12752
rect 74638 12692 74644 12752
rect 74704 12692 74710 12752
rect 75154 12692 75160 12752
rect 75220 12692 75226 12752
rect 74140 12434 74200 12692
rect 74636 12480 74642 12540
rect 74702 12480 74708 12540
rect 73922 12428 74410 12434
rect 73922 12394 73934 12428
rect 74398 12394 74410 12428
rect 73922 12388 74410 12394
rect 72656 11768 72662 12310
rect 73626 12302 73640 12344
rect 73634 11810 73640 12302
rect 72616 11756 72662 11768
rect 73626 11768 73640 11810
rect 73674 12302 73686 12344
rect 74642 12344 74702 12480
rect 75160 12434 75220 12692
rect 74940 12428 75428 12434
rect 74940 12394 74952 12428
rect 75416 12394 75428 12428
rect 74940 12388 75428 12394
rect 73674 11810 73680 12302
rect 74642 12282 74658 12344
rect 73674 11768 73686 11810
rect 71886 11718 72374 11724
rect 71886 11684 71898 11718
rect 72362 11684 72374 11718
rect 71886 11678 72374 11684
rect 72904 11718 73392 11724
rect 72904 11684 72916 11718
rect 73380 11684 73392 11718
rect 72904 11678 73392 11684
rect 72084 11650 72144 11678
rect 73110 11650 73170 11678
rect 72078 11590 72084 11650
rect 72144 11590 72150 11650
rect 73104 11590 73110 11650
rect 73170 11590 73176 11650
rect 71578 11486 71584 11546
rect 71644 11486 71650 11546
rect 71584 11252 71590 11312
rect 71650 11252 71656 11312
rect 70866 11194 71354 11200
rect 70866 11160 70878 11194
rect 71342 11160 71354 11194
rect 70866 11154 71354 11160
rect 69600 10534 69606 11084
rect 70572 11078 70584 11110
rect 70578 10574 70584 11078
rect 69560 10522 69606 10534
rect 70570 10534 70584 10574
rect 70618 11078 70632 11110
rect 71590 11110 71650 11252
rect 72084 11200 72144 11590
rect 72598 11486 72604 11546
rect 72664 11486 72670 11546
rect 71884 11194 72372 11200
rect 71884 11160 71896 11194
rect 72360 11160 72372 11194
rect 71884 11154 72372 11160
rect 71590 11080 71602 11110
rect 70618 10574 70624 11078
rect 70618 10534 70630 10574
rect 68830 10484 69318 10490
rect 68830 10450 68842 10484
rect 69306 10450 69318 10484
rect 68830 10444 69318 10450
rect 69848 10484 70336 10490
rect 69848 10450 69860 10484
rect 70324 10450 70336 10484
rect 69848 10444 70336 10450
rect 67392 10322 67398 10382
rect 67458 10322 67464 10382
rect 68530 10322 68536 10382
rect 68596 10322 68602 10382
rect 67280 10122 67286 10182
rect 67346 10122 67352 10182
rect 67174 10020 67180 10080
rect 67240 10020 67246 10080
rect 67180 6590 67240 10020
rect 67286 8946 67346 10122
rect 67280 8886 67286 8946
rect 67346 8886 67352 8946
rect 67174 6530 67180 6590
rect 67240 6530 67246 6590
rect 67180 5286 67240 6530
rect 67286 6344 67346 8886
rect 67398 7608 67458 10322
rect 68528 10122 68534 10182
rect 68594 10122 68600 10182
rect 68534 10078 68594 10122
rect 67518 10018 68594 10078
rect 67518 10016 68082 10018
rect 67518 9876 67578 10016
rect 68022 9966 68082 10016
rect 67812 9960 68300 9966
rect 67812 9926 67824 9960
rect 68288 9926 68300 9960
rect 67812 9920 68300 9926
rect 67518 9844 67530 9876
rect 67524 9300 67530 9844
rect 67564 9844 67578 9876
rect 68534 9876 68594 10018
rect 69038 9966 69098 10444
rect 69546 10242 69552 10302
rect 69612 10242 69618 10302
rect 68830 9960 69318 9966
rect 68830 9926 68842 9960
rect 69306 9926 69318 9960
rect 68830 9920 69318 9926
rect 67564 9300 67570 9844
rect 68534 9840 68548 9876
rect 67524 9288 67570 9300
rect 68542 9300 68548 9840
rect 68582 9840 68594 9876
rect 69552 9876 69612 10242
rect 70066 10188 70126 10444
rect 70570 10406 70630 10534
rect 71596 10534 71602 11080
rect 71636 11080 71650 11110
rect 72604 11110 72664 11486
rect 73110 11200 73170 11590
rect 73626 11546 73686 11768
rect 74652 11768 74658 12282
rect 74692 12282 74702 12344
rect 75658 12344 75718 12802
rect 76180 12752 76240 12910
rect 76680 12864 76740 13000
rect 76976 12950 77464 12956
rect 76976 12916 76988 12950
rect 77452 12916 77464 12950
rect 76976 12910 77464 12916
rect 76680 12804 76858 12864
rect 76174 12692 76180 12752
rect 76240 12692 76246 12752
rect 76676 12692 76682 12752
rect 76742 12692 76748 12752
rect 76180 12434 76240 12692
rect 75958 12428 76446 12434
rect 75958 12394 75970 12428
rect 76434 12394 76446 12428
rect 75958 12388 76446 12394
rect 76682 12344 76742 12692
rect 76798 12540 76858 12804
rect 77176 12692 77182 12752
rect 77242 12692 77248 12752
rect 76798 12474 76858 12480
rect 77182 12434 77242 12692
rect 77322 12648 77382 12910
rect 77694 12862 77754 13000
rect 78716 13000 78730 13026
rect 78764 13542 78774 13576
rect 79742 13576 79788 13588
rect 78764 13026 78770 13542
rect 79742 13060 79748 13576
rect 78764 13000 78776 13026
rect 77994 12950 78482 12956
rect 77994 12916 78006 12950
rect 78470 12916 78482 12950
rect 77994 12910 78482 12916
rect 77688 12802 77694 12862
rect 77754 12802 77760 12862
rect 77316 12588 77322 12648
rect 77382 12588 77388 12648
rect 76976 12428 77464 12434
rect 76976 12394 76988 12428
rect 77452 12394 77464 12428
rect 76976 12388 77464 12394
rect 75658 12288 75676 12344
rect 74692 11768 74698 12282
rect 75670 11810 75676 12288
rect 74652 11756 74698 11768
rect 75662 11768 75676 11810
rect 75710 12288 75718 12344
rect 76678 12292 76694 12344
rect 75710 11810 75716 12288
rect 76688 11816 76694 12292
rect 75710 11768 75722 11810
rect 73922 11718 74410 11724
rect 73922 11684 73934 11718
rect 74398 11684 74410 11718
rect 73922 11678 74410 11684
rect 74940 11718 75428 11724
rect 74940 11684 74952 11718
rect 75416 11684 75428 11718
rect 74940 11678 75428 11684
rect 75662 11546 75722 11768
rect 76680 11768 76694 11816
rect 76728 12300 76742 12344
rect 77694 12344 77754 12802
rect 78202 12692 78208 12752
rect 78268 12692 78274 12752
rect 78208 12434 78268 12692
rect 78330 12648 78390 12910
rect 78716 12864 78776 13000
rect 79730 13000 79748 13060
rect 79782 13060 79788 13576
rect 80752 13576 80812 13732
rect 81262 13666 81322 13732
rect 82278 13732 82850 13792
rect 82278 13666 82338 13732
rect 81048 13660 81536 13666
rect 81048 13626 81060 13660
rect 81524 13626 81536 13660
rect 81048 13620 81536 13626
rect 82066 13660 82554 13666
rect 82066 13626 82078 13660
rect 82542 13626 82554 13660
rect 82066 13620 82554 13626
rect 80752 13536 80766 13576
rect 80760 13066 80766 13536
rect 79782 13000 79790 13060
rect 79012 12950 79500 12956
rect 79012 12916 79024 12950
rect 79488 12916 79500 12950
rect 79012 12910 79500 12916
rect 78522 12804 78776 12864
rect 78324 12588 78330 12648
rect 78390 12588 78396 12648
rect 78522 12538 78582 12804
rect 78712 12692 78718 12752
rect 78778 12692 78784 12752
rect 79220 12692 79226 12752
rect 79286 12692 79292 12752
rect 78522 12472 78582 12478
rect 77994 12428 78482 12434
rect 77994 12394 78006 12428
rect 78470 12394 78482 12428
rect 77994 12388 78482 12394
rect 78718 12344 78778 12692
rect 79226 12434 79286 12692
rect 79372 12648 79432 12910
rect 79730 12862 79790 13000
rect 80756 13000 80766 13066
rect 80800 13536 80812 13576
rect 81778 13576 81824 13588
rect 80800 13066 80806 13536
rect 80800 13000 80816 13066
rect 81778 13050 81784 13576
rect 80030 12950 80518 12956
rect 80030 12916 80042 12950
rect 80506 12916 80518 12950
rect 80030 12910 80518 12916
rect 79724 12802 79730 12862
rect 79790 12802 79796 12862
rect 79366 12588 79372 12648
rect 79432 12588 79438 12648
rect 79012 12428 79500 12434
rect 79012 12394 79024 12428
rect 79488 12394 79500 12428
rect 79012 12388 79500 12394
rect 79730 12344 79790 12802
rect 80234 12752 80294 12910
rect 80756 12752 80816 13000
rect 81768 13000 81784 13050
rect 81818 13050 81824 13576
rect 82790 13576 82850 13732
rect 83084 13660 83572 13666
rect 83084 13626 83096 13660
rect 83560 13626 83572 13660
rect 83084 13620 83572 13626
rect 84102 13660 84590 13666
rect 84102 13626 84114 13660
rect 84578 13626 84590 13660
rect 84102 13620 84590 13626
rect 82790 13550 82802 13576
rect 82796 13056 82802 13550
rect 81818 13000 81828 13050
rect 82788 13000 82802 13056
rect 82836 13550 82850 13576
rect 83814 13576 83860 13588
rect 82836 13056 82842 13550
rect 82836 13054 82848 13056
rect 82836 13000 82850 13054
rect 83814 13036 83820 13576
rect 81246 12956 81306 12958
rect 81048 12950 81536 12956
rect 81048 12916 81060 12950
rect 81524 12916 81536 12950
rect 81048 12910 81536 12916
rect 81246 12752 81306 12910
rect 81768 12862 81828 13000
rect 82278 12956 82338 12958
rect 82066 12950 82554 12956
rect 82066 12916 82078 12950
rect 82542 12916 82554 12950
rect 82066 12910 82554 12916
rect 81762 12802 81768 12862
rect 81828 12802 81834 12862
rect 80228 12692 80234 12752
rect 80294 12692 80300 12752
rect 80750 12692 80756 12752
rect 80816 12692 80822 12752
rect 81240 12692 81246 12752
rect 81306 12692 81312 12752
rect 80234 12434 80294 12692
rect 80750 12480 80756 12540
rect 80816 12480 80822 12540
rect 80030 12428 80518 12434
rect 80030 12394 80042 12428
rect 80506 12394 80518 12428
rect 80030 12388 80518 12394
rect 76728 12292 76738 12300
rect 77694 12296 77712 12344
rect 76728 11816 76734 12292
rect 77706 11816 77712 12296
rect 76728 11768 76740 11816
rect 75958 11718 76446 11724
rect 75958 11684 75970 11718
rect 76434 11684 76446 11718
rect 75958 11678 76446 11684
rect 76162 11618 76222 11678
rect 76680 11618 76740 11768
rect 77700 11768 77712 11816
rect 77746 12296 77754 12344
rect 78714 12304 78730 12344
rect 77746 11816 77752 12296
rect 77746 11768 77760 11816
rect 78724 11786 78730 12304
rect 76976 11718 77464 11724
rect 76976 11684 76988 11718
rect 77452 11684 77464 11718
rect 76976 11678 77464 11684
rect 77182 11618 77242 11678
rect 76162 11558 77242 11618
rect 77700 11546 77760 11768
rect 78718 11768 78730 11786
rect 78764 12306 78780 12344
rect 78764 12304 78778 12306
rect 78764 11786 78770 12304
rect 79730 12298 79748 12344
rect 79742 11822 79748 12298
rect 78764 11768 78778 11786
rect 77994 11718 78482 11724
rect 77994 11684 78006 11718
rect 78470 11684 78482 11718
rect 77994 11678 78482 11684
rect 78206 11622 78266 11678
rect 78718 11622 78778 11768
rect 79730 11768 79748 11822
rect 79782 12298 79790 12344
rect 80756 12344 80816 12480
rect 81246 12434 81306 12692
rect 81048 12428 81536 12434
rect 81048 12394 81060 12428
rect 81524 12394 81536 12428
rect 81048 12388 81536 12394
rect 80756 12302 80766 12344
rect 79782 11822 79788 12298
rect 79782 11768 79790 11822
rect 79012 11718 79500 11724
rect 79012 11684 79024 11718
rect 79488 11684 79500 11718
rect 79012 11678 79500 11684
rect 79208 11622 79268 11678
rect 78206 11562 79268 11622
rect 79730 11546 79790 11768
rect 80760 11768 80766 12302
rect 80800 12302 80816 12344
rect 81768 12344 81828 12802
rect 82278 12752 82338 12910
rect 82790 12752 82850 13000
rect 83806 13000 83820 13036
rect 83854 13036 83860 13576
rect 84824 13576 84884 13934
rect 85328 13666 85388 14144
rect 85844 14092 85904 14234
rect 86862 14234 86874 14810
rect 86908 14234 86922 14810
rect 87886 14810 87932 14822
rect 87886 14288 87892 14810
rect 86138 14184 86626 14190
rect 86138 14150 86150 14184
rect 86614 14150 86626 14184
rect 86138 14144 86626 14150
rect 85838 14032 85844 14092
rect 85904 14032 85910 14092
rect 85120 13660 85608 13666
rect 85120 13626 85132 13660
rect 85596 13626 85608 13660
rect 85120 13620 85608 13626
rect 84824 13536 84838 13576
rect 83854 13000 83866 13036
rect 83084 12950 83572 12956
rect 83084 12916 83096 12950
rect 83560 12916 83572 12950
rect 83084 12910 83572 12916
rect 83292 12862 83352 12910
rect 83806 12862 83866 13000
rect 84832 13000 84838 13536
rect 84872 13536 84884 13576
rect 85844 13576 85904 14032
rect 86354 13666 86414 14144
rect 86862 13994 86922 14234
rect 87874 14234 87892 14288
rect 87926 14288 87932 14810
rect 89766 14470 89878 15256
rect 87926 14234 87934 14288
rect 87156 14184 87644 14190
rect 87156 14150 87168 14184
rect 87632 14150 87644 14184
rect 87156 14144 87644 14150
rect 86856 13934 86862 13994
rect 86922 13934 86928 13994
rect 86138 13660 86626 13666
rect 86138 13626 86150 13660
rect 86614 13626 86626 13660
rect 86138 13620 86626 13626
rect 85844 13544 85856 13576
rect 84872 13000 84878 13536
rect 84832 12988 84878 13000
rect 85850 13000 85856 13544
rect 85890 13544 85904 13576
rect 86862 13576 86922 13934
rect 87376 13666 87436 14144
rect 87874 14092 87934 14234
rect 87868 14032 87874 14092
rect 87934 14032 87940 14092
rect 87156 13660 87644 13666
rect 87156 13626 87168 13660
rect 87632 13626 87644 13660
rect 87156 13620 87644 13626
rect 86862 13548 86874 13576
rect 85890 13000 85896 13544
rect 85850 12988 85896 13000
rect 86868 13000 86874 13548
rect 86908 13548 86922 13576
rect 87874 13576 87934 14032
rect 88592 13934 88598 13994
rect 88658 13934 88664 13994
rect 87874 13550 87892 13576
rect 86908 13000 86914 13548
rect 86868 12988 86914 13000
rect 87886 13000 87892 13550
rect 87926 13550 87934 13576
rect 87926 13000 87932 13550
rect 87886 12988 87932 13000
rect 84102 12950 84590 12956
rect 84102 12916 84114 12950
rect 84578 12916 84590 12950
rect 84102 12910 84590 12916
rect 85120 12950 85608 12956
rect 85120 12916 85132 12950
rect 85596 12916 85608 12950
rect 85120 12910 85608 12916
rect 86138 12950 86626 12956
rect 86138 12916 86150 12950
rect 86614 12916 86626 12950
rect 86138 12910 86626 12916
rect 87156 12950 87644 12956
rect 87156 12916 87168 12950
rect 87632 12916 87644 12950
rect 87156 12910 87644 12916
rect 84314 12862 84374 12910
rect 83800 12802 83806 12862
rect 83866 12802 83872 12862
rect 84308 12802 84314 12862
rect 84374 12802 84380 12862
rect 83292 12796 83352 12802
rect 82272 12692 82278 12752
rect 82338 12692 82344 12752
rect 82784 12692 82790 12752
rect 82850 12692 82856 12752
rect 82258 12588 82264 12648
rect 82324 12588 82330 12648
rect 83296 12588 83302 12648
rect 83362 12588 83368 12648
rect 82264 12434 82324 12588
rect 82782 12480 82788 12540
rect 82848 12480 82854 12540
rect 82066 12428 82554 12434
rect 82066 12394 82078 12428
rect 82542 12394 82554 12428
rect 82066 12388 82554 12394
rect 80800 11768 80806 12302
rect 80760 11756 80806 11768
rect 81768 11768 81784 12344
rect 81818 11768 81828 12344
rect 82788 12344 82848 12480
rect 83302 12434 83362 12588
rect 83084 12428 83572 12434
rect 83084 12394 83096 12428
rect 83560 12394 83572 12428
rect 83084 12388 83572 12394
rect 82788 12302 82802 12344
rect 80030 11718 80518 11724
rect 80030 11684 80042 11718
rect 80506 11684 80518 11718
rect 80030 11678 80518 11684
rect 81048 11718 81536 11724
rect 81048 11684 81060 11718
rect 81524 11684 81536 11718
rect 81048 11678 81536 11684
rect 80254 11576 81316 11636
rect 73620 11486 73626 11546
rect 73686 11486 73692 11546
rect 75656 11486 75662 11546
rect 75722 11486 75728 11546
rect 77694 11486 77700 11546
rect 77760 11486 77766 11546
rect 79724 11486 79730 11546
rect 79790 11486 79796 11546
rect 74640 11364 74646 11424
rect 74706 11364 74712 11424
rect 76674 11364 76680 11424
rect 76740 11364 76746 11424
rect 78704 11364 78710 11424
rect 78770 11364 78776 11424
rect 72902 11194 73390 11200
rect 72902 11160 72914 11194
rect 73378 11160 73390 11194
rect 72902 11154 73390 11160
rect 73920 11194 74408 11200
rect 73920 11160 73932 11194
rect 74396 11160 74408 11194
rect 73920 11154 74408 11160
rect 71636 10534 71642 11080
rect 72604 11066 72620 11110
rect 72614 10584 72620 11066
rect 71596 10522 71642 10534
rect 72606 10534 72620 10584
rect 72654 11066 72664 11110
rect 73632 11110 73678 11122
rect 72654 10584 72660 11066
rect 72654 10534 72666 10584
rect 73632 10570 73638 11110
rect 70866 10484 71354 10490
rect 70866 10450 70878 10484
rect 71342 10450 71354 10484
rect 70866 10444 71354 10450
rect 71884 10484 72372 10490
rect 71884 10450 71896 10484
rect 72360 10450 72372 10484
rect 71884 10444 72372 10450
rect 70564 10346 70570 10406
rect 70630 10346 70636 10406
rect 70060 10128 70066 10188
rect 70126 10128 70132 10188
rect 70066 9966 70126 10128
rect 69848 9960 70336 9966
rect 69848 9926 69860 9960
rect 70324 9926 70336 9960
rect 69848 9920 70336 9926
rect 68582 9300 68588 9840
rect 69552 9834 69566 9876
rect 69560 9358 69566 9834
rect 68542 9288 68588 9300
rect 69554 9300 69566 9358
rect 69600 9834 69612 9876
rect 70570 9876 70630 10346
rect 71068 10194 71128 10444
rect 71586 10242 71592 10302
rect 71652 10242 71658 10302
rect 71068 10188 71130 10194
rect 71068 10128 71070 10188
rect 71068 10122 71130 10128
rect 71068 9966 71128 10122
rect 70866 9960 71354 9966
rect 70866 9926 70878 9960
rect 71342 9926 71354 9960
rect 70866 9920 71354 9926
rect 69600 9358 69606 9834
rect 70570 9832 70584 9876
rect 69600 9300 69614 9358
rect 70578 9348 70584 9832
rect 67812 9250 68300 9256
rect 67812 9216 67824 9250
rect 68288 9216 68300 9250
rect 67812 9210 68300 9216
rect 68830 9250 69318 9256
rect 68830 9216 68842 9250
rect 69306 9216 69318 9250
rect 68830 9210 69318 9216
rect 68528 9090 68534 9150
rect 68594 9090 68600 9150
rect 67812 8728 68300 8734
rect 67812 8694 67824 8728
rect 68288 8694 68300 8728
rect 67812 8688 68300 8694
rect 67524 8644 67570 8656
rect 67524 8114 67530 8644
rect 67514 8068 67530 8114
rect 67564 8114 67570 8644
rect 68534 8644 68594 9090
rect 69040 9048 69100 9210
rect 69034 8988 69040 9048
rect 69100 8988 69106 9048
rect 69554 8846 69614 9300
rect 70572 9300 70584 9348
rect 70618 9832 70630 9876
rect 71592 9876 71652 10242
rect 72084 10194 72144 10444
rect 72606 10406 72666 10534
rect 73624 10534 73638 10570
rect 73672 10570 73678 11110
rect 74646 11110 74706 11364
rect 74938 11194 75426 11200
rect 74938 11160 74950 11194
rect 75414 11160 75426 11194
rect 74938 11154 75426 11160
rect 75956 11194 76444 11200
rect 75956 11160 75968 11194
rect 76432 11160 76444 11194
rect 75956 11154 76444 11160
rect 74646 11054 74656 11110
rect 73672 10534 73684 10570
rect 72902 10484 73390 10490
rect 72902 10450 72914 10484
rect 73378 10450 73390 10484
rect 72902 10444 73390 10450
rect 72600 10346 72606 10406
rect 72666 10346 72672 10406
rect 72082 10188 72144 10194
rect 72142 10128 72144 10188
rect 72082 10122 72144 10128
rect 72084 9966 72144 10122
rect 71884 9960 72372 9966
rect 71884 9926 71896 9960
rect 72360 9926 72372 9960
rect 71884 9920 72372 9926
rect 71592 9834 71602 9876
rect 70618 9348 70624 9832
rect 70618 9300 70632 9348
rect 69848 9250 70336 9256
rect 69848 9216 69860 9250
rect 70324 9216 70336 9250
rect 69848 9210 70336 9216
rect 70572 9150 70632 9300
rect 71596 9300 71602 9834
rect 71636 9834 71652 9876
rect 72606 9876 72666 10346
rect 73102 10188 73162 10444
rect 73624 10302 73684 10534
rect 74650 10534 74656 11054
rect 74690 11054 74706 11110
rect 75668 11110 75714 11122
rect 74690 10534 74696 11054
rect 75668 10564 75674 11110
rect 74650 10522 74696 10534
rect 75658 10534 75674 10564
rect 75708 10564 75714 11110
rect 76680 11110 76740 11364
rect 76974 11194 77462 11200
rect 76974 11160 76986 11194
rect 77450 11160 77462 11194
rect 76974 11154 77462 11160
rect 77992 11194 78480 11200
rect 77992 11160 78004 11194
rect 78468 11160 78480 11194
rect 77992 11154 78480 11160
rect 76680 11060 76692 11110
rect 75708 10534 75718 10564
rect 73920 10484 74408 10490
rect 73920 10450 73932 10484
rect 74396 10450 74408 10484
rect 73920 10444 74408 10450
rect 74938 10484 75426 10490
rect 74938 10450 74950 10484
rect 75414 10450 75426 10484
rect 74938 10444 75426 10450
rect 73618 10242 73624 10302
rect 73684 10242 73690 10302
rect 74114 10246 74174 10444
rect 75156 10246 75216 10444
rect 75658 10302 75718 10534
rect 76686 10534 76692 11060
rect 76726 11060 76740 11110
rect 77704 11110 77750 11122
rect 76726 10534 76732 11060
rect 77704 10576 77710 11110
rect 76686 10522 76732 10534
rect 77698 10534 77710 10576
rect 77744 10576 77750 11110
rect 78710 11110 78770 11364
rect 80254 11200 80314 11576
rect 80744 11486 80750 11546
rect 80810 11486 80816 11546
rect 79010 11194 79498 11200
rect 79010 11160 79022 11194
rect 79486 11160 79498 11194
rect 79010 11154 79498 11160
rect 80028 11194 80516 11200
rect 80028 11160 80040 11194
rect 80504 11160 80516 11194
rect 80028 11154 80516 11160
rect 78710 11066 78728 11110
rect 77744 10534 77758 10576
rect 75956 10484 76444 10490
rect 75956 10450 75968 10484
rect 76432 10450 76444 10484
rect 75956 10444 76444 10450
rect 76974 10484 77462 10490
rect 76974 10450 76986 10484
rect 77450 10450 77462 10484
rect 76974 10444 77462 10450
rect 73618 10130 73624 10190
rect 73684 10130 73690 10190
rect 74114 10186 75216 10246
rect 75652 10242 75658 10302
rect 75718 10242 75724 10302
rect 73102 9966 73162 10128
rect 72902 9960 73390 9966
rect 72902 9926 72914 9960
rect 73378 9926 73390 9960
rect 72902 9920 73390 9926
rect 71636 9300 71642 9834
rect 72606 9828 72620 9876
rect 72614 9350 72620 9828
rect 71596 9288 71642 9300
rect 72608 9300 72620 9350
rect 72654 9828 72666 9876
rect 73624 9876 73684 10130
rect 74114 9966 74174 10186
rect 74636 10020 74642 10080
rect 74702 10020 74708 10080
rect 73920 9960 74408 9966
rect 73920 9926 73932 9960
rect 74396 9926 74408 9960
rect 73920 9920 74408 9926
rect 72654 9350 72660 9828
rect 73624 9818 73638 9876
rect 72654 9300 72668 9350
rect 70866 9250 71354 9256
rect 70866 9216 70878 9250
rect 71342 9216 71354 9250
rect 70866 9210 71354 9216
rect 71884 9250 72372 9256
rect 71884 9216 71896 9250
rect 72360 9216 72372 9250
rect 71884 9210 72372 9216
rect 70566 9090 70572 9150
rect 70632 9090 70638 9150
rect 70564 8886 70570 8946
rect 70630 8886 70636 8946
rect 71078 8940 71138 9210
rect 72100 8940 72160 9210
rect 72608 9150 72668 9300
rect 73632 9300 73638 9818
rect 73672 9818 73684 9876
rect 74642 9876 74702 10020
rect 75156 9966 75216 10186
rect 75654 10130 75660 10190
rect 75720 10130 75726 10190
rect 74938 9960 75426 9966
rect 74938 9926 74950 9960
rect 75414 9926 75426 9960
rect 74938 9920 75426 9926
rect 74642 9830 74656 9876
rect 73672 9300 73678 9818
rect 73632 9288 73678 9300
rect 74650 9300 74656 9830
rect 74690 9830 74702 9876
rect 75660 9876 75720 10130
rect 76156 9966 76216 10444
rect 76670 10020 76676 10080
rect 76736 10020 76742 10080
rect 75956 9960 76444 9966
rect 75956 9926 75968 9960
rect 76432 9926 76444 9960
rect 75956 9920 76444 9926
rect 74690 9300 74696 9830
rect 75660 9808 75674 9876
rect 74650 9288 74696 9300
rect 75668 9300 75674 9808
rect 75708 9808 75720 9876
rect 76676 9876 76736 10020
rect 77190 9966 77250 10444
rect 77698 10302 77758 10534
rect 78722 10534 78728 11066
rect 78762 11066 78770 11110
rect 79740 11110 79786 11122
rect 78762 10534 78768 11066
rect 79740 10586 79746 11110
rect 78722 10522 78768 10534
rect 79732 10534 79746 10586
rect 79780 10586 79786 11110
rect 80750 11110 80810 11486
rect 81256 11370 81316 11576
rect 81768 11546 81828 11768
rect 82796 11768 82802 12302
rect 82836 12302 82848 12344
rect 83806 12344 83866 12802
rect 85328 12692 85334 12752
rect 85394 12692 85400 12752
rect 86348 12692 86354 12752
rect 86414 12692 86420 12752
rect 84296 12588 84302 12648
rect 84362 12588 84368 12648
rect 84302 12434 84362 12588
rect 84814 12480 84820 12540
rect 84880 12480 84886 12540
rect 84102 12428 84590 12434
rect 84102 12394 84114 12428
rect 84578 12394 84590 12428
rect 84102 12388 84590 12394
rect 84302 12376 84362 12388
rect 82836 11768 82842 12302
rect 83806 12286 83820 12344
rect 83814 11816 83820 12286
rect 82796 11756 82842 11768
rect 83804 11768 83820 11816
rect 83854 12286 83866 12344
rect 84820 12344 84880 12480
rect 85334 12434 85394 12692
rect 86354 12434 86414 12692
rect 86856 12480 86862 12540
rect 86922 12480 86928 12540
rect 87360 12480 87366 12540
rect 87426 12480 87432 12540
rect 87870 12480 87876 12540
rect 87936 12480 87942 12540
rect 85120 12428 85608 12434
rect 85120 12394 85132 12428
rect 85596 12394 85608 12428
rect 85120 12388 85608 12394
rect 86138 12428 86626 12434
rect 86138 12394 86150 12428
rect 86614 12394 86626 12428
rect 86138 12388 86626 12394
rect 84820 12298 84838 12344
rect 83854 11816 83860 12286
rect 83854 11768 83864 11816
rect 82066 11718 82554 11724
rect 82066 11684 82078 11718
rect 82542 11684 82554 11718
rect 82066 11678 82554 11684
rect 83084 11718 83572 11724
rect 83084 11684 83096 11718
rect 83560 11684 83572 11718
rect 83084 11678 83572 11684
rect 82268 11650 82328 11678
rect 83302 11650 83362 11678
rect 82260 11590 82266 11650
rect 82326 11590 82332 11650
rect 83296 11590 83302 11650
rect 83362 11590 83368 11650
rect 81762 11486 81768 11546
rect 81828 11486 81834 11546
rect 82268 11370 82328 11590
rect 82782 11486 82788 11546
rect 82848 11486 82854 11546
rect 81256 11310 82328 11370
rect 81256 11200 81316 11310
rect 82268 11200 82328 11310
rect 81046 11194 81534 11200
rect 81046 11160 81058 11194
rect 81522 11160 81534 11194
rect 81046 11154 81534 11160
rect 82064 11194 82552 11200
rect 82064 11160 82076 11194
rect 82540 11160 82552 11194
rect 82064 11154 82552 11160
rect 80750 11062 80764 11110
rect 79780 10534 79792 10586
rect 80758 10566 80764 11062
rect 77992 10484 78480 10490
rect 77992 10450 78004 10484
rect 78468 10450 78480 10484
rect 77992 10444 78480 10450
rect 79010 10484 79498 10490
rect 79010 10450 79022 10484
rect 79486 10450 79498 10484
rect 79010 10444 79498 10450
rect 77692 10242 77698 10302
rect 77758 10242 77764 10302
rect 78212 10246 78272 10444
rect 79220 10246 79280 10444
rect 79732 10302 79792 10534
rect 80750 10534 80764 10566
rect 80798 11062 80810 11110
rect 81776 11110 81822 11122
rect 80798 10566 80804 11062
rect 81776 10570 81782 11110
rect 80798 10534 80810 10566
rect 80028 10484 80516 10490
rect 80028 10450 80040 10484
rect 80504 10450 80516 10484
rect 80028 10444 80516 10450
rect 77690 10130 77696 10190
rect 77756 10130 77762 10190
rect 78212 10186 79280 10246
rect 79726 10242 79732 10302
rect 79792 10242 79798 10302
rect 79922 10238 79928 10298
rect 79988 10238 79994 10298
rect 76974 9960 77462 9966
rect 76974 9926 76986 9960
rect 77450 9926 77462 9960
rect 76974 9920 77462 9926
rect 76676 9828 76692 9876
rect 75708 9300 75714 9808
rect 75668 9288 75714 9300
rect 76686 9300 76692 9828
rect 76726 9828 76736 9876
rect 77696 9876 77756 10130
rect 78212 9966 78272 10186
rect 78710 10020 78716 10080
rect 78776 10020 78782 10080
rect 77992 9960 78480 9966
rect 77992 9926 78004 9960
rect 78468 9926 78480 9960
rect 77992 9920 78480 9926
rect 76726 9300 76732 9828
rect 77696 9826 77710 9876
rect 76686 9288 76732 9300
rect 77704 9300 77710 9826
rect 77744 9826 77756 9876
rect 78716 9876 78776 10020
rect 79220 9966 79280 10186
rect 79726 10130 79732 10190
rect 79792 10130 79798 10190
rect 79010 9960 79498 9966
rect 79010 9926 79022 9960
rect 79486 9926 79498 9960
rect 79010 9920 79498 9926
rect 78716 9838 78728 9876
rect 77744 9300 77750 9826
rect 78722 9346 78728 9838
rect 77704 9288 77750 9300
rect 78716 9300 78728 9346
rect 78762 9838 78776 9876
rect 79732 9876 79792 10130
rect 79928 10080 79988 10238
rect 80222 10082 80282 10444
rect 80750 10406 80810 10534
rect 81766 10534 81782 10570
rect 81816 10570 81822 11110
rect 82788 11110 82848 11486
rect 83302 11362 83362 11590
rect 83804 11546 83864 11768
rect 84832 11768 84838 12298
rect 84872 12298 84880 12344
rect 85850 12344 85896 12356
rect 84872 11768 84878 12298
rect 85850 11826 85856 12344
rect 84832 11756 84878 11768
rect 85840 11768 85856 11826
rect 85890 11826 85896 12344
rect 86862 12344 86922 12480
rect 87366 12434 87426 12480
rect 87156 12428 87644 12434
rect 87156 12394 87168 12428
rect 87632 12394 87644 12428
rect 87156 12388 87644 12394
rect 86862 12288 86874 12344
rect 85890 11768 85900 11826
rect 84102 11718 84590 11724
rect 84102 11684 84114 11718
rect 84578 11684 84590 11718
rect 84102 11678 84590 11684
rect 85120 11718 85608 11724
rect 85120 11684 85132 11718
rect 85596 11684 85608 11718
rect 85120 11678 85608 11684
rect 84318 11650 84378 11678
rect 84312 11590 84318 11650
rect 84378 11590 84384 11650
rect 85840 11546 85900 11768
rect 86868 11768 86874 12288
rect 86908 12288 86922 12344
rect 87876 12344 87936 12480
rect 87876 12308 87892 12344
rect 86908 11768 86914 12288
rect 86868 11756 86914 11768
rect 87886 11768 87892 12308
rect 87926 12308 87936 12344
rect 87926 11768 87932 12308
rect 87886 11756 87932 11768
rect 86138 11718 86626 11724
rect 86138 11684 86150 11718
rect 86614 11684 86626 11718
rect 86138 11678 86626 11684
rect 87156 11718 87644 11724
rect 87156 11684 87168 11718
rect 87632 11684 87644 11718
rect 87156 11678 87644 11684
rect 83798 11486 83804 11546
rect 83864 11486 83870 11546
rect 85834 11486 85840 11546
rect 85900 11486 85906 11546
rect 83302 11302 86390 11362
rect 83302 11200 83362 11302
rect 86330 11200 86390 11302
rect 87368 11276 87936 11336
rect 87368 11200 87428 11276
rect 83082 11194 83570 11200
rect 83082 11160 83094 11194
rect 83558 11160 83570 11194
rect 83082 11154 83570 11160
rect 84100 11194 84588 11200
rect 84100 11160 84112 11194
rect 84576 11160 84588 11194
rect 84100 11154 84588 11160
rect 85118 11194 85606 11200
rect 85118 11160 85130 11194
rect 85594 11160 85606 11194
rect 85118 11154 85606 11160
rect 86136 11194 86624 11200
rect 86136 11160 86148 11194
rect 86612 11160 86624 11194
rect 86136 11154 86624 11160
rect 87154 11194 87642 11200
rect 87154 11160 87166 11194
rect 87630 11160 87642 11194
rect 87154 11154 87642 11160
rect 82788 11052 82800 11110
rect 82794 10580 82800 11052
rect 81816 10534 81826 10570
rect 81046 10484 81534 10490
rect 81046 10450 81058 10484
rect 81522 10450 81534 10484
rect 81046 10444 81534 10450
rect 80744 10346 80750 10406
rect 80810 10346 80816 10406
rect 79922 10020 79928 10080
rect 79988 10020 79994 10080
rect 80216 10022 80222 10082
rect 80282 10022 80288 10082
rect 80222 9966 80282 10022
rect 80028 9960 80516 9966
rect 80028 9926 80040 9960
rect 80504 9926 80516 9960
rect 80028 9920 80516 9926
rect 78762 9346 78768 9838
rect 79732 9832 79746 9876
rect 78762 9300 78776 9346
rect 72902 9250 73390 9256
rect 72902 9216 72914 9250
rect 73378 9216 73390 9250
rect 72902 9210 73390 9216
rect 73920 9250 74408 9256
rect 73920 9216 73932 9250
rect 74396 9216 74408 9250
rect 73920 9210 74408 9216
rect 74938 9250 75426 9256
rect 74938 9216 74950 9250
rect 75414 9216 75426 9250
rect 74938 9210 75426 9216
rect 75956 9250 76444 9256
rect 75956 9216 75968 9250
rect 76432 9216 76444 9250
rect 75956 9210 76444 9216
rect 76974 9250 77462 9256
rect 76974 9216 76986 9250
rect 77450 9216 77462 9250
rect 76974 9210 77462 9216
rect 77992 9250 78480 9256
rect 77992 9216 78004 9250
rect 78468 9216 78480 9250
rect 77992 9210 78480 9216
rect 72602 9090 72608 9150
rect 72668 9090 72674 9150
rect 69548 8786 69554 8846
rect 69614 8786 69620 8846
rect 68830 8728 69318 8734
rect 68830 8694 68842 8728
rect 69306 8694 69318 8728
rect 68830 8688 69318 8694
rect 68534 8606 68548 8644
rect 67564 8068 67574 8114
rect 68542 8110 68548 8606
rect 67514 7906 67574 8068
rect 68532 8068 68548 8110
rect 68582 8606 68594 8644
rect 69554 8644 69614 8786
rect 69848 8728 70336 8734
rect 69848 8694 69860 8728
rect 70324 8694 70336 8728
rect 69848 8688 70336 8694
rect 68582 8110 68588 8606
rect 69554 8604 69566 8644
rect 68582 8068 68592 8110
rect 67812 8018 68300 8024
rect 67812 7984 67824 8018
rect 68288 7984 68300 8018
rect 67812 7978 68300 7984
rect 68026 7906 68086 7978
rect 68532 7906 68592 8068
rect 69560 8068 69566 8604
rect 69600 8604 69614 8644
rect 70570 8644 70630 8886
rect 71072 8880 71078 8940
rect 71138 8880 71144 8940
rect 72094 8880 72100 8940
rect 72160 8880 72166 8940
rect 71582 8786 71588 8846
rect 71648 8786 71654 8846
rect 70866 8728 71354 8734
rect 70866 8694 70878 8728
rect 71342 8694 71354 8728
rect 70866 8688 71354 8694
rect 69600 8068 69606 8604
rect 70570 8592 70584 8644
rect 69560 8056 69606 8068
rect 70578 8068 70584 8592
rect 70618 8592 70630 8644
rect 71588 8644 71648 8786
rect 72100 8734 72160 8880
rect 71884 8728 72372 8734
rect 71884 8694 71896 8728
rect 72360 8694 72372 8728
rect 71884 8688 72372 8694
rect 71588 8600 71602 8644
rect 70618 8068 70624 8592
rect 71596 8104 71602 8600
rect 70578 8056 70624 8068
rect 71588 8068 71602 8104
rect 71636 8600 71648 8644
rect 72608 8644 72668 9090
rect 73114 8940 73174 9210
rect 74132 9048 74192 9210
rect 75152 9160 75212 9210
rect 76152 9160 76212 9210
rect 77190 9160 77250 9210
rect 78218 9160 78278 9210
rect 74634 9090 74640 9150
rect 74700 9090 74706 9150
rect 75152 9100 78278 9160
rect 74126 8988 74132 9048
rect 74192 8988 74198 9048
rect 73108 8880 73114 8940
rect 73174 8880 73180 8940
rect 74126 8880 74132 8940
rect 74192 8880 74198 8940
rect 73114 8734 73174 8880
rect 73618 8786 73624 8846
rect 73684 8786 73690 8846
rect 72902 8728 73390 8734
rect 72902 8694 72914 8728
rect 73378 8694 73390 8728
rect 72902 8688 73390 8694
rect 71636 8104 71642 8600
rect 71636 8068 71648 8104
rect 68830 8018 69318 8024
rect 68830 7984 68842 8018
rect 69306 7984 69318 8018
rect 68830 7978 69318 7984
rect 69848 8018 70336 8024
rect 69848 7984 69860 8018
rect 70324 7984 70336 8018
rect 69848 7978 70336 7984
rect 70866 8018 71354 8024
rect 70866 7984 70878 8018
rect 71342 7984 71354 8018
rect 70866 7978 71354 7984
rect 69036 7922 69096 7978
rect 67514 7846 68592 7906
rect 69030 7862 69036 7922
rect 69096 7862 69102 7922
rect 69940 7862 69946 7922
rect 70006 7862 70012 7922
rect 69030 7646 69036 7706
rect 69096 7646 69102 7706
rect 69036 7640 69098 7646
rect 67398 7602 67460 7608
rect 67398 7542 67400 7602
rect 67398 7536 67460 7542
rect 67280 6284 67286 6344
rect 67346 6284 67352 6344
rect 67180 5280 67244 5286
rect 67180 5228 67192 5280
rect 67180 5222 67244 5228
rect 67180 4100 67240 5222
rect 67286 4226 67346 6284
rect 67398 5358 67458 7536
rect 69038 7500 69098 7640
rect 69946 7500 70006 7862
rect 70074 7706 70134 7978
rect 70942 7862 70948 7922
rect 71008 7862 71014 7922
rect 70074 7640 70134 7646
rect 70948 7500 71008 7862
rect 71088 7706 71148 7978
rect 71588 7820 71648 8068
rect 72608 8068 72620 8644
rect 72654 8068 72668 8644
rect 73624 8644 73684 8786
rect 74132 8734 74192 8880
rect 73920 8728 74408 8734
rect 73920 8694 73932 8728
rect 74396 8694 74408 8728
rect 73920 8688 74408 8694
rect 73624 8608 73638 8644
rect 71884 8018 72372 8024
rect 71884 7984 71896 8018
rect 72360 7984 72372 8018
rect 71884 7978 72372 7984
rect 72100 7922 72160 7978
rect 72094 7862 72100 7922
rect 72160 7862 72166 7922
rect 71582 7760 71588 7820
rect 71648 7760 71654 7820
rect 71082 7646 71088 7706
rect 71148 7646 71154 7706
rect 72100 7500 72160 7862
rect 67812 7494 68300 7500
rect 67812 7460 67824 7494
rect 68288 7460 68300 7494
rect 67812 7454 68300 7460
rect 68830 7494 69318 7500
rect 68830 7460 68842 7494
rect 69306 7460 69318 7494
rect 68830 7454 69318 7460
rect 69848 7494 70336 7500
rect 69848 7460 69860 7494
rect 70324 7460 70336 7494
rect 69848 7454 70336 7460
rect 70866 7494 71354 7500
rect 70866 7460 70878 7494
rect 71342 7460 71354 7494
rect 70866 7454 71354 7460
rect 71884 7494 72372 7500
rect 71884 7460 71896 7494
rect 72360 7460 72372 7494
rect 71884 7454 72372 7460
rect 67524 7410 67570 7422
rect 67524 6872 67530 7410
rect 67518 6834 67530 6872
rect 67564 6872 67570 7410
rect 68542 7410 68588 7422
rect 68542 6872 68548 7410
rect 67564 6834 67578 6872
rect 67518 6704 67578 6834
rect 68536 6834 68548 6872
rect 68582 6872 68588 7410
rect 69560 7410 69606 7422
rect 69560 6884 69566 7410
rect 68582 6834 68596 6872
rect 67812 6784 68300 6790
rect 67812 6750 67824 6784
rect 68288 6750 68300 6784
rect 67812 6744 68300 6750
rect 68016 6704 68076 6744
rect 68536 6704 68596 6834
rect 69552 6834 69566 6884
rect 69600 6884 69606 7410
rect 70578 7410 70624 7422
rect 70578 6892 70584 7410
rect 69600 6834 69612 6884
rect 68830 6784 69318 6790
rect 68830 6750 68842 6784
rect 69306 6750 69318 6784
rect 68830 6744 69318 6750
rect 67518 6644 68596 6704
rect 68536 6590 68596 6644
rect 69028 6634 69034 6694
rect 69094 6634 69100 6694
rect 68530 6530 68536 6590
rect 68596 6530 68602 6590
rect 68526 6320 68532 6380
rect 68592 6320 68598 6380
rect 67812 6260 68300 6266
rect 67812 6226 67824 6260
rect 68288 6226 68300 6260
rect 67812 6220 68300 6226
rect 67524 6176 67570 6188
rect 67524 5634 67530 6176
rect 67514 5600 67530 5634
rect 67564 5634 67570 6176
rect 68532 6176 68592 6320
rect 69034 6266 69094 6634
rect 69552 6478 69612 6834
rect 70570 6834 70584 6892
rect 70618 6892 70624 7410
rect 71596 7410 71642 7422
rect 70618 6834 70630 6892
rect 71596 6880 71602 7410
rect 69848 6784 70336 6790
rect 69848 6750 69860 6784
rect 70324 6750 70336 6784
rect 69848 6744 70336 6750
rect 70042 6694 70102 6744
rect 70036 6634 70042 6694
rect 70102 6634 70108 6694
rect 69546 6418 69552 6478
rect 69612 6418 69618 6478
rect 70570 6380 70630 6834
rect 71590 6834 71602 6880
rect 71636 6880 71642 7410
rect 72608 7410 72668 8068
rect 73632 8068 73638 8608
rect 73672 8608 73684 8644
rect 74640 8644 74700 9090
rect 75146 8880 75152 8940
rect 75212 8880 75218 8940
rect 78218 8924 78278 9100
rect 78716 9034 78776 9300
rect 79740 9300 79746 9832
rect 79780 9832 79792 9876
rect 80750 9876 80810 10346
rect 81252 10088 81312 10444
rect 81766 10190 81826 10534
rect 82786 10534 82800 10580
rect 82834 11052 82848 11110
rect 83812 11110 83858 11122
rect 82834 10580 82840 11052
rect 83812 10590 83818 11110
rect 82834 10534 82846 10580
rect 82064 10484 82552 10490
rect 82064 10450 82076 10484
rect 82540 10450 82552 10484
rect 82064 10444 82552 10450
rect 81760 10130 81766 10190
rect 81826 10130 81832 10190
rect 81250 10082 81312 10088
rect 81310 10022 81312 10082
rect 81250 10016 81312 10022
rect 81762 10016 81768 10076
rect 81828 10016 81834 10076
rect 81252 9966 81312 10016
rect 81046 9960 81534 9966
rect 81046 9926 81058 9960
rect 81522 9926 81534 9960
rect 81046 9920 81534 9926
rect 80750 9832 80764 9876
rect 79780 9300 79786 9832
rect 79740 9288 79786 9300
rect 80758 9300 80764 9832
rect 80798 9832 80810 9876
rect 81768 9876 81828 10016
rect 82276 9966 82336 10444
rect 82786 10406 82846 10534
rect 83804 10534 83818 10590
rect 83852 10590 83858 11110
rect 84830 11110 84876 11122
rect 83852 10534 83864 10590
rect 84830 10578 84836 11110
rect 83082 10484 83570 10490
rect 83082 10450 83094 10484
rect 83558 10450 83570 10484
rect 83082 10444 83570 10450
rect 82780 10346 82786 10406
rect 82846 10346 82852 10406
rect 82064 9960 82552 9966
rect 82064 9926 82076 9960
rect 82540 9926 82552 9960
rect 82064 9920 82552 9926
rect 81768 9846 81782 9876
rect 80798 9300 80804 9832
rect 81776 9340 81782 9846
rect 80758 9288 80804 9300
rect 81768 9300 81782 9340
rect 81816 9846 81828 9876
rect 82786 9876 82846 10346
rect 83302 9966 83362 10444
rect 83804 10190 83864 10534
rect 84820 10534 84836 10578
rect 84870 10578 84876 11110
rect 85848 11110 85894 11122
rect 85848 10578 85854 11110
rect 84870 10534 84880 10578
rect 84100 10484 84588 10490
rect 84100 10450 84112 10484
rect 84576 10450 84588 10484
rect 84100 10444 84588 10450
rect 83798 10130 83804 10190
rect 83864 10130 83870 10190
rect 84310 10140 84370 10444
rect 84820 10298 84880 10534
rect 85844 10534 85854 10578
rect 85888 10578 85894 11110
rect 86866 11110 86912 11122
rect 86866 10584 86872 11110
rect 85888 10534 85904 10578
rect 85118 10484 85606 10490
rect 85118 10450 85130 10484
rect 85594 10450 85606 10484
rect 85118 10444 85606 10450
rect 85326 10300 85386 10444
rect 84814 10238 84820 10298
rect 84880 10238 84886 10298
rect 85324 10294 85386 10300
rect 85384 10234 85386 10294
rect 85324 10228 85386 10234
rect 85326 10140 85386 10228
rect 85844 10190 85904 10534
rect 86860 10534 86872 10584
rect 86906 10584 86912 11110
rect 87876 11110 87936 11276
rect 87978 11252 87984 11312
rect 88044 11252 88050 11312
rect 87876 11082 87890 11110
rect 87884 10592 87890 11082
rect 86906 10534 86920 10584
rect 86136 10484 86624 10490
rect 86136 10450 86148 10484
rect 86612 10450 86624 10484
rect 86136 10444 86624 10450
rect 84310 10080 85386 10140
rect 85838 10130 85844 10190
rect 85904 10130 85910 10190
rect 83798 10016 83804 10076
rect 83864 10016 83870 10076
rect 83082 9960 83570 9966
rect 83082 9926 83094 9960
rect 83558 9926 83570 9960
rect 83082 9920 83570 9926
rect 81816 9340 81822 9846
rect 82786 9836 82800 9876
rect 81816 9300 81828 9340
rect 82794 9334 82800 9836
rect 79010 9250 79498 9256
rect 79010 9216 79022 9250
rect 79486 9216 79498 9250
rect 79010 9210 79498 9216
rect 80028 9250 80516 9256
rect 80028 9216 80040 9250
rect 80504 9216 80516 9250
rect 80028 9210 80516 9216
rect 81046 9250 81534 9256
rect 81046 9216 81058 9250
rect 81522 9216 81534 9250
rect 81046 9210 81534 9216
rect 79222 9162 79282 9210
rect 78710 8974 78716 9034
rect 78776 8974 78782 9034
rect 79222 8924 79282 9102
rect 75152 8734 75212 8880
rect 78218 8864 79282 8924
rect 80746 8776 80752 8836
rect 80812 8776 80818 8836
rect 74938 8728 75426 8734
rect 74938 8694 74950 8728
rect 75414 8694 75426 8728
rect 74938 8688 75426 8694
rect 75956 8728 76444 8734
rect 75956 8694 75968 8728
rect 76432 8694 76444 8728
rect 75956 8688 76444 8694
rect 76974 8728 77462 8734
rect 76974 8694 76986 8728
rect 77450 8694 77462 8728
rect 76974 8688 77462 8694
rect 77992 8728 78480 8734
rect 77992 8694 78004 8728
rect 78468 8694 78480 8728
rect 77992 8688 78480 8694
rect 79010 8728 79498 8734
rect 79010 8694 79022 8728
rect 79486 8694 79498 8728
rect 79010 8688 79498 8694
rect 80028 8728 80516 8734
rect 80028 8694 80040 8728
rect 80504 8694 80516 8728
rect 80028 8688 80516 8694
rect 73672 8068 73678 8608
rect 74640 8606 74656 8644
rect 73632 8056 73678 8068
rect 74650 8068 74656 8606
rect 74690 8606 74700 8644
rect 75668 8644 75714 8656
rect 74690 8068 74696 8606
rect 75668 8110 75674 8644
rect 74650 8056 74696 8068
rect 75660 8068 75674 8110
rect 75708 8110 75714 8644
rect 76686 8644 76732 8656
rect 75708 8068 75720 8110
rect 76686 8106 76692 8644
rect 72902 8018 73390 8024
rect 72902 7984 72914 8018
rect 73378 7984 73390 8018
rect 72902 7978 73390 7984
rect 73920 8018 74408 8024
rect 73920 7984 73932 8018
rect 74396 7984 74408 8018
rect 73920 7978 74408 7984
rect 74938 8018 75426 8024
rect 74938 7984 74950 8018
rect 75414 7984 75426 8018
rect 74938 7978 75426 7984
rect 73110 7922 73170 7978
rect 74116 7922 74176 7978
rect 75160 7922 75220 7978
rect 75660 7928 75720 8068
rect 76680 8068 76692 8106
rect 76726 8106 76732 8644
rect 77704 8644 77750 8656
rect 76726 8068 76740 8106
rect 77704 8100 77710 8644
rect 75956 8018 76444 8024
rect 75956 7984 75968 8018
rect 76432 7984 76444 8018
rect 75956 7978 76444 7984
rect 73104 7862 73110 7922
rect 73170 7862 73176 7922
rect 74110 7862 74116 7922
rect 74176 7862 74182 7922
rect 75154 7862 75160 7922
rect 75220 7862 75226 7922
rect 75654 7868 75660 7928
rect 75720 7868 75726 7928
rect 73110 7500 73170 7862
rect 74108 7646 74114 7706
rect 74174 7646 74180 7706
rect 75148 7646 75154 7706
rect 75214 7646 75220 7706
rect 74114 7500 74174 7646
rect 74632 7542 74638 7602
rect 74698 7542 74704 7602
rect 72902 7494 73390 7500
rect 72902 7460 72914 7494
rect 73378 7460 73390 7494
rect 72902 7454 73390 7460
rect 73920 7494 74408 7500
rect 73920 7460 73932 7494
rect 74396 7460 74408 7494
rect 73920 7454 74408 7460
rect 72608 7328 72620 7410
rect 72614 6880 72620 7328
rect 71636 6834 71650 6880
rect 70866 6784 71354 6790
rect 70866 6750 70878 6784
rect 71342 6750 71354 6784
rect 70866 6744 71354 6750
rect 71056 6694 71116 6744
rect 71050 6634 71056 6694
rect 71116 6634 71122 6694
rect 71590 6478 71650 6834
rect 72610 6834 72620 6880
rect 72654 7328 72668 7410
rect 73632 7410 73678 7422
rect 72654 6880 72660 7328
rect 72654 6834 72670 6880
rect 73632 6878 73638 7410
rect 71884 6784 72372 6790
rect 71884 6750 71896 6784
rect 72360 6750 72372 6784
rect 71884 6744 72372 6750
rect 72094 6694 72154 6744
rect 72088 6634 72094 6694
rect 72154 6634 72160 6694
rect 71584 6418 71590 6478
rect 71650 6418 71656 6478
rect 70564 6320 70570 6380
rect 70630 6320 70636 6380
rect 72094 6266 72154 6634
rect 72610 6380 72670 6834
rect 73628 6834 73638 6878
rect 73672 6878 73678 7410
rect 74638 7410 74698 7542
rect 75154 7500 75214 7646
rect 74938 7494 75426 7500
rect 74938 7460 74950 7494
rect 75414 7460 75426 7494
rect 74938 7454 75426 7460
rect 74638 7346 74656 7410
rect 73672 6834 73688 6878
rect 72902 6784 73390 6790
rect 72902 6750 72914 6784
rect 73378 6750 73390 6784
rect 72902 6744 73390 6750
rect 73112 6694 73172 6744
rect 73628 6700 73688 6834
rect 74650 6834 74656 7346
rect 74690 7346 74698 7410
rect 75660 7410 75720 7868
rect 76168 7706 76228 7978
rect 76162 7646 76168 7706
rect 76228 7646 76234 7706
rect 76168 7500 76228 7646
rect 76680 7602 76740 8068
rect 77696 8068 77710 8100
rect 77744 8100 77750 8644
rect 78722 8644 78768 8656
rect 78722 8102 78728 8644
rect 77744 8068 77756 8100
rect 76974 8018 77462 8024
rect 76974 7984 76986 8018
rect 77450 7984 77462 8018
rect 76974 7978 77462 7984
rect 77176 7706 77236 7978
rect 77696 7928 77756 8068
rect 78718 8068 78728 8102
rect 78762 8102 78768 8644
rect 79740 8644 79786 8656
rect 78762 8068 78778 8102
rect 79740 8100 79746 8644
rect 77992 8018 78480 8024
rect 77992 7984 78004 8018
rect 78468 7984 78480 8018
rect 77992 7978 78480 7984
rect 77690 7868 77696 7928
rect 77756 7868 77762 7928
rect 78220 7706 78280 7978
rect 77170 7646 77176 7706
rect 77236 7646 77242 7706
rect 78214 7646 78220 7706
rect 78280 7646 78286 7706
rect 76674 7542 76680 7602
rect 76740 7542 76746 7602
rect 75956 7494 76444 7500
rect 75956 7460 75968 7494
rect 76432 7460 76444 7494
rect 75956 7454 76444 7460
rect 75660 7374 75674 7410
rect 74690 6834 74696 7346
rect 75668 6892 75674 7374
rect 74650 6822 74696 6834
rect 75664 6834 75674 6892
rect 75708 7374 75720 7410
rect 76680 7410 76740 7542
rect 77176 7500 77236 7646
rect 78220 7500 78280 7646
rect 78718 7602 78778 8068
rect 79732 8068 79746 8100
rect 79780 8100 79786 8644
rect 80752 8644 80812 8776
rect 81046 8728 81534 8734
rect 81046 8694 81058 8728
rect 81522 8694 81534 8728
rect 81046 8688 81534 8694
rect 79780 8068 79792 8100
rect 79010 8018 79498 8024
rect 79010 7984 79022 8018
rect 79486 7984 79498 8018
rect 79010 7978 79498 7984
rect 79210 7706 79270 7978
rect 79732 7928 79792 8068
rect 80752 8068 80764 8644
rect 80798 8068 80812 8644
rect 81768 8644 81828 9300
rect 82788 9300 82800 9334
rect 82834 9836 82846 9876
rect 83804 9876 83864 10016
rect 84310 9966 84370 10080
rect 85326 9966 85386 10080
rect 85836 10016 85842 10076
rect 85902 10016 85908 10076
rect 84100 9960 84588 9966
rect 84100 9926 84112 9960
rect 84576 9926 84588 9960
rect 84100 9920 84588 9926
rect 85118 9960 85606 9966
rect 85118 9926 85130 9960
rect 85594 9926 85606 9960
rect 85118 9920 85606 9926
rect 82834 9334 82840 9836
rect 83804 9834 83818 9876
rect 82834 9300 82848 9334
rect 82064 9250 82552 9256
rect 82064 9216 82076 9250
rect 82540 9216 82552 9250
rect 82064 9210 82552 9216
rect 82264 8940 82324 9210
rect 82258 8880 82264 8940
rect 82324 8880 82330 8940
rect 82264 8734 82324 8880
rect 82064 8728 82552 8734
rect 82064 8694 82076 8728
rect 82540 8694 82552 8728
rect 82064 8688 82552 8694
rect 81768 8604 81782 8644
rect 81776 8100 81782 8604
rect 80028 8018 80516 8024
rect 80028 7984 80040 8018
rect 80504 7984 80516 8018
rect 80028 7978 80516 7984
rect 79726 7868 79732 7928
rect 79792 7868 79798 7928
rect 80228 7706 80288 7978
rect 79204 7646 79210 7706
rect 79270 7646 79276 7706
rect 80222 7646 80228 7706
rect 80288 7646 80294 7706
rect 78712 7542 78718 7602
rect 78778 7542 78784 7602
rect 76974 7494 77462 7500
rect 76974 7460 76986 7494
rect 77450 7460 77462 7494
rect 76974 7454 77462 7460
rect 77992 7494 78480 7500
rect 77992 7460 78004 7494
rect 78468 7460 78480 7494
rect 77992 7454 78480 7460
rect 75708 6892 75714 7374
rect 76680 7372 76692 7410
rect 75708 6834 75724 6892
rect 73920 6784 74408 6790
rect 73920 6750 73932 6784
rect 74396 6750 74408 6784
rect 73920 6744 74408 6750
rect 74938 6784 75426 6790
rect 74938 6750 74950 6784
rect 75414 6750 75426 6784
rect 74938 6744 75426 6750
rect 75664 6700 75724 6834
rect 76686 6834 76692 7372
rect 76726 7372 76740 7410
rect 77704 7410 77750 7422
rect 76726 6834 76732 7372
rect 77704 6884 77710 7410
rect 76686 6822 76732 6834
rect 77696 6834 77710 6884
rect 77744 6884 77750 7410
rect 78718 7410 78778 7542
rect 79210 7500 79270 7646
rect 80752 7602 80812 8068
rect 81770 8068 81782 8100
rect 81816 8604 81828 8644
rect 82788 8644 82848 9300
rect 83812 9300 83818 9834
rect 83852 9834 83864 9876
rect 84830 9876 84876 9888
rect 83852 9300 83858 9834
rect 84830 9358 84836 9876
rect 83812 9288 83858 9300
rect 84822 9300 84836 9358
rect 84870 9358 84876 9876
rect 85842 9876 85902 10016
rect 86344 9966 86404 10444
rect 86860 10406 86920 10534
rect 87878 10534 87890 10592
rect 87924 11082 87936 11110
rect 87924 10592 87930 11082
rect 87924 10534 87938 10592
rect 87154 10484 87642 10490
rect 87154 10450 87166 10484
rect 87630 10450 87642 10484
rect 87154 10444 87642 10450
rect 87878 10424 87938 10534
rect 86854 10346 86860 10406
rect 86920 10346 86926 10406
rect 87872 10364 87878 10424
rect 87938 10364 87944 10424
rect 86860 10128 86920 10346
rect 86860 10068 87934 10128
rect 87984 10076 88044 11252
rect 88472 10234 88478 10294
rect 88538 10234 88544 10294
rect 88222 10130 88228 10190
rect 88288 10130 88294 10190
rect 86136 9960 86624 9966
rect 86136 9926 86148 9960
rect 86612 9926 86624 9960
rect 86136 9920 86624 9926
rect 85842 9834 85854 9876
rect 84870 9300 84882 9358
rect 83294 9256 83354 9258
rect 83082 9250 83570 9256
rect 83082 9216 83094 9250
rect 83558 9216 83570 9250
rect 83082 9210 83570 9216
rect 84100 9250 84588 9256
rect 84100 9216 84112 9250
rect 84576 9216 84588 9250
rect 84100 9210 84588 9216
rect 83294 8940 83354 9210
rect 84316 9162 84376 9210
rect 84310 9102 84316 9162
rect 84376 9102 84382 9162
rect 84448 9106 84454 9166
rect 84514 9106 84520 9166
rect 84454 8940 84514 9106
rect 84822 8940 84882 9300
rect 85848 9300 85854 9834
rect 85888 9834 85902 9876
rect 86860 9876 86920 10068
rect 87364 9966 87424 10068
rect 87154 9960 87642 9966
rect 87154 9926 87166 9960
rect 87630 9926 87642 9960
rect 87154 9920 87642 9926
rect 86860 9842 86872 9876
rect 85888 9300 85894 9834
rect 86866 9340 86872 9842
rect 85848 9288 85894 9300
rect 86860 9300 86872 9340
rect 86906 9842 86920 9876
rect 87874 9876 87934 10068
rect 87978 10016 87984 10076
rect 88044 10016 88050 10076
rect 87874 9852 87890 9876
rect 86906 9340 86912 9842
rect 86906 9300 86920 9340
rect 85118 9250 85606 9256
rect 85118 9216 85130 9250
rect 85594 9216 85606 9250
rect 85118 9210 85606 9216
rect 86136 9250 86624 9256
rect 86136 9216 86148 9250
rect 86612 9216 86624 9250
rect 86136 9210 86624 9216
rect 86342 9166 86402 9210
rect 85330 9106 85336 9166
rect 85396 9106 85402 9166
rect 86336 9106 86342 9166
rect 86402 9106 86408 9166
rect 86860 9162 86920 9300
rect 87884 9300 87890 9852
rect 87924 9852 87934 9876
rect 87924 9300 87930 9852
rect 87884 9288 87930 9300
rect 87154 9250 87642 9256
rect 87154 9216 87166 9250
rect 87630 9216 87642 9250
rect 87154 9210 87642 9216
rect 83288 8880 83294 8940
rect 83354 8880 83360 8940
rect 84448 8880 84454 8940
rect 84514 8880 84520 8940
rect 84816 8880 84822 8940
rect 84882 8880 84888 8940
rect 83294 8734 83354 8880
rect 84454 8734 84514 8880
rect 84822 8836 84882 8880
rect 84816 8776 84822 8836
rect 84882 8776 84888 8836
rect 85336 8734 85396 9106
rect 86854 9102 86860 9162
rect 86920 9102 86926 9162
rect 86854 8974 86860 9034
rect 86920 8974 86926 9034
rect 85832 8778 85838 8838
rect 85898 8778 85904 8838
rect 83082 8728 83570 8734
rect 83082 8694 83094 8728
rect 83558 8694 83570 8728
rect 83082 8688 83570 8694
rect 84100 8728 84588 8734
rect 84100 8694 84112 8728
rect 84576 8694 84588 8728
rect 84100 8688 84588 8694
rect 85118 8728 85606 8734
rect 85118 8694 85130 8728
rect 85594 8694 85606 8728
rect 85118 8688 85606 8694
rect 85336 8686 85396 8688
rect 81816 8100 81822 8604
rect 82788 8598 82800 8644
rect 82794 8112 82800 8598
rect 81816 8068 81830 8100
rect 81046 8018 81534 8024
rect 81046 7984 81058 8018
rect 81522 7984 81534 8018
rect 81046 7978 81534 7984
rect 81262 7706 81322 7978
rect 81770 7928 81830 8068
rect 82786 8068 82800 8112
rect 82834 8598 82848 8644
rect 83812 8644 83858 8656
rect 82834 8112 82840 8598
rect 82834 8068 82846 8112
rect 83812 8108 83818 8644
rect 82064 8018 82552 8024
rect 82064 7984 82076 8018
rect 82540 7984 82552 8018
rect 82064 7978 82552 7984
rect 81764 7868 81770 7928
rect 81830 7868 81836 7928
rect 81756 7760 81762 7820
rect 81822 7760 81828 7820
rect 81256 7646 81262 7706
rect 81322 7646 81328 7706
rect 80746 7542 80752 7602
rect 80812 7542 80818 7602
rect 81258 7538 81264 7598
rect 81324 7538 81330 7598
rect 81264 7500 81324 7538
rect 79010 7494 79498 7500
rect 79010 7460 79022 7494
rect 79486 7460 79498 7494
rect 79010 7454 79498 7460
rect 80028 7494 80516 7500
rect 80028 7460 80040 7494
rect 80504 7460 80516 7494
rect 80028 7454 80516 7460
rect 81046 7494 81534 7500
rect 81046 7460 81058 7494
rect 81522 7460 81534 7494
rect 81046 7454 81534 7460
rect 78718 7374 78728 7410
rect 77744 6834 77756 6884
rect 75956 6784 76444 6790
rect 75956 6750 75968 6784
rect 76432 6750 76444 6784
rect 75956 6744 76444 6750
rect 76974 6784 77462 6790
rect 76974 6750 76986 6784
rect 77450 6750 77462 6784
rect 76974 6744 77462 6750
rect 77696 6700 77756 6834
rect 78722 6834 78728 7374
rect 78762 7374 78778 7410
rect 79740 7410 79786 7422
rect 78762 6834 78768 7374
rect 79740 6896 79746 7410
rect 78722 6822 78768 6834
rect 79730 6834 79746 6896
rect 79780 6896 79786 7410
rect 80758 7410 80804 7422
rect 79780 6834 79790 6896
rect 80758 6876 80764 7410
rect 77992 6784 78480 6790
rect 77992 6750 78004 6784
rect 78468 6750 78480 6784
rect 77992 6744 78480 6750
rect 79010 6784 79498 6790
rect 79010 6750 79022 6784
rect 79486 6750 79498 6784
rect 79010 6744 79498 6750
rect 79730 6700 79790 6834
rect 80752 6834 80764 6876
rect 80798 6876 80804 7410
rect 81762 7410 81822 7760
rect 82286 7598 82346 7978
rect 82786 7604 82846 8068
rect 83806 8068 83818 8108
rect 83852 8108 83858 8644
rect 84830 8644 84876 8656
rect 84830 8112 84836 8644
rect 83852 8068 83866 8108
rect 83082 8018 83570 8024
rect 83082 7984 83094 8018
rect 83558 7984 83570 8018
rect 83082 7978 83570 7984
rect 82280 7538 82286 7598
rect 82346 7538 82352 7598
rect 82780 7544 82786 7604
rect 82846 7544 82852 7604
rect 82286 7500 82346 7538
rect 82064 7494 82552 7500
rect 82064 7460 82076 7494
rect 82540 7460 82552 7494
rect 82064 7454 82552 7460
rect 81762 7374 81782 7410
rect 80798 6834 80812 6876
rect 80028 6784 80516 6790
rect 80028 6750 80040 6784
rect 80504 6750 80516 6784
rect 80028 6744 80516 6750
rect 73106 6634 73112 6694
rect 73172 6634 73178 6694
rect 73622 6640 73628 6700
rect 73688 6640 73694 6700
rect 77690 6640 77696 6700
rect 77756 6640 77762 6700
rect 79724 6640 79730 6700
rect 79790 6640 79796 6700
rect 72604 6320 72610 6380
rect 72670 6320 72676 6380
rect 68830 6260 69318 6266
rect 68830 6226 68842 6260
rect 69306 6226 69318 6260
rect 68830 6220 69318 6226
rect 69848 6260 70336 6266
rect 69848 6226 69860 6260
rect 70324 6226 70336 6260
rect 69848 6220 70336 6226
rect 70866 6260 71354 6266
rect 70866 6226 70878 6260
rect 71342 6226 71354 6260
rect 70866 6220 71354 6226
rect 71884 6260 72372 6266
rect 71884 6226 71896 6260
rect 72360 6226 72372 6260
rect 71884 6220 72372 6226
rect 68532 6122 68548 6176
rect 67564 5600 67574 5634
rect 68542 5630 68548 6122
rect 67514 5468 67574 5600
rect 68538 5600 68548 5630
rect 68582 6122 68592 6176
rect 69560 6176 69606 6188
rect 68582 5630 68588 6122
rect 69560 5646 69566 6176
rect 68582 5600 68598 5630
rect 67812 5550 68300 5556
rect 67812 5516 67824 5550
rect 68288 5516 68300 5550
rect 67812 5510 68300 5516
rect 68034 5468 68094 5510
rect 68538 5468 68598 5600
rect 69552 5600 69566 5646
rect 69600 5646 69606 6176
rect 70578 6176 70624 6188
rect 69600 5600 69612 5646
rect 70578 5630 70584 6176
rect 68830 5550 69318 5556
rect 68830 5516 68842 5550
rect 69306 5516 69318 5550
rect 68830 5510 69318 5516
rect 67514 5408 68598 5468
rect 67392 5298 67398 5358
rect 67458 5298 67464 5358
rect 68538 5262 68598 5408
rect 67514 5202 68598 5262
rect 67514 4944 67574 5202
rect 68026 5034 68086 5202
rect 68538 5142 68598 5202
rect 68532 5082 68538 5142
rect 68598 5082 68604 5142
rect 67812 5028 68300 5034
rect 67812 4994 67824 5028
rect 68288 4994 68300 5028
rect 67812 4988 68300 4994
rect 67514 4908 67530 4944
rect 67524 4368 67530 4908
rect 67564 4908 67574 4944
rect 68538 4944 68598 5082
rect 69030 5034 69090 5510
rect 69552 5456 69612 5600
rect 70570 5600 70584 5630
rect 70618 5630 70624 6176
rect 71596 6176 71642 6188
rect 71596 5642 71602 6176
rect 70618 5600 70630 5630
rect 69848 5550 70336 5556
rect 69848 5516 69860 5550
rect 70324 5516 70336 5550
rect 69848 5510 70336 5516
rect 69546 5396 69552 5456
rect 69612 5396 69618 5456
rect 69550 5202 69556 5262
rect 69616 5202 69622 5262
rect 68830 5028 69318 5034
rect 68830 4994 68842 5028
rect 69306 4994 69318 5028
rect 68830 4988 69318 4994
rect 67564 4368 67570 4908
rect 68538 4904 68548 4944
rect 67524 4356 67570 4368
rect 68542 4368 68548 4904
rect 68582 4904 68598 4944
rect 69556 4944 69616 5202
rect 70050 5198 70110 5510
rect 70570 5358 70630 5600
rect 71588 5600 71602 5642
rect 71636 5642 71642 6176
rect 72610 6176 72670 6320
rect 73112 6266 73172 6634
rect 72902 6260 73390 6266
rect 72902 6226 72914 6260
rect 73378 6226 73390 6260
rect 72902 6220 73390 6226
rect 72610 6146 72620 6176
rect 72614 5664 72620 6146
rect 71636 5600 71648 5642
rect 70866 5550 71354 5556
rect 70866 5516 70878 5550
rect 71342 5516 71354 5550
rect 70866 5510 71354 5516
rect 70564 5298 70570 5358
rect 70630 5298 70636 5358
rect 71084 5198 71144 5510
rect 71588 5456 71648 5600
rect 72606 5600 72620 5664
rect 72654 6146 72670 6176
rect 73628 6176 73688 6640
rect 75664 6634 75724 6640
rect 76674 6530 76680 6590
rect 76740 6530 76746 6590
rect 78710 6530 78716 6590
rect 78776 6530 78782 6590
rect 75656 6418 75662 6478
rect 75722 6418 75728 6478
rect 74640 6320 74646 6380
rect 74706 6320 74712 6380
rect 73920 6260 74408 6266
rect 73920 6226 73932 6260
rect 74396 6226 74408 6260
rect 73920 6220 74408 6226
rect 72654 5664 72660 6146
rect 73628 6134 73638 6176
rect 72654 5600 72666 5664
rect 73632 5640 73638 6134
rect 71884 5550 72372 5556
rect 71884 5516 71896 5550
rect 72360 5516 72372 5550
rect 71884 5510 72372 5516
rect 71582 5396 71588 5456
rect 71648 5396 71654 5456
rect 72094 5358 72154 5510
rect 72088 5298 72094 5358
rect 72154 5298 72160 5358
rect 71586 5202 71592 5262
rect 71652 5202 71658 5262
rect 70050 5138 71144 5198
rect 70050 5034 70110 5138
rect 71084 5034 71144 5138
rect 69848 5028 70336 5034
rect 69848 4994 69860 5028
rect 70324 4994 70336 5028
rect 69848 4988 70336 4994
rect 70866 5028 71354 5034
rect 70866 4994 70878 5028
rect 71342 4994 71354 5028
rect 70866 4988 71354 4994
rect 68582 4368 68588 4904
rect 69556 4900 69566 4944
rect 68542 4356 68588 4368
rect 69560 4368 69566 4900
rect 69600 4900 69616 4944
rect 70578 4944 70624 4956
rect 69600 4368 69606 4900
rect 70578 4410 70584 4944
rect 69560 4356 69606 4368
rect 70570 4368 70584 4410
rect 70618 4410 70624 4944
rect 71592 4944 71652 5202
rect 72094 5034 72154 5298
rect 72606 5142 72666 5600
rect 73626 5600 73638 5640
rect 73672 6134 73688 6176
rect 74646 6176 74706 6320
rect 74938 6260 75426 6266
rect 74938 6226 74950 6260
rect 75414 6226 75426 6260
rect 74938 6220 75426 6226
rect 74646 6140 74656 6176
rect 73672 5640 73678 6134
rect 73672 5600 73686 5640
rect 74650 5634 74656 6140
rect 72902 5550 73390 5556
rect 72902 5516 72914 5550
rect 73378 5516 73390 5550
rect 72902 5510 73390 5516
rect 73116 5358 73176 5510
rect 73626 5456 73686 5600
rect 74640 5600 74656 5634
rect 74690 6140 74706 6176
rect 75662 6176 75722 6418
rect 75956 6260 76444 6266
rect 75956 6226 75968 6260
rect 76432 6226 76444 6260
rect 75956 6220 76444 6226
rect 75662 6150 75674 6176
rect 74690 5634 74696 6140
rect 75668 5656 75674 6150
rect 74690 5600 74700 5634
rect 73920 5550 74408 5556
rect 73920 5516 73932 5550
rect 74396 5516 74408 5550
rect 73920 5510 74408 5516
rect 73620 5396 73626 5456
rect 73686 5396 73692 5456
rect 74140 5364 74200 5510
rect 72600 5082 72606 5142
rect 72666 5082 72672 5142
rect 71884 5028 72372 5034
rect 71884 4994 71896 5028
rect 72360 4994 72372 5028
rect 71884 4988 72372 4994
rect 71592 4892 71602 4944
rect 70618 4368 70630 4410
rect 67812 4318 68300 4324
rect 67812 4284 67824 4318
rect 68288 4284 68300 4318
rect 67812 4278 68300 4284
rect 68830 4318 69318 4324
rect 68830 4284 68842 4318
rect 69306 4284 69318 4318
rect 68830 4278 69318 4284
rect 69848 4318 70336 4324
rect 69848 4284 69860 4318
rect 70324 4284 70336 4318
rect 69848 4278 70336 4284
rect 67280 4166 67286 4226
rect 67346 4166 67352 4226
rect 70570 4100 70630 4368
rect 71596 4368 71602 4892
rect 71636 4892 71652 4944
rect 72606 4944 72666 5082
rect 73116 5034 73176 5298
rect 74138 5358 74200 5364
rect 74198 5298 74200 5358
rect 74138 5292 74200 5298
rect 73614 5202 73620 5262
rect 73680 5202 73686 5262
rect 72902 5028 73390 5034
rect 72902 4994 72914 5028
rect 73378 4994 73390 5028
rect 72902 4988 73390 4994
rect 72606 4904 72620 4944
rect 71636 4368 71642 4892
rect 72614 4422 72620 4904
rect 71596 4356 71642 4368
rect 72608 4368 72620 4422
rect 72654 4904 72666 4944
rect 73620 4944 73680 5202
rect 74140 5034 74200 5292
rect 74640 5142 74700 5600
rect 75658 5600 75674 5656
rect 75708 6150 75722 6176
rect 76680 6176 76740 6530
rect 76974 6260 77462 6266
rect 76974 6226 76986 6260
rect 77450 6226 77462 6260
rect 76974 6220 77462 6226
rect 77992 6260 78480 6266
rect 77992 6226 78004 6260
rect 78468 6226 78480 6260
rect 77992 6220 78480 6226
rect 75708 5656 75714 6150
rect 76680 6144 76692 6176
rect 75708 5600 75718 5656
rect 74938 5550 75426 5556
rect 74938 5516 74950 5550
rect 75414 5516 75426 5550
rect 74938 5510 75426 5516
rect 75142 5358 75202 5510
rect 75488 5476 75548 5482
rect 75658 5476 75718 5600
rect 76686 5600 76692 6144
rect 76726 6144 76740 6176
rect 77704 6176 77750 6188
rect 76726 5600 76732 6144
rect 77704 5670 77710 6176
rect 76686 5588 76732 5600
rect 77700 5600 77710 5670
rect 77744 5670 77750 6176
rect 78716 6176 78776 6530
rect 80258 6492 80318 6744
rect 80752 6702 80812 6834
rect 81776 6834 81782 7374
rect 81816 6834 81822 7410
rect 82786 7410 82846 7544
rect 83264 7500 83324 7978
rect 83806 7928 83866 8068
rect 84820 8068 84836 8112
rect 84870 8112 84876 8644
rect 85838 8644 85898 8778
rect 86136 8728 86624 8734
rect 86136 8694 86148 8728
rect 86612 8694 86624 8728
rect 86136 8688 86624 8694
rect 85838 8594 85854 8644
rect 84870 8068 84880 8112
rect 85848 8096 85854 8594
rect 84100 8018 84588 8024
rect 84100 7984 84112 8018
rect 84576 7984 84588 8018
rect 84100 7978 84588 7984
rect 83800 7868 83806 7928
rect 83866 7868 83872 7928
rect 83796 7760 83802 7820
rect 83862 7760 83868 7820
rect 83082 7494 83570 7500
rect 83082 7460 83094 7494
rect 83558 7460 83570 7494
rect 83082 7454 83570 7460
rect 82786 7316 82800 7410
rect 82794 6876 82800 7316
rect 81776 6822 81822 6834
rect 82786 6834 82800 6876
rect 82834 7316 82846 7410
rect 83802 7410 83862 7760
rect 84288 7646 84294 7706
rect 84354 7646 84360 7706
rect 84294 7500 84354 7646
rect 84820 7604 84880 8068
rect 85844 8068 85854 8096
rect 85888 8594 85898 8644
rect 86860 8644 86920 8974
rect 87154 8728 87642 8734
rect 87154 8694 87166 8728
rect 87630 8694 87642 8728
rect 87154 8688 87642 8694
rect 85888 8096 85894 8594
rect 86860 8592 86872 8644
rect 86866 8096 86872 8592
rect 85888 8068 85904 8096
rect 85118 8018 85606 8024
rect 85118 7984 85130 8018
rect 85594 7984 85606 8018
rect 85118 7978 85606 7984
rect 85844 7928 85904 8068
rect 86860 8068 86872 8096
rect 86906 8592 86920 8644
rect 87884 8644 87930 8656
rect 86906 8096 86912 8592
rect 87884 8102 87890 8644
rect 86906 8068 86920 8096
rect 86136 8018 86624 8024
rect 86136 7984 86148 8018
rect 86612 7984 86624 8018
rect 86136 7978 86624 7984
rect 85838 7868 85844 7928
rect 85904 7868 85910 7928
rect 85834 7760 85840 7820
rect 85900 7760 85906 7820
rect 85326 7646 85332 7706
rect 85392 7646 85398 7706
rect 84814 7544 84820 7604
rect 84880 7544 84886 7604
rect 85332 7500 85392 7646
rect 84100 7494 84588 7500
rect 84100 7460 84112 7494
rect 84576 7460 84588 7494
rect 84100 7454 84588 7460
rect 85118 7494 85606 7500
rect 85118 7460 85130 7494
rect 85594 7460 85606 7494
rect 85118 7454 85606 7460
rect 83802 7344 83818 7410
rect 82834 6876 82840 7316
rect 82834 6834 82846 6876
rect 81046 6784 81534 6790
rect 81046 6750 81058 6784
rect 81522 6750 81534 6784
rect 81046 6744 81534 6750
rect 82064 6784 82552 6790
rect 82064 6750 82076 6784
rect 82540 6750 82552 6784
rect 82064 6744 82552 6750
rect 80746 6642 80752 6702
rect 80812 6642 80818 6702
rect 81100 6642 81106 6702
rect 81166 6642 81172 6702
rect 80742 6530 80748 6590
rect 80808 6530 80814 6590
rect 80252 6432 80258 6492
rect 80318 6432 80324 6492
rect 79010 6260 79498 6266
rect 79010 6226 79022 6260
rect 79486 6226 79498 6260
rect 79010 6220 79498 6226
rect 80028 6260 80516 6266
rect 80028 6226 80040 6260
rect 80504 6226 80516 6260
rect 80028 6220 80516 6226
rect 78716 6138 78728 6176
rect 77744 5600 77760 5670
rect 75956 5550 76444 5556
rect 75956 5516 75968 5550
rect 76432 5516 76444 5550
rect 75956 5510 76444 5516
rect 76974 5550 77462 5556
rect 76974 5516 76986 5550
rect 77450 5516 77462 5550
rect 76974 5510 77462 5516
rect 75652 5416 75658 5476
rect 75718 5416 75724 5476
rect 75136 5298 75142 5358
rect 75202 5298 75208 5358
rect 74634 5082 74640 5142
rect 74700 5082 74706 5142
rect 73920 5028 74408 5034
rect 73920 4994 73932 5028
rect 74396 4994 74408 5028
rect 73920 4988 74408 4994
rect 72654 4422 72660 4904
rect 73620 4884 73638 4944
rect 72654 4368 72668 4422
rect 70866 4318 71354 4324
rect 70866 4284 70878 4318
rect 71342 4284 71354 4318
rect 70866 4278 71354 4284
rect 71884 4318 72372 4324
rect 71884 4284 71896 4318
rect 72360 4284 72372 4318
rect 71884 4278 72372 4284
rect 71090 4112 71150 4278
rect 67174 4040 67180 4100
rect 67240 4040 67246 4100
rect 70564 4040 70570 4100
rect 70630 4040 70636 4100
rect 71084 4052 71090 4112
rect 71150 4052 71156 4112
rect 69546 3930 69552 3990
rect 69612 3930 69618 3990
rect 71582 3930 71588 3990
rect 71648 3930 71654 3990
rect 67812 3794 68300 3800
rect 67812 3760 67824 3794
rect 68288 3760 68300 3794
rect 67812 3754 68300 3760
rect 68830 3794 69318 3800
rect 68830 3760 68842 3794
rect 69306 3760 69318 3794
rect 68830 3754 69318 3760
rect 67524 3710 67570 3722
rect 67524 3160 67530 3710
rect 67518 3134 67530 3160
rect 67564 3160 67570 3710
rect 68542 3710 68588 3722
rect 68542 3188 68548 3710
rect 67564 3134 67578 3160
rect 67518 2996 67578 3134
rect 68530 3134 68548 3188
rect 68582 3188 68588 3710
rect 69552 3710 69612 3930
rect 71200 3836 71206 3896
rect 71266 3836 71272 3896
rect 71206 3800 71266 3836
rect 69848 3794 70336 3800
rect 69848 3760 69860 3794
rect 70324 3760 70336 3794
rect 69848 3754 70336 3760
rect 70866 3794 71354 3800
rect 70866 3760 70878 3794
rect 71342 3760 71354 3794
rect 70866 3754 71354 3760
rect 69552 3650 69566 3710
rect 68582 3134 68590 3188
rect 67812 3084 68300 3090
rect 67812 3050 67824 3084
rect 68288 3050 68300 3084
rect 67812 3044 68300 3050
rect 68032 2996 68092 3044
rect 68530 2996 68590 3134
rect 69560 3134 69566 3650
rect 69600 3650 69612 3710
rect 70578 3710 70624 3722
rect 69600 3134 69606 3650
rect 70578 3178 70584 3710
rect 69560 3122 69606 3134
rect 70572 3134 70584 3178
rect 70618 3178 70624 3710
rect 71588 3710 71648 3930
rect 72090 3896 72150 4278
rect 72608 3990 72668 4368
rect 73632 4368 73638 4884
rect 73672 4884 73680 4944
rect 74640 4944 74700 5082
rect 75142 5034 75202 5298
rect 75488 5262 75548 5416
rect 75482 5202 75488 5262
rect 75548 5202 75554 5262
rect 75658 5208 75664 5268
rect 75724 5208 75730 5268
rect 74938 5028 75426 5034
rect 74938 4994 74950 5028
rect 75414 4994 75426 5028
rect 74938 4988 75426 4994
rect 74640 4904 74656 4944
rect 73672 4368 73678 4884
rect 74650 4434 74656 4904
rect 73632 4356 73678 4368
rect 74644 4368 74656 4434
rect 74690 4904 74700 4944
rect 75664 4944 75724 5208
rect 76180 5206 76240 5510
rect 77194 5370 77254 5510
rect 77700 5476 77760 5600
rect 78722 5600 78728 6138
rect 78762 6138 78776 6176
rect 79740 6176 79786 6188
rect 78762 5600 78768 6138
rect 79740 5670 79746 6176
rect 78722 5588 78768 5600
rect 79732 5600 79746 5670
rect 79780 5670 79786 6176
rect 80748 6176 80808 6530
rect 81106 6384 81166 6642
rect 81296 6492 81356 6744
rect 82272 6492 82332 6744
rect 81290 6432 81296 6492
rect 81356 6432 81362 6492
rect 82266 6432 82272 6492
rect 82332 6432 82338 6492
rect 82786 6380 82846 6834
rect 83812 6834 83818 7344
rect 83852 7344 83862 7410
rect 84830 7410 84876 7422
rect 83852 6834 83858 7344
rect 84830 6878 84836 7410
rect 83812 6822 83858 6834
rect 84824 6834 84836 6878
rect 84870 6878 84876 7410
rect 85840 7410 85900 7760
rect 86358 7706 86418 7978
rect 86860 7886 86920 8068
rect 87874 8068 87890 8102
rect 87924 8102 87930 8644
rect 87924 8068 87934 8102
rect 87154 8018 87642 8024
rect 87154 7984 87166 8018
rect 87630 7984 87642 8018
rect 87154 7978 87642 7984
rect 87368 7886 87428 7978
rect 87874 7886 87934 8068
rect 86860 7826 87934 7886
rect 86352 7646 86358 7706
rect 86418 7646 86424 7706
rect 86856 7544 86862 7604
rect 86922 7544 86928 7604
rect 86136 7494 86624 7500
rect 86136 7460 86148 7494
rect 86612 7460 86624 7494
rect 86136 7454 86624 7460
rect 85840 7358 85854 7410
rect 85848 6884 85854 7358
rect 84870 6834 84884 6878
rect 83082 6784 83570 6790
rect 83082 6750 83094 6784
rect 83558 6750 83570 6784
rect 83082 6744 83570 6750
rect 84100 6784 84588 6790
rect 84100 6750 84112 6784
rect 84576 6750 84588 6784
rect 84100 6744 84588 6750
rect 83288 6492 83348 6744
rect 84824 6702 84884 6834
rect 85842 6834 85854 6884
rect 85888 7358 85900 7410
rect 86862 7410 86922 7544
rect 87154 7494 87642 7500
rect 87154 7460 87166 7494
rect 87630 7460 87642 7494
rect 87154 7454 87642 7460
rect 86862 7376 86872 7410
rect 85888 6884 85894 7358
rect 85888 6834 85902 6884
rect 86866 6878 86872 7376
rect 85118 6784 85606 6790
rect 85118 6750 85130 6784
rect 85594 6750 85606 6784
rect 85118 6744 85606 6750
rect 84818 6642 84824 6702
rect 84884 6642 84890 6702
rect 83282 6432 83288 6492
rect 83348 6432 83354 6492
rect 85308 6432 85314 6492
rect 85374 6432 85380 6492
rect 81106 6318 81166 6324
rect 82780 6320 82786 6380
rect 82846 6320 82852 6380
rect 84816 6320 84822 6380
rect 84882 6320 84888 6380
rect 81046 6260 81534 6266
rect 81046 6226 81058 6260
rect 81522 6226 81534 6260
rect 81046 6220 81534 6226
rect 82064 6260 82552 6266
rect 82064 6226 82076 6260
rect 82540 6226 82552 6260
rect 82064 6220 82552 6226
rect 80748 6134 80764 6176
rect 79780 5600 79792 5670
rect 77992 5550 78480 5556
rect 77992 5516 78004 5550
rect 78468 5516 78480 5550
rect 77992 5510 78480 5516
rect 79010 5550 79498 5556
rect 79010 5516 79022 5550
rect 79486 5516 79498 5550
rect 79010 5510 79498 5516
rect 77694 5416 77700 5476
rect 77760 5416 77766 5476
rect 78216 5370 78276 5510
rect 79230 5370 79290 5510
rect 79732 5476 79792 5600
rect 80758 5600 80764 6134
rect 80798 6134 80808 6176
rect 81776 6176 81822 6188
rect 80798 5600 80804 6134
rect 81776 5636 81782 6176
rect 80758 5588 80804 5600
rect 81772 5600 81782 5636
rect 81816 5636 81822 6176
rect 82786 6176 82846 6320
rect 83082 6260 83570 6266
rect 83082 6226 83094 6260
rect 83558 6226 83570 6260
rect 83082 6220 83570 6226
rect 84100 6260 84588 6266
rect 84100 6226 84112 6260
rect 84576 6226 84588 6260
rect 84100 6220 84588 6226
rect 82786 6138 82800 6176
rect 82794 5652 82800 6138
rect 81816 5600 81832 5636
rect 80028 5550 80516 5556
rect 80028 5516 80040 5550
rect 80504 5516 80516 5550
rect 80028 5510 80516 5516
rect 81046 5550 81534 5556
rect 81046 5516 81058 5550
rect 81522 5516 81534 5550
rect 81046 5510 81534 5516
rect 79726 5416 79732 5476
rect 79792 5416 79798 5476
rect 80232 5470 80292 5510
rect 81258 5470 81318 5510
rect 81772 5476 81832 5600
rect 82790 5600 82800 5652
rect 82834 6138 82846 6176
rect 83812 6176 83858 6188
rect 82834 5652 82840 6138
rect 82834 5600 82850 5652
rect 83812 5644 83818 6176
rect 82064 5550 82552 5556
rect 82064 5516 82076 5550
rect 82540 5516 82552 5550
rect 82064 5510 82552 5516
rect 80232 5410 81318 5470
rect 81766 5416 81772 5476
rect 81832 5416 81838 5476
rect 80232 5370 80292 5410
rect 77194 5310 80292 5370
rect 80744 5318 80750 5378
rect 80810 5318 80816 5378
rect 77194 5206 77254 5310
rect 77686 5208 77692 5268
rect 77752 5208 77758 5268
rect 76180 5146 77254 5206
rect 76180 5034 76240 5146
rect 77194 5034 77254 5146
rect 75956 5028 76444 5034
rect 75956 4994 75968 5028
rect 76432 4994 76444 5028
rect 75956 4988 76444 4994
rect 76974 5028 77462 5034
rect 76974 4994 76986 5028
rect 77450 4994 77462 5028
rect 76974 4988 77462 4994
rect 74690 4434 74696 4904
rect 75664 4900 75674 4944
rect 74690 4368 74704 4434
rect 72902 4318 73390 4324
rect 72902 4284 72914 4318
rect 73378 4284 73390 4318
rect 72902 4278 73390 4284
rect 73920 4318 74408 4324
rect 73920 4284 73932 4318
rect 74396 4284 74408 4318
rect 73920 4278 74408 4284
rect 72602 3930 72608 3990
rect 72668 3930 72674 3990
rect 73112 3896 73172 4278
rect 74644 3990 74704 4368
rect 75668 4368 75674 4900
rect 75708 4900 75724 4944
rect 76686 4944 76732 4956
rect 75708 4368 75714 4900
rect 76686 4420 76692 4944
rect 75668 4356 75714 4368
rect 76674 4368 76692 4420
rect 76726 4420 76732 4944
rect 77692 4944 77752 5208
rect 78216 5034 78276 5310
rect 79230 5034 79290 5310
rect 79730 5208 79736 5268
rect 79796 5208 79802 5268
rect 77992 5028 78480 5034
rect 77992 4994 78004 5028
rect 78468 4994 78480 5028
rect 77992 4988 78480 4994
rect 79010 5028 79498 5034
rect 79010 4994 79022 5028
rect 79486 4994 79498 5028
rect 79010 4988 79498 4994
rect 77692 4900 77710 4944
rect 76726 4368 76734 4420
rect 74938 4318 75426 4324
rect 74938 4284 74950 4318
rect 75414 4284 75426 4318
rect 74938 4278 75426 4284
rect 75956 4318 76444 4324
rect 75956 4284 75968 4318
rect 76432 4284 76444 4318
rect 75956 4278 76444 4284
rect 73618 3930 73624 3990
rect 73684 3930 73690 3990
rect 74638 3930 74644 3990
rect 74704 3930 74710 3990
rect 72084 3836 72090 3896
rect 72150 3836 72156 3896
rect 73106 3836 73112 3896
rect 73172 3836 73178 3896
rect 72090 3800 72150 3836
rect 73112 3800 73172 3836
rect 71884 3794 72372 3800
rect 71884 3760 71896 3794
rect 72360 3760 72372 3794
rect 71884 3754 72372 3760
rect 72902 3794 73390 3800
rect 72902 3760 72914 3794
rect 73378 3760 73390 3794
rect 72902 3754 73390 3760
rect 71588 3660 71602 3710
rect 71596 3196 71602 3660
rect 70618 3134 70632 3178
rect 68830 3084 69318 3090
rect 68830 3050 68842 3084
rect 69306 3050 69318 3084
rect 68830 3044 69318 3050
rect 69848 3084 70336 3090
rect 69848 3050 69860 3084
rect 70324 3050 70336 3084
rect 69848 3044 70336 3050
rect 67512 2936 67518 2996
rect 67578 2936 67584 2996
rect 68026 2936 68032 2996
rect 68092 2936 68098 2996
rect 68524 2936 68530 2996
rect 68590 2936 68596 2996
rect 69046 2778 69106 3044
rect 70068 2778 70128 3044
rect 70572 2996 70632 3134
rect 71586 3134 71602 3196
rect 71636 3660 71648 3710
rect 72614 3710 72660 3722
rect 71636 3196 71642 3660
rect 71636 3134 71646 3196
rect 72614 3174 72620 3710
rect 70866 3084 71354 3090
rect 70866 3050 70878 3084
rect 71342 3050 71354 3084
rect 70866 3044 71354 3050
rect 70566 2936 70572 2996
rect 70632 2936 70638 2996
rect 71080 2884 71140 3044
rect 71074 2824 71080 2884
rect 71140 2824 71146 2884
rect 67054 2718 67060 2778
rect 67120 2718 67126 2778
rect 69040 2718 69046 2778
rect 69106 2718 69112 2778
rect 70062 2718 70068 2778
rect 70128 2718 70134 2778
rect 71586 2674 71646 3134
rect 72604 3134 72620 3174
rect 72654 3174 72660 3710
rect 73624 3710 73684 3930
rect 75154 3896 75214 4278
rect 76170 4112 76230 4278
rect 76674 4226 76734 4368
rect 77704 4368 77710 4900
rect 77744 4900 77752 4944
rect 78722 4944 78768 4956
rect 77744 4368 77750 4900
rect 78722 4420 78728 4944
rect 77704 4356 77750 4368
rect 78716 4368 78728 4420
rect 78762 4420 78768 4944
rect 79736 4944 79796 5208
rect 80232 5034 80292 5310
rect 80028 5028 80516 5034
rect 80028 4994 80040 5028
rect 80504 4994 80516 5028
rect 80028 4988 80516 4994
rect 79736 4896 79746 4944
rect 78762 4368 78776 4420
rect 76974 4318 77462 4324
rect 76974 4284 76986 4318
rect 77450 4284 77462 4318
rect 76974 4278 77462 4284
rect 77992 4318 78480 4324
rect 77992 4284 78004 4318
rect 78468 4284 78480 4318
rect 77992 4278 78480 4284
rect 78716 4226 78776 4368
rect 79740 4368 79746 4896
rect 79780 4896 79796 4944
rect 80750 4944 80810 5318
rect 81258 5034 81318 5410
rect 81758 5208 81764 5268
rect 81824 5208 81830 5268
rect 81046 5028 81534 5034
rect 81046 4994 81058 5028
rect 81522 4994 81534 5028
rect 81046 4988 81534 4994
rect 80750 4908 80764 4944
rect 79780 4368 79786 4896
rect 80758 4412 80764 4908
rect 79740 4356 79786 4368
rect 80752 4368 80764 4412
rect 80798 4908 80810 4944
rect 81764 4944 81824 5208
rect 82278 5034 82338 5510
rect 82790 5142 82850 5600
rect 83802 5600 83818 5644
rect 83852 5644 83858 6176
rect 84822 6176 84882 6320
rect 85314 6266 85374 6432
rect 85118 6260 85606 6266
rect 85118 6226 85130 6260
rect 85594 6226 85606 6260
rect 85118 6220 85606 6226
rect 84822 6118 84836 6176
rect 83852 5600 83862 5644
rect 84830 5640 84836 6118
rect 83082 5550 83570 5556
rect 83082 5516 83094 5550
rect 83558 5516 83570 5550
rect 83082 5510 83570 5516
rect 82784 5082 82790 5142
rect 82850 5082 82856 5142
rect 82064 5028 82552 5034
rect 82064 4994 82076 5028
rect 82540 4994 82552 5028
rect 82064 4988 82552 4994
rect 80798 4412 80804 4908
rect 81764 4896 81782 4944
rect 80798 4368 80812 4412
rect 79010 4318 79498 4324
rect 79010 4284 79022 4318
rect 79486 4284 79498 4318
rect 79010 4278 79498 4284
rect 80028 4318 80516 4324
rect 80028 4284 80040 4318
rect 80504 4284 80516 4318
rect 80028 4278 80516 4284
rect 80752 4226 80812 4368
rect 81776 4368 81782 4896
rect 81816 4896 81824 4944
rect 82790 4944 82850 5082
rect 83294 5034 83354 5510
rect 83802 5268 83862 5600
rect 84820 5600 84836 5640
rect 84870 6118 84882 6176
rect 85842 6176 85902 6834
rect 86858 6834 86872 6878
rect 86906 7376 86922 7410
rect 87884 7410 87930 7422
rect 86906 6878 86912 7376
rect 86906 6834 86918 6878
rect 87884 6864 87890 7410
rect 86136 6784 86624 6790
rect 86136 6750 86148 6784
rect 86612 6750 86624 6784
rect 86136 6744 86624 6750
rect 86344 6492 86404 6744
rect 86858 6652 86918 6834
rect 87874 6834 87890 6864
rect 87924 6864 87930 7410
rect 87924 6834 87934 6864
rect 87154 6784 87642 6790
rect 87154 6750 87166 6784
rect 87630 6750 87642 6784
rect 87154 6744 87642 6750
rect 87364 6652 87424 6744
rect 87874 6652 87934 6834
rect 86858 6592 87934 6652
rect 86338 6432 86344 6492
rect 86404 6432 86410 6492
rect 86858 6380 86918 6592
rect 86852 6320 86858 6380
rect 86918 6320 86924 6380
rect 86136 6260 86624 6266
rect 86136 6226 86148 6260
rect 86612 6226 86624 6260
rect 86136 6220 86624 6226
rect 87154 6260 87642 6266
rect 87154 6226 87166 6260
rect 87630 6226 87642 6260
rect 87154 6220 87642 6226
rect 85842 6134 85854 6176
rect 84870 5640 84876 6118
rect 85848 5654 85854 6134
rect 84870 5600 84880 5640
rect 84100 5550 84588 5556
rect 84100 5516 84112 5550
rect 84576 5516 84588 5550
rect 84100 5510 84588 5516
rect 83796 5208 83802 5268
rect 83862 5208 83868 5268
rect 84328 5034 84388 5510
rect 84820 5142 84880 5600
rect 85842 5600 85854 5654
rect 85888 6134 85902 6176
rect 86866 6176 86912 6188
rect 85888 5654 85894 6134
rect 85888 5600 85902 5654
rect 86866 5646 86872 6176
rect 85118 5550 85606 5556
rect 85118 5516 85130 5550
rect 85594 5516 85606 5550
rect 85118 5510 85606 5516
rect 85346 5144 85406 5510
rect 85842 5268 85902 5600
rect 86856 5600 86872 5646
rect 86906 5646 86912 6176
rect 87884 6176 87930 6188
rect 86906 5600 86916 5646
rect 87884 5628 87890 6176
rect 86136 5550 86624 5556
rect 86136 5516 86148 5550
rect 86612 5516 86624 5550
rect 86136 5510 86624 5516
rect 86360 5272 86420 5510
rect 86856 5474 86916 5600
rect 87876 5600 87890 5628
rect 87924 5628 87930 6176
rect 87924 5600 87936 5628
rect 87154 5550 87642 5556
rect 87154 5516 87166 5550
rect 87630 5516 87642 5550
rect 87154 5510 87642 5516
rect 87362 5476 87422 5510
rect 87876 5476 87936 5600
rect 87362 5474 87936 5476
rect 86856 5414 87936 5474
rect 86856 5378 86916 5414
rect 86850 5318 86856 5378
rect 86916 5318 86922 5378
rect 85836 5208 85842 5268
rect 85902 5208 85908 5268
rect 86354 5212 86360 5272
rect 86420 5212 86426 5272
rect 84814 5082 84820 5142
rect 84880 5082 84886 5142
rect 83082 5028 83570 5034
rect 83082 4994 83094 5028
rect 83558 4994 83570 5028
rect 83082 4988 83570 4994
rect 84100 5028 84588 5034
rect 84100 4994 84112 5028
rect 84576 4994 84588 5028
rect 84100 4988 84588 4994
rect 82790 4898 82800 4944
rect 81816 4368 81822 4896
rect 82794 4428 82800 4898
rect 81776 4356 81822 4368
rect 82788 4368 82800 4428
rect 82834 4898 82850 4944
rect 83812 4944 83858 4956
rect 82834 4428 82840 4898
rect 82834 4368 82848 4428
rect 83812 4412 83818 4944
rect 81046 4318 81534 4324
rect 81046 4284 81058 4318
rect 81522 4284 81534 4318
rect 81046 4278 81534 4284
rect 82064 4318 82552 4324
rect 82064 4284 82076 4318
rect 82540 4284 82552 4318
rect 82064 4278 82552 4284
rect 76668 4166 76674 4226
rect 76734 4166 76740 4226
rect 78710 4166 78716 4226
rect 78776 4166 78782 4226
rect 80746 4166 80752 4226
rect 80812 4166 80818 4226
rect 81258 4116 81318 4278
rect 76164 4052 76170 4112
rect 76230 4052 76236 4112
rect 81252 4056 81258 4116
rect 81318 4056 81324 4116
rect 75656 3930 75662 3990
rect 75722 3930 75728 3990
rect 77686 3930 77692 3990
rect 77752 3930 77758 3990
rect 79724 3930 79730 3990
rect 79790 3930 79796 3990
rect 81760 3930 81766 3990
rect 81826 3930 81832 3990
rect 75148 3836 75154 3896
rect 75214 3836 75220 3896
rect 73920 3794 74408 3800
rect 73920 3760 73932 3794
rect 74396 3760 74408 3794
rect 73920 3754 74408 3760
rect 74938 3794 75426 3800
rect 74938 3760 74950 3794
rect 75414 3760 75426 3794
rect 74938 3754 75426 3760
rect 72654 3134 72664 3174
rect 71884 3084 72372 3090
rect 71884 3050 71896 3084
rect 72360 3050 72372 3084
rect 71884 3044 72372 3050
rect 72092 2884 72152 3044
rect 72604 2996 72664 3134
rect 73624 3134 73638 3710
rect 73672 3134 73684 3710
rect 74650 3710 74696 3722
rect 74650 3174 74656 3710
rect 72902 3084 73390 3090
rect 72902 3050 72914 3084
rect 73378 3050 73390 3084
rect 72902 3044 73390 3050
rect 72598 2936 72604 2996
rect 72664 2936 72670 2996
rect 73106 2884 73166 3044
rect 72086 2824 72092 2884
rect 72152 2824 72158 2884
rect 73100 2824 73106 2884
rect 73166 2824 73172 2884
rect 72600 2718 72606 2778
rect 72666 2718 72672 2778
rect 73112 2718 73118 2778
rect 73178 2718 73184 2778
rect 66648 2614 66654 2674
rect 66714 2614 66720 2674
rect 71076 2614 71082 2674
rect 71142 2614 71148 2674
rect 71580 2614 71586 2674
rect 71646 2614 71652 2674
rect 72096 2614 72102 2674
rect 72162 2614 72168 2674
rect 66020 1566 66026 1626
rect 66086 1566 66092 1626
rect 62818 540 62824 600
rect 62884 540 62890 600
rect 64006 540 64012 600
rect 64072 540 64078 600
rect 65202 540 65208 600
rect 65268 540 65274 600
rect 65896 540 65902 600
rect 65962 540 65968 600
rect 66654 110 66714 2614
rect 71082 2566 71142 2614
rect 67812 2560 68300 2566
rect 67812 2526 67824 2560
rect 68288 2526 68300 2560
rect 67812 2520 68300 2526
rect 68830 2560 69318 2566
rect 68830 2526 68842 2560
rect 69306 2526 69318 2560
rect 68830 2520 69318 2526
rect 69848 2560 70336 2566
rect 69848 2526 69860 2560
rect 70324 2526 70336 2560
rect 69848 2520 70336 2526
rect 70866 2560 71354 2566
rect 70866 2526 70878 2560
rect 71342 2526 71354 2560
rect 70866 2520 71354 2526
rect 67524 2476 67570 2488
rect 67524 1926 67530 2476
rect 67518 1900 67530 1926
rect 67564 1926 67570 2476
rect 68542 2476 68588 2488
rect 68542 1928 68548 2476
rect 67564 1900 67578 1926
rect 67518 1444 67578 1900
rect 68530 1900 68548 1928
rect 68582 1928 68588 2476
rect 69560 2476 69606 2488
rect 69560 1932 69566 2476
rect 68582 1900 68590 1928
rect 67812 1850 68300 1856
rect 67812 1816 67824 1850
rect 68288 1816 68300 1850
rect 67812 1810 68300 1816
rect 67512 1384 67518 1444
rect 67578 1384 67584 1444
rect 67518 1244 67578 1384
rect 68016 1334 68076 1810
rect 68530 1542 68590 1900
rect 69548 1900 69566 1932
rect 69600 1932 69606 2476
rect 70578 2476 70624 2488
rect 70578 1940 70584 2476
rect 69600 1900 69608 1932
rect 68830 1850 69318 1856
rect 68830 1816 68842 1850
rect 69306 1816 69318 1850
rect 68830 1810 69318 1816
rect 68524 1482 68530 1542
rect 68590 1482 68596 1542
rect 67812 1328 68300 1334
rect 67812 1294 67824 1328
rect 68288 1294 68300 1328
rect 67812 1288 68300 1294
rect 67518 1188 67530 1244
rect 67524 668 67530 1188
rect 67564 1188 67578 1244
rect 68530 1244 68590 1482
rect 69038 1334 69098 1810
rect 69548 1444 69608 1900
rect 70568 1900 70584 1940
rect 70618 1940 70624 2476
rect 71586 2476 71646 2614
rect 72102 2566 72162 2614
rect 71884 2560 72372 2566
rect 71884 2526 71896 2560
rect 72360 2526 72372 2560
rect 71884 2520 72372 2526
rect 72606 2476 72666 2718
rect 73118 2566 73178 2718
rect 73624 2674 73684 3134
rect 74636 3134 74656 3174
rect 74690 3134 74696 3710
rect 75662 3710 75722 3930
rect 76168 3854 77238 3914
rect 76168 3800 76228 3854
rect 75956 3794 76444 3800
rect 75956 3760 75968 3794
rect 76432 3760 76444 3794
rect 75956 3754 76444 3760
rect 75662 3654 75674 3710
rect 75668 3186 75674 3654
rect 73920 3084 74408 3090
rect 73920 3050 73932 3084
rect 74396 3050 74408 3084
rect 73920 3044 74408 3050
rect 74136 2778 74196 3044
rect 74636 2996 74696 3134
rect 75662 3134 75674 3186
rect 75708 3654 75722 3710
rect 76680 3710 76740 3854
rect 77178 3800 77238 3854
rect 76974 3794 77462 3800
rect 76974 3760 76986 3794
rect 77450 3760 77462 3794
rect 76974 3754 77462 3760
rect 76680 3674 76692 3710
rect 75708 3186 75714 3654
rect 75708 3134 75722 3186
rect 76686 3178 76692 3674
rect 76678 3170 76692 3178
rect 76672 3134 76692 3170
rect 76726 3674 76740 3710
rect 77692 3710 77752 3930
rect 78192 3858 79280 3918
rect 78192 3800 78252 3858
rect 77992 3794 78480 3800
rect 77992 3760 78004 3794
rect 78468 3760 78480 3794
rect 77992 3754 78480 3760
rect 76726 3178 76732 3674
rect 77692 3660 77710 3710
rect 77704 3184 77710 3660
rect 76726 3134 76738 3178
rect 74938 3084 75426 3090
rect 74938 3050 74950 3084
rect 75414 3050 75426 3084
rect 74938 3044 75426 3050
rect 74630 2936 74636 2996
rect 74696 2936 74702 2996
rect 75148 2778 75208 3044
rect 74130 2718 74136 2778
rect 74196 2718 74202 2778
rect 74636 2718 74642 2778
rect 74702 2718 74708 2778
rect 75142 2718 75148 2778
rect 75208 2718 75214 2778
rect 73618 2614 73624 2674
rect 73684 2614 73690 2674
rect 72902 2560 73390 2566
rect 72902 2526 72914 2560
rect 73378 2526 73390 2560
rect 72902 2520 73390 2526
rect 71586 2424 71602 2476
rect 70618 1900 70628 1940
rect 69848 1850 70336 1856
rect 69848 1816 69860 1850
rect 70324 1816 70336 1850
rect 69848 1810 70336 1816
rect 69542 1384 69548 1444
rect 69608 1384 69614 1444
rect 68830 1328 69318 1334
rect 68830 1294 68842 1328
rect 69306 1294 69318 1328
rect 68830 1288 69318 1294
rect 68530 1206 68548 1244
rect 67564 668 67570 1188
rect 68542 718 68548 1206
rect 67524 656 67570 668
rect 68532 668 68548 718
rect 68582 1206 68590 1244
rect 69548 1244 69608 1384
rect 70064 1334 70124 1810
rect 70568 1542 70628 1900
rect 71596 1900 71602 2424
rect 71636 2424 71646 2476
rect 71636 1900 71642 2424
rect 72604 2420 72620 2476
rect 72614 1942 72620 2420
rect 71596 1888 71642 1900
rect 72604 1900 72620 1942
rect 72654 2424 72666 2476
rect 73624 2476 73684 2614
rect 74136 2566 74196 2718
rect 73920 2560 74408 2566
rect 73920 2526 73932 2560
rect 74396 2526 74408 2560
rect 73920 2520 74408 2526
rect 74642 2476 74702 2718
rect 75148 2566 75208 2718
rect 75662 2674 75722 3134
rect 75956 3084 76444 3090
rect 75956 3050 75968 3084
rect 76432 3050 76444 3084
rect 75956 3044 76444 3050
rect 76012 2824 76018 2884
rect 76078 2824 76084 2884
rect 75656 2614 75662 2674
rect 75722 2614 75728 2674
rect 74938 2560 75426 2566
rect 74938 2526 74950 2560
rect 75414 2526 75426 2560
rect 74938 2520 75426 2526
rect 73624 2426 73638 2476
rect 72654 2420 72664 2424
rect 72654 1942 72660 2420
rect 72654 1900 72664 1942
rect 70866 1850 71354 1856
rect 70866 1816 70878 1850
rect 71342 1816 71354 1850
rect 70866 1810 71354 1816
rect 71884 1850 72372 1856
rect 71884 1816 71896 1850
rect 72360 1816 72372 1850
rect 71884 1810 72372 1816
rect 72604 1756 72664 1900
rect 73632 1900 73638 2426
rect 73672 2426 73684 2476
rect 73672 1900 73678 2426
rect 74636 2410 74656 2476
rect 74650 1934 74656 2410
rect 73632 1888 73678 1900
rect 74642 1900 74656 1934
rect 74690 2436 74702 2476
rect 75662 2476 75722 2614
rect 76018 2566 76078 2824
rect 76160 2778 76220 3044
rect 76540 2996 76600 3002
rect 76154 2718 76160 2778
rect 76220 2718 76226 2778
rect 76540 2766 76600 2936
rect 76678 2886 76738 3134
rect 77698 3134 77710 3184
rect 77744 3660 77752 3710
rect 78716 3710 78776 3858
rect 79220 3800 79280 3858
rect 79010 3794 79498 3800
rect 79010 3760 79022 3794
rect 79486 3760 79498 3794
rect 79010 3754 79498 3760
rect 78716 3678 78728 3710
rect 77744 3184 77750 3660
rect 78722 3188 78728 3678
rect 77744 3134 77758 3184
rect 76974 3084 77462 3090
rect 76974 3050 76986 3084
rect 77450 3050 77462 3084
rect 76974 3044 77462 3050
rect 76672 2826 76678 2886
rect 76738 2826 76744 2886
rect 77180 2778 77240 3044
rect 77300 2822 77306 2882
rect 77366 2822 77372 2882
rect 76540 2706 76740 2766
rect 77174 2718 77180 2778
rect 77240 2718 77246 2778
rect 75956 2560 76444 2566
rect 75956 2526 75968 2560
rect 76432 2526 76444 2560
rect 75956 2520 76444 2526
rect 74690 1934 74696 2436
rect 75662 2416 75674 2476
rect 74690 1900 74702 1934
rect 72902 1850 73390 1856
rect 72902 1816 72914 1850
rect 73378 1816 73390 1850
rect 72902 1810 73390 1816
rect 73920 1850 74408 1856
rect 73920 1816 73932 1850
rect 74396 1816 74408 1850
rect 73920 1810 74408 1816
rect 73108 1756 73168 1810
rect 72604 1696 73168 1756
rect 74124 1748 74184 1810
rect 74642 1748 74702 1900
rect 75668 1900 75674 2416
rect 75708 2416 75722 2476
rect 76680 2476 76740 2706
rect 77306 2566 77366 2822
rect 77698 2674 77758 3134
rect 78714 3134 78728 3188
rect 78762 3678 78776 3710
rect 79730 3710 79790 3930
rect 80028 3794 80516 3800
rect 80028 3760 80040 3794
rect 80504 3760 80516 3794
rect 80028 3754 80516 3760
rect 81046 3794 81534 3800
rect 81046 3760 81058 3794
rect 81522 3760 81534 3794
rect 81046 3754 81534 3760
rect 78762 3188 78768 3678
rect 79730 3666 79746 3710
rect 78762 3134 78774 3188
rect 79740 3172 79746 3666
rect 77992 3084 78480 3090
rect 77992 3050 78004 3084
rect 78468 3050 78480 3084
rect 77992 3044 78480 3050
rect 78202 2778 78262 3044
rect 78346 2822 78352 2882
rect 78412 2822 78418 2882
rect 78196 2718 78202 2778
rect 78262 2718 78268 2778
rect 77692 2614 77698 2674
rect 77758 2614 77764 2674
rect 76974 2560 77462 2566
rect 76974 2526 76986 2560
rect 77450 2526 77462 2560
rect 76974 2520 77462 2526
rect 76680 2448 76692 2476
rect 75708 1900 75714 2416
rect 76686 1924 76692 2448
rect 75668 1888 75714 1900
rect 76680 1900 76692 1924
rect 76726 2448 76740 2476
rect 77698 2476 77758 2614
rect 78352 2566 78412 2822
rect 78714 2778 78774 3134
rect 79734 3134 79746 3172
rect 79780 3666 79790 3710
rect 80758 3710 80804 3722
rect 79780 3172 79786 3666
rect 80758 3194 80764 3710
rect 79780 3134 79794 3172
rect 79010 3084 79498 3090
rect 79010 3050 79022 3084
rect 79486 3050 79498 3084
rect 79010 3044 79498 3050
rect 78900 2998 78960 3004
rect 78708 2718 78714 2778
rect 78774 2718 78780 2778
rect 78900 2670 78960 2938
rect 79220 2778 79280 3044
rect 79214 2718 79220 2778
rect 79280 2718 79286 2778
rect 78716 2610 78960 2670
rect 77992 2560 78480 2566
rect 77992 2526 78004 2560
rect 78468 2526 78480 2560
rect 77992 2520 78480 2526
rect 76726 1924 76732 2448
rect 77698 2410 77710 2476
rect 76726 1900 76740 1924
rect 74938 1850 75426 1856
rect 74938 1816 74950 1850
rect 75414 1816 75426 1850
rect 74938 1810 75426 1816
rect 75956 1850 76444 1856
rect 75956 1816 75968 1850
rect 76432 1816 76444 1850
rect 75956 1810 76444 1816
rect 75150 1748 75210 1810
rect 74124 1688 75210 1748
rect 76170 1638 76230 1810
rect 76680 1742 76740 1900
rect 77704 1900 77710 2410
rect 77744 2410 77758 2476
rect 78716 2476 78776 2610
rect 79220 2566 79280 2718
rect 79734 2674 79794 3134
rect 80750 3134 80764 3194
rect 80798 3194 80804 3710
rect 81766 3710 81826 3930
rect 82276 3896 82336 4278
rect 82788 3990 82848 4368
rect 83806 4368 83818 4412
rect 83852 4412 83858 4944
rect 84820 4944 84880 5082
rect 85346 5034 85406 5084
rect 86360 5034 86420 5212
rect 86858 5144 87936 5202
rect 86852 5084 86858 5144
rect 86918 5142 87936 5144
rect 86918 5084 86924 5142
rect 85118 5028 85606 5034
rect 85118 4994 85130 5028
rect 85594 4994 85606 5028
rect 85118 4988 85606 4994
rect 86136 5028 86624 5034
rect 86136 4994 86148 5028
rect 86612 4994 86624 5028
rect 86136 4988 86624 4994
rect 84820 4898 84836 4944
rect 84830 4416 84836 4898
rect 83852 4368 83866 4412
rect 83082 4318 83570 4324
rect 83082 4284 83094 4318
rect 83558 4284 83570 4318
rect 83082 4278 83570 4284
rect 82782 3930 82788 3990
rect 82848 3930 82854 3990
rect 83296 3896 83356 4278
rect 83806 4226 83866 4368
rect 84822 4368 84836 4416
rect 84870 4898 84880 4944
rect 85848 4944 85894 4956
rect 84870 4416 84876 4898
rect 84870 4368 84882 4416
rect 85848 4412 85854 4944
rect 84100 4318 84588 4324
rect 84100 4284 84112 4318
rect 84576 4284 84588 4318
rect 84100 4278 84588 4284
rect 83800 4166 83806 4226
rect 83866 4166 83872 4226
rect 83802 3930 83808 3990
rect 83868 3930 83874 3990
rect 82270 3836 82276 3896
rect 82336 3836 82342 3896
rect 83290 3836 83296 3896
rect 83356 3836 83362 3896
rect 82276 3800 82336 3836
rect 83296 3800 83356 3836
rect 82064 3794 82552 3800
rect 82064 3760 82076 3794
rect 82540 3760 82552 3794
rect 82064 3754 82552 3760
rect 83082 3794 83570 3800
rect 83082 3760 83094 3794
rect 83558 3760 83570 3794
rect 83082 3754 83570 3760
rect 81766 3666 81782 3710
rect 80798 3134 80810 3194
rect 81776 3188 81782 3666
rect 80028 3084 80516 3090
rect 80028 3050 80040 3084
rect 80504 3050 80516 3084
rect 80028 3044 80516 3050
rect 80238 2778 80298 3044
rect 80750 2996 80810 3134
rect 81766 3134 81782 3188
rect 81816 3666 81826 3710
rect 82794 3710 82840 3722
rect 81816 3188 81822 3666
rect 81816 3134 81826 3188
rect 82794 3166 82800 3710
rect 81046 3084 81534 3090
rect 81046 3050 81058 3084
rect 81522 3050 81534 3084
rect 81046 3044 81534 3050
rect 80744 2936 80750 2996
rect 80810 2936 80816 2996
rect 81258 2778 81318 3044
rect 80232 2718 80238 2778
rect 80298 2718 80304 2778
rect 80744 2718 80750 2778
rect 80810 2718 80816 2778
rect 81252 2718 81258 2778
rect 81318 2718 81324 2778
rect 79728 2614 79734 2674
rect 79794 2614 79800 2674
rect 79010 2560 79498 2566
rect 79010 2526 79022 2560
rect 79486 2526 79498 2560
rect 79010 2520 79498 2526
rect 78716 2442 78728 2476
rect 77744 1900 77750 2410
rect 78722 1966 78728 2442
rect 77704 1888 77750 1900
rect 78716 1900 78728 1966
rect 78762 2442 78776 2476
rect 79734 2476 79794 2614
rect 80238 2566 80298 2718
rect 80028 2560 80516 2566
rect 80028 2526 80040 2560
rect 80504 2526 80516 2560
rect 80028 2520 80516 2526
rect 80750 2476 80810 2718
rect 81258 2566 81318 2718
rect 81766 2674 81826 3134
rect 82784 3134 82800 3166
rect 82834 3166 82840 3710
rect 83808 3710 83868 3930
rect 84310 3896 84370 4278
rect 84822 3990 84882 4368
rect 85838 4368 85854 4412
rect 85888 4412 85894 4944
rect 86858 4944 86918 5084
rect 87360 5034 87420 5142
rect 87154 5028 87642 5034
rect 87154 4994 87166 5028
rect 87630 4994 87642 5028
rect 87154 4988 87642 4994
rect 86858 4910 86872 4944
rect 85888 4368 85898 4412
rect 85118 4318 85606 4324
rect 85118 4284 85130 4318
rect 85594 4284 85606 4318
rect 85118 4278 85606 4284
rect 84816 3930 84822 3990
rect 84882 3930 84888 3990
rect 85346 3896 85406 4278
rect 85838 4226 85898 4368
rect 86866 4368 86872 4910
rect 86906 4910 86918 4944
rect 87876 4944 87936 5142
rect 86906 4368 86912 4910
rect 87876 4906 87890 4944
rect 86866 4356 86912 4368
rect 87884 4368 87890 4906
rect 87924 4906 87936 4944
rect 87924 4368 87930 4906
rect 87884 4356 87930 4368
rect 86136 4318 86624 4324
rect 86136 4284 86148 4318
rect 86612 4284 86624 4318
rect 86136 4278 86624 4284
rect 87154 4318 87642 4324
rect 87154 4284 87166 4318
rect 87630 4284 87642 4318
rect 87154 4278 87642 4284
rect 85832 4166 85838 4226
rect 85898 4166 85904 4226
rect 86358 4116 86418 4278
rect 87984 4226 88044 10016
rect 88106 9102 88112 9162
rect 88172 9102 88178 9162
rect 88112 7604 88172 9102
rect 88228 8838 88288 10130
rect 88344 8880 88350 8940
rect 88410 8880 88416 8940
rect 88222 8778 88228 8838
rect 88288 8778 88294 8838
rect 88106 7544 88112 7604
rect 88172 7544 88178 7604
rect 88102 6642 88108 6702
rect 88168 6642 88174 6702
rect 88108 5378 88168 6642
rect 88228 5476 88288 8778
rect 88222 5416 88228 5476
rect 88288 5416 88294 5476
rect 88102 5318 88108 5378
rect 88168 5318 88174 5378
rect 88350 5144 88410 8880
rect 88478 7712 88538 10234
rect 88476 7706 88538 7712
rect 88536 7646 88538 7706
rect 88476 7640 88538 7646
rect 88478 5272 88538 7640
rect 88472 5212 88478 5272
rect 88538 5212 88544 5272
rect 88344 5084 88350 5144
rect 88410 5084 88416 5144
rect 87978 4166 87984 4226
rect 88044 4166 88050 4226
rect 86352 4056 86358 4116
rect 86418 4056 86424 4116
rect 86358 3992 86418 4056
rect 85838 3930 85844 3990
rect 85904 3930 85910 3990
rect 86358 3932 88104 3992
rect 84304 3836 84310 3896
rect 84370 3836 84376 3896
rect 85340 3836 85346 3896
rect 85406 3836 85412 3896
rect 84310 3800 84370 3836
rect 84100 3794 84588 3800
rect 84100 3760 84112 3794
rect 84576 3760 84588 3794
rect 84100 3754 84588 3760
rect 85118 3794 85606 3800
rect 85118 3760 85130 3794
rect 85594 3760 85606 3794
rect 85118 3754 85606 3760
rect 84318 3750 84378 3754
rect 83808 3644 83818 3710
rect 83812 3182 83818 3644
rect 82834 3134 82844 3166
rect 82064 3084 82552 3090
rect 82064 3050 82076 3084
rect 82540 3050 82552 3084
rect 82064 3044 82552 3050
rect 82280 2882 82340 3044
rect 82784 2996 82844 3134
rect 83804 3134 83818 3182
rect 83852 3644 83868 3710
rect 84830 3710 84876 3722
rect 83852 3182 83858 3644
rect 84830 3184 84836 3710
rect 83852 3134 83864 3182
rect 83082 3084 83570 3090
rect 83082 3050 83094 3084
rect 83558 3050 83570 3084
rect 83082 3044 83570 3050
rect 82778 2936 82784 2996
rect 82844 2936 82850 2996
rect 83298 2882 83358 3044
rect 82274 2822 82280 2882
rect 82340 2822 82346 2882
rect 83292 2822 83298 2882
rect 83358 2822 83364 2882
rect 83804 2674 83864 3134
rect 84818 3134 84836 3184
rect 84870 3184 84876 3710
rect 85844 3710 85904 3930
rect 86136 3794 86624 3800
rect 86136 3760 86148 3794
rect 86612 3760 86624 3794
rect 86136 3754 86624 3760
rect 87154 3794 87642 3800
rect 87154 3760 87166 3794
rect 87630 3760 87642 3794
rect 87154 3754 87642 3760
rect 85844 3650 85854 3710
rect 84870 3134 84878 3184
rect 84100 3084 84588 3090
rect 84100 3050 84112 3084
rect 84576 3050 84588 3084
rect 84100 3044 84588 3050
rect 84306 2888 84366 3044
rect 84818 2996 84878 3134
rect 85848 3134 85854 3650
rect 85888 3650 85904 3710
rect 86866 3710 86912 3722
rect 85888 3134 85894 3650
rect 86866 3178 86872 3710
rect 85848 3122 85894 3134
rect 86860 3134 86872 3178
rect 86906 3178 86912 3710
rect 87884 3710 87930 3722
rect 86906 3134 86920 3178
rect 87884 3176 87890 3710
rect 85118 3084 85606 3090
rect 85118 3050 85130 3084
rect 85594 3050 85606 3084
rect 85118 3044 85606 3050
rect 86136 3084 86624 3090
rect 86136 3050 86148 3084
rect 86612 3050 86624 3084
rect 86136 3044 86624 3050
rect 84812 2936 84818 2996
rect 84878 2936 84884 2996
rect 84306 2882 84368 2888
rect 84306 2822 84308 2882
rect 84306 2816 84368 2822
rect 81760 2614 81766 2674
rect 81826 2614 81832 2674
rect 82282 2614 82288 2674
rect 82348 2614 82354 2674
rect 82782 2614 82788 2674
rect 82848 2614 82854 2674
rect 83290 2614 83296 2674
rect 83356 2614 83362 2674
rect 83798 2614 83804 2674
rect 83864 2614 83870 2674
rect 84148 2614 84154 2674
rect 84214 2614 84220 2674
rect 84306 2672 84366 2816
rect 85330 2778 85390 3044
rect 86332 2778 86392 3044
rect 86860 2996 86920 3134
rect 87878 3134 87890 3176
rect 87924 3176 87930 3710
rect 87924 3134 87938 3176
rect 87154 3084 87642 3090
rect 87154 3050 87166 3084
rect 87630 3050 87642 3084
rect 87154 3044 87642 3050
rect 87372 2996 87432 3044
rect 87878 2996 87938 3134
rect 86854 2936 86860 2996
rect 86920 2936 86926 2996
rect 87366 2936 87372 2996
rect 87432 2936 87438 2996
rect 87872 2936 87878 2996
rect 87938 2936 87944 2996
rect 85324 2718 85330 2778
rect 85390 2718 85396 2778
rect 86326 2718 86332 2778
rect 86392 2718 86398 2778
rect 81046 2560 81534 2566
rect 81046 2526 81058 2560
rect 81522 2526 81534 2560
rect 81046 2520 81534 2526
rect 78762 1966 78768 2442
rect 79734 2400 79746 2476
rect 78762 1900 78776 1966
rect 76974 1850 77462 1856
rect 76974 1816 76986 1850
rect 77450 1816 77462 1850
rect 76974 1810 77462 1816
rect 77992 1850 78480 1856
rect 77992 1816 78004 1850
rect 78468 1816 78480 1850
rect 77992 1810 78480 1816
rect 76674 1682 76680 1742
rect 76740 1682 76746 1742
rect 77182 1638 77242 1810
rect 78208 1638 78268 1810
rect 78716 1742 78776 1900
rect 79740 1900 79746 2400
rect 79780 2400 79794 2476
rect 80746 2426 80764 2476
rect 79780 1900 79786 2400
rect 80758 1932 80764 2426
rect 79740 1888 79786 1900
rect 80748 1900 80764 1932
rect 80798 2428 80810 2476
rect 81766 2476 81826 2614
rect 82288 2566 82348 2614
rect 82064 2560 82552 2566
rect 82064 2526 82076 2560
rect 82540 2526 82552 2560
rect 82064 2520 82552 2526
rect 82288 2514 82348 2520
rect 82788 2476 82848 2614
rect 83296 2566 83356 2614
rect 83082 2560 83570 2566
rect 83082 2526 83094 2560
rect 83558 2526 83570 2560
rect 83082 2520 83570 2526
rect 80798 2426 80806 2428
rect 80798 1932 80804 2426
rect 81766 2420 81782 2476
rect 80798 1900 80808 1932
rect 79010 1850 79498 1856
rect 79010 1816 79022 1850
rect 79486 1816 79498 1850
rect 79010 1810 79498 1816
rect 80028 1850 80516 1856
rect 80028 1816 80040 1850
rect 80504 1816 80516 1850
rect 80028 1810 80516 1816
rect 80236 1750 80296 1810
rect 80748 1750 80808 1900
rect 81776 1900 81782 2420
rect 81816 2420 81826 2476
rect 81816 1900 81822 2420
rect 82782 2416 82800 2476
rect 82794 1938 82800 2416
rect 82784 1900 82800 1938
rect 82834 2416 82848 2476
rect 83804 2476 83864 2614
rect 84154 2566 84214 2614
rect 84306 2612 84884 2672
rect 84100 2560 84588 2566
rect 84100 2526 84112 2560
rect 84576 2526 84588 2560
rect 84100 2520 84588 2526
rect 83804 2442 83818 2476
rect 82834 1938 82840 2416
rect 82834 1900 82844 1938
rect 83812 1900 83818 2442
rect 83852 2442 83864 2476
rect 84824 2476 84884 2612
rect 88044 2610 88104 3932
rect 85118 2560 85606 2566
rect 85118 2526 85130 2560
rect 85594 2526 85606 2560
rect 85118 2520 85606 2526
rect 86136 2560 86624 2566
rect 86136 2526 86148 2560
rect 86612 2526 86624 2560
rect 86136 2520 86624 2526
rect 87154 2560 87642 2566
rect 87154 2526 87166 2560
rect 87630 2526 87642 2560
rect 87154 2520 87642 2526
rect 87884 2550 88104 2610
rect 83852 1900 83858 2442
rect 84824 2438 84836 2476
rect 81776 1888 81822 1900
rect 82794 1888 82840 1900
rect 83812 1888 83858 1900
rect 84830 1900 84836 2438
rect 84870 2438 84884 2476
rect 85848 2476 85894 2488
rect 84870 1900 84876 2438
rect 85848 1932 85854 2476
rect 84830 1888 84876 1900
rect 85838 1900 85854 1932
rect 85888 1932 85894 2476
rect 86866 2476 86912 2488
rect 86866 1948 86872 2476
rect 85888 1900 85898 1932
rect 81046 1850 81534 1856
rect 81046 1816 81058 1850
rect 81522 1816 81534 1850
rect 81046 1810 81534 1816
rect 82064 1850 82552 1856
rect 82064 1816 82076 1850
rect 82540 1816 82552 1850
rect 82064 1810 82552 1816
rect 83082 1850 83570 1856
rect 83082 1816 83094 1850
rect 83558 1816 83570 1850
rect 83082 1810 83570 1816
rect 84100 1850 84588 1856
rect 84100 1816 84112 1850
rect 84576 1816 84588 1850
rect 84100 1810 84588 1816
rect 85118 1850 85606 1856
rect 85118 1816 85130 1850
rect 85594 1816 85606 1850
rect 85118 1810 85606 1816
rect 81254 1750 81314 1810
rect 78710 1682 78716 1742
rect 78776 1682 78782 1742
rect 80236 1690 81314 1750
rect 76170 1578 78268 1638
rect 70562 1482 70568 1542
rect 70628 1482 70634 1542
rect 72600 1482 72606 1542
rect 72666 1482 72672 1542
rect 74632 1482 74638 1542
rect 74698 1482 74704 1542
rect 76670 1482 76676 1542
rect 76736 1482 76742 1542
rect 78704 1482 78710 1542
rect 78770 1482 78776 1542
rect 80744 1482 80750 1542
rect 80810 1482 80816 1542
rect 82778 1482 82784 1542
rect 82844 1482 82850 1542
rect 84812 1482 84818 1542
rect 84878 1482 84884 1542
rect 69848 1328 70336 1334
rect 69848 1294 69860 1328
rect 70324 1294 70336 1328
rect 69848 1288 70336 1294
rect 68582 718 68588 1206
rect 69548 1196 69566 1244
rect 68582 668 68592 718
rect 67812 618 68300 624
rect 67812 584 67824 618
rect 68288 584 68300 618
rect 67812 578 68300 584
rect 68016 512 68076 578
rect 68532 512 68592 668
rect 69560 668 69566 1196
rect 69600 1196 69608 1244
rect 70568 1244 70628 1482
rect 71580 1384 71586 1444
rect 71646 1384 71652 1444
rect 70866 1328 71354 1334
rect 70866 1294 70878 1328
rect 71342 1294 71354 1328
rect 70866 1288 71354 1294
rect 70568 1212 70584 1244
rect 69600 668 69606 1196
rect 70578 696 70584 1212
rect 69560 656 69606 668
rect 70570 668 70584 696
rect 70618 1212 70628 1244
rect 71586 1244 71646 1384
rect 71884 1328 72372 1334
rect 71884 1294 71896 1328
rect 72360 1294 72372 1328
rect 71884 1288 72372 1294
rect 70618 696 70624 1212
rect 71586 1188 71602 1244
rect 70618 668 70630 696
rect 68830 618 69318 624
rect 68830 584 68842 618
rect 69306 584 69318 618
rect 68830 578 69318 584
rect 69848 618 70336 624
rect 69848 584 69860 618
rect 70324 584 70336 618
rect 69848 578 70336 584
rect 69064 512 69124 578
rect 70054 512 70114 578
rect 70570 512 70630 668
rect 71596 668 71602 1188
rect 71636 1188 71646 1244
rect 72606 1244 72666 1482
rect 73616 1384 73622 1444
rect 73682 1384 73688 1444
rect 72902 1328 73390 1334
rect 72902 1294 72914 1328
rect 73378 1294 73390 1328
rect 72902 1288 73390 1294
rect 72606 1198 72620 1244
rect 71636 668 71642 1188
rect 72614 696 72620 1198
rect 71596 656 71642 668
rect 72606 668 72620 696
rect 72654 1198 72666 1244
rect 73622 1244 73682 1384
rect 73920 1328 74408 1334
rect 73920 1294 73932 1328
rect 74396 1294 74408 1328
rect 73920 1288 74408 1294
rect 72654 696 72660 1198
rect 73622 1194 73638 1244
rect 72654 668 72666 696
rect 70866 618 71354 624
rect 70866 584 70878 618
rect 71342 584 71354 618
rect 70866 578 71354 584
rect 71884 618 72372 624
rect 71884 584 71896 618
rect 72360 584 72372 618
rect 71884 578 72372 584
rect 71076 512 71136 578
rect 72098 512 72158 578
rect 72606 512 72666 668
rect 73632 668 73638 1194
rect 73672 1194 73682 1244
rect 74638 1244 74698 1482
rect 75652 1384 75658 1444
rect 75718 1384 75724 1444
rect 74938 1328 75426 1334
rect 74938 1294 74950 1328
rect 75414 1294 75426 1328
rect 74938 1288 75426 1294
rect 73672 668 73678 1194
rect 74638 1188 74656 1244
rect 74650 702 74656 1188
rect 73632 656 73678 668
rect 74640 668 74656 702
rect 74690 1188 74698 1244
rect 75658 1244 75718 1384
rect 75956 1328 76444 1334
rect 75956 1294 75968 1328
rect 76432 1294 76444 1328
rect 75956 1288 76444 1294
rect 75658 1196 75674 1244
rect 74690 702 74696 1188
rect 74690 668 74700 702
rect 72902 618 73390 624
rect 72902 584 72914 618
rect 73378 584 73390 618
rect 72902 578 73390 584
rect 73920 618 74408 624
rect 73920 584 73932 618
rect 74396 584 74408 618
rect 73920 578 74408 584
rect 73120 512 73180 578
rect 74130 512 74190 578
rect 74640 512 74700 668
rect 75668 668 75674 1196
rect 75708 1196 75718 1244
rect 76676 1244 76736 1482
rect 77688 1384 77694 1444
rect 77754 1384 77760 1444
rect 76974 1328 77462 1334
rect 76974 1294 76986 1328
rect 77450 1294 77462 1328
rect 76974 1288 77462 1294
rect 76676 1200 76692 1244
rect 75708 668 75714 1196
rect 76686 726 76692 1200
rect 75668 656 75714 668
rect 76680 668 76692 726
rect 76726 1200 76736 1244
rect 77694 1244 77754 1384
rect 77992 1328 78480 1334
rect 77992 1294 78004 1328
rect 78468 1294 78480 1328
rect 77992 1288 78480 1294
rect 77694 1202 77710 1244
rect 76726 726 76732 1200
rect 76726 668 76740 726
rect 74938 618 75426 624
rect 74938 584 74950 618
rect 75414 584 75426 618
rect 74938 578 75426 584
rect 75956 618 76444 624
rect 75956 584 75968 618
rect 76432 584 76444 618
rect 75956 578 76444 584
rect 75158 512 75218 578
rect 76176 512 76236 578
rect 76680 512 76740 668
rect 77704 668 77710 1202
rect 77744 1202 77754 1244
rect 78710 1244 78770 1482
rect 79722 1384 79728 1444
rect 79788 1384 79794 1444
rect 79010 1328 79498 1334
rect 79010 1294 79022 1328
rect 79486 1294 79498 1328
rect 79010 1288 79498 1294
rect 77744 668 77750 1202
rect 78710 1188 78728 1244
rect 78722 698 78728 1188
rect 77704 656 77750 668
rect 78718 668 78728 698
rect 78762 1188 78770 1244
rect 79728 1244 79788 1384
rect 80028 1328 80516 1334
rect 80028 1294 80040 1328
rect 80504 1294 80516 1328
rect 80028 1288 80516 1294
rect 79728 1202 79746 1244
rect 78762 698 78768 1188
rect 78762 668 78778 698
rect 76974 618 77462 624
rect 76974 584 76986 618
rect 77450 584 77462 618
rect 76974 578 77462 584
rect 77992 618 78480 624
rect 77992 584 78004 618
rect 78468 584 78480 618
rect 77992 578 78480 584
rect 77192 512 77252 578
rect 78214 512 78274 578
rect 78718 512 78778 668
rect 79740 668 79746 1202
rect 79780 1202 79788 1244
rect 80750 1244 80810 1482
rect 81758 1384 81764 1444
rect 81824 1384 81830 1444
rect 81046 1328 81534 1334
rect 81046 1294 81058 1328
rect 81522 1294 81534 1328
rect 81046 1288 81534 1294
rect 79780 668 79786 1202
rect 80750 1198 80764 1244
rect 80758 712 80764 1198
rect 79740 656 79786 668
rect 80752 668 80764 712
rect 80798 1198 80810 1244
rect 81764 1244 81824 1384
rect 82064 1328 82552 1334
rect 82064 1294 82076 1328
rect 82540 1294 82552 1328
rect 82064 1288 82552 1294
rect 81764 1198 81782 1244
rect 80798 712 80804 1198
rect 80798 668 80812 712
rect 79010 618 79498 624
rect 79010 584 79022 618
rect 79486 584 79498 618
rect 79010 578 79498 584
rect 80028 618 80516 624
rect 80028 584 80040 618
rect 80504 584 80516 618
rect 80028 578 80516 584
rect 79236 512 79296 578
rect 80244 512 80304 578
rect 80752 512 80812 668
rect 81776 668 81782 1198
rect 81816 1198 81824 1244
rect 82784 1244 82844 1482
rect 83798 1384 83804 1444
rect 83864 1384 83870 1444
rect 83082 1328 83570 1334
rect 83082 1294 83094 1328
rect 83558 1294 83570 1328
rect 83082 1288 83570 1294
rect 81816 668 81822 1198
rect 82784 1186 82800 1244
rect 82794 708 82800 1186
rect 81776 656 81822 668
rect 82788 668 82800 708
rect 82834 1186 82844 1244
rect 83804 1244 83864 1384
rect 84100 1328 84588 1334
rect 84100 1294 84112 1328
rect 84576 1294 84588 1328
rect 84100 1288 84588 1294
rect 83804 1212 83818 1244
rect 82834 708 82840 1186
rect 82834 668 82848 708
rect 81248 624 81308 626
rect 81046 618 81534 624
rect 81046 584 81058 618
rect 81522 584 81534 618
rect 81046 578 81534 584
rect 82064 618 82552 624
rect 82064 584 82076 618
rect 82540 584 82552 618
rect 82064 578 82552 584
rect 81248 512 81308 578
rect 82294 512 82354 578
rect 82788 512 82848 668
rect 83812 668 83818 1212
rect 83852 1212 83864 1244
rect 84818 1244 84878 1482
rect 85316 1334 85376 1810
rect 85838 1444 85898 1900
rect 86856 1900 86872 1948
rect 86906 1948 86912 2476
rect 87884 2476 87944 2550
rect 86906 1900 86916 1948
rect 87884 1934 87890 2476
rect 86136 1850 86624 1856
rect 86136 1816 86148 1850
rect 86612 1816 86624 1850
rect 86136 1810 86624 1816
rect 85832 1384 85838 1444
rect 85898 1384 85904 1444
rect 85118 1328 85606 1334
rect 85118 1294 85130 1328
rect 85594 1294 85606 1328
rect 85118 1288 85606 1294
rect 83852 668 83858 1212
rect 84818 1202 84836 1244
rect 84830 702 84836 1202
rect 83812 656 83858 668
rect 84826 668 84836 702
rect 84870 1202 84878 1244
rect 85838 1244 85898 1384
rect 86344 1334 86404 1810
rect 86856 1542 86916 1900
rect 87874 1900 87890 1934
rect 87924 2400 87944 2476
rect 87924 1934 87930 2400
rect 87924 1900 87934 1934
rect 87154 1850 87642 1856
rect 87154 1816 87166 1850
rect 87630 1816 87642 1850
rect 87154 1810 87642 1816
rect 86850 1482 86856 1542
rect 86916 1482 86922 1542
rect 86136 1328 86624 1334
rect 86136 1294 86148 1328
rect 86612 1294 86624 1328
rect 86136 1288 86624 1294
rect 85838 1204 85854 1244
rect 84870 702 84876 1202
rect 84870 668 84886 702
rect 83082 618 83570 624
rect 83082 584 83094 618
rect 83558 584 83570 618
rect 83082 578 83570 584
rect 84100 618 84588 624
rect 84100 584 84112 618
rect 84576 584 84588 618
rect 84100 578 84588 584
rect 83292 512 83352 578
rect 84304 512 84364 578
rect 84826 512 84886 668
rect 85848 668 85854 1204
rect 85888 1204 85898 1244
rect 86856 1244 86916 1482
rect 87336 1334 87396 1810
rect 87874 1444 87934 1900
rect 88598 1542 88658 13934
rect 88750 2614 88756 2674
rect 88816 2614 88822 2674
rect 88592 1482 88598 1542
rect 88658 1482 88664 1542
rect 87868 1384 87874 1444
rect 87934 1384 87940 1444
rect 87154 1328 87642 1334
rect 87154 1294 87166 1328
rect 87630 1294 87642 1328
rect 87154 1288 87642 1294
rect 87336 1286 87396 1288
rect 86856 1214 86872 1244
rect 85888 668 85894 1204
rect 86866 696 86872 1214
rect 85848 656 85894 668
rect 86854 668 86872 696
rect 86906 1214 86916 1244
rect 87874 1244 87934 1384
rect 86906 696 86912 1214
rect 87874 1208 87890 1244
rect 86906 668 86914 696
rect 85118 618 85606 624
rect 85118 584 85130 618
rect 85594 584 85606 618
rect 85118 578 85606 584
rect 86136 618 86624 624
rect 86136 584 86148 618
rect 86612 584 86624 618
rect 86136 578 86624 584
rect 85326 512 85386 578
rect 86392 512 86452 578
rect 86854 512 86914 668
rect 87884 668 87890 1208
rect 87924 1208 87934 1244
rect 87924 668 87930 1208
rect 87884 656 87930 668
rect 87154 618 87642 624
rect 87154 584 87166 618
rect 87630 584 87642 618
rect 87154 578 87642 584
rect 87354 512 87414 578
rect 68016 452 87414 512
rect 88756 110 88816 2614
rect 89766 210 89772 14470
rect 89872 210 89878 14470
rect 57432 64 88918 110
rect 57432 -90 57478 64
rect 88878 -90 88918 64
rect 57432 -136 88918 -90
rect 53334 -576 53344 -276
rect 89156 -576 89166 -276
rect 89766 -576 89878 210
rect 52622 -582 89878 -576
rect 52622 -682 52728 -582
rect 89772 -682 89878 -582
rect 52622 -688 89878 -682
<< via1 >>
rect -1414 27582 -1354 27642
rect 11434 27856 12034 28156
rect 35066 27856 35666 28156
rect 15011 27560 31796 27774
rect 15106 21978 15166 22038
rect 15218 21978 15278 22038
rect 15328 21978 15388 22038
rect 14442 21266 14502 21326
rect 14782 21266 14842 21326
rect 14892 21266 14952 21326
rect 13060 20320 13120 20380
rect 15978 21978 16038 22038
rect 16088 21978 16148 22038
rect 16196 21978 16256 22038
rect 15542 21266 15602 21326
rect 15654 21266 15714 21326
rect 15762 21266 15822 21326
rect 18936 27364 18996 27424
rect 20018 27364 20078 27424
rect 20976 27364 21036 27424
rect 19462 27118 19522 27178
rect 22012 27364 22072 27424
rect 23018 27364 23078 27424
rect 21498 27118 21558 27178
rect 17280 26186 17340 26246
rect 18444 26186 18504 26246
rect 17150 25982 17210 26042
rect 18444 25982 18504 26042
rect 22516 27230 22576 27290
rect 24040 27364 24100 27424
rect 25058 27364 25118 27424
rect 23536 27120 23596 27180
rect 20480 26082 20540 26142
rect 26082 27364 26142 27424
rect 27094 27364 27154 27424
rect 25566 27120 25626 27180
rect 22516 26082 22576 26142
rect 19460 25048 19520 25108
rect 28112 27364 28172 27424
rect 29124 27364 29184 27424
rect 27608 27122 27668 27182
rect 24554 26186 24614 26246
rect 24550 25982 24610 26042
rect 21496 25048 21556 25108
rect 20478 24952 20538 25012
rect 21182 24946 21246 25010
rect 22354 24946 22418 25010
rect 22516 24842 22576 24902
rect 19460 23910 19520 23970
rect 28620 27230 28680 27290
rect 30152 27364 30212 27424
rect 31164 27364 31224 27424
rect 29640 27122 29700 27182
rect 26588 26186 26648 26246
rect 26586 25982 26646 26042
rect 23530 25048 23590 25108
rect 20476 23796 20540 23860
rect 18438 23658 18502 23722
rect 17280 23512 17340 23572
rect 18262 23512 18322 23572
rect 17866 23176 17926 23236
rect 16998 21978 17058 22038
rect 16414 21266 16474 21326
rect 16524 21266 16584 21326
rect 14998 21160 15058 21220
rect 15434 21160 15494 21220
rect 15872 21160 15932 21220
rect 16306 21160 16366 21220
rect 15218 21044 15278 21104
rect 14782 20320 14842 20380
rect 14998 20216 15058 20276
rect 14892 20118 14952 20178
rect 15216 20320 15276 20380
rect 15106 20118 15166 20178
rect 14442 19482 14502 19542
rect 16088 21044 16148 21104
rect 15434 20216 15494 20276
rect 15326 20118 15386 20178
rect 14782 19382 14842 19442
rect 15652 20320 15712 20380
rect 15872 20216 15932 20276
rect 15544 20118 15604 20178
rect 15654 20118 15714 20178
rect 15760 20118 15820 20178
rect 16088 20320 16148 20380
rect 15978 20118 16038 20178
rect 16882 21044 16942 21104
rect 16306 20216 16366 20276
rect 16196 20118 16256 20178
rect 15652 19382 15712 19442
rect 16526 20320 16586 20380
rect 16412 20118 16472 20178
rect 16526 19382 16586 19442
rect 16882 19382 16942 19442
rect 14998 19284 15058 19344
rect 15434 19284 15494 19344
rect 15872 19284 15932 19344
rect 16306 19284 16366 19344
rect 14442 19166 14502 19226
rect 15108 19166 15168 19226
rect 15216 19166 15276 19226
rect 15324 19166 15384 19226
rect 15970 19166 16030 19226
rect 16088 19166 16148 19226
rect 16197 19166 16255 19224
rect 17752 20872 17812 20932
rect 32182 27364 32242 27424
rect 31676 27122 31736 27182
rect 28622 26082 28682 26142
rect 25568 25046 25628 25106
rect 21496 23910 21556 23970
rect 20476 23362 20540 23426
rect 18262 23076 18322 23136
rect 19428 23076 19488 23136
rect 17994 22030 18054 22090
rect 17866 20768 17926 20828
rect 14782 18446 14842 18506
rect 14892 18446 14952 18506
rect 15546 18446 15606 18506
rect 15652 18446 15712 18506
rect 15762 18446 15822 18506
rect 16414 18446 16474 18506
rect 16526 18446 16586 18506
rect 16998 18446 17058 18506
rect 18130 21932 18190 21992
rect 17994 18358 18054 18418
rect 28764 25978 28824 26038
rect 26588 24948 26648 25008
rect 30656 26082 30716 26142
rect 30658 25978 30718 26038
rect 27604 25046 27664 25106
rect 22990 23906 23050 23966
rect 22514 23176 22574 23236
rect 21464 23076 21524 23136
rect 23530 23968 23590 23970
rect 23498 23910 23590 23968
rect 23990 23910 24050 23970
rect 23498 23908 23558 23910
rect 19432 21822 19492 21882
rect 28622 24842 28682 24902
rect 25034 23912 25094 23972
rect 24548 23658 24612 23722
rect 24548 23374 24612 23438
rect 25536 23968 25596 23972
rect 25536 23912 25628 23968
rect 25568 23908 25628 23912
rect 26050 23912 26110 23972
rect 20446 22128 20506 22188
rect 20446 21932 20506 21992
rect 21466 21934 21526 21994
rect 21466 21822 21526 21882
rect 32696 26186 32756 26246
rect 33834 26186 33894 26246
rect 29640 25046 29700 25106
rect 30658 24842 30718 24902
rect 31674 25044 31734 25104
rect 27078 23912 27138 23972
rect 26584 23658 26648 23722
rect 27604 23966 27664 23968
rect 27572 23908 27664 23966
rect 27572 23906 27632 23908
rect 28100 23902 28160 23962
rect 28588 23906 28648 23966
rect 32696 24948 32756 25008
rect 29100 23902 29160 23962
rect 29640 23906 29700 23966
rect 31674 23906 31734 23966
rect 30656 23796 30720 23860
rect 32692 23658 32756 23722
rect 32664 23382 32724 23442
rect 33834 23376 33894 23436
rect 29610 23076 29670 23136
rect 31644 23076 31704 23136
rect 22482 22128 22542 22188
rect 24522 21820 24582 21880
rect 20448 20768 20508 20828
rect 20448 20564 20508 20624
rect 26556 21820 26616 21880
rect 22484 20768 22544 20828
rect 22482 20666 22542 20726
rect 22482 20564 22542 20624
rect 19430 19616 19490 19676
rect 18262 19408 18322 19468
rect 20444 19306 20504 19366
rect 24518 20872 24578 20932
rect 25538 20872 25598 20932
rect 25538 20566 25598 20626
rect 21466 19616 21526 19676
rect 21466 19508 21526 19568
rect 29612 21820 29672 21880
rect 26556 20566 26616 20626
rect 34088 23076 34148 23136
rect 30626 22128 30686 22188
rect 31646 21820 31706 21880
rect 32662 22128 32722 22188
rect 33928 21934 33988 21994
rect 27574 20872 27634 20932
rect 27572 20566 27632 20626
rect 22478 19306 22538 19366
rect 22682 19312 22742 19372
rect 19426 18358 19486 18418
rect 24520 19618 24580 19678
rect 29608 20768 29668 20828
rect 30476 20886 30536 20946
rect 30624 20776 30684 20836
rect 30476 20566 30536 20626
rect 30628 20568 30688 20628
rect 26556 19618 26616 19678
rect 31644 20666 31704 20726
rect 32664 20776 32724 20836
rect 33796 20776 33856 20836
rect 32662 20568 32722 20628
rect 24516 19312 24576 19372
rect 25536 19308 25596 19368
rect 27570 19308 27630 19368
rect 21462 18358 21522 18418
rect 18130 18228 18190 18288
rect 13060 18088 13120 18148
rect 12904 17982 12964 18042
rect 27784 19304 27844 19364
rect 29610 19620 29670 19680
rect 30120 19304 30180 19364
rect 30632 19306 30692 19366
rect 31646 19620 31706 19680
rect 33928 20568 33988 20628
rect 33796 19508 33856 19568
rect 32666 19306 32726 19366
rect 29614 18358 29674 18418
rect 31650 18358 31710 18418
rect 22484 18088 22544 18148
rect 47824 27564 48000 27680
rect 48306 27564 48462 27680
rect 65434 27856 66034 28156
rect 89066 27856 89666 28156
rect 48528 25370 48588 25430
rect 47880 24604 47940 24664
rect 47622 24455 47682 24515
rect 48398 24604 48458 24664
rect 48138 24455 48198 24515
rect 49201 24586 49261 24592
rect 49201 24538 49207 24586
rect 49207 24538 49255 24586
rect 49255 24538 49261 24586
rect 49201 24532 49261 24538
rect 49519 24554 49579 24614
rect 48656 24455 48716 24515
rect 47250 23874 47310 23934
rect 48526 23907 48586 23967
rect 48528 23370 48588 23430
rect 47880 22604 47940 22664
rect 47622 22455 47682 22515
rect 48398 22604 48458 22664
rect 48138 22455 48198 22515
rect 49201 22586 49261 22592
rect 49201 22538 49207 22586
rect 49207 22538 49255 22586
rect 49255 22538 49261 22586
rect 49201 22532 49261 22538
rect 49519 22554 49579 22614
rect 48656 22455 48716 22515
rect 46978 21860 47038 21920
rect 48526 21907 48586 21967
rect 34088 18088 34148 18148
rect 12134 17864 12194 17924
rect -8742 16348 -8682 16408
rect -1414 16348 -1354 16408
rect -11830 16240 -11770 16300
rect -12478 15474 -12418 15534
rect -12736 15325 -12676 15385
rect -11960 15474 -11900 15534
rect -12220 15325 -12160 15385
rect -9230 16240 -9170 16300
rect -11157 15456 -11097 15462
rect -11157 15408 -11151 15456
rect -11151 15408 -11103 15456
rect -11103 15408 -11097 15456
rect -11157 15402 -11097 15408
rect -10839 15424 -10779 15484
rect -9878 15474 -9818 15534
rect -11702 15325 -11642 15385
rect -12478 14896 -12418 14956
rect -10136 15325 -10076 15385
rect -11832 14777 -11772 14837
rect -9360 15474 -9300 15534
rect -9620 15325 -9560 15385
rect -8557 15456 -8497 15462
rect -8557 15408 -8551 15456
rect -8551 15408 -8503 15456
rect -8503 15408 -8497 15456
rect -8557 15402 -8497 15408
rect -8239 15424 -8179 15484
rect -9102 15325 -9042 15385
rect 5912 15362 6012 15364
rect 8512 15362 8612 15364
rect 10316 15362 10416 15364
rect -9878 14892 -9818 14952
rect -1082 15262 -982 15362
rect 712 15262 812 15362
rect 3312 15262 3412 15362
rect 5912 15264 6012 15362
rect 8512 15264 8612 15362
rect 10316 15264 10416 15362
rect -10006 14777 -9946 14837
rect -9232 14777 -9172 14837
rect 12904 15132 12964 15192
rect 13060 15132 13120 15192
rect -8750 14652 -8690 14712
rect -1792 14652 -1732 14712
rect 12134 14146 12194 14206
rect 12800 14032 12860 14092
rect 13286 15124 13346 15184
rect 13062 12692 13122 12752
rect 12926 12480 12986 12540
rect 12800 11578 12860 11638
rect 11640 7592 11700 7652
rect 7974 6320 8034 6380
rect 3564 4880 3624 4940
rect 5604 4880 5664 4940
rect 1412 3976 1472 4036
rect 2550 3976 2610 4036
rect 3564 3880 3624 3940
rect 4586 3764 4646 3824
rect 5604 3880 5664 3940
rect 2696 2864 2756 2924
rect 2548 2756 2608 2816
rect 6624 3976 6684 4036
rect 10136 7356 10196 7416
rect 11048 7356 11108 7416
rect 9266 7246 9326 7306
rect 8352 7138 8412 7198
rect 8482 7030 8542 7090
rect 10030 7138 10090 7198
rect 9812 7030 9872 7090
rect 8940 6530 9000 6590
rect 9048 6430 9108 6490
rect 9050 6320 9110 6380
rect 9596 6530 9656 6590
rect 9486 6430 9546 6490
rect 9484 6320 9544 6380
rect 9158 6210 9218 6270
rect 9378 6210 9438 6270
rect 8482 5706 8542 5766
rect 8352 5584 8412 5644
rect 8940 5706 9000 5766
rect 9158 5584 9218 5644
rect 8832 5460 8892 5520
rect 10928 7246 10988 7306
rect 10248 7138 10308 7198
rect 10466 7030 10526 7090
rect 10466 6530 10526 6590
rect 9812 6320 9872 6380
rect 9922 6320 9982 6380
rect 10358 6320 10418 6380
rect 10032 6210 10092 6270
rect 10248 6210 10308 6270
rect 9596 5706 9656 5766
rect 9376 5584 9436 5644
rect 9270 5334 9330 5394
rect 10928 6756 10988 6816
rect 10576 6410 10636 6470
rect 10140 5706 10200 5766
rect 9812 5586 9872 5646
rect 10468 5586 10528 5646
rect 10928 5706 10988 5766
rect 9702 5460 9762 5520
rect 10574 5460 10634 5520
rect 11170 6530 11230 6590
rect 11170 6284 11230 6344
rect 11048 5334 11108 5394
rect 9604 5228 9656 5280
rect 8280 5144 8340 5204
rect 11902 7622 11962 7682
rect 8280 4900 8340 4960
rect 3566 2644 3626 2704
rect 7748 3764 7808 3824
rect 4582 2864 4642 2924
rect 4584 2756 4644 2816
rect 5604 2644 5664 2704
rect 2550 1660 2610 1720
rect 1412 1554 1472 1614
rect 6452 2864 6512 2924
rect 6620 2756 6680 2816
rect 3568 1762 3628 1822
rect 4584 1554 4644 1614
rect 5598 1762 5658 1822
rect 3054 610 3114 670
rect 8828 5000 8888 5060
rect 10018 5000 10078 5060
rect 11212 5000 11272 5060
rect 11902 5000 11962 5060
rect 9272 4900 9332 4960
rect 9570 4900 9630 4960
rect 8408 3866 8468 3926
rect 8824 3866 8884 3926
rect 10466 4900 10526 4960
rect 10762 4900 10822 4960
rect 9121 3999 9179 4057
rect 8976 3758 9036 3818
rect 9725 3999 9783 4057
rect 9418 3866 9478 3926
rect 9274 3758 9334 3818
rect 9574 3758 9634 3818
rect 8280 2860 8340 2920
rect 6618 1660 6678 1720
rect 7748 1660 7808 1720
rect 4080 610 4140 670
rect 5104 610 5164 670
rect 8974 2860 9034 2920
rect 10016 3866 10076 3926
rect 9868 3758 9928 3818
rect 10316 3999 10374 4057
rect 10164 3758 10224 3818
rect 10913 3999 10971 4057
rect 10610 3866 10670 3926
rect 10464 3758 10524 3818
rect 10766 3758 10826 3818
rect 9420 2752 9480 2812
rect 11208 3866 11268 3926
rect 11056 3758 11116 3818
rect 11509 3999 11567 4057
rect 11360 3758 11420 3818
rect 9870 2860 9930 2920
rect 10164 2860 10224 2920
rect 10614 2752 10674 2812
rect 9122 1768 9182 1828
rect 8524 1674 8584 1734
rect 8972 1566 9032 1626
rect 9416 1674 9476 1734
rect 9270 1566 9330 1626
rect 9716 1768 9776 1828
rect 9566 1566 9626 1626
rect 11058 2860 11118 2920
rect 11360 2860 11420 2920
rect 10316 1768 10376 1828
rect 10014 1674 10074 1734
rect 9870 1566 9930 1626
rect 10166 1566 10226 1626
rect 10612 1674 10672 1734
rect 10464 1566 10524 1626
rect 11902 2752 11962 2812
rect 10910 1768 10970 1828
rect 10760 1566 10820 1626
rect 11504 1768 11564 1828
rect 11212 1674 11272 1734
rect 11056 1566 11116 1626
rect 11360 1566 11420 1626
rect 6004 610 6064 670
rect 8280 640 8340 700
rect 9270 640 9330 700
rect 9568 640 9628 700
rect 10464 640 10524 700
rect 10766 640 10826 700
rect 12026 3758 12086 3818
rect 12926 2936 12986 2996
rect 13518 14032 13578 14092
rect 14536 13934 14596 13994
rect 15554 14032 15614 14092
rect 17588 14032 17648 14092
rect 19628 14032 19688 14092
rect 21664 14032 21724 14092
rect 23698 14032 23758 14092
rect 25734 14032 25794 14092
rect 27770 14032 27830 14092
rect 29806 14032 29866 14092
rect 16574 13934 16634 13994
rect 18608 13934 18668 13994
rect 20642 13934 20702 13994
rect 22682 13934 22742 13994
rect 24716 13934 24776 13994
rect 26754 13934 26814 13994
rect 28786 13934 28846 13994
rect 30824 13934 30884 13994
rect 22682 13722 22742 13782
rect 24714 13722 24774 13782
rect 17222 12802 17282 12862
rect 17592 12802 17652 12862
rect 18094 12802 18154 12862
rect 18606 12802 18666 12862
rect 19134 12802 19194 12862
rect 19626 12802 19686 12862
rect 15046 12692 15106 12752
rect 16068 12692 16128 12752
rect 13522 12480 13582 12540
rect 14020 12480 14080 12540
rect 14532 12480 14592 12540
rect 17088 12588 17148 12648
rect 16574 12480 16634 12540
rect 15036 11578 15096 11638
rect 13286 11364 13346 11424
rect 18088 12588 18148 12648
rect 19108 12588 19168 12648
rect 18608 12480 18668 12540
rect 16052 11590 16112 11650
rect 17072 11590 17132 11650
rect 15548 11486 15608 11546
rect 15554 11252 15614 11312
rect 16572 11486 16632 11546
rect 21658 12802 21718 12862
rect 20140 12692 20200 12752
rect 20644 12692 20704 12752
rect 21160 12692 21220 12752
rect 20642 12480 20702 12540
rect 18084 11590 18144 11650
rect 19110 11590 19170 11650
rect 17584 11486 17644 11546
rect 17590 11252 17650 11312
rect 18604 11486 18664 11546
rect 13398 10322 13458 10382
rect 14536 10322 14596 10382
rect 13286 10122 13346 10182
rect 13180 10020 13240 10080
rect 13286 8886 13346 8946
rect 13180 6530 13240 6590
rect 14534 10122 14594 10182
rect 15552 10242 15612 10302
rect 22180 12692 22240 12752
rect 22682 12692 22742 12752
rect 23182 12692 23242 12752
rect 22798 12480 22858 12540
rect 23694 12802 23754 12862
rect 23322 12588 23382 12648
rect 24208 12692 24268 12752
rect 24330 12588 24390 12648
rect 24718 12692 24778 12752
rect 25226 12692 25286 12752
rect 24522 12478 24582 12538
rect 25730 12802 25790 12862
rect 25372 12588 25432 12648
rect 27768 12802 27828 12862
rect 26234 12692 26294 12752
rect 26756 12692 26816 12752
rect 27246 12692 27306 12752
rect 26756 12480 26816 12540
rect 31844 14032 31904 14092
rect 32862 13934 32922 13994
rect 33874 14032 33934 14092
rect 34598 13934 34658 13994
rect 29292 12802 29352 12862
rect 29806 12802 29866 12862
rect 30314 12802 30374 12862
rect 28278 12692 28338 12752
rect 28790 12692 28850 12752
rect 28264 12588 28324 12648
rect 29302 12588 29362 12648
rect 28788 12480 28848 12540
rect 19626 11486 19686 11546
rect 21662 11486 21722 11546
rect 23700 11486 23760 11546
rect 25730 11486 25790 11546
rect 20646 11364 20706 11424
rect 22680 11364 22740 11424
rect 24710 11364 24770 11424
rect 16570 10346 16630 10406
rect 16066 10128 16126 10188
rect 17592 10242 17652 10302
rect 17070 10128 17130 10188
rect 14534 9090 14594 9150
rect 15040 8988 15100 9048
rect 18606 10346 18666 10406
rect 18082 10128 18142 10188
rect 19624 10242 19684 10302
rect 26750 11486 26810 11546
rect 19102 10128 19162 10188
rect 19624 10130 19684 10190
rect 21658 10242 21718 10302
rect 20642 10020 20702 10080
rect 16572 9090 16632 9150
rect 16570 8886 16630 8946
rect 21660 10130 21720 10190
rect 22676 10020 22736 10080
rect 31334 12692 31394 12752
rect 32354 12692 32414 12752
rect 30302 12588 30362 12648
rect 30820 12480 30880 12540
rect 32862 12480 32922 12540
rect 33366 12480 33426 12540
rect 33876 12480 33936 12540
rect 28266 11590 28326 11650
rect 29302 11590 29362 11650
rect 27768 11486 27828 11546
rect 28788 11486 28848 11546
rect 23698 10242 23758 10302
rect 23696 10130 23756 10190
rect 25732 10242 25792 10302
rect 25928 10238 25988 10298
rect 24716 10020 24776 10080
rect 25732 10130 25792 10190
rect 30318 11590 30378 11650
rect 29804 11486 29864 11546
rect 31840 11486 31900 11546
rect 26750 10346 26810 10406
rect 25928 10020 25988 10080
rect 26222 10022 26282 10082
rect 18608 9090 18668 9150
rect 15554 8786 15614 8846
rect 17078 8880 17138 8940
rect 18100 8880 18160 8940
rect 17588 8786 17648 8846
rect 20640 9090 20700 9150
rect 20132 8988 20192 9048
rect 19114 8880 19174 8940
rect 20132 8880 20192 8940
rect 19624 8786 19684 8846
rect 15036 7862 15096 7922
rect 15946 7862 16006 7922
rect 15036 7646 15096 7706
rect 13400 7542 13460 7602
rect 13286 6284 13346 6344
rect 13192 5228 13244 5280
rect 16948 7862 17008 7922
rect 16074 7646 16134 7706
rect 18100 7862 18160 7922
rect 17588 7760 17648 7820
rect 17088 7646 17148 7706
rect 15034 6634 15094 6694
rect 14536 6530 14596 6590
rect 14532 6320 14592 6380
rect 16042 6634 16102 6694
rect 15552 6418 15612 6478
rect 21152 8880 21212 8940
rect 27766 10130 27826 10190
rect 27250 10022 27310 10082
rect 27768 10016 27828 10076
rect 28786 10346 28846 10406
rect 29804 10130 29864 10190
rect 30820 10238 30880 10298
rect 31324 10234 31384 10294
rect 33984 11252 34044 11312
rect 31844 10130 31904 10190
rect 29804 10016 29864 10076
rect 25222 9102 25282 9162
rect 24716 8974 24776 9034
rect 26752 8776 26812 8836
rect 19110 7862 19170 7922
rect 20116 7862 20176 7922
rect 21160 7862 21220 7922
rect 21660 7868 21720 7928
rect 20114 7646 20174 7706
rect 21154 7646 21214 7706
rect 20638 7542 20698 7602
rect 17056 6634 17116 6694
rect 18094 6634 18154 6694
rect 17590 6418 17650 6478
rect 16570 6320 16630 6380
rect 22168 7646 22228 7706
rect 23696 7868 23756 7928
rect 23176 7646 23236 7706
rect 24220 7646 24280 7706
rect 22680 7542 22740 7602
rect 31842 10016 31902 10076
rect 28264 8880 28324 8940
rect 25732 7868 25792 7928
rect 25210 7646 25270 7706
rect 26228 7646 26288 7706
rect 24718 7542 24778 7602
rect 32860 10346 32920 10406
rect 33878 10364 33938 10424
rect 34478 10234 34538 10294
rect 34228 10130 34288 10190
rect 30316 9102 30376 9162
rect 30454 9106 30514 9166
rect 33984 10016 34044 10076
rect 31336 9106 31396 9166
rect 32342 9106 32402 9166
rect 29294 8880 29354 8940
rect 30454 8880 30514 8940
rect 30822 8880 30882 8940
rect 30822 8776 30882 8836
rect 32860 9102 32920 9162
rect 32860 8974 32920 9034
rect 31838 8778 31898 8838
rect 27770 7868 27830 7928
rect 27762 7760 27822 7820
rect 27262 7646 27322 7706
rect 26752 7542 26812 7602
rect 27264 7538 27324 7598
rect 28286 7538 28346 7598
rect 28786 7544 28846 7604
rect 19112 6634 19172 6694
rect 19628 6640 19688 6700
rect 21664 6640 21724 6700
rect 23696 6640 23756 6700
rect 25730 6640 25790 6700
rect 18610 6320 18670 6380
rect 13398 5298 13458 5358
rect 14538 5082 14598 5142
rect 15552 5396 15612 5456
rect 15556 5202 15616 5262
rect 16570 5298 16630 5358
rect 22680 6530 22740 6590
rect 24716 6530 24776 6590
rect 21662 6418 21722 6478
rect 20646 6320 20706 6380
rect 17588 5396 17648 5456
rect 18094 5298 18154 5358
rect 17592 5202 17652 5262
rect 19626 5396 19686 5456
rect 19116 5298 19176 5358
rect 18606 5082 18666 5142
rect 13286 4166 13346 4226
rect 20138 5298 20198 5358
rect 19620 5202 19680 5262
rect 29806 7868 29866 7928
rect 29802 7760 29862 7820
rect 30294 7646 30354 7706
rect 31844 7868 31904 7928
rect 31840 7760 31900 7820
rect 31332 7646 31392 7706
rect 30820 7544 30880 7604
rect 26752 6642 26812 6702
rect 27106 6642 27166 6702
rect 26748 6530 26808 6590
rect 26258 6432 26318 6492
rect 21488 5416 21548 5476
rect 21658 5416 21718 5476
rect 21142 5298 21202 5358
rect 20640 5082 20700 5142
rect 13180 4040 13240 4100
rect 16570 4040 16630 4100
rect 17090 4052 17150 4112
rect 15552 3930 15612 3990
rect 17588 3930 17648 3990
rect 17206 3836 17266 3896
rect 21488 5202 21548 5262
rect 21664 5208 21724 5268
rect 27296 6432 27356 6492
rect 28272 6432 28332 6492
rect 27106 6324 27166 6384
rect 32358 7646 32418 7706
rect 32862 7544 32922 7604
rect 30824 6642 30884 6702
rect 29288 6432 29348 6492
rect 31314 6432 31374 6492
rect 28786 6320 28846 6380
rect 30822 6320 30882 6380
rect 23700 5416 23760 5476
rect 25732 5416 25792 5476
rect 27772 5416 27832 5476
rect 26750 5318 26810 5378
rect 23692 5208 23752 5268
rect 18608 3930 18668 3990
rect 25736 5208 25796 5268
rect 19624 3930 19684 3990
rect 20644 3930 20704 3990
rect 18090 3836 18150 3896
rect 19112 3836 19172 3896
rect 13518 2936 13578 2996
rect 14032 2936 14092 2996
rect 14530 2936 14590 2996
rect 16572 2936 16632 2996
rect 17080 2824 17140 2884
rect 13060 2718 13120 2778
rect 15046 2718 15106 2778
rect 16068 2718 16128 2778
rect 27764 5208 27824 5268
rect 28790 5082 28850 5142
rect 32344 6432 32404 6492
rect 32858 6320 32918 6380
rect 29802 5208 29862 5268
rect 32856 5318 32916 5378
rect 31842 5208 31902 5268
rect 32360 5212 32420 5272
rect 30820 5082 30880 5142
rect 31346 5084 31406 5144
rect 22674 4166 22734 4226
rect 24716 4166 24776 4226
rect 26752 4166 26812 4226
rect 22170 4052 22230 4112
rect 27258 4056 27318 4116
rect 21662 3930 21722 3990
rect 23692 3930 23752 3990
rect 25730 3930 25790 3990
rect 27766 3930 27826 3990
rect 21154 3836 21214 3896
rect 18604 2936 18664 2996
rect 18092 2824 18152 2884
rect 19106 2824 19166 2884
rect 18606 2718 18666 2778
rect 19118 2718 19178 2778
rect 12654 2614 12714 2674
rect 17082 2614 17142 2674
rect 17586 2614 17646 2674
rect 18102 2614 18162 2674
rect 12026 1566 12086 1626
rect 8824 540 8884 600
rect 10012 540 10072 600
rect 11208 540 11268 600
rect 11902 540 11962 600
rect 13518 1384 13578 1444
rect 14530 1482 14590 1542
rect 20636 2936 20696 2996
rect 20136 2718 20196 2778
rect 20642 2718 20702 2778
rect 21148 2718 21208 2778
rect 19624 2614 19684 2674
rect 15548 1384 15608 1444
rect 22018 2824 22078 2884
rect 21662 2614 21722 2674
rect 22540 2936 22600 2996
rect 22160 2718 22220 2778
rect 22678 2826 22738 2886
rect 23306 2822 23366 2882
rect 23180 2718 23240 2778
rect 24352 2822 24412 2882
rect 24202 2718 24262 2778
rect 23698 2614 23758 2674
rect 24900 2938 24960 2998
rect 24714 2718 24774 2778
rect 25220 2718 25280 2778
rect 32858 5084 32918 5144
rect 28788 3930 28848 3990
rect 29806 4166 29866 4226
rect 29808 3930 29868 3990
rect 28276 3836 28336 3896
rect 29296 3836 29356 3896
rect 26750 2936 26810 2996
rect 26238 2718 26298 2778
rect 26750 2718 26810 2778
rect 27258 2718 27318 2778
rect 25734 2614 25794 2674
rect 30822 3930 30882 3990
rect 31838 4166 31898 4226
rect 34112 9102 34172 9162
rect 34350 8880 34410 8940
rect 34228 8778 34288 8838
rect 34112 7544 34172 7604
rect 34108 6642 34168 6702
rect 34228 5416 34288 5476
rect 34108 5318 34168 5378
rect 34476 7646 34536 7706
rect 34478 5212 34538 5272
rect 34350 5084 34410 5144
rect 33984 4166 34044 4226
rect 32358 4056 32418 4116
rect 31844 3930 31904 3990
rect 30310 3836 30370 3896
rect 31346 3836 31406 3896
rect 28784 2936 28844 2996
rect 28280 2822 28340 2882
rect 29298 2822 29358 2882
rect 30818 2936 30878 2996
rect 30308 2822 30368 2882
rect 27766 2614 27826 2674
rect 28288 2614 28348 2674
rect 28788 2614 28848 2674
rect 29296 2614 29356 2674
rect 29804 2614 29864 2674
rect 30154 2614 30214 2674
rect 32860 2936 32920 2996
rect 33372 2936 33432 2996
rect 33878 2936 33938 2996
rect 31330 2718 31390 2778
rect 32332 2718 32392 2778
rect 22680 1682 22740 1742
rect 24716 1682 24776 1742
rect 16568 1482 16628 1542
rect 18606 1482 18666 1542
rect 20638 1482 20698 1542
rect 22676 1482 22736 1542
rect 24710 1482 24770 1542
rect 26750 1482 26810 1542
rect 28784 1482 28844 1542
rect 30818 1482 30878 1542
rect 17586 1384 17646 1444
rect 19622 1384 19682 1444
rect 21658 1384 21718 1444
rect 23694 1384 23754 1444
rect 25728 1384 25788 1444
rect 27764 1384 27824 1444
rect 29804 1384 29864 1444
rect 31838 1384 31898 1444
rect 32856 1482 32916 1542
rect 34756 2614 34816 2674
rect 34598 1482 34658 1542
rect 33874 1384 33934 1444
rect 69011 27560 85796 27774
rect 69106 21978 69166 22038
rect 69218 21978 69278 22038
rect 69328 21978 69388 22038
rect 68442 21266 68502 21326
rect 68782 21266 68842 21326
rect 68892 21266 68952 21326
rect 67060 20320 67120 20380
rect 69978 21978 70038 22038
rect 70088 21978 70148 22038
rect 70196 21978 70256 22038
rect 69542 21266 69602 21326
rect 69654 21266 69714 21326
rect 69762 21266 69822 21326
rect 72936 27364 72996 27424
rect 74018 27364 74078 27424
rect 74976 27364 75036 27424
rect 73462 27118 73522 27178
rect 76012 27364 76072 27424
rect 77018 27364 77078 27424
rect 75498 27118 75558 27178
rect 71280 26186 71340 26246
rect 72444 26186 72504 26246
rect 71150 25982 71210 26042
rect 72444 25982 72504 26042
rect 76516 27230 76576 27290
rect 78040 27364 78100 27424
rect 79058 27364 79118 27424
rect 77536 27120 77596 27180
rect 74480 26082 74540 26142
rect 80082 27364 80142 27424
rect 81094 27364 81154 27424
rect 79566 27120 79626 27180
rect 76516 26082 76576 26142
rect 73460 25048 73520 25108
rect 82112 27364 82172 27424
rect 83124 27364 83184 27424
rect 81608 27122 81668 27182
rect 78554 26186 78614 26246
rect 78550 25982 78610 26042
rect 75496 25048 75556 25108
rect 74478 24952 74538 25012
rect 75182 24946 75246 25010
rect 76354 24946 76418 25010
rect 76516 24842 76576 24902
rect 73460 23910 73520 23970
rect 82620 27230 82680 27290
rect 84152 27364 84212 27424
rect 85164 27364 85224 27424
rect 83640 27122 83700 27182
rect 80588 26186 80648 26246
rect 80586 25982 80646 26042
rect 77530 25048 77590 25108
rect 74476 23796 74540 23860
rect 72438 23658 72502 23722
rect 71280 23512 71340 23572
rect 72262 23512 72322 23572
rect 71866 23176 71926 23236
rect 70998 21978 71058 22038
rect 70414 21266 70474 21326
rect 70524 21266 70584 21326
rect 68998 21160 69058 21220
rect 69434 21160 69494 21220
rect 69872 21160 69932 21220
rect 70306 21160 70366 21220
rect 69218 21044 69278 21104
rect 68782 20320 68842 20380
rect 68998 20216 69058 20276
rect 68892 20118 68952 20178
rect 69216 20320 69276 20380
rect 69106 20118 69166 20178
rect 68442 19482 68502 19542
rect 70088 21044 70148 21104
rect 69434 20216 69494 20276
rect 69326 20118 69386 20178
rect 68782 19382 68842 19442
rect 69652 20320 69712 20380
rect 69872 20216 69932 20276
rect 69544 20118 69604 20178
rect 69654 20118 69714 20178
rect 69760 20118 69820 20178
rect 70088 20320 70148 20380
rect 69978 20118 70038 20178
rect 70882 21044 70942 21104
rect 70306 20216 70366 20276
rect 70196 20118 70256 20178
rect 69652 19382 69712 19442
rect 70526 20320 70586 20380
rect 70412 20118 70472 20178
rect 70526 19382 70586 19442
rect 70882 19382 70942 19442
rect 68998 19284 69058 19344
rect 69434 19284 69494 19344
rect 69872 19284 69932 19344
rect 70306 19284 70366 19344
rect 68442 19166 68502 19226
rect 69108 19166 69168 19226
rect 69216 19166 69276 19226
rect 69324 19166 69384 19226
rect 69970 19166 70030 19226
rect 70088 19166 70148 19226
rect 70197 19166 70255 19224
rect 71752 20872 71812 20932
rect 86182 27364 86242 27424
rect 85676 27122 85736 27182
rect 82622 26082 82682 26142
rect 79568 25046 79628 25106
rect 75496 23910 75556 23970
rect 74476 23362 74540 23426
rect 72262 23076 72322 23136
rect 73428 23076 73488 23136
rect 71994 22030 72054 22090
rect 71866 20768 71926 20828
rect 68782 18446 68842 18506
rect 68892 18446 68952 18506
rect 69546 18446 69606 18506
rect 69652 18446 69712 18506
rect 69762 18446 69822 18506
rect 70414 18446 70474 18506
rect 70526 18446 70586 18506
rect 70998 18446 71058 18506
rect 72130 21932 72190 21992
rect 71994 18358 72054 18418
rect 82764 25978 82824 26038
rect 80588 24948 80648 25008
rect 84656 26082 84716 26142
rect 84658 25978 84718 26038
rect 81604 25046 81664 25106
rect 76990 23906 77050 23966
rect 76514 23176 76574 23236
rect 75464 23076 75524 23136
rect 77530 23968 77590 23970
rect 77498 23910 77590 23968
rect 77990 23910 78050 23970
rect 77498 23908 77558 23910
rect 73432 21822 73492 21882
rect 82622 24842 82682 24902
rect 79034 23912 79094 23972
rect 78548 23658 78612 23722
rect 78548 23374 78612 23438
rect 79536 23968 79596 23972
rect 79536 23912 79628 23968
rect 79568 23908 79628 23912
rect 80050 23912 80110 23972
rect 74446 22128 74506 22188
rect 74446 21932 74506 21992
rect 75466 21934 75526 21994
rect 75466 21822 75526 21882
rect 86696 26186 86756 26246
rect 87834 26186 87894 26246
rect 83640 25046 83700 25106
rect 84658 24842 84718 24902
rect 85674 25044 85734 25104
rect 81078 23912 81138 23972
rect 80584 23658 80648 23722
rect 81604 23966 81664 23968
rect 81572 23908 81664 23966
rect 81572 23906 81632 23908
rect 82100 23902 82160 23962
rect 82588 23906 82648 23966
rect 86696 24948 86756 25008
rect 83100 23902 83160 23962
rect 83640 23906 83700 23966
rect 85674 23906 85734 23966
rect 84656 23796 84720 23860
rect 86692 23658 86756 23722
rect 86664 23382 86724 23442
rect 87834 23376 87894 23436
rect 83610 23076 83670 23136
rect 85644 23076 85704 23136
rect 76482 22128 76542 22188
rect 78522 21820 78582 21880
rect 74448 20768 74508 20828
rect 74448 20564 74508 20624
rect 80556 21820 80616 21880
rect 76484 20768 76544 20828
rect 76482 20666 76542 20726
rect 76482 20564 76542 20624
rect 73430 19616 73490 19676
rect 72262 19408 72322 19468
rect 74444 19306 74504 19366
rect 78518 20872 78578 20932
rect 79538 20872 79598 20932
rect 79538 20566 79598 20626
rect 75466 19616 75526 19676
rect 75466 19508 75526 19568
rect 83612 21820 83672 21880
rect 80556 20566 80616 20626
rect 88088 23076 88148 23136
rect 84626 22128 84686 22188
rect 85646 21820 85706 21880
rect 86662 22128 86722 22188
rect 87928 21934 87988 21994
rect 81574 20872 81634 20932
rect 81572 20566 81632 20626
rect 76478 19306 76538 19366
rect 76682 19312 76742 19372
rect 73426 18358 73486 18418
rect 78520 19618 78580 19678
rect 83608 20768 83668 20828
rect 84476 20886 84536 20946
rect 84624 20776 84684 20836
rect 84476 20566 84536 20626
rect 84628 20568 84688 20628
rect 80556 19618 80616 19678
rect 85644 20666 85704 20726
rect 86664 20776 86724 20836
rect 87796 20776 87856 20836
rect 86662 20568 86722 20628
rect 78516 19312 78576 19372
rect 79536 19308 79596 19368
rect 81570 19308 81630 19368
rect 75462 18358 75522 18418
rect 72130 18228 72190 18288
rect 67060 18088 67120 18148
rect 66904 17982 66964 18042
rect 81784 19304 81844 19364
rect 83610 19620 83670 19680
rect 84120 19304 84180 19364
rect 84632 19306 84692 19366
rect 85646 19620 85706 19680
rect 87928 20568 87988 20628
rect 87796 19508 87856 19568
rect 86666 19306 86726 19366
rect 83614 18358 83674 18418
rect 85650 18358 85710 18418
rect 76484 18088 76544 18148
rect 88088 18088 88148 18148
rect 66134 17864 66194 17924
rect 59912 15362 60012 15364
rect 62512 15362 62612 15364
rect 64316 15362 64416 15364
rect 52918 15262 53018 15362
rect 54712 15262 54812 15362
rect 57312 15262 57412 15362
rect 59912 15264 60012 15362
rect 62512 15264 62612 15362
rect 64316 15264 64416 15362
rect 66904 15132 66964 15192
rect 67060 15132 67120 15192
rect 50944 9048 51004 9108
rect 48364 7491 48424 7551
rect 49954 8406 50014 8466
rect 49306 7640 49366 7700
rect 49048 7491 49108 7551
rect 49824 7640 49884 7700
rect 49564 7491 49624 7551
rect 50627 7622 50687 7628
rect 50627 7574 50633 7622
rect 50633 7574 50681 7622
rect 50681 7574 50687 7622
rect 50627 7568 50687 7574
rect 50945 7590 51005 7650
rect 50082 7491 50142 7551
rect 49952 6943 50012 7003
rect 48364 6116 48424 6176
rect 49954 6442 50014 6502
rect 49306 5676 49366 5736
rect 49048 5527 49108 5587
rect 49824 5676 49884 5736
rect 49564 5527 49624 5587
rect 50627 5658 50687 5664
rect 50627 5610 50633 5658
rect 50633 5610 50681 5658
rect 50681 5610 50687 5658
rect 50627 5604 50687 5610
rect 50945 5626 51005 5686
rect 50082 5527 50142 5587
rect 49952 4979 50012 5039
rect 49954 4442 50014 4502
rect 49306 3676 49366 3736
rect 49048 3527 49108 3587
rect 49824 3676 49884 3736
rect 49564 3527 49624 3587
rect 50627 3658 50687 3664
rect 50627 3610 50633 3658
rect 50633 3610 50681 3658
rect 50681 3610 50687 3658
rect 50627 3604 50687 3610
rect 50945 3626 51005 3686
rect 50082 3527 50142 3587
rect 49952 2979 50012 3039
rect 49954 2352 50014 2412
rect 49306 1586 49366 1646
rect 49048 1437 49108 1497
rect 49824 1586 49884 1646
rect 49564 1437 49624 1497
rect 50627 1568 50687 1574
rect 50627 1520 50633 1568
rect 50633 1520 50681 1568
rect 50681 1520 50687 1568
rect 50627 1514 50687 1520
rect 50945 1536 51005 1596
rect 50082 1437 50142 1497
rect 49952 889 50012 949
rect 3478 -90 34878 64
rect -1266 -576 -666 -276
rect 35166 -576 35766 -276
rect 66134 14146 66194 14206
rect 66800 14032 66860 14092
rect 67286 15124 67346 15184
rect 67062 12692 67122 12752
rect 66926 12480 66986 12540
rect 66800 11578 66860 11638
rect 65640 7592 65700 7652
rect 61974 6320 62034 6380
rect 57564 4880 57624 4940
rect 59604 4880 59664 4940
rect 55412 3976 55472 4036
rect 56550 3976 56610 4036
rect 57564 3880 57624 3940
rect 58586 3764 58646 3824
rect 59604 3880 59664 3940
rect 56696 2864 56756 2924
rect 56548 2756 56608 2816
rect 60624 3976 60684 4036
rect 64136 7356 64196 7416
rect 65048 7356 65108 7416
rect 63266 7246 63326 7306
rect 62352 7138 62412 7198
rect 62482 7030 62542 7090
rect 64030 7138 64090 7198
rect 63812 7030 63872 7090
rect 62940 6530 63000 6590
rect 63048 6430 63108 6490
rect 63050 6320 63110 6380
rect 63596 6530 63656 6590
rect 63486 6430 63546 6490
rect 63484 6320 63544 6380
rect 63158 6210 63218 6270
rect 63378 6210 63438 6270
rect 62482 5706 62542 5766
rect 62352 5584 62412 5644
rect 62940 5706 63000 5766
rect 63158 5584 63218 5644
rect 62832 5460 62892 5520
rect 64928 7246 64988 7306
rect 64248 7138 64308 7198
rect 64466 7030 64526 7090
rect 64466 6530 64526 6590
rect 63812 6320 63872 6380
rect 63922 6320 63982 6380
rect 64358 6320 64418 6380
rect 64032 6210 64092 6270
rect 64248 6210 64308 6270
rect 63596 5706 63656 5766
rect 63376 5584 63436 5644
rect 63270 5334 63330 5394
rect 64928 6756 64988 6816
rect 64576 6410 64636 6470
rect 64140 5706 64200 5766
rect 63812 5586 63872 5646
rect 64468 5586 64528 5646
rect 64928 5706 64988 5766
rect 63702 5460 63762 5520
rect 64574 5460 64634 5520
rect 65170 6530 65230 6590
rect 65170 6284 65230 6344
rect 65048 5334 65108 5394
rect 63604 5228 63656 5280
rect 65902 7622 65962 7682
rect 62280 4900 62340 4960
rect 57566 2644 57626 2704
rect 61748 3764 61808 3824
rect 58582 2864 58642 2924
rect 58584 2756 58644 2816
rect 59604 2644 59664 2704
rect 56550 1660 56610 1720
rect 55412 1554 55472 1614
rect 60452 2864 60512 2924
rect 60620 2756 60680 2816
rect 57568 1762 57628 1822
rect 58584 1554 58644 1614
rect 59598 1762 59658 1822
rect 57054 610 57114 670
rect 62828 5000 62888 5060
rect 64018 5000 64078 5060
rect 65212 5000 65272 5060
rect 65902 5000 65962 5060
rect 63272 4900 63332 4960
rect 63570 4900 63630 4960
rect 62408 3866 62468 3926
rect 62824 3866 62884 3926
rect 64466 4900 64526 4960
rect 64762 4900 64822 4960
rect 63121 3999 63179 4057
rect 62976 3758 63036 3818
rect 63725 3999 63783 4057
rect 63418 3866 63478 3926
rect 63274 3758 63334 3818
rect 63574 3758 63634 3818
rect 62280 2860 62340 2920
rect 60618 1660 60678 1720
rect 61748 1660 61808 1720
rect 58080 610 58140 670
rect 59104 610 59164 670
rect 62974 2860 63034 2920
rect 64016 3866 64076 3926
rect 63868 3758 63928 3818
rect 64316 3999 64374 4057
rect 64164 3758 64224 3818
rect 64913 3999 64971 4057
rect 64610 3866 64670 3926
rect 64464 3758 64524 3818
rect 64766 3758 64826 3818
rect 63420 2752 63480 2812
rect 65208 3866 65268 3926
rect 65056 3758 65116 3818
rect 65509 3999 65567 4057
rect 65360 3758 65420 3818
rect 63870 2860 63930 2920
rect 64164 2860 64224 2920
rect 64614 2752 64674 2812
rect 63122 1768 63182 1828
rect 62524 1674 62584 1734
rect 62972 1566 63032 1626
rect 63416 1674 63476 1734
rect 63270 1566 63330 1626
rect 63716 1768 63776 1828
rect 63566 1566 63626 1626
rect 65058 2860 65118 2920
rect 65360 2860 65420 2920
rect 64316 1768 64376 1828
rect 64014 1674 64074 1734
rect 63870 1566 63930 1626
rect 64166 1566 64226 1626
rect 64612 1674 64672 1734
rect 64464 1566 64524 1626
rect 65902 2752 65962 2812
rect 64910 1768 64970 1828
rect 64760 1566 64820 1626
rect 65504 1768 65564 1828
rect 65212 1674 65272 1734
rect 65056 1566 65116 1626
rect 65360 1566 65420 1626
rect 60004 610 60064 670
rect 62280 640 62340 700
rect 63270 640 63330 700
rect 63568 640 63628 700
rect 64464 640 64524 700
rect 64766 640 64826 700
rect 66026 3758 66086 3818
rect 66926 2936 66986 2996
rect 67518 14032 67578 14092
rect 68536 13934 68596 13994
rect 69554 14032 69614 14092
rect 71588 14032 71648 14092
rect 73628 14032 73688 14092
rect 75664 14032 75724 14092
rect 77698 14032 77758 14092
rect 79734 14032 79794 14092
rect 81770 14032 81830 14092
rect 83806 14032 83866 14092
rect 70574 13934 70634 13994
rect 72608 13934 72668 13994
rect 74642 13934 74702 13994
rect 76682 13934 76742 13994
rect 78716 13934 78776 13994
rect 80754 13934 80814 13994
rect 82786 13934 82846 13994
rect 84824 13934 84884 13994
rect 76682 13722 76742 13782
rect 78714 13722 78774 13782
rect 71222 12802 71282 12862
rect 71592 12802 71652 12862
rect 72094 12802 72154 12862
rect 72606 12802 72666 12862
rect 73134 12802 73194 12862
rect 73626 12802 73686 12862
rect 69046 12692 69106 12752
rect 70068 12692 70128 12752
rect 67522 12480 67582 12540
rect 68020 12480 68080 12540
rect 68532 12480 68592 12540
rect 71088 12588 71148 12648
rect 70574 12480 70634 12540
rect 69036 11578 69096 11638
rect 67286 11364 67346 11424
rect 72088 12588 72148 12648
rect 73108 12588 73168 12648
rect 72608 12480 72668 12540
rect 70052 11590 70112 11650
rect 71072 11590 71132 11650
rect 69548 11486 69608 11546
rect 69554 11252 69614 11312
rect 70572 11486 70632 11546
rect 75658 12802 75718 12862
rect 74140 12692 74200 12752
rect 74644 12692 74704 12752
rect 75160 12692 75220 12752
rect 74642 12480 74702 12540
rect 72084 11590 72144 11650
rect 73110 11590 73170 11650
rect 71584 11486 71644 11546
rect 71590 11252 71650 11312
rect 72604 11486 72664 11546
rect 67398 10322 67458 10382
rect 68536 10322 68596 10382
rect 67286 10122 67346 10182
rect 67180 10020 67240 10080
rect 67286 8886 67346 8946
rect 67180 6530 67240 6590
rect 68534 10122 68594 10182
rect 69552 10242 69612 10302
rect 76180 12692 76240 12752
rect 76682 12692 76742 12752
rect 77182 12692 77242 12752
rect 76798 12480 76858 12540
rect 77694 12802 77754 12862
rect 77322 12588 77382 12648
rect 78208 12692 78268 12752
rect 78330 12588 78390 12648
rect 78718 12692 78778 12752
rect 79226 12692 79286 12752
rect 78522 12478 78582 12538
rect 79730 12802 79790 12862
rect 79372 12588 79432 12648
rect 81768 12802 81828 12862
rect 80234 12692 80294 12752
rect 80756 12692 80816 12752
rect 81246 12692 81306 12752
rect 80756 12480 80816 12540
rect 85844 14032 85904 14092
rect 86862 13934 86922 13994
rect 87874 14032 87934 14092
rect 88598 13934 88658 13994
rect 83292 12802 83352 12862
rect 83806 12802 83866 12862
rect 84314 12802 84374 12862
rect 82278 12692 82338 12752
rect 82790 12692 82850 12752
rect 82264 12588 82324 12648
rect 83302 12588 83362 12648
rect 82788 12480 82848 12540
rect 73626 11486 73686 11546
rect 75662 11486 75722 11546
rect 77700 11486 77760 11546
rect 79730 11486 79790 11546
rect 74646 11364 74706 11424
rect 76680 11364 76740 11424
rect 78710 11364 78770 11424
rect 70570 10346 70630 10406
rect 70066 10128 70126 10188
rect 71592 10242 71652 10302
rect 71070 10128 71130 10188
rect 68534 9090 68594 9150
rect 69040 8988 69100 9048
rect 72606 10346 72666 10406
rect 72082 10128 72142 10188
rect 73624 10242 73684 10302
rect 80750 11486 80810 11546
rect 73102 10128 73162 10188
rect 73624 10130 73684 10190
rect 75658 10242 75718 10302
rect 74642 10020 74702 10080
rect 70572 9090 70632 9150
rect 70570 8886 70630 8946
rect 75660 10130 75720 10190
rect 76676 10020 76736 10080
rect 85334 12692 85394 12752
rect 86354 12692 86414 12752
rect 84302 12588 84362 12648
rect 84820 12480 84880 12540
rect 86862 12480 86922 12540
rect 87366 12480 87426 12540
rect 87876 12480 87936 12540
rect 82266 11590 82326 11650
rect 83302 11590 83362 11650
rect 81768 11486 81828 11546
rect 82788 11486 82848 11546
rect 77698 10242 77758 10302
rect 77696 10130 77756 10190
rect 79732 10242 79792 10302
rect 79928 10238 79988 10298
rect 78716 10020 78776 10080
rect 79732 10130 79792 10190
rect 84318 11590 84378 11650
rect 83804 11486 83864 11546
rect 85840 11486 85900 11546
rect 80750 10346 80810 10406
rect 79928 10020 79988 10080
rect 80222 10022 80282 10082
rect 72608 9090 72668 9150
rect 69554 8786 69614 8846
rect 71078 8880 71138 8940
rect 72100 8880 72160 8940
rect 71588 8786 71648 8846
rect 74640 9090 74700 9150
rect 74132 8988 74192 9048
rect 73114 8880 73174 8940
rect 74132 8880 74192 8940
rect 73624 8786 73684 8846
rect 69036 7862 69096 7922
rect 69946 7862 70006 7922
rect 69036 7646 69096 7706
rect 67400 7542 67460 7602
rect 67286 6284 67346 6344
rect 67192 5228 67244 5280
rect 70948 7862 71008 7922
rect 70074 7646 70134 7706
rect 72100 7862 72160 7922
rect 71588 7760 71648 7820
rect 71088 7646 71148 7706
rect 69034 6634 69094 6694
rect 68536 6530 68596 6590
rect 68532 6320 68592 6380
rect 70042 6634 70102 6694
rect 69552 6418 69612 6478
rect 75152 8880 75212 8940
rect 81766 10130 81826 10190
rect 81250 10022 81310 10082
rect 81768 10016 81828 10076
rect 82786 10346 82846 10406
rect 83804 10130 83864 10190
rect 84820 10238 84880 10298
rect 85324 10234 85384 10294
rect 87984 11252 88044 11312
rect 85844 10130 85904 10190
rect 83804 10016 83864 10076
rect 79222 9102 79282 9162
rect 78716 8974 78776 9034
rect 80752 8776 80812 8836
rect 73110 7862 73170 7922
rect 74116 7862 74176 7922
rect 75160 7862 75220 7922
rect 75660 7868 75720 7928
rect 74114 7646 74174 7706
rect 75154 7646 75214 7706
rect 74638 7542 74698 7602
rect 71056 6634 71116 6694
rect 72094 6634 72154 6694
rect 71590 6418 71650 6478
rect 70570 6320 70630 6380
rect 76168 7646 76228 7706
rect 77696 7868 77756 7928
rect 77176 7646 77236 7706
rect 78220 7646 78280 7706
rect 76680 7542 76740 7602
rect 85842 10016 85902 10076
rect 82264 8880 82324 8940
rect 79732 7868 79792 7928
rect 79210 7646 79270 7706
rect 80228 7646 80288 7706
rect 78718 7542 78778 7602
rect 86860 10346 86920 10406
rect 87878 10364 87938 10424
rect 88478 10234 88538 10294
rect 88228 10130 88288 10190
rect 84316 9102 84376 9162
rect 84454 9106 84514 9166
rect 87984 10016 88044 10076
rect 85336 9106 85396 9166
rect 86342 9106 86402 9166
rect 83294 8880 83354 8940
rect 84454 8880 84514 8940
rect 84822 8880 84882 8940
rect 84822 8776 84882 8836
rect 86860 9102 86920 9162
rect 86860 8974 86920 9034
rect 85838 8778 85898 8838
rect 81770 7868 81830 7928
rect 81762 7760 81822 7820
rect 81262 7646 81322 7706
rect 80752 7542 80812 7602
rect 81264 7538 81324 7598
rect 82286 7538 82346 7598
rect 82786 7544 82846 7604
rect 73112 6634 73172 6694
rect 73628 6640 73688 6700
rect 75664 6640 75724 6700
rect 77696 6640 77756 6700
rect 79730 6640 79790 6700
rect 72610 6320 72670 6380
rect 67398 5298 67458 5358
rect 68538 5082 68598 5142
rect 69552 5396 69612 5456
rect 69556 5202 69616 5262
rect 70570 5298 70630 5358
rect 76680 6530 76740 6590
rect 78716 6530 78776 6590
rect 75662 6418 75722 6478
rect 74646 6320 74706 6380
rect 71588 5396 71648 5456
rect 72094 5298 72154 5358
rect 71592 5202 71652 5262
rect 73626 5396 73686 5456
rect 73116 5298 73176 5358
rect 72606 5082 72666 5142
rect 67286 4166 67346 4226
rect 74138 5298 74198 5358
rect 73620 5202 73680 5262
rect 83806 7868 83866 7928
rect 83802 7760 83862 7820
rect 84294 7646 84354 7706
rect 85844 7868 85904 7928
rect 85840 7760 85900 7820
rect 85332 7646 85392 7706
rect 84820 7544 84880 7604
rect 80752 6642 80812 6702
rect 81106 6642 81166 6702
rect 80748 6530 80808 6590
rect 80258 6432 80318 6492
rect 75488 5416 75548 5476
rect 75658 5416 75718 5476
rect 75142 5298 75202 5358
rect 74640 5082 74700 5142
rect 67180 4040 67240 4100
rect 70570 4040 70630 4100
rect 71090 4052 71150 4112
rect 69552 3930 69612 3990
rect 71588 3930 71648 3990
rect 71206 3836 71266 3896
rect 75488 5202 75548 5262
rect 75664 5208 75724 5268
rect 81296 6432 81356 6492
rect 82272 6432 82332 6492
rect 81106 6324 81166 6384
rect 86358 7646 86418 7706
rect 86862 7544 86922 7604
rect 84824 6642 84884 6702
rect 83288 6432 83348 6492
rect 85314 6432 85374 6492
rect 82786 6320 82846 6380
rect 84822 6320 84882 6380
rect 77700 5416 77760 5476
rect 79732 5416 79792 5476
rect 81772 5416 81832 5476
rect 80750 5318 80810 5378
rect 77692 5208 77752 5268
rect 72608 3930 72668 3990
rect 79736 5208 79796 5268
rect 73624 3930 73684 3990
rect 74644 3930 74704 3990
rect 72090 3836 72150 3896
rect 73112 3836 73172 3896
rect 67518 2936 67578 2996
rect 68032 2936 68092 2996
rect 68530 2936 68590 2996
rect 70572 2936 70632 2996
rect 71080 2824 71140 2884
rect 67060 2718 67120 2778
rect 69046 2718 69106 2778
rect 70068 2718 70128 2778
rect 81764 5208 81824 5268
rect 82790 5082 82850 5142
rect 86344 6432 86404 6492
rect 86858 6320 86918 6380
rect 83802 5208 83862 5268
rect 86856 5318 86916 5378
rect 85842 5208 85902 5268
rect 86360 5212 86420 5272
rect 84820 5082 84880 5142
rect 85346 5084 85406 5144
rect 76674 4166 76734 4226
rect 78716 4166 78776 4226
rect 80752 4166 80812 4226
rect 76170 4052 76230 4112
rect 81258 4056 81318 4116
rect 75662 3930 75722 3990
rect 77692 3930 77752 3990
rect 79730 3930 79790 3990
rect 81766 3930 81826 3990
rect 75154 3836 75214 3896
rect 72604 2936 72664 2996
rect 72092 2824 72152 2884
rect 73106 2824 73166 2884
rect 72606 2718 72666 2778
rect 73118 2718 73178 2778
rect 66654 2614 66714 2674
rect 71082 2614 71142 2674
rect 71586 2614 71646 2674
rect 72102 2614 72162 2674
rect 66026 1566 66086 1626
rect 62824 540 62884 600
rect 64012 540 64072 600
rect 65208 540 65268 600
rect 65902 540 65962 600
rect 67518 1384 67578 1444
rect 68530 1482 68590 1542
rect 74636 2936 74696 2996
rect 74136 2718 74196 2778
rect 74642 2718 74702 2778
rect 75148 2718 75208 2778
rect 73624 2614 73684 2674
rect 69548 1384 69608 1444
rect 76018 2824 76078 2884
rect 75662 2614 75722 2674
rect 76540 2936 76600 2996
rect 76160 2718 76220 2778
rect 76678 2826 76738 2886
rect 77306 2822 77366 2882
rect 77180 2718 77240 2778
rect 78352 2822 78412 2882
rect 78202 2718 78262 2778
rect 77698 2614 77758 2674
rect 78900 2938 78960 2998
rect 78714 2718 78774 2778
rect 79220 2718 79280 2778
rect 86858 5084 86918 5144
rect 82788 3930 82848 3990
rect 83806 4166 83866 4226
rect 83808 3930 83868 3990
rect 82276 3836 82336 3896
rect 83296 3836 83356 3896
rect 80750 2936 80810 2996
rect 80238 2718 80298 2778
rect 80750 2718 80810 2778
rect 81258 2718 81318 2778
rect 79734 2614 79794 2674
rect 84822 3930 84882 3990
rect 85838 4166 85898 4226
rect 88112 9102 88172 9162
rect 88350 8880 88410 8940
rect 88228 8778 88288 8838
rect 88112 7544 88172 7604
rect 88108 6642 88168 6702
rect 88228 5416 88288 5476
rect 88108 5318 88168 5378
rect 88476 7646 88536 7706
rect 88478 5212 88538 5272
rect 88350 5084 88410 5144
rect 87984 4166 88044 4226
rect 86358 4056 86418 4116
rect 85844 3930 85904 3990
rect 84310 3836 84370 3896
rect 85346 3836 85406 3896
rect 82784 2936 82844 2996
rect 82280 2822 82340 2882
rect 83298 2822 83358 2882
rect 84818 2936 84878 2996
rect 84308 2822 84368 2882
rect 81766 2614 81826 2674
rect 82288 2614 82348 2674
rect 82788 2614 82848 2674
rect 83296 2614 83356 2674
rect 83804 2614 83864 2674
rect 84154 2614 84214 2674
rect 86860 2936 86920 2996
rect 87372 2936 87432 2996
rect 87878 2936 87938 2996
rect 85330 2718 85390 2778
rect 86332 2718 86392 2778
rect 76680 1682 76740 1742
rect 78716 1682 78776 1742
rect 70568 1482 70628 1542
rect 72606 1482 72666 1542
rect 74638 1482 74698 1542
rect 76676 1482 76736 1542
rect 78710 1482 78770 1542
rect 80750 1482 80810 1542
rect 82784 1482 82844 1542
rect 84818 1482 84878 1542
rect 71586 1384 71646 1444
rect 73622 1384 73682 1444
rect 75658 1384 75718 1444
rect 77694 1384 77754 1444
rect 79728 1384 79788 1444
rect 81764 1384 81824 1444
rect 83804 1384 83864 1444
rect 85838 1384 85898 1444
rect 86856 1482 86916 1542
rect 88756 2614 88816 2674
rect 88598 1482 88658 1542
rect 87874 1384 87934 1444
rect 57478 -90 88878 64
rect 52734 -576 53334 -276
rect 89166 -576 89766 -276
<< metal2 >>
rect 11434 28156 12034 28166
rect 11434 27846 12034 27856
rect 35066 28156 35666 28166
rect 35066 27846 35666 27856
rect 65434 28156 66034 28166
rect 65434 27846 66034 27856
rect 89066 28156 89666 28166
rect 89066 27846 89666 27856
rect 14948 27774 31828 27806
rect -1414 27642 -1354 27651
rect -1420 27582 -1414 27642
rect -1354 27582 -1348 27642
rect -1414 27573 -1354 27582
rect 14948 27560 15011 27774
rect 31796 27560 31828 27774
rect 68948 27774 85828 27806
rect 14948 27540 31828 27560
rect 47796 27680 48490 27702
rect 47796 27564 47824 27680
rect 48462 27564 48490 27680
rect 14948 27538 19302 27540
rect 47796 27536 48490 27564
rect 68948 27560 69011 27774
rect 85796 27560 85828 27774
rect 68948 27540 85828 27560
rect 68948 27538 73302 27540
rect 18936 27424 18996 27430
rect 20018 27424 20078 27430
rect 20976 27424 21036 27430
rect 22012 27424 22072 27430
rect 23018 27424 23078 27430
rect 24040 27424 24100 27430
rect 25058 27424 25118 27430
rect 26082 27424 26142 27430
rect 27094 27424 27154 27430
rect 28112 27424 28172 27430
rect 29124 27424 29184 27430
rect 30152 27424 30212 27430
rect 31164 27424 31224 27430
rect 32182 27424 32242 27430
rect 18996 27364 20018 27424
rect 20078 27364 20976 27424
rect 21036 27364 22012 27424
rect 22072 27364 23018 27424
rect 23078 27364 24040 27424
rect 24100 27364 25058 27424
rect 25118 27364 26082 27424
rect 26142 27364 27094 27424
rect 27154 27364 28112 27424
rect 28172 27364 29124 27424
rect 29184 27364 30152 27424
rect 30212 27364 31164 27424
rect 31224 27364 32182 27424
rect 18936 27358 18996 27364
rect 20018 27358 20078 27364
rect 20976 27358 21036 27364
rect 22012 27358 22072 27364
rect 23018 27358 23078 27364
rect 24040 27358 24100 27364
rect 25058 27358 25118 27364
rect 26082 27358 26142 27364
rect 27094 27358 27154 27364
rect 28112 27358 28172 27364
rect 29124 27358 29184 27364
rect 30152 27358 30212 27364
rect 31164 27358 31224 27364
rect 32182 27358 32242 27364
rect 72936 27424 72996 27430
rect 74018 27424 74078 27430
rect 74976 27424 75036 27430
rect 76012 27424 76072 27430
rect 77018 27424 77078 27430
rect 78040 27424 78100 27430
rect 79058 27424 79118 27430
rect 80082 27424 80142 27430
rect 81094 27424 81154 27430
rect 82112 27424 82172 27430
rect 83124 27424 83184 27430
rect 84152 27424 84212 27430
rect 85164 27424 85224 27430
rect 86182 27424 86242 27430
rect 72996 27364 74018 27424
rect 74078 27364 74976 27424
rect 75036 27364 76012 27424
rect 76072 27364 77018 27424
rect 77078 27364 78040 27424
rect 78100 27364 79058 27424
rect 79118 27364 80082 27424
rect 80142 27364 81094 27424
rect 81154 27364 82112 27424
rect 82172 27364 83124 27424
rect 83184 27364 84152 27424
rect 84212 27364 85164 27424
rect 85224 27364 86182 27424
rect 72936 27358 72996 27364
rect 74018 27358 74078 27364
rect 74976 27358 75036 27364
rect 76012 27358 76072 27364
rect 77018 27358 77078 27364
rect 78040 27358 78100 27364
rect 79058 27358 79118 27364
rect 80082 27358 80142 27364
rect 81094 27358 81154 27364
rect 82112 27358 82172 27364
rect 83124 27358 83184 27364
rect 84152 27358 84212 27364
rect 85164 27358 85224 27364
rect 86182 27358 86242 27364
rect 22516 27290 22576 27296
rect 28620 27290 28680 27296
rect 22576 27230 28620 27290
rect 22516 27224 22576 27230
rect 28620 27224 28680 27230
rect 76516 27290 76576 27296
rect 82620 27290 82680 27296
rect 76576 27230 82620 27290
rect 76516 27224 76576 27230
rect 82620 27224 82680 27230
rect 19462 27178 19522 27184
rect 21498 27178 21558 27184
rect 23536 27180 23596 27186
rect 25566 27180 25626 27186
rect 27608 27182 27668 27188
rect 29640 27182 29700 27188
rect 31676 27182 31736 27188
rect 19522 27118 21498 27178
rect 21558 27120 23536 27178
rect 23596 27120 25566 27180
rect 25626 27122 27608 27180
rect 27668 27122 29640 27182
rect 29700 27122 31676 27182
rect 25626 27120 27806 27122
rect 21558 27118 23718 27120
rect 19462 27112 19522 27118
rect 21498 27112 21558 27118
rect 23536 27114 23596 27118
rect 25566 27114 25626 27120
rect 27608 27116 27668 27120
rect 29640 27116 29700 27122
rect 31676 27116 31736 27122
rect 73462 27178 73522 27184
rect 75498 27178 75558 27184
rect 77536 27180 77596 27186
rect 79566 27180 79626 27186
rect 81608 27182 81668 27188
rect 83640 27182 83700 27188
rect 85676 27182 85736 27188
rect 73522 27118 75498 27178
rect 75558 27120 77536 27178
rect 77596 27120 79566 27180
rect 79626 27122 81608 27180
rect 81668 27122 83640 27182
rect 83700 27122 85676 27182
rect 79626 27120 81806 27122
rect 75558 27118 77718 27120
rect 73462 27112 73522 27118
rect 75498 27112 75558 27118
rect 77536 27114 77596 27118
rect 79566 27114 79626 27120
rect 81608 27116 81668 27120
rect 83640 27116 83700 27122
rect 85676 27116 85736 27122
rect 17280 26246 17340 26252
rect 18444 26246 18504 26252
rect 24554 26246 24614 26252
rect 17340 26186 18444 26246
rect 18504 26186 24554 26246
rect 17280 26180 17340 26186
rect 18444 26180 18504 26186
rect 24554 26180 24614 26186
rect 26588 26246 26648 26252
rect 32696 26246 32756 26252
rect 33834 26246 33894 26252
rect 26648 26186 32696 26246
rect 32756 26186 33834 26246
rect 26588 26180 26648 26186
rect 32696 26180 32756 26186
rect 33834 26180 33894 26186
rect 71280 26246 71340 26252
rect 72444 26246 72504 26252
rect 78554 26246 78614 26252
rect 71340 26186 72444 26246
rect 72504 26186 78554 26246
rect 71280 26180 71340 26186
rect 72444 26180 72504 26186
rect 78554 26180 78614 26186
rect 80588 26246 80648 26252
rect 86696 26246 86756 26252
rect 87834 26246 87894 26252
rect 80648 26186 86696 26246
rect 86756 26186 87834 26246
rect 80588 26180 80648 26186
rect 86696 26180 86756 26186
rect 87834 26180 87894 26186
rect 20480 26142 20540 26148
rect 22516 26142 22576 26148
rect 28622 26142 28682 26148
rect 30656 26142 30716 26148
rect 20540 26082 22516 26142
rect 22576 26134 22994 26142
rect 23210 26134 28622 26142
rect 22576 26088 28622 26134
rect 22576 26084 25010 26088
rect 22576 26082 23984 26084
rect 24222 26082 25010 26084
rect 25226 26082 28622 26088
rect 28682 26082 30656 26142
rect 20480 26076 20540 26082
rect 22516 26076 22576 26082
rect 28622 26076 28682 26082
rect 30656 26076 30716 26082
rect 74480 26142 74540 26148
rect 76516 26142 76576 26148
rect 82622 26142 82682 26148
rect 84656 26142 84716 26148
rect 74540 26082 76516 26142
rect 76576 26134 76994 26142
rect 77210 26134 82622 26142
rect 76576 26088 82622 26134
rect 76576 26084 79010 26088
rect 76576 26082 77984 26084
rect 78222 26082 79010 26084
rect 79226 26082 82622 26088
rect 82682 26082 84656 26142
rect 74480 26076 74540 26082
rect 76516 26076 76576 26082
rect 82622 26076 82682 26082
rect 84656 26076 84716 26082
rect 17150 26042 17210 26048
rect 18444 26042 18504 26048
rect 24550 26042 24610 26048
rect 26586 26042 26646 26048
rect 17210 25982 18444 26042
rect 18504 25982 24550 26042
rect 24610 25982 26586 26042
rect 17150 25976 17210 25982
rect 18444 25976 18504 25982
rect 24550 25976 24610 25982
rect 26586 25976 26646 25982
rect 28764 26038 28824 26044
rect 30658 26038 30718 26044
rect 28824 25978 30658 26038
rect 28764 25972 28824 25978
rect 30658 25972 30718 25978
rect 71150 26042 71210 26048
rect 72444 26042 72504 26048
rect 78550 26042 78610 26048
rect 80586 26042 80646 26048
rect 71210 25982 72444 26042
rect 72504 25982 78550 26042
rect 78610 25982 80586 26042
rect 71150 25976 71210 25982
rect 72444 25976 72504 25982
rect 78550 25976 78610 25982
rect 80586 25976 80646 25982
rect 82764 26038 82824 26044
rect 84658 26038 84718 26044
rect 82824 25978 84658 26038
rect 82764 25972 82824 25978
rect 84658 25972 84718 25978
rect 48522 25370 48528 25430
rect 48588 25370 49187 25430
rect 19460 25108 19520 25114
rect 21496 25108 21556 25114
rect 23530 25108 23590 25114
rect 25568 25108 25628 25112
rect 19520 25048 21496 25108
rect 21556 25048 23530 25108
rect 23590 25106 25772 25108
rect 27604 25106 27664 25112
rect 29640 25106 29700 25112
rect 23590 25048 25568 25106
rect 19460 25042 19520 25048
rect 21496 25042 21556 25048
rect 23530 25042 23590 25048
rect 25628 25046 27604 25106
rect 27664 25046 29640 25106
rect 29700 25104 30510 25106
rect 31674 25104 31734 25110
rect 29700 25046 31674 25104
rect 25568 25040 25628 25046
rect 27604 25040 27664 25046
rect 29539 25044 30054 25046
rect 30304 25044 31674 25046
rect 29640 25040 29700 25044
rect 31674 25038 31734 25044
rect 20478 25012 20538 25018
rect 20538 24952 21050 25012
rect 20478 24946 20538 24952
rect 20990 24902 21050 24952
rect 21182 25010 21246 25016
rect 22354 25010 22418 25016
rect 21246 24946 22354 25010
rect 21182 24940 21246 24946
rect 22354 24940 22418 24946
rect 26588 25008 26648 25014
rect 32696 25008 32756 25014
rect 26648 24948 32696 25008
rect 26588 24942 26648 24948
rect 32696 24942 32756 24948
rect 22516 24902 22576 24908
rect 28622 24902 28682 24908
rect 30658 24902 30718 24908
rect 20990 24842 22516 24902
rect 22576 24842 28622 24902
rect 28682 24842 30658 24902
rect 22516 24836 22576 24842
rect 28622 24836 28682 24842
rect 30658 24836 30718 24842
rect 47880 24664 47940 24670
rect 48398 24664 48458 24670
rect 47940 24604 48398 24664
rect 48458 24604 48467 24664
rect 47880 24598 47940 24604
rect 48398 24598 48458 24604
rect 49127 24592 49187 25370
rect 73460 25108 73520 25114
rect 75496 25108 75556 25114
rect 77530 25108 77590 25114
rect 79568 25108 79628 25112
rect 73520 25048 75496 25108
rect 75556 25048 77530 25108
rect 77590 25106 79772 25108
rect 81604 25106 81664 25112
rect 83640 25106 83700 25112
rect 77590 25048 79568 25106
rect 73460 25042 73520 25048
rect 75496 25042 75556 25048
rect 77530 25042 77590 25048
rect 79628 25046 81604 25106
rect 81664 25046 83640 25106
rect 83700 25104 84510 25106
rect 85674 25104 85734 25110
rect 83700 25046 85674 25104
rect 79568 25040 79628 25046
rect 81604 25040 81664 25046
rect 83539 25044 84054 25046
rect 84304 25044 85674 25046
rect 83640 25040 83700 25044
rect 85674 25038 85734 25044
rect 74478 25012 74538 25018
rect 74538 24952 75050 25012
rect 74478 24946 74538 24952
rect 74990 24902 75050 24952
rect 75182 25010 75246 25016
rect 76354 25010 76418 25016
rect 75246 24946 76354 25010
rect 75182 24940 75246 24946
rect 76354 24940 76418 24946
rect 80588 25008 80648 25014
rect 86696 25008 86756 25014
rect 80648 24948 86696 25008
rect 80588 24942 80648 24948
rect 86696 24942 86756 24948
rect 76516 24902 76576 24908
rect 82622 24902 82682 24908
rect 84658 24902 84718 24908
rect 74990 24842 76516 24902
rect 76576 24842 82622 24902
rect 82682 24842 84658 24902
rect 76516 24836 76576 24842
rect 82622 24836 82682 24842
rect 84658 24836 84718 24842
rect 49127 24532 49201 24592
rect 49261 24532 49267 24592
rect 49513 24554 49519 24614
rect 49579 24554 49585 24614
rect 47622 24515 47682 24521
rect 48138 24515 48198 24521
rect 47611 24455 47622 24515
rect 47684 24455 48138 24515
rect 48198 24455 48656 24515
rect 48716 24455 48722 24515
rect 47622 24449 47682 24455
rect 48138 24449 48198 24455
rect 19460 23970 19520 23976
rect 21496 23970 21556 23976
rect 23530 23970 23590 23976
rect 23990 23970 24050 23976
rect 25568 23972 25628 23974
rect 25028 23970 25034 23972
rect 19520 23910 21496 23970
rect 21556 23968 23530 23970
rect 21556 23966 23498 23968
rect 21556 23910 22990 23966
rect 19460 23904 19520 23910
rect 21496 23904 21556 23910
rect 22984 23906 22990 23910
rect 23050 23910 23498 23966
rect 23590 23910 23990 23970
rect 24050 23912 25034 23970
rect 25094 23970 25100 23972
rect 25530 23970 25536 23972
rect 25094 23912 25536 23970
rect 25596 23970 25628 23972
rect 26044 23970 26050 23972
rect 25596 23968 26050 23970
rect 25628 23912 26050 23968
rect 26110 23970 26116 23972
rect 27072 23970 27078 23972
rect 26110 23912 27078 23970
rect 27138 23970 27144 23972
rect 27138 23968 27450 23970
rect 27604 23968 27664 23974
rect 29640 23968 29700 23972
rect 27138 23966 27604 23968
rect 27664 23966 29828 23968
rect 31674 23966 31734 23972
rect 27138 23912 27572 23966
rect 24050 23910 25568 23912
rect 23050 23906 23056 23910
rect 23492 23908 23498 23910
rect 23558 23908 23590 23910
rect 23530 23904 23590 23908
rect 23990 23904 24050 23910
rect 25628 23910 27572 23912
rect 25628 23908 26016 23910
rect 26222 23908 27036 23910
rect 27242 23908 27572 23910
rect 27664 23962 28588 23966
rect 27664 23908 28100 23962
rect 25568 23902 25628 23908
rect 27566 23906 27572 23908
rect 27632 23906 27664 23908
rect 27604 23902 27664 23906
rect 28094 23902 28100 23908
rect 28160 23908 28588 23962
rect 28160 23902 28166 23908
rect 28582 23906 28588 23908
rect 28648 23962 29640 23966
rect 28648 23908 29100 23962
rect 28648 23906 28654 23908
rect 29094 23902 29100 23908
rect 29160 23908 29640 23962
rect 29160 23902 29166 23908
rect 29700 23906 31674 23966
rect 48526 23967 48586 23973
rect 49519 23968 49579 24554
rect 49033 23967 49579 23968
rect 47250 23934 47310 23940
rect 29640 23900 29700 23906
rect 31674 23900 31734 23906
rect 42781 23874 42790 23934
rect 42850 23874 47250 23934
rect 48586 23908 49579 23967
rect 48586 23907 49137 23908
rect 48526 23901 48586 23907
rect 47250 23868 47310 23874
rect 20476 23860 20540 23866
rect 30656 23860 30720 23866
rect 38874 23861 38964 23866
rect 20540 23796 30656 23860
rect 30720 23796 34304 23860
rect 20476 23790 20540 23796
rect 30656 23790 30720 23796
rect 18438 23722 18502 23728
rect 24548 23722 24612 23728
rect 18502 23658 24548 23722
rect 18438 23652 18502 23658
rect 24548 23652 24612 23658
rect 26584 23722 26648 23728
rect 32692 23722 32756 23728
rect 26648 23714 29024 23722
rect 29406 23714 32692 23722
rect 26648 23658 32692 23714
rect 26584 23652 26648 23658
rect 17280 23572 17340 23578
rect 26788 23572 26848 23658
rect 32692 23652 32756 23658
rect 17340 23512 18262 23572
rect 18322 23512 26848 23572
rect 17280 23506 17340 23512
rect 32658 23440 32664 23442
rect 24548 23438 32664 23440
rect 20476 23426 20540 23432
rect 11640 23362 20476 23426
rect 24542 23374 24548 23438
rect 24612 23382 32664 23438
rect 32724 23440 32730 23442
rect 32724 23436 33894 23440
rect 32724 23382 33834 23436
rect 24612 23376 33834 23382
rect 33894 23376 33900 23436
rect 24612 23374 24618 23376
rect 11206 18913 11306 18918
rect 11202 18823 11211 18913
rect 11301 18823 11310 18913
rect -1414 16408 -1354 16414
rect -8748 16348 -8742 16408
rect -8682 16348 -1414 16408
rect -1414 16342 -1354 16348
rect 10953 16318 10962 16418
rect 11062 16318 11071 16418
rect -11836 16240 -11830 16300
rect -11770 16240 -11171 16300
rect -9236 16240 -9230 16300
rect -9170 16240 -8571 16300
rect -12478 15534 -12418 15540
rect -11960 15534 -11900 15540
rect -12418 15474 -11960 15534
rect -12478 15468 -12418 15474
rect -11960 15468 -11900 15474
rect -11231 15462 -11171 16240
rect -9878 15534 -9818 15540
rect -9360 15534 -9300 15540
rect -11231 15402 -11157 15462
rect -11097 15402 -11091 15462
rect -10845 15424 -10839 15484
rect -10779 15424 -10773 15484
rect -9818 15474 -9360 15534
rect -9878 15468 -9818 15474
rect -9360 15468 -9300 15474
rect -8631 15462 -8571 16240
rect -12736 15385 -12676 15391
rect -12220 15385 -12160 15391
rect -13295 15325 -13286 15385
rect -13226 15325 -12736 15385
rect -12676 15325 -12220 15385
rect -12160 15325 -11702 15385
rect -11642 15325 -11636 15385
rect -12736 15319 -12676 15325
rect -12220 15319 -12160 15325
rect -12478 14956 -12418 14962
rect -13467 14610 -13377 14614
rect -12478 14610 -12418 14896
rect -11832 14837 -11772 14843
rect -10839 14838 -10779 15424
rect -8631 15402 -8557 15462
rect -8497 15402 -8491 15462
rect -8245 15424 -8239 15484
rect -8179 15424 -8173 15484
rect -10136 15385 -10076 15391
rect -9620 15385 -9560 15391
rect -10629 15325 -10620 15385
rect -10560 15325 -10136 15385
rect -10076 15325 -9620 15385
rect -9560 15325 -9102 15385
rect -9042 15325 -9036 15385
rect -10136 15319 -10076 15325
rect -9620 15319 -9560 15325
rect -11325 14837 -10779 14838
rect -9878 14952 -9818 14958
rect -11772 14778 -10006 14837
rect -11772 14777 -11221 14778
rect -10838 14777 -10006 14778
rect -9946 14777 -9940 14837
rect -11832 14771 -11772 14777
rect -13472 14605 -12418 14610
rect -13472 14515 -13467 14605
rect -13377 14515 -12418 14605
rect -13472 14510 -12418 14515
rect -13467 14506 -13377 14510
rect -9878 13120 -9818 14892
rect -9232 14837 -9172 14843
rect -8239 14838 -8179 15424
rect -1082 15362 -982 15368
rect 712 15362 812 15368
rect 3312 15362 3412 15368
rect 5912 15364 6012 15370
rect 8512 15364 8612 15370
rect 10316 15364 10416 15370
rect -1086 15267 -1082 15357
rect -982 15267 -978 15357
rect 708 15267 712 15357
rect 812 15267 816 15357
rect 3308 15267 3312 15357
rect 3412 15267 3416 15357
rect 5908 15269 5912 15359
rect 6012 15269 6016 15359
rect 8508 15269 8512 15359
rect 8612 15269 8616 15359
rect 10312 15269 10316 15359
rect 10416 15269 10420 15359
rect -1082 15256 -982 15262
rect 712 15256 812 15262
rect 3312 15256 3412 15262
rect 5912 15258 6012 15264
rect 8512 15258 8612 15264
rect 10316 15258 10416 15264
rect -1933 15092 -1924 15152
rect -1864 15092 -1855 15152
rect -1924 14838 -1864 15092
rect 10962 14983 11062 16318
rect 11206 15882 11306 18823
rect 11197 15782 11206 15882
rect 11306 15782 11315 15882
rect 10958 14893 10967 14983
rect 11057 14893 11066 14983
rect 10962 14888 11062 14893
rect -8725 14837 -1864 14838
rect -9172 14778 -1864 14837
rect 11206 14812 11306 15782
rect -9172 14777 -8621 14778
rect -9232 14771 -9172 14777
rect 11197 14712 11206 14812
rect 11306 14712 11315 14812
rect -8756 14652 -8750 14712
rect -8690 14652 -1792 14712
rect -1732 14652 -1726 14712
rect -9878 13051 -9818 13060
rect -9960 11043 -9846 11048
rect -9964 10939 -9955 11043
rect -9851 10939 -9842 11043
rect -5826 11027 -5720 11032
rect -9960 10871 -9846 10939
rect -5830 10931 -5821 11027
rect -5725 10931 -5716 11027
rect -5826 10891 -5720 10931
rect -9960 10757 -8667 10871
rect -5826 10785 -4683 10891
rect -8781 10725 -8667 10757
rect -8781 10602 -8667 10611
rect -4789 10715 -4683 10785
rect -4789 10600 -4683 10609
rect 11640 7652 11700 23362
rect 20476 23356 20540 23362
rect 22514 23236 22574 23242
rect 11902 23176 17866 23236
rect 17926 23176 22514 23236
rect 11902 7682 11962 23176
rect 22514 23170 22574 23176
rect 18262 23136 18322 23142
rect 19428 23136 19488 23142
rect 21464 23136 21524 23142
rect 18322 23076 19428 23136
rect 19488 23076 21464 23136
rect 18262 23070 18322 23076
rect 19428 23070 19488 23076
rect 21464 23070 21524 23076
rect 29610 23136 29670 23142
rect 31644 23136 31704 23142
rect 34088 23136 34148 23142
rect 29670 23076 31644 23136
rect 31704 23076 34088 23136
rect 29610 23070 29670 23076
rect 31644 23070 31704 23076
rect 34088 23070 34148 23076
rect 20446 22188 20506 22194
rect 22482 22188 22542 22194
rect 20506 22128 22482 22188
rect 20446 22122 20506 22128
rect 22482 22122 22542 22128
rect 30626 22188 30686 22194
rect 32662 22188 32722 22194
rect 30686 22128 32662 22188
rect 30626 22122 30686 22128
rect 17994 22090 18054 22096
rect 30734 22090 30794 22128
rect 32662 22122 32722 22128
rect 15106 22038 15166 22044
rect 15218 22038 15278 22044
rect 15328 22038 15388 22044
rect 15978 22038 16038 22044
rect 16088 22038 16148 22044
rect 16196 22038 16256 22044
rect 16998 22038 17058 22044
rect 12280 21978 15106 22038
rect 15166 21978 15218 22038
rect 15278 21978 15328 22038
rect 15388 21978 15978 22038
rect 16038 21978 16088 22038
rect 16148 21978 16196 22038
rect 16256 21978 16998 22038
rect 18054 22030 30794 22090
rect 17994 22024 18054 22030
rect 12128 17864 12134 17924
rect 12194 17864 12200 17924
rect 12134 14206 12194 17864
rect 12128 14146 12134 14206
rect 12194 14146 12200 14206
rect 11634 7592 11640 7652
rect 11700 7592 11706 7652
rect 11896 7622 11902 7682
rect 11962 7622 11968 7682
rect 10136 7416 10196 7422
rect 11048 7416 11108 7422
rect 12280 7416 12340 21978
rect 15106 21972 15166 21978
rect 15218 21972 15278 21978
rect 15328 21972 15388 21978
rect 15978 21972 16038 21978
rect 16088 21972 16148 21978
rect 16196 21972 16256 21978
rect 16998 21972 17058 21978
rect 18130 21992 18190 21998
rect 20446 21992 20506 21998
rect 18190 21932 20446 21992
rect 18130 21926 18190 21932
rect 20446 21926 20506 21932
rect 21466 21994 21526 22000
rect 33928 21994 33988 22000
rect 21526 21934 33928 21994
rect 21466 21928 21526 21934
rect 33928 21928 33988 21934
rect 19432 21882 19492 21888
rect 21466 21882 21526 21888
rect 19492 21822 21466 21882
rect 19432 21816 19492 21822
rect 21466 21816 21526 21822
rect 24522 21880 24582 21886
rect 26556 21880 26616 21886
rect 24582 21820 26556 21880
rect 24522 21814 24582 21820
rect 26556 21814 26616 21820
rect 29612 21880 29672 21886
rect 31646 21882 31706 21886
rect 34240 21882 34304 23796
rect 38870 23781 38879 23861
rect 38959 23781 38968 23861
rect 38874 23705 38964 23781
rect 38874 23615 41091 23705
rect 41001 23527 41091 23615
rect 41001 23428 41091 23437
rect 48522 23370 48528 23430
rect 48588 23370 49187 23430
rect 47880 22664 47940 22670
rect 48398 22664 48458 22670
rect 47867 22604 47876 22664
rect 47940 22604 48398 22664
rect 47880 22598 47940 22604
rect 48398 22598 48458 22604
rect 49127 22592 49187 23370
rect 49519 22614 49579 23908
rect 73460 23970 73520 23976
rect 75496 23970 75556 23976
rect 77530 23970 77590 23976
rect 77990 23970 78050 23976
rect 79568 23972 79628 23974
rect 79028 23970 79034 23972
rect 73520 23910 75496 23970
rect 75556 23968 77530 23970
rect 75556 23966 77498 23968
rect 75556 23910 76990 23966
rect 73460 23904 73520 23910
rect 75496 23904 75556 23910
rect 76984 23906 76990 23910
rect 77050 23910 77498 23966
rect 77590 23910 77990 23970
rect 78050 23912 79034 23970
rect 79094 23970 79100 23972
rect 79530 23970 79536 23972
rect 79094 23912 79536 23970
rect 79596 23970 79628 23972
rect 80044 23970 80050 23972
rect 79596 23968 80050 23970
rect 79628 23912 80050 23968
rect 80110 23970 80116 23972
rect 81072 23970 81078 23972
rect 80110 23912 81078 23970
rect 81138 23970 81144 23972
rect 81138 23968 81450 23970
rect 81604 23968 81664 23974
rect 83640 23968 83700 23972
rect 81138 23966 81604 23968
rect 81664 23966 83828 23968
rect 85674 23966 85734 23972
rect 81138 23912 81572 23966
rect 78050 23910 79568 23912
rect 77050 23906 77056 23910
rect 77492 23908 77498 23910
rect 77558 23908 77590 23910
rect 77530 23904 77590 23908
rect 77990 23904 78050 23910
rect 79628 23910 81572 23912
rect 79628 23908 80016 23910
rect 80222 23908 81036 23910
rect 81242 23908 81572 23910
rect 81664 23962 82588 23966
rect 81664 23908 82100 23962
rect 79568 23902 79628 23908
rect 81566 23906 81572 23908
rect 81632 23906 81664 23908
rect 81604 23902 81664 23906
rect 82094 23902 82100 23908
rect 82160 23908 82588 23962
rect 82160 23902 82166 23908
rect 82582 23906 82588 23908
rect 82648 23962 83640 23966
rect 82648 23908 83100 23962
rect 82648 23906 82654 23908
rect 83094 23902 83100 23908
rect 83160 23908 83640 23962
rect 83160 23902 83166 23908
rect 83700 23906 85674 23966
rect 83640 23900 83700 23906
rect 85674 23900 85734 23906
rect 74476 23860 74540 23866
rect 84656 23860 84720 23866
rect 74540 23796 84656 23860
rect 84720 23796 88304 23860
rect 74476 23790 74540 23796
rect 84656 23790 84720 23796
rect 72438 23722 72502 23728
rect 78548 23722 78612 23728
rect 72502 23658 78548 23722
rect 72438 23652 72502 23658
rect 78548 23652 78612 23658
rect 80584 23722 80648 23728
rect 86692 23722 86756 23728
rect 80648 23714 83024 23722
rect 83406 23714 86692 23722
rect 80648 23658 86692 23714
rect 80584 23652 80648 23658
rect 71280 23572 71340 23578
rect 80788 23572 80848 23658
rect 86692 23652 86756 23658
rect 71340 23512 72262 23572
rect 72322 23512 80848 23572
rect 71280 23506 71340 23512
rect 86658 23440 86664 23442
rect 78548 23438 86664 23440
rect 74476 23426 74540 23432
rect 65640 23362 74476 23426
rect 78542 23374 78548 23438
rect 78612 23382 86664 23438
rect 86724 23440 86730 23442
rect 86724 23436 87894 23440
rect 86724 23382 87834 23436
rect 78612 23376 87834 23382
rect 87894 23376 87900 23436
rect 78612 23374 78618 23376
rect 49127 22532 49201 22592
rect 49261 22532 49267 22592
rect 49513 22554 49519 22614
rect 49579 22554 49585 22614
rect 47622 22515 47682 22521
rect 48138 22515 48198 22521
rect 47611 22455 47622 22515
rect 47682 22455 48138 22515
rect 48198 22455 48656 22515
rect 48716 22455 48725 22515
rect 47622 22449 47682 22455
rect 48138 22449 48198 22455
rect 48526 21967 48586 21973
rect 49519 21968 49579 22554
rect 49033 21967 49579 21968
rect 46978 21920 47038 21926
rect 31578 21880 34304 21882
rect 29672 21820 31646 21880
rect 31706 21820 34304 21880
rect 42791 21860 42800 21920
rect 42860 21860 46978 21920
rect 48586 21908 49579 21967
rect 48586 21907 49137 21908
rect 48526 21901 48586 21907
rect 46978 21854 47038 21860
rect 29612 21814 29672 21820
rect 31578 21818 34304 21820
rect 31646 21814 31706 21818
rect 40228 21414 40328 21423
rect 14442 21326 14502 21332
rect 14782 21326 14842 21332
rect 14892 21326 14952 21332
rect 15542 21326 15602 21332
rect 15654 21326 15714 21332
rect 15762 21326 15822 21332
rect 16414 21326 16474 21332
rect 16524 21326 16584 21332
rect 14502 21266 14782 21326
rect 14842 21266 14892 21326
rect 14952 21266 15542 21326
rect 15602 21266 15654 21326
rect 15714 21266 15762 21326
rect 15822 21266 16414 21326
rect 16474 21266 16524 21326
rect 14442 21260 14502 21266
rect 14782 21260 14842 21266
rect 14892 21260 14952 21266
rect 15542 21260 15602 21266
rect 15654 21260 15714 21266
rect 15762 21260 15822 21266
rect 16414 21260 16474 21266
rect 16524 21260 16584 21266
rect 36254 21314 40228 21414
rect 14998 21220 15058 21226
rect 15434 21220 15494 21226
rect 15872 21220 15932 21226
rect 16306 21220 16366 21226
rect 15058 21160 15434 21220
rect 15494 21160 15872 21220
rect 15932 21160 16306 21220
rect 14998 21154 15058 21160
rect 15434 21154 15494 21160
rect 15872 21154 15932 21160
rect 16306 21154 16366 21160
rect 15218 21104 15278 21110
rect 16088 21104 16148 21110
rect 16882 21104 16942 21110
rect 15278 21044 16088 21104
rect 16148 21044 16882 21104
rect 15218 21038 15278 21044
rect 16088 21038 16148 21044
rect 16882 21038 16942 21044
rect 30476 20946 30536 20952
rect 17752 20932 17812 20938
rect 24518 20932 24578 20938
rect 25538 20932 25598 20938
rect 27574 20932 27634 20938
rect 17812 20872 24518 20932
rect 24578 20872 25538 20932
rect 25598 20872 27574 20932
rect 30536 20886 34898 20946
rect 30476 20880 30536 20886
rect 17752 20866 17812 20872
rect 24518 20866 24578 20872
rect 25538 20866 25598 20872
rect 27574 20866 27634 20872
rect 30624 20836 30684 20842
rect 32664 20836 32724 20842
rect 33796 20836 33856 20842
rect 17866 20828 17926 20834
rect 22484 20828 22544 20834
rect 29608 20828 29668 20834
rect 17926 20768 20448 20828
rect 20508 20768 22484 20828
rect 22544 20768 29608 20828
rect 30684 20776 32664 20836
rect 32724 20776 33796 20836
rect 30624 20770 30684 20776
rect 32664 20770 32724 20776
rect 33796 20770 33856 20776
rect 17866 20762 17926 20768
rect 22484 20762 22544 20768
rect 29608 20762 29668 20768
rect 22482 20726 22542 20732
rect 31644 20726 31704 20732
rect 22542 20666 31644 20726
rect 22482 20660 22542 20666
rect 31644 20660 31704 20666
rect 20448 20624 20508 20630
rect 22482 20624 22542 20630
rect 20508 20564 22482 20624
rect 20448 20558 20508 20564
rect 22482 20558 22542 20564
rect 25538 20626 25598 20632
rect 26556 20626 26616 20632
rect 27572 20626 27632 20632
rect 30476 20626 30536 20632
rect 25598 20566 26556 20626
rect 26616 20566 27572 20626
rect 27632 20566 30476 20626
rect 25538 20560 25598 20566
rect 26556 20560 26616 20566
rect 27572 20560 27632 20566
rect 30476 20560 30536 20566
rect 30628 20628 30688 20634
rect 32662 20628 32722 20634
rect 33928 20628 33988 20634
rect 30688 20568 32662 20628
rect 32722 20568 33928 20628
rect 33988 20568 34770 20628
rect 30628 20562 30688 20568
rect 32662 20562 32722 20568
rect 33928 20562 33988 20568
rect 13060 20380 13120 20386
rect 14782 20380 14842 20386
rect 15216 20380 15276 20386
rect 15652 20380 15712 20386
rect 16088 20380 16148 20386
rect 16526 20380 16586 20386
rect 13120 20320 14782 20380
rect 14842 20320 15216 20380
rect 15276 20320 15652 20380
rect 15712 20320 16088 20380
rect 16148 20320 16526 20380
rect 13060 20314 13120 20320
rect 14782 20314 14842 20320
rect 15216 20314 15276 20320
rect 15652 20314 15712 20320
rect 16088 20314 16148 20320
rect 16526 20314 16586 20320
rect 14998 20276 15058 20282
rect 15434 20276 15494 20282
rect 15872 20276 15932 20282
rect 16306 20276 16366 20282
rect 15058 20216 15434 20276
rect 15494 20216 15872 20276
rect 15932 20216 16306 20276
rect 14998 20210 15058 20216
rect 15434 20210 15494 20216
rect 15872 20210 15932 20216
rect 16306 20210 16366 20216
rect 14892 20178 14952 20184
rect 15106 20178 15166 20184
rect 15326 20178 15386 20184
rect 15544 20178 15604 20184
rect 15654 20178 15714 20184
rect 15760 20178 15820 20184
rect 15978 20178 16038 20184
rect 16196 20178 16256 20184
rect 16412 20178 16472 20184
rect 14952 20118 15106 20178
rect 15166 20118 15326 20178
rect 15386 20118 15544 20178
rect 15604 20118 15654 20178
rect 15714 20118 15760 20178
rect 15820 20118 15978 20178
rect 16038 20118 16196 20178
rect 16256 20118 16412 20178
rect 14892 20112 14952 20118
rect 15106 20112 15166 20118
rect 15326 20112 15386 20118
rect 15544 20112 15604 20118
rect 15654 20112 15714 20118
rect 15760 20112 15820 20118
rect 15978 20112 16038 20118
rect 16196 20112 16256 20118
rect 16412 20112 16472 20118
rect 19430 19676 19490 19682
rect 21466 19676 21526 19682
rect 17864 19616 19430 19676
rect 19490 19616 21466 19676
rect 10196 7356 11048 7416
rect 11108 7356 12340 7416
rect 12418 19482 14442 19542
rect 14502 19482 14508 19542
rect 10136 7350 10196 7356
rect 11048 7350 11108 7356
rect 9266 7306 9326 7312
rect 10928 7306 10988 7312
rect 9326 7246 10928 7306
rect 9266 7240 9326 7246
rect 10928 7240 10988 7246
rect 8352 7198 8412 7204
rect 10030 7198 10090 7204
rect 10248 7198 10308 7204
rect 11382 7198 11442 7207
rect 8412 7138 10030 7198
rect 10090 7138 10248 7198
rect 10308 7138 11382 7198
rect 8352 7132 8412 7138
rect 10030 7132 10090 7138
rect 10248 7132 10308 7138
rect 11382 7129 11442 7138
rect 8482 7090 8542 7096
rect 9812 7090 9872 7096
rect 10466 7090 10526 7096
rect 8542 7030 9812 7090
rect 9872 7030 10466 7090
rect 8482 7024 8542 7030
rect 9812 7024 9872 7030
rect 10466 7024 10526 7030
rect 12418 6816 12478 19482
rect 14782 19442 14842 19448
rect 15652 19442 15712 19448
rect 16526 19442 16586 19448
rect 16882 19442 16942 19448
rect 10922 6756 10928 6816
rect 10988 6756 12478 6816
rect 12536 19382 14782 19442
rect 14842 19382 15652 19442
rect 15712 19382 16526 19442
rect 16586 19382 16882 19442
rect 8940 6590 9000 6596
rect 9596 6590 9656 6596
rect 10466 6590 10526 6596
rect 11170 6590 11230 6596
rect 9000 6530 9596 6590
rect 9656 6530 10466 6590
rect 10526 6530 11170 6590
rect 8940 6524 9000 6530
rect 9596 6524 9656 6530
rect 10466 6524 10526 6530
rect 11170 6524 11230 6530
rect 9048 6490 9108 6496
rect 9486 6490 9546 6496
rect 7854 6430 9048 6490
rect 9108 6430 9486 6490
rect 9546 6430 9982 6490
rect 3564 4940 3624 4946
rect 5604 4940 5664 4946
rect 3624 4880 5604 4940
rect 3564 4874 3624 4880
rect 5604 4874 5664 4880
rect 1412 4036 1472 4042
rect 2550 4036 2610 4042
rect 6624 4036 6684 4042
rect 1472 3976 2550 4036
rect 2610 3976 6624 4036
rect 1412 3970 1472 3976
rect 2550 3970 2610 3976
rect 6624 3970 6684 3976
rect 3564 3940 3624 3946
rect 5604 3940 5664 3946
rect 3624 3880 5604 3940
rect 3564 3874 3624 3880
rect 5604 3874 5664 3880
rect -10820 3835 -10716 3840
rect -10824 3741 -10815 3835
rect -10721 3741 -10712 3835
rect -6742 3827 -6642 3832
rect -10820 3688 -10716 3741
rect -6746 3737 -6737 3827
rect -6647 3737 -6638 3827
rect 4586 3824 4646 3830
rect 7748 3824 7808 3830
rect 4646 3764 7748 3824
rect 4586 3758 4646 3764
rect 7748 3758 7808 3764
rect -10820 3584 -8906 3688
rect -6742 3686 -6642 3737
rect -6742 3586 -4536 3686
rect -9010 3514 -8906 3584
rect -9010 3401 -8906 3410
rect -4636 3510 -4536 3586
rect -4636 3401 -4536 3410
rect 2696 2924 2756 2930
rect 4582 2924 4642 2930
rect 6452 2924 6512 2930
rect 7854 2924 7914 6430
rect 9048 6424 9108 6430
rect 9486 6424 9546 6430
rect 7974 6380 8034 6386
rect 9050 6380 9110 6386
rect 9484 6380 9544 6386
rect 9812 6380 9872 6386
rect 8034 6320 9050 6380
rect 9110 6320 9484 6380
rect 9544 6320 9812 6380
rect 7974 6314 8034 6320
rect 9050 6314 9110 6320
rect 9484 6314 9544 6320
rect 9812 6314 9872 6320
rect 9922 6380 9982 6430
rect 10576 6470 10636 6476
rect 12536 6470 12596 19382
rect 14782 19376 14842 19382
rect 15652 19376 15712 19382
rect 16526 19376 16586 19382
rect 16882 19376 16942 19382
rect 14998 19344 15058 19350
rect 15434 19344 15494 19350
rect 15872 19344 15932 19350
rect 16306 19344 16366 19350
rect 15058 19284 15434 19344
rect 15494 19284 15872 19344
rect 15932 19284 16306 19344
rect 14998 19278 15058 19284
rect 15434 19278 15494 19284
rect 15872 19278 15932 19284
rect 16306 19278 16366 19284
rect 14442 19226 14502 19232
rect 15108 19226 15168 19232
rect 15216 19226 15276 19232
rect 15324 19226 15384 19232
rect 15970 19226 16030 19232
rect 16088 19226 16148 19232
rect 14502 19166 15108 19226
rect 15168 19166 15216 19226
rect 15276 19166 15324 19226
rect 15384 19166 15970 19226
rect 16030 19166 16088 19226
rect 16197 19224 16255 19230
rect 16148 19166 16197 19224
rect 14442 19160 14502 19166
rect 15108 19160 15168 19166
rect 15216 19160 15276 19166
rect 15324 19160 15384 19166
rect 15970 19160 16030 19166
rect 16088 19160 16148 19166
rect 16197 19160 16255 19166
rect 13268 18823 13277 18913
rect 13367 18823 13376 18913
rect 13060 18148 13120 18154
rect 12898 17982 12904 18042
rect 12964 17982 12970 18042
rect 12646 16327 12655 16417
rect 12745 16327 12754 16417
rect 12670 15064 12730 16327
rect 12904 15192 12964 17982
rect 12904 15126 12964 15132
rect 13060 15192 13120 18088
rect 13286 15184 13346 18823
rect 14782 18506 14842 18512
rect 14892 18506 14952 18512
rect 15546 18506 15606 18512
rect 15652 18506 15712 18512
rect 15762 18506 15822 18512
rect 16414 18506 16474 18512
rect 16526 18506 16586 18512
rect 16998 18506 17058 18512
rect 14842 18446 14892 18506
rect 14952 18446 15546 18506
rect 15606 18446 15652 18506
rect 15712 18446 15762 18506
rect 15822 18446 16414 18506
rect 16474 18446 16526 18506
rect 16586 18446 16998 18506
rect 14782 18440 14842 18446
rect 14892 18440 14952 18446
rect 15546 18440 15606 18446
rect 15652 18440 15712 18446
rect 15762 18440 15822 18446
rect 16414 18440 16474 18446
rect 16526 18440 16586 18446
rect 16998 18440 17058 18446
rect 13060 15126 13120 15132
rect 13280 15124 13286 15184
rect 13346 15124 13352 15184
rect 17864 15064 17924 19616
rect 19430 19610 19490 19616
rect 21466 19610 21526 19616
rect 24520 19678 24580 19684
rect 26556 19678 26616 19684
rect 24580 19618 26556 19678
rect 24520 19612 24580 19618
rect 26556 19612 26616 19618
rect 29610 19680 29670 19686
rect 31646 19680 31706 19686
rect 29670 19620 31646 19680
rect 29610 19614 29670 19620
rect 31646 19614 31706 19620
rect 21466 19568 21526 19574
rect 33796 19568 33856 19574
rect 21526 19508 33796 19568
rect 21466 19502 21526 19508
rect 33796 19502 33856 19508
rect 18262 19468 18322 19474
rect 18322 19408 30846 19468
rect 18262 19402 18322 19408
rect 22682 19372 22742 19378
rect 20444 19366 20504 19372
rect 22478 19366 22538 19372
rect 20504 19306 22478 19366
rect 22742 19312 24516 19372
rect 24576 19312 24582 19372
rect 25536 19368 25596 19374
rect 27570 19368 27630 19374
rect 22682 19306 22742 19312
rect 25596 19308 27570 19368
rect 20444 19300 20504 19306
rect 22478 19300 22538 19306
rect 25536 19302 25596 19308
rect 27570 19302 27630 19308
rect 27784 19364 27844 19370
rect 30632 19366 30692 19372
rect 30786 19366 30846 19408
rect 32666 19366 32726 19372
rect 27844 19304 30120 19364
rect 30180 19304 30186 19364
rect 30692 19306 32666 19366
rect 27784 19298 27844 19304
rect 30632 19300 30692 19306
rect 32666 19300 32726 19306
rect 17994 18418 18054 18424
rect 19426 18418 19486 18424
rect 21462 18418 21522 18424
rect 18054 18358 19426 18418
rect 19486 18358 21462 18418
rect 17994 18352 18054 18358
rect 19426 18352 19486 18358
rect 21462 18352 21522 18358
rect 29614 18418 29674 18424
rect 31650 18418 31710 18424
rect 29674 18358 31650 18418
rect 29614 18352 29674 18358
rect 18130 18288 18190 18294
rect 29744 18288 29804 18358
rect 31650 18352 31710 18358
rect 18190 18228 29804 18288
rect 18130 18222 18190 18228
rect 22484 18148 22544 18154
rect 34088 18148 34148 18154
rect 22544 18088 34088 18148
rect 22484 18082 22544 18088
rect 12670 15004 17924 15064
rect 12670 10080 12730 15004
rect 12800 14092 12860 14098
rect 13518 14092 13578 14098
rect 15554 14092 15614 14098
rect 17588 14092 17648 14098
rect 19628 14092 19688 14098
rect 21664 14092 21724 14098
rect 23698 14092 23758 14098
rect 25734 14092 25794 14098
rect 27770 14092 27830 14098
rect 29806 14092 29866 14098
rect 31844 14092 31904 14098
rect 33874 14092 33934 14098
rect 12860 14032 13518 14092
rect 13578 14032 15554 14092
rect 15614 14032 17588 14092
rect 17648 14032 19628 14092
rect 19688 14032 21664 14092
rect 21724 14032 23698 14092
rect 23758 14032 25734 14092
rect 25794 14032 27770 14092
rect 27830 14032 29806 14092
rect 29866 14032 31844 14092
rect 31904 14032 33874 14092
rect 12800 14026 12860 14032
rect 13518 14026 13578 14032
rect 15554 14026 15614 14032
rect 17588 14026 17648 14032
rect 19628 14026 19688 14032
rect 21664 14026 21724 14032
rect 23698 14026 23758 14032
rect 25734 14026 25794 14032
rect 27770 14026 27830 14032
rect 29806 14026 29866 14032
rect 31844 14026 31904 14032
rect 33874 14026 33934 14032
rect 14536 13994 14596 14000
rect 16574 13994 16634 14000
rect 18608 13994 18668 14000
rect 20642 13994 20702 14000
rect 22682 13994 22742 14000
rect 24716 13994 24776 14000
rect 26754 13994 26814 14000
rect 28786 13994 28846 14000
rect 30824 13994 30884 14000
rect 32862 13994 32922 14000
rect 33996 13994 34056 18088
rect 34088 18082 34148 18088
rect 34598 13994 34658 14000
rect 14596 13934 16574 13994
rect 16634 13934 18608 13994
rect 18668 13934 20642 13994
rect 20702 13934 22682 13994
rect 22742 13934 24716 13994
rect 24776 13934 26754 13994
rect 26814 13934 28786 13994
rect 28846 13934 30824 13994
rect 30884 13934 32862 13994
rect 32922 13934 34598 13994
rect 14536 13928 14596 13934
rect 16574 13928 16634 13934
rect 18608 13928 18668 13934
rect 20642 13928 20702 13934
rect 22682 13928 22742 13934
rect 24716 13928 24776 13934
rect 26754 13928 26814 13934
rect 28786 13928 28846 13934
rect 30824 13928 30884 13934
rect 32862 13928 32922 13934
rect 34598 13928 34658 13934
rect 22682 13782 22742 13788
rect 24714 13782 24774 13788
rect 22742 13722 24714 13782
rect 22682 13716 22742 13722
rect 24714 13716 24774 13722
rect 17222 12862 17282 12868
rect 17592 12862 17652 12868
rect 18094 12862 18154 12868
rect 18606 12862 18666 12868
rect 19134 12862 19194 12868
rect 19626 12862 19686 12868
rect 21658 12862 21718 12868
rect 23694 12862 23754 12868
rect 25730 12862 25790 12868
rect 27768 12862 27828 12868
rect 29806 12862 29866 12868
rect 30314 12862 30374 12868
rect 17282 12802 17592 12862
rect 17652 12802 18094 12862
rect 18154 12802 18606 12862
rect 18666 12802 19134 12862
rect 19194 12802 19626 12862
rect 19686 12802 21658 12862
rect 21718 12802 23694 12862
rect 23754 12802 25730 12862
rect 25790 12802 27768 12862
rect 27828 12802 29292 12862
rect 29352 12802 29806 12862
rect 29866 12802 30314 12862
rect 17222 12796 17282 12802
rect 17592 12796 17652 12802
rect 18094 12796 18154 12802
rect 18606 12796 18666 12802
rect 19134 12796 19194 12802
rect 19626 12796 19686 12802
rect 21658 12796 21718 12802
rect 23694 12796 23754 12802
rect 25730 12796 25790 12802
rect 27768 12796 27828 12802
rect 29806 12796 29866 12802
rect 30314 12796 30374 12802
rect 15046 12752 15106 12758
rect 16068 12752 16128 12758
rect 20140 12752 20200 12758
rect 20644 12752 20704 12758
rect 21160 12752 21220 12758
rect 22180 12752 22240 12758
rect 22682 12752 22742 12758
rect 23182 12752 23242 12758
rect 24208 12752 24268 12758
rect 24718 12752 24778 12758
rect 25226 12752 25286 12758
rect 26234 12752 26294 12758
rect 26756 12752 26816 12758
rect 27246 12752 27306 12758
rect 28278 12752 28338 12758
rect 28790 12752 28850 12758
rect 31334 12752 31394 12758
rect 32354 12752 32414 12758
rect 13056 12692 13062 12752
rect 13122 12692 15046 12752
rect 15106 12692 16068 12752
rect 16128 12692 20140 12752
rect 20200 12692 20644 12752
rect 20704 12692 21160 12752
rect 21220 12692 22180 12752
rect 22240 12692 22682 12752
rect 22742 12692 23182 12752
rect 23242 12692 24208 12752
rect 24268 12692 24718 12752
rect 24778 12692 25226 12752
rect 25286 12692 26234 12752
rect 26294 12692 26756 12752
rect 26816 12692 27246 12752
rect 27306 12692 28278 12752
rect 28338 12692 28790 12752
rect 28850 12692 31334 12752
rect 31394 12692 32354 12752
rect 15046 12686 15106 12692
rect 16068 12686 16128 12692
rect 20140 12686 20200 12692
rect 20644 12686 20704 12692
rect 21160 12686 21220 12692
rect 22180 12686 22240 12692
rect 22682 12686 22742 12692
rect 23182 12686 23242 12692
rect 24208 12686 24268 12692
rect 24718 12686 24778 12692
rect 25226 12686 25286 12692
rect 26234 12686 26294 12692
rect 26756 12686 26816 12692
rect 27246 12686 27306 12692
rect 28278 12686 28338 12692
rect 28790 12686 28850 12692
rect 31334 12686 31394 12692
rect 32354 12686 32414 12692
rect 18088 12648 18148 12654
rect 19108 12648 19168 12654
rect 23322 12648 23382 12654
rect 24330 12648 24390 12654
rect 25372 12648 25432 12654
rect 28264 12648 28324 12654
rect 29302 12648 29362 12654
rect 30302 12648 30362 12654
rect 17082 12588 17088 12648
rect 17148 12588 18088 12648
rect 18148 12588 19108 12648
rect 19168 12588 23322 12648
rect 23382 12588 24330 12648
rect 24390 12588 25372 12648
rect 25432 12588 28264 12648
rect 28324 12588 29302 12648
rect 29362 12588 30302 12648
rect 18088 12582 18148 12588
rect 19108 12582 19168 12588
rect 23322 12582 23382 12588
rect 24330 12582 24390 12588
rect 25372 12582 25432 12588
rect 28264 12582 28324 12588
rect 29302 12582 29362 12588
rect 30302 12582 30362 12588
rect 12926 12540 12986 12546
rect 13522 12540 13582 12546
rect 14020 12540 14080 12546
rect 14532 12540 14592 12546
rect 16574 12540 16634 12546
rect 18608 12540 18668 12546
rect 20642 12540 20702 12546
rect 26756 12540 26816 12546
rect 28788 12540 28848 12546
rect 30820 12540 30880 12546
rect 32862 12540 32922 12546
rect 33366 12540 33426 12546
rect 33876 12540 33936 12546
rect 12986 12480 13522 12540
rect 13582 12480 14020 12540
rect 14080 12480 14532 12540
rect 14592 12480 16574 12540
rect 16634 12480 18608 12540
rect 18668 12480 20642 12540
rect 20702 12480 22798 12540
rect 22858 12538 26756 12540
rect 22858 12480 24522 12538
rect 12926 12474 12986 12480
rect 13522 12474 13582 12480
rect 14020 12474 14080 12480
rect 14532 12474 14592 12480
rect 16574 12474 16634 12480
rect 18608 12474 18668 12480
rect 20642 12474 20702 12480
rect 24516 12478 24522 12480
rect 24582 12480 26756 12538
rect 26816 12480 28788 12540
rect 28848 12480 30820 12540
rect 30880 12480 32862 12540
rect 32922 12480 33366 12540
rect 33426 12480 33876 12540
rect 24582 12478 24588 12480
rect 26756 12474 26816 12480
rect 28788 12474 28848 12480
rect 30820 12474 30880 12480
rect 32862 12474 32922 12480
rect 33366 12474 33426 12480
rect 33876 12474 33936 12480
rect 16052 11650 16112 11656
rect 17072 11650 17132 11656
rect 18084 11650 18144 11656
rect 19110 11650 19170 11656
rect 28266 11650 28326 11656
rect 29302 11650 29362 11656
rect 30318 11650 30378 11656
rect 12800 11638 12860 11644
rect 15036 11638 15096 11644
rect 12860 11578 15036 11638
rect 16112 11590 17072 11650
rect 17132 11590 18084 11650
rect 18144 11590 19110 11650
rect 19170 11590 28266 11650
rect 28326 11590 29302 11650
rect 29362 11590 30318 11650
rect 16052 11584 16112 11590
rect 17072 11584 17132 11590
rect 18084 11584 18144 11590
rect 19110 11584 19170 11590
rect 28266 11584 28326 11590
rect 29302 11584 29362 11590
rect 30318 11584 30378 11590
rect 12800 11572 12860 11578
rect 15036 11572 15096 11578
rect 15548 11546 15608 11552
rect 16572 11546 16632 11552
rect 17584 11546 17644 11552
rect 18604 11546 18664 11552
rect 19626 11546 19686 11552
rect 21662 11546 21722 11552
rect 23700 11546 23760 11552
rect 25730 11546 25790 11552
rect 26750 11546 26810 11552
rect 27768 11546 27828 11552
rect 28788 11546 28848 11552
rect 29804 11546 29864 11552
rect 31840 11546 31900 11552
rect 15608 11486 16572 11546
rect 16632 11486 17584 11546
rect 17644 11486 18604 11546
rect 18664 11486 19626 11546
rect 19686 11486 21662 11546
rect 21722 11486 23700 11546
rect 23760 11486 25730 11546
rect 25790 11486 26750 11546
rect 26810 11486 27768 11546
rect 27828 11486 28788 11546
rect 28848 11486 29804 11546
rect 29864 11486 31840 11546
rect 15548 11480 15608 11486
rect 16572 11480 16632 11486
rect 17584 11480 17644 11486
rect 18604 11480 18664 11486
rect 19626 11480 19686 11486
rect 21662 11480 21722 11486
rect 23700 11480 23760 11486
rect 25730 11480 25790 11486
rect 26750 11480 26810 11486
rect 27768 11480 27828 11486
rect 28788 11480 28848 11486
rect 29804 11480 29864 11486
rect 31840 11480 31900 11486
rect 13286 11424 13346 11430
rect 20646 11424 20706 11430
rect 22680 11424 22740 11430
rect 24710 11424 24770 11430
rect 34710 11424 34770 20568
rect 13346 11364 20646 11424
rect 20706 11364 22680 11424
rect 22740 11364 24710 11424
rect 24770 11364 34770 11424
rect 13286 11358 13346 11364
rect 20646 11358 20706 11364
rect 22680 11358 22740 11364
rect 24710 11358 24770 11364
rect 15554 11312 15614 11318
rect 17590 11312 17650 11318
rect 33984 11312 34044 11318
rect 15614 11252 17590 11312
rect 17650 11252 33984 11312
rect 15554 11246 15614 11252
rect 17590 11246 17650 11252
rect 33984 11246 34044 11252
rect 33878 10424 33938 10430
rect 34838 10424 34898 20886
rect 36254 16193 36354 21314
rect 40228 21305 40328 21314
rect 65088 18913 65188 18918
rect 65084 18823 65093 18913
rect 65183 18823 65192 18913
rect 43134 17841 43262 17846
rect 38968 17829 39076 17834
rect 38964 17731 38973 17829
rect 39071 17731 39080 17829
rect 38968 17668 39076 17731
rect 43130 17723 43139 17841
rect 43257 17723 43266 17841
rect 47326 17831 47436 17836
rect 47322 17731 47331 17831
rect 47431 17731 47440 17831
rect 43134 17694 43262 17723
rect 38968 17560 41102 17668
rect 43134 17566 45316 17694
rect 40994 17516 41102 17560
rect 40994 17399 41102 17408
rect 45188 17526 45316 17566
rect 47326 17669 47436 17731
rect 47326 17559 49393 17669
rect 45188 17389 45316 17398
rect 49283 17507 49393 17559
rect 49283 17388 49393 17397
rect 36250 16103 36259 16193
rect 36349 16103 36358 16193
rect 36254 16098 36354 16103
rect 52918 15362 53018 15368
rect 54712 15362 54812 15368
rect 57312 15362 57412 15368
rect 59912 15364 60012 15370
rect 62512 15364 62612 15370
rect 64316 15364 64416 15370
rect 52914 15267 52918 15357
rect 53018 15267 53022 15357
rect 54708 15267 54712 15357
rect 54812 15267 54816 15357
rect 57308 15267 57312 15357
rect 57412 15267 57416 15357
rect 59908 15269 59912 15359
rect 60012 15269 60016 15359
rect 62508 15269 62512 15359
rect 62612 15269 62616 15359
rect 64312 15269 64316 15359
rect 64416 15269 64420 15359
rect 52918 15256 53018 15262
rect 54712 15256 54812 15262
rect 57312 15256 57412 15262
rect 59912 15258 60012 15264
rect 62512 15258 62612 15264
rect 64316 15258 64416 15264
rect 65088 14738 65188 18823
rect 65079 14638 65088 14738
rect 65188 14638 65197 14738
rect 36456 13814 36556 13823
rect 39253 13814 39343 13818
rect 36556 13809 39348 13814
rect 36556 13719 39253 13809
rect 39343 13719 39348 13809
rect 36556 13714 39348 13719
rect 36456 13705 36556 13714
rect 39253 13710 39343 13714
rect 42994 11727 43130 11732
rect 38844 11711 38950 11716
rect 38840 11615 38849 11711
rect 38945 11615 38954 11711
rect 38844 11553 38950 11615
rect 42990 11597 42999 11727
rect 43125 11597 43134 11727
rect 42994 11590 43134 11597
rect 38844 11447 40991 11553
rect 42994 11454 45158 11590
rect 40885 11381 40991 11447
rect 45050 11392 45158 11454
rect 45050 11275 45158 11284
rect 40885 11266 40991 11275
rect 16570 10406 16630 10412
rect 18606 10406 18666 10412
rect 26750 10406 26810 10412
rect 28786 10406 28846 10412
rect 32860 10406 32920 10412
rect 13398 10382 13458 10388
rect 14536 10382 14596 10388
rect 13458 10322 14536 10382
rect 14596 10322 15418 10382
rect 16630 10346 18606 10406
rect 18666 10346 26750 10406
rect 26810 10346 28786 10406
rect 28846 10346 32860 10406
rect 33938 10364 34898 10424
rect 33878 10358 33938 10364
rect 16570 10340 16630 10346
rect 18606 10340 18666 10346
rect 26750 10340 26810 10346
rect 28786 10340 28846 10346
rect 32860 10340 32920 10346
rect 13398 10316 13458 10322
rect 14536 10316 14596 10322
rect 13286 10182 13346 10188
rect 14534 10182 14594 10188
rect 13346 10122 14534 10182
rect 15358 10186 15418 10322
rect 15552 10302 15612 10308
rect 17592 10302 17652 10308
rect 19624 10302 19684 10308
rect 21658 10302 21718 10308
rect 23698 10302 23758 10308
rect 25732 10302 25792 10308
rect 15612 10242 17592 10302
rect 17652 10242 19624 10302
rect 19684 10242 21658 10302
rect 21718 10242 23698 10302
rect 23758 10242 25732 10302
rect 15552 10236 15612 10242
rect 17592 10236 17652 10242
rect 19624 10236 19684 10242
rect 21658 10236 21718 10242
rect 23698 10236 23758 10242
rect 25732 10236 25792 10242
rect 25928 10298 25988 10304
rect 30820 10298 30880 10304
rect 25988 10238 30820 10298
rect 34478 10294 34538 10300
rect 25928 10232 25988 10238
rect 30820 10232 30880 10238
rect 31318 10234 31324 10294
rect 31384 10234 34478 10294
rect 34478 10228 34538 10234
rect 16066 10188 16126 10194
rect 19624 10190 19684 10196
rect 21660 10190 21720 10196
rect 23696 10190 23756 10196
rect 25732 10190 25792 10196
rect 27766 10190 27826 10196
rect 29804 10190 29864 10196
rect 31844 10190 31904 10196
rect 34228 10190 34288 10196
rect 15358 10128 16066 10186
rect 16126 10128 17070 10188
rect 17130 10128 18082 10188
rect 18142 10128 19102 10188
rect 19162 10128 19168 10188
rect 19684 10130 21660 10190
rect 21720 10130 23696 10190
rect 23756 10130 25732 10190
rect 25792 10130 27766 10190
rect 27826 10130 29804 10190
rect 29864 10130 31844 10190
rect 31904 10130 34228 10190
rect 15358 10126 16408 10128
rect 16066 10122 16126 10126
rect 19624 10124 19684 10130
rect 21660 10124 21720 10130
rect 23696 10124 23756 10130
rect 25732 10124 25792 10130
rect 27766 10124 27826 10130
rect 29804 10124 29864 10130
rect 31844 10124 31904 10130
rect 34228 10124 34288 10130
rect 13286 10116 13346 10122
rect 14534 10116 14594 10122
rect 13180 10080 13240 10086
rect 20642 10080 20702 10086
rect 22676 10080 22736 10086
rect 24716 10080 24776 10086
rect 25928 10080 25988 10086
rect 12670 10020 13180 10080
rect 13240 10020 20642 10080
rect 20702 10020 22676 10080
rect 22736 10020 24716 10080
rect 24776 10020 25928 10080
rect 13180 10014 13240 10020
rect 20642 10014 20702 10020
rect 22676 10014 22736 10020
rect 24716 10014 24776 10020
rect 25928 10014 25988 10020
rect 26222 10082 26282 10088
rect 26282 10022 27250 10082
rect 27310 10022 27316 10082
rect 27768 10076 27828 10082
rect 29804 10076 29864 10082
rect 31842 10076 31902 10082
rect 33984 10076 34044 10082
rect 26222 10016 26282 10022
rect 27828 10016 29804 10076
rect 29864 10016 31842 10076
rect 31902 10016 33984 10076
rect 27768 10010 27828 10016
rect 29804 10010 29864 10016
rect 31842 10010 31902 10016
rect 33984 10010 34044 10016
rect 36060 9306 36160 9315
rect 39009 9306 39099 9310
rect 36056 9206 36060 9306
rect 36160 9301 39104 9306
rect 36160 9211 39009 9301
rect 39099 9211 39104 9301
rect 36160 9206 39104 9211
rect 36060 9197 36160 9206
rect 39009 9202 39099 9206
rect 30316 9162 30376 9168
rect 14534 9150 14594 9156
rect 16572 9150 16632 9156
rect 18608 9150 18668 9156
rect 20640 9150 20700 9156
rect 14594 9090 16572 9150
rect 16632 9090 18608 9150
rect 18668 9090 20640 9150
rect 25216 9102 25222 9162
rect 25282 9102 30316 9162
rect 30316 9096 30376 9102
rect 30454 9166 30514 9172
rect 31336 9166 31396 9172
rect 32342 9166 32402 9172
rect 30514 9106 31336 9166
rect 31396 9106 32342 9166
rect 30454 9100 30514 9106
rect 31336 9100 31396 9106
rect 32342 9100 32402 9106
rect 32860 9162 32920 9168
rect 34112 9162 34172 9168
rect 32920 9102 34112 9162
rect 35833 9132 35935 9136
rect 32860 9096 32920 9102
rect 34112 9096 34172 9102
rect 35828 9127 51026 9132
rect 14534 9084 14594 9090
rect 16572 9084 16632 9090
rect 18608 9084 18668 9090
rect 20640 9084 20700 9090
rect 15040 9048 15100 9054
rect 20132 9048 20192 9054
rect 15100 8988 20132 9048
rect 15040 8982 15100 8988
rect 20132 8982 20192 8988
rect 24716 9034 24776 9040
rect 32860 9034 32920 9040
rect 24776 8974 32860 9034
rect 35828 9025 35833 9127
rect 35935 9108 51026 9127
rect 35935 9048 50944 9108
rect 51004 9048 51026 9108
rect 35935 9025 51026 9048
rect 35828 9020 51026 9025
rect 35833 9016 35935 9020
rect 24716 8968 24776 8974
rect 32860 8968 32920 8974
rect 13286 8946 13346 8952
rect 16570 8946 16630 8952
rect 13346 8886 16570 8946
rect 13286 8880 13346 8886
rect 16570 8880 16630 8886
rect 17078 8940 17138 8946
rect 18100 8940 18160 8946
rect 19114 8940 19174 8946
rect 20132 8940 20192 8946
rect 21152 8940 21212 8946
rect 28264 8940 28324 8946
rect 29294 8940 29354 8946
rect 30454 8940 30514 8946
rect 17138 8880 18100 8940
rect 18160 8880 19114 8940
rect 19174 8880 20132 8940
rect 20192 8880 21152 8940
rect 21212 8880 28264 8940
rect 28324 8880 29294 8940
rect 29354 8880 30454 8940
rect 17078 8874 17138 8880
rect 18100 8874 18160 8880
rect 19114 8874 19174 8880
rect 20132 8874 20192 8880
rect 21152 8874 21212 8880
rect 28264 8874 28324 8880
rect 29294 8874 29354 8880
rect 30454 8874 30514 8880
rect 30822 8940 30882 8946
rect 34350 8940 34410 8946
rect 30882 8880 34350 8940
rect 30822 8874 30882 8880
rect 34350 8874 34410 8880
rect 15554 8846 15614 8852
rect 17588 8846 17648 8852
rect 19624 8846 19684 8852
rect 15614 8786 17588 8846
rect 17648 8786 19624 8846
rect 15554 8780 15614 8786
rect 17588 8780 17648 8786
rect 19624 8780 19684 8786
rect 26752 8836 26812 8842
rect 30822 8836 30882 8842
rect 26812 8776 30822 8836
rect 26752 8770 26812 8776
rect 30822 8770 30882 8776
rect 31838 8838 31898 8844
rect 34228 8838 34288 8844
rect 31898 8778 34228 8838
rect 31838 8772 31898 8778
rect 34228 8772 34288 8778
rect 49948 8406 49954 8466
rect 50014 8406 50613 8466
rect 21660 7928 21720 7934
rect 23696 7928 23756 7934
rect 25732 7928 25792 7934
rect 27770 7928 27830 7934
rect 15036 7922 15096 7928
rect 15946 7922 16006 7928
rect 16948 7922 17008 7928
rect 18100 7922 18160 7928
rect 19110 7922 19170 7928
rect 20116 7922 20176 7928
rect 21160 7922 21220 7928
rect 15096 7862 15946 7922
rect 16006 7862 16948 7922
rect 17008 7862 18100 7922
rect 18160 7862 19110 7922
rect 19170 7862 20116 7922
rect 20176 7862 21160 7922
rect 21720 7868 23696 7928
rect 23756 7868 25732 7928
rect 25792 7868 27770 7928
rect 21660 7862 21720 7868
rect 23696 7862 23756 7868
rect 25732 7862 25792 7868
rect 27770 7862 27830 7868
rect 29806 7928 29866 7934
rect 31844 7928 31904 7934
rect 29866 7868 31844 7928
rect 29806 7862 29866 7868
rect 31844 7862 31904 7868
rect 15036 7856 15096 7862
rect 15946 7856 16006 7862
rect 16948 7856 17008 7862
rect 18100 7856 18160 7862
rect 19110 7856 19170 7862
rect 20116 7856 20176 7862
rect 21160 7856 21220 7862
rect 17588 7820 17648 7826
rect 27762 7820 27822 7826
rect 29802 7820 29862 7826
rect 31840 7820 31900 7826
rect 17648 7760 27762 7820
rect 27822 7760 29802 7820
rect 29862 7760 31840 7820
rect 17588 7754 17648 7760
rect 27762 7754 27822 7760
rect 29802 7754 29862 7760
rect 31840 7754 31900 7760
rect 15036 7706 15096 7712
rect 17088 7706 17148 7712
rect 20114 7706 20174 7712
rect 21154 7706 21214 7712
rect 22168 7706 22228 7712
rect 23176 7706 23236 7712
rect 24220 7706 24280 7712
rect 25210 7706 25270 7712
rect 26228 7706 26288 7712
rect 27262 7706 27322 7712
rect 30294 7706 30354 7712
rect 31332 7706 31392 7712
rect 32358 7706 32418 7712
rect 15096 7646 16074 7706
rect 16134 7646 17088 7706
rect 17148 7646 20114 7706
rect 20174 7646 21154 7706
rect 21214 7646 22168 7706
rect 22228 7646 23176 7706
rect 23236 7646 24220 7706
rect 24280 7646 25210 7706
rect 25270 7646 26228 7706
rect 26288 7646 27262 7706
rect 27322 7646 30294 7706
rect 30354 7646 31332 7706
rect 31392 7646 32358 7706
rect 32418 7646 34476 7706
rect 34536 7646 34542 7706
rect 49306 7700 49366 7706
rect 49824 7700 49884 7706
rect 15036 7640 15096 7646
rect 17088 7640 17148 7646
rect 20114 7640 20174 7646
rect 21154 7640 21214 7646
rect 22168 7640 22228 7646
rect 23176 7640 23236 7646
rect 24220 7640 24280 7646
rect 25210 7640 25270 7646
rect 26228 7640 26288 7646
rect 27262 7640 27322 7646
rect 30294 7640 30354 7646
rect 31332 7640 31392 7646
rect 32358 7640 32418 7646
rect 49366 7640 49822 7700
rect 49884 7640 49891 7700
rect 49306 7634 49366 7640
rect 49824 7634 49884 7640
rect 50553 7628 50613 8406
rect 65640 7652 65700 23362
rect 74476 23356 74540 23362
rect 76514 23236 76574 23242
rect 65902 23176 71866 23236
rect 71926 23176 76514 23236
rect 65902 7682 65962 23176
rect 76514 23170 76574 23176
rect 72262 23136 72322 23142
rect 73428 23136 73488 23142
rect 75464 23136 75524 23142
rect 72322 23076 73428 23136
rect 73488 23076 75464 23136
rect 72262 23070 72322 23076
rect 73428 23070 73488 23076
rect 75464 23070 75524 23076
rect 83610 23136 83670 23142
rect 85644 23136 85704 23142
rect 88088 23136 88148 23142
rect 83670 23076 85644 23136
rect 85704 23076 88088 23136
rect 83610 23070 83670 23076
rect 85644 23070 85704 23076
rect 88088 23070 88148 23076
rect 74446 22188 74506 22194
rect 76482 22188 76542 22194
rect 74506 22128 76482 22188
rect 74446 22122 74506 22128
rect 76482 22122 76542 22128
rect 84626 22188 84686 22194
rect 86662 22188 86722 22194
rect 84686 22128 86662 22188
rect 84626 22122 84686 22128
rect 71994 22090 72054 22096
rect 84734 22090 84794 22128
rect 86662 22122 86722 22128
rect 69106 22038 69166 22044
rect 69218 22038 69278 22044
rect 69328 22038 69388 22044
rect 69978 22038 70038 22044
rect 70088 22038 70148 22044
rect 70196 22038 70256 22044
rect 70998 22038 71058 22044
rect 66280 21978 69106 22038
rect 69166 21978 69218 22038
rect 69278 21978 69328 22038
rect 69388 21978 69978 22038
rect 70038 21978 70088 22038
rect 70148 21978 70196 22038
rect 70256 21978 70998 22038
rect 72054 22030 84794 22090
rect 71994 22024 72054 22030
rect 66128 17864 66134 17924
rect 66194 17864 66200 17924
rect 66134 14206 66194 17864
rect 66128 14146 66134 14206
rect 66194 14146 66200 14206
rect 20638 7602 20698 7608
rect 22680 7602 22740 7608
rect 24718 7602 24778 7608
rect 26752 7602 26812 7608
rect 28786 7604 28846 7610
rect 30820 7604 30880 7610
rect 32862 7604 32922 7610
rect 34112 7604 34172 7610
rect 13394 7542 13400 7602
rect 13460 7542 20638 7602
rect 20698 7542 22680 7602
rect 22740 7542 24718 7602
rect 24778 7542 26752 7602
rect 20638 7536 20698 7542
rect 22680 7536 22740 7542
rect 24718 7536 24778 7542
rect 26752 7536 26812 7542
rect 27264 7598 27324 7604
rect 28286 7598 28346 7604
rect 27324 7538 28286 7598
rect 28846 7544 30820 7604
rect 30880 7544 32862 7604
rect 32922 7544 34112 7604
rect 50553 7568 50627 7628
rect 50687 7568 50693 7628
rect 50939 7590 50945 7650
rect 51005 7590 51011 7650
rect 65634 7592 65640 7652
rect 65700 7592 65706 7652
rect 65896 7622 65902 7682
rect 65962 7622 65968 7682
rect 28786 7538 28846 7544
rect 30820 7538 30880 7544
rect 32862 7538 32922 7544
rect 34112 7538 34172 7544
rect 48364 7551 48424 7557
rect 49048 7551 49108 7557
rect 49564 7551 49624 7557
rect 27264 7532 27324 7538
rect 28286 7532 28346 7538
rect 48424 7491 49048 7551
rect 49108 7491 49564 7551
rect 49624 7491 50082 7551
rect 50142 7491 50148 7551
rect 48364 7485 48424 7491
rect 49048 7485 49108 7491
rect 49564 7485 49624 7491
rect 49952 7003 50012 7009
rect 50945 7004 51005 7590
rect 64136 7416 64196 7422
rect 65048 7416 65108 7422
rect 66280 7416 66340 21978
rect 69106 21972 69166 21978
rect 69218 21972 69278 21978
rect 69328 21972 69388 21978
rect 69978 21972 70038 21978
rect 70088 21972 70148 21978
rect 70196 21972 70256 21978
rect 70998 21972 71058 21978
rect 72130 21992 72190 21998
rect 74446 21992 74506 21998
rect 72190 21932 74446 21992
rect 72130 21926 72190 21932
rect 74446 21926 74506 21932
rect 75466 21994 75526 22000
rect 87928 21994 87988 22000
rect 75526 21934 87928 21994
rect 75466 21928 75526 21934
rect 87928 21928 87988 21934
rect 73432 21882 73492 21888
rect 75466 21882 75526 21888
rect 73492 21822 75466 21882
rect 73432 21816 73492 21822
rect 75466 21816 75526 21822
rect 78522 21880 78582 21886
rect 80556 21880 80616 21886
rect 78582 21820 80556 21880
rect 78522 21814 78582 21820
rect 80556 21814 80616 21820
rect 83612 21880 83672 21886
rect 85646 21882 85706 21886
rect 88240 21882 88304 23796
rect 85578 21880 88304 21882
rect 83672 21820 85646 21880
rect 85706 21820 88304 21880
rect 83612 21814 83672 21820
rect 85578 21818 88304 21820
rect 85646 21814 85706 21818
rect 68442 21326 68502 21332
rect 68782 21326 68842 21332
rect 68892 21326 68952 21332
rect 69542 21326 69602 21332
rect 69654 21326 69714 21332
rect 69762 21326 69822 21332
rect 70414 21326 70474 21332
rect 70524 21326 70584 21332
rect 68502 21266 68782 21326
rect 68842 21266 68892 21326
rect 68952 21266 69542 21326
rect 69602 21266 69654 21326
rect 69714 21266 69762 21326
rect 69822 21266 70414 21326
rect 70474 21266 70524 21326
rect 68442 21260 68502 21266
rect 68782 21260 68842 21266
rect 68892 21260 68952 21266
rect 69542 21260 69602 21266
rect 69654 21260 69714 21266
rect 69762 21260 69822 21266
rect 70414 21260 70474 21266
rect 70524 21260 70584 21266
rect 68998 21220 69058 21226
rect 69434 21220 69494 21226
rect 69872 21220 69932 21226
rect 70306 21220 70366 21226
rect 69058 21160 69434 21220
rect 69494 21160 69872 21220
rect 69932 21160 70306 21220
rect 68998 21154 69058 21160
rect 69434 21154 69494 21160
rect 69872 21154 69932 21160
rect 70306 21154 70366 21160
rect 69218 21104 69278 21110
rect 70088 21104 70148 21110
rect 70882 21104 70942 21110
rect 69278 21044 70088 21104
rect 70148 21044 70882 21104
rect 69218 21038 69278 21044
rect 70088 21038 70148 21044
rect 70882 21038 70942 21044
rect 84476 20946 84536 20952
rect 71752 20932 71812 20938
rect 78518 20932 78578 20938
rect 79538 20932 79598 20938
rect 81574 20932 81634 20938
rect 71812 20872 78518 20932
rect 78578 20872 79538 20932
rect 79598 20872 81574 20932
rect 84536 20886 88898 20946
rect 84476 20880 84536 20886
rect 71752 20866 71812 20872
rect 78518 20866 78578 20872
rect 79538 20866 79598 20872
rect 81574 20866 81634 20872
rect 84624 20836 84684 20842
rect 86664 20836 86724 20842
rect 87796 20836 87856 20842
rect 71866 20828 71926 20834
rect 76484 20828 76544 20834
rect 83608 20828 83668 20834
rect 71926 20768 74448 20828
rect 74508 20768 76484 20828
rect 76544 20768 83608 20828
rect 84684 20776 86664 20836
rect 86724 20776 87796 20836
rect 84624 20770 84684 20776
rect 86664 20770 86724 20776
rect 87796 20770 87856 20776
rect 71866 20762 71926 20768
rect 76484 20762 76544 20768
rect 83608 20762 83668 20768
rect 76482 20726 76542 20732
rect 85644 20726 85704 20732
rect 76542 20666 85644 20726
rect 76482 20660 76542 20666
rect 85644 20660 85704 20666
rect 74448 20624 74508 20630
rect 76482 20624 76542 20630
rect 74508 20564 76482 20624
rect 74448 20558 74508 20564
rect 76482 20558 76542 20564
rect 79538 20626 79598 20632
rect 80556 20626 80616 20632
rect 81572 20626 81632 20632
rect 84476 20626 84536 20632
rect 79598 20566 80556 20626
rect 80616 20566 81572 20626
rect 81632 20566 84476 20626
rect 79538 20560 79598 20566
rect 80556 20560 80616 20566
rect 81572 20560 81632 20566
rect 84476 20560 84536 20566
rect 84628 20628 84688 20634
rect 86662 20628 86722 20634
rect 87928 20628 87988 20634
rect 84688 20568 86662 20628
rect 86722 20568 87928 20628
rect 87988 20568 88770 20628
rect 84628 20562 84688 20568
rect 86662 20562 86722 20568
rect 87928 20562 87988 20568
rect 67060 20380 67120 20386
rect 68782 20380 68842 20386
rect 69216 20380 69276 20386
rect 69652 20380 69712 20386
rect 70088 20380 70148 20386
rect 70526 20380 70586 20386
rect 67120 20320 68782 20380
rect 68842 20320 69216 20380
rect 69276 20320 69652 20380
rect 69712 20320 70088 20380
rect 70148 20320 70526 20380
rect 67060 20314 67120 20320
rect 68782 20314 68842 20320
rect 69216 20314 69276 20320
rect 69652 20314 69712 20320
rect 70088 20314 70148 20320
rect 70526 20314 70586 20320
rect 68998 20276 69058 20282
rect 69434 20276 69494 20282
rect 69872 20276 69932 20282
rect 70306 20276 70366 20282
rect 69058 20216 69434 20276
rect 69494 20216 69872 20276
rect 69932 20216 70306 20276
rect 68998 20210 69058 20216
rect 69434 20210 69494 20216
rect 69872 20210 69932 20216
rect 70306 20210 70366 20216
rect 68892 20178 68952 20184
rect 69106 20178 69166 20184
rect 69326 20178 69386 20184
rect 69544 20178 69604 20184
rect 69654 20178 69714 20184
rect 69760 20178 69820 20184
rect 69978 20178 70038 20184
rect 70196 20178 70256 20184
rect 70412 20178 70472 20184
rect 68952 20118 69106 20178
rect 69166 20118 69326 20178
rect 69386 20118 69544 20178
rect 69604 20118 69654 20178
rect 69714 20118 69760 20178
rect 69820 20118 69978 20178
rect 70038 20118 70196 20178
rect 70256 20118 70412 20178
rect 68892 20112 68952 20118
rect 69106 20112 69166 20118
rect 69326 20112 69386 20118
rect 69544 20112 69604 20118
rect 69654 20112 69714 20118
rect 69760 20112 69820 20118
rect 69978 20112 70038 20118
rect 70196 20112 70256 20118
rect 70412 20112 70472 20118
rect 73430 19676 73490 19682
rect 75466 19676 75526 19682
rect 71864 19616 73430 19676
rect 73490 19616 75466 19676
rect 64196 7356 65048 7416
rect 65108 7356 66340 7416
rect 66418 19482 68442 19542
rect 68502 19482 68508 19542
rect 64136 7350 64196 7356
rect 65048 7350 65108 7356
rect 63266 7306 63326 7312
rect 64928 7306 64988 7312
rect 63326 7246 64928 7306
rect 63266 7240 63326 7246
rect 64928 7240 64988 7246
rect 62352 7198 62412 7204
rect 64030 7198 64090 7204
rect 64248 7198 64308 7204
rect 62341 7138 62350 7198
rect 62412 7138 64030 7198
rect 64090 7138 64248 7198
rect 62352 7132 62412 7138
rect 64030 7132 64090 7138
rect 64248 7132 64308 7138
rect 62482 7090 62542 7096
rect 63812 7090 63872 7096
rect 64466 7090 64526 7096
rect 62542 7030 63812 7090
rect 63872 7030 64466 7090
rect 62482 7024 62542 7030
rect 63812 7024 63872 7030
rect 64466 7024 64526 7030
rect 50459 7003 51160 7004
rect 50012 6944 51160 7003
rect 50012 6943 50563 6944
rect 49952 6937 50012 6943
rect 19628 6700 19688 6706
rect 23696 6700 23756 6706
rect 25730 6700 25790 6706
rect 15034 6694 15094 6700
rect 16042 6694 16102 6700
rect 17056 6694 17116 6700
rect 18094 6694 18154 6700
rect 19112 6694 19172 6700
rect 15094 6634 16042 6694
rect 16102 6634 17056 6694
rect 17116 6634 18094 6694
rect 18154 6634 19112 6694
rect 19688 6640 21664 6700
rect 21724 6640 23696 6700
rect 23756 6640 25730 6700
rect 19628 6634 19688 6640
rect 23696 6634 23756 6640
rect 25730 6634 25790 6640
rect 26752 6702 26812 6708
rect 27106 6702 27166 6708
rect 26812 6642 27106 6702
rect 26752 6636 26812 6642
rect 27106 6636 27166 6642
rect 30824 6702 30884 6708
rect 34108 6702 34168 6708
rect 30884 6642 34108 6702
rect 30824 6636 30884 6642
rect 34108 6636 34168 6642
rect 15034 6628 15094 6634
rect 16042 6628 16102 6634
rect 17056 6628 17116 6634
rect 18094 6628 18154 6634
rect 19112 6628 19172 6634
rect 13180 6590 13240 6596
rect 14536 6590 14596 6596
rect 22680 6590 22740 6596
rect 24716 6590 24776 6596
rect 26748 6590 26808 6596
rect 13240 6530 14536 6590
rect 14596 6530 22680 6590
rect 22740 6530 24716 6590
rect 24776 6530 26748 6590
rect 13180 6524 13240 6530
rect 14536 6524 14596 6530
rect 22680 6524 22740 6530
rect 24716 6524 24776 6530
rect 26748 6524 26808 6530
rect 26258 6492 26318 6498
rect 27296 6492 27356 6498
rect 28272 6492 28332 6498
rect 29288 6492 29348 6498
rect 31314 6492 31374 6498
rect 32344 6492 32404 6498
rect 10636 6410 12596 6470
rect 15552 6478 15612 6484
rect 17590 6478 17650 6484
rect 21662 6478 21722 6484
rect 15612 6418 17590 6478
rect 17650 6418 21662 6478
rect 26318 6432 27296 6492
rect 27356 6432 28272 6492
rect 28332 6432 29288 6492
rect 29348 6432 31314 6492
rect 31374 6432 32344 6492
rect 49948 6442 49954 6502
rect 50014 6442 50613 6502
rect 26258 6426 26318 6432
rect 27296 6426 27356 6432
rect 28272 6426 28332 6432
rect 29288 6426 29348 6432
rect 31314 6426 31374 6432
rect 32344 6426 32404 6432
rect 15552 6412 15612 6418
rect 17590 6412 17650 6418
rect 21662 6412 21722 6418
rect 10576 6404 10636 6410
rect 10358 6380 10418 6386
rect 9982 6320 10358 6380
rect 14532 6380 14592 6386
rect 16570 6380 16630 6386
rect 18610 6380 18670 6386
rect 20646 6380 20706 6386
rect 26750 6380 26810 6386
rect 27100 6380 27106 6384
rect 13286 6344 13346 6350
rect 9922 6314 9982 6320
rect 10358 6314 10418 6320
rect 11164 6284 11170 6344
rect 11230 6284 13286 6344
rect 14592 6320 16570 6380
rect 16630 6320 18610 6380
rect 18670 6320 20646 6380
rect 20706 6324 27106 6380
rect 27166 6380 27172 6384
rect 28786 6380 28846 6386
rect 30822 6380 30882 6386
rect 32858 6380 32918 6386
rect 27166 6324 28786 6380
rect 20706 6320 28786 6324
rect 28846 6320 30822 6380
rect 30882 6320 32858 6380
rect 14532 6314 14592 6320
rect 16570 6314 16630 6320
rect 18610 6314 18670 6320
rect 20646 6314 20706 6320
rect 26750 6314 26810 6320
rect 28786 6314 28846 6320
rect 30822 6314 30882 6320
rect 32858 6314 32918 6320
rect 13286 6278 13346 6284
rect 9158 6270 9218 6276
rect 9378 6270 9438 6276
rect 10032 6270 10092 6276
rect 10248 6270 10308 6276
rect 9218 6210 9378 6270
rect 9438 6210 10032 6270
rect 10092 6210 10248 6270
rect 9158 6204 9218 6210
rect 9378 6204 9438 6210
rect 10032 6204 10092 6210
rect 10248 6204 10308 6210
rect 45907 6098 45916 6198
rect 46016 6176 48434 6198
rect 46016 6116 48364 6176
rect 48424 6116 48434 6176
rect 46016 6098 48434 6116
rect 8482 5766 8542 5772
rect 8940 5766 9000 5772
rect 9596 5766 9656 5772
rect 8542 5706 8940 5766
rect 9000 5706 9596 5766
rect 8482 5700 8542 5706
rect 8940 5700 9000 5706
rect 9596 5700 9656 5706
rect 10140 5766 10200 5772
rect 10928 5766 10988 5772
rect 10200 5706 10928 5766
rect 49306 5736 49366 5742
rect 49824 5736 49884 5742
rect 10140 5700 10200 5706
rect 10928 5700 10988 5706
rect 49297 5676 49306 5736
rect 49366 5676 49824 5736
rect 49306 5670 49366 5676
rect 49824 5670 49884 5676
rect 50553 5664 50613 6442
rect 8352 5644 8412 5650
rect 9158 5644 9218 5650
rect 9376 5644 9436 5650
rect 8412 5584 9158 5644
rect 9218 5584 9376 5644
rect 8352 5578 8412 5584
rect 9158 5578 9218 5584
rect 9376 5578 9436 5584
rect 9812 5646 9872 5652
rect 10468 5646 10528 5652
rect 9872 5586 10468 5646
rect 50553 5604 50627 5664
rect 50687 5604 50693 5664
rect 50939 5626 50945 5686
rect 51005 5626 51011 5686
rect 49048 5587 49108 5593
rect 49564 5587 49624 5593
rect 9812 5580 9872 5586
rect 10468 5580 10528 5586
rect 49037 5527 49048 5587
rect 49108 5527 49564 5587
rect 49624 5527 49940 5587
rect 50000 5527 50082 5587
rect 50142 5527 50148 5587
rect 8832 5520 8892 5526
rect 9702 5520 9762 5526
rect 10574 5520 10634 5526
rect 49048 5521 49108 5527
rect 49564 5521 49624 5527
rect 8892 5460 9702 5520
rect 9762 5460 10574 5520
rect 21658 5476 21718 5482
rect 23700 5476 23760 5482
rect 25732 5476 25792 5482
rect 27772 5476 27832 5482
rect 34228 5476 34288 5482
rect 8832 5454 8892 5460
rect 9702 5454 9762 5460
rect 10574 5454 10634 5460
rect 15552 5456 15612 5462
rect 17588 5456 17648 5462
rect 19626 5456 19686 5462
rect 9270 5394 9330 5400
rect 11048 5394 11108 5400
rect 9330 5334 11048 5394
rect 15612 5396 17588 5456
rect 17648 5396 19626 5456
rect 21482 5416 21488 5476
rect 21548 5416 21658 5476
rect 21718 5416 23700 5476
rect 23760 5416 25732 5476
rect 25792 5416 27772 5476
rect 27832 5416 34228 5476
rect 21658 5410 21718 5416
rect 23700 5410 23760 5416
rect 25732 5410 25792 5416
rect 27772 5410 27832 5416
rect 34228 5410 34288 5416
rect 15552 5390 15612 5396
rect 17588 5390 17648 5396
rect 19626 5390 19686 5396
rect 26750 5378 26810 5384
rect 32856 5378 32916 5384
rect 34108 5378 34168 5384
rect 9270 5328 9330 5334
rect 11048 5328 11108 5334
rect 13398 5358 13458 5364
rect 16570 5358 16630 5364
rect 13458 5298 16570 5358
rect 13398 5292 13458 5298
rect 16570 5292 16630 5298
rect 18094 5358 18154 5364
rect 21142 5358 21202 5364
rect 18154 5298 19116 5358
rect 19176 5298 20138 5358
rect 20198 5298 21142 5358
rect 26810 5318 32856 5378
rect 32916 5318 34108 5378
rect 26750 5312 26810 5318
rect 32856 5312 32916 5318
rect 34108 5312 34168 5318
rect 18094 5292 18154 5298
rect 21142 5292 21202 5298
rect 9604 5280 9656 5286
rect 13186 5278 13192 5280
rect 9656 5230 13192 5278
rect 13186 5228 13192 5230
rect 13244 5228 13250 5280
rect 21664 5268 21724 5274
rect 23692 5268 23752 5274
rect 25736 5268 25796 5274
rect 27764 5268 27824 5274
rect 29802 5268 29862 5274
rect 31842 5268 31902 5274
rect 15556 5262 15616 5268
rect 17592 5262 17652 5268
rect 19620 5262 19680 5268
rect 21488 5262 21548 5268
rect 9604 5222 9656 5228
rect 8280 5204 8340 5210
rect 8271 5144 8280 5204
rect 8340 5144 8349 5204
rect 15616 5202 17592 5262
rect 17652 5202 19620 5262
rect 19680 5202 21488 5262
rect 21724 5208 23692 5268
rect 23752 5208 25736 5268
rect 25796 5208 27764 5268
rect 27824 5208 29802 5268
rect 29862 5208 31842 5268
rect 21664 5202 21724 5208
rect 23692 5202 23752 5208
rect 25736 5202 25796 5208
rect 27764 5202 27824 5208
rect 29802 5202 29862 5208
rect 31842 5202 31902 5208
rect 32360 5272 32420 5278
rect 34478 5272 34538 5278
rect 32420 5212 34478 5272
rect 32360 5206 32420 5212
rect 34478 5206 34538 5212
rect 15556 5196 15616 5202
rect 17592 5196 17652 5202
rect 19620 5196 19680 5202
rect 21488 5196 21548 5202
rect 8280 5138 8340 5144
rect 14538 5142 14598 5148
rect 18606 5142 18666 5148
rect 20640 5142 20700 5148
rect 28790 5142 28850 5148
rect 30820 5142 30880 5148
rect 32858 5144 32918 5150
rect 34350 5144 34410 5150
rect 14598 5082 18606 5142
rect 18666 5082 20640 5142
rect 20700 5082 28790 5142
rect 28850 5082 30820 5142
rect 31340 5084 31346 5144
rect 31406 5084 32858 5144
rect 32918 5084 34350 5144
rect 14538 5076 14598 5082
rect 18606 5076 18666 5082
rect 20640 5076 20700 5082
rect 28790 5076 28850 5082
rect 30820 5076 30880 5082
rect 32858 5078 32918 5084
rect 34350 5078 34410 5084
rect 10018 5060 10078 5066
rect 11212 5060 11272 5066
rect 11902 5060 11962 5066
rect 8822 5000 8828 5060
rect 8888 5000 10018 5060
rect 10078 5000 11212 5060
rect 11272 5000 11902 5060
rect 10018 4994 10078 5000
rect 11212 4994 11272 5000
rect 11902 4994 11962 5000
rect 49952 5039 50012 5045
rect 50945 5040 51005 5626
rect 50459 5039 51005 5040
rect 50012 4980 51005 5039
rect 50012 4979 50563 4980
rect 49952 4973 50012 4979
rect 8280 4960 8340 4966
rect 9272 4960 9332 4966
rect 9570 4960 9630 4966
rect 10466 4960 10526 4966
rect 10762 4960 10822 4966
rect 8340 4900 9272 4960
rect 9332 4900 9570 4960
rect 9630 4900 10466 4960
rect 10526 4900 10762 4960
rect 8280 4894 8340 4900
rect 9272 4894 9332 4900
rect 9570 4894 9630 4900
rect 10466 4894 10526 4900
rect 10762 4894 10822 4900
rect 49948 4442 49954 4502
rect 50014 4442 50613 4502
rect 13286 4226 13346 4232
rect 22674 4226 22734 4232
rect 24716 4226 24776 4232
rect 26752 4226 26812 4232
rect 13346 4166 22674 4226
rect 22734 4166 24716 4226
rect 24776 4166 26752 4226
rect 13286 4160 13346 4166
rect 22674 4160 22734 4166
rect 24716 4160 24776 4166
rect 26752 4160 26812 4166
rect 29806 4226 29866 4232
rect 31838 4226 31898 4232
rect 33984 4226 34044 4232
rect 29866 4166 31838 4226
rect 31898 4166 33984 4226
rect 29806 4160 29866 4166
rect 31838 4160 31898 4166
rect 33984 4160 34044 4166
rect 17090 4112 17150 4118
rect 22170 4112 22230 4118
rect 13180 4100 13240 4106
rect 16570 4100 16630 4106
rect 9121 4057 9179 4063
rect 9725 4057 9783 4063
rect 10316 4057 10374 4063
rect 9179 3999 9725 4057
rect 9783 3999 10316 4057
rect 10374 3999 10913 4057
rect 10971 3999 11509 4057
rect 11567 3999 11573 4057
rect 13240 4040 16570 4100
rect 17150 4052 22170 4112
rect 17090 4046 17150 4052
rect 22170 4046 22230 4052
rect 27258 4116 27318 4122
rect 32358 4116 32418 4122
rect 27318 4056 32358 4116
rect 38910 4099 39020 4104
rect 27258 4050 27318 4056
rect 32358 4050 32418 4056
rect 13180 4034 13240 4040
rect 16570 4034 16630 4040
rect 38906 3999 38915 4099
rect 39015 3999 39024 4099
rect 43082 4097 43192 4102
rect 9121 3993 9179 3999
rect 9725 3993 9783 3999
rect 10316 3993 10374 3999
rect 15552 3990 15612 3996
rect 17588 3990 17648 3996
rect 18608 3990 18668 3996
rect 19624 3990 19684 3996
rect 20644 3990 20704 3996
rect 21662 3990 21722 3996
rect 23692 3990 23752 3996
rect 25730 3990 25790 3996
rect 27766 3990 27826 3996
rect 28788 3990 28848 3996
rect 29808 3990 29868 3996
rect 30822 3990 30882 3996
rect 31844 3990 31904 3996
rect 8408 3926 8468 3932
rect 9418 3926 9478 3932
rect 10016 3926 10076 3932
rect 10610 3926 10670 3932
rect 11208 3926 11268 3932
rect 8468 3866 8824 3926
rect 8884 3866 9418 3926
rect 9478 3866 10016 3926
rect 10076 3866 10610 3926
rect 10670 3866 11208 3926
rect 15612 3930 17588 3990
rect 17648 3930 18608 3990
rect 18668 3930 19624 3990
rect 19684 3930 20644 3990
rect 20704 3930 21662 3990
rect 21722 3930 23692 3990
rect 23752 3930 25730 3990
rect 25790 3930 27766 3990
rect 27826 3930 28788 3990
rect 28848 3930 29808 3990
rect 29868 3930 30822 3990
rect 30882 3930 31844 3990
rect 15552 3924 15612 3930
rect 17588 3924 17648 3930
rect 18608 3924 18668 3930
rect 19624 3924 19684 3930
rect 20644 3924 20704 3930
rect 21662 3924 21722 3930
rect 23692 3924 23752 3930
rect 25730 3924 25790 3930
rect 27766 3924 27826 3930
rect 28788 3924 28848 3930
rect 29808 3924 29868 3930
rect 30822 3924 30882 3930
rect 31844 3924 31904 3930
rect 38910 3971 39020 3999
rect 43078 3997 43087 4097
rect 43187 3997 43196 4097
rect 8408 3860 8468 3866
rect 9418 3860 9478 3866
rect 10016 3860 10076 3866
rect 10610 3860 10670 3866
rect 11208 3860 11268 3866
rect 17206 3896 17266 3902
rect 18090 3896 18150 3902
rect 19112 3896 19172 3902
rect 21154 3896 21214 3902
rect 17266 3836 18090 3896
rect 18150 3836 19112 3896
rect 19172 3836 21154 3896
rect 17206 3830 17266 3836
rect 18090 3830 18150 3836
rect 19112 3830 19172 3836
rect 21154 3830 21214 3836
rect 28276 3896 28336 3902
rect 29296 3896 29356 3902
rect 30310 3896 30370 3902
rect 31346 3896 31406 3902
rect 28336 3836 29296 3896
rect 29356 3836 30310 3896
rect 30370 3836 31346 3896
rect 38910 3861 40895 3971
rect 28276 3830 28336 3836
rect 29296 3830 29356 3836
rect 30310 3830 30370 3836
rect 31346 3830 31406 3836
rect 8976 3818 9036 3824
rect 9274 3818 9334 3824
rect 9574 3818 9634 3824
rect 9868 3818 9928 3824
rect 10164 3818 10224 3824
rect 10464 3818 10524 3824
rect 10766 3818 10826 3824
rect 11056 3818 11116 3824
rect 11360 3818 11420 3824
rect 9036 3758 9274 3818
rect 9334 3758 9574 3818
rect 9634 3758 9868 3818
rect 9928 3758 10164 3818
rect 10224 3758 10464 3818
rect 10524 3758 10766 3818
rect 10826 3758 11056 3818
rect 11116 3758 11360 3818
rect 11420 3758 12026 3818
rect 12086 3758 12092 3818
rect 40785 3799 40895 3861
rect 43082 3957 43192 3997
rect 43082 3847 45171 3957
rect 8976 3752 9036 3758
rect 9274 3752 9334 3758
rect 9574 3752 9634 3758
rect 9868 3752 9928 3758
rect 10164 3752 10224 3758
rect 10464 3752 10524 3758
rect 10766 3752 10826 3758
rect 11056 3752 11116 3758
rect 11360 3752 11420 3758
rect 40785 3680 40895 3689
rect 45061 3787 45171 3847
rect 49306 3736 49366 3742
rect 49824 3736 49884 3742
rect 45061 3668 45171 3677
rect 49293 3676 49302 3736
rect 49366 3676 49824 3736
rect 49306 3670 49366 3676
rect 49824 3670 49884 3676
rect 50553 3664 50613 4442
rect 50945 3686 51005 4980
rect 50553 3604 50627 3664
rect 50687 3604 50693 3664
rect 50939 3626 50945 3686
rect 51005 3626 51011 3686
rect 49048 3587 49108 3593
rect 49564 3587 49624 3593
rect 49037 3527 49048 3587
rect 49108 3527 49564 3587
rect 49624 3527 50082 3587
rect 50142 3527 50151 3587
rect 49048 3521 49108 3527
rect 49564 3521 49624 3527
rect 49952 3039 50012 3045
rect 50945 3040 51005 3626
rect 50459 3039 51005 3040
rect 12926 2996 12986 3002
rect 13518 2996 13578 3002
rect 14032 2996 14092 3002
rect 14530 2996 14590 3002
rect 16572 2996 16632 3002
rect 18604 2996 18664 3002
rect 20636 2996 20696 3002
rect 24894 2996 24900 2998
rect 12494 2994 12926 2996
rect 12350 2936 12926 2994
rect 12986 2936 13518 2996
rect 13578 2936 14032 2996
rect 14092 2936 14530 2996
rect 14590 2936 16572 2996
rect 16632 2936 18604 2996
rect 18664 2936 20636 2996
rect 20696 2936 22540 2996
rect 22600 2938 24900 2996
rect 24960 2996 24966 2998
rect 26750 2996 26810 3002
rect 28784 2996 28844 3002
rect 30818 2996 30878 3002
rect 32860 2996 32920 3002
rect 33372 2996 33432 3002
rect 33878 2996 33938 3002
rect 24960 2938 26750 2996
rect 22600 2936 26750 2938
rect 26810 2936 28784 2996
rect 28844 2936 30818 2996
rect 30878 2936 32860 2996
rect 32920 2936 33372 2996
rect 33432 2936 33878 2996
rect 50012 2980 51005 3039
rect 50012 2979 50563 2980
rect 49952 2973 50012 2979
rect 12350 2934 12586 2936
rect 2756 2864 4582 2924
rect 4642 2864 6452 2924
rect 6512 2864 7914 2924
rect 8280 2920 8340 2926
rect 8974 2920 9034 2926
rect 9870 2920 9930 2926
rect 10164 2920 10224 2926
rect 11058 2920 11118 2926
rect 11360 2920 11420 2926
rect 2696 2858 2756 2864
rect 4582 2858 4642 2864
rect 6452 2858 6512 2864
rect 8340 2860 8974 2920
rect 9034 2860 9870 2920
rect 9930 2860 10164 2920
rect 10224 2860 11058 2920
rect 11118 2860 11360 2920
rect 8280 2854 8340 2860
rect 8974 2854 9034 2860
rect 9870 2854 9930 2860
rect 10164 2854 10224 2860
rect 11058 2854 11118 2860
rect 11360 2854 11420 2860
rect 2548 2816 2608 2822
rect 4584 2816 4644 2822
rect 6620 2816 6680 2822
rect 2608 2756 4584 2816
rect 4644 2756 6620 2816
rect 2548 2750 2608 2756
rect 4584 2750 4644 2756
rect 6620 2750 6680 2756
rect 9420 2812 9480 2818
rect 10614 2812 10674 2818
rect 9480 2752 10614 2812
rect 10674 2752 11902 2812
rect 11962 2752 11968 2812
rect 9420 2746 9480 2752
rect 10614 2746 10674 2752
rect 3566 2704 3626 2710
rect 3626 2644 5604 2704
rect 5664 2644 5670 2704
rect 3566 2638 3626 2644
rect 9122 1828 9182 1834
rect 9716 1828 9776 1834
rect 10316 1828 10376 1834
rect 10910 1828 10970 1834
rect 11504 1828 11564 1834
rect 12350 1828 12410 2934
rect 12926 2930 12986 2936
rect 13518 2930 13578 2936
rect 14032 2930 14092 2936
rect 14530 2930 14590 2936
rect 16572 2930 16632 2936
rect 18604 2930 18664 2936
rect 20636 2930 20696 2936
rect 26750 2930 26810 2936
rect 28784 2930 28844 2936
rect 30818 2930 30878 2936
rect 32860 2930 32920 2936
rect 33372 2930 33432 2936
rect 33878 2930 33938 2936
rect 17080 2884 17140 2890
rect 18092 2884 18152 2890
rect 19106 2884 19166 2890
rect 22018 2884 22078 2890
rect 17140 2824 18092 2884
rect 18152 2824 19106 2884
rect 19166 2824 22018 2884
rect 17080 2818 17140 2824
rect 18092 2818 18152 2824
rect 19106 2818 19166 2824
rect 22018 2818 22078 2824
rect 22678 2886 22738 2892
rect 13060 2778 13120 2784
rect 15046 2778 15106 2784
rect 16068 2778 16128 2784
rect 18606 2778 18666 2784
rect 19118 2778 19178 2784
rect 20136 2778 20196 2784
rect 20642 2778 20702 2784
rect 21148 2778 21208 2784
rect 22160 2778 22220 2784
rect 22678 2778 22738 2826
rect 23306 2882 23366 2888
rect 24352 2882 24412 2888
rect 28280 2882 28340 2888
rect 29298 2882 29358 2888
rect 23366 2822 24352 2882
rect 24412 2822 28280 2882
rect 28340 2822 29298 2882
rect 29358 2822 30308 2882
rect 30368 2822 30374 2882
rect 23306 2816 23366 2822
rect 24352 2816 24412 2822
rect 28280 2816 28340 2822
rect 29298 2816 29358 2822
rect 23180 2778 23240 2784
rect 24202 2778 24262 2784
rect 24714 2778 24774 2784
rect 25220 2778 25280 2784
rect 26238 2778 26298 2784
rect 26750 2778 26810 2784
rect 27258 2778 27318 2784
rect 31330 2778 31390 2784
rect 32332 2778 32392 2784
rect 13120 2718 15046 2778
rect 15106 2718 16068 2778
rect 16128 2718 18606 2778
rect 18666 2718 19118 2778
rect 19178 2718 20136 2778
rect 20196 2718 20642 2778
rect 20702 2718 21148 2778
rect 21208 2718 22160 2778
rect 22220 2718 23180 2778
rect 23240 2718 24202 2778
rect 24262 2718 24714 2778
rect 24774 2718 25220 2778
rect 25280 2718 26238 2778
rect 26298 2718 26750 2778
rect 26810 2718 27258 2778
rect 27318 2718 31330 2778
rect 31390 2718 32332 2778
rect 13060 2712 13120 2718
rect 15046 2712 15106 2718
rect 16068 2712 16128 2718
rect 18606 2712 18666 2718
rect 19118 2712 19178 2718
rect 20136 2712 20196 2718
rect 20642 2712 20702 2718
rect 21148 2712 21208 2718
rect 22160 2712 22220 2718
rect 23180 2712 23240 2718
rect 24202 2712 24262 2718
rect 24714 2712 24774 2718
rect 25220 2712 25280 2718
rect 26238 2712 26298 2718
rect 26750 2712 26810 2718
rect 27258 2712 27318 2718
rect 31330 2712 31390 2718
rect 32332 2712 32392 2718
rect 12654 2674 12714 2680
rect 17082 2674 17142 2680
rect 17586 2674 17646 2680
rect 18102 2674 18162 2680
rect 19624 2674 19684 2680
rect 21662 2674 21722 2680
rect 23698 2674 23758 2680
rect 25734 2674 25794 2680
rect 27766 2674 27826 2680
rect 28288 2674 28348 2680
rect 28788 2674 28848 2680
rect 29296 2674 29356 2680
rect 29804 2674 29864 2680
rect 30154 2674 30214 2680
rect 34756 2674 34816 2680
rect 12714 2614 17082 2674
rect 17142 2614 17586 2674
rect 17646 2614 18102 2674
rect 18162 2614 19624 2674
rect 19684 2614 21662 2674
rect 21722 2614 23698 2674
rect 23758 2614 25734 2674
rect 25794 2614 27766 2674
rect 27826 2614 28288 2674
rect 28348 2614 28788 2674
rect 28848 2614 29296 2674
rect 29356 2614 29804 2674
rect 29864 2614 30154 2674
rect 30214 2614 34756 2674
rect 12654 2608 12714 2614
rect 17082 2608 17142 2614
rect 17586 2608 17646 2614
rect 18102 2608 18162 2614
rect 19624 2608 19684 2614
rect 21662 2608 21722 2614
rect 23698 2608 23758 2614
rect 25734 2608 25794 2614
rect 27766 2608 27826 2614
rect 28288 2608 28348 2614
rect 28788 2608 28848 2614
rect 29296 2608 29356 2614
rect 29804 2608 29864 2614
rect 30154 2608 30214 2614
rect 34756 2608 34816 2614
rect 49948 2352 49954 2412
rect 50014 2352 50613 2412
rect 3568 1822 3628 1828
rect 3628 1762 5598 1822
rect 5658 1762 5664 1822
rect 9182 1768 9716 1828
rect 9776 1768 10316 1828
rect 10376 1768 10910 1828
rect 10970 1768 11504 1828
rect 11564 1768 12410 1828
rect 9122 1762 9182 1768
rect 9716 1762 9776 1768
rect 10316 1762 10376 1768
rect 10910 1762 10970 1768
rect 11504 1762 11564 1768
rect 3568 1756 3628 1762
rect 22680 1742 22740 1748
rect 24716 1742 24776 1748
rect 9416 1734 9476 1740
rect 10014 1734 10074 1740
rect 10612 1734 10672 1740
rect 11212 1734 11272 1740
rect 2550 1720 2610 1726
rect 6618 1720 6678 1726
rect 7748 1720 7808 1726
rect 2610 1660 6618 1720
rect 6678 1660 7748 1720
rect 8518 1674 8524 1734
rect 8584 1674 9416 1734
rect 9476 1674 10014 1734
rect 10074 1674 10612 1734
rect 10672 1674 11212 1734
rect 22740 1682 24716 1742
rect 22680 1676 22740 1682
rect 24716 1676 24776 1682
rect 9416 1668 9476 1674
rect 10014 1668 10074 1674
rect 10612 1668 10672 1674
rect 11212 1668 11272 1674
rect 2550 1654 2610 1660
rect 6618 1654 6678 1660
rect 7748 1654 7808 1660
rect 8972 1626 9032 1632
rect 9270 1626 9330 1632
rect 9566 1626 9626 1632
rect 9870 1626 9930 1632
rect 10166 1626 10226 1632
rect 10464 1626 10524 1632
rect 10760 1626 10820 1632
rect 11056 1626 11116 1632
rect 11360 1626 11420 1632
rect 12026 1626 12086 1632
rect 1412 1614 1472 1620
rect 4584 1614 4644 1620
rect 1472 1554 4584 1614
rect 1412 1548 1472 1554
rect 4584 1548 4644 1554
rect 8042 1566 8972 1626
rect 9032 1566 9270 1626
rect 9330 1566 9566 1626
rect 9626 1566 9870 1626
rect 9930 1566 10166 1626
rect 10226 1566 10464 1626
rect 10524 1566 10760 1626
rect 10820 1566 11056 1626
rect 11116 1566 11360 1626
rect 11420 1566 12026 1626
rect 46079 1610 46088 1670
rect 46148 1610 46157 1670
rect 49306 1646 49366 1652
rect 49824 1646 49884 1652
rect 3054 670 3114 676
rect 4080 670 4140 676
rect 5104 670 5164 676
rect 3114 610 4080 670
rect 4140 610 5104 670
rect 5164 610 6004 670
rect 6064 610 6070 670
rect 3054 604 3114 610
rect 4080 604 4140 610
rect 5104 604 5164 610
rect 8042 582 8102 1566
rect 8972 1560 9032 1566
rect 9270 1560 9330 1566
rect 9566 1560 9626 1566
rect 9870 1560 9930 1566
rect 10166 1560 10226 1566
rect 10464 1560 10524 1566
rect 10760 1560 10820 1566
rect 11056 1560 11116 1566
rect 11360 1560 11420 1566
rect 12026 1560 12086 1566
rect 14530 1542 14590 1548
rect 16568 1542 16628 1548
rect 18606 1542 18666 1548
rect 20638 1542 20698 1548
rect 22676 1542 22736 1548
rect 24710 1542 24770 1548
rect 26750 1542 26810 1548
rect 28784 1542 28844 1548
rect 30818 1542 30878 1548
rect 32856 1542 32916 1548
rect 34598 1542 34658 1548
rect 14590 1482 16568 1542
rect 16628 1482 18606 1542
rect 18666 1482 20638 1542
rect 20698 1482 22676 1542
rect 22736 1482 24710 1542
rect 24770 1482 26750 1542
rect 26810 1482 28784 1542
rect 28844 1482 30818 1542
rect 30878 1482 32856 1542
rect 32916 1482 34598 1542
rect 14530 1476 14590 1482
rect 16568 1476 16628 1482
rect 18606 1476 18666 1482
rect 20638 1476 20698 1482
rect 22676 1476 22736 1482
rect 24710 1476 24770 1482
rect 26750 1476 26810 1482
rect 28784 1476 28844 1482
rect 30818 1476 30878 1482
rect 32856 1476 32916 1482
rect 34598 1476 34658 1482
rect 46088 1497 46148 1610
rect 49366 1586 49824 1646
rect 49888 1586 49897 1646
rect 49306 1580 49366 1586
rect 49824 1580 49884 1586
rect 50553 1574 50613 2352
rect 51100 1596 51160 6944
rect 66418 6816 66478 19482
rect 68782 19442 68842 19448
rect 69652 19442 69712 19448
rect 70526 19442 70586 19448
rect 70882 19442 70942 19448
rect 64922 6756 64928 6816
rect 64988 6756 66478 6816
rect 66536 19382 68782 19442
rect 68842 19382 69652 19442
rect 69712 19382 70526 19442
rect 70586 19382 70882 19442
rect 62940 6590 63000 6596
rect 63596 6590 63656 6596
rect 64466 6590 64526 6596
rect 65170 6590 65230 6596
rect 63000 6530 63596 6590
rect 63656 6530 64466 6590
rect 64526 6530 65170 6590
rect 62940 6524 63000 6530
rect 63596 6524 63656 6530
rect 64466 6524 64526 6530
rect 65170 6524 65230 6530
rect 63048 6490 63108 6496
rect 63486 6490 63546 6496
rect 61854 6430 63048 6490
rect 63108 6430 63486 6490
rect 63546 6430 63982 6490
rect 57564 4940 57624 4946
rect 59604 4940 59664 4946
rect 57624 4880 59604 4940
rect 57564 4874 57624 4880
rect 59604 4874 59664 4880
rect 55412 4036 55472 4042
rect 56550 4036 56610 4042
rect 60624 4036 60684 4042
rect 55472 3976 56550 4036
rect 56610 3976 60624 4036
rect 55412 3970 55472 3976
rect 56550 3970 56610 3976
rect 60624 3970 60684 3976
rect 57564 3940 57624 3946
rect 59604 3940 59664 3946
rect 57624 3880 59604 3940
rect 57564 3874 57624 3880
rect 59604 3874 59664 3880
rect 58586 3824 58646 3830
rect 61748 3824 61808 3830
rect 58646 3764 61748 3824
rect 58586 3758 58646 3764
rect 61748 3758 61808 3764
rect 56696 2924 56756 2930
rect 58582 2924 58642 2930
rect 60452 2924 60512 2930
rect 61854 2924 61914 6430
rect 63048 6424 63108 6430
rect 63486 6424 63546 6430
rect 61974 6380 62034 6386
rect 63050 6380 63110 6386
rect 63484 6380 63544 6386
rect 63812 6380 63872 6386
rect 62034 6320 63050 6380
rect 63110 6320 63484 6380
rect 63544 6320 63812 6380
rect 61974 6314 62034 6320
rect 63050 6314 63110 6320
rect 63484 6314 63544 6320
rect 63812 6314 63872 6320
rect 63922 6380 63982 6430
rect 64576 6470 64636 6476
rect 66536 6470 66596 19382
rect 68782 19376 68842 19382
rect 69652 19376 69712 19382
rect 70526 19376 70586 19382
rect 70882 19376 70942 19382
rect 68998 19344 69058 19350
rect 69434 19344 69494 19350
rect 69872 19344 69932 19350
rect 70306 19344 70366 19350
rect 69058 19284 69434 19344
rect 69494 19284 69872 19344
rect 69932 19284 70306 19344
rect 68998 19278 69058 19284
rect 69434 19278 69494 19284
rect 69872 19278 69932 19284
rect 70306 19278 70366 19284
rect 68442 19226 68502 19232
rect 69108 19226 69168 19232
rect 69216 19226 69276 19232
rect 69324 19226 69384 19232
rect 69970 19226 70030 19232
rect 70088 19226 70148 19232
rect 68502 19166 69108 19226
rect 69168 19166 69216 19226
rect 69276 19166 69324 19226
rect 69384 19166 69970 19226
rect 70030 19166 70088 19226
rect 70197 19224 70255 19230
rect 70148 19166 70197 19224
rect 68442 19160 68502 19166
rect 69108 19160 69168 19166
rect 69216 19160 69276 19166
rect 69324 19160 69384 19166
rect 69970 19160 70030 19166
rect 70088 19160 70148 19166
rect 70197 19160 70255 19166
rect 67268 18823 67277 18913
rect 67367 18823 67376 18913
rect 67060 18148 67120 18154
rect 66898 17982 66904 18042
rect 66964 17982 66970 18042
rect 66646 16327 66655 16417
rect 66745 16327 66754 16417
rect 66670 15064 66730 16327
rect 66904 15192 66964 17982
rect 66904 15126 66964 15132
rect 67060 15192 67120 18088
rect 67286 15184 67346 18823
rect 68782 18506 68842 18512
rect 68892 18506 68952 18512
rect 69546 18506 69606 18512
rect 69652 18506 69712 18512
rect 69762 18506 69822 18512
rect 70414 18506 70474 18512
rect 70526 18506 70586 18512
rect 70998 18506 71058 18512
rect 68842 18446 68892 18506
rect 68952 18446 69546 18506
rect 69606 18446 69652 18506
rect 69712 18446 69762 18506
rect 69822 18446 70414 18506
rect 70474 18446 70526 18506
rect 70586 18446 70998 18506
rect 68782 18440 68842 18446
rect 68892 18440 68952 18446
rect 69546 18440 69606 18446
rect 69652 18440 69712 18446
rect 69762 18440 69822 18446
rect 70414 18440 70474 18446
rect 70526 18440 70586 18446
rect 70998 18440 71058 18446
rect 67060 15126 67120 15132
rect 67280 15124 67286 15184
rect 67346 15124 67352 15184
rect 71864 15064 71924 19616
rect 73430 19610 73490 19616
rect 75466 19610 75526 19616
rect 78520 19678 78580 19684
rect 80556 19678 80616 19684
rect 78580 19618 80556 19678
rect 78520 19612 78580 19618
rect 80556 19612 80616 19618
rect 83610 19680 83670 19686
rect 85646 19680 85706 19686
rect 83670 19620 85646 19680
rect 83610 19614 83670 19620
rect 85646 19614 85706 19620
rect 75466 19568 75526 19574
rect 87796 19568 87856 19574
rect 75526 19508 87796 19568
rect 75466 19502 75526 19508
rect 87796 19502 87856 19508
rect 72262 19468 72322 19474
rect 72322 19408 84846 19468
rect 72262 19402 72322 19408
rect 76682 19372 76742 19378
rect 74444 19366 74504 19372
rect 76478 19366 76538 19372
rect 74504 19306 76478 19366
rect 76742 19312 78516 19372
rect 78576 19312 78582 19372
rect 79536 19368 79596 19374
rect 81570 19368 81630 19374
rect 76682 19306 76742 19312
rect 79596 19308 81570 19368
rect 74444 19300 74504 19306
rect 76478 19300 76538 19306
rect 79536 19302 79596 19308
rect 81570 19302 81630 19308
rect 81784 19364 81844 19370
rect 84632 19366 84692 19372
rect 84786 19366 84846 19408
rect 86666 19366 86726 19372
rect 81844 19304 84120 19364
rect 84180 19304 84186 19364
rect 84692 19306 86666 19366
rect 81784 19298 81844 19304
rect 84632 19300 84692 19306
rect 86666 19300 86726 19306
rect 71994 18418 72054 18424
rect 73426 18418 73486 18424
rect 75462 18418 75522 18424
rect 72054 18358 73426 18418
rect 73486 18358 75462 18418
rect 71994 18352 72054 18358
rect 73426 18352 73486 18358
rect 75462 18352 75522 18358
rect 83614 18418 83674 18424
rect 85650 18418 85710 18424
rect 83674 18358 85650 18418
rect 83614 18352 83674 18358
rect 72130 18288 72190 18294
rect 83744 18288 83804 18358
rect 85650 18352 85710 18358
rect 72190 18228 83804 18288
rect 72130 18222 72190 18228
rect 76484 18148 76544 18154
rect 88088 18148 88148 18154
rect 76544 18088 88088 18148
rect 76484 18082 76544 18088
rect 66670 15004 71924 15064
rect 66670 10080 66730 15004
rect 66800 14092 66860 14098
rect 67518 14092 67578 14098
rect 69554 14092 69614 14098
rect 71588 14092 71648 14098
rect 73628 14092 73688 14098
rect 75664 14092 75724 14098
rect 77698 14092 77758 14098
rect 79734 14092 79794 14098
rect 81770 14092 81830 14098
rect 83806 14092 83866 14098
rect 85844 14092 85904 14098
rect 87874 14092 87934 14098
rect 66860 14032 67518 14092
rect 67578 14032 69554 14092
rect 69614 14032 71588 14092
rect 71648 14032 73628 14092
rect 73688 14032 75664 14092
rect 75724 14032 77698 14092
rect 77758 14032 79734 14092
rect 79794 14032 81770 14092
rect 81830 14032 83806 14092
rect 83866 14032 85844 14092
rect 85904 14032 87874 14092
rect 66800 14026 66860 14032
rect 67518 14026 67578 14032
rect 69554 14026 69614 14032
rect 71588 14026 71648 14032
rect 73628 14026 73688 14032
rect 75664 14026 75724 14032
rect 77698 14026 77758 14032
rect 79734 14026 79794 14032
rect 81770 14026 81830 14032
rect 83806 14026 83866 14032
rect 85844 14026 85904 14032
rect 87874 14026 87934 14032
rect 68536 13994 68596 14000
rect 70574 13994 70634 14000
rect 72608 13994 72668 14000
rect 74642 13994 74702 14000
rect 76682 13994 76742 14000
rect 78716 13994 78776 14000
rect 80754 13994 80814 14000
rect 82786 13994 82846 14000
rect 84824 13994 84884 14000
rect 86862 13994 86922 14000
rect 87996 13994 88056 18088
rect 88088 18082 88148 18088
rect 88598 13994 88658 14000
rect 68596 13934 70574 13994
rect 70634 13934 72608 13994
rect 72668 13934 74642 13994
rect 74702 13934 76682 13994
rect 76742 13934 78716 13994
rect 78776 13934 80754 13994
rect 80814 13934 82786 13994
rect 82846 13934 84824 13994
rect 84884 13934 86862 13994
rect 86922 13934 88598 13994
rect 68536 13928 68596 13934
rect 70574 13928 70634 13934
rect 72608 13928 72668 13934
rect 74642 13928 74702 13934
rect 76682 13928 76742 13934
rect 78716 13928 78776 13934
rect 80754 13928 80814 13934
rect 82786 13928 82846 13934
rect 84824 13928 84884 13934
rect 86862 13928 86922 13934
rect 88598 13928 88658 13934
rect 76682 13782 76742 13788
rect 78714 13782 78774 13788
rect 76742 13722 78714 13782
rect 76682 13716 76742 13722
rect 78714 13716 78774 13722
rect 71222 12862 71282 12868
rect 71592 12862 71652 12868
rect 72094 12862 72154 12868
rect 72606 12862 72666 12868
rect 73134 12862 73194 12868
rect 73626 12862 73686 12868
rect 75658 12862 75718 12868
rect 77694 12862 77754 12868
rect 79730 12862 79790 12868
rect 81768 12862 81828 12868
rect 83806 12862 83866 12868
rect 84314 12862 84374 12868
rect 71282 12802 71592 12862
rect 71652 12802 72094 12862
rect 72154 12802 72606 12862
rect 72666 12802 73134 12862
rect 73194 12802 73626 12862
rect 73686 12802 75658 12862
rect 75718 12802 77694 12862
rect 77754 12802 79730 12862
rect 79790 12802 81768 12862
rect 81828 12802 83292 12862
rect 83352 12802 83806 12862
rect 83866 12802 84314 12862
rect 71222 12796 71282 12802
rect 71592 12796 71652 12802
rect 72094 12796 72154 12802
rect 72606 12796 72666 12802
rect 73134 12796 73194 12802
rect 73626 12796 73686 12802
rect 75658 12796 75718 12802
rect 77694 12796 77754 12802
rect 79730 12796 79790 12802
rect 81768 12796 81828 12802
rect 83806 12796 83866 12802
rect 84314 12796 84374 12802
rect 69046 12752 69106 12758
rect 70068 12752 70128 12758
rect 74140 12752 74200 12758
rect 74644 12752 74704 12758
rect 75160 12752 75220 12758
rect 76180 12752 76240 12758
rect 76682 12752 76742 12758
rect 77182 12752 77242 12758
rect 78208 12752 78268 12758
rect 78718 12752 78778 12758
rect 79226 12752 79286 12758
rect 80234 12752 80294 12758
rect 80756 12752 80816 12758
rect 81246 12752 81306 12758
rect 82278 12752 82338 12758
rect 82790 12752 82850 12758
rect 85334 12752 85394 12758
rect 86354 12752 86414 12758
rect 67056 12692 67062 12752
rect 67122 12692 69046 12752
rect 69106 12692 70068 12752
rect 70128 12692 74140 12752
rect 74200 12692 74644 12752
rect 74704 12692 75160 12752
rect 75220 12692 76180 12752
rect 76240 12692 76682 12752
rect 76742 12692 77182 12752
rect 77242 12692 78208 12752
rect 78268 12692 78718 12752
rect 78778 12692 79226 12752
rect 79286 12692 80234 12752
rect 80294 12692 80756 12752
rect 80816 12692 81246 12752
rect 81306 12692 82278 12752
rect 82338 12692 82790 12752
rect 82850 12692 85334 12752
rect 85394 12692 86354 12752
rect 69046 12686 69106 12692
rect 70068 12686 70128 12692
rect 74140 12686 74200 12692
rect 74644 12686 74704 12692
rect 75160 12686 75220 12692
rect 76180 12686 76240 12692
rect 76682 12686 76742 12692
rect 77182 12686 77242 12692
rect 78208 12686 78268 12692
rect 78718 12686 78778 12692
rect 79226 12686 79286 12692
rect 80234 12686 80294 12692
rect 80756 12686 80816 12692
rect 81246 12686 81306 12692
rect 82278 12686 82338 12692
rect 82790 12686 82850 12692
rect 85334 12686 85394 12692
rect 86354 12686 86414 12692
rect 72088 12648 72148 12654
rect 73108 12648 73168 12654
rect 77322 12648 77382 12654
rect 78330 12648 78390 12654
rect 79372 12648 79432 12654
rect 82264 12648 82324 12654
rect 83302 12648 83362 12654
rect 84302 12648 84362 12654
rect 71082 12588 71088 12648
rect 71148 12588 72088 12648
rect 72148 12588 73108 12648
rect 73168 12588 77322 12648
rect 77382 12588 78330 12648
rect 78390 12588 79372 12648
rect 79432 12588 82264 12648
rect 82324 12588 83302 12648
rect 83362 12588 84302 12648
rect 72088 12582 72148 12588
rect 73108 12582 73168 12588
rect 77322 12582 77382 12588
rect 78330 12582 78390 12588
rect 79372 12582 79432 12588
rect 82264 12582 82324 12588
rect 83302 12582 83362 12588
rect 84302 12582 84362 12588
rect 66926 12540 66986 12546
rect 67522 12540 67582 12546
rect 68020 12540 68080 12546
rect 68532 12540 68592 12546
rect 70574 12540 70634 12546
rect 72608 12540 72668 12546
rect 74642 12540 74702 12546
rect 80756 12540 80816 12546
rect 82788 12540 82848 12546
rect 84820 12540 84880 12546
rect 86862 12540 86922 12546
rect 87366 12540 87426 12546
rect 87876 12540 87936 12546
rect 66986 12480 67522 12540
rect 67582 12480 68020 12540
rect 68080 12480 68532 12540
rect 68592 12480 70574 12540
rect 70634 12480 72608 12540
rect 72668 12480 74642 12540
rect 74702 12480 76798 12540
rect 76858 12538 80756 12540
rect 76858 12480 78522 12538
rect 66926 12474 66986 12480
rect 67522 12474 67582 12480
rect 68020 12474 68080 12480
rect 68532 12474 68592 12480
rect 70574 12474 70634 12480
rect 72608 12474 72668 12480
rect 74642 12474 74702 12480
rect 78516 12478 78522 12480
rect 78582 12480 80756 12538
rect 80816 12480 82788 12540
rect 82848 12480 84820 12540
rect 84880 12480 86862 12540
rect 86922 12480 87366 12540
rect 87426 12480 87876 12540
rect 78582 12478 78588 12480
rect 80756 12474 80816 12480
rect 82788 12474 82848 12480
rect 84820 12474 84880 12480
rect 86862 12474 86922 12480
rect 87366 12474 87426 12480
rect 87876 12474 87936 12480
rect 70052 11650 70112 11656
rect 71072 11650 71132 11656
rect 72084 11650 72144 11656
rect 73110 11650 73170 11656
rect 82266 11650 82326 11656
rect 83302 11650 83362 11656
rect 84318 11650 84378 11656
rect 66800 11638 66860 11644
rect 69036 11638 69096 11644
rect 66860 11578 69036 11638
rect 70112 11590 71072 11650
rect 71132 11590 72084 11650
rect 72144 11590 73110 11650
rect 73170 11590 82266 11650
rect 82326 11590 83302 11650
rect 83362 11590 84318 11650
rect 70052 11584 70112 11590
rect 71072 11584 71132 11590
rect 72084 11584 72144 11590
rect 73110 11584 73170 11590
rect 82266 11584 82326 11590
rect 83302 11584 83362 11590
rect 84318 11584 84378 11590
rect 66800 11572 66860 11578
rect 69036 11572 69096 11578
rect 69548 11546 69608 11552
rect 70572 11546 70632 11552
rect 71584 11546 71644 11552
rect 72604 11546 72664 11552
rect 73626 11546 73686 11552
rect 75662 11546 75722 11552
rect 77700 11546 77760 11552
rect 79730 11546 79790 11552
rect 80750 11546 80810 11552
rect 81768 11546 81828 11552
rect 82788 11546 82848 11552
rect 83804 11546 83864 11552
rect 85840 11546 85900 11552
rect 69608 11486 70572 11546
rect 70632 11486 71584 11546
rect 71644 11486 72604 11546
rect 72664 11486 73626 11546
rect 73686 11486 75662 11546
rect 75722 11486 77700 11546
rect 77760 11486 79730 11546
rect 79790 11486 80750 11546
rect 80810 11486 81768 11546
rect 81828 11486 82788 11546
rect 82848 11486 83804 11546
rect 83864 11486 85840 11546
rect 69548 11480 69608 11486
rect 70572 11480 70632 11486
rect 71584 11480 71644 11486
rect 72604 11480 72664 11486
rect 73626 11480 73686 11486
rect 75662 11480 75722 11486
rect 77700 11480 77760 11486
rect 79730 11480 79790 11486
rect 80750 11480 80810 11486
rect 81768 11480 81828 11486
rect 82788 11480 82848 11486
rect 83804 11480 83864 11486
rect 85840 11480 85900 11486
rect 67286 11424 67346 11430
rect 74646 11424 74706 11430
rect 76680 11424 76740 11430
rect 78710 11424 78770 11430
rect 88710 11424 88770 20568
rect 67346 11364 74646 11424
rect 74706 11364 76680 11424
rect 76740 11364 78710 11424
rect 78770 11364 88770 11424
rect 67286 11358 67346 11364
rect 74646 11358 74706 11364
rect 76680 11358 76740 11364
rect 78710 11358 78770 11364
rect 69554 11312 69614 11318
rect 71590 11312 71650 11318
rect 87984 11312 88044 11318
rect 69614 11252 71590 11312
rect 71650 11252 87984 11312
rect 69554 11246 69614 11252
rect 71590 11246 71650 11252
rect 87984 11246 88044 11252
rect 87878 10424 87938 10430
rect 88838 10424 88898 20886
rect 70570 10406 70630 10412
rect 72606 10406 72666 10412
rect 80750 10406 80810 10412
rect 82786 10406 82846 10412
rect 86860 10406 86920 10412
rect 67398 10382 67458 10388
rect 68536 10382 68596 10388
rect 67458 10322 68536 10382
rect 68596 10322 69418 10382
rect 70630 10346 72606 10406
rect 72666 10346 80750 10406
rect 80810 10346 82786 10406
rect 82846 10346 86860 10406
rect 87938 10364 88898 10424
rect 87878 10358 87938 10364
rect 70570 10340 70630 10346
rect 72606 10340 72666 10346
rect 80750 10340 80810 10346
rect 82786 10340 82846 10346
rect 86860 10340 86920 10346
rect 67398 10316 67458 10322
rect 68536 10316 68596 10322
rect 67286 10182 67346 10188
rect 68534 10182 68594 10188
rect 67346 10122 68534 10182
rect 69358 10186 69418 10322
rect 69552 10302 69612 10308
rect 71592 10302 71652 10308
rect 73624 10302 73684 10308
rect 75658 10302 75718 10308
rect 77698 10302 77758 10308
rect 79732 10302 79792 10308
rect 69612 10242 71592 10302
rect 71652 10242 73624 10302
rect 73684 10242 75658 10302
rect 75718 10242 77698 10302
rect 77758 10242 79732 10302
rect 69552 10236 69612 10242
rect 71592 10236 71652 10242
rect 73624 10236 73684 10242
rect 75658 10236 75718 10242
rect 77698 10236 77758 10242
rect 79732 10236 79792 10242
rect 79928 10298 79988 10304
rect 84820 10298 84880 10304
rect 79988 10238 84820 10298
rect 88478 10294 88538 10300
rect 79928 10232 79988 10238
rect 84820 10232 84880 10238
rect 85318 10234 85324 10294
rect 85384 10234 88478 10294
rect 88478 10228 88538 10234
rect 70066 10188 70126 10194
rect 73624 10190 73684 10196
rect 75660 10190 75720 10196
rect 77696 10190 77756 10196
rect 79732 10190 79792 10196
rect 81766 10190 81826 10196
rect 83804 10190 83864 10196
rect 85844 10190 85904 10196
rect 88228 10190 88288 10196
rect 69358 10128 70066 10186
rect 70126 10128 71070 10188
rect 71130 10128 72082 10188
rect 72142 10128 73102 10188
rect 73162 10128 73168 10188
rect 73684 10130 75660 10190
rect 75720 10130 77696 10190
rect 77756 10130 79732 10190
rect 79792 10130 81766 10190
rect 81826 10130 83804 10190
rect 83864 10130 85844 10190
rect 85904 10130 88228 10190
rect 69358 10126 70408 10128
rect 70066 10122 70126 10126
rect 73624 10124 73684 10130
rect 75660 10124 75720 10130
rect 77696 10124 77756 10130
rect 79732 10124 79792 10130
rect 81766 10124 81826 10130
rect 83804 10124 83864 10130
rect 85844 10124 85904 10130
rect 88228 10124 88288 10130
rect 67286 10116 67346 10122
rect 68534 10116 68594 10122
rect 67180 10080 67240 10086
rect 74642 10080 74702 10086
rect 76676 10080 76736 10086
rect 78716 10080 78776 10086
rect 79928 10080 79988 10086
rect 66670 10020 67180 10080
rect 67240 10020 74642 10080
rect 74702 10020 76676 10080
rect 76736 10020 78716 10080
rect 78776 10020 79928 10080
rect 67180 10014 67240 10020
rect 74642 10014 74702 10020
rect 76676 10014 76736 10020
rect 78716 10014 78776 10020
rect 79928 10014 79988 10020
rect 80222 10082 80282 10088
rect 80282 10022 81250 10082
rect 81310 10022 81316 10082
rect 81768 10076 81828 10082
rect 83804 10076 83864 10082
rect 85842 10076 85902 10082
rect 87984 10076 88044 10082
rect 80222 10016 80282 10022
rect 81828 10016 83804 10076
rect 83864 10016 85842 10076
rect 85902 10016 87984 10076
rect 81768 10010 81828 10016
rect 83804 10010 83864 10016
rect 85842 10010 85902 10016
rect 87984 10010 88044 10016
rect 84316 9162 84376 9168
rect 68534 9150 68594 9156
rect 70572 9150 70632 9156
rect 72608 9150 72668 9156
rect 74640 9150 74700 9156
rect 68594 9090 70572 9150
rect 70632 9090 72608 9150
rect 72668 9090 74640 9150
rect 79216 9102 79222 9162
rect 79282 9102 84316 9162
rect 84316 9096 84376 9102
rect 84454 9166 84514 9172
rect 85336 9166 85396 9172
rect 86342 9166 86402 9172
rect 84514 9106 85336 9166
rect 85396 9106 86342 9166
rect 84454 9100 84514 9106
rect 85336 9100 85396 9106
rect 86342 9100 86402 9106
rect 86860 9162 86920 9168
rect 88112 9162 88172 9168
rect 86920 9102 88112 9162
rect 86860 9096 86920 9102
rect 88112 9096 88172 9102
rect 68534 9084 68594 9090
rect 70572 9084 70632 9090
rect 72608 9084 72668 9090
rect 74640 9084 74700 9090
rect 69040 9048 69100 9054
rect 74132 9048 74192 9054
rect 69100 8988 74132 9048
rect 69040 8982 69100 8988
rect 74132 8982 74192 8988
rect 78716 9034 78776 9040
rect 86860 9034 86920 9040
rect 78776 8974 86860 9034
rect 78716 8968 78776 8974
rect 86860 8968 86920 8974
rect 67286 8946 67346 8952
rect 70570 8946 70630 8952
rect 67346 8886 70570 8946
rect 67286 8880 67346 8886
rect 70570 8880 70630 8886
rect 71078 8940 71138 8946
rect 72100 8940 72160 8946
rect 73114 8940 73174 8946
rect 74132 8940 74192 8946
rect 75152 8940 75212 8946
rect 82264 8940 82324 8946
rect 83294 8940 83354 8946
rect 84454 8940 84514 8946
rect 71138 8880 72100 8940
rect 72160 8880 73114 8940
rect 73174 8880 74132 8940
rect 74192 8880 75152 8940
rect 75212 8880 82264 8940
rect 82324 8880 83294 8940
rect 83354 8880 84454 8940
rect 71078 8874 71138 8880
rect 72100 8874 72160 8880
rect 73114 8874 73174 8880
rect 74132 8874 74192 8880
rect 75152 8874 75212 8880
rect 82264 8874 82324 8880
rect 83294 8874 83354 8880
rect 84454 8874 84514 8880
rect 84822 8940 84882 8946
rect 88350 8940 88410 8946
rect 84882 8880 88350 8940
rect 84822 8874 84882 8880
rect 88350 8874 88410 8880
rect 69554 8846 69614 8852
rect 71588 8846 71648 8852
rect 73624 8846 73684 8852
rect 69614 8786 71588 8846
rect 71648 8786 73624 8846
rect 69554 8780 69614 8786
rect 71588 8780 71648 8786
rect 73624 8780 73684 8786
rect 80752 8836 80812 8842
rect 84822 8836 84882 8842
rect 80812 8776 84822 8836
rect 80752 8770 80812 8776
rect 84822 8770 84882 8776
rect 85838 8838 85898 8844
rect 88228 8838 88288 8844
rect 85898 8778 88228 8838
rect 85838 8772 85898 8778
rect 88228 8772 88288 8778
rect 75660 7928 75720 7934
rect 77696 7928 77756 7934
rect 79732 7928 79792 7934
rect 81770 7928 81830 7934
rect 69036 7922 69096 7928
rect 69946 7922 70006 7928
rect 70948 7922 71008 7928
rect 72100 7922 72160 7928
rect 73110 7922 73170 7928
rect 74116 7922 74176 7928
rect 75160 7922 75220 7928
rect 69096 7862 69946 7922
rect 70006 7862 70948 7922
rect 71008 7862 72100 7922
rect 72160 7862 73110 7922
rect 73170 7862 74116 7922
rect 74176 7862 75160 7922
rect 75720 7868 77696 7928
rect 77756 7868 79732 7928
rect 79792 7868 81770 7928
rect 75660 7862 75720 7868
rect 77696 7862 77756 7868
rect 79732 7862 79792 7868
rect 81770 7862 81830 7868
rect 83806 7928 83866 7934
rect 85844 7928 85904 7934
rect 83866 7868 85844 7928
rect 83806 7862 83866 7868
rect 85844 7862 85904 7868
rect 69036 7856 69096 7862
rect 69946 7856 70006 7862
rect 70948 7856 71008 7862
rect 72100 7856 72160 7862
rect 73110 7856 73170 7862
rect 74116 7856 74176 7862
rect 75160 7856 75220 7862
rect 71588 7820 71648 7826
rect 81762 7820 81822 7826
rect 83802 7820 83862 7826
rect 85840 7820 85900 7826
rect 71648 7760 81762 7820
rect 81822 7760 83802 7820
rect 83862 7760 85840 7820
rect 71588 7754 71648 7760
rect 81762 7754 81822 7760
rect 83802 7754 83862 7760
rect 85840 7754 85900 7760
rect 69036 7706 69096 7712
rect 71088 7706 71148 7712
rect 74114 7706 74174 7712
rect 75154 7706 75214 7712
rect 76168 7706 76228 7712
rect 77176 7706 77236 7712
rect 78220 7706 78280 7712
rect 79210 7706 79270 7712
rect 80228 7706 80288 7712
rect 81262 7706 81322 7712
rect 84294 7706 84354 7712
rect 85332 7706 85392 7712
rect 86358 7706 86418 7712
rect 69096 7646 70074 7706
rect 70134 7646 71088 7706
rect 71148 7646 74114 7706
rect 74174 7646 75154 7706
rect 75214 7646 76168 7706
rect 76228 7646 77176 7706
rect 77236 7646 78220 7706
rect 78280 7646 79210 7706
rect 79270 7646 80228 7706
rect 80288 7646 81262 7706
rect 81322 7646 84294 7706
rect 84354 7646 85332 7706
rect 85392 7646 86358 7706
rect 86418 7646 88476 7706
rect 88536 7646 88542 7706
rect 69036 7640 69096 7646
rect 71088 7640 71148 7646
rect 74114 7640 74174 7646
rect 75154 7640 75214 7646
rect 76168 7640 76228 7646
rect 77176 7640 77236 7646
rect 78220 7640 78280 7646
rect 79210 7640 79270 7646
rect 80228 7640 80288 7646
rect 81262 7640 81322 7646
rect 84294 7640 84354 7646
rect 85332 7640 85392 7646
rect 86358 7640 86418 7646
rect 74638 7602 74698 7608
rect 76680 7602 76740 7608
rect 78718 7602 78778 7608
rect 80752 7602 80812 7608
rect 82786 7604 82846 7610
rect 84820 7604 84880 7610
rect 86862 7604 86922 7610
rect 88112 7604 88172 7610
rect 67394 7542 67400 7602
rect 67460 7542 74638 7602
rect 74698 7542 76680 7602
rect 76740 7542 78718 7602
rect 78778 7542 80752 7602
rect 74638 7536 74698 7542
rect 76680 7536 76740 7542
rect 78718 7536 78778 7542
rect 80752 7536 80812 7542
rect 81264 7598 81324 7604
rect 82286 7598 82346 7604
rect 81324 7538 82286 7598
rect 82846 7544 84820 7604
rect 84880 7544 86862 7604
rect 86922 7544 88112 7604
rect 82786 7538 82846 7544
rect 84820 7538 84880 7544
rect 86862 7538 86922 7544
rect 88112 7538 88172 7544
rect 81264 7532 81324 7538
rect 82286 7532 82346 7538
rect 73628 6700 73688 6706
rect 77696 6700 77756 6706
rect 79730 6700 79790 6706
rect 69034 6694 69094 6700
rect 70042 6694 70102 6700
rect 71056 6694 71116 6700
rect 72094 6694 72154 6700
rect 73112 6694 73172 6700
rect 69094 6634 70042 6694
rect 70102 6634 71056 6694
rect 71116 6634 72094 6694
rect 72154 6634 73112 6694
rect 73688 6640 75664 6700
rect 75724 6640 77696 6700
rect 77756 6640 79730 6700
rect 73628 6634 73688 6640
rect 77696 6634 77756 6640
rect 79730 6634 79790 6640
rect 80752 6702 80812 6708
rect 81106 6702 81166 6708
rect 80812 6642 81106 6702
rect 80752 6636 80812 6642
rect 81106 6636 81166 6642
rect 84824 6702 84884 6708
rect 88108 6702 88168 6708
rect 84884 6642 88108 6702
rect 84824 6636 84884 6642
rect 88108 6636 88168 6642
rect 69034 6628 69094 6634
rect 70042 6628 70102 6634
rect 71056 6628 71116 6634
rect 72094 6628 72154 6634
rect 73112 6628 73172 6634
rect 67180 6590 67240 6596
rect 68536 6590 68596 6596
rect 76680 6590 76740 6596
rect 78716 6590 78776 6596
rect 80748 6590 80808 6596
rect 67240 6530 68536 6590
rect 68596 6530 76680 6590
rect 76740 6530 78716 6590
rect 78776 6530 80748 6590
rect 67180 6524 67240 6530
rect 68536 6524 68596 6530
rect 76680 6524 76740 6530
rect 78716 6524 78776 6530
rect 80748 6524 80808 6530
rect 80258 6492 80318 6498
rect 81296 6492 81356 6498
rect 82272 6492 82332 6498
rect 83288 6492 83348 6498
rect 85314 6492 85374 6498
rect 86344 6492 86404 6498
rect 64636 6410 66596 6470
rect 69552 6478 69612 6484
rect 71590 6478 71650 6484
rect 75662 6478 75722 6484
rect 69612 6418 71590 6478
rect 71650 6418 75662 6478
rect 80318 6432 81296 6492
rect 81356 6432 82272 6492
rect 82332 6432 83288 6492
rect 83348 6432 85314 6492
rect 85374 6432 86344 6492
rect 80258 6426 80318 6432
rect 81296 6426 81356 6432
rect 82272 6426 82332 6432
rect 83288 6426 83348 6432
rect 85314 6426 85374 6432
rect 86344 6426 86404 6432
rect 69552 6412 69612 6418
rect 71590 6412 71650 6418
rect 75662 6412 75722 6418
rect 64576 6404 64636 6410
rect 64358 6380 64418 6386
rect 63982 6320 64358 6380
rect 68532 6380 68592 6386
rect 70570 6380 70630 6386
rect 72610 6380 72670 6386
rect 74646 6380 74706 6386
rect 80750 6380 80810 6386
rect 81100 6380 81106 6384
rect 67286 6344 67346 6350
rect 63922 6314 63982 6320
rect 64358 6314 64418 6320
rect 65164 6284 65170 6344
rect 65230 6284 67286 6344
rect 68592 6320 70570 6380
rect 70630 6320 72610 6380
rect 72670 6320 74646 6380
rect 74706 6324 81106 6380
rect 81166 6380 81172 6384
rect 82786 6380 82846 6386
rect 84822 6380 84882 6386
rect 86858 6380 86918 6386
rect 81166 6324 82786 6380
rect 74706 6320 82786 6324
rect 82846 6320 84822 6380
rect 84882 6320 86858 6380
rect 68532 6314 68592 6320
rect 70570 6314 70630 6320
rect 72610 6314 72670 6320
rect 74646 6314 74706 6320
rect 80750 6314 80810 6320
rect 82786 6314 82846 6320
rect 84822 6314 84882 6320
rect 86858 6314 86918 6320
rect 67286 6278 67346 6284
rect 63158 6270 63218 6276
rect 63378 6270 63438 6276
rect 64032 6270 64092 6276
rect 64248 6270 64308 6276
rect 63218 6210 63378 6270
rect 63438 6210 64032 6270
rect 64092 6210 64248 6270
rect 63158 6204 63218 6210
rect 63378 6204 63438 6210
rect 64032 6204 64092 6210
rect 64248 6204 64308 6210
rect 62482 5766 62542 5772
rect 62940 5766 63000 5772
rect 63596 5766 63656 5772
rect 62542 5706 62940 5766
rect 63000 5706 63596 5766
rect 62482 5700 62542 5706
rect 62940 5700 63000 5706
rect 63596 5700 63656 5706
rect 64140 5766 64200 5772
rect 64928 5766 64988 5772
rect 64200 5706 64928 5766
rect 64140 5700 64200 5706
rect 64928 5700 64988 5706
rect 62352 5644 62412 5650
rect 63158 5644 63218 5650
rect 63376 5644 63436 5650
rect 62412 5584 63158 5644
rect 63218 5584 63376 5644
rect 62352 5578 62412 5584
rect 63158 5578 63218 5584
rect 63376 5578 63436 5584
rect 63812 5646 63872 5652
rect 64468 5646 64528 5652
rect 63872 5586 64468 5646
rect 63812 5580 63872 5586
rect 64468 5580 64528 5586
rect 62832 5520 62892 5526
rect 63702 5520 63762 5526
rect 64574 5520 64634 5526
rect 62892 5460 63702 5520
rect 63762 5460 64574 5520
rect 75658 5476 75718 5482
rect 77700 5476 77760 5482
rect 79732 5476 79792 5482
rect 81772 5476 81832 5482
rect 88228 5476 88288 5482
rect 62832 5454 62892 5460
rect 63702 5454 63762 5460
rect 64574 5454 64634 5460
rect 69552 5456 69612 5462
rect 71588 5456 71648 5462
rect 73626 5456 73686 5462
rect 63270 5394 63330 5400
rect 65048 5394 65108 5400
rect 63330 5334 65048 5394
rect 69612 5396 71588 5456
rect 71648 5396 73626 5456
rect 75482 5416 75488 5476
rect 75548 5416 75658 5476
rect 75718 5416 77700 5476
rect 77760 5416 79732 5476
rect 79792 5416 81772 5476
rect 81832 5416 88228 5476
rect 75658 5410 75718 5416
rect 77700 5410 77760 5416
rect 79732 5410 79792 5416
rect 81772 5410 81832 5416
rect 88228 5410 88288 5416
rect 69552 5390 69612 5396
rect 71588 5390 71648 5396
rect 73626 5390 73686 5396
rect 80750 5378 80810 5384
rect 86856 5378 86916 5384
rect 88108 5378 88168 5384
rect 63270 5328 63330 5334
rect 65048 5328 65108 5334
rect 67398 5358 67458 5364
rect 70570 5358 70630 5364
rect 67458 5298 70570 5358
rect 67398 5292 67458 5298
rect 70570 5292 70630 5298
rect 72094 5358 72154 5364
rect 75142 5358 75202 5364
rect 72154 5298 73116 5358
rect 73176 5298 74138 5358
rect 74198 5298 75142 5358
rect 80810 5318 86856 5378
rect 86916 5318 88108 5378
rect 80750 5312 80810 5318
rect 86856 5312 86916 5318
rect 88108 5312 88168 5318
rect 72094 5292 72154 5298
rect 75142 5292 75202 5298
rect 63604 5280 63656 5286
rect 67186 5278 67192 5280
rect 63656 5230 67192 5278
rect 67186 5228 67192 5230
rect 67244 5228 67250 5280
rect 75664 5268 75724 5274
rect 77692 5268 77752 5274
rect 79736 5268 79796 5274
rect 81764 5268 81824 5274
rect 83802 5268 83862 5274
rect 85842 5268 85902 5274
rect 69556 5262 69616 5268
rect 71592 5262 71652 5268
rect 73620 5262 73680 5268
rect 75488 5262 75548 5268
rect 63604 5222 63656 5228
rect 69616 5202 71592 5262
rect 71652 5202 73620 5262
rect 73680 5202 75488 5262
rect 75724 5208 77692 5268
rect 77752 5208 79736 5268
rect 79796 5208 81764 5268
rect 81824 5208 83802 5268
rect 83862 5208 85842 5268
rect 75664 5202 75724 5208
rect 77692 5202 77752 5208
rect 79736 5202 79796 5208
rect 81764 5202 81824 5208
rect 83802 5202 83862 5208
rect 85842 5202 85902 5208
rect 86360 5272 86420 5278
rect 88478 5272 88538 5278
rect 86420 5212 88478 5272
rect 86360 5206 86420 5212
rect 88478 5206 88538 5212
rect 69556 5196 69616 5202
rect 71592 5196 71652 5202
rect 73620 5196 73680 5202
rect 75488 5196 75548 5202
rect 68538 5142 68598 5148
rect 72606 5142 72666 5148
rect 74640 5142 74700 5148
rect 82790 5142 82850 5148
rect 84820 5142 84880 5148
rect 86858 5144 86918 5150
rect 88350 5144 88410 5150
rect 68598 5082 72606 5142
rect 72666 5082 74640 5142
rect 74700 5082 82790 5142
rect 82850 5082 84820 5142
rect 85340 5084 85346 5144
rect 85406 5084 86858 5144
rect 86918 5084 88350 5144
rect 68538 5076 68598 5082
rect 72606 5076 72666 5082
rect 74640 5076 74700 5082
rect 82790 5076 82850 5082
rect 84820 5076 84880 5082
rect 86858 5078 86918 5084
rect 88350 5078 88410 5084
rect 64018 5060 64078 5066
rect 65212 5060 65272 5066
rect 65902 5060 65962 5066
rect 62822 5000 62828 5060
rect 62888 5000 64018 5060
rect 64078 5000 65212 5060
rect 65272 5000 65902 5060
rect 64018 4994 64078 5000
rect 65212 4994 65272 5000
rect 65902 4994 65962 5000
rect 62280 4960 62340 4966
rect 63272 4960 63332 4966
rect 63570 4960 63630 4966
rect 64466 4960 64526 4966
rect 64762 4960 64822 4966
rect 62340 4900 63272 4960
rect 63332 4900 63570 4960
rect 63630 4900 64466 4960
rect 64526 4900 64762 4960
rect 62280 4894 62340 4900
rect 63272 4894 63332 4900
rect 63570 4894 63630 4900
rect 64466 4894 64526 4900
rect 64762 4894 64822 4900
rect 66017 4876 66026 4936
rect 66086 4876 66095 4936
rect 63121 4057 63179 4063
rect 63725 4057 63783 4063
rect 64316 4057 64374 4063
rect 63179 3999 63725 4057
rect 63783 3999 64316 4057
rect 64374 3999 64913 4057
rect 64971 3999 65509 4057
rect 65567 3999 65573 4057
rect 63121 3993 63179 3999
rect 63725 3993 63783 3999
rect 64316 3993 64374 3999
rect 62408 3926 62468 3932
rect 63418 3926 63478 3932
rect 64016 3926 64076 3932
rect 64610 3926 64670 3932
rect 65208 3926 65268 3932
rect 62468 3866 62824 3926
rect 62884 3866 63418 3926
rect 63478 3866 64016 3926
rect 64076 3866 64610 3926
rect 64670 3866 65208 3926
rect 62408 3860 62468 3866
rect 63418 3860 63478 3866
rect 64016 3860 64076 3866
rect 64610 3860 64670 3866
rect 65208 3860 65268 3866
rect 62976 3818 63036 3824
rect 63274 3818 63334 3824
rect 63574 3818 63634 3824
rect 63868 3818 63928 3824
rect 64164 3818 64224 3824
rect 64464 3818 64524 3824
rect 64766 3818 64826 3824
rect 65056 3818 65116 3824
rect 65360 3818 65420 3824
rect 66026 3818 66086 4876
rect 67286 4226 67346 4232
rect 76674 4226 76734 4232
rect 78716 4226 78776 4232
rect 80752 4226 80812 4232
rect 67346 4166 76674 4226
rect 76734 4166 78716 4226
rect 78776 4166 80752 4226
rect 67286 4160 67346 4166
rect 76674 4160 76734 4166
rect 78716 4160 78776 4166
rect 80752 4160 80812 4166
rect 83806 4226 83866 4232
rect 85838 4226 85898 4232
rect 87984 4226 88044 4232
rect 83866 4166 85838 4226
rect 85898 4166 87984 4226
rect 83806 4160 83866 4166
rect 85838 4160 85898 4166
rect 87984 4160 88044 4166
rect 71090 4112 71150 4118
rect 76170 4112 76230 4118
rect 67180 4100 67240 4106
rect 70570 4100 70630 4106
rect 67240 4040 70570 4100
rect 71150 4052 76170 4112
rect 71090 4046 71150 4052
rect 76170 4046 76230 4052
rect 81258 4116 81318 4122
rect 86358 4116 86418 4122
rect 81318 4056 86358 4116
rect 81258 4050 81318 4056
rect 86358 4050 86418 4056
rect 67180 4034 67240 4040
rect 70570 4034 70630 4040
rect 69552 3990 69612 3996
rect 71588 3990 71648 3996
rect 72608 3990 72668 3996
rect 73624 3990 73684 3996
rect 74644 3990 74704 3996
rect 75662 3990 75722 3996
rect 77692 3990 77752 3996
rect 79730 3990 79790 3996
rect 81766 3990 81826 3996
rect 82788 3990 82848 3996
rect 83808 3990 83868 3996
rect 84822 3990 84882 3996
rect 85844 3990 85904 3996
rect 69612 3930 71588 3990
rect 71648 3930 72608 3990
rect 72668 3930 73624 3990
rect 73684 3930 74644 3990
rect 74704 3930 75662 3990
rect 75722 3930 77692 3990
rect 77752 3930 79730 3990
rect 79790 3930 81766 3990
rect 81826 3930 82788 3990
rect 82848 3930 83808 3990
rect 83868 3930 84822 3990
rect 84882 3930 85844 3990
rect 69552 3924 69612 3930
rect 71588 3924 71648 3930
rect 72608 3924 72668 3930
rect 73624 3924 73684 3930
rect 74644 3924 74704 3930
rect 75662 3924 75722 3930
rect 77692 3924 77752 3930
rect 79730 3924 79790 3930
rect 81766 3924 81826 3930
rect 82788 3924 82848 3930
rect 83808 3924 83868 3930
rect 84822 3924 84882 3930
rect 85844 3924 85904 3930
rect 71206 3896 71266 3902
rect 72090 3896 72150 3902
rect 73112 3896 73172 3902
rect 75154 3896 75214 3902
rect 71266 3836 72090 3896
rect 72150 3836 73112 3896
rect 73172 3836 75154 3896
rect 71206 3830 71266 3836
rect 72090 3830 72150 3836
rect 73112 3830 73172 3836
rect 75154 3830 75214 3836
rect 82276 3896 82336 3902
rect 83296 3896 83356 3902
rect 84310 3896 84370 3902
rect 85346 3896 85406 3902
rect 82336 3836 83296 3896
rect 83356 3836 84310 3896
rect 84370 3836 85346 3896
rect 82276 3830 82336 3836
rect 83296 3830 83356 3836
rect 84310 3830 84370 3836
rect 85346 3830 85406 3836
rect 63036 3758 63274 3818
rect 63334 3758 63574 3818
rect 63634 3758 63868 3818
rect 63928 3758 64164 3818
rect 64224 3758 64464 3818
rect 64524 3758 64766 3818
rect 64826 3758 65056 3818
rect 65116 3758 65360 3818
rect 65420 3758 66026 3818
rect 66086 3758 66092 3818
rect 62976 3752 63036 3758
rect 63274 3752 63334 3758
rect 63574 3752 63634 3758
rect 63868 3752 63928 3758
rect 64164 3752 64224 3758
rect 64464 3752 64524 3758
rect 64766 3752 64826 3758
rect 65056 3752 65116 3758
rect 65360 3752 65420 3758
rect 66926 2996 66986 3002
rect 67518 2996 67578 3002
rect 68032 2996 68092 3002
rect 68530 2996 68590 3002
rect 70572 2996 70632 3002
rect 72604 2996 72664 3002
rect 74636 2996 74696 3002
rect 78894 2996 78900 2998
rect 66494 2994 66926 2996
rect 56756 2864 58582 2924
rect 58642 2864 60452 2924
rect 60512 2864 61914 2924
rect 62153 2933 62243 2942
rect 56696 2858 56756 2864
rect 58582 2858 58642 2864
rect 60452 2858 60512 2864
rect 66350 2936 66926 2994
rect 66986 2936 67518 2996
rect 67578 2936 68032 2996
rect 68092 2936 68530 2996
rect 68590 2936 70572 2996
rect 70632 2936 72604 2996
rect 72664 2936 74636 2996
rect 74696 2936 76540 2996
rect 76600 2938 78900 2996
rect 78960 2996 78966 2998
rect 80750 2996 80810 3002
rect 82784 2996 82844 3002
rect 84818 2996 84878 3002
rect 86860 2996 86920 3002
rect 87372 2996 87432 3002
rect 87878 2996 87938 3002
rect 78960 2938 80750 2996
rect 76600 2936 80750 2938
rect 80810 2936 82784 2996
rect 82844 2936 84818 2996
rect 84878 2936 86860 2996
rect 86920 2936 87372 2996
rect 87432 2936 87878 2996
rect 66350 2934 66586 2936
rect 62280 2920 62340 2926
rect 62974 2920 63034 2926
rect 63870 2920 63930 2926
rect 64164 2920 64224 2926
rect 65058 2920 65118 2926
rect 65360 2920 65420 2926
rect 62243 2860 62280 2920
rect 62340 2860 62974 2920
rect 63034 2860 63870 2920
rect 63930 2860 64164 2920
rect 64224 2860 65058 2920
rect 65118 2860 65360 2920
rect 62280 2854 62340 2860
rect 62974 2854 63034 2860
rect 63870 2854 63930 2860
rect 64164 2854 64224 2860
rect 65058 2854 65118 2860
rect 65360 2854 65420 2860
rect 62153 2834 62243 2843
rect 56548 2816 56608 2822
rect 58584 2816 58644 2822
rect 60620 2816 60680 2822
rect 56608 2756 58584 2816
rect 58644 2756 60620 2816
rect 56548 2750 56608 2756
rect 58584 2750 58644 2756
rect 60620 2750 60680 2756
rect 63420 2812 63480 2818
rect 64614 2812 64674 2818
rect 63480 2752 64614 2812
rect 64674 2752 65902 2812
rect 65962 2752 65968 2812
rect 63420 2746 63480 2752
rect 64614 2746 64674 2752
rect 57566 2704 57626 2710
rect 57626 2644 59604 2704
rect 59664 2644 59670 2704
rect 57566 2638 57626 2644
rect 63122 1828 63182 1834
rect 63716 1828 63776 1834
rect 64316 1828 64376 1834
rect 64910 1828 64970 1834
rect 65504 1828 65564 1834
rect 66350 1828 66410 2934
rect 66926 2930 66986 2936
rect 67518 2930 67578 2936
rect 68032 2930 68092 2936
rect 68530 2930 68590 2936
rect 70572 2930 70632 2936
rect 72604 2930 72664 2936
rect 74636 2930 74696 2936
rect 80750 2930 80810 2936
rect 82784 2930 82844 2936
rect 84818 2930 84878 2936
rect 86860 2930 86920 2936
rect 87372 2930 87432 2936
rect 87878 2930 87938 2936
rect 71080 2884 71140 2890
rect 72092 2884 72152 2890
rect 73106 2884 73166 2890
rect 76018 2884 76078 2890
rect 71140 2824 72092 2884
rect 72152 2824 73106 2884
rect 73166 2824 76018 2884
rect 71080 2818 71140 2824
rect 72092 2818 72152 2824
rect 73106 2818 73166 2824
rect 76018 2818 76078 2824
rect 76678 2886 76738 2892
rect 67060 2778 67120 2784
rect 69046 2778 69106 2784
rect 70068 2778 70128 2784
rect 72606 2778 72666 2784
rect 73118 2778 73178 2784
rect 74136 2778 74196 2784
rect 74642 2778 74702 2784
rect 75148 2778 75208 2784
rect 76160 2778 76220 2784
rect 76678 2778 76738 2826
rect 77306 2882 77366 2888
rect 78352 2882 78412 2888
rect 82280 2882 82340 2888
rect 83298 2882 83358 2888
rect 77366 2822 78352 2882
rect 78412 2822 82280 2882
rect 82340 2822 83298 2882
rect 83358 2822 84308 2882
rect 84368 2822 84374 2882
rect 77306 2816 77366 2822
rect 78352 2816 78412 2822
rect 82280 2816 82340 2822
rect 83298 2816 83358 2822
rect 77180 2778 77240 2784
rect 78202 2778 78262 2784
rect 78714 2778 78774 2784
rect 79220 2778 79280 2784
rect 80238 2778 80298 2784
rect 80750 2778 80810 2784
rect 81258 2778 81318 2784
rect 85330 2778 85390 2784
rect 86332 2778 86392 2784
rect 67120 2718 69046 2778
rect 69106 2718 70068 2778
rect 70128 2718 72606 2778
rect 72666 2718 73118 2778
rect 73178 2718 74136 2778
rect 74196 2718 74642 2778
rect 74702 2718 75148 2778
rect 75208 2718 76160 2778
rect 76220 2718 77180 2778
rect 77240 2718 78202 2778
rect 78262 2718 78714 2778
rect 78774 2718 79220 2778
rect 79280 2718 80238 2778
rect 80298 2718 80750 2778
rect 80810 2718 81258 2778
rect 81318 2718 85330 2778
rect 85390 2718 86332 2778
rect 67060 2712 67120 2718
rect 69046 2712 69106 2718
rect 70068 2712 70128 2718
rect 72606 2712 72666 2718
rect 73118 2712 73178 2718
rect 74136 2712 74196 2718
rect 74642 2712 74702 2718
rect 75148 2712 75208 2718
rect 76160 2712 76220 2718
rect 77180 2712 77240 2718
rect 78202 2712 78262 2718
rect 78714 2712 78774 2718
rect 79220 2712 79280 2718
rect 80238 2712 80298 2718
rect 80750 2712 80810 2718
rect 81258 2712 81318 2718
rect 85330 2712 85390 2718
rect 86332 2712 86392 2718
rect 66654 2674 66714 2680
rect 71082 2674 71142 2680
rect 71586 2674 71646 2680
rect 72102 2674 72162 2680
rect 73624 2674 73684 2680
rect 75662 2674 75722 2680
rect 77698 2674 77758 2680
rect 79734 2674 79794 2680
rect 81766 2674 81826 2680
rect 82288 2674 82348 2680
rect 82788 2674 82848 2680
rect 83296 2674 83356 2680
rect 83804 2674 83864 2680
rect 84154 2674 84214 2680
rect 88756 2674 88816 2680
rect 66714 2614 71082 2674
rect 71142 2614 71586 2674
rect 71646 2614 72102 2674
rect 72162 2614 73624 2674
rect 73684 2614 75662 2674
rect 75722 2614 77698 2674
rect 77758 2614 79734 2674
rect 79794 2614 81766 2674
rect 81826 2614 82288 2674
rect 82348 2614 82788 2674
rect 82848 2614 83296 2674
rect 83356 2614 83804 2674
rect 83864 2614 84154 2674
rect 84214 2614 88756 2674
rect 66654 2608 66714 2614
rect 71082 2608 71142 2614
rect 71586 2608 71646 2614
rect 72102 2608 72162 2614
rect 73624 2608 73684 2614
rect 75662 2608 75722 2614
rect 77698 2608 77758 2614
rect 79734 2608 79794 2614
rect 81766 2608 81826 2614
rect 82288 2608 82348 2614
rect 82788 2608 82848 2614
rect 83296 2608 83356 2614
rect 83804 2608 83864 2614
rect 84154 2608 84214 2614
rect 88756 2608 88816 2614
rect 57568 1822 57628 1828
rect 57628 1762 59598 1822
rect 59658 1762 59664 1822
rect 63182 1768 63716 1828
rect 63776 1768 64316 1828
rect 64376 1768 64910 1828
rect 64970 1768 65504 1828
rect 65564 1768 66410 1828
rect 63122 1762 63182 1768
rect 63716 1762 63776 1768
rect 64316 1762 64376 1768
rect 64910 1762 64970 1768
rect 65504 1762 65564 1768
rect 57568 1756 57628 1762
rect 76680 1742 76740 1748
rect 78716 1742 78776 1748
rect 63416 1734 63476 1740
rect 64014 1734 64074 1740
rect 64612 1734 64672 1740
rect 65212 1734 65272 1740
rect 56550 1720 56610 1726
rect 60618 1720 60678 1726
rect 61748 1720 61808 1726
rect 56610 1660 60618 1720
rect 60678 1660 61748 1720
rect 62518 1674 62524 1734
rect 62584 1674 63416 1734
rect 63476 1674 64014 1734
rect 64074 1674 64612 1734
rect 64672 1674 65212 1734
rect 76740 1682 78716 1742
rect 76680 1676 76740 1682
rect 78716 1676 78776 1682
rect 63416 1668 63476 1674
rect 64014 1668 64074 1674
rect 64612 1668 64672 1674
rect 65212 1668 65272 1674
rect 56550 1654 56610 1660
rect 60618 1654 60678 1660
rect 61748 1654 61808 1660
rect 62972 1626 63032 1632
rect 63270 1626 63330 1632
rect 63566 1626 63626 1632
rect 63870 1626 63930 1632
rect 64166 1626 64226 1632
rect 64464 1626 64524 1632
rect 64760 1626 64820 1632
rect 65056 1626 65116 1632
rect 65360 1626 65420 1632
rect 66026 1626 66086 1632
rect 50553 1514 50627 1574
rect 50687 1514 50693 1574
rect 50939 1536 50945 1596
rect 51005 1536 51160 1596
rect 55412 1614 55472 1620
rect 58584 1614 58644 1620
rect 55472 1554 58584 1614
rect 63032 1566 63270 1626
rect 63330 1566 63566 1626
rect 63626 1566 63870 1626
rect 63930 1566 64166 1626
rect 64226 1566 64464 1626
rect 64524 1566 64760 1626
rect 64820 1566 65056 1626
rect 65116 1566 65360 1626
rect 65420 1566 66026 1626
rect 62972 1560 63032 1566
rect 63270 1560 63330 1566
rect 63566 1560 63626 1566
rect 63870 1560 63930 1566
rect 64166 1560 64226 1566
rect 64464 1560 64524 1566
rect 64760 1560 64820 1566
rect 65056 1560 65116 1566
rect 65360 1560 65420 1566
rect 66026 1560 66086 1566
rect 55412 1548 55472 1554
rect 58584 1548 58644 1554
rect 68530 1542 68590 1548
rect 70568 1542 70628 1548
rect 72606 1542 72666 1548
rect 74638 1542 74698 1548
rect 76676 1542 76736 1548
rect 78710 1542 78770 1548
rect 80750 1542 80810 1548
rect 82784 1542 82844 1548
rect 84818 1542 84878 1548
rect 86856 1542 86916 1548
rect 88598 1542 88658 1548
rect 49048 1497 49108 1503
rect 49564 1497 49624 1503
rect 13518 1444 13578 1450
rect 15548 1444 15608 1450
rect 17586 1444 17646 1450
rect 19622 1444 19682 1450
rect 21658 1444 21718 1450
rect 23694 1444 23754 1450
rect 25728 1444 25788 1450
rect 27764 1444 27824 1450
rect 29804 1444 29864 1450
rect 31838 1444 31898 1450
rect 33874 1444 33934 1450
rect 13578 1384 15548 1444
rect 15608 1384 17586 1444
rect 17646 1384 19622 1444
rect 19682 1384 21658 1444
rect 21718 1384 23694 1444
rect 23754 1384 25728 1444
rect 25788 1384 27764 1444
rect 27824 1384 29804 1444
rect 29864 1384 31838 1444
rect 31898 1384 33874 1444
rect 46088 1437 49048 1497
rect 49108 1437 49564 1497
rect 49624 1437 50082 1497
rect 50142 1437 50148 1497
rect 49048 1431 49108 1437
rect 49564 1431 49624 1437
rect 13518 1378 13578 1384
rect 15548 1378 15608 1384
rect 17586 1378 17646 1384
rect 19622 1378 19682 1384
rect 21658 1378 21718 1384
rect 23694 1378 23754 1384
rect 25728 1378 25788 1384
rect 27764 1378 27824 1384
rect 29804 1378 29864 1384
rect 31838 1378 31898 1384
rect 33874 1378 33934 1384
rect 49952 949 50012 955
rect 50945 950 51005 1536
rect 68590 1482 70568 1542
rect 70628 1482 72606 1542
rect 72666 1482 74638 1542
rect 74698 1482 76676 1542
rect 76736 1482 78710 1542
rect 78770 1482 80750 1542
rect 80810 1482 82784 1542
rect 82844 1482 84818 1542
rect 84878 1482 86856 1542
rect 86916 1482 88598 1542
rect 68530 1476 68590 1482
rect 70568 1476 70628 1482
rect 72606 1476 72666 1482
rect 74638 1476 74698 1482
rect 76676 1476 76736 1482
rect 78710 1476 78770 1482
rect 80750 1476 80810 1482
rect 82784 1476 82844 1482
rect 84818 1476 84878 1482
rect 86856 1476 86916 1482
rect 88598 1476 88658 1482
rect 67518 1444 67578 1450
rect 69548 1444 69608 1450
rect 71586 1444 71646 1450
rect 73622 1444 73682 1450
rect 75658 1444 75718 1450
rect 77694 1444 77754 1450
rect 79728 1444 79788 1450
rect 81764 1444 81824 1450
rect 83804 1444 83864 1450
rect 85838 1444 85898 1450
rect 87874 1444 87934 1450
rect 67578 1384 69548 1444
rect 69608 1384 71586 1444
rect 71646 1384 73622 1444
rect 73682 1384 75658 1444
rect 75718 1384 77694 1444
rect 77754 1384 79728 1444
rect 79788 1384 81764 1444
rect 81824 1384 83804 1444
rect 83864 1384 85838 1444
rect 85898 1384 87874 1444
rect 67518 1378 67578 1384
rect 69548 1378 69608 1384
rect 71586 1378 71646 1384
rect 73622 1378 73682 1384
rect 75658 1378 75718 1384
rect 77694 1378 77754 1384
rect 79728 1378 79788 1384
rect 81764 1378 81824 1384
rect 83804 1378 83864 1384
rect 85838 1378 85898 1384
rect 87874 1378 87934 1384
rect 50459 949 51005 950
rect 50012 890 51005 949
rect 50012 889 50563 890
rect 49952 883 50012 889
rect 8280 700 8340 706
rect 9270 700 9330 706
rect 9568 700 9628 706
rect 10464 700 10524 706
rect 10766 700 10826 706
rect 8340 640 9270 700
rect 9330 640 9568 700
rect 9628 640 10464 700
rect 10524 640 10766 700
rect 62280 700 62340 706
rect 63270 700 63330 706
rect 63568 700 63628 706
rect 64464 700 64524 706
rect 64766 700 64826 706
rect 8280 634 8340 640
rect 9270 634 9330 640
rect 9568 634 9628 640
rect 10464 634 10524 640
rect 10766 634 10826 640
rect 57054 670 57114 676
rect 58080 670 58140 676
rect 59104 670 59164 676
rect 57114 610 58080 670
rect 58140 610 59104 670
rect 59164 610 60004 670
rect 60064 610 60070 670
rect 62340 640 63270 700
rect 63330 640 63568 700
rect 63628 640 64464 700
rect 64524 640 64766 700
rect 62280 634 62340 640
rect 63270 634 63330 640
rect 63568 634 63628 640
rect 64464 634 64524 640
rect 64766 634 64826 640
rect 8824 600 8884 606
rect 10012 600 10072 606
rect 11208 600 11268 606
rect 11902 600 11962 606
rect 57054 604 57114 610
rect 58080 604 58140 610
rect 59104 604 59164 610
rect 8033 522 8042 582
rect 8102 522 8111 582
rect 8884 540 10012 600
rect 10072 540 11208 600
rect 11268 540 11902 600
rect 8824 534 8884 540
rect 10012 534 10072 540
rect 11208 534 11268 540
rect 11902 534 11962 540
rect 62824 600 62884 606
rect 64012 600 64072 606
rect 65208 600 65268 606
rect 65902 600 65962 606
rect 62884 540 64012 600
rect 64072 540 65208 600
rect 65268 540 65902 600
rect 62824 534 62884 540
rect 64012 534 64072 540
rect 65208 534 65268 540
rect 65902 534 65962 540
rect 3432 64 34918 110
rect 3432 -90 3478 64
rect 34878 -90 34918 64
rect 3432 -136 34918 -90
rect 57432 64 88918 110
rect 57432 -90 57478 64
rect 88878 -90 88918 64
rect 57432 -136 88918 -90
rect -1266 -276 -666 -266
rect -1266 -586 -666 -576
rect 35166 -276 35766 -266
rect 35166 -586 35766 -576
rect 52734 -276 53334 -266
rect 52734 -586 53334 -576
rect 89166 -276 89766 -266
rect 89166 -586 89766 -576
<< via2 >>
rect 11434 27856 12034 28156
rect 35066 27856 35666 28156
rect 65434 27856 66034 28156
rect 89066 27856 89666 28156
rect -1414 27582 -1354 27642
rect 15011 27560 31796 27774
rect 47824 27564 48000 27680
rect 48000 27564 48306 27680
rect 48306 27564 48462 27680
rect 69011 27560 85796 27774
rect 48398 24604 48458 24664
rect 47624 24455 47682 24515
rect 47682 24455 47684 24515
rect 42790 23874 42850 23934
rect 11211 18823 11301 18913
rect 10962 16318 11062 16418
rect -13286 15325 -13226 15385
rect -10620 15325 -10560 15385
rect -13467 14515 -13377 14605
rect -1077 15267 -987 15357
rect 717 15267 807 15357
rect 3317 15267 3407 15357
rect 5917 15269 6007 15359
rect 8517 15269 8607 15359
rect 10321 15269 10411 15359
rect -1924 15092 -1864 15152
rect 11206 15782 11306 15882
rect 10967 14893 11057 14983
rect 11206 14712 11306 14812
rect -9878 13060 -9818 13120
rect -9955 10939 -9851 11043
rect -5821 10931 -5725 11027
rect -8781 10611 -8667 10725
rect -4789 10609 -4683 10715
rect 38879 23781 38959 23861
rect 41001 23437 41091 23527
rect 47876 22604 47880 22664
rect 47880 22604 47936 22664
rect 48656 22455 48716 22515
rect 42800 21860 42860 21920
rect 40228 21314 40328 21414
rect 11382 7138 11442 7198
rect -10815 3741 -10721 3835
rect -6737 3737 -6647 3827
rect -9010 3410 -8906 3514
rect -4636 3410 -4536 3510
rect 13277 18823 13367 18913
rect 12655 16327 12745 16417
rect 65093 18823 65183 18913
rect 38973 17731 39071 17829
rect 43139 17723 43257 17841
rect 47331 17731 47431 17831
rect 40994 17408 41102 17516
rect 45188 17398 45316 17526
rect 49283 17397 49393 17507
rect 36259 16103 36349 16193
rect 52923 15267 53013 15357
rect 54717 15267 54807 15357
rect 57317 15267 57407 15357
rect 59917 15269 60007 15359
rect 62517 15269 62607 15359
rect 64321 15269 64411 15359
rect 65088 14638 65188 14738
rect 36456 13714 36556 13814
rect 39253 13719 39343 13809
rect 38849 11615 38945 11711
rect 42999 11597 43125 11727
rect 40885 11275 40991 11381
rect 45050 11284 45158 11392
rect 36060 9206 36160 9306
rect 39009 9211 39099 9301
rect 35833 9025 35935 9127
rect 49822 7640 49824 7700
rect 49824 7640 49882 7700
rect 62350 7138 62352 7198
rect 62352 7138 62410 7198
rect 45916 6098 46016 6198
rect 49306 5676 49366 5736
rect 49940 5527 50000 5587
rect 8280 5144 8340 5204
rect 38915 3999 39015 4099
rect 43087 3997 43187 4097
rect 40785 3689 40895 3799
rect 45061 3677 45171 3787
rect 49302 3676 49306 3736
rect 49306 3676 49362 3736
rect 50082 3527 50142 3587
rect 46088 1610 46148 1670
rect 49828 1586 49884 1646
rect 49884 1586 49888 1646
rect 67277 18823 67367 18913
rect 66655 16327 66745 16417
rect 66026 4876 66086 4936
rect 62153 2843 62243 2933
rect 8042 522 8102 582
rect 3478 -90 34878 64
rect 57478 -90 88878 64
rect -1266 -576 -666 -276
rect 35166 -576 35766 -276
rect 52734 -576 53334 -276
rect 89166 -576 89766 -276
<< metal3 >>
rect 11424 28156 12044 28161
rect 11424 27856 11434 28156
rect 12034 27856 12044 28156
rect 11424 27851 12044 27856
rect 35056 28156 35676 28161
rect 35056 27856 35066 28156
rect 35666 27856 35676 28156
rect 35056 27851 35676 27856
rect 65424 28156 66044 28161
rect 65424 27856 65434 28156
rect 66034 27856 66044 28156
rect 65424 27851 66044 27856
rect 89056 28156 89676 28161
rect 89056 27856 89066 28156
rect 89666 27856 89676 28156
rect 89056 27851 89676 27856
rect 14948 27774 31828 27806
rect -1436 27647 -1330 27668
rect -1436 27583 -1419 27647
rect -1349 27583 -1330 27647
rect -1436 27582 -1414 27583
rect -1354 27582 -1330 27583
rect -1436 27562 -1330 27582
rect 14948 27560 15011 27774
rect 31796 27560 31828 27774
rect 68948 27774 85828 27806
rect 14948 27540 31828 27560
rect 47796 27680 48490 27702
rect 47796 27564 47824 27680
rect 48462 27564 48490 27680
rect 14948 27538 19302 27540
rect 47796 27536 48490 27564
rect 68948 27560 69011 27774
rect 85796 27560 85828 27774
rect 68948 27540 85828 27560
rect 68948 27538 73302 27540
rect -1328 27092 -629 27120
rect -1328 26548 -713 27092
rect -649 26548 -629 27092
rect -1328 26520 -629 26548
rect -334 27093 1965 27121
rect -334 26549 1881 27093
rect 1945 26549 1965 27093
rect -334 26521 1965 26549
rect 2266 27093 4565 27121
rect 2266 26549 4481 27093
rect 4545 26549 4565 27093
rect 2266 26521 4565 26549
rect 4866 27093 7165 27121
rect 4866 26549 7081 27093
rect 7145 26549 7165 27093
rect 4866 26521 7165 26549
rect 7466 27093 9765 27121
rect 7466 26549 9681 27093
rect 9745 26549 9765 27093
rect 7466 26521 9765 26549
rect 10066 27092 10765 27120
rect 10066 26548 10681 27092
rect 10745 26548 10765 27092
rect 52672 27092 53371 27120
rect 712 26220 812 26521
rect 3312 26220 3412 26521
rect 5912 26220 6012 26521
rect 8512 26220 8612 26521
rect 10066 26520 10765 26548
rect 38430 26568 38578 26574
rect 37160 26420 38430 26494
rect 41348 26568 41506 26574
rect 38578 26420 41348 26494
rect 37160 26410 41348 26420
rect 52672 26548 53287 27092
rect 53351 26548 53371 27092
rect 52672 26520 53371 26548
rect 53666 27093 55965 27121
rect 53666 26549 55881 27093
rect 55945 26549 55965 27093
rect 53666 26521 55965 26549
rect 56266 27093 58565 27121
rect 56266 26549 58481 27093
rect 58545 26549 58565 27093
rect 56266 26521 58565 26549
rect 58866 27093 61165 27121
rect 58866 26549 61081 27093
rect 61145 26549 61165 27093
rect 58866 26521 61165 26549
rect 61466 27093 63765 27121
rect 61466 26549 63681 27093
rect 63745 26549 63765 27093
rect 61466 26521 63765 26549
rect 64066 27092 64765 27120
rect 64066 26548 64681 27092
rect 64745 26548 64765 27092
rect 41506 26410 42865 26494
rect -1330 26192 -631 26220
rect -1330 24048 -715 26192
rect -651 25162 -631 26192
rect -333 26192 1966 26220
rect -333 25162 1882 26192
rect -651 25062 1882 25162
rect -651 24048 -631 25062
rect -1330 24020 -631 24048
rect -333 24048 1882 25062
rect 1946 25162 1966 26192
rect 2267 26192 4566 26220
rect 2267 25162 4482 26192
rect 1946 25062 4482 25162
rect 1946 24048 1966 25062
rect -333 24020 1966 24048
rect 2267 24048 4482 25062
rect 4546 25162 4566 26192
rect 4867 26192 7166 26220
rect 4867 25162 7082 26192
rect 4546 25062 7082 25162
rect 4546 24048 4566 25062
rect 2267 24020 4566 24048
rect 4867 24048 7082 25062
rect 7146 25162 7166 26192
rect 7467 26192 9766 26220
rect 7467 25162 9682 26192
rect 7146 25062 9682 25162
rect 7146 24048 7166 25062
rect 4867 24020 7166 24048
rect 7467 24048 9682 25062
rect 9746 25162 9766 26192
rect 10064 26192 10763 26220
rect 10064 25162 10679 26192
rect 9746 25062 10679 25162
rect 9746 24048 9766 25062
rect 7467 24020 9766 24048
rect 10064 24048 10679 25062
rect 10743 24048 10763 26192
rect 37160 25893 42865 26410
rect 54712 26220 54812 26521
rect 57312 26220 57412 26521
rect 59912 26220 60012 26521
rect 62512 26220 62612 26521
rect 64066 26520 64765 26548
rect 37160 25880 39750 25893
rect 40168 25880 42865 25893
rect 37160 24776 37761 25880
rect 37044 24644 37050 24776
rect 37182 24644 37761 24776
rect 10064 24020 10763 24048
rect -1330 23692 -631 23720
rect 712 23719 812 24020
rect 3312 23719 3412 24020
rect 5912 23719 6012 24020
rect 8512 23719 8612 24020
rect -1330 21548 -715 23692
rect -651 22662 -631 23692
rect -333 23691 1966 23719
rect -333 22662 1882 23691
rect -651 22562 1882 22662
rect -651 21548 -631 22562
rect -1330 21520 -631 21548
rect -333 21547 1882 22562
rect 1946 22662 1966 23691
rect 2267 23691 4566 23719
rect 2267 22662 4482 23691
rect 1946 22562 4482 22662
rect 1946 21547 1966 22562
rect -333 21519 1966 21547
rect 2267 21547 4482 22562
rect 4546 22662 4566 23691
rect 4867 23691 7166 23719
rect 4867 22662 7082 23691
rect 4546 22562 7082 22662
rect 4546 21547 4566 22562
rect 2267 21519 4566 21547
rect 4867 21547 7082 22562
rect 7146 22662 7166 23691
rect 7467 23691 9766 23719
rect 7467 22662 9682 23691
rect 7146 22562 9682 22662
rect 7146 21547 7166 22562
rect 4867 21519 7166 21547
rect 7467 21547 9682 22562
rect 9746 22662 9766 23691
rect 10064 23692 10763 23720
rect 10064 22662 10679 23692
rect 9746 22562 10679 22662
rect 9746 21547 9766 22562
rect 7467 21519 9766 21547
rect 10064 21548 10679 22562
rect 10743 21548 10763 23692
rect 36462 23470 36468 23570
rect 36568 23470 36574 23570
rect 10064 21520 10763 21548
rect -1330 21192 -631 21220
rect 712 21219 812 21519
rect 3312 21219 3412 21519
rect 5912 21219 6012 21519
rect 8512 21219 8612 21519
rect -1330 19048 -715 21192
rect -651 20162 -631 21192
rect -333 21191 1966 21219
rect -333 20162 1882 21191
rect -651 20062 1882 20162
rect -651 19048 -631 20062
rect -1330 19020 -631 19048
rect -333 19047 1882 20062
rect 1946 20162 1966 21191
rect 2267 21191 4566 21219
rect 2267 20162 4482 21191
rect 1946 20062 4482 20162
rect 1946 19047 1966 20062
rect -333 19019 1966 19047
rect 2267 19047 4482 20062
rect 4546 20162 4566 21191
rect 4867 21191 7166 21219
rect 4867 20162 7082 21191
rect 4546 20062 7082 20162
rect 4546 19047 4566 20062
rect 2267 19019 4566 19047
rect 4867 19047 7082 20062
rect 7146 20162 7166 21191
rect 7467 21191 9766 21219
rect 7467 20162 9682 21191
rect 7146 20062 9682 20162
rect 7146 19047 7166 20062
rect 4867 19019 7166 19047
rect 7467 19047 9682 20062
rect 9746 20162 9766 21191
rect 10064 21192 10763 21220
rect 10064 20162 10679 21192
rect 9746 20062 10679 20162
rect 9746 19047 9766 20062
rect 7467 19019 9766 19047
rect 10064 19048 10679 20062
rect 10743 19048 10763 21192
rect 36468 20168 36568 23470
rect 37160 22676 37761 24644
rect 38018 23861 39806 25612
rect 38018 23812 38879 23861
rect 38874 23781 38879 23812
rect 38959 23812 39806 23861
rect 40048 23870 41836 25612
rect 40048 23812 40402 23870
rect 38959 23781 38964 23812
rect 38874 23776 38964 23781
rect 40396 23770 40402 23812
rect 40502 23812 41836 23870
rect 42251 24768 42865 25880
rect 52670 26192 53369 26220
rect 42251 24632 42912 24768
rect 43048 24632 43054 24768
rect 48378 24664 51894 24688
rect 42251 23934 42865 24632
rect 48378 24604 48398 24664
rect 48458 24604 51894 24664
rect 48378 24588 51894 24604
rect 46576 24534 46676 24540
rect 46676 24515 47704 24534
rect 46676 24455 47624 24515
rect 47684 24455 47704 24515
rect 46676 24434 47704 24455
rect 46576 24428 46676 24434
rect 42251 23874 42790 23934
rect 42850 23874 42865 23934
rect 40502 23770 40508 23812
rect 40401 23769 40503 23770
rect 41563 23712 41661 23717
rect 42030 23712 42130 23718
rect 41562 23711 42030 23712
rect 41562 23613 41563 23711
rect 41661 23613 42030 23711
rect 41562 23612 42030 23613
rect 41563 23607 41661 23612
rect 42030 23606 42130 23612
rect 39492 23567 39592 23568
rect 39487 23512 39493 23567
rect 37070 22556 37076 22676
rect 37196 22556 37761 22676
rect 37160 21038 37761 22556
rect 38018 23469 39493 23512
rect 39591 23512 39597 23567
rect 40996 23527 41096 23532
rect 40996 23512 41001 23527
rect 39591 23469 39806 23512
rect 38018 21712 39806 23469
rect 40048 23437 41001 23512
rect 41091 23512 41096 23527
rect 41091 23437 41836 23512
rect 40048 21712 41836 23437
rect 42251 22658 42865 23874
rect 46404 22664 47952 22684
rect 42251 22518 42864 22658
rect 43004 22518 43010 22658
rect 46404 22604 47876 22664
rect 47936 22604 47952 22664
rect 46404 22584 47952 22604
rect 42251 21920 42865 22518
rect 42251 21860 42800 21920
rect 42860 21860 42865 21920
rect 40228 21419 40328 21712
rect 40223 21414 40333 21419
rect 40223 21314 40228 21414
rect 40328 21314 40333 21414
rect 40223 21309 40333 21314
rect 42251 21038 42865 21860
rect 46404 21381 46504 22584
rect 48640 22515 49860 22532
rect 48640 22455 48656 22515
rect 48716 22455 49860 22515
rect 48640 22432 49860 22455
rect 49760 21700 49860 22432
rect 49760 21594 49860 21600
rect 46399 21283 46405 21381
rect 46503 21283 46509 21381
rect 46404 21282 46504 21283
rect 51794 21066 51894 24588
rect 52670 24048 53285 26192
rect 53349 25162 53369 26192
rect 53667 26192 55966 26220
rect 53667 25162 55882 26192
rect 53349 25062 55882 25162
rect 53349 24048 53369 25062
rect 52670 24020 53369 24048
rect 53667 24048 55882 25062
rect 55946 25162 55966 26192
rect 56267 26192 58566 26220
rect 56267 25162 58482 26192
rect 55946 25062 58482 25162
rect 55946 24048 55966 25062
rect 53667 24020 55966 24048
rect 56267 24048 58482 25062
rect 58546 25162 58566 26192
rect 58867 26192 61166 26220
rect 58867 25162 61082 26192
rect 58546 25062 61082 25162
rect 58546 24048 58566 25062
rect 56267 24020 58566 24048
rect 58867 24048 61082 25062
rect 61146 25162 61166 26192
rect 61467 26192 63766 26220
rect 61467 25162 63682 26192
rect 61146 25062 63682 25162
rect 61146 24048 61166 25062
rect 58867 24020 61166 24048
rect 61467 24048 63682 25062
rect 63746 25162 63766 26192
rect 64064 26192 64763 26220
rect 64064 25162 64679 26192
rect 63746 25062 64679 25162
rect 63746 24048 63766 25062
rect 61467 24020 63766 24048
rect 64064 24048 64679 25062
rect 64743 24048 64763 26192
rect 64064 24020 64763 24048
rect 52138 23614 52144 23714
rect 52244 23614 52250 23714
rect 52670 23692 53369 23720
rect 54712 23719 54812 24020
rect 57312 23719 57412 24020
rect 59912 23719 60012 24020
rect 62512 23719 62612 24020
rect 37160 20490 51393 21038
rect 51788 20966 51794 21066
rect 51894 20966 51900 21066
rect 37160 20437 38494 20490
rect 37279 20420 38494 20437
rect 36468 19925 36572 20168
rect 36467 19827 36473 19925
rect 36571 19827 36577 19925
rect 10064 19020 10763 19048
rect -1330 18692 -631 18720
rect 712 18719 812 19019
rect 3312 18719 3412 19019
rect 5912 18719 6012 19019
rect 8512 18719 8612 19019
rect 9201 18918 9299 18923
rect 9200 18917 13372 18918
rect 9200 18819 9201 18917
rect 9299 18913 13372 18917
rect 9299 18823 11211 18913
rect 11301 18823 13277 18913
rect 13367 18823 13372 18913
rect 9299 18819 13372 18823
rect 9200 18818 13372 18819
rect 9201 18813 9299 18818
rect -1330 16548 -715 18692
rect -651 17662 -631 18692
rect -333 18691 1966 18719
rect -333 17662 1882 18691
rect -651 17562 1882 17662
rect -651 16548 -631 17562
rect -1330 16520 -631 16548
rect -333 16547 1882 17562
rect 1946 17662 1966 18691
rect 2267 18691 4566 18719
rect 2267 17662 4482 18691
rect 1946 17562 4482 17662
rect 1946 16547 1966 17562
rect -333 16519 1966 16547
rect 2267 16547 4482 17562
rect 4546 17662 4566 18691
rect 4867 18691 7166 18719
rect 4867 17662 7082 18691
rect 4546 17562 7082 17662
rect 4546 16547 4566 17562
rect 2267 16519 4566 16547
rect 4867 16547 7082 17562
rect 7146 17662 7166 18691
rect 7467 18691 9766 18719
rect 7467 17662 9682 18691
rect 7146 17562 9682 17662
rect 7146 16547 7166 17562
rect 4867 16519 7166 16547
rect 7467 16547 9682 17562
rect 9746 17662 9766 18691
rect 10064 18692 10763 18720
rect 10064 17662 10679 18692
rect 9746 17562 10679 17662
rect 9746 16547 9766 17562
rect 7467 16519 9766 16547
rect 10064 16548 10679 17562
rect 10743 16548 10763 18692
rect 36468 17152 36572 19827
rect 37279 19649 37879 20420
rect 38672 20420 40894 20490
rect 38494 20306 38672 20312
rect 41072 20420 43294 20490
rect 40894 20306 41072 20312
rect 43472 20420 45420 20490
rect 43294 20306 43472 20312
rect 45598 20420 47594 20490
rect 45420 20306 45598 20312
rect 47772 20420 49994 20490
rect 47594 20306 47772 20312
rect 50172 20420 51393 20490
rect 49994 20306 50172 20312
rect 39072 19826 39078 19926
rect 39178 19826 46764 19926
rect 37279 18790 37881 19649
rect 39682 19574 39782 19826
rect 42460 19574 42560 19826
rect 46664 19574 46764 19826
rect 37144 18582 37150 18790
rect 37358 18582 37881 18790
rect 36468 17048 36852 17152
rect 10064 16520 10763 16548
rect -1332 16194 -633 16222
rect 712 16221 812 16519
rect 3312 16221 3412 16519
rect 5912 16221 6012 16519
rect 8512 16221 8612 16519
rect 9861 16422 9959 16427
rect 10957 16422 11067 16423
rect 9860 16421 36558 16422
rect 9860 16323 9861 16421
rect 9959 16418 36558 16421
rect 9959 16323 10962 16418
rect 9860 16322 10962 16323
rect 9861 16317 9959 16322
rect 10957 16318 10962 16322
rect 11062 16417 36558 16418
rect 11062 16327 12655 16417
rect 12745 16327 36558 16417
rect 11062 16322 36558 16327
rect 11062 16318 11067 16322
rect 10957 16313 11067 16318
rect -1332 15650 -717 16194
rect -653 15650 -633 16194
rect -1332 15622 -633 15650
rect -334 16193 1965 16221
rect -334 15649 1881 16193
rect 1945 15649 1965 16193
rect -13304 15385 -13204 15396
rect -13304 15325 -13286 15385
rect -13226 15325 -13204 15385
rect -13304 14732 -13204 15325
rect -10642 15385 -10542 15410
rect -10642 15325 -10620 15385
rect -10560 15325 -10542 15385
rect -10642 14732 -10542 15325
rect -1082 15357 -982 15622
rect -334 15621 1965 15649
rect 2266 16193 4565 16221
rect 2266 15649 4481 16193
rect 4545 15649 4565 16193
rect 2266 15621 4565 15649
rect 4866 16193 7165 16221
rect 4866 15649 7081 16193
rect 7145 15649 7165 16193
rect 4866 15621 7165 15649
rect 7466 16193 9765 16221
rect 7466 15649 9681 16193
rect 9745 15649 9765 16193
rect 7466 15621 9765 15649
rect 10066 16194 10765 16222
rect 10066 15650 10681 16194
rect 10745 15650 10765 16194
rect 36254 16193 36354 16198
rect 36254 16103 36259 16193
rect 36349 16103 36354 16193
rect 11201 15882 11311 15887
rect 11201 15782 11206 15882
rect 11306 15782 36158 15882
rect 11201 15777 11311 15782
rect 10066 15622 10765 15650
rect -1082 15267 -1077 15357
rect -987 15267 -982 15357
rect -1082 15262 -982 15267
rect 712 15357 812 15621
rect 712 15267 717 15357
rect 807 15267 812 15357
rect 712 15262 812 15267
rect 3312 15357 3412 15621
rect 3312 15267 3317 15357
rect 3407 15267 3412 15357
rect 3312 15262 3412 15267
rect 5912 15359 6012 15621
rect 5912 15269 5917 15359
rect 6007 15269 6012 15359
rect 5912 15264 6012 15269
rect 8512 15359 8612 15621
rect 8512 15269 8517 15359
rect 8607 15269 8612 15359
rect 8512 15264 8612 15269
rect 10316 15359 10416 15622
rect 10316 15269 10321 15359
rect 10411 15269 10416 15359
rect 10316 15264 10416 15269
rect -1950 15152 35940 15182
rect -1950 15092 -1924 15152
rect -1864 15092 35940 15152
rect -1950 15070 35940 15092
rect -13304 14632 -10542 14732
rect -2396 14983 11062 14988
rect -2396 14893 10967 14983
rect 11057 14893 11062 14983
rect -2396 14888 11062 14893
rect -13472 14605 -13372 14610
rect -13472 14515 -13467 14605
rect -13377 14515 -13372 14605
rect -13472 10731 -13372 14515
rect -13477 10633 -13471 10731
rect -13373 10633 -13367 10731
rect -13472 10632 -13372 10633
rect -13304 3537 -13204 14632
rect -8836 14174 -8646 14180
rect -11154 14168 -11008 14174
rect -11154 14002 -11008 14022
rect -12476 13984 -8836 14002
rect -3940 14168 -3782 14174
rect -6346 14150 -6170 14156
rect -8646 13984 -6346 14002
rect -12476 13974 -6346 13984
rect -3940 14002 -3782 14010
rect -6170 13974 -2606 14002
rect -12476 13400 -2606 13974
rect -12476 13398 -7666 13400
rect -13108 13137 -13008 13138
rect -13113 13039 -13107 13137
rect -13009 13039 -13003 13137
rect -13108 12772 -13006 13039
rect -13106 9154 -13006 12772
rect -12476 11974 -11875 13398
rect -10580 13038 -10574 13138
rect -10474 13120 -7214 13138
rect -10474 13060 -9878 13120
rect -9818 13060 -7214 13120
rect -10474 13038 -7214 13060
rect -9994 12784 -9894 13038
rect -7314 12784 -7214 13038
rect -12630 11880 -12624 11974
rect -12530 11880 -11875 11974
rect -12476 10010 -11875 11880
rect -11628 11043 -9840 12784
rect -11628 10984 -9955 11043
rect -9960 10939 -9955 10984
rect -9851 10984 -9840 11043
rect -9598 11029 -7810 12784
rect -9598 10984 -9225 11029
rect -9851 10939 -9846 10984
rect -9960 10934 -9846 10939
rect -9231 10931 -9225 10984
rect -9127 10984 -7810 11029
rect -7438 11027 -5650 12784
rect -7438 10984 -5821 11027
rect -9127 10931 -9121 10984
rect -5826 10931 -5821 10984
rect -5725 10984 -5650 11027
rect -5398 11029 -3610 12784
rect -5398 10984 -5269 11029
rect -5725 10931 -5720 10984
rect -5275 10931 -5269 10984
rect -5171 10984 -3610 11029
rect -3207 12166 -2606 13400
rect -2396 12904 -2296 14888
rect 11201 14812 11311 14817
rect 10974 14810 11206 14812
rect -1756 14712 11206 14810
rect 11306 14712 11311 14812
rect -1756 14710 11311 14712
rect -2402 12804 -2396 12904
rect -2296 12804 -2290 12904
rect -3207 11856 -2604 12166
rect -3207 11764 -2524 11856
rect -2432 11764 -2426 11856
rect -3207 11566 -2604 11764
rect -5171 10931 -5165 10984
rect -9226 10930 -9126 10931
rect -5826 10926 -5720 10931
rect -5270 10930 -5170 10931
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10881 -7570 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -7570 10881
rect -8102 10782 -7570 10783
rect -3901 10880 -3803 10885
rect -3392 10880 -3292 10886
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -3902 10879 -3392 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3392 10879
rect -3902 10780 -3392 10781
rect -3292 10780 -3288 10880
rect -3901 10775 -3803 10780
rect -3392 10774 -3292 10780
rect -6556 10733 -6456 10734
rect -10356 10731 -10256 10732
rect -10361 10684 -10355 10731
rect -12640 9930 -12634 10010
rect -12554 9930 -11875 10010
rect -13106 9054 -12632 9154
rect -13100 8619 -13000 8620
rect -13105 8521 -13099 8619
rect -13001 8521 -12995 8619
rect -13309 3439 -13303 3537
rect -13205 3439 -13199 3537
rect -13304 3438 -13204 3439
rect -13100 1627 -13000 8521
rect -12732 5665 -12632 9054
rect -12476 8262 -11875 9930
rect -11628 10633 -10355 10684
rect -10257 10684 -10251 10731
rect -8786 10725 -8662 10730
rect -8786 10684 -8781 10725
rect -10257 10633 -9840 10684
rect -11628 8884 -9840 10633
rect -9598 10611 -8781 10684
rect -8667 10684 -8662 10725
rect -6561 10684 -6555 10733
rect -8667 10611 -7810 10684
rect -9598 8884 -7810 10611
rect -7438 10635 -6555 10684
rect -6457 10684 -6451 10733
rect -4794 10715 -4678 10720
rect -4794 10684 -4789 10715
rect -6457 10635 -5650 10684
rect -7438 8884 -5650 10635
rect -5398 10609 -4789 10684
rect -4683 10684 -4678 10715
rect -4683 10609 -3610 10684
rect -5398 8884 -3610 10609
rect -3207 9848 -2606 11566
rect -1756 11018 -1656 14710
rect 11201 14707 11311 14710
rect -3207 9742 -2518 9848
rect -2412 9742 -2406 9848
rect -10132 8620 -10032 8884
rect -7192 8620 -7092 8884
rect -10540 8520 -10534 8620
rect -10434 8520 -7092 8620
rect -3207 8264 -2606 9742
rect -1758 8863 -1656 11018
rect 35828 9127 35940 15070
rect 36058 9716 36158 15782
rect 36254 15375 36354 16103
rect 36249 15277 36255 15375
rect 36353 15277 36359 15375
rect 35828 9025 35833 9127
rect 35935 9025 35940 9127
rect 35828 9020 35940 9025
rect 36054 9311 36158 9716
rect 36254 9541 36354 15277
rect 36458 13819 36558 16322
rect 36451 13814 36561 13819
rect 36451 13714 36456 13814
rect 36556 13714 36561 13814
rect 36451 13709 36561 13714
rect 36249 9443 36255 9541
rect 36353 9443 36359 9541
rect 36254 9442 36354 9443
rect 36054 9306 36165 9311
rect 36054 9206 36060 9306
rect 36160 9206 36165 9306
rect 36054 9201 36165 9206
rect -1761 8765 -1755 8863
rect -1657 8765 -1651 8863
rect -7140 8262 -2606 8264
rect -12476 7662 -2606 8262
rect 35229 7738 35327 7743
rect 11362 7737 35328 7738
rect -12476 7660 -6020 7662
rect -4183 7660 -3581 7662
rect -11204 7646 -10950 7660
rect -11204 7406 -11197 7646
rect -10957 7556 -10950 7646
rect -8792 7646 -8538 7660
rect -10957 7406 -10951 7556
rect -8792 7406 -8785 7646
rect -8545 7556 -8538 7646
rect -6380 7646 -6126 7660
rect -8545 7406 -8539 7556
rect -6380 7406 -6373 7646
rect -6133 7556 -6126 7646
rect -3968 7646 -3714 7660
rect -6133 7406 -6127 7556
rect -3968 7406 -3961 7646
rect -3721 7556 -3714 7646
rect 11362 7639 35229 7737
rect 35327 7639 35328 7737
rect 11362 7638 35328 7639
rect -3721 7406 -3715 7556
rect -11204 7056 -10954 7406
rect -11204 6814 -11198 7056
rect -10956 6814 -10954 7056
rect -11204 6812 -10954 6814
rect -8792 7056 -8542 7406
rect -8792 6814 -8786 7056
rect -8544 6814 -8542 7056
rect -8792 6812 -8542 6814
rect -6380 7056 -6130 7406
rect -6380 6814 -6374 7056
rect -6132 6814 -6130 7056
rect -6380 6812 -6130 6814
rect -3968 7056 -3718 7406
rect 11362 7198 11462 7638
rect 35229 7633 35327 7638
rect 11362 7138 11382 7198
rect 11442 7138 11462 7198
rect 11362 7102 11462 7138
rect -3968 6814 -3962 7056
rect -3720 6814 -3718 7056
rect -3968 6812 -3718 6814
rect -12474 6798 -2604 6812
rect -12475 6712 -2604 6798
rect -12475 6198 -2607 6712
rect -12737 5567 -12731 5665
rect -12633 5567 -12627 5665
rect -12732 5566 -12632 5567
rect -12475 4766 -11875 6198
rect -9948 5852 -7198 5952
rect -9948 5584 -9848 5852
rect -7298 5584 -7198 5852
rect -12592 4616 -12586 4766
rect -12436 4616 -11875 4766
rect -12475 2650 -11875 4616
rect -11628 3835 -9840 5584
rect -11628 3784 -10815 3835
rect -10820 3741 -10815 3784
rect -10721 3784 -9840 3835
rect -9598 3827 -7810 5584
rect -9598 3784 -9365 3827
rect -10721 3741 -10716 3784
rect -10820 3736 -10716 3741
rect -9371 3729 -9365 3784
rect -9267 3784 -7810 3827
rect -7438 3827 -5650 5584
rect -7438 3784 -6737 3827
rect -9267 3729 -9261 3784
rect -6742 3737 -6737 3784
rect -6647 3784 -5650 3827
rect -5398 3839 -3610 5584
rect -5398 3784 -5143 3839
rect -6647 3737 -6642 3784
rect -6742 3732 -6642 3737
rect -9366 3728 -9266 3729
rect -5149 3725 -5143 3784
rect -5029 3784 -3610 3839
rect -3207 4716 -2607 6198
rect -2426 5665 -2322 5666
rect -2427 5567 -2421 5665
rect -2323 5567 -2317 5665
rect -2426 5228 -2322 5567
rect -2426 5226 8314 5228
rect -2426 5204 8366 5226
rect -2426 5144 8280 5204
rect 8340 5144 8366 5204
rect -2426 5126 8366 5144
rect -2426 5124 8314 5126
rect -3207 4562 -2660 4716
rect -2506 4562 -2500 4716
rect -5029 3725 -5023 3784
rect -5144 3724 -5028 3725
rect -8085 3682 -7987 3687
rect -7554 3682 -7454 3688
rect -3885 3684 -3787 3689
rect -3382 3684 -3282 3690
rect -8086 3681 -7554 3682
rect -8086 3583 -8085 3681
rect -7987 3583 -7554 3681
rect -8086 3582 -7554 3583
rect -3886 3683 -3382 3684
rect -3886 3585 -3885 3683
rect -3787 3585 -3382 3683
rect -3886 3584 -3382 3585
rect -8085 3577 -7987 3582
rect -7554 3576 -7454 3582
rect -3885 3579 -3787 3584
rect -3382 3578 -3282 3584
rect -10168 3537 -10068 3538
rect -10173 3484 -10167 3537
rect -12586 2524 -12580 2650
rect -12454 2524 -11875 2650
rect -13103 1529 -13097 1627
rect -12999 1529 -12993 1627
rect -13100 1528 -13000 1529
rect -12475 1062 -11875 2524
rect -11628 3439 -10167 3484
rect -10069 3484 -10063 3537
rect -9015 3514 -8901 3519
rect -9015 3484 -9010 3514
rect -10069 3439 -9840 3484
rect -11628 1684 -9840 3439
rect -9598 3410 -9010 3484
rect -8906 3484 -8901 3514
rect -5914 3484 -5908 3542
rect -8906 3410 -7810 3484
rect -9598 1684 -7810 3410
rect -7438 3426 -5908 3484
rect -5792 3484 -5786 3542
rect -4641 3510 -4531 3515
rect -4641 3484 -4636 3510
rect -5792 3426 -5650 3484
rect -7438 1684 -5650 3426
rect -5398 3410 -4636 3484
rect -4536 3484 -4531 3510
rect -4536 3410 -3610 3484
rect -5398 1684 -3610 3410
rect -3207 3060 -2607 4562
rect -3207 2664 -2608 3060
rect -3207 2504 -2666 2664
rect -2506 2504 -2500 2664
rect -3207 2202 -2608 2504
rect 36054 2238 36158 9201
rect 36458 6197 36558 13709
rect 36748 13581 36852 17048
rect 37279 16650 37881 18582
rect 38126 17829 39914 19574
rect 38126 17774 38973 17829
rect 38968 17731 38973 17774
rect 39071 17774 39914 17829
rect 40156 17829 41944 19574
rect 40156 17774 40417 17829
rect 39071 17731 39076 17774
rect 40411 17731 40417 17774
rect 40515 17774 41944 17829
rect 42316 17841 44104 19574
rect 42316 17774 43139 17841
rect 40515 17731 40521 17774
rect 38968 17726 39076 17731
rect 40416 17730 40516 17731
rect 43134 17723 43139 17774
rect 43257 17774 44104 17841
rect 44356 17817 46144 19574
rect 44356 17774 44643 17817
rect 43257 17723 43262 17774
rect 43134 17718 43262 17723
rect 44637 17719 44643 17774
rect 44741 17774 46144 17817
rect 46512 17831 48300 19574
rect 46512 17774 47331 17831
rect 44741 17719 44747 17774
rect 47326 17731 47331 17774
rect 47431 17774 48300 17831
rect 48552 17827 50340 19574
rect 48552 17774 48765 17827
rect 47431 17731 47436 17774
rect 47326 17726 47436 17731
rect 48759 17729 48765 17774
rect 48863 17774 50340 17827
rect 50792 18732 51393 20420
rect 50792 18570 51338 18732
rect 51500 18570 51506 18732
rect 48863 17729 48869 17774
rect 48764 17728 48864 17729
rect 44642 17718 44742 17719
rect 41673 17678 41771 17683
rect 42204 17678 42304 17684
rect 45873 17678 45971 17683
rect 46404 17678 46504 17684
rect 50073 17678 50171 17683
rect 50604 17678 50704 17684
rect 41672 17677 42204 17678
rect 41672 17579 41673 17677
rect 41771 17579 42204 17677
rect 41672 17578 42204 17579
rect 45872 17677 46404 17678
rect 45872 17579 45873 17677
rect 45971 17579 46404 17677
rect 45872 17578 46404 17579
rect 50072 17677 50604 17678
rect 50072 17579 50073 17677
rect 50171 17579 50604 17677
rect 50072 17578 50604 17579
rect 41673 17573 41771 17578
rect 42204 17572 42304 17578
rect 45873 17573 45971 17578
rect 46404 17572 46504 17578
rect 50073 17573 50171 17578
rect 50604 17572 50704 17578
rect 45183 17526 45321 17531
rect 39618 17523 39718 17524
rect 43818 17523 43918 17524
rect 39613 17474 39619 17523
rect 37073 16464 37079 16650
rect 37265 16464 37881 16650
rect 37279 14870 37881 16464
rect 38126 17425 39619 17474
rect 39717 17474 39723 17523
rect 40989 17516 41107 17521
rect 40989 17474 40994 17516
rect 39717 17425 39914 17474
rect 38126 15674 39914 17425
rect 40156 17408 40994 17474
rect 41102 17474 41107 17516
rect 43813 17474 43819 17523
rect 41102 17408 41944 17474
rect 40156 15674 41944 17408
rect 42316 17425 43819 17474
rect 43917 17474 43923 17523
rect 45183 17474 45188 17526
rect 43917 17425 44104 17474
rect 42316 15674 44104 17425
rect 44356 17398 45188 17474
rect 45316 17474 45321 17526
rect 48018 17521 48118 17522
rect 48013 17474 48019 17521
rect 45316 17398 46144 17474
rect 44356 15674 46144 17398
rect 46512 17423 48019 17474
rect 48117 17474 48123 17521
rect 49278 17507 49398 17512
rect 49278 17474 49283 17507
rect 48117 17423 48300 17474
rect 46512 15674 48300 17423
rect 48552 17397 49283 17474
rect 49393 17474 49398 17507
rect 49393 17397 50340 17474
rect 48552 15674 50340 17397
rect 50792 16638 51393 18570
rect 50792 16470 51364 16638
rect 51532 16470 51538 16638
rect 39672 15376 39772 15674
rect 42582 15376 42682 15674
rect 46660 15376 46760 15674
rect 39292 15276 39298 15376
rect 39398 15276 46760 15376
rect 50792 14870 51393 16470
rect 37131 14316 51393 14870
rect 52144 14738 52244 23614
rect 52670 21548 53285 23692
rect 53349 22662 53369 23692
rect 53667 23691 55966 23719
rect 53667 22662 55882 23691
rect 53349 22562 55882 22662
rect 53349 21548 53369 22562
rect 52670 21520 53369 21548
rect 53667 21547 55882 22562
rect 55946 22662 55966 23691
rect 56267 23691 58566 23719
rect 56267 22662 58482 23691
rect 55946 22562 58482 22662
rect 55946 21547 55966 22562
rect 53667 21519 55966 21547
rect 56267 21547 58482 22562
rect 58546 22662 58566 23691
rect 58867 23691 61166 23719
rect 58867 22662 61082 23691
rect 58546 22562 61082 22662
rect 58546 21547 58566 22562
rect 56267 21519 58566 21547
rect 58867 21547 61082 22562
rect 61146 22662 61166 23691
rect 61467 23691 63766 23719
rect 61467 22662 63682 23691
rect 61146 22562 63682 22662
rect 61146 21547 61166 22562
rect 58867 21519 61166 21547
rect 61467 21547 63682 22562
rect 63746 22662 63766 23691
rect 64064 23692 64763 23720
rect 64064 22662 64679 23692
rect 63746 22562 64679 22662
rect 63746 21547 63766 22562
rect 61467 21519 63766 21547
rect 64064 21548 64679 22562
rect 64743 21548 64763 23692
rect 64064 21520 64763 21548
rect 52670 21192 53369 21220
rect 54712 21219 54812 21519
rect 57312 21219 57412 21519
rect 59912 21219 60012 21519
rect 62512 21219 62612 21519
rect 52670 19048 53285 21192
rect 53349 20162 53369 21192
rect 53667 21191 55966 21219
rect 53667 20162 55882 21191
rect 53349 20062 55882 20162
rect 53349 19048 53369 20062
rect 52670 19020 53369 19048
rect 53667 19047 55882 20062
rect 55946 20162 55966 21191
rect 56267 21191 58566 21219
rect 56267 20162 58482 21191
rect 55946 20062 58482 20162
rect 55946 19047 55966 20062
rect 53667 19019 55966 19047
rect 56267 19047 58482 20062
rect 58546 20162 58566 21191
rect 58867 21191 61166 21219
rect 58867 20162 61082 21191
rect 58546 20062 61082 20162
rect 58546 19047 58566 20062
rect 56267 19019 58566 19047
rect 58867 19047 61082 20062
rect 61146 20162 61166 21191
rect 61467 21191 63766 21219
rect 61467 20162 63682 21191
rect 61146 20062 63682 20162
rect 61146 19047 61166 20062
rect 58867 19019 61166 19047
rect 61467 19047 63682 20062
rect 63746 20162 63766 21191
rect 64064 21192 64763 21220
rect 64064 20162 64679 21192
rect 63746 20062 64679 20162
rect 63746 19047 63766 20062
rect 61467 19019 63766 19047
rect 64064 19048 64679 20062
rect 64743 19048 64763 21192
rect 64064 19020 64763 19048
rect 52670 18692 53369 18720
rect 54712 18719 54812 19019
rect 57312 18719 57412 19019
rect 59912 18719 60012 19019
rect 62512 18719 62612 19019
rect 63201 18918 63299 18923
rect 63200 18917 67372 18918
rect 63200 18819 63201 18917
rect 63299 18913 67372 18917
rect 63299 18823 65093 18913
rect 65183 18823 67277 18913
rect 67367 18823 67372 18913
rect 63299 18819 67372 18823
rect 63200 18818 67372 18819
rect 63201 18813 63299 18818
rect 52670 16548 53285 18692
rect 53349 17662 53369 18692
rect 53667 18691 55966 18719
rect 53667 17662 55882 18691
rect 53349 17562 55882 17662
rect 53349 16548 53369 17562
rect 52670 16520 53369 16548
rect 53667 16547 55882 17562
rect 55946 17662 55966 18691
rect 56267 18691 58566 18719
rect 56267 17662 58482 18691
rect 55946 17562 58482 17662
rect 55946 16547 55966 17562
rect 53667 16519 55966 16547
rect 56267 16547 58482 17562
rect 58546 17662 58566 18691
rect 58867 18691 61166 18719
rect 58867 17662 61082 18691
rect 58546 17562 61082 17662
rect 58546 16547 58566 17562
rect 56267 16519 58566 16547
rect 58867 16547 61082 17562
rect 61146 17662 61166 18691
rect 61467 18691 63766 18719
rect 61467 17662 63682 18691
rect 61146 17562 63682 17662
rect 61146 16547 61166 17562
rect 58867 16519 61166 16547
rect 61467 16547 63682 17562
rect 63746 17662 63766 18691
rect 64064 18692 64763 18720
rect 64064 17662 64679 18692
rect 63746 17562 64679 17662
rect 63746 16547 63766 17562
rect 61467 16519 63766 16547
rect 64064 16548 64679 17562
rect 64743 16548 64763 18692
rect 64064 16520 64763 16548
rect 52668 16194 53367 16222
rect 54712 16221 54812 16519
rect 57312 16221 57412 16519
rect 59912 16221 60012 16519
rect 62512 16221 62612 16519
rect 63861 16422 63959 16427
rect 63860 16421 66750 16422
rect 63860 16323 63861 16421
rect 63959 16417 66750 16421
rect 63959 16327 66655 16417
rect 66745 16327 66750 16417
rect 63959 16323 66750 16327
rect 63860 16322 66750 16323
rect 63861 16317 63959 16322
rect 52668 15650 53283 16194
rect 53347 15650 53367 16194
rect 52668 15622 53367 15650
rect 53666 16193 55965 16221
rect 53666 15649 55881 16193
rect 55945 15649 55965 16193
rect 52918 15357 53018 15622
rect 53666 15621 55965 15649
rect 56266 16193 58565 16221
rect 56266 15649 58481 16193
rect 58545 15649 58565 16193
rect 56266 15621 58565 15649
rect 58866 16193 61165 16221
rect 58866 15649 61081 16193
rect 61145 15649 61165 16193
rect 58866 15621 61165 15649
rect 61466 16193 63765 16221
rect 61466 15649 63681 16193
rect 63745 15649 63765 16193
rect 61466 15621 63765 15649
rect 64066 16194 64765 16222
rect 64066 15650 64681 16194
rect 64745 15650 64765 16194
rect 64066 15622 64765 15650
rect 52918 15267 52923 15357
rect 53013 15267 53018 15357
rect 52918 15262 53018 15267
rect 54712 15357 54812 15621
rect 54712 15267 54717 15357
rect 54807 15267 54812 15357
rect 54712 15262 54812 15267
rect 57312 15357 57412 15621
rect 57312 15267 57317 15357
rect 57407 15267 57412 15357
rect 57312 15262 57412 15267
rect 59912 15359 60012 15621
rect 59912 15269 59917 15359
rect 60007 15269 60012 15359
rect 59912 15264 60012 15269
rect 62512 15359 62612 15621
rect 62512 15269 62517 15359
rect 62607 15269 62612 15359
rect 62512 15264 62612 15269
rect 64316 15359 64416 15622
rect 64316 15269 64321 15359
rect 64411 15269 64416 15359
rect 64316 15264 64416 15269
rect 52380 15100 52480 15106
rect 64976 15100 65076 16322
rect 52480 15000 65076 15100
rect 52380 14994 52480 15000
rect 65083 14738 65193 14743
rect 52144 14638 65088 14738
rect 65188 14638 65193 14738
rect 65083 14633 65193 14638
rect 37131 14260 38478 14316
rect 36743 13483 36749 13581
rect 36847 13483 36853 13581
rect 37131 13527 37731 14260
rect 38636 14260 40890 14316
rect 38478 14152 38636 14158
rect 41048 14260 43290 14316
rect 40890 14152 41048 14158
rect 43448 14260 45690 14316
rect 43290 14152 43448 14158
rect 45848 14268 47690 14316
rect 45848 14260 46992 14268
rect 45690 14152 45848 14158
rect 39248 13809 42430 13814
rect 39248 13719 39253 13809
rect 39343 13719 42430 13809
rect 39248 13714 42430 13719
rect 36748 13480 36852 13483
rect 37131 12668 37733 13527
rect 39568 13452 39668 13714
rect 42330 13452 42430 13714
rect 46399 13454 46992 14260
rect 47848 14268 50090 14316
rect 47690 14152 47848 14158
rect 50248 14268 51393 14316
rect 50792 14264 51393 14268
rect 50090 14152 50248 14158
rect 36996 12460 37002 12668
rect 37210 12460 37733 12668
rect 37131 10528 37733 12460
rect 37978 11711 39766 13452
rect 37978 11652 38849 11711
rect 38844 11615 38849 11652
rect 38945 11652 39766 11711
rect 40008 11709 41796 13452
rect 40008 11652 40293 11709
rect 38945 11615 38950 11652
rect 38844 11610 38950 11615
rect 40287 11611 40293 11652
rect 40391 11652 41796 11709
rect 42168 11727 43956 13452
rect 42168 11652 42999 11727
rect 40391 11611 40397 11652
rect 40292 11610 40392 11611
rect 42994 11597 42999 11652
rect 43125 11652 43956 11727
rect 44208 11709 45996 13452
rect 44208 11652 44513 11709
rect 43125 11597 43130 11652
rect 44507 11611 44513 11652
rect 44611 11652 45996 11709
rect 46399 12734 46998 13454
rect 46399 12610 46999 12734
rect 46399 12448 47030 12610
rect 47192 12448 47198 12610
rect 46399 12380 46999 12448
rect 46399 11654 46998 12380
rect 44611 11611 44617 11652
rect 44512 11610 44612 11611
rect 42994 11592 43130 11597
rect 41543 11560 41641 11565
rect 42074 11560 42174 11566
rect 45743 11560 45841 11565
rect 46218 11560 46318 11566
rect 41542 11559 42074 11560
rect 41542 11461 41543 11559
rect 41641 11461 42074 11559
rect 41542 11460 42074 11461
rect 45742 11559 46218 11560
rect 45742 11461 45743 11559
rect 45841 11461 46218 11559
rect 45742 11460 46218 11461
rect 41543 11455 41641 11460
rect 42074 11454 42174 11460
rect 45743 11455 45841 11460
rect 46218 11454 46318 11460
rect 39488 11411 39588 11412
rect 39483 11352 39489 11411
rect 36925 10342 36931 10528
rect 37117 10342 37733 10528
rect 37131 8932 37733 10342
rect 37978 11313 39489 11352
rect 39587 11352 39593 11411
rect 43688 11393 43788 11394
rect 40880 11381 40996 11386
rect 40880 11352 40885 11381
rect 39587 11313 39766 11352
rect 37978 9552 39766 11313
rect 40008 11275 40885 11352
rect 40991 11352 40996 11381
rect 43683 11352 43689 11393
rect 40991 11275 41796 11352
rect 40008 9552 41796 11275
rect 42168 11295 43689 11352
rect 43787 11352 43793 11393
rect 45045 11392 45163 11397
rect 45045 11352 45050 11392
rect 43787 11295 43956 11352
rect 42168 9552 43956 11295
rect 44208 11284 45050 11352
rect 45158 11352 45163 11392
rect 45158 11284 45996 11352
rect 44208 9552 45996 11284
rect 46399 11350 46992 11654
rect 46399 10634 46998 11350
rect 46399 10510 46999 10634
rect 46399 10342 46992 10510
rect 47160 10342 47166 10510
rect 46399 9958 46999 10342
rect 39542 9306 39642 9552
rect 42452 9306 42552 9552
rect 39004 9301 42552 9306
rect 39004 9211 39009 9301
rect 39099 9211 42552 9301
rect 39004 9206 42552 9211
rect 46399 9218 47037 9958
rect 46399 8932 46999 9218
rect 37131 8400 46999 8932
rect 37131 8330 38476 8400
rect 37131 8328 37731 8330
rect 38704 8398 46999 8400
rect 38704 8328 40888 8398
rect 40886 8312 40888 8328
rect 38476 8166 38704 8172
rect 41116 8328 43232 8398
rect 43230 8312 43232 8328
rect 40888 8164 41116 8170
rect 43460 8330 45620 8398
rect 43460 8328 44542 8330
rect 43232 8164 43460 8170
rect 45848 8332 46999 8398
rect 45848 8330 46992 8332
rect 45848 8310 45850 8330
rect 45620 8164 45848 8170
rect 36990 7638 36996 7738
rect 37096 7638 47596 7738
rect 53050 7722 53150 7728
rect 47496 7222 47596 7638
rect 49800 7700 53050 7722
rect 49800 7640 49822 7700
rect 49882 7640 53050 7700
rect 49800 7622 53050 7640
rect 53050 7616 53150 7622
rect 47494 7198 62432 7222
rect 38428 7174 38610 7180
rect 37150 7064 38428 7078
rect 37149 6992 38428 7064
rect 40828 7174 41010 7180
rect 38610 6992 40828 7078
rect 43240 7174 43422 7180
rect 41010 6992 43240 7078
rect 45640 7174 45822 7180
rect 43422 6992 45640 7078
rect 47494 7138 62350 7198
rect 62410 7138 62432 7198
rect 47494 7122 62432 7138
rect 45822 6992 47017 7078
rect 37149 6464 47017 6992
rect 36453 6099 36459 6197
rect 36557 6099 36563 6197
rect 36458 6098 36558 6099
rect 37149 5066 37749 6464
rect 45911 6198 46021 6203
rect 39048 6098 39054 6198
rect 39154 6098 45916 6198
rect 46016 6098 46021 6198
rect 39368 5850 39468 6098
rect 42330 5850 42430 6098
rect 45911 6093 46021 6098
rect 37014 4858 37020 5066
rect 37228 4858 37749 5066
rect 37149 2926 37749 4858
rect 37996 4099 39784 5850
rect 37996 4050 38915 4099
rect 38910 3999 38915 4050
rect 39015 4050 39784 4099
rect 40026 4105 41814 5850
rect 40026 4050 40279 4105
rect 39015 3999 39020 4050
rect 40273 4007 40279 4050
rect 40377 4050 41814 4105
rect 42186 4097 43974 5850
rect 42186 4050 43087 4097
rect 40377 4007 40383 4050
rect 40278 4006 40378 4007
rect 38910 3994 39020 3999
rect 43082 3997 43087 4050
rect 43187 4050 43974 4097
rect 44226 4089 46014 5850
rect 44226 4050 44491 4089
rect 43187 3997 43192 4050
rect 43082 3992 43192 3997
rect 44485 3991 44491 4050
rect 44589 4050 46014 4089
rect 46417 5008 47017 6464
rect 48476 5981 48576 5982
rect 48471 5883 48477 5981
rect 48575 5883 48581 5981
rect 48476 5758 48576 5883
rect 48476 5736 49388 5758
rect 48476 5676 49306 5736
rect 49366 5676 49388 5736
rect 48476 5658 49388 5676
rect 53048 5604 53148 5610
rect 49924 5587 53048 5604
rect 49924 5527 49940 5587
rect 50000 5527 53048 5587
rect 49924 5504 53048 5527
rect 53048 5498 53148 5504
rect 46417 4846 47048 5008
rect 47210 4846 47216 5008
rect 52183 4956 52281 4961
rect 52183 4955 66110 4956
rect 52281 4936 66110 4955
rect 52281 4876 66026 4936
rect 66086 4876 66110 4936
rect 52281 4857 66110 4876
rect 52183 4856 66110 4857
rect 52183 4851 52281 4856
rect 44589 3991 44595 4050
rect 44490 3990 44590 3991
rect 41543 3960 41641 3965
rect 42074 3960 42174 3966
rect 45743 3960 45841 3965
rect 46238 3960 46338 3966
rect 41542 3959 42074 3960
rect 41542 3861 41543 3959
rect 41641 3861 42074 3959
rect 41542 3860 42074 3861
rect 45742 3959 46238 3960
rect 45742 3861 45743 3959
rect 45841 3861 46238 3959
rect 45742 3860 46238 3861
rect 41543 3855 41641 3860
rect 42074 3854 42174 3860
rect 45743 3855 45841 3860
rect 46238 3854 46338 3860
rect 40780 3799 40900 3804
rect 43688 3799 43788 3800
rect 39488 3797 39588 3798
rect 39483 3750 39489 3797
rect 36943 2740 36949 2926
rect 37135 2740 37749 2926
rect -10086 1422 -9986 1684
rect -7176 1422 -7076 1684
rect -10086 1322 -7076 1422
rect -3207 1064 -2607 2202
rect 36054 1691 36154 2238
rect -2334 1625 -2234 1626
rect -2339 1527 -2333 1625
rect -2235 1527 -2229 1625
rect 36049 1593 36055 1691
rect 36153 1593 36159 1691
rect 36054 1592 36154 1593
rect -7140 1062 -2607 1064
rect -12475 512 -2607 1062
rect -12475 460 -11156 512
rect -10918 460 -8744 512
rect -11156 268 -10918 274
rect -8506 460 -6332 512
rect -8744 268 -8506 274
rect -6094 462 -3920 512
rect -6094 460 -5990 462
rect -3978 460 -3920 462
rect -6332 268 -6094 274
rect -3682 462 -2607 512
rect -2334 602 -2230 1527
rect 37149 1330 37749 2740
rect 37996 3699 39489 3750
rect 39587 3750 39593 3797
rect 40780 3750 40785 3799
rect 39587 3699 39784 3750
rect 37996 1950 39784 3699
rect 40026 3689 40785 3750
rect 40895 3750 40900 3799
rect 43683 3750 43689 3799
rect 40895 3689 41814 3750
rect 40026 1950 41814 3689
rect 42186 3701 43689 3750
rect 43787 3750 43793 3799
rect 45056 3787 45176 3792
rect 45056 3750 45061 3787
rect 43787 3701 43974 3750
rect 42186 1950 43974 3701
rect 44226 3677 45061 3750
rect 45171 3750 45176 3787
rect 45171 3677 46014 3750
rect 44226 1950 46014 3677
rect 46417 2908 47017 4846
rect 48482 3756 48582 3762
rect 48582 3736 49378 3756
rect 48582 3676 49302 3736
rect 49362 3676 49378 3736
rect 48582 3656 49378 3676
rect 48482 3650 48582 3656
rect 52181 3605 52283 3611
rect 50066 3587 52181 3604
rect 50066 3527 50082 3587
rect 50142 3527 52181 3587
rect 50066 3504 52181 3527
rect 52181 3497 52283 3503
rect 61918 2933 62248 2938
rect 46417 2740 47010 2908
rect 47178 2740 47184 2908
rect 61918 2843 62153 2933
rect 62243 2843 62248 2933
rect 53051 2834 53149 2839
rect 61918 2838 62248 2843
rect 61918 2834 62018 2838
rect 53051 2833 62018 2834
rect 39542 1692 39642 1950
rect 42452 1692 42552 1950
rect 39160 1592 39166 1692
rect 39266 1670 46162 1692
rect 39266 1610 46088 1670
rect 46148 1610 46162 1670
rect 39266 1592 46162 1610
rect 46417 1330 47017 2740
rect 53149 2735 62018 2833
rect 53051 2734 62018 2735
rect 53051 2729 53149 2734
rect 52177 1672 52287 1678
rect 49806 1646 52177 1672
rect 49806 1586 49828 1646
rect 49888 1586 52177 1646
rect 49806 1562 52177 1586
rect 52177 1556 52287 1562
rect 37149 798 47017 1330
rect 37149 728 38494 798
rect 37149 726 37749 728
rect -2334 582 8126 602
rect -2334 522 8042 582
rect 8102 522 8126 582
rect 38722 796 47017 798
rect 38722 726 40906 796
rect 40904 710 40906 726
rect 38494 564 38722 570
rect 41134 726 43250 796
rect 43248 710 43250 726
rect 40906 562 41134 568
rect 43478 728 45638 796
rect 43478 726 44560 728
rect 43250 562 43478 568
rect 45866 730 47017 796
rect 45866 728 47016 730
rect 45866 708 45868 728
rect 45638 562 45866 568
rect -2334 502 8126 522
rect -2334 500 -2234 502
rect -3682 460 -3578 462
rect -3920 268 -3682 274
rect 3432 64 34918 110
rect 3432 -90 3478 64
rect 34878 -90 34918 64
rect 3432 -136 34918 -90
rect 57432 64 88918 110
rect 57432 -90 57478 64
rect 88878 -90 88918 64
rect 57432 -136 88918 -90
rect -1276 -276 -656 -271
rect -1276 -576 -1266 -276
rect -666 -576 -656 -276
rect -1276 -581 -656 -576
rect 35156 -276 35776 -271
rect 35156 -576 35166 -276
rect 35766 -576 35776 -276
rect 35156 -581 35776 -576
rect 52724 -276 53344 -271
rect 52724 -576 52734 -276
rect 53334 -576 53344 -276
rect 52724 -581 53344 -576
rect 89156 -276 89776 -271
rect 89156 -576 89166 -276
rect 89766 -576 89776 -276
rect 89156 -581 89776 -576
<< via3 >>
rect 11434 27856 12034 28156
rect 35066 27856 35666 28156
rect 65434 27856 66034 28156
rect 89066 27856 89666 28156
rect -1419 27642 -1349 27647
rect -1419 27583 -1414 27642
rect -1414 27583 -1354 27642
rect -1354 27583 -1349 27642
rect 15011 27560 31796 27774
rect 47824 27564 48462 27680
rect 69011 27560 85796 27774
rect -713 26548 -649 27092
rect 1881 26549 1945 27093
rect 4481 26549 4545 27093
rect 7081 26549 7145 27093
rect 9681 26549 9745 27093
rect 10681 26548 10745 27092
rect 38430 26420 38578 26568
rect 41348 26410 41506 26568
rect 53287 26548 53351 27092
rect 55881 26549 55945 27093
rect 58481 26549 58545 27093
rect 61081 26549 61145 27093
rect 63681 26549 63745 27093
rect 64681 26548 64745 27092
rect -715 24048 -651 26192
rect 1882 24048 1946 26192
rect 4482 24048 4546 26192
rect 7082 24048 7146 26192
rect 9682 24048 9746 26192
rect 10679 24048 10743 26192
rect 37050 24644 37182 24776
rect -715 21548 -651 23692
rect 1882 21547 1946 23691
rect 4482 21547 4546 23691
rect 7082 21547 7146 23691
rect 9682 21547 9746 23691
rect 10679 21548 10743 23692
rect 36468 23470 36568 23570
rect -715 19048 -651 21192
rect 1882 19047 1946 21191
rect 4482 19047 4546 21191
rect 7082 19047 7146 21191
rect 9682 19047 9746 21191
rect 10679 19048 10743 21192
rect 40402 23770 40502 23870
rect 42912 24632 43048 24768
rect 46576 24434 46676 24534
rect 41563 23613 41661 23711
rect 42030 23612 42130 23712
rect 37076 22556 37196 22676
rect 39493 23469 39591 23567
rect 42864 22518 43004 22658
rect 49760 21600 49860 21700
rect 46405 21283 46503 21381
rect 53285 24048 53349 26192
rect 55882 24048 55946 26192
rect 58482 24048 58546 26192
rect 61082 24048 61146 26192
rect 63682 24048 63746 26192
rect 64679 24048 64743 26192
rect 52144 23614 52244 23714
rect 51794 20966 51894 21066
rect 36473 19827 36571 19925
rect 9201 18819 9299 18917
rect -715 16548 -651 18692
rect 1882 16547 1946 18691
rect 4482 16547 4546 18691
rect 7082 16547 7146 18691
rect 9682 16547 9746 18691
rect 10679 16548 10743 18692
rect 38494 20312 38672 20490
rect 40894 20312 41072 20490
rect 43294 20312 43472 20490
rect 45420 20312 45598 20490
rect 47594 20312 47772 20490
rect 49994 20312 50172 20490
rect 39078 19826 39178 19926
rect 37150 18582 37358 18790
rect 9861 16323 9959 16421
rect -717 15650 -653 16194
rect 1881 15649 1945 16193
rect 4481 15649 4545 16193
rect 7081 15649 7145 16193
rect 9681 15649 9745 16193
rect 10681 15650 10745 16194
rect -13471 10633 -13373 10731
rect -11154 14022 -11008 14168
rect -8836 13984 -8646 14174
rect -6346 13974 -6170 14150
rect -3940 14010 -3782 14168
rect -13107 13039 -13009 13137
rect -10574 13038 -10474 13138
rect -12624 11880 -12530 11974
rect -9225 10931 -9127 11029
rect -5269 10931 -5171 11029
rect -2396 12804 -2296 12904
rect -2524 11764 -2432 11856
rect -8101 10783 -8003 10881
rect -7570 10782 -7470 10882
rect -3901 10781 -3803 10879
rect -3392 10780 -3292 10880
rect -12634 9930 -12554 10010
rect -13099 8521 -13001 8619
rect -13303 3439 -13205 3537
rect -10355 10633 -10257 10731
rect -6555 10635 -6457 10733
rect -2518 9742 -2412 9848
rect -10534 8520 -10434 8620
rect 36255 15277 36353 15375
rect 36255 9443 36353 9541
rect -1755 8765 -1657 8863
rect -11197 7406 -10957 7646
rect -8785 7406 -8545 7646
rect -6373 7406 -6133 7646
rect -3961 7406 -3721 7646
rect 35229 7639 35327 7737
rect -11198 6814 -10956 7056
rect -8786 6814 -8544 7056
rect -6374 6814 -6132 7056
rect -3962 6814 -3720 7056
rect -12731 5567 -12633 5665
rect -12586 4616 -12436 4766
rect -9365 3729 -9267 3827
rect -5143 3725 -5029 3839
rect -2421 5567 -2323 5665
rect -2660 4562 -2506 4716
rect -8085 3583 -7987 3681
rect -7554 3582 -7454 3682
rect -3885 3585 -3787 3683
rect -3382 3584 -3282 3684
rect -12580 2524 -12454 2650
rect -13097 1529 -12999 1627
rect -10167 3439 -10069 3537
rect -5908 3426 -5792 3542
rect -2666 2504 -2506 2664
rect 40417 17731 40515 17829
rect 44643 17719 44741 17817
rect 48765 17729 48863 17827
rect 51338 18570 51500 18732
rect 41673 17579 41771 17677
rect 42204 17578 42304 17678
rect 45873 17579 45971 17677
rect 46404 17578 46504 17678
rect 50073 17579 50171 17677
rect 50604 17578 50704 17678
rect 37079 16464 37265 16650
rect 39619 17425 39717 17523
rect 43819 17425 43917 17523
rect 48019 17423 48117 17521
rect 51364 16470 51532 16638
rect 39298 15276 39398 15376
rect 53285 21548 53349 23692
rect 55882 21547 55946 23691
rect 58482 21547 58546 23691
rect 61082 21547 61146 23691
rect 63682 21547 63746 23691
rect 64679 21548 64743 23692
rect 53285 19048 53349 21192
rect 55882 19047 55946 21191
rect 58482 19047 58546 21191
rect 61082 19047 61146 21191
rect 63682 19047 63746 21191
rect 64679 19048 64743 21192
rect 63201 18819 63299 18917
rect 53285 16548 53349 18692
rect 55882 16547 55946 18691
rect 58482 16547 58546 18691
rect 61082 16547 61146 18691
rect 63682 16547 63746 18691
rect 64679 16548 64743 18692
rect 63861 16323 63959 16421
rect 53283 15650 53347 16194
rect 55881 15649 55945 16193
rect 58481 15649 58545 16193
rect 61081 15649 61145 16193
rect 63681 15649 63745 16193
rect 64681 15650 64745 16194
rect 52380 15000 52480 15100
rect 36749 13483 36847 13581
rect 38478 14158 38636 14316
rect 40890 14158 41048 14316
rect 43290 14158 43448 14316
rect 45690 14158 45848 14316
rect 47690 14158 47848 14316
rect 50090 14158 50248 14316
rect 37002 12460 37210 12668
rect 40293 11611 40391 11709
rect 44513 11611 44611 11709
rect 47030 12448 47192 12610
rect 41543 11461 41641 11559
rect 42074 11460 42174 11560
rect 45743 11461 45841 11559
rect 46218 11460 46318 11560
rect 36931 10342 37117 10528
rect 39489 11313 39587 11411
rect 43689 11295 43787 11393
rect 46992 10342 47160 10510
rect 38476 8172 38704 8400
rect 40888 8170 41116 8398
rect 43232 8170 43460 8398
rect 45620 8170 45848 8398
rect 36996 7638 37096 7738
rect 53050 7622 53150 7722
rect 38428 6992 38610 7174
rect 40828 6992 41010 7174
rect 43240 6992 43422 7174
rect 45640 6992 45822 7174
rect 36459 6099 36557 6197
rect 39054 6098 39154 6198
rect 37020 4858 37228 5066
rect 40279 4007 40377 4105
rect 44491 3991 44589 4089
rect 48477 5883 48575 5981
rect 53048 5504 53148 5604
rect 47048 4846 47210 5008
rect 52183 4857 52281 4955
rect 41543 3861 41641 3959
rect 42074 3860 42174 3960
rect 45743 3861 45841 3959
rect 46238 3860 46338 3960
rect 36949 2740 37135 2926
rect -2333 1527 -2235 1625
rect 36055 1593 36153 1691
rect -11156 274 -10918 512
rect -8744 274 -8506 512
rect -6332 274 -6094 512
rect -3920 274 -3682 512
rect 39489 3699 39587 3797
rect 43689 3701 43787 3799
rect 48482 3656 48582 3756
rect 52181 3503 52283 3605
rect 47010 2740 47178 2908
rect 39166 1592 39266 1692
rect 53051 2735 53149 2833
rect 52177 1562 52287 1672
rect 38494 570 38722 798
rect 40906 568 41134 796
rect 43250 568 43478 796
rect 45638 568 45866 796
rect 3478 -90 34878 64
rect 57478 -90 88878 64
rect -1266 -576 -666 -276
rect 35166 -576 35766 -276
rect 52734 -576 53334 -276
rect 89166 -576 89766 -276
<< mimcap >>
rect -1228 26980 -828 27020
rect -1228 26660 -1188 26980
rect -868 26660 -828 26980
rect -1228 26620 -828 26660
rect -234 26981 1766 27021
rect -234 26661 -194 26981
rect 1726 26661 1766 26981
rect -234 26621 1766 26661
rect 2366 26981 4366 27021
rect 2366 26661 2406 26981
rect 4326 26661 4366 26981
rect 2366 26621 4366 26661
rect 4966 26981 6966 27021
rect 4966 26661 5006 26981
rect 6926 26661 6966 26981
rect 4966 26621 6966 26661
rect 7566 26981 9566 27021
rect 7566 26661 7606 26981
rect 9526 26661 9566 26981
rect 7566 26621 9566 26661
rect 10166 26980 10566 27020
rect 10166 26660 10206 26980
rect 10526 26660 10566 26980
rect 10166 26620 10566 26660
rect 52772 26980 53172 27020
rect 52772 26660 52812 26980
rect 53132 26660 53172 26980
rect 52772 26620 53172 26660
rect 53766 26981 55766 27021
rect 53766 26661 53806 26981
rect 55726 26661 55766 26981
rect 53766 26621 55766 26661
rect 56366 26981 58366 27021
rect 56366 26661 56406 26981
rect 58326 26661 58366 26981
rect 56366 26621 58366 26661
rect 58966 26981 60966 27021
rect 58966 26661 59006 26981
rect 60926 26661 60966 26981
rect 58966 26621 60966 26661
rect 61566 26981 63566 27021
rect 61566 26661 61606 26981
rect 63526 26661 63566 26981
rect 61566 26621 63566 26661
rect 64166 26980 64566 27020
rect 64166 26660 64206 26980
rect 64526 26660 64566 26980
rect 64166 26620 64566 26660
rect 37250 26340 39650 26380
rect -1230 26080 -830 26120
rect -1230 24160 -1190 26080
rect -870 24160 -830 26080
rect -1230 24120 -830 24160
rect -233 26080 1767 26120
rect -233 24160 -193 26080
rect 1727 24160 1767 26080
rect -233 24120 1767 24160
rect 2367 26080 4367 26120
rect 2367 24160 2407 26080
rect 4327 24160 4367 26080
rect 2367 24120 4367 24160
rect 4967 26080 6967 26120
rect 4967 24160 5007 26080
rect 6927 24160 6967 26080
rect 4967 24120 6967 24160
rect 7567 26080 9567 26120
rect 7567 24160 7607 26080
rect 9527 24160 9567 26080
rect 7567 24120 9567 24160
rect 10164 26080 10564 26120
rect 10164 24160 10204 26080
rect 10524 24160 10564 26080
rect 37250 26020 37290 26340
rect 39610 26020 39650 26340
rect 37250 25980 39650 26020
rect 40250 26340 42650 26380
rect 40250 26020 40290 26340
rect 42610 26020 42650 26340
rect 40250 25980 42650 26020
rect 52770 26080 53170 26120
rect 10164 24120 10564 24160
rect 37266 25476 37666 25516
rect 37266 23956 37306 25476
rect 37626 23956 37666 25476
rect 37266 23916 37666 23956
rect 38118 25472 39718 25512
rect 38118 23952 38158 25472
rect 39678 23952 39718 25472
rect 38118 23912 39718 23952
rect 40148 25472 41748 25512
rect 40148 23952 40188 25472
rect 41708 23952 41748 25472
rect 40148 23912 41748 23952
rect 42366 25476 42766 25516
rect 42366 23956 42406 25476
rect 42726 23956 42766 25476
rect 52770 24160 52810 26080
rect 53130 24160 53170 26080
rect 52770 24120 53170 24160
rect 53767 26080 55767 26120
rect 53767 24160 53807 26080
rect 55727 24160 55767 26080
rect 53767 24120 55767 24160
rect 56367 26080 58367 26120
rect 56367 24160 56407 26080
rect 58327 24160 58367 26080
rect 56367 24120 58367 24160
rect 58967 26080 60967 26120
rect 58967 24160 59007 26080
rect 60927 24160 60967 26080
rect 58967 24120 60967 24160
rect 61567 26080 63567 26120
rect 61567 24160 61607 26080
rect 63527 24160 63567 26080
rect 61567 24120 63567 24160
rect 64164 26080 64564 26120
rect 64164 24160 64204 26080
rect 64524 24160 64564 26080
rect 64164 24120 64564 24160
rect 42366 23916 42766 23956
rect -1230 23580 -830 23620
rect -1230 21660 -1190 23580
rect -870 21660 -830 23580
rect -1230 21620 -830 21660
rect -233 23579 1767 23619
rect -233 21659 -193 23579
rect 1727 21659 1767 23579
rect -233 21619 1767 21659
rect 2367 23579 4367 23619
rect 2367 21659 2407 23579
rect 4327 21659 4367 23579
rect 2367 21619 4367 21659
rect 4967 23579 6967 23619
rect 4967 21659 5007 23579
rect 6927 21659 6967 23579
rect 4967 21619 6967 21659
rect 7567 23579 9567 23619
rect 7567 21659 7607 23579
rect 9527 21659 9567 23579
rect 7567 21619 9567 21659
rect 10164 23580 10564 23620
rect 10164 21660 10204 23580
rect 10524 21660 10564 23580
rect 52770 23580 53170 23620
rect 37266 23372 37666 23412
rect 37266 21852 37306 23372
rect 37626 21852 37666 23372
rect 37266 21812 37666 21852
rect 38118 23372 39718 23412
rect 38118 21852 38158 23372
rect 39678 21852 39718 23372
rect 38118 21812 39718 21852
rect 40148 23372 41748 23412
rect 40148 21852 40188 23372
rect 41708 21852 41748 23372
rect 40148 21812 41748 21852
rect 42366 23372 42766 23412
rect 42366 21852 42406 23372
rect 42726 21852 42766 23372
rect 42366 21812 42766 21852
rect 10164 21620 10564 21660
rect 52770 21660 52810 23580
rect 53130 21660 53170 23580
rect 52770 21620 53170 21660
rect 53767 23579 55767 23619
rect 53767 21659 53807 23579
rect 55727 21659 55767 23579
rect 53767 21619 55767 21659
rect 56367 23579 58367 23619
rect 56367 21659 56407 23579
rect 58327 21659 58367 23579
rect 56367 21619 58367 21659
rect 58967 23579 60967 23619
rect 58967 21659 59007 23579
rect 60927 21659 60967 23579
rect 58967 21619 60967 21659
rect 61567 23579 63567 23619
rect 61567 21659 61607 23579
rect 63527 21659 63567 23579
rect 61567 21619 63567 21659
rect 64164 23580 64564 23620
rect 64164 21660 64204 23580
rect 64524 21660 64564 23580
rect 64164 21620 64564 21660
rect -1230 21080 -830 21120
rect -1230 19160 -1190 21080
rect -870 19160 -830 21080
rect -1230 19120 -830 19160
rect -233 21079 1767 21119
rect -233 19159 -193 21079
rect 1727 19159 1767 21079
rect -233 19119 1767 19159
rect 2367 21079 4367 21119
rect 2367 19159 2407 21079
rect 4327 19159 4367 21079
rect 2367 19119 4367 19159
rect 4967 21079 6967 21119
rect 4967 19159 5007 21079
rect 6927 19159 6967 21079
rect 4967 19119 6967 19159
rect 7567 21079 9567 21119
rect 7567 19159 7607 21079
rect 9527 19159 9567 21079
rect 7567 19119 9567 19159
rect 10164 21080 10564 21120
rect 10164 19160 10204 21080
rect 10524 19160 10564 21080
rect 52770 21080 53170 21120
rect 37363 20886 39763 20926
rect 37363 20566 37403 20886
rect 39723 20566 39763 20886
rect 37363 20526 39763 20566
rect 40146 20886 41746 20926
rect 40146 20566 40186 20886
rect 41706 20566 41746 20886
rect 40146 20526 41746 20566
rect 42534 20888 44134 20928
rect 42534 20568 42574 20888
rect 44094 20568 44134 20888
rect 42534 20528 44134 20568
rect 44642 20888 46242 20928
rect 44642 20568 44682 20888
rect 46202 20568 46242 20888
rect 44642 20528 46242 20568
rect 46928 20888 48528 20928
rect 46928 20568 46968 20888
rect 48488 20568 48528 20888
rect 46928 20528 48528 20568
rect 48911 20888 51311 20928
rect 48911 20568 48951 20888
rect 51271 20568 51311 20888
rect 48911 20528 51311 20568
rect 10164 19120 10564 19160
rect 37380 19434 37780 19474
rect -1230 18580 -830 18620
rect -1230 16660 -1190 18580
rect -870 16660 -830 18580
rect -1230 16620 -830 16660
rect -233 18579 1767 18619
rect -233 16659 -193 18579
rect 1727 16659 1767 18579
rect -233 16619 1767 16659
rect 2367 18579 4367 18619
rect 2367 16659 2407 18579
rect 4327 16659 4367 18579
rect 2367 16619 4367 16659
rect 4967 18579 6967 18619
rect 4967 16659 5007 18579
rect 6927 16659 6967 18579
rect 4967 16619 6967 16659
rect 7567 18579 9567 18619
rect 7567 16659 7607 18579
rect 9527 16659 9567 18579
rect 7567 16619 9567 16659
rect 10164 18580 10564 18620
rect 10164 16660 10204 18580
rect 10524 16660 10564 18580
rect 37380 17914 37420 19434
rect 37740 17914 37780 19434
rect 37380 17874 37780 17914
rect 38226 19434 39826 19474
rect 38226 17914 38266 19434
rect 39786 17914 39826 19434
rect 38226 17874 39826 17914
rect 40256 19434 41856 19474
rect 40256 17914 40296 19434
rect 41816 17914 41856 19434
rect 40256 17874 41856 17914
rect 42416 19434 44016 19474
rect 42416 17914 42456 19434
rect 43976 17914 44016 19434
rect 42416 17874 44016 17914
rect 44456 19434 46056 19474
rect 44456 17914 44496 19434
rect 46016 17914 46056 19434
rect 44456 17874 46056 17914
rect 46612 19434 48212 19474
rect 46612 17914 46652 19434
rect 48172 17914 48212 19434
rect 46612 17874 48212 17914
rect 48652 19434 50252 19474
rect 48652 17914 48692 19434
rect 50212 17914 50252 19434
rect 48652 17874 50252 17914
rect 50892 19434 51292 19474
rect 50892 17914 50932 19434
rect 51252 17914 51292 19434
rect 52770 19160 52810 21080
rect 53130 19160 53170 21080
rect 52770 19120 53170 19160
rect 53767 21079 55767 21119
rect 53767 19159 53807 21079
rect 55727 19159 55767 21079
rect 53767 19119 55767 19159
rect 56367 21079 58367 21119
rect 56367 19159 56407 21079
rect 58327 19159 58367 21079
rect 56367 19119 58367 19159
rect 58967 21079 60967 21119
rect 58967 19159 59007 21079
rect 60927 19159 60967 21079
rect 58967 19119 60967 19159
rect 61567 21079 63567 21119
rect 61567 19159 61607 21079
rect 63527 19159 63567 21079
rect 61567 19119 63567 19159
rect 64164 21080 64564 21120
rect 64164 19160 64204 21080
rect 64524 19160 64564 21080
rect 64164 19120 64564 19160
rect 50892 17874 51292 17914
rect 52770 18580 53170 18620
rect 10164 16620 10564 16660
rect 37380 17330 37780 17370
rect -1232 16082 -832 16122
rect -1232 15762 -1192 16082
rect -872 15762 -832 16082
rect -1232 15722 -832 15762
rect -234 16081 1766 16121
rect -234 15761 -194 16081
rect 1726 15761 1766 16081
rect -234 15721 1766 15761
rect 2366 16081 4366 16121
rect 2366 15761 2406 16081
rect 4326 15761 4366 16081
rect 2366 15721 4366 15761
rect 4966 16081 6966 16121
rect 4966 15761 5006 16081
rect 6926 15761 6966 16081
rect 4966 15721 6966 15761
rect 7566 16081 9566 16121
rect 7566 15761 7606 16081
rect 9526 15761 9566 16081
rect 7566 15721 9566 15761
rect 10166 16082 10566 16122
rect 10166 15762 10206 16082
rect 10526 15762 10566 16082
rect 37380 15810 37420 17330
rect 37740 15810 37780 17330
rect 37380 15770 37780 15810
rect 38226 17334 39826 17374
rect 38226 15814 38266 17334
rect 39786 15814 39826 17334
rect 38226 15774 39826 15814
rect 40256 17334 41856 17374
rect 40256 15814 40296 17334
rect 41816 15814 41856 17334
rect 40256 15774 41856 15814
rect 42416 17334 44016 17374
rect 42416 15814 42456 17334
rect 43976 15814 44016 17334
rect 42416 15774 44016 15814
rect 44456 17334 46056 17374
rect 44456 15814 44496 17334
rect 46016 15814 46056 17334
rect 44456 15774 46056 15814
rect 46612 17334 48212 17374
rect 46612 15814 46652 17334
rect 48172 15814 48212 17334
rect 46612 15774 48212 15814
rect 48652 17334 50252 17374
rect 48652 15814 48692 17334
rect 50212 15814 50252 17334
rect 48652 15774 50252 15814
rect 50892 17330 51292 17370
rect 50892 15810 50932 17330
rect 51252 15810 51292 17330
rect 52770 16660 52810 18580
rect 53130 16660 53170 18580
rect 52770 16620 53170 16660
rect 53767 18579 55767 18619
rect 53767 16659 53807 18579
rect 55727 16659 55767 18579
rect 53767 16619 55767 16659
rect 56367 18579 58367 18619
rect 56367 16659 56407 18579
rect 58327 16659 58367 18579
rect 56367 16619 58367 16659
rect 58967 18579 60967 18619
rect 58967 16659 59007 18579
rect 60927 16659 60967 18579
rect 58967 16619 60967 16659
rect 61567 18579 63567 18619
rect 61567 16659 61607 18579
rect 63527 16659 63567 18579
rect 61567 16619 63567 16659
rect 64164 18580 64564 18620
rect 64164 16660 64204 18580
rect 64524 16660 64564 18580
rect 64164 16620 64564 16660
rect 50892 15770 51292 15810
rect 52768 16082 53168 16122
rect 10166 15722 10566 15762
rect 52768 15762 52808 16082
rect 53128 15762 53168 16082
rect 52768 15722 53168 15762
rect 53766 16081 55766 16121
rect 53766 15761 53806 16081
rect 55726 15761 55766 16081
rect 53766 15721 55766 15761
rect 56366 16081 58366 16121
rect 56366 15761 56406 16081
rect 58326 15761 58366 16081
rect 56366 15721 58366 15761
rect 58966 16081 60966 16121
rect 58966 15761 59006 16081
rect 60926 15761 60966 16081
rect 58966 15721 60966 15761
rect 61566 16081 63566 16121
rect 61566 15761 61606 16081
rect 63526 15761 63566 16081
rect 61566 15721 63566 15761
rect 64166 16082 64566 16122
rect 64166 15762 64206 16082
rect 64526 15762 64566 16082
rect 64166 15722 64566 15762
rect 37363 14726 39763 14766
rect 37363 14406 37403 14726
rect 39723 14406 39763 14726
rect 37363 14366 39763 14406
rect 40146 14726 41746 14766
rect 40146 14406 40186 14726
rect 41706 14406 41746 14726
rect 40146 14366 41746 14406
rect 42534 14728 44134 14768
rect 42534 14408 42574 14728
rect 44094 14408 44134 14728
rect 42534 14368 44134 14408
rect 44816 14728 46416 14768
rect 44816 14408 44856 14728
rect 46376 14408 46416 14728
rect 44816 14368 46416 14408
rect 46928 14728 48528 14768
rect 46928 14408 46968 14728
rect 48488 14408 48528 14728
rect 46928 14368 48528 14408
rect 48911 14728 51311 14768
rect 48911 14408 48951 14728
rect 51271 14408 51311 14728
rect 48911 14368 51311 14408
rect -12243 13858 -9843 13898
rect -12243 13538 -12203 13858
rect -9883 13538 -9843 13858
rect -12243 13498 -9843 13538
rect -9460 13858 -7860 13898
rect -9460 13538 -9420 13858
rect -7900 13538 -7860 13858
rect -9460 13498 -7860 13538
rect -7072 13860 -5472 13900
rect -7072 13540 -7032 13860
rect -5512 13540 -5472 13860
rect -7072 13500 -5472 13540
rect -5089 13860 -2689 13900
rect -5089 13540 -5049 13860
rect -2729 13540 -2689 13860
rect -5089 13500 -2689 13540
rect 37232 13312 37632 13352
rect -12374 12644 -11974 12684
rect -12374 11124 -12334 12644
rect -12014 11124 -11974 12644
rect -12374 11084 -11974 11124
rect -11528 12644 -9928 12684
rect -11528 11124 -11488 12644
rect -9968 11124 -9928 12644
rect -11528 11084 -9928 11124
rect -9498 12644 -7898 12684
rect -9498 11124 -9458 12644
rect -7938 11124 -7898 12644
rect -9498 11084 -7898 11124
rect -7338 12644 -5738 12684
rect -7338 11124 -7298 12644
rect -5778 11124 -5738 12644
rect -7338 11084 -5738 11124
rect -5298 12644 -3698 12684
rect -5298 11124 -5258 12644
rect -3738 11124 -3698 12644
rect -5298 11084 -3698 11124
rect -3108 12646 -2708 12686
rect -3108 11126 -3068 12646
rect -2748 11126 -2708 12646
rect 37232 11792 37272 13312
rect 37592 11792 37632 13312
rect 37232 11752 37632 11792
rect 38078 13312 39678 13352
rect 38078 11792 38118 13312
rect 39638 11792 39678 13312
rect 38078 11752 39678 11792
rect 40108 13312 41708 13352
rect 40108 11792 40148 13312
rect 41668 11792 41708 13312
rect 40108 11752 41708 11792
rect 42268 13312 43868 13352
rect 42268 11792 42308 13312
rect 43828 11792 43868 13312
rect 42268 11752 43868 11792
rect 44308 13312 45908 13352
rect 44308 11792 44348 13312
rect 45868 11792 45908 13312
rect 44308 11752 45908 11792
rect 46498 13314 46898 13354
rect 46498 11794 46538 13314
rect 46858 11794 46898 13314
rect 46498 11754 46898 11794
rect -3108 11086 -2708 11126
rect 37232 11208 37632 11248
rect -12374 10540 -11974 10580
rect -12374 9020 -12334 10540
rect -12014 9020 -11974 10540
rect -12374 8980 -11974 9020
rect -11528 10544 -9928 10584
rect -11528 9024 -11488 10544
rect -9968 9024 -9928 10544
rect -11528 8984 -9928 9024
rect -9498 10544 -7898 10584
rect -9498 9024 -9458 10544
rect -7938 9024 -7898 10544
rect -9498 8984 -7898 9024
rect -7338 10544 -5738 10584
rect -7338 9024 -7298 10544
rect -5778 9024 -5738 10544
rect -7338 8984 -5738 9024
rect -5298 10544 -3698 10584
rect -5298 9024 -5258 10544
rect -3738 9024 -3698 10544
rect -5298 8984 -3698 9024
rect -3108 10542 -2708 10582
rect -3108 9022 -3068 10542
rect -2748 9022 -2708 10542
rect 37232 9688 37272 11208
rect 37592 9688 37632 11208
rect 37232 9648 37632 9688
rect 38078 11212 39678 11252
rect 38078 9692 38118 11212
rect 39638 9692 39678 11212
rect 38078 9652 39678 9692
rect 40108 11212 41708 11252
rect 40108 9692 40148 11212
rect 41668 9692 41708 11212
rect 40108 9652 41708 9692
rect 42268 11212 43868 11252
rect 42268 9692 42308 11212
rect 43828 9692 43868 11212
rect 42268 9652 43868 9692
rect 44308 11212 45908 11252
rect 44308 9692 44348 11212
rect 45868 9692 45908 11212
rect 44308 9652 45908 9692
rect 46498 11210 46898 11250
rect 46498 9690 46538 11210
rect 46858 9690 46898 11210
rect 46498 9650 46898 9690
rect -3108 8982 -2708 9022
rect 37363 8790 39763 8830
rect 37363 8470 37403 8790
rect 39723 8470 39763 8790
rect 37363 8430 39763 8470
rect 40146 8790 41746 8830
rect 40146 8470 40186 8790
rect 41706 8470 41746 8790
rect 40146 8430 41746 8470
rect 42534 8792 44134 8832
rect 42534 8472 42574 8792
rect 44094 8472 44134 8792
rect 42534 8432 44134 8472
rect 44517 8792 46917 8832
rect 44517 8472 44557 8792
rect 46877 8472 46917 8792
rect 44517 8432 46917 8472
rect -12243 8122 -9843 8162
rect -12243 7802 -12203 8122
rect -9883 7802 -9843 8122
rect -12243 7762 -9843 7802
rect -9460 8122 -7860 8162
rect -9460 7802 -9420 8122
rect -7900 7802 -7860 8122
rect -9460 7762 -7860 7802
rect -7072 8124 -5472 8164
rect -7072 7804 -7032 8124
rect -5512 7804 -5472 8124
rect -7072 7764 -5472 7804
rect -5089 8124 -2689 8164
rect -5089 7804 -5049 8124
rect -2729 7804 -2689 8124
rect -5089 7764 -2689 7804
rect 37381 6924 39781 6964
rect -12243 6658 -9843 6698
rect -12243 6338 -12203 6658
rect -9883 6338 -9843 6658
rect -12243 6298 -9843 6338
rect -9460 6658 -7860 6698
rect -9460 6338 -9420 6658
rect -7900 6338 -7860 6658
rect -9460 6298 -7860 6338
rect -7072 6660 -5472 6700
rect -7072 6340 -7032 6660
rect -5512 6340 -5472 6660
rect -7072 6300 -5472 6340
rect -5089 6660 -2689 6700
rect -5089 6340 -5049 6660
rect -2729 6340 -2689 6660
rect 37381 6604 37421 6924
rect 39741 6604 39781 6924
rect 37381 6564 39781 6604
rect 40164 6924 41764 6964
rect 40164 6604 40204 6924
rect 41724 6604 41764 6924
rect 40164 6564 41764 6604
rect 42552 6926 44152 6966
rect 42552 6606 42592 6926
rect 44112 6606 44152 6926
rect 42552 6566 44152 6606
rect 44535 6926 46935 6966
rect 44535 6606 44575 6926
rect 46895 6606 46935 6926
rect 44535 6566 46935 6606
rect -5089 6300 -2689 6340
rect 37250 5710 37650 5750
rect -12374 5444 -11974 5484
rect -12374 3924 -12334 5444
rect -12014 3924 -11974 5444
rect -12374 3884 -11974 3924
rect -11528 5444 -9928 5484
rect -11528 3924 -11488 5444
rect -9968 3924 -9928 5444
rect -11528 3884 -9928 3924
rect -9498 5444 -7898 5484
rect -9498 3924 -9458 5444
rect -7938 3924 -7898 5444
rect -9498 3884 -7898 3924
rect -7338 5444 -5738 5484
rect -7338 3924 -7298 5444
rect -5778 3924 -5738 5444
rect -7338 3884 -5738 3924
rect -5298 5444 -3698 5484
rect -5298 3924 -5258 5444
rect -3738 3924 -3698 5444
rect -5298 3884 -3698 3924
rect -3108 5446 -2708 5486
rect -3108 3926 -3068 5446
rect -2748 3926 -2708 5446
rect 37250 4190 37290 5710
rect 37610 4190 37650 5710
rect 37250 4150 37650 4190
rect 38096 5710 39696 5750
rect 38096 4190 38136 5710
rect 39656 4190 39696 5710
rect 38096 4150 39696 4190
rect 40126 5710 41726 5750
rect 40126 4190 40166 5710
rect 41686 4190 41726 5710
rect 40126 4150 41726 4190
rect 42286 5710 43886 5750
rect 42286 4190 42326 5710
rect 43846 4190 43886 5710
rect 42286 4150 43886 4190
rect 44326 5710 45926 5750
rect 44326 4190 44366 5710
rect 45886 4190 45926 5710
rect 44326 4150 45926 4190
rect 46516 5712 46916 5752
rect 46516 4192 46556 5712
rect 46876 4192 46916 5712
rect 46516 4152 46916 4192
rect -3108 3886 -2708 3926
rect 37250 3606 37650 3646
rect -12374 3340 -11974 3380
rect -12374 1820 -12334 3340
rect -12014 1820 -11974 3340
rect -12374 1780 -11974 1820
rect -11528 3344 -9928 3384
rect -11528 1824 -11488 3344
rect -9968 1824 -9928 3344
rect -11528 1784 -9928 1824
rect -9498 3344 -7898 3384
rect -9498 1824 -9458 3344
rect -7938 1824 -7898 3344
rect -9498 1784 -7898 1824
rect -7338 3344 -5738 3384
rect -7338 1824 -7298 3344
rect -5778 1824 -5738 3344
rect -7338 1784 -5738 1824
rect -5298 3344 -3698 3384
rect -5298 1824 -5258 3344
rect -3738 1824 -3698 3344
rect -5298 1784 -3698 1824
rect -3108 3342 -2708 3382
rect -3108 1822 -3068 3342
rect -2748 1822 -2708 3342
rect 37250 2086 37290 3606
rect 37610 2086 37650 3606
rect 37250 2046 37650 2086
rect 38096 3610 39696 3650
rect 38096 2090 38136 3610
rect 39656 2090 39696 3610
rect 38096 2050 39696 2090
rect 40126 3610 41726 3650
rect 40126 2090 40166 3610
rect 41686 2090 41726 3610
rect 40126 2050 41726 2090
rect 42286 3610 43886 3650
rect 42286 2090 42326 3610
rect 43846 2090 43886 3610
rect 42286 2050 43886 2090
rect 44326 3610 45926 3650
rect 44326 2090 44366 3610
rect 45886 2090 45926 3610
rect 44326 2050 45926 2090
rect 46516 3608 46916 3648
rect 46516 2088 46556 3608
rect 46876 2088 46916 3608
rect 46516 2048 46916 2088
rect -3108 1782 -2708 1822
rect 37381 1188 39781 1228
rect -12243 922 -9843 962
rect -12243 602 -12203 922
rect -9883 602 -9843 922
rect -12243 562 -9843 602
rect -9460 922 -7860 962
rect -9460 602 -9420 922
rect -7900 602 -7860 922
rect -9460 562 -7860 602
rect -7072 924 -5472 964
rect -7072 604 -7032 924
rect -5512 604 -5472 924
rect -7072 564 -5472 604
rect -5089 924 -2689 964
rect -5089 604 -5049 924
rect -2729 604 -2689 924
rect 37381 868 37421 1188
rect 39741 868 39781 1188
rect 37381 828 39781 868
rect 40164 1188 41764 1228
rect 40164 868 40204 1188
rect 41724 868 41764 1188
rect 40164 828 41764 868
rect 42552 1190 44152 1230
rect 42552 870 42592 1190
rect 44112 870 44152 1190
rect 42552 830 44152 870
rect 44535 1190 46935 1230
rect 44535 870 44575 1190
rect 46895 870 46935 1190
rect 44535 830 46935 870
rect -5089 564 -2689 604
<< mimcapcontact >>
rect -1188 26660 -868 26980
rect -194 26661 1726 26981
rect 2406 26661 4326 26981
rect 5006 26661 6926 26981
rect 7606 26661 9526 26981
rect 10206 26660 10526 26980
rect 52812 26660 53132 26980
rect 53806 26661 55726 26981
rect 56406 26661 58326 26981
rect 59006 26661 60926 26981
rect 61606 26661 63526 26981
rect 64206 26660 64526 26980
rect -1190 24160 -870 26080
rect -193 24160 1727 26080
rect 2407 24160 4327 26080
rect 5007 24160 6927 26080
rect 7607 24160 9527 26080
rect 10204 24160 10524 26080
rect 37290 26020 39610 26340
rect 40290 26020 42610 26340
rect 37306 23956 37626 25476
rect 38158 23952 39678 25472
rect 40188 23952 41708 25472
rect 42406 23956 42726 25476
rect 52810 24160 53130 26080
rect 53807 24160 55727 26080
rect 56407 24160 58327 26080
rect 59007 24160 60927 26080
rect 61607 24160 63527 26080
rect 64204 24160 64524 26080
rect -1190 21660 -870 23580
rect -193 21659 1727 23579
rect 2407 21659 4327 23579
rect 5007 21659 6927 23579
rect 7607 21659 9527 23579
rect 10204 21660 10524 23580
rect 37306 21852 37626 23372
rect 38158 21852 39678 23372
rect 40188 21852 41708 23372
rect 42406 21852 42726 23372
rect 52810 21660 53130 23580
rect 53807 21659 55727 23579
rect 56407 21659 58327 23579
rect 59007 21659 60927 23579
rect 61607 21659 63527 23579
rect 64204 21660 64524 23580
rect -1190 19160 -870 21080
rect -193 19159 1727 21079
rect 2407 19159 4327 21079
rect 5007 19159 6927 21079
rect 7607 19159 9527 21079
rect 10204 19160 10524 21080
rect 37403 20566 39723 20886
rect 40186 20566 41706 20886
rect 42574 20568 44094 20888
rect 44682 20568 46202 20888
rect 46968 20568 48488 20888
rect 48951 20568 51271 20888
rect -1190 16660 -870 18580
rect -193 16659 1727 18579
rect 2407 16659 4327 18579
rect 5007 16659 6927 18579
rect 7607 16659 9527 18579
rect 10204 16660 10524 18580
rect 37420 17914 37740 19434
rect 38266 17914 39786 19434
rect 40296 17914 41816 19434
rect 42456 17914 43976 19434
rect 44496 17914 46016 19434
rect 46652 17914 48172 19434
rect 48692 17914 50212 19434
rect 50932 17914 51252 19434
rect 52810 19160 53130 21080
rect 53807 19159 55727 21079
rect 56407 19159 58327 21079
rect 59007 19159 60927 21079
rect 61607 19159 63527 21079
rect 64204 19160 64524 21080
rect -1192 15762 -872 16082
rect -194 15761 1726 16081
rect 2406 15761 4326 16081
rect 5006 15761 6926 16081
rect 7606 15761 9526 16081
rect 10206 15762 10526 16082
rect 37420 15810 37740 17330
rect 38266 15814 39786 17334
rect 40296 15814 41816 17334
rect 42456 15814 43976 17334
rect 44496 15814 46016 17334
rect 46652 15814 48172 17334
rect 48692 15814 50212 17334
rect 50932 15810 51252 17330
rect 52810 16660 53130 18580
rect 53807 16659 55727 18579
rect 56407 16659 58327 18579
rect 59007 16659 60927 18579
rect 61607 16659 63527 18579
rect 64204 16660 64524 18580
rect 52808 15762 53128 16082
rect 53806 15761 55726 16081
rect 56406 15761 58326 16081
rect 59006 15761 60926 16081
rect 61606 15761 63526 16081
rect 64206 15762 64526 16082
rect 37403 14406 39723 14726
rect 40186 14406 41706 14726
rect 42574 14408 44094 14728
rect 44856 14408 46376 14728
rect 46968 14408 48488 14728
rect 48951 14408 51271 14728
rect -12203 13538 -9883 13858
rect -9420 13538 -7900 13858
rect -7032 13540 -5512 13860
rect -5049 13540 -2729 13860
rect -12334 11124 -12014 12644
rect -11488 11124 -9968 12644
rect -9458 11124 -7938 12644
rect -7298 11124 -5778 12644
rect -5258 11124 -3738 12644
rect -3068 11126 -2748 12646
rect 37272 11792 37592 13312
rect 38118 11792 39638 13312
rect 40148 11792 41668 13312
rect 42308 11792 43828 13312
rect 44348 11792 45868 13312
rect 46538 11794 46858 13314
rect -12334 9020 -12014 10540
rect -11488 9024 -9968 10544
rect -9458 9024 -7938 10544
rect -7298 9024 -5778 10544
rect -5258 9024 -3738 10544
rect -3068 9022 -2748 10542
rect 37272 9688 37592 11208
rect 38118 9692 39638 11212
rect 40148 9692 41668 11212
rect 42308 9692 43828 11212
rect 44348 9692 45868 11212
rect 46538 9690 46858 11210
rect 37403 8470 39723 8790
rect 40186 8470 41706 8790
rect 42574 8472 44094 8792
rect 44557 8472 46877 8792
rect -12203 7802 -9883 8122
rect -9420 7802 -7900 8122
rect -7032 7804 -5512 8124
rect -5049 7804 -2729 8124
rect -12203 6338 -9883 6658
rect -9420 6338 -7900 6658
rect -7032 6340 -5512 6660
rect -5049 6340 -2729 6660
rect 37421 6604 39741 6924
rect 40204 6604 41724 6924
rect 42592 6606 44112 6926
rect 44575 6606 46895 6926
rect -12334 3924 -12014 5444
rect -11488 3924 -9968 5444
rect -9458 3924 -7938 5444
rect -7298 3924 -5778 5444
rect -5258 3924 -3738 5444
rect -3068 3926 -2748 5446
rect 37290 4190 37610 5710
rect 38136 4190 39656 5710
rect 40166 4190 41686 5710
rect 42326 4190 43846 5710
rect 44366 4190 45886 5710
rect 46556 4192 46876 5712
rect -12334 1820 -12014 3340
rect -11488 1824 -9968 3344
rect -9458 1824 -7938 3344
rect -7298 1824 -5778 3344
rect -5258 1824 -3738 3344
rect -3068 1822 -2748 3342
rect 37290 2086 37610 3606
rect 38136 2090 39656 3610
rect 40166 2090 41686 3610
rect 42326 2090 43846 3610
rect 44366 2090 45886 3610
rect 46556 2088 46876 3608
rect -12203 602 -9883 922
rect -9420 602 -7900 922
rect -7032 604 -5512 924
rect -5049 604 -2729 924
rect 37421 868 39741 1188
rect 40204 868 41724 1188
rect 42592 870 44112 1190
rect 44575 870 46895 1190
<< metal4 >>
rect -1450 28156 89950 28340
rect -1450 27856 11434 28156
rect 12034 27856 35066 28156
rect 35666 27856 65434 28156
rect 66034 27856 89066 28156
rect 89666 27856 89950 28156
rect -1450 27774 89950 27856
rect -1450 27647 15011 27774
rect -1450 27583 -1419 27647
rect -1349 27583 15011 27647
rect -1450 27560 15011 27583
rect 31796 27680 69011 27774
rect 31796 27564 47824 27680
rect 48462 27564 69011 27680
rect 31796 27560 69011 27564
rect 85796 27560 89950 27774
rect -1450 27540 89950 27560
rect -729 27092 -633 27108
rect -1189 26980 -867 26981
rect -1189 26660 -1188 26980
rect -868 26866 -867 26980
rect -729 26866 -713 27092
rect -868 26766 -713 26866
rect -868 26660 -867 26766
rect -1189 26659 -867 26660
rect -1082 26081 -982 26659
rect -730 26548 -713 26766
rect -649 26866 -633 27092
rect 1865 27093 1961 27109
rect -195 26981 1727 26982
rect -195 26866 -194 26981
rect -649 26766 -194 26866
rect -649 26548 -630 26766
rect -195 26661 -194 26766
rect 1726 26866 1727 26981
rect 1865 26866 1881 27093
rect 1726 26766 1881 26866
rect 1726 26661 1727 26766
rect -195 26660 1727 26661
rect -730 26208 -630 26548
rect 1865 26549 1881 26766
rect 1945 26866 1961 27093
rect 4465 27093 4561 27109
rect 2405 26981 4327 26982
rect 2405 26866 2406 26981
rect 1945 26766 2406 26866
rect 1945 26549 1961 26766
rect 2405 26661 2406 26766
rect 4326 26866 4327 26981
rect 4465 26866 4481 27093
rect 4326 26766 4481 26866
rect 4326 26661 4327 26766
rect 2405 26660 4327 26661
rect 1865 26533 1961 26549
rect 4465 26549 4481 26766
rect 4545 26866 4561 27093
rect 7065 27093 7161 27109
rect 5005 26981 6927 26982
rect 5005 26866 5006 26981
rect 4545 26766 5006 26866
rect 4545 26549 4561 26766
rect 5005 26661 5006 26766
rect 6926 26866 6927 26981
rect 7065 26866 7081 27093
rect 6926 26766 7081 26866
rect 6926 26661 6927 26766
rect 5005 26660 6927 26661
rect 4465 26533 4561 26549
rect 7065 26549 7081 26766
rect 7145 26866 7161 27093
rect 9665 27093 9761 27109
rect 7605 26981 9527 26982
rect 7605 26866 7606 26981
rect 7145 26766 7606 26866
rect 7145 26549 7161 26766
rect 7605 26661 7606 26766
rect 9526 26866 9527 26981
rect 9665 26866 9681 27093
rect 9526 26766 9681 26866
rect 9526 26661 9527 26766
rect 7605 26660 9527 26661
rect 7065 26533 7161 26549
rect 9665 26549 9681 26766
rect 9745 26866 9761 27093
rect 10665 27092 10761 27108
rect 10205 26980 10527 26981
rect 10205 26866 10206 26980
rect 9745 26766 10206 26866
rect 9745 26549 9761 26766
rect 10205 26660 10206 26766
rect 10526 26866 10527 26980
rect 10665 26866 10681 27092
rect 10526 26766 10681 26866
rect 10526 26660 10527 26766
rect 10205 26659 10527 26660
rect 9665 26533 9761 26549
rect -731 26192 -630 26208
rect -1191 26080 -869 26081
rect -1191 24160 -1190 26080
rect -870 24160 -869 26080
rect -1191 24159 -869 24160
rect -1082 23581 -982 24159
rect -731 24048 -715 26192
rect -651 24048 -630 26192
rect 720 26320 9958 26420
rect 720 26081 820 26320
rect 1866 26192 1962 26208
rect -194 26080 1728 26081
rect -194 24160 -193 26080
rect 1727 24160 1728 26080
rect -194 24159 1728 24160
rect -731 24032 -630 24048
rect 1866 24048 1882 26192
rect 1946 24048 1962 26192
rect 4466 26192 4562 26208
rect 2406 26080 4328 26081
rect 2406 24160 2407 26080
rect 4327 24160 4328 26080
rect 2406 24159 4328 24160
rect 1866 24032 1962 24048
rect -730 23708 -630 24032
rect 3342 23918 3442 24159
rect 4466 24048 4482 26192
rect 4546 24048 4562 26192
rect 5950 26081 6050 26320
rect 7066 26192 7162 26208
rect 5006 26080 6928 26081
rect 5006 24160 5007 26080
rect 6927 24160 6928 26080
rect 5006 24159 6928 24160
rect 4466 24032 4562 24048
rect 7066 24048 7082 26192
rect 7146 24048 7162 26192
rect 9666 26192 9762 26208
rect 7606 26080 9528 26081
rect 7606 24160 7607 26080
rect 9527 24160 9528 26080
rect 7606 24159 9528 24160
rect 7066 24032 7162 24048
rect 8526 23918 8626 24159
rect 9666 24048 9682 26192
rect 9746 24048 9762 26192
rect 9666 24032 9762 24048
rect -731 23692 -630 23708
rect -1191 23580 -869 23581
rect -1191 21660 -1190 23580
rect -870 21660 -869 23580
rect -1191 21659 -869 21660
rect -1082 21081 -982 21659
rect -731 21548 -715 23692
rect -651 21548 -630 23692
rect -731 21532 -630 21548
rect -730 21208 -630 21532
rect -731 21192 -630 21208
rect -1191 21080 -869 21081
rect -1191 19160 -1190 21080
rect -870 19160 -869 21080
rect -1191 19159 -869 19160
rect -1082 18581 -982 19159
rect -731 19048 -715 21192
rect -651 19048 -630 21192
rect -731 19032 -630 19048
rect -730 18708 -630 19032
rect -528 23818 8626 23918
rect -528 18918 -428 23818
rect 712 23580 812 23818
rect 1866 23691 1962 23707
rect -194 23579 1728 23580
rect -194 21659 -193 23579
rect 1727 21659 1728 23579
rect -194 21658 1728 21659
rect 1866 21547 1882 23691
rect 1946 21547 1962 23691
rect 4466 23691 4562 23707
rect 2406 23579 4328 23580
rect 2406 21659 2407 23579
rect 4327 21659 4328 23579
rect 2406 21658 4328 21659
rect 1866 21531 1962 21547
rect 3328 21418 3428 21658
rect 4466 21547 4482 23691
rect 4546 21547 4562 23691
rect 5950 23580 6050 23818
rect 7066 23691 7162 23707
rect 5006 23579 6928 23580
rect 5006 21659 5007 23579
rect 6927 21659 6928 23579
rect 5006 21658 6928 21659
rect 4466 21531 4562 21547
rect 7066 21547 7082 23691
rect 7146 21547 7162 23691
rect 9666 23691 9762 23707
rect 7606 23579 9528 23580
rect 7606 21659 7607 23579
rect 9527 21659 9528 23579
rect 7606 21658 9528 21659
rect 7066 21531 7162 21547
rect 8518 21418 8618 21658
rect 9666 21547 9682 23691
rect 9746 21547 9762 23691
rect 9666 21531 9762 21547
rect 9858 21418 9958 26320
rect 10314 26081 10414 26659
rect 10664 26548 10681 26766
rect 10745 26866 10761 27092
rect 53271 27092 53367 27108
rect 52811 26980 53133 26981
rect 10745 26548 10764 26866
rect 52811 26660 52812 26980
rect 53132 26866 53133 26980
rect 53271 26866 53287 27092
rect 53132 26766 53287 26866
rect 53132 26660 53133 26766
rect 52811 26659 53133 26660
rect 10664 26208 10764 26548
rect 38429 26568 38579 26569
rect 38429 26420 38430 26568
rect 38578 26420 38579 26568
rect 38429 26419 38579 26420
rect 41347 26568 41507 26569
rect 38430 26341 38578 26419
rect 41347 26410 41348 26568
rect 41506 26410 41507 26568
rect 41347 26409 41507 26410
rect 41348 26341 41506 26409
rect 10663 26192 10764 26208
rect 10203 26080 10525 26081
rect 10203 24160 10204 26080
rect 10524 24160 10525 26080
rect 10203 24159 10525 24160
rect 10314 23581 10414 24159
rect 10663 24048 10679 26192
rect 10743 24048 10764 26192
rect 37289 26340 39611 26341
rect 37289 26020 37290 26340
rect 39610 26020 39611 26340
rect 37289 26019 39611 26020
rect 40289 26340 42611 26341
rect 40289 26020 40290 26340
rect 42610 26020 42611 26340
rect 52918 26081 53018 26659
rect 53270 26548 53287 26766
rect 53351 26866 53367 27092
rect 55865 27093 55961 27109
rect 53805 26981 55727 26982
rect 53805 26866 53806 26981
rect 53351 26766 53806 26866
rect 53351 26548 53370 26766
rect 53805 26661 53806 26766
rect 55726 26866 55727 26981
rect 55865 26866 55881 27093
rect 55726 26766 55881 26866
rect 55726 26661 55727 26766
rect 53805 26660 55727 26661
rect 53270 26208 53370 26548
rect 55865 26549 55881 26766
rect 55945 26866 55961 27093
rect 58465 27093 58561 27109
rect 56405 26981 58327 26982
rect 56405 26866 56406 26981
rect 55945 26766 56406 26866
rect 55945 26549 55961 26766
rect 56405 26661 56406 26766
rect 58326 26866 58327 26981
rect 58465 26866 58481 27093
rect 58326 26766 58481 26866
rect 58326 26661 58327 26766
rect 56405 26660 58327 26661
rect 55865 26533 55961 26549
rect 58465 26549 58481 26766
rect 58545 26866 58561 27093
rect 61065 27093 61161 27109
rect 59005 26981 60927 26982
rect 59005 26866 59006 26981
rect 58545 26766 59006 26866
rect 58545 26549 58561 26766
rect 59005 26661 59006 26766
rect 60926 26866 60927 26981
rect 61065 26866 61081 27093
rect 60926 26766 61081 26866
rect 60926 26661 60927 26766
rect 59005 26660 60927 26661
rect 58465 26533 58561 26549
rect 61065 26549 61081 26766
rect 61145 26866 61161 27093
rect 63665 27093 63761 27109
rect 61605 26981 63527 26982
rect 61605 26866 61606 26981
rect 61145 26766 61606 26866
rect 61145 26549 61161 26766
rect 61605 26661 61606 26766
rect 63526 26866 63527 26981
rect 63665 26866 63681 27093
rect 63526 26766 63681 26866
rect 63526 26661 63527 26766
rect 61605 26660 63527 26661
rect 61065 26533 61161 26549
rect 63665 26549 63681 26766
rect 63745 26866 63761 27093
rect 64665 27092 64761 27108
rect 64205 26980 64527 26981
rect 64205 26866 64206 26980
rect 63745 26766 64206 26866
rect 63745 26549 63761 26766
rect 64205 26660 64206 26766
rect 64526 26866 64527 26980
rect 64665 26866 64681 27092
rect 64526 26766 64681 26866
rect 64526 26660 64527 26766
rect 64205 26659 64527 26660
rect 63665 26533 63761 26549
rect 53269 26192 53370 26208
rect 40289 26019 42611 26020
rect 52809 26080 53131 26081
rect 39530 25634 46676 25734
rect 37305 25476 37627 25477
rect 37049 24776 37183 24777
rect 37305 24776 37306 25476
rect 37049 24644 37050 24776
rect 37182 24644 37306 24776
rect 37049 24643 37183 24644
rect 10663 24032 10764 24048
rect 10664 23708 10764 24032
rect 37305 23956 37306 24644
rect 37626 23956 37627 25476
rect 39530 25473 39630 25634
rect 37305 23955 37627 23956
rect 38157 25472 39679 25473
rect 38157 23952 38158 25472
rect 39678 23952 39679 25472
rect 38157 23951 39679 23952
rect 40187 25472 41709 25473
rect 40187 23952 40188 25472
rect 41708 24714 41709 25472
rect 41708 24614 41928 24714
rect 41708 23952 41709 24614
rect 40187 23951 41709 23952
rect 10663 23692 10764 23708
rect 10203 23580 10525 23581
rect 10203 21660 10204 23580
rect 10524 21660 10525 23580
rect 10203 21659 10525 21660
rect 704 21318 9958 21418
rect 704 21080 804 21318
rect 1866 21191 1962 21207
rect -194 21079 1728 21080
rect -194 19159 -193 21079
rect 1727 19159 1728 21079
rect -194 19158 1728 19159
rect 1866 19047 1882 21191
rect 1946 19047 1962 21191
rect 4466 21191 4562 21207
rect 2406 21079 4328 21080
rect 2406 19159 2407 21079
rect 4327 19159 4328 21079
rect 2406 19158 4328 19159
rect 1866 19031 1962 19047
rect 3320 18918 3420 19158
rect 4466 19047 4482 21191
rect 4546 19047 4562 21191
rect 5942 21080 6042 21318
rect 7066 21191 7162 21207
rect 5006 21079 6928 21080
rect 5006 19159 5007 21079
rect 6927 19159 6928 21079
rect 5006 19158 6928 19159
rect 4466 19031 4562 19047
rect 7066 19047 7082 21191
rect 7146 19047 7162 21191
rect 9666 21191 9762 21207
rect 7606 21079 9528 21080
rect 7606 19159 7607 21079
rect 9527 19159 9528 21079
rect 7606 19158 9528 19159
rect 7066 19031 7162 19047
rect 8510 18918 8610 19158
rect 9666 19047 9682 21191
rect 9746 19047 9762 21191
rect 9666 19031 9762 19047
rect -528 18917 9300 18918
rect -528 18819 9201 18917
rect 9299 18819 9300 18917
rect -528 18818 9300 18819
rect -731 18692 -630 18708
rect -1191 18580 -869 18581
rect -1191 16660 -1190 18580
rect -870 16660 -869 18580
rect -1191 16659 -869 16660
rect -1082 16083 -982 16659
rect -731 16548 -715 18692
rect -651 16548 -630 18692
rect 696 18580 796 18818
rect 1866 18691 1962 18707
rect -194 18579 1728 18580
rect -194 16659 -193 18579
rect 1727 16659 1728 18579
rect -194 16658 1728 16659
rect -731 16532 -630 16548
rect -730 16210 -630 16532
rect 1866 16547 1882 18691
rect 1946 16547 1962 18691
rect 4466 18691 4562 18707
rect 2406 18579 4328 18580
rect 2406 16659 2407 18579
rect 4327 16659 4328 18579
rect 2406 16658 4328 16659
rect 1866 16531 1962 16547
rect 3304 16422 3404 16658
rect 4466 16547 4482 18691
rect 4546 16547 4562 18691
rect 5942 18580 6042 18818
rect 7066 18691 7162 18707
rect 5006 18579 6928 18580
rect 5006 16659 5007 18579
rect 6927 16659 6928 18579
rect 5006 16658 6928 16659
rect 4466 16531 4562 16547
rect 7066 16547 7082 18691
rect 7146 16547 7162 18691
rect 9666 18691 9762 18707
rect 7606 18579 9528 18580
rect 7606 16659 7607 18579
rect 9527 16659 9528 18579
rect 7606 16658 9528 16659
rect 7066 16531 7162 16547
rect 8510 16422 8610 16658
rect 9666 16547 9682 18691
rect 9746 16547 9762 18691
rect 9666 16531 9762 16547
rect 9858 16422 9958 21318
rect 10314 21081 10414 21659
rect 10663 21548 10679 23692
rect 10743 21548 10764 23692
rect 40401 23870 40503 23871
rect 40401 23770 40402 23870
rect 40502 23770 40503 23870
rect 36467 23570 36569 23571
rect 36467 23568 36468 23570
rect 36462 23470 36468 23568
rect 36568 23568 36569 23570
rect 40401 23568 40503 23770
rect 36568 23567 40503 23568
rect 36568 23470 39493 23567
rect 36462 23469 39493 23470
rect 39591 23469 40503 23567
rect 36462 23468 40503 23469
rect 40401 23467 40503 23468
rect 41562 23711 41662 23712
rect 41562 23613 41563 23711
rect 41661 23613 41662 23711
rect 41562 23373 41662 23613
rect 37305 23372 37627 23373
rect 37075 22676 37197 22677
rect 37305 22676 37306 23372
rect 37075 22556 37076 22676
rect 37196 22556 37306 22676
rect 37075 22555 37197 22556
rect 37305 21852 37306 22556
rect 37626 21852 37627 23372
rect 37305 21851 37627 21852
rect 38157 23372 39679 23373
rect 38157 21852 38158 23372
rect 39678 21852 39679 23372
rect 38157 21851 39679 21852
rect 40187 23372 41709 23373
rect 40187 21852 40188 23372
rect 41708 21852 41709 23372
rect 40187 21851 41709 21852
rect 39512 21694 39612 21851
rect 41828 21694 41928 24614
rect 42030 23714 42130 25634
rect 42405 25476 42727 25477
rect 42405 23956 42406 25476
rect 42726 24768 42727 25476
rect 42911 24768 43049 24769
rect 42726 24632 42912 24768
rect 43048 24632 43049 24768
rect 42726 23956 42727 24632
rect 42911 24631 43049 24632
rect 46576 24535 46676 25634
rect 46575 24534 46677 24535
rect 46575 24434 46576 24534
rect 46676 24434 46677 24534
rect 46575 24433 46677 24434
rect 52809 24160 52810 26080
rect 53130 24160 53131 26080
rect 52809 24159 53131 24160
rect 42405 23955 42727 23956
rect 52143 23714 52245 23715
rect 42030 23713 52144 23714
rect 42029 23712 52144 23713
rect 42029 23612 42030 23712
rect 42130 23614 52144 23712
rect 52244 23614 52245 23714
rect 42130 23612 42131 23614
rect 52143 23613 52245 23614
rect 42029 23611 42131 23612
rect 52918 23581 53018 24159
rect 53269 24048 53285 26192
rect 53349 24048 53370 26192
rect 54720 26320 63958 26420
rect 54720 26081 54820 26320
rect 55866 26192 55962 26208
rect 53806 26080 55728 26081
rect 53806 24160 53807 26080
rect 55727 24160 55728 26080
rect 53806 24159 55728 24160
rect 53269 24032 53370 24048
rect 55866 24048 55882 26192
rect 55946 24048 55962 26192
rect 58466 26192 58562 26208
rect 56406 26080 58328 26081
rect 56406 24160 56407 26080
rect 58327 24160 58328 26080
rect 56406 24159 58328 24160
rect 55866 24032 55962 24048
rect 53270 23708 53370 24032
rect 57342 23918 57442 24159
rect 58466 24048 58482 26192
rect 58546 24048 58562 26192
rect 59950 26081 60050 26320
rect 61066 26192 61162 26208
rect 59006 26080 60928 26081
rect 59006 24160 59007 26080
rect 60927 24160 60928 26080
rect 59006 24159 60928 24160
rect 58466 24032 58562 24048
rect 61066 24048 61082 26192
rect 61146 24048 61162 26192
rect 63666 26192 63762 26208
rect 61606 26080 63528 26081
rect 61606 24160 61607 26080
rect 63527 24160 63528 26080
rect 61606 24159 63528 24160
rect 61066 24032 61162 24048
rect 62526 23918 62626 24159
rect 63666 24048 63682 26192
rect 63746 24048 63762 26192
rect 63666 24032 63762 24048
rect 53269 23692 53370 23708
rect 52809 23580 53131 23581
rect 42405 23372 42727 23373
rect 42405 21852 42406 23372
rect 42726 22658 42727 23372
rect 42863 22658 43005 22659
rect 42726 22518 42864 22658
rect 43004 22518 43005 22658
rect 42726 21852 42727 22518
rect 42863 22517 43005 22518
rect 42405 21851 42727 21852
rect 49759 21700 49861 21701
rect 49759 21694 49760 21700
rect 39512 21600 49760 21694
rect 49860 21694 49861 21700
rect 52380 21694 52480 21696
rect 49860 21600 52480 21694
rect 52809 21660 52810 23580
rect 53130 21660 53131 23580
rect 52809 21659 53131 21660
rect 39512 21594 52480 21600
rect 10663 21532 10764 21548
rect 10664 21208 10764 21532
rect 10663 21192 10764 21208
rect 10203 21080 10525 21081
rect 10203 19160 10204 21080
rect 10524 19160 10525 21080
rect 10203 19159 10525 19160
rect 10314 18581 10414 19159
rect 10663 19048 10679 21192
rect 10743 19048 10764 21192
rect 46404 21381 46504 21382
rect 46404 21283 46405 21381
rect 46503 21283 46504 21381
rect 42573 20888 44095 20889
rect 37402 20886 39724 20887
rect 37402 20566 37403 20886
rect 39723 20566 39724 20886
rect 37402 20565 39724 20566
rect 40185 20886 41707 20887
rect 40185 20566 40186 20886
rect 41706 20566 41707 20886
rect 42573 20568 42574 20888
rect 44094 20568 44095 20888
rect 42573 20567 44095 20568
rect 44681 20888 46203 20889
rect 44681 20568 44682 20888
rect 46202 20568 46203 20888
rect 44681 20567 46203 20568
rect 40185 20565 41707 20566
rect 38494 20491 38672 20565
rect 40894 20491 41072 20565
rect 43294 20491 43472 20567
rect 45420 20491 45598 20567
rect 38493 20490 38673 20491
rect 38493 20312 38494 20490
rect 38672 20312 38673 20490
rect 38493 20311 38673 20312
rect 40893 20490 41073 20491
rect 40893 20312 40894 20490
rect 41072 20312 41073 20490
rect 40893 20311 41073 20312
rect 43293 20490 43473 20491
rect 43293 20312 43294 20490
rect 43472 20312 43473 20490
rect 43293 20311 43473 20312
rect 45419 20490 45599 20491
rect 45419 20312 45420 20490
rect 45598 20312 45599 20490
rect 45419 20311 45599 20312
rect 39077 19926 39179 19927
rect 36472 19925 39078 19926
rect 36472 19827 36473 19925
rect 36571 19827 39078 19925
rect 36472 19826 39078 19827
rect 39178 19826 39179 19926
rect 39077 19825 39179 19826
rect 46404 19700 46504 21283
rect 51793 21066 51895 21067
rect 51793 20966 51794 21066
rect 51894 20966 52248 21066
rect 51793 20965 51895 20966
rect 46967 20888 48489 20889
rect 46967 20568 46968 20888
rect 48488 20568 48489 20888
rect 46967 20567 48489 20568
rect 48950 20888 51272 20889
rect 48950 20568 48951 20888
rect 51271 20568 51272 20888
rect 48950 20567 51272 20568
rect 47594 20491 47772 20567
rect 49994 20491 50172 20567
rect 47593 20490 47773 20491
rect 47593 20312 47594 20490
rect 47772 20312 47773 20490
rect 47593 20311 47773 20312
rect 49993 20490 50173 20491
rect 49993 20312 49994 20490
rect 50172 20312 50173 20490
rect 49993 20311 50173 20312
rect 39640 19600 50704 19700
rect 39640 19435 39740 19600
rect 10663 19032 10764 19048
rect 10664 18708 10764 19032
rect 37419 19434 37741 19435
rect 10663 18692 10764 18708
rect 10203 18580 10525 18581
rect 10203 16660 10204 18580
rect 10524 16660 10525 18580
rect 10203 16659 10525 16660
rect 3304 16421 9960 16422
rect 3304 16323 9861 16421
rect 9959 16323 9960 16421
rect 3304 16322 9960 16323
rect -733 16194 -630 16210
rect -1193 16082 -871 16083
rect -1193 15762 -1192 16082
rect -872 15974 -871 16082
rect -733 15974 -717 16194
rect -872 15874 -717 15974
rect -872 15762 -871 15874
rect -1193 15761 -871 15762
rect -733 15650 -717 15874
rect -653 15974 -630 16194
rect 1865 16193 1961 16209
rect -195 16081 1727 16082
rect -195 15974 -194 16081
rect -653 15874 -194 15974
rect -653 15872 -630 15874
rect -653 15650 -637 15872
rect -195 15761 -194 15874
rect 1726 15974 1727 16081
rect 1865 15974 1881 16193
rect 1726 15874 1881 15974
rect 1726 15761 1727 15874
rect -195 15760 1727 15761
rect -733 15634 -637 15650
rect 1865 15649 1881 15874
rect 1945 15974 1961 16193
rect 4465 16193 4561 16209
rect 2405 16081 4327 16082
rect 2405 15974 2406 16081
rect 1945 15874 2406 15974
rect 1945 15649 1961 15874
rect 2405 15761 2406 15874
rect 4326 15974 4327 16081
rect 4465 15974 4481 16193
rect 4326 15874 4481 15974
rect 4326 15761 4327 15874
rect 2405 15760 4327 15761
rect 1865 15633 1961 15649
rect 4465 15649 4481 15874
rect 4545 15974 4561 16193
rect 7065 16193 7161 16209
rect 5005 16081 6927 16082
rect 5005 15974 5006 16081
rect 4545 15874 5006 15974
rect 4545 15649 4561 15874
rect 5005 15761 5006 15874
rect 6926 15974 6927 16081
rect 7065 15974 7081 16193
rect 6926 15874 7081 15974
rect 6926 15761 6927 15874
rect 5005 15760 6927 15761
rect 4465 15633 4561 15649
rect 7065 15649 7081 15874
rect 7145 15974 7161 16193
rect 9665 16193 9761 16209
rect 7605 16081 9527 16082
rect 7605 15974 7606 16081
rect 7145 15874 7606 15974
rect 7145 15649 7161 15874
rect 7605 15761 7606 15874
rect 9526 15974 9527 16081
rect 9665 15974 9681 16193
rect 9526 15874 9681 15974
rect 9526 15761 9527 15874
rect 7605 15760 9527 15761
rect 7065 15633 7161 15649
rect 9665 15649 9681 15874
rect 9745 15974 9761 16193
rect 10314 16083 10414 16659
rect 10663 16548 10679 18692
rect 10743 16548 10764 18692
rect 37149 18790 37359 18791
rect 37419 18790 37420 19434
rect 37149 18582 37150 18790
rect 37358 18582 37420 18790
rect 37149 18581 37359 18582
rect 37419 17914 37420 18582
rect 37740 17914 37741 19434
rect 37419 17913 37741 17914
rect 38265 19434 39787 19435
rect 38265 17914 38266 19434
rect 39786 17914 39787 19434
rect 38265 17913 39787 17914
rect 40295 19434 41817 19435
rect 40295 17914 40296 19434
rect 41816 18680 41817 19434
rect 41816 18580 42068 18680
rect 41816 17914 41817 18580
rect 40295 17913 41817 17914
rect 40416 17829 40516 17830
rect 40416 17731 40417 17829
rect 40515 17731 40516 17829
rect 40416 17524 40516 17731
rect 39618 17523 40516 17524
rect 39618 17425 39619 17523
rect 39717 17425 40516 17523
rect 39618 17424 40516 17425
rect 41672 17677 41772 17678
rect 41672 17579 41673 17677
rect 41771 17579 41772 17677
rect 41672 17335 41772 17579
rect 38265 17334 39787 17335
rect 37419 17330 37741 17331
rect 10663 16532 10764 16548
rect 10664 16194 10764 16532
rect 37078 16650 37266 16651
rect 37419 16650 37420 17330
rect 37078 16464 37079 16650
rect 37265 16464 37420 16650
rect 37078 16463 37266 16464
rect 10205 16082 10527 16083
rect 10205 15974 10206 16082
rect 9745 15874 10206 15974
rect 9745 15649 9761 15874
rect 10205 15762 10206 15874
rect 10526 15974 10527 16082
rect 10664 15974 10681 16194
rect 10526 15874 10681 15974
rect 10526 15762 10527 15874
rect 10664 15872 10681 15874
rect 10205 15761 10527 15762
rect 9665 15633 9761 15649
rect 10665 15650 10681 15872
rect 10745 15872 10764 16194
rect 10745 15650 10761 15872
rect 37419 15810 37420 16464
rect 37740 15810 37741 17330
rect 38265 15814 38266 17334
rect 39786 15814 39787 17334
rect 38265 15813 39787 15814
rect 40295 17334 41817 17335
rect 40295 15814 40296 17334
rect 41816 15814 41817 17334
rect 40295 15813 41817 15814
rect 37419 15809 37741 15810
rect 10665 15634 10761 15650
rect 39622 15660 39722 15813
rect 41968 15660 42068 18580
rect 42204 17679 42304 19600
rect 43840 19435 43940 19600
rect 42455 19434 43977 19435
rect 42455 17914 42456 19434
rect 43976 17914 43977 19434
rect 42455 17913 43977 17914
rect 44495 19434 46017 19435
rect 44495 17914 44496 19434
rect 46016 18680 46017 19434
rect 46016 18580 46268 18680
rect 46016 17914 46017 18580
rect 44495 17913 46017 17914
rect 44642 17817 44742 17818
rect 44642 17719 44643 17817
rect 44741 17719 44742 17817
rect 42203 17678 42305 17679
rect 42203 17578 42204 17678
rect 42304 17578 42305 17678
rect 42203 17577 42305 17578
rect 44642 17524 44742 17719
rect 43818 17523 44742 17524
rect 43818 17425 43819 17523
rect 43917 17425 44742 17523
rect 43818 17424 44742 17425
rect 45872 17677 45972 17678
rect 45872 17579 45873 17677
rect 45971 17579 45972 17677
rect 45872 17335 45972 17579
rect 42455 17334 43977 17335
rect 42455 15814 42456 17334
rect 43976 15814 43977 17334
rect 42455 15813 43977 15814
rect 44495 17334 46017 17335
rect 44495 15814 44496 17334
rect 46016 15814 46017 17334
rect 44495 15813 46017 15814
rect 43822 15660 43922 15813
rect 46168 15660 46268 18580
rect 46404 17679 46504 19600
rect 48040 19435 48140 19600
rect 46651 19434 48173 19435
rect 46651 17914 46652 19434
rect 48172 17914 48173 19434
rect 46651 17913 48173 17914
rect 48691 19434 50213 19435
rect 48691 17914 48692 19434
rect 50212 18680 50213 19434
rect 50212 18580 50468 18680
rect 50212 17914 50213 18580
rect 48691 17913 50213 17914
rect 48764 17827 48864 17828
rect 48764 17729 48765 17827
rect 48863 17729 48864 17827
rect 46403 17678 46505 17679
rect 46403 17578 46404 17678
rect 46504 17578 46505 17678
rect 46403 17577 46505 17578
rect 48764 17522 48864 17729
rect 48018 17521 48864 17522
rect 48018 17423 48019 17521
rect 48117 17423 48864 17521
rect 48018 17422 48864 17423
rect 50072 17677 50172 17678
rect 50072 17579 50073 17677
rect 50171 17579 50172 17677
rect 50072 17335 50172 17579
rect 46651 17334 48173 17335
rect 46651 15814 46652 17334
rect 48172 15814 48173 17334
rect 46651 15813 48173 15814
rect 48691 17334 50213 17335
rect 48691 15814 48692 17334
rect 50212 15814 50213 17334
rect 48691 15813 50213 15814
rect 48022 15660 48122 15813
rect 50368 15660 50468 18580
rect 50604 17679 50704 19600
rect 50931 19434 51253 19435
rect 50931 17914 50932 19434
rect 51252 18732 51253 19434
rect 51337 18732 51501 18733
rect 51252 18570 51338 18732
rect 51500 18570 51501 18732
rect 51252 17914 51253 18570
rect 51337 18569 51501 18570
rect 50931 17913 51253 17914
rect 50603 17678 50705 17679
rect 50603 17578 50604 17678
rect 50704 17578 50705 17678
rect 50603 17577 50705 17578
rect 50931 17330 51253 17331
rect 50931 15810 50932 17330
rect 51252 16638 51253 17330
rect 51363 16638 51533 16639
rect 51252 16470 51364 16638
rect 51532 16470 51533 16638
rect 51252 15810 51253 16470
rect 51363 16469 51533 16470
rect 50931 15809 51253 15810
rect 52148 15660 52248 20966
rect 39622 15560 52248 15660
rect 39297 15376 39399 15377
rect 36254 15375 39298 15376
rect 36254 15277 36255 15375
rect 36353 15277 39298 15375
rect 36254 15276 39298 15277
rect 39398 15276 39399 15376
rect 39297 15275 39399 15276
rect 52380 15101 52480 21594
rect 52918 21081 53018 21659
rect 53269 21548 53285 23692
rect 53349 21548 53370 23692
rect 53269 21532 53370 21548
rect 53270 21208 53370 21532
rect 53269 21192 53370 21208
rect 52809 21080 53131 21081
rect 52809 19160 52810 21080
rect 53130 19160 53131 21080
rect 52809 19159 53131 19160
rect 52918 18581 53018 19159
rect 53269 19048 53285 21192
rect 53349 19048 53370 21192
rect 53269 19032 53370 19048
rect 53270 18708 53370 19032
rect 53472 23818 62626 23918
rect 53472 18918 53572 23818
rect 54712 23580 54812 23818
rect 55866 23691 55962 23707
rect 53806 23579 55728 23580
rect 53806 21659 53807 23579
rect 55727 21659 55728 23579
rect 53806 21658 55728 21659
rect 55866 21547 55882 23691
rect 55946 21547 55962 23691
rect 58466 23691 58562 23707
rect 56406 23579 58328 23580
rect 56406 21659 56407 23579
rect 58327 21659 58328 23579
rect 56406 21658 58328 21659
rect 55866 21531 55962 21547
rect 57328 21418 57428 21658
rect 58466 21547 58482 23691
rect 58546 21547 58562 23691
rect 59950 23580 60050 23818
rect 61066 23691 61162 23707
rect 59006 23579 60928 23580
rect 59006 21659 59007 23579
rect 60927 21659 60928 23579
rect 59006 21658 60928 21659
rect 58466 21531 58562 21547
rect 61066 21547 61082 23691
rect 61146 21547 61162 23691
rect 63666 23691 63762 23707
rect 61606 23579 63528 23580
rect 61606 21659 61607 23579
rect 63527 21659 63528 23579
rect 61606 21658 63528 21659
rect 61066 21531 61162 21547
rect 62518 21418 62618 21658
rect 63666 21547 63682 23691
rect 63746 21547 63762 23691
rect 63666 21531 63762 21547
rect 63858 21418 63958 26320
rect 64314 26081 64414 26659
rect 64664 26548 64681 26766
rect 64745 26866 64761 27092
rect 64745 26548 64764 26866
rect 64664 26208 64764 26548
rect 64663 26192 64764 26208
rect 64203 26080 64525 26081
rect 64203 24160 64204 26080
rect 64524 24160 64525 26080
rect 64203 24159 64525 24160
rect 64314 23581 64414 24159
rect 64663 24048 64679 26192
rect 64743 24048 64764 26192
rect 64663 24032 64764 24048
rect 64664 23708 64764 24032
rect 64663 23692 64764 23708
rect 64203 23580 64525 23581
rect 64203 21660 64204 23580
rect 64524 21660 64525 23580
rect 64203 21659 64525 21660
rect 54704 21318 63958 21418
rect 54704 21080 54804 21318
rect 55866 21191 55962 21207
rect 53806 21079 55728 21080
rect 53806 19159 53807 21079
rect 55727 19159 55728 21079
rect 53806 19158 55728 19159
rect 55866 19047 55882 21191
rect 55946 19047 55962 21191
rect 58466 21191 58562 21207
rect 56406 21079 58328 21080
rect 56406 19159 56407 21079
rect 58327 19159 58328 21079
rect 56406 19158 58328 19159
rect 55866 19031 55962 19047
rect 57320 18918 57420 19158
rect 58466 19047 58482 21191
rect 58546 19047 58562 21191
rect 59942 21080 60042 21318
rect 61066 21191 61162 21207
rect 59006 21079 60928 21080
rect 59006 19159 59007 21079
rect 60927 19159 60928 21079
rect 59006 19158 60928 19159
rect 58466 19031 58562 19047
rect 61066 19047 61082 21191
rect 61146 19047 61162 21191
rect 63666 21191 63762 21207
rect 61606 21079 63528 21080
rect 61606 19159 61607 21079
rect 63527 19159 63528 21079
rect 61606 19158 63528 19159
rect 61066 19031 61162 19047
rect 62510 18918 62610 19158
rect 63666 19047 63682 21191
rect 63746 19047 63762 21191
rect 63666 19031 63762 19047
rect 53472 18917 63300 18918
rect 53472 18819 63201 18917
rect 63299 18819 63300 18917
rect 53472 18818 63300 18819
rect 53269 18692 53370 18708
rect 52809 18580 53131 18581
rect 52809 16660 52810 18580
rect 53130 16660 53131 18580
rect 52809 16659 53131 16660
rect 52918 16083 53018 16659
rect 53269 16548 53285 18692
rect 53349 16548 53370 18692
rect 54696 18580 54796 18818
rect 55866 18691 55962 18707
rect 53806 18579 55728 18580
rect 53806 16659 53807 18579
rect 55727 16659 55728 18579
rect 53806 16658 55728 16659
rect 53269 16532 53370 16548
rect 53270 16210 53370 16532
rect 55866 16547 55882 18691
rect 55946 16547 55962 18691
rect 58466 18691 58562 18707
rect 56406 18579 58328 18580
rect 56406 16659 56407 18579
rect 58327 16659 58328 18579
rect 56406 16658 58328 16659
rect 55866 16531 55962 16547
rect 57304 16422 57404 16658
rect 58466 16547 58482 18691
rect 58546 16547 58562 18691
rect 59942 18580 60042 18818
rect 61066 18691 61162 18707
rect 59006 18579 60928 18580
rect 59006 16659 59007 18579
rect 60927 16659 60928 18579
rect 59006 16658 60928 16659
rect 58466 16531 58562 16547
rect 61066 16547 61082 18691
rect 61146 16547 61162 18691
rect 63666 18691 63762 18707
rect 61606 18579 63528 18580
rect 61606 16659 61607 18579
rect 63527 16659 63528 18579
rect 61606 16658 63528 16659
rect 61066 16531 61162 16547
rect 62510 16422 62610 16658
rect 63666 16547 63682 18691
rect 63746 16547 63762 18691
rect 63666 16531 63762 16547
rect 63858 16422 63958 21318
rect 64314 21081 64414 21659
rect 64663 21548 64679 23692
rect 64743 21548 64764 23692
rect 64663 21532 64764 21548
rect 64664 21208 64764 21532
rect 64663 21192 64764 21208
rect 64203 21080 64525 21081
rect 64203 19160 64204 21080
rect 64524 19160 64525 21080
rect 64203 19159 64525 19160
rect 64314 18581 64414 19159
rect 64663 19048 64679 21192
rect 64743 19048 64764 21192
rect 64663 19032 64764 19048
rect 64664 18708 64764 19032
rect 64663 18692 64764 18708
rect 64203 18580 64525 18581
rect 64203 16660 64204 18580
rect 64524 16660 64525 18580
rect 64203 16659 64525 16660
rect 57304 16421 63960 16422
rect 57304 16323 63861 16421
rect 63959 16323 63960 16421
rect 57304 16322 63960 16323
rect 53267 16194 53370 16210
rect 52807 16082 53129 16083
rect 52807 15762 52808 16082
rect 53128 15974 53129 16082
rect 53267 15974 53283 16194
rect 53128 15874 53283 15974
rect 53128 15762 53129 15874
rect 52807 15761 53129 15762
rect 53267 15650 53283 15874
rect 53347 15974 53370 16194
rect 55865 16193 55961 16209
rect 53805 16081 55727 16082
rect 53805 15974 53806 16081
rect 53347 15874 53806 15974
rect 53347 15872 53370 15874
rect 53347 15650 53363 15872
rect 53805 15761 53806 15874
rect 55726 15974 55727 16081
rect 55865 15974 55881 16193
rect 55726 15874 55881 15974
rect 55726 15761 55727 15874
rect 53805 15760 55727 15761
rect 53267 15634 53363 15650
rect 55865 15649 55881 15874
rect 55945 15974 55961 16193
rect 58465 16193 58561 16209
rect 56405 16081 58327 16082
rect 56405 15974 56406 16081
rect 55945 15874 56406 15974
rect 55945 15649 55961 15874
rect 56405 15761 56406 15874
rect 58326 15974 58327 16081
rect 58465 15974 58481 16193
rect 58326 15874 58481 15974
rect 58326 15761 58327 15874
rect 56405 15760 58327 15761
rect 55865 15633 55961 15649
rect 58465 15649 58481 15874
rect 58545 15974 58561 16193
rect 61065 16193 61161 16209
rect 59005 16081 60927 16082
rect 59005 15974 59006 16081
rect 58545 15874 59006 15974
rect 58545 15649 58561 15874
rect 59005 15761 59006 15874
rect 60926 15974 60927 16081
rect 61065 15974 61081 16193
rect 60926 15874 61081 15974
rect 60926 15761 60927 15874
rect 59005 15760 60927 15761
rect 58465 15633 58561 15649
rect 61065 15649 61081 15874
rect 61145 15974 61161 16193
rect 63665 16193 63761 16209
rect 61605 16081 63527 16082
rect 61605 15974 61606 16081
rect 61145 15874 61606 15974
rect 61145 15649 61161 15874
rect 61605 15761 61606 15874
rect 63526 15974 63527 16081
rect 63665 15974 63681 16193
rect 63526 15874 63681 15974
rect 63526 15761 63527 15874
rect 61605 15760 63527 15761
rect 61065 15633 61161 15649
rect 63665 15649 63681 15874
rect 63745 15974 63761 16193
rect 64314 16083 64414 16659
rect 64663 16548 64679 18692
rect 64743 16548 64764 18692
rect 64663 16532 64764 16548
rect 64664 16194 64764 16532
rect 64205 16082 64527 16083
rect 64205 15974 64206 16082
rect 63745 15874 64206 15974
rect 63745 15649 63761 15874
rect 64205 15762 64206 15874
rect 64526 15974 64527 16082
rect 64664 15974 64681 16194
rect 64526 15874 64681 15974
rect 64526 15762 64527 15874
rect 64664 15872 64681 15874
rect 64205 15761 64527 15762
rect 63665 15633 63761 15649
rect 64665 15650 64681 15872
rect 64745 15872 64764 16194
rect 64745 15650 64761 15872
rect 64665 15634 64761 15650
rect 52379 15100 52481 15101
rect 52379 15000 52380 15100
rect 52480 15000 52481 15100
rect 52379 14999 52481 15000
rect 42573 14728 44095 14729
rect 37402 14726 39724 14727
rect 37402 14406 37403 14726
rect 39723 14406 39724 14726
rect 37402 14405 39724 14406
rect 40185 14726 41707 14727
rect 40185 14406 40186 14726
rect 41706 14406 41707 14726
rect 42573 14408 42574 14728
rect 44094 14408 44095 14728
rect 42573 14407 44095 14408
rect 44855 14728 46377 14729
rect 44855 14408 44856 14728
rect 46376 14408 46377 14728
rect 44855 14407 46377 14408
rect 46967 14728 48489 14729
rect 46967 14408 46968 14728
rect 48488 14408 48489 14728
rect 46967 14407 48489 14408
rect 48950 14728 51272 14729
rect 48950 14408 48951 14728
rect 51271 14408 51272 14728
rect 48950 14407 51272 14408
rect 40185 14405 41707 14406
rect 38478 14317 38636 14405
rect 40890 14317 41048 14405
rect 43290 14317 43448 14407
rect 45690 14317 45848 14407
rect 47690 14317 47848 14407
rect 50090 14317 50248 14407
rect 38477 14316 38637 14317
rect -8837 14174 -8645 14175
rect -11155 14168 -11007 14169
rect -11155 14022 -11154 14168
rect -11008 14022 -11007 14168
rect -11155 14021 -11007 14022
rect -11154 13859 -11008 14021
rect -8837 13984 -8836 14174
rect -8646 13984 -8645 14174
rect -3941 14168 -3781 14169
rect -8837 13983 -8645 13984
rect -6347 14150 -6169 14151
rect -8836 13859 -8646 13983
rect -6347 13974 -6346 14150
rect -6170 13974 -6169 14150
rect -3941 14010 -3940 14168
rect -3782 14010 -3781 14168
rect 38477 14158 38478 14316
rect 38636 14158 38637 14316
rect 38477 14157 38637 14158
rect 40889 14316 41049 14317
rect 40889 14158 40890 14316
rect 41048 14158 41049 14316
rect 40889 14157 41049 14158
rect 43289 14316 43449 14317
rect 43289 14158 43290 14316
rect 43448 14158 43449 14316
rect 43289 14157 43449 14158
rect 45689 14316 45849 14317
rect 45689 14158 45690 14316
rect 45848 14158 45849 14316
rect 45689 14157 45849 14158
rect 47689 14316 47849 14317
rect 47689 14158 47690 14316
rect 47848 14158 47849 14316
rect 47689 14157 47849 14158
rect 50089 14316 50249 14317
rect 50089 14158 50090 14316
rect 50248 14158 50249 14316
rect 50089 14157 50249 14158
rect -3941 14009 -3781 14010
rect -6347 13973 -6169 13974
rect -6346 13861 -6170 13973
rect -3940 13861 -3782 14009
rect -7033 13860 -5511 13861
rect -12204 13858 -9882 13859
rect -12204 13538 -12203 13858
rect -9883 13538 -9882 13858
rect -12204 13537 -9882 13538
rect -9421 13858 -7899 13859
rect -9421 13538 -9420 13858
rect -7900 13538 -7899 13858
rect -7033 13540 -7032 13860
rect -5512 13540 -5511 13860
rect -7033 13539 -5511 13540
rect -5050 13860 -2728 13861
rect -5050 13540 -5049 13860
rect -2729 13540 -2728 13860
rect -5050 13539 -2728 13540
rect 36748 13581 46318 13582
rect -9421 13537 -7899 13538
rect 36748 13483 36749 13581
rect 36847 13483 46318 13581
rect 36748 13482 46318 13483
rect 39510 13313 39610 13482
rect 37271 13312 37593 13313
rect -10575 13138 -10473 13139
rect -13108 13137 -10574 13138
rect -13108 13039 -13107 13137
rect -13009 13039 -10574 13137
rect -13108 13038 -10574 13039
rect -10474 13038 -10473 13138
rect -10575 13037 -10473 13038
rect -2397 12904 -2295 12905
rect -10164 12804 -2396 12904
rect -2296 12804 -2295 12904
rect -10164 12645 -10064 12804
rect -12335 12644 -12013 12645
rect -12625 11974 -12529 11975
rect -12335 11974 -12334 12644
rect -12625 11880 -12624 11974
rect -12530 11880 -12334 11974
rect -12625 11879 -12529 11880
rect -12335 11124 -12334 11880
rect -12014 11124 -12013 12644
rect -12335 11123 -12013 11124
rect -11489 12644 -9967 12645
rect -11489 11124 -11488 12644
rect -9968 11124 -9967 12644
rect -11489 11123 -9967 11124
rect -9459 12644 -7937 12645
rect -9459 11124 -9458 12644
rect -7938 11884 -7937 12644
rect -7938 11784 -7706 11884
rect -7938 11124 -7937 11784
rect -9459 11123 -7937 11124
rect -9226 11029 -9126 11030
rect -9226 10931 -9225 11029
rect -9127 10931 -9126 11029
rect -9226 10732 -9126 10931
rect -13472 10731 -9126 10732
rect -13472 10633 -13471 10731
rect -13373 10633 -10355 10731
rect -10257 10633 -9126 10731
rect -13472 10632 -9126 10633
rect -8102 10881 -8002 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -8002 10881
rect -8102 10545 -8002 10783
rect -11489 10544 -9967 10545
rect -12335 10540 -12013 10541
rect -12635 10010 -12553 10011
rect -12335 10010 -12334 10540
rect -12635 9930 -12634 10010
rect -12554 9930 -12334 10010
rect -12635 9929 -12553 9930
rect -12335 9020 -12334 9930
rect -12014 9020 -12013 10540
rect -11489 9024 -11488 10544
rect -9968 9024 -9967 10544
rect -11489 9023 -9967 9024
rect -9459 10544 -7937 10545
rect -9459 9024 -9458 10544
rect -7938 9024 -7937 10544
rect -9459 9023 -7937 9024
rect -12335 9019 -12013 9020
rect -10182 8864 -10082 9023
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12645 -5834 12804
rect -7299 12644 -5777 12645
rect -7299 11124 -7298 12644
rect -5778 11124 -5777 12644
rect -7299 11123 -5777 11124
rect -5259 12644 -3737 12645
rect -5259 11124 -5258 12644
rect -3738 11884 -3737 12644
rect -3738 11784 -3506 11884
rect -3738 11124 -3737 11784
rect -5259 11123 -3737 11124
rect -5270 11029 -5170 11030
rect -5270 10931 -5269 11029
rect -5171 10931 -5170 11029
rect -7571 10882 -7469 10883
rect -7571 10782 -7570 10882
rect -7470 10782 -7469 10882
rect -7571 10781 -7469 10782
rect -5270 10734 -5170 10931
rect -6556 10733 -5170 10734
rect -6556 10635 -6555 10733
rect -6457 10635 -5170 10733
rect -6556 10634 -5170 10635
rect -3902 10879 -3802 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3802 10879
rect -3902 10545 -3802 10781
rect -7299 10544 -5777 10545
rect -7299 9024 -7298 10544
rect -5778 9024 -5777 10544
rect -7299 9023 -5777 9024
rect -5259 10544 -3737 10545
rect -5259 9024 -5258 10544
rect -3738 9024 -3737 10544
rect -5259 9023 -3737 9024
rect -5952 8864 -5852 9023
rect -3606 8864 -3506 11784
rect -3392 10881 -3292 12804
rect -2397 12803 -2295 12804
rect 37001 12668 37211 12669
rect 37271 12668 37272 13312
rect -3069 12646 -2747 12647
rect -3069 11126 -3068 12646
rect -2748 11856 -2747 12646
rect 37001 12460 37002 12668
rect 37210 12460 37272 12668
rect 37001 12459 37211 12460
rect -2525 11856 -2431 11857
rect -2748 11764 -2524 11856
rect -2432 11764 -2431 11856
rect 37271 11792 37272 12460
rect 37592 11792 37593 13312
rect 37271 11791 37593 11792
rect 38117 13312 39639 13313
rect 38117 11792 38118 13312
rect 39638 11792 39639 13312
rect 38117 11791 39639 11792
rect 40147 13312 41669 13313
rect 40147 11792 40148 13312
rect 41668 12562 41669 13312
rect 41668 12462 41938 12562
rect 41668 11792 41669 12462
rect 40147 11791 41669 11792
rect -2748 11126 -2747 11764
rect -2525 11763 -2431 11764
rect 40292 11709 40392 11710
rect 40292 11611 40293 11709
rect 40391 11611 40392 11709
rect 40292 11412 40392 11611
rect 39488 11411 40392 11412
rect 39488 11313 39489 11411
rect 39587 11313 40392 11411
rect 39488 11312 40392 11313
rect 41542 11559 41642 11560
rect 41542 11461 41543 11559
rect 41641 11461 41642 11559
rect 41542 11213 41642 11461
rect 38117 11212 39639 11213
rect -3069 11125 -2747 11126
rect 37271 11208 37593 11209
rect -3393 10880 -3291 10881
rect -3393 10780 -3392 10880
rect -3292 10780 -3291 10880
rect -3393 10779 -3291 10780
rect -3392 10776 -3292 10779
rect -3069 10542 -2747 10543
rect -3069 9022 -3068 10542
rect -2748 9848 -2747 10542
rect 36930 10528 37118 10529
rect 37271 10528 37272 11208
rect 36930 10342 36931 10528
rect 37117 10342 37272 10528
rect 36930 10341 37118 10342
rect -2519 9848 -2411 9849
rect -2748 9742 -2518 9848
rect -2412 9742 -2411 9848
rect -2748 9022 -2747 9742
rect -2519 9741 -2411 9742
rect 37271 9688 37272 10342
rect 37592 9688 37593 11208
rect 38117 9692 38118 11212
rect 39638 9692 39639 11212
rect 38117 9691 39639 9692
rect 40147 11212 41669 11213
rect 40147 9692 40148 11212
rect 41668 9692 41669 11212
rect 40147 9691 41669 9692
rect 37271 9687 37593 9688
rect 39492 9542 39592 9691
rect 41838 9542 41938 12462
rect 42074 11561 42174 13482
rect 43710 13313 43810 13482
rect 42307 13312 43829 13313
rect 42307 11792 42308 13312
rect 43828 11792 43829 13312
rect 42307 11791 43829 11792
rect 44347 13312 45869 13313
rect 44347 11792 44348 13312
rect 45868 12562 45869 13312
rect 45868 12462 46138 12562
rect 45868 11792 45869 12462
rect 44347 11791 45869 11792
rect 44512 11709 44612 11710
rect 44512 11611 44513 11709
rect 44611 11611 44612 11709
rect 42073 11560 42175 11561
rect 42073 11460 42074 11560
rect 42174 11460 42175 11560
rect 42073 11459 42175 11460
rect 44512 11394 44612 11611
rect 43688 11393 44612 11394
rect 43688 11295 43689 11393
rect 43787 11295 44612 11393
rect 43688 11294 44612 11295
rect 45742 11559 45842 11560
rect 45742 11461 45743 11559
rect 45841 11461 45842 11559
rect 45742 11213 45842 11461
rect 42307 11212 43829 11213
rect 42307 9692 42308 11212
rect 43828 9692 43829 11212
rect 42307 9691 43829 9692
rect 44347 11212 45869 11213
rect 44347 9692 44348 11212
rect 45868 9692 45869 11212
rect 44347 9691 45869 9692
rect 43692 9542 43792 9691
rect 46038 9542 46138 12462
rect 46218 11561 46318 13482
rect 46537 13314 46859 13315
rect 46537 11794 46538 13314
rect 46858 12610 46859 13314
rect 47029 12610 47193 12611
rect 46858 12448 47030 12610
rect 47192 12448 47193 12610
rect 46858 11794 46859 12448
rect 47029 12447 47193 12448
rect 46537 11793 46859 11794
rect 46217 11560 46319 11561
rect 46217 11460 46218 11560
rect 46318 11556 46319 11560
rect 46318 11460 53150 11556
rect 46217 11459 53150 11460
rect 46218 11456 53150 11459
rect 46537 11210 46859 11211
rect 46537 9690 46538 11210
rect 46858 10510 46859 11210
rect 46991 10510 47161 10511
rect 46858 10342 46992 10510
rect 47160 10342 47161 10510
rect 46858 9690 46859 10342
rect 46991 10341 47161 10342
rect 46537 9689 46859 9690
rect 36254 9541 52282 9542
rect 36254 9443 36255 9541
rect 36353 9443 52282 9541
rect 36254 9442 52282 9443
rect -3069 9021 -2747 9022
rect -10182 8863 -1656 8864
rect -10182 8765 -1755 8863
rect -1657 8765 -1656 8863
rect 42573 8792 44095 8793
rect -10182 8764 -1656 8765
rect 37402 8790 39724 8791
rect -10535 8620 -10433 8621
rect -13100 8619 -10534 8620
rect -13100 8521 -13099 8619
rect -13001 8521 -10534 8619
rect -13100 8520 -10534 8521
rect -10434 8520 -10433 8620
rect -10535 8519 -10433 8520
rect 37402 8470 37403 8790
rect 39723 8470 39724 8790
rect 37402 8469 39724 8470
rect 40185 8790 41707 8791
rect 40185 8470 40186 8790
rect 41706 8470 41707 8790
rect 42573 8472 42574 8792
rect 44094 8472 44095 8792
rect 42573 8471 44095 8472
rect 44556 8792 46878 8793
rect 44556 8472 44557 8792
rect 46877 8472 46878 8792
rect 44556 8471 46878 8472
rect 40185 8469 41707 8470
rect 38394 8400 38748 8469
rect 38394 8172 38476 8400
rect 38704 8172 38748 8400
rect -7033 8124 -5511 8125
rect -12204 8122 -9882 8123
rect -12204 7802 -12203 8122
rect -9883 7802 -9882 8122
rect -12204 7801 -9882 7802
rect -9421 8122 -7899 8123
rect -9421 7802 -9420 8122
rect -7900 7802 -7899 8122
rect -7033 7804 -7032 8124
rect -5512 7804 -5511 8124
rect -7033 7803 -5511 7804
rect -5050 8124 -2728 8125
rect -5050 7804 -5049 8124
rect -2729 7804 -2728 8124
rect -5050 7803 -2728 7804
rect -9421 7801 -7899 7802
rect -11198 7646 -10956 7801
rect -11198 7406 -11197 7646
rect -10957 7406 -10956 7646
rect -11198 7057 -10956 7406
rect -8786 7646 -8544 7801
rect -8786 7406 -8785 7646
rect -8545 7406 -8544 7646
rect -8786 7057 -8544 7406
rect -6374 7646 -6132 7803
rect -6374 7406 -6373 7646
rect -6133 7406 -6132 7646
rect -6374 7057 -6132 7406
rect -3962 7646 -3720 7803
rect 36995 7738 37097 7739
rect -3962 7406 -3961 7646
rect -3721 7406 -3720 7646
rect 35228 7737 36996 7738
rect 35228 7639 35229 7737
rect 35327 7639 36996 7737
rect 35228 7638 36996 7639
rect 37096 7638 37097 7738
rect 36995 7637 37097 7638
rect -3962 7057 -3720 7406
rect 38394 7174 38748 8172
rect -11199 7056 -10955 7057
rect -11199 6814 -11198 7056
rect -10956 6814 -10955 7056
rect -11199 6813 -10955 6814
rect -8787 7056 -8543 7057
rect -8787 6814 -8786 7056
rect -8544 6814 -8543 7056
rect -8787 6813 -8543 6814
rect -6375 7056 -6131 7057
rect -6375 6814 -6374 7056
rect -6132 6814 -6131 7056
rect -6375 6813 -6131 6814
rect -3963 7056 -3719 7057
rect -3963 6814 -3962 7056
rect -3720 6814 -3719 7056
rect 38394 6992 38428 7174
rect 38610 6992 38748 7174
rect 38394 6925 38748 6992
rect 40796 8398 41150 8469
rect 40796 8170 40888 8398
rect 41116 8170 41150 8398
rect 40796 7174 41150 8170
rect 40796 6992 40828 7174
rect 41010 6992 41150 7174
rect 40796 6925 41150 6992
rect 43168 8398 43504 8471
rect 43168 8170 43232 8398
rect 43460 8170 43504 8398
rect 43168 7174 43504 8170
rect 43168 6992 43240 7174
rect 43422 6992 43504 7174
rect 43168 6927 43504 6992
rect 45576 8398 45872 8471
rect 45576 8170 45620 8398
rect 45848 8170 45872 8398
rect 45576 7174 45872 8170
rect 45576 6992 45640 7174
rect 45822 6992 45872 7174
rect 45576 6927 45872 6992
rect 42591 6926 44113 6927
rect -3963 6813 -3719 6814
rect 37420 6924 39742 6925
rect -11198 6659 -10956 6813
rect -8786 6659 -8544 6813
rect -6374 6661 -6132 6813
rect -3962 6661 -3720 6813
rect -7033 6660 -5511 6661
rect -12204 6658 -9882 6659
rect -12204 6338 -12203 6658
rect -9883 6338 -9882 6658
rect -12204 6337 -9882 6338
rect -9421 6658 -7899 6659
rect -9421 6338 -9420 6658
rect -7900 6338 -7899 6658
rect -7033 6340 -7032 6660
rect -5512 6340 -5511 6660
rect -7033 6339 -5511 6340
rect -5050 6660 -2728 6661
rect -5050 6340 -5049 6660
rect -2729 6340 -2728 6660
rect 37420 6604 37421 6924
rect 39741 6604 39742 6924
rect 37420 6603 39742 6604
rect 40203 6924 41725 6925
rect 40203 6604 40204 6924
rect 41724 6604 41725 6924
rect 42591 6606 42592 6926
rect 44112 6606 44113 6926
rect 42591 6605 44113 6606
rect 44574 6926 46896 6927
rect 44574 6606 44575 6926
rect 46895 6606 46896 6926
rect 44574 6605 46896 6606
rect 40203 6603 41725 6604
rect -5050 6339 -2728 6340
rect -9421 6337 -7899 6338
rect 39053 6198 39155 6199
rect 36458 6197 39054 6198
rect 36458 6099 36459 6197
rect 36557 6099 39054 6197
rect 36458 6098 39054 6099
rect 39154 6098 39155 6198
rect 39053 6097 39155 6098
rect 39510 5981 48576 5982
rect 39510 5883 48477 5981
rect 48575 5883 48576 5981
rect 39510 5882 48576 5883
rect 39510 5711 39610 5882
rect 37289 5710 37611 5711
rect -12732 5665 -2322 5666
rect -12732 5567 -12731 5665
rect -12633 5567 -2421 5665
rect -2323 5567 -2322 5665
rect -12732 5566 -2322 5567
rect -10118 5445 -10018 5566
rect -12335 5444 -12013 5445
rect -12587 4766 -12435 4767
rect -12335 4766 -12334 5444
rect -12587 4616 -12586 4766
rect -12436 4616 -12334 4766
rect -12587 4615 -12435 4616
rect -12335 3924 -12334 4616
rect -12014 3924 -12013 5444
rect -12335 3923 -12013 3924
rect -11489 5444 -9967 5445
rect -11489 3924 -11488 5444
rect -9968 3924 -9967 5444
rect -11489 3923 -9967 3924
rect -9459 5444 -7937 5445
rect -9459 3924 -9458 5444
rect -7938 4646 -7937 5444
rect -7938 4546 -7690 4646
rect -7938 3924 -7937 4546
rect -9459 3923 -7937 3924
rect -9366 3827 -9266 3828
rect -9366 3729 -9365 3827
rect -9267 3729 -9266 3827
rect -9366 3538 -9266 3729
rect -13304 3537 -9266 3538
rect -13304 3439 -13303 3537
rect -13205 3439 -10167 3537
rect -10069 3439 -9266 3537
rect -13304 3438 -9266 3439
rect -8086 3681 -7986 3682
rect -8086 3583 -8085 3681
rect -7987 3583 -7986 3681
rect -8086 3345 -7986 3583
rect -11489 3344 -9967 3345
rect -12335 3340 -12013 3341
rect -12581 2650 -12453 2651
rect -12335 2650 -12334 3340
rect -12581 2524 -12580 2650
rect -12454 2524 -12334 2650
rect -12581 2523 -12453 2524
rect -12335 1820 -12334 2524
rect -12014 1820 -12013 3340
rect -11489 1824 -11488 3344
rect -9968 1824 -9967 3344
rect -11489 1823 -9967 1824
rect -9459 3344 -7937 3345
rect -9459 1824 -9458 3344
rect -7938 1824 -7937 3344
rect -9459 1823 -7937 1824
rect -12335 1819 -12013 1820
rect -10136 1628 -10036 1823
rect -13098 1627 -9512 1628
rect -13098 1529 -13097 1627
rect -12999 1626 -9512 1627
rect -7790 1626 -7690 4546
rect -7554 3683 -7454 5566
rect -5918 5445 -5818 5566
rect -7299 5444 -5777 5445
rect -7299 3924 -7298 5444
rect -5778 3924 -5777 5444
rect -7299 3923 -5777 3924
rect -5259 5444 -3737 5445
rect -5259 3924 -5258 5444
rect -3738 4646 -3737 5444
rect -3738 4546 -3490 4646
rect -3738 3924 -3737 4546
rect -5259 3923 -3737 3924
rect -5144 3839 -5028 3840
rect -5144 3725 -5143 3839
rect -5029 3725 -5028 3839
rect -7555 3682 -7453 3683
rect -7555 3582 -7554 3682
rect -7454 3582 -7453 3682
rect -7555 3581 -7453 3582
rect -5909 3542 -5791 3543
rect -5144 3542 -5028 3725
rect -5909 3426 -5908 3542
rect -5792 3426 -5028 3542
rect -3886 3683 -3786 3684
rect -3886 3585 -3885 3683
rect -3787 3585 -3786 3683
rect -5909 3425 -5791 3426
rect -3886 3345 -3786 3585
rect -7299 3344 -5777 3345
rect -7299 1824 -7298 3344
rect -5778 1824 -5777 3344
rect -7299 1823 -5777 1824
rect -5259 3344 -3737 3345
rect -5259 1824 -5258 3344
rect -3738 1824 -3737 3344
rect -5259 1823 -3737 1824
rect -5936 1626 -5836 1823
rect -3590 1626 -3490 4546
rect -3382 3685 -3282 5566
rect -3069 5446 -2747 5447
rect -3069 3926 -3068 5446
rect -2748 4716 -2747 5446
rect 37019 5066 37229 5067
rect 37289 5066 37290 5710
rect 37019 4858 37020 5066
rect 37228 4858 37290 5066
rect 37019 4857 37229 4858
rect -2661 4716 -2505 4717
rect -2748 4562 -2660 4716
rect -2506 4562 -2505 4716
rect -2748 3926 -2747 4562
rect -2661 4561 -2505 4562
rect 37289 4190 37290 4858
rect 37610 4190 37611 5710
rect 37289 4189 37611 4190
rect 38135 5710 39657 5711
rect 38135 4190 38136 5710
rect 39656 4190 39657 5710
rect 38135 4189 39657 4190
rect 40165 5710 41687 5711
rect 40165 4190 40166 5710
rect 41686 4962 41687 5710
rect 41686 4862 41938 4962
rect 41686 4190 41687 4862
rect 40165 4189 41687 4190
rect -3069 3925 -2747 3926
rect 40278 4105 40378 4106
rect 40278 4007 40279 4105
rect 40377 4007 40378 4105
rect 40278 3798 40378 4007
rect 39488 3797 40378 3798
rect 39488 3699 39489 3797
rect 39587 3699 40378 3797
rect 39488 3698 40378 3699
rect 41542 3959 41642 3960
rect 41542 3861 41543 3959
rect 41641 3861 41642 3959
rect -3383 3684 -3281 3685
rect -3383 3584 -3382 3684
rect -3282 3584 -3281 3684
rect 41542 3611 41642 3861
rect 38135 3610 39657 3611
rect -3383 3583 -3281 3584
rect 37289 3606 37611 3607
rect -3069 3342 -2747 3343
rect -3069 1822 -3068 3342
rect -2748 2664 -2747 3342
rect 36948 2926 37136 2927
rect 37289 2926 37290 3606
rect 36948 2740 36949 2926
rect 37135 2740 37290 2926
rect 36948 2739 37136 2740
rect -2667 2664 -2505 2665
rect -2748 2504 -2666 2664
rect -2506 2504 -2505 2664
rect -2748 1822 -2747 2504
rect -2667 2503 -2505 2504
rect 37289 2086 37290 2740
rect 37610 2086 37611 3606
rect 38135 2090 38136 3610
rect 39656 2090 39657 3610
rect 38135 2089 39657 2090
rect 40165 3610 41687 3611
rect 40165 2090 40166 3610
rect 41686 2090 41687 3610
rect 40165 2089 41687 2090
rect 37289 2085 37611 2086
rect 39492 1942 39592 2089
rect 41838 1942 41938 4862
rect 42074 3961 42174 5882
rect 43710 5711 43810 5882
rect 42325 5710 43847 5711
rect 42325 4190 42326 5710
rect 43846 4190 43847 5710
rect 42325 4189 43847 4190
rect 44365 5710 45887 5711
rect 44365 4190 44366 5710
rect 45886 4962 45887 5710
rect 45886 4862 46138 4962
rect 45886 4190 45887 4862
rect 44365 4189 45887 4190
rect 44490 4089 44590 4090
rect 44490 3991 44491 4089
rect 44589 3991 44590 4089
rect 42073 3960 42175 3961
rect 42073 3860 42074 3960
rect 42174 3860 42175 3960
rect 42073 3859 42175 3860
rect 44490 3800 44590 3991
rect 43688 3799 44590 3800
rect 43688 3701 43689 3799
rect 43787 3701 44590 3799
rect 43688 3700 44590 3701
rect 45742 3959 45842 3960
rect 45742 3861 45743 3959
rect 45841 3861 45842 3959
rect 45742 3611 45842 3861
rect 42325 3610 43847 3611
rect 42325 2090 42326 3610
rect 43846 2090 43847 3610
rect 42325 2089 43847 2090
rect 44365 3610 45887 3611
rect 44365 2090 44366 3610
rect 45886 2090 45887 3610
rect 44365 2089 45887 2090
rect 43692 1942 43792 2089
rect 46038 1942 46138 4862
rect 46238 3961 46338 5882
rect 46555 5712 46877 5713
rect 46555 4192 46556 5712
rect 46876 5008 46877 5712
rect 47047 5008 47211 5009
rect 46876 4846 47048 5008
rect 47210 4846 47211 5008
rect 46876 4192 46877 4846
rect 47047 4845 47211 4846
rect 52182 4955 52282 9442
rect 53050 7723 53150 11456
rect 53049 7722 53151 7723
rect 53049 7622 53050 7722
rect 53150 7622 53151 7722
rect 53049 7621 53151 7622
rect 53050 5605 53150 7621
rect 53047 5604 53150 5605
rect 53047 5504 53048 5604
rect 53148 5504 53150 5604
rect 53047 5503 53150 5504
rect 52182 4857 52183 4955
rect 52281 4857 52282 4955
rect 46555 4191 46877 4192
rect 52182 4087 52282 4857
rect 46237 3960 46339 3961
rect 46237 3860 46238 3960
rect 46338 3860 46339 3960
rect 46237 3859 46339 3860
rect 48481 3756 48583 3757
rect 48481 3656 48482 3756
rect 48582 3656 48583 3756
rect 48481 3655 48583 3656
rect 46555 3608 46877 3609
rect 46555 2088 46556 3608
rect 46876 2908 46877 3608
rect 47009 2908 47179 2909
rect 46876 2740 47010 2908
rect 47178 2740 47179 2908
rect 46876 2088 46877 2740
rect 47009 2739 47179 2740
rect 46555 2087 46877 2088
rect 48482 1942 48582 3655
rect 52181 3606 52283 4087
rect 52180 3605 52284 3606
rect 52180 3503 52181 3605
rect 52283 3503 52284 3605
rect 52180 3502 52284 3503
rect 39492 1842 48582 1942
rect 52181 1897 52283 3502
rect 53050 2833 53150 5503
rect 53050 2735 53051 2833
rect 53149 2735 53150 2833
rect 53050 2734 53150 2735
rect -3069 1821 -2747 1822
rect 39165 1692 39267 1693
rect 36054 1691 39166 1692
rect -12999 1625 -2234 1626
rect -12999 1529 -2333 1625
rect -13098 1528 -2333 1529
rect -10136 1527 -2333 1528
rect -2235 1527 -2234 1625
rect 36054 1593 36055 1691
rect 36153 1593 39166 1691
rect 36054 1592 39166 1593
rect 39266 1592 39267 1692
rect 52177 1673 52287 1897
rect 39165 1591 39267 1592
rect 52176 1672 52288 1673
rect 52176 1562 52177 1672
rect 52287 1562 52288 1672
rect 52176 1561 52288 1562
rect -10136 1526 -2234 1527
rect 42591 1190 44113 1191
rect 37420 1188 39742 1189
rect -7033 924 -5511 925
rect -12204 922 -9882 923
rect -12204 602 -12203 922
rect -9883 602 -9882 922
rect -12204 601 -9882 602
rect -9421 922 -7899 923
rect -9421 602 -9420 922
rect -7900 602 -7899 922
rect -7033 604 -7032 924
rect -5512 604 -5511 924
rect -7033 603 -5511 604
rect -5050 924 -2728 925
rect -5050 604 -5049 924
rect -2729 604 -2728 924
rect 37420 868 37421 1188
rect 39741 868 39742 1188
rect 37420 867 39742 868
rect 40203 1188 41725 1189
rect 40203 868 40204 1188
rect 41724 868 41725 1188
rect 42591 870 42592 1190
rect 44112 870 44113 1190
rect 42591 869 44113 870
rect 44574 1190 46896 1191
rect 44574 870 44575 1190
rect 46895 870 46896 1190
rect 44574 869 46896 870
rect 40203 867 41725 868
rect 38494 799 38722 867
rect -5050 603 -2728 604
rect 38493 798 38723 799
rect -9421 601 -7899 602
rect -11156 513 -10918 601
rect -8744 513 -8506 601
rect -6332 513 -6094 603
rect -3920 513 -3682 603
rect 38493 570 38494 798
rect 38722 570 38723 798
rect 40906 797 41134 867
rect 43250 797 43478 869
rect 45638 797 45866 869
rect 38493 569 38723 570
rect 40905 796 41135 797
rect -11157 512 -10917 513
rect -11157 274 -11156 512
rect -10918 274 -10917 512
rect -11157 273 -10917 274
rect -8745 512 -8505 513
rect -8745 274 -8744 512
rect -8506 274 -8505 512
rect -8745 273 -8505 274
rect -6333 512 -6093 513
rect -6333 274 -6332 512
rect -6094 274 -6093 512
rect -6333 273 -6093 274
rect -3921 512 -3681 513
rect -3921 274 -3920 512
rect -3682 274 -3681 512
rect -3921 273 -3681 274
rect -11156 140 -10918 273
rect -8744 140 -8506 273
rect -6332 140 -6094 273
rect -3920 140 -3682 273
rect 38494 140 38722 569
rect 40905 568 40906 796
rect 41134 568 41135 796
rect 40905 567 41135 568
rect 43249 796 43479 797
rect 43249 568 43250 796
rect 43478 568 43479 796
rect 43249 567 43479 568
rect 45637 796 45867 797
rect 45637 568 45638 796
rect 45866 568 45867 796
rect 45637 567 45867 568
rect 40906 140 41134 567
rect 43250 140 43478 567
rect 45638 140 45866 567
rect -13292 64 90192 140
rect -13292 -90 3478 64
rect 34878 -90 57478 64
rect 88878 -90 90192 64
rect -13292 -276 90192 -90
rect -13292 -576 -1266 -276
rect -666 -576 35166 -276
rect 35766 -576 52734 -276
rect 53334 -576 89166 -276
rect 89766 -576 90192 -276
rect -13292 -660 90192 -576
<< labels >>
flabel metal4 -9700 5602 -9690 5614 1 FreeSans 480 0 0 0 vip1
flabel metal4 -9752 1570 -9732 1586 1 FreeSans 480 0 0 0 vim1
flabel metal4 -5616 -342 -5562 -296 1 FreeSans 480 0 0 0 VSS
port 2 n ground bidirectional
flabel metal4 39914 1890 39924 1898 1 FreeSans 480 0 0 0 venp1
flabel metal4 39912 5932 39922 5950 1 FreeSans 480 0 0 0 venm1
flabel metal4 39872 9472 39892 9486 1 FreeSans 480 0 0 0 vim2
flabel metal4 39942 13524 39962 13540 1 FreeSans 480 0 0 0 vip2
flabel metal4 40082 15590 40102 15606 1 FreeSans 480 0 0 0 venp2
flabel metal4 40024 19636 40048 19656 1 FreeSans 480 0 0 0 venm2
flabel metal4 40068 25698 40084 25712 1 FreeSans 480 0 0 0 vop
port 10 n
flabel metal4 49508 27900 49618 28008 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel metal2 50956 4528 50982 4554 1 FreeSans 480 0 0 0 gain_ctrl_0
port 5 n
flabel metal2 49538 23440 49558 23458 1 FreeSans 480 0 0 0 gain_ctrl_1
port 6 n
flabel metal4 36296 7672 36328 7702 1 FreeSans 480 0 0 0 vocm
port 7 n
flabel metal1 3968 4954 3982 4962 1 FreeSans 480 0 0 0 ibiasn1
port 8 n
flabel metal1 57962 4966 57978 4972 1 FreeSans 480 0 0 0 ibiasn2
port 11 n
flabel metal1 -7768 15456 -7762 15460 1 FreeSans 480 0 0 0 rst_n
port 12 n
flabel metal1 -8136 15450 -8128 15458 1 FreeSans 480 0 0 0 rst
flabel metal3 -9694 13074 -9674 13090 1 FreeSans 480 0 0 0 vip1
flabel metal4 -9728 8802 -9684 8828 1 FreeSans 480 0 0 0 vop1
flabel metal4 -9734 12846 -9714 12872 1 FreeSans 480 0 0 0 vom1
flabel metal3 -9770 8556 -9744 8576 1 FreeSans 480 0 0 0 vim1
flabel metal3 -9338 5886 -9298 5918 1 FreeSans 480 0 0 0 vhpf
port 4 n
flabel metal3 -9718 1372 -9700 1386 1 FreeSans 480 0 0 0 vincm
port 3 n
flabel metal3 39912 1630 39926 1644 1 FreeSans 480 0 0 0 vop1
flabel metal3 39900 6144 39910 6156 1 FreeSans 480 0 0 0 vom1
flabel metal3 39848 9234 39866 9256 1 FreeSans 480 0 0 0 vop1
flabel metal3 39924 13774 39940 13786 1 FreeSans 480 0 0 0 vom1
flabel metal3 40106 19872 40122 19884 1 FreeSans 480 0 0 0 vip2
flabel metal3 40076 15316 40096 15328 1 FreeSans 480 0 0 0 vim2
flabel metal2 40896 23642 40916 23660 1 FreeSans 480 0 0 0 vim2
flabel metal4 39646 23514 39664 23536 1 FreeSans 480 0 0 0 vip2
flabel metal4 41878 23258 41900 23278 1 FreeSans 480 0 0 0 vom
port 9 n
flabel locali -8032 15507 -7998 15541 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -8032 15439 -7998 15473 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7940 15439 -7906 15473 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell -7897 15745 -7863 15779 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -7897 15201 -7863 15235 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -7897 15201 -7863 15235 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -7897 15745 -7863 15779 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -7834 15218 -7834 15218 6 sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -10899 15446 -10891 15452 1 FreeSans 480 0 0 0 txgate_4/tx
flabel metal1 -12717 15426 -12707 15434 1 FreeSans 480 0 0 0 txgate_4/out
flabel metal1 -12455 15432 -12445 15440 1 FreeSans 480 0 0 0 txgate_4/in
flabel metal1 -12201 16374 -12191 16384 1 FreeSans 480 0 0 0 txgate_4/VDD
flabel metal1 -12203 14684 -12195 14690 1 FreeSans 480 0 0 0 txgate_4/VSS
flabel metal2 -11201 15948 -11191 15956 1 FreeSans 480 0 0 0 txgate_4/txb
flabel locali -11132 15507 -11098 15541 0 FreeSans 340 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -11132 15439 -11098 15473 0 FreeSans 340 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -11040 15439 -11006 15473 0 FreeSans 340 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -10997 15745 -10963 15779 0 FreeSans 200 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -10997 15201 -10963 15235 0 FreeSans 200 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -10997 15201 -10963 15235 0 FreeSans 200 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -10997 15745 -10963 15779 0 FreeSans 200 0 0 0 txgate_4/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -10934 15218 -10934 15218 6 txgate_4/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -8299 15446 -8291 15452 1 FreeSans 480 0 0 0 txgate_5/tx
flabel metal1 -10117 15426 -10107 15434 1 FreeSans 480 0 0 0 txgate_5/out
flabel metal1 -9855 15432 -9845 15440 1 FreeSans 480 0 0 0 txgate_5/in
flabel metal1 -9601 16374 -9591 16384 1 FreeSans 480 0 0 0 txgate_5/VDD
flabel metal1 -9603 14684 -9595 14690 1 FreeSans 480 0 0 0 txgate_5/VSS
flabel metal2 -8601 15948 -8591 15956 1 FreeSans 480 0 0 0 txgate_5/txb
flabel locali -8532 15507 -8498 15541 0 FreeSans 340 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -8532 15439 -8498 15473 0 FreeSans 340 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -8440 15439 -8406 15473 0 FreeSans 340 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -8397 15745 -8363 15779 0 FreeSans 200 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -8397 15201 -8363 15235 0 FreeSans 200 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -8397 15201 -8363 15235 0 FreeSans 200 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -8397 15745 -8363 15779 0 FreeSans 200 0 0 0 txgate_5/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -8334 15218 -8334 15218 6 txgate_5/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal2 20874 23830 20874 23830 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vfoldm
flabel metal1 17306 26040 17306 26040 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M1d
flabel metal1 18470 23856 18470 23856 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M2d
flabel metal2 18748 26016 18748 26016 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M6d
flabel metal1 18290 22924 18290 22924 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M1d
flabel metal2 18568 21958 18568 21958 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias1
flabel metal2 18464 18386 18464 18386 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M2d
flabel metal2 27422 20892 27422 20892 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M6d
flabel metal1 27618 20540 27618 20540 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M13d
flabel metal2 22822 18108 22822 18108 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M3d
flabel metal1 31676 20922 31676 20922 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vfoldm
flabel metal2 31548 19646 31548 19646 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vfoldp
flabel metal2 22780 27256 22780 27256 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vfoldp
flabel metal2 14914 20354 14914 20354 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmc_casc
flabel metal2 16750 19406 16750 19406 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmcn_casc
flabel metal1 17030 18870 17030 18870 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmcn2_casc
flabel metal1 14474 19284 14474 19284 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmcn1_casc
flabel metal2 19274 27390 19274 27390 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias1
flabel metal2 33336 20798 33368 20814 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vom
flabel metal1 33524 19640 33566 19662 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vop
flabel metal2 20252 27128 20282 27156 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/VDD
flabel metal2 8452 7148 8526 7182 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vocm
flabel metal1 4602 4954 4634 4974 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/ibiasn
flabel metal1 13198 9466 13220 9494 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vom
flabel metal2 23354 11380 23386 11398 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vop
flabel metal1 34130 8502 34154 8532 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/VSS
flabel metal1 5620 1544 5656 1580 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/VSS
flabel metal1 34506 9350 34506 9350 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias3
flabel metal1 13094 13808 13094 13808 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmc_casc
flabel metal1 8010 5912 8010 5912 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmn_casc_tail2
flabel metal2 7882 6324 7882 6324 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmn_casc_tail1
flabel metal1 11082 6918 11082 6918 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmcn2_casc
flabel metal1 10612 6396 10612 6396 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmcn_casc
flabel metal1 10968 7052 10968 7052 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmcn1_casc
flabel metal2 9836 5024 9836 5024 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vfoldp
flabel metal1 8294 3038 8328 3070 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vip
flabel metal1 12046 3246 12072 3276 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vim
flabel metal1 15598 10104 15598 10104 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcascnp
flabel metal1 34250 9556 34250 9556 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcascnm
flabel metal1 34386 5324 34386 5324 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias4
flabel metal1 12956 12056 12956 12056 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vtail_casc
flabel metal1 34628 13722 34628 13726 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M3d
flabel metal1 33904 11204 33904 11204 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/M13d
flabel metal1 11542 3792 11542 3792 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vtail_casc
flabel metal1 8858 2724 8858 2724 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vfoldm
flabel metal1 1444 3634 1444 3634 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmn_casc_tail2
flabel metal1 2586 2904 2586 2904 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias2
flabel metal1 6658 2676 6658 2676 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vcmn_casc_tail1
flabel metal1 2872 14188 2872 14188 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias1
flabel metal1 4744 7514 4744 7514 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vbias2
flabel metal4 9608 21342 9684 21384 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vom
flabel metal4 130 23836 194 23876 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vop
flabel metal1 8500 6614 8528 6650 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vom
flabel metal2 10182 6550 10214 6572 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/vop
flabel metal1 28460 22146 28496 22174 1 FreeSans 480 0 0 0 diff_fold_casc_ota_0/VDD
flabel metal4 -1450 27540 -1450 28340 3 FreeSans 3200 0 0 0 diff_fold_casc_ota_0/VDD
flabel metal4 -1450 -660 -1450 140 3 FreeSans 3200 0 0 0 diff_fold_casc_ota_0/VSS
flabel metal1 50885 1558 50893 1564 1 FreeSans 480 0 0 0 txgate_6/tx
flabel metal1 49067 1538 49077 1546 1 FreeSans 480 0 0 0 txgate_6/out
flabel metal1 49329 1544 49339 1552 1 FreeSans 480 0 0 0 txgate_6/in
flabel metal1 49583 2486 49593 2496 1 FreeSans 480 0 0 0 txgate_6/VDD
flabel metal1 49581 796 49589 802 1 FreeSans 480 0 0 0 txgate_6/VSS
flabel metal2 50583 2060 50593 2068 1 FreeSans 480 0 0 0 txgate_6/txb
flabel locali 50652 1619 50686 1653 0 FreeSans 340 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50652 1551 50686 1585 0 FreeSans 340 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50744 1551 50778 1585 0 FreeSans 340 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 50787 1857 50821 1891 0 FreeSans 200 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 50787 1313 50821 1347 0 FreeSans 200 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 50787 1313 50821 1347 0 FreeSans 200 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 50787 1857 50821 1891 0 FreeSans 200 0 0 0 txgate_6/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 50850 1330 50850 1330 6 txgate_6/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 50885 3648 50893 3654 1 FreeSans 480 0 0 0 txgate_1/tx
flabel metal1 49067 3628 49077 3636 1 FreeSans 480 0 0 0 txgate_1/out
flabel metal1 49329 3634 49339 3642 1 FreeSans 480 0 0 0 txgate_1/in
flabel metal1 49583 4576 49593 4586 1 FreeSans 480 0 0 0 txgate_1/VDD
flabel metal1 49581 2886 49589 2892 1 FreeSans 480 0 0 0 txgate_1/VSS
flabel metal2 50583 4150 50593 4158 1 FreeSans 480 0 0 0 txgate_1/txb
flabel locali 50652 3709 50686 3743 0 FreeSans 340 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50652 3641 50686 3675 0 FreeSans 340 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50744 3641 50778 3675 0 FreeSans 340 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 50787 3947 50821 3981 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 50787 3403 50821 3437 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 50787 3403 50821 3437 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 50787 3947 50821 3981 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 50850 3420 50850 3420 6 txgate_1/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 50885 5648 50893 5654 1 FreeSans 480 0 0 0 txgate_0/tx
flabel metal1 49067 5628 49077 5636 1 FreeSans 480 0 0 0 txgate_0/out
flabel metal1 49329 5634 49339 5642 1 FreeSans 480 0 0 0 txgate_0/in
flabel metal1 49583 6576 49593 6586 1 FreeSans 480 0 0 0 txgate_0/VDD
flabel metal1 49581 4886 49589 4892 1 FreeSans 480 0 0 0 txgate_0/VSS
flabel metal2 50583 6150 50593 6158 1 FreeSans 480 0 0 0 txgate_0/txb
flabel locali 50652 5709 50686 5743 0 FreeSans 340 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50652 5641 50686 5675 0 FreeSans 340 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50744 5641 50778 5675 0 FreeSans 340 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 50787 5947 50821 5981 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 50787 5403 50821 5437 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 50787 5403 50821 5437 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 50787 5947 50821 5981 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 50850 5420 50850 5420 6 txgate_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 50885 7612 50893 7618 1 FreeSans 480 0 0 0 txgate_7/tx
flabel metal1 49067 7592 49077 7600 1 FreeSans 480 0 0 0 txgate_7/out
flabel metal1 49329 7598 49339 7606 1 FreeSans 480 0 0 0 txgate_7/in
flabel metal1 49583 8540 49593 8550 1 FreeSans 480 0 0 0 txgate_7/VDD
flabel metal1 49581 6850 49589 6856 1 FreeSans 480 0 0 0 txgate_7/VSS
flabel metal2 50583 8114 50593 8122 1 FreeSans 480 0 0 0 txgate_7/txb
flabel locali 50652 7673 50686 7707 0 FreeSans 340 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50652 7605 50686 7639 0 FreeSans 340 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 50744 7605 50778 7639 0 FreeSans 340 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 50787 7911 50821 7945 0 FreeSans 200 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 50787 7367 50821 7401 0 FreeSans 200 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 50787 7367 50821 7401 0 FreeSans 200 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 50787 7911 50821 7945 0 FreeSans 200 0 0 0 txgate_7/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 50850 7384 50850 7384 6 txgate_7/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 49459 22576 49467 22582 1 FreeSans 480 0 0 0 txgate_2/tx
flabel metal1 47641 22556 47651 22564 1 FreeSans 480 0 0 0 txgate_2/out
flabel metal1 47903 22562 47913 22570 1 FreeSans 480 0 0 0 txgate_2/in
flabel metal1 48157 23504 48167 23514 1 FreeSans 480 0 0 0 txgate_2/VDD
flabel metal1 48155 21814 48163 21820 1 FreeSans 480 0 0 0 txgate_2/VSS
flabel metal2 49157 23078 49167 23086 1 FreeSans 480 0 0 0 txgate_2/txb
flabel locali 49226 22637 49260 22671 0 FreeSans 340 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 49226 22569 49260 22603 0 FreeSans 340 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 49318 22569 49352 22603 0 FreeSans 340 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 49361 22875 49395 22909 0 FreeSans 200 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 49361 22331 49395 22365 0 FreeSans 200 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 49361 22331 49395 22365 0 FreeSans 200 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 49361 22875 49395 22909 0 FreeSans 200 0 0 0 txgate_2/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 49424 22348 49424 22348 6 txgate_2/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 49459 24576 49467 24582 1 FreeSans 480 0 0 0 txgate_3/tx
flabel metal1 47641 24556 47651 24564 1 FreeSans 480 0 0 0 txgate_3/out
flabel metal1 47903 24562 47913 24570 1 FreeSans 480 0 0 0 txgate_3/in
flabel metal1 48157 25504 48167 25514 1 FreeSans 480 0 0 0 txgate_3/VDD
flabel metal1 48155 23814 48163 23820 1 FreeSans 480 0 0 0 txgate_3/VSS
flabel metal2 49157 25078 49167 25086 1 FreeSans 480 0 0 0 txgate_3/txb
flabel locali 49226 24637 49260 24671 0 FreeSans 340 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 49226 24569 49260 24603 0 FreeSans 340 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 49318 24569 49352 24603 0 FreeSans 340 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 49361 24875 49395 24909 0 FreeSans 200 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 49361 24331 49395 24365 0 FreeSans 200 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 49361 24331 49395 24365 0 FreeSans 200 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 49361 24875 49395 24909 0 FreeSans 200 0 0 0 txgate_3/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 49424 24348 49424 24348 6 txgate_3/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal2 74874 23830 74874 23830 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vfoldm
flabel metal1 71306 26040 71306 26040 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M1d
flabel metal1 72470 23856 72470 23856 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M2d
flabel metal2 72748 26016 72748 26016 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M6d
flabel metal1 72290 22924 72290 22924 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M1d
flabel metal2 72568 21958 72568 21958 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias1
flabel metal2 72464 18386 72464 18386 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M2d
flabel metal2 81422 20892 81422 20892 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M6d
flabel metal1 81618 20540 81618 20540 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M13d
flabel metal2 76822 18108 76822 18108 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M3d
flabel metal1 85676 20922 85676 20922 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vfoldm
flabel metal2 85548 19646 85548 19646 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vfoldp
flabel metal2 76780 27256 76780 27256 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vfoldp
flabel metal2 68914 20354 68914 20354 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmc_casc
flabel metal2 70750 19406 70750 19406 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmcn_casc
flabel metal1 71030 18870 71030 18870 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmcn2_casc
flabel metal1 68474 19284 68474 19284 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmcn1_casc
flabel metal2 73274 27390 73274 27390 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias1
flabel metal2 87336 20798 87368 20814 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vom
flabel metal1 87524 19640 87566 19662 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vop
flabel metal2 74252 27128 74282 27156 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/VDD
flabel metal2 62452 7148 62526 7182 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vocm
flabel metal1 58602 4954 58634 4974 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/ibiasn
flabel metal1 67198 9466 67220 9494 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vom
flabel metal2 77354 11380 77386 11398 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vop
flabel metal1 88130 8502 88154 8532 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/VSS
flabel metal1 59620 1544 59656 1580 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/VSS
flabel metal1 88506 9350 88506 9350 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias3
flabel metal1 67094 13808 67094 13808 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmc_casc
flabel metal1 62010 5912 62010 5912 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmn_casc_tail2
flabel metal2 61882 6324 61882 6324 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmn_casc_tail1
flabel metal1 65082 6918 65082 6918 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmcn2_casc
flabel metal1 64612 6396 64612 6396 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmcn_casc
flabel metal1 64968 7052 64968 7052 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmcn1_casc
flabel metal2 63836 5024 63836 5024 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vfoldp
flabel metal1 62294 3038 62328 3070 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vip
flabel metal1 66046 3246 66072 3276 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vim
flabel metal1 69598 10104 69598 10104 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcascnp
flabel metal1 88250 9556 88250 9556 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcascnm
flabel metal1 88386 5324 88386 5324 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias4
flabel metal1 66956 12056 66956 12056 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vtail_casc
flabel metal1 88628 13722 88628 13726 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M3d
flabel metal1 87904 11204 87904 11204 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/M13d
flabel metal1 65542 3792 65542 3792 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vtail_casc
flabel metal1 62858 2724 62858 2724 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vfoldm
flabel metal1 55444 3634 55444 3634 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmn_casc_tail2
flabel metal1 56586 2904 56586 2904 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias2
flabel metal1 60658 2676 60658 2676 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vcmn_casc_tail1
flabel metal1 56872 14188 56872 14188 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias1
flabel metal1 58744 7514 58744 7514 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vbias2
flabel metal4 63608 21342 63684 21384 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vom
flabel metal4 54130 23836 54194 23876 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vop
flabel metal1 62500 6614 62528 6650 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vom
flabel metal2 64182 6550 64214 6572 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/vop
flabel metal1 82460 22146 82496 22174 1 FreeSans 480 0 0 0 diff_fold_casc_ota_1/VDD
flabel metal4 52550 27540 52550 28340 3 FreeSans 3200 0 0 0 diff_fold_casc_ota_1/VDD
flabel metal4 52550 -660 52550 140 3 FreeSans 3200 0 0 0 diff_fold_casc_ota_1/VSS
<< end >>
