magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< nwell >>
rect -2000 400 2000 2400
rect -2400 -400 2400 -40
rect -2400 -2400 -2000 -400
rect 2000 -2400 2400 -400
rect -2400 -2800 2400 -2400
<< pwell >>
rect -2400 2400 2400 2800
rect -2400 400 -2000 2400
rect 2000 400 2400 2400
rect -2400 40 2400 400
rect -2000 -2400 2000 -400
<< mvpsubdiff >>
rect -2334 2722 2334 2734
rect -2334 2562 -2100 2722
rect 2100 2562 2334 2722
rect -2334 2550 2334 2562
rect -2334 2500 -2150 2550
rect -2334 340 -2322 2500
rect -2162 340 -2150 2500
rect 2150 2500 2334 2550
rect -2334 290 -2150 340
rect 2150 340 2162 2500
rect 2322 340 2334 2500
rect 2150 290 2334 340
rect -2334 278 2334 290
rect -2334 118 -2100 278
rect 2100 118 2334 278
rect -2334 106 2334 118
rect -1934 -478 1934 -466
rect -1934 -638 -1700 -478
rect 1700 -638 1934 -478
rect -1934 -650 1934 -638
rect -1934 -700 -1750 -650
rect -1934 -2100 -1922 -700
rect -1762 -2100 -1750 -700
rect -1934 -2150 -1750 -2100
rect 1750 -700 1934 -650
rect 1750 -2100 1762 -700
rect 1922 -2100 1934 -700
rect 1750 -2150 1934 -2100
rect -1934 -2162 1934 -2150
rect -1934 -2322 -1700 -2162
rect 1700 -2322 1934 -2162
rect -1934 -2334 1934 -2322
<< mvnsubdiff >>
rect -1934 2322 1934 2334
rect -1934 2162 -1700 2322
rect 1700 2162 1934 2322
rect -1934 2150 1934 2162
rect -1934 2100 -1750 2150
rect -1934 700 -1922 2100
rect -1762 700 -1750 2100
rect -1934 650 -1750 700
rect 1750 2100 1934 2150
rect 1750 700 1762 2100
rect 1922 700 1934 2100
rect 1750 650 1934 700
rect -1934 638 1934 650
rect -1934 478 -1700 638
rect 1700 478 1934 638
rect -1934 466 1934 478
rect -2334 -118 2334 -106
rect -2334 -278 -2100 -118
rect 2100 -278 2334 -118
rect -2334 -290 2334 -278
rect -2334 -340 -2150 -290
rect -2334 -2500 -2322 -340
rect -2162 -2500 -2150 -340
rect 2150 -340 2334 -290
rect -2334 -2550 -2150 -2500
rect 2150 -2500 2162 -340
rect 2322 -2500 2334 -340
rect 2150 -2550 2334 -2500
rect -2334 -2562 2334 -2550
rect -2334 -2722 -2100 -2562
rect 2100 -2722 2334 -2562
rect -2334 -2734 2334 -2722
<< mvpsubdiffcont >>
rect -2100 2562 2100 2722
rect -2322 340 -2162 2500
rect 2162 340 2322 2500
rect -2100 118 2100 278
rect -1700 -638 1700 -478
rect -1922 -2100 -1762 -700
rect 1762 -2100 1922 -700
rect -1700 -2322 1700 -2162
<< mvnsubdiffcont >>
rect -1700 2162 1700 2322
rect -1922 700 -1762 2100
rect 1762 700 1922 2100
rect -1700 478 1700 638
rect -2100 -278 2100 -118
rect -2322 -2500 -2162 -340
rect 2162 -2500 2322 -340
rect -2100 -2722 2100 -2562
<< locali >>
rect -2322 2500 -2162 2722
rect 2162 2500 2322 2722
rect -1922 2100 -1762 2322
rect 1762 2100 1922 2322
rect -1922 478 -1762 700
rect 1762 478 1922 700
rect -2322 118 -2162 340
rect 2162 118 2322 340
rect -2322 -340 -2162 -118
rect 2162 -340 2322 -118
rect -1922 -700 -1762 -478
rect 1762 -700 1922 -478
rect -1922 -2322 -1762 -2100
rect 1762 -2322 1922 -2100
rect -2322 -2722 -2162 -2500
rect 2162 -2722 2322 -2500
<< viali >>
rect -2162 2562 -2100 2722
rect -2100 2562 2100 2722
rect 2100 2562 2162 2722
rect -2322 392 -2162 2448
rect -1762 2162 -1700 2322
rect -1700 2162 1700 2322
rect 1700 2162 1762 2322
rect -1922 714 -1762 2086
rect -1603 1947 1603 1981
rect 1762 714 1922 2086
rect -1762 478 -1700 638
rect -1700 478 1700 638
rect 1700 478 1762 638
rect 2162 392 2322 2448
rect -2162 118 -2100 278
rect -2100 118 2100 278
rect 2100 118 2162 278
rect -2162 -278 -2100 -118
rect -2100 -278 2100 -118
rect 2100 -278 2162 -118
rect -2322 -2448 -2162 -392
rect -1762 -638 -1700 -478
rect -1700 -638 1700 -478
rect 1700 -638 1762 -478
rect -1922 -2086 -1762 -714
rect -1603 -1972 1603 -1938
rect 1762 -2086 1922 -714
rect -1762 -2322 -1700 -2162
rect -1700 -2322 1700 -2162
rect 1700 -2322 1762 -2162
rect 2162 -2448 2322 -392
rect -2162 -2722 -2100 -2562
rect -2100 -2722 2100 -2562
rect 2100 -2722 2162 -2562
<< metal1 >>
rect -2400 3118 2400 3178
rect -2400 2838 -2340 3118
rect 2340 2838 2400 3118
rect -2400 2824 2400 2838
rect -2328 2722 2328 2728
rect -2328 2562 -2162 2722
rect 2162 2562 2328 2722
rect -2328 2460 2328 2562
rect -2328 2448 -2060 2460
rect -2328 392 -2322 2448
rect -2162 392 -2060 2448
rect 2061 2448 2328 2460
rect -2000 2328 2000 2400
rect -2000 2156 -1928 2328
rect 1928 2156 2000 2328
rect -2000 2086 -1756 2156
rect -2000 714 -1922 2086
rect -1762 714 -1756 2086
rect -1603 1987 -1557 2156
rect -1287 1987 -1241 2156
rect -971 1987 -925 2156
rect -655 1987 -609 2156
rect -339 1987 -293 2156
rect -23 1987 23 2156
rect 293 1987 339 2156
rect 609 1987 655 2156
rect 925 1987 971 2156
rect 1241 1987 1287 2156
rect 1557 1987 1603 2156
rect 1756 2086 2000 2156
rect -1615 1981 1615 1987
rect -1615 1947 -1603 1981
rect 1603 1947 1615 1981
rect -1615 1941 1615 1947
rect -1603 1900 -1557 1941
rect -1287 1900 -1241 1941
rect -971 1900 -925 1941
rect -655 1900 -609 1941
rect -339 1900 -293 1941
rect -23 1900 23 1941
rect 293 1900 339 1941
rect 609 1900 655 1941
rect 925 1900 971 1941
rect 1241 1900 1287 1941
rect 1557 1900 1603 1941
rect -1445 860 -1399 900
rect -1129 860 -1083 900
rect -813 860 -767 900
rect -497 860 -451 900
rect -181 860 -135 900
rect 135 860 181 900
rect 451 860 497 900
rect 767 860 813 900
rect 1083 860 1129 900
rect 1399 860 1445 900
rect -2000 644 -1756 714
rect -1455 700 -1445 860
rect -1045 700 1045 860
rect 1445 700 1455 860
rect 1756 714 1762 2086
rect 1922 714 2000 2086
rect 1756 644 2000 714
rect -2000 638 35 644
rect 955 638 2000 644
rect -2000 478 -1762 638
rect 1762 478 2000 638
rect -2000 472 35 478
rect 955 472 2000 478
rect -2000 400 2000 472
rect -2328 340 -2060 392
rect 2061 392 2162 2448
rect 2322 392 2328 2448
rect 2061 340 2328 392
rect -2328 284 2328 340
rect -2328 278 -965 284
rect -45 278 2328 284
rect -2328 118 -2162 278
rect 2162 118 2328 278
rect -2328 112 -965 118
rect -45 112 2328 118
rect -2328 40 2328 112
rect -2360 -112 2360 -40
rect -2360 -118 35 -112
rect 955 -118 2360 -112
rect -2360 -278 -2162 -118
rect 2162 -278 2360 -118
rect -2360 -284 35 -278
rect 955 -284 2360 -278
rect -2360 -340 2360 -284
rect -2360 -392 -2060 -340
rect -2360 -2448 -2322 -392
rect -2162 -2448 -2060 -392
rect 2060 -392 2360 -340
rect -2000 -472 2000 -400
rect -2000 -478 -965 -472
rect -45 -478 2000 -472
rect -2000 -638 -1762 -478
rect 1762 -638 2000 -478
rect -2000 -644 -965 -638
rect -45 -644 2000 -638
rect -2000 -714 -1750 -644
rect -2000 -2086 -1922 -714
rect -1762 -2086 -1750 -714
rect -1455 -860 -1445 -700
rect -1045 -860 1045 -700
rect 1445 -860 1455 -700
rect 1756 -714 2000 -644
rect -1445 -900 -1399 -860
rect -1129 -900 -1083 -860
rect -813 -900 -767 -860
rect -497 -900 -451 -860
rect -181 -900 -135 -860
rect 135 -900 181 -860
rect 451 -900 497 -860
rect 767 -900 813 -860
rect 1083 -900 1129 -860
rect 1399 -900 1445 -860
rect -1603 -1932 -1557 -1900
rect -1287 -1932 -1241 -1900
rect -971 -1932 -925 -1900
rect -655 -1932 -609 -1900
rect -339 -1932 -293 -1900
rect -23 -1932 23 -1900
rect 293 -1932 339 -1900
rect 609 -1932 655 -1900
rect 925 -1932 971 -1900
rect 1241 -1932 1287 -1900
rect 1557 -1932 1603 -1900
rect -1615 -1938 1615 -1932
rect -1615 -1972 -1603 -1938
rect 1603 -1972 1615 -1938
rect -1615 -1978 1615 -1972
rect -2000 -2156 -1750 -2086
rect -1603 -2156 -1557 -1978
rect -1287 -2156 -1241 -1978
rect -971 -2156 -925 -1978
rect -655 -2156 -609 -1978
rect -339 -2156 -293 -1978
rect -23 -2156 23 -1978
rect 293 -2156 339 -1978
rect 609 -2156 655 -1978
rect 925 -2156 971 -1978
rect 1241 -2156 1287 -1978
rect 1557 -2156 1603 -1978
rect 1756 -2086 1762 -714
rect 1922 -2086 2000 -714
rect 1756 -2156 2000 -2086
rect -2000 -2328 -1928 -2156
rect 1928 -2328 2000 -2156
rect -2000 -2400 2000 -2328
rect -2360 -2460 -2060 -2448
rect 2060 -2448 2162 -392
rect 2322 -2448 2360 -392
rect 2060 -2460 2360 -2448
rect -2360 -2562 2360 -2460
rect -2360 -2722 -2162 -2562
rect 2162 -2722 2360 -2562
rect -2360 -2728 2360 -2722
rect -2400 -2838 2400 -2825
rect -2400 -3118 -2340 -2838
rect 2340 -3118 2400 -2838
rect -2400 -3178 2400 -3118
<< via1 >>
rect -2340 2838 2340 3118
rect -1928 2322 1928 2328
rect -1928 2162 -1762 2322
rect -1762 2162 1762 2322
rect 1762 2162 1928 2322
rect -1928 2156 1928 2162
rect -1445 700 -1045 860
rect 1045 700 1445 860
rect 35 638 955 644
rect 35 478 955 638
rect 35 472 955 478
rect -965 278 -45 284
rect -965 118 -45 278
rect -965 112 -45 118
rect 35 -118 955 -112
rect 35 -278 955 -118
rect 35 -284 955 -278
rect -965 -478 -45 -472
rect -965 -638 -45 -478
rect -965 -644 -45 -638
rect -1445 -860 -1045 -700
rect 1045 -860 1445 -700
rect -1928 -2162 1928 -2156
rect -1928 -2322 -1762 -2162
rect -1762 -2322 1762 -2162
rect 1762 -2322 1928 -2162
rect -1928 -2328 1928 -2322
rect -2340 -3118 2340 -2838
<< metal2 >>
rect -2400 3118 2400 3178
rect -2400 2838 -2340 3118
rect 2340 2838 2400 3118
rect -2400 2328 2400 2838
rect -2400 2156 -1928 2328
rect 1928 2156 2400 2328
rect -2400 2150 2400 2156
rect -1928 2146 1928 2150
rect -1445 860 -1045 870
rect -1445 284 -1045 700
rect 1045 860 1445 870
rect 35 644 955 654
rect -2400 -284 -1045 284
rect -1445 -700 -1045 -284
rect -965 284 -45 294
rect -965 -472 -45 112
rect 35 -112 955 472
rect 35 -294 955 -284
rect 1045 284 1445 700
rect 1045 -284 2400 284
rect -965 -654 -45 -644
rect -1445 -870 -1045 -860
rect 1045 -700 1445 -284
rect 1045 -870 1445 -860
rect -1928 -2150 1928 -2146
rect -2400 -2156 2400 -2150
rect -2400 -2328 -1928 -2156
rect 1928 -2328 2400 -2156
rect -2400 -2838 2400 -2328
rect -2400 -3118 -2340 -2838
rect 2340 -3118 2400 -2838
rect -2400 -3178 2400 -3118
use sky130_fd_pr__pfet_g5v0d10v5_Q5DL9H  xm2
timestamp 1624477805
transform 1 0 0 0 1 1400
box -1675 -600 1675 600
use sky130_fd_pr__nfet_g5v0d10v5_ZGGKXL  xm1
timestamp 1624477805
transform 1 0 0 0 1 -1400
box -1609 -588 1609 588
<< labels >>
flabel metal2 -2400 -284 -2397 284 3 FreeSans 400 0 0 0 clamp
flabel metal2 -2392 -2814 -2386 -2808 1 FreeSans 480 0 0 0 VSS
flabel metal2 -2376 2812 -2370 2816 1 FreeSans 480 0 0 0 VDD
<< properties >>
string FIXED_BBOX -1842 -2242 1842 -558
<< end >>
