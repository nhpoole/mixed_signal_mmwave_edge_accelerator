* NGSPICE file created from diff_fold_casc_ota_flat.ext - technology: sky130A

.subckt diff_fold_casc_ota_flat vop vom vip vim vocm ibiasn VDD VSS
X0 vom vbias2 vfoldm VDD sky130_fd_pr__pfet_01v8 ad=5.22e+12p pd=3.948e+07u as=8.7e+12p ps=6.58e+07u w=3e+06u l=4.8e+06u
X1 vop vbias2 vfoldp VDD sky130_fd_pr__pfet_01v8 ad=5.22e+12p pd=3.948e+07u as=8.7e+12p ps=6.58e+07u w=3e+06u l=4.8e+06u
X2 VDD vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=4.147e+13p pd=3.1674e+08u as=4.06e+12p ps=3.206e+07u w=2e+06u l=800000u
X3 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=1.044e+13p pd=7.896e+07u as=4.176e+13p ps=3.1584e+08u w=3e+06u l=1.2e+06u
X4 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=2.61e+13p pd=1.974e+08u as=2.262e+13p ps=1.7108e+08u w=3e+06u l=4.8e+06u
X5 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=3.915e+13p pd=2.961e+08u as=3.48e+13p ps=2.632e+08u w=3e+06u l=4.8e+06u
X6 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=6.699e+13p pd=5.0666e+08u as=0p ps=0u w=3e+06u l=4.8e+06u
X7 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X8 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X9 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X10 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.044e+13p ps=7.896e+07u w=3e+06u l=1.2e+06u
X11 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X12 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X13 M13d M13d VSS VSS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=4.8e+06u
X14 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X15 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X16 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X17 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X18 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X19 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X20 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X21 vbias1 vbias2 M1d VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.632e+07u as=1.044e+13p ps=7.896e+07u w=3e+06u l=4.8e+06u
X22 VDD vcmcn_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=800000u
X23 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=1.044e+13p pd=7.896e+07u as=1.566e+13p ps=1.1844e+08u w=3e+06u l=4.8e+06u
X24 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=1.566e+13p pd=1.1844e+08u as=1.044e+13p ps=7.896e+07u w=3e+06u l=4.8e+06u
X25 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X26 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=8.7e+12p pd=6.58e+07u as=0p ps=0u w=3e+06u l=4.8e+06u
X27 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X28 M3d vbias2 M2d VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.632e+07u as=1.044e+13p ps=7.896e+07u w=3e+06u l=4.8e+06u
X29 vbias3 M3d vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+13p ps=9.212e+07u w=3e+06u l=4.8e+06u
X30 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X31 VDD vbias1 vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X32 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.566e+13p ps=1.1844e+08u w=3e+06u l=4.8e+06u
X33 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X34 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X35 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X36 vcmcn1_casc vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X37 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X38 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X39 vcmn_casc_tail1 vcmn_casc_tail1 vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=5.51e+12p pd=4.322e+07u as=0p ps=0u w=3e+06u l=4.8e+06u
X40 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X41 vcmc_casc vcmc_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X42 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X43 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X44 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X45 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X46 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X47 vom vom vom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X48 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X49 VDD vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=800000u
X50 vop vop vop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X51 vop vop vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X52 VDD vbias1 vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X53 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X54 VDD vbias1 vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X55 vcmc_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X56 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X57 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X58 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X59 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X60 VDD vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X61 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X62 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X63 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X64 VSS VSS vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X65 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X66 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X67 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X68 M1d M1d M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X69 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X70 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X71 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X72 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X73 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X74 VSS ibiasn vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.51e+12p ps=4.322e+07u w=3e+06u l=4.8e+06u
X75 VDD VDD M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X76 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X77 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X78 vcmc_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X79 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X80 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.29e+07u w=3e+06u l=4.8e+06u
X81 M2d M2d M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X82 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X83 vcmcn2_casc vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X84 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X85 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X86 VDD vbias1 vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X87 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X88 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X89 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X90 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X91 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X92 vcmcn_casc vom vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.58e+07u as=0p ps=0u w=1e+06u l=800000u
X93 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X94 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X95 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X96 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X97 vcmcn2_casc vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X98 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X99 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X100 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X101 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X102 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X103 vcmn_casc_tail1 vocm vcmcn1_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=800000u
X104 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X105 vcmcn_casc vcmcn_casc vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X106 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X107 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X108 VDD vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=800000u
X109 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X110 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X111 vcmn_casc_tail1 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X112 M1d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X113 VDD vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X114 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X115 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X116 VDD vbias1 M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=8.7e+12p ps=6.58e+07u w=3e+06u l=4.8e+06u
X117 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X118 vcmn_casc_tail1 vcmn_casc_tail1 vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X119 VDD vbias1 M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X120 vbias1 vbias2 M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X121 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X122 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X123 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X124 vcmcn2_casc vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X125 vcmn_casc_tail1 vop vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X126 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X127 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X128 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X129 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X130 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X131 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X132 vbias2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X133 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X134 M6d M6d M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X135 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X136 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X137 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X138 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X139 M1d M1d M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X140 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X141 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X142 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X143 M6d vbias2 M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.632e+07u w=3e+06u l=4.8e+06u
X144 vcmcn1_casc vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X145 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X146 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X147 M13d vbias2 M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X148 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X149 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X150 vcmn_casc_tail2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X151 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X152 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X153 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X154 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X155 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X156 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X157 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X158 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X159 vbias4 M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X160 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X161 M6d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X162 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X163 M6d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X164 M1d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X165 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X166 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X167 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X168 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X169 M2d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X170 vom vbias2 vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X171 vcmcn2_casc vocm vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=800000u
X172 M2d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X173 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X174 vop vbias2 vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X175 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X176 M1d vbias2 vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X177 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X178 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X179 VSS ibiasn vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X180 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X181 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X182 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X183 vcmcn1_casc vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X184 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X185 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X186 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X187 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X188 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X189 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X190 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X191 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X192 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X193 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X194 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X195 M2d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X196 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X197 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X198 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X199 VSS VSS M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X200 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X201 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X202 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X203 vcmcn_casc vcmcn_casc vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X204 M3d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X205 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X206 VDD vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X207 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X208 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X209 M13d vbias2 M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X210 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X211 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X212 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X213 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X214 M6d vbias2 M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X215 vcmcn_casc vom vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X216 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X217 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X218 vcmn_casc_tail2 vom vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X219 M2d vbias2 M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X220 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X221 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X222 VDD vbias1 M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X223 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X224 VDD vbias1 M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X225 VDD vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X226 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X227 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X228 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X229 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X230 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X231 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X232 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X233 vcmcn1_casc vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X234 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X235 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X236 vfoldm vbias2 vom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X237 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X238 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X239 vfoldp vbias2 vop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X240 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X241 vcmcn_casc vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X242 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X243 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X244 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X245 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X246 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X247 vfoldp vbias2 vop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X248 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X249 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X250 VSS vbias4 vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X251 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X252 vfoldm vbias2 vom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X253 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X254 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X255 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X256 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X257 VDD vbias1 M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X258 vcmn_casc_tail2 vocm vcmcn2_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X259 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X260 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X261 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X262 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X263 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X264 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X265 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X266 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X267 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X268 vcmcn1_casc vocm vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X269 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X270 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X271 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X272 vcmcn_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X273 M6d vbias2 M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X274 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X275 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X276 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X277 M13d vbias2 M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X278 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X279 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X280 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X281 M2d M2d M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X282 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X283 vbias4 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X284 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X285 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X286 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X287 vcmcn_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X288 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X289 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X290 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X291 M3d vbias2 M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X292 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X293 M2d M2d M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X294 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X295 vcmcn2_casc vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X296 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X297 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X298 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X299 vom vom vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X300 VDD vcmcn_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X301 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X302 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X303 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X304 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X305 VDD VDD vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X306 VDD vbias1 M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X307 VDD VDD vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X308 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X309 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X310 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X311 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X312 vop vop vop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X313 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X314 VDD vcmcn_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X315 vom vom vom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X316 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X317 VDD vbias1 vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X318 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X319 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X320 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X321 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X322 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X323 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X324 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X325 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X326 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X327 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X328 ibiasn ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X329 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X330 VDD VDD M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X331 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X332 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X333 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X334 VDD VDD M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X335 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X336 vcmn_casc_tail2 vcmn_casc_tail2 vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X337 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X338 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X339 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X340 vcmc_casc vcmc_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X341 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X342 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X343 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X344 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X345 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X346 M2d vbias2 M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X347 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X348 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X349 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X350 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X351 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X352 vcmc_casc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X353 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X354 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X355 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X356 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X357 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X358 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X359 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X360 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X361 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X362 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X363 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X364 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X365 vcmcn_casc vop vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X366 VDD vbias1 M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X367 vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X368 vcmc_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X369 VSS ibiasn vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X370 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X371 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X372 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X373 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X374 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X375 vcmn_casc_tail2 vocm vcmcn2_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X376 vcmcn_casc vcmcn_casc vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X377 M1d vbias2 vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X378 M6d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X379 M1d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X380 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X381 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X382 VDD vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X383 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X384 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X385 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X386 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X387 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X388 VSS ibiasn vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X389 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X390 M2d vbias2 M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X391 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X392 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X393 ibiasn ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X394 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X395 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X396 vcmn_casc_tail2 vcmn_casc_tail2 vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X397 vcmcn2_casc vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X398 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X399 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X400 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X401 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X402 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X403 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X404 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X405 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X406 VDD vcmcn_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X407 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X408 VDD vbias1 vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X409 VDD vbias1 vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X410 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X411 VDD vbias1 vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X412 VDD vbias1 vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X413 vcmn_casc_tail2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X414 M1d M1d M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X415 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X416 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X417 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X418 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X419 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X420 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X421 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X422 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X423 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X424 vfoldp vfoldp vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X425 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X426 VDD vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X427 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X428 vcmcn1_casc vocm vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X429 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X430 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X431 vbias2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X432 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X433 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X434 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X435 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X436 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X437 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X438 vcmcn2_casc vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X439 VDD vbias1 vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X440 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X441 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X442 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X443 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X444 VDD vbias1 vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X445 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X446 M3d vbias2 M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X447 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X448 vcmc_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X449 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X450 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X451 vcmcn_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X452 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X453 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X454 VSS ibiasn vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X455 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X456 vbias1 vbias2 M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X457 vcmcn1_casc vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X458 M6d M6d M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X459 vcmn_casc_tail2 vom vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X460 vcmn_casc_tail1 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X461 M2d M2d M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X462 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X463 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X464 vop VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X465 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X466 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X467 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X468 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X469 VDD vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X470 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X471 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X472 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X473 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X474 VDD vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X475 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X476 VSS ibiasn vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X477 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X478 VSS vbias4 vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X479 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X480 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X481 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X482 vfoldp vbias2 vop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X483 vtail_casc vim vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X484 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X485 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X486 vfoldm vbias2 vom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X487 vcmcn1_casc vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X488 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X489 a_4604_n20952# vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X490 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X491 vcmn_casc_tail1 vocm vcmcn1_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X492 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X493 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X494 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X495 VSS vcmc_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X496 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X497 VSS VSS vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X498 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X499 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X500 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X501 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X502 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X503 VDD vbias1 M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X504 VDD VDD vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X505 vcmcn2_casc vocm vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X506 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X507 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X508 VDD vbias1 M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X509 vcmcn_casc vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X510 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X511 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X512 M1d M1d M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X513 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X514 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X515 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X516 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X517 vcascnm vbias3 vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X518 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X519 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X520 VDD vbias1 vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X521 VDD vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X522 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X523 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X524 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X525 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X526 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X527 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X528 vcmcn_casc vcmcn_casc vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X529 vbias4 vbias4 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X530 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X531 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X532 vfoldm vfoldm vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X533 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X534 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X535 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X536 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X537 vcmcn_casc vop vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X538 vcmn_casc_tail1 vop vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X539 M1d vbias2 vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X540 vop vbias2 vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X541 vcmcn_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X542 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X543 VSS vbias4 vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X544 vcascnp vbias3 vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X545 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X546 M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X547 vom vbias2 vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X548 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X549 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X550 vom VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X551 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X552 M6d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X553 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X554 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X555 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X556 vtail_casc vip vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X557 vom vom vom VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X558 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X559 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X560 VSS vbias4 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X561 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X562 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X563 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X564 vbias3 M3d M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X565 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X566 vbias4 vbias4 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X567 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X568 a_4604_n20952# vbias3 vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X569 vfoldm vfoldm vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X570 VSS vcmc_casc vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X571 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X572 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X573 vfoldm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X574 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X575 vbias4 vbias3 a_4604_n20952# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X576 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X577 vfoldp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X578 vbias2 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X579 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X580 vfoldp vfoldp vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X581 M3d VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X582 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X583 vop vop vop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
C0 vfoldm M6d 10.15fF
C1 vfoldm vbias1 2.33fF
C2 M13d vtail_casc 0.04fF
C3 vcmcn1_casc vcmcn2_casc 13.41fF
C4 vbias3 vbias1 0.02fF
C5 M13d vfoldp 1.62fF
C6 vcmc_casc VDD 5.11fF
C7 M1d M3d 2.62fF
C8 vip vtail_casc 3.62fF
C9 vom vcascnp 3.37fF
C10 vbias2 M1d 6.85fF
C11 vfoldm vim 7.27fF
C12 vip vfoldp 9.23fF
C13 vop M13d 9.72fF
C14 VDD vfoldp 16.44fF
C15 vcmcn2_casc vom 2.96fF
C16 vcmcn1_casc vfoldm 0.08fF
C17 a_4604_n20952# vcascnp 6.65fF
C18 vcmcn1_casc vbias3 0.02fF
C19 vop VDD 5.44fF
C20 vcmc_casc vtail_casc 23.17fF
C21 M2d M6d 2.00fF
C22 vcmcn2_casc vcmcn_casc 6.63fF
C23 M2d vbias1 11.84fF
C24 vfoldm vom 2.33fF
C25 vop vocm 1.19fF
C26 vcmcn2_casc vbias2 2.34fF
C27 vcmn_casc_tail2 vcmcn2_casc 0.37fF
C28 vom vbias4 28.62fF
C29 vbias3 vom 5.67fF
C30 vtail_casc vfoldp 8.06fF
C31 VDD M1d 9.43fF
C32 vop vcmc_casc 4.23fF
C33 vop vtail_casc 1.62fF
C34 vbias3 a_4604_n20952# 7.49fF
C35 a_4604_n20952# vbias4 14.02fF
C36 vop vfoldp 0.18fF
C37 M6d vbias1 1.84fF
C38 vfoldm vcmcn_casc 0.12fF
C39 vfoldm M3d 0.12fF
C40 vfoldm vbias2 1.45fF
C41 vcmn_casc_tail2 vfoldm 0.03fF
C42 vbias3 vcmcn_casc 0.04fF
C43 vbias3 M3d 60.63fF
C44 vbias4 M3d 1.53fF
C45 vcmcn2_casc vip 0.22fF
C46 M1d vfoldp 6.26fF
C47 vcmcn2_casc VDD 5.31fF
C48 M2d vom 0.38fF
C49 vcascnm vom 18.97fF
C50 vcmcn1_casc vbias1 0.09fF
C51 vfoldm M13d 6.93fF
C52 vcmcn1_casc vcmn_casc_tail1 0.36fF
C53 vcmcn2_casc vocm 1.38fF
C54 vbias3 M13d 0.48fF
C55 M13d vbias4 0.04fF
C56 vop M1d 0.54fF
C57 vfoldm vip 3.11fF
C58 vcascnm a_4604_n20952# 9.83fF
C59 vcmcn2_casc vcmc_casc 0.16fF
C60 M6d vom 2.11fF
C61 vfoldm VDD 19.14fF
C62 vbias1 vom 0.93fF
C63 M2d M3d 1.87fF
C64 vbias2 M2d 1.06fF
C65 vcmn_casc_tail1 vom 0.10fF
C66 vcascnm M3d 0.69fF
C67 vcmcn2_casc vfoldp 2.70fF
C68 ibiasn vcmn_casc_tail1 1.79fF
C69 vfoldm vocm 0.02fF
C70 vop vcascnp 7.04fF
C71 vcmcn2_casc vop 0.60fF
C72 vbias1 vcmcn_casc 0.55fF
C73 vbias3 vcmc_casc 1.29fF
C74 vcmc_casc vbias4 36.08fF
C75 vbias2 M6d 1.00fF
C76 vbias1 M3d 5.14fF
C77 vcmcn1_casc vom 2.27fF
C78 vbias2 vbias1 11.85fF
C79 vcmn_casc_tail1 vcmcn_casc 0.97fF
C80 M2d M13d 0.70fF
C81 vfoldm vtail_casc 10.25fF
C82 vfoldm vfoldp 23.11fF
C83 vcascnm M13d 0.12fF
C84 vcmn_casc_tail1 vbias2 5.47fF
C85 vcmn_casc_tail2 vcmn_casc_tail1 3.28fF
C86 vbias3 vtail_casc 2.12fF
C87 vbias4 vtail_casc 28.15fF
C88 M2d VDD 8.52fF
C89 vfoldm vop 5.90fF
C90 vop vbias3 11.45fF
C91 vop vbias4 14.85fF
C92 vcmcn1_casc vcmcn_casc 16.79fF
C93 M6d M13d 0.56fF
C94 vcmcn1_casc vbias2 0.96fF
C95 a_4604_n20952# vom 8.05fF
C96 vfoldm M1d 13.09fF
C97 M6d VDD 10.55fF
C98 vcmn_casc_tail1 vip 0.02fF
C99 vcmcn_casc vom 7.09fF
C100 vbias1 VDD 19.60fF
C101 vom M3d 3.23fF
C102 vbias2 vom 5.46fF
C103 vcmn_casc_tail2 vom 0.45fF
C104 ibiasn vbias2 1.60fF
C105 vcmn_casc_tail2 ibiasn 3.91fF
C106 M2d vfoldp 1.90fF
C107 vim vip 3.15fF
C108 vcmn_casc_tail1 vocm 2.06fF
C109 vbias1 vcmc_casc 2.10fF
C110 vop M2d 14.54fF
C111 vop vcascnm 11.77fF
C112 vbias2 vcmcn_casc 0.63fF
C113 vbias4 vcascnp 17.91fF
C114 vcmn_casc_tail2 vcmcn_casc 1.11fF
C115 vcmcn1_casc VDD 8.62fF
C116 vbias3 vcascnp 18.64fF
C117 M13d vom 3.51fF
C118 vbias2 M3d 0.61fF
C119 M6d vfoldp 18.03fF
C120 vcmn_casc_tail2 vbias2 2.21fF
C121 vbias1 vfoldp 6.84fF
C122 vfoldm vcmcn2_casc 0.15fF
C123 vcmcn1_casc vocm 1.53fF
C124 vip vom 0.24fF
C125 M2d M1d 8.30fF
C126 vim vtail_casc 8.59fF
C127 vop M6d 0.31fF
C128 a_4604_n20952# M13d 1.44fF
C129 VDD vom 2.36fF
C130 vim vfoldp 3.14fF
C131 vop vbias1 2.53fF
C132 vcmcn1_casc vcmc_casc 0.86fF
C133 vop vcmn_casc_tail1 2.44fF
C134 M13d M3d 0.18fF
C135 vom vocm 4.79fF
C136 vbias2 M13d 1.61fF
C137 vcmcn1_casc vfoldp 0.08fF
C138 vbias3 vbias4 36.54fF
C139 M6d M1d 5.96fF
C140 vcmc_casc vom 5.06fF
C141 vbias2 vip 0.42fF
C142 vbias1 M1d 2.72fF
C143 VDD vcmcn_casc 15.75fF
C144 vcascnm vcascnp 12.37fF
C145 VDD M3d 1.56fF
C146 vbias2 VDD 11.06fF
C147 vcmcn1_casc vop 0.86fF
C148 vom vtail_casc 1.58fF
C149 vom vfoldp 2.90fF
C150 vcmcn_casc vocm 1.38fF
C151 vbias2 vocm 0.42fF
C152 vcmn_casc_tail2 vocm 2.22fF
C153 vcmc_casc vcmcn_casc 6.12fF
C154 vop vom 23.66fF
C155 vcmc_casc M3d 0.64fF
C156 vbias2 vcmc_casc 0.10fF
C157 VDD M13d 1.24fF
C158 vcmcn_casc vtail_casc 0.01fF
C159 vcmcn_casc vfoldp 0.12fF
C160 vtail_casc M3d 1.56fF
C161 vfoldm M2d 10.45fF
C162 vcmcn2_casc vbias1 0.08fF
C163 vbias2 vfoldp 2.32fF
C164 vbias3 vcascnm 10.63fF
C165 vcascnm vbias4 16.60fF
C166 vop a_4604_n20952# 19.89fF
C167 M1d vom 14.05fF
C168 vop vcmcn_casc 4.62fF
C169 vop M3d 0.98fF
C170 vop vbias2 1.14fF
C171 vcmn_casc_tail2 vop 0.69fF
.ends

