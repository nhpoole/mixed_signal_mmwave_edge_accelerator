magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -36 679 2240 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 2204 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 1998 1130 2032 1397
rect 2102 1322 2136 1397
rect 64 674 98 740
rect 1030 724 1064 1096
rect 1030 690 1081 724
rect 1030 318 1064 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 1998 17 2032 218
rect 2102 17 2136 92
rect 0 -17 2204 17
use nmos_m18_w2_000_sli_dli_da_p  nmos_m18_w2_000_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 51
box -26 -26 2012 456
use pmos_m18_w2_000_sli_dli_da_p  pmos_m18_w2_000_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 963
box -59 -56 2045 454
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 48 0 1 674
box 0 0 66 66
use contact_28  contact_28_0
timestamp 1624494425
transform 1 0 2094 0 1 51
box -26 -26 76 108
use contact_27  contact_27_0
timestamp 1624494425
transform 1 0 2094 0 1 1281
box -59 -43 109 125
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 1064 707 1064 707 4 Z
rlabel locali s 1102 0 1102 0 4 gnd
rlabel locali s 1102 1414 1102 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2204 1414
<< end >>
