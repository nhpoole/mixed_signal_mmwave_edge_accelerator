magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -11495 -1648 11495 1648
<< pwell >>
rect -10235 -326 10235 326
<< nmos >>
rect -10151 -300 -9191 300
rect -9133 -300 -8173 300
rect -8115 -300 -7155 300
rect -7097 -300 -6137 300
rect -6079 -300 -5119 300
rect -5061 -300 -4101 300
rect -4043 -300 -3083 300
rect -3025 -300 -2065 300
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
rect 2065 -300 3025 300
rect 3083 -300 4043 300
rect 4101 -300 5061 300
rect 5119 -300 6079 300
rect 6137 -300 7097 300
rect 7155 -300 8115 300
rect 8173 -300 9133 300
rect 9191 -300 10151 300
<< ndiff >>
rect -10209 255 -10151 300
rect -10209 221 -10197 255
rect -10163 221 -10151 255
rect -10209 187 -10151 221
rect -10209 153 -10197 187
rect -10163 153 -10151 187
rect -10209 119 -10151 153
rect -10209 85 -10197 119
rect -10163 85 -10151 119
rect -10209 51 -10151 85
rect -10209 17 -10197 51
rect -10163 17 -10151 51
rect -10209 -17 -10151 17
rect -10209 -51 -10197 -17
rect -10163 -51 -10151 -17
rect -10209 -85 -10151 -51
rect -10209 -119 -10197 -85
rect -10163 -119 -10151 -85
rect -10209 -153 -10151 -119
rect -10209 -187 -10197 -153
rect -10163 -187 -10151 -153
rect -10209 -221 -10151 -187
rect -10209 -255 -10197 -221
rect -10163 -255 -10151 -221
rect -10209 -300 -10151 -255
rect -9191 255 -9133 300
rect -9191 221 -9179 255
rect -9145 221 -9133 255
rect -9191 187 -9133 221
rect -9191 153 -9179 187
rect -9145 153 -9133 187
rect -9191 119 -9133 153
rect -9191 85 -9179 119
rect -9145 85 -9133 119
rect -9191 51 -9133 85
rect -9191 17 -9179 51
rect -9145 17 -9133 51
rect -9191 -17 -9133 17
rect -9191 -51 -9179 -17
rect -9145 -51 -9133 -17
rect -9191 -85 -9133 -51
rect -9191 -119 -9179 -85
rect -9145 -119 -9133 -85
rect -9191 -153 -9133 -119
rect -9191 -187 -9179 -153
rect -9145 -187 -9133 -153
rect -9191 -221 -9133 -187
rect -9191 -255 -9179 -221
rect -9145 -255 -9133 -221
rect -9191 -300 -9133 -255
rect -8173 255 -8115 300
rect -8173 221 -8161 255
rect -8127 221 -8115 255
rect -8173 187 -8115 221
rect -8173 153 -8161 187
rect -8127 153 -8115 187
rect -8173 119 -8115 153
rect -8173 85 -8161 119
rect -8127 85 -8115 119
rect -8173 51 -8115 85
rect -8173 17 -8161 51
rect -8127 17 -8115 51
rect -8173 -17 -8115 17
rect -8173 -51 -8161 -17
rect -8127 -51 -8115 -17
rect -8173 -85 -8115 -51
rect -8173 -119 -8161 -85
rect -8127 -119 -8115 -85
rect -8173 -153 -8115 -119
rect -8173 -187 -8161 -153
rect -8127 -187 -8115 -153
rect -8173 -221 -8115 -187
rect -8173 -255 -8161 -221
rect -8127 -255 -8115 -221
rect -8173 -300 -8115 -255
rect -7155 255 -7097 300
rect -7155 221 -7143 255
rect -7109 221 -7097 255
rect -7155 187 -7097 221
rect -7155 153 -7143 187
rect -7109 153 -7097 187
rect -7155 119 -7097 153
rect -7155 85 -7143 119
rect -7109 85 -7097 119
rect -7155 51 -7097 85
rect -7155 17 -7143 51
rect -7109 17 -7097 51
rect -7155 -17 -7097 17
rect -7155 -51 -7143 -17
rect -7109 -51 -7097 -17
rect -7155 -85 -7097 -51
rect -7155 -119 -7143 -85
rect -7109 -119 -7097 -85
rect -7155 -153 -7097 -119
rect -7155 -187 -7143 -153
rect -7109 -187 -7097 -153
rect -7155 -221 -7097 -187
rect -7155 -255 -7143 -221
rect -7109 -255 -7097 -221
rect -7155 -300 -7097 -255
rect -6137 255 -6079 300
rect -6137 221 -6125 255
rect -6091 221 -6079 255
rect -6137 187 -6079 221
rect -6137 153 -6125 187
rect -6091 153 -6079 187
rect -6137 119 -6079 153
rect -6137 85 -6125 119
rect -6091 85 -6079 119
rect -6137 51 -6079 85
rect -6137 17 -6125 51
rect -6091 17 -6079 51
rect -6137 -17 -6079 17
rect -6137 -51 -6125 -17
rect -6091 -51 -6079 -17
rect -6137 -85 -6079 -51
rect -6137 -119 -6125 -85
rect -6091 -119 -6079 -85
rect -6137 -153 -6079 -119
rect -6137 -187 -6125 -153
rect -6091 -187 -6079 -153
rect -6137 -221 -6079 -187
rect -6137 -255 -6125 -221
rect -6091 -255 -6079 -221
rect -6137 -300 -6079 -255
rect -5119 255 -5061 300
rect -5119 221 -5107 255
rect -5073 221 -5061 255
rect -5119 187 -5061 221
rect -5119 153 -5107 187
rect -5073 153 -5061 187
rect -5119 119 -5061 153
rect -5119 85 -5107 119
rect -5073 85 -5061 119
rect -5119 51 -5061 85
rect -5119 17 -5107 51
rect -5073 17 -5061 51
rect -5119 -17 -5061 17
rect -5119 -51 -5107 -17
rect -5073 -51 -5061 -17
rect -5119 -85 -5061 -51
rect -5119 -119 -5107 -85
rect -5073 -119 -5061 -85
rect -5119 -153 -5061 -119
rect -5119 -187 -5107 -153
rect -5073 -187 -5061 -153
rect -5119 -221 -5061 -187
rect -5119 -255 -5107 -221
rect -5073 -255 -5061 -221
rect -5119 -300 -5061 -255
rect -4101 255 -4043 300
rect -4101 221 -4089 255
rect -4055 221 -4043 255
rect -4101 187 -4043 221
rect -4101 153 -4089 187
rect -4055 153 -4043 187
rect -4101 119 -4043 153
rect -4101 85 -4089 119
rect -4055 85 -4043 119
rect -4101 51 -4043 85
rect -4101 17 -4089 51
rect -4055 17 -4043 51
rect -4101 -17 -4043 17
rect -4101 -51 -4089 -17
rect -4055 -51 -4043 -17
rect -4101 -85 -4043 -51
rect -4101 -119 -4089 -85
rect -4055 -119 -4043 -85
rect -4101 -153 -4043 -119
rect -4101 -187 -4089 -153
rect -4055 -187 -4043 -153
rect -4101 -221 -4043 -187
rect -4101 -255 -4089 -221
rect -4055 -255 -4043 -221
rect -4101 -300 -4043 -255
rect -3083 255 -3025 300
rect -3083 221 -3071 255
rect -3037 221 -3025 255
rect -3083 187 -3025 221
rect -3083 153 -3071 187
rect -3037 153 -3025 187
rect -3083 119 -3025 153
rect -3083 85 -3071 119
rect -3037 85 -3025 119
rect -3083 51 -3025 85
rect -3083 17 -3071 51
rect -3037 17 -3025 51
rect -3083 -17 -3025 17
rect -3083 -51 -3071 -17
rect -3037 -51 -3025 -17
rect -3083 -85 -3025 -51
rect -3083 -119 -3071 -85
rect -3037 -119 -3025 -85
rect -3083 -153 -3025 -119
rect -3083 -187 -3071 -153
rect -3037 -187 -3025 -153
rect -3083 -221 -3025 -187
rect -3083 -255 -3071 -221
rect -3037 -255 -3025 -221
rect -3083 -300 -3025 -255
rect -2065 255 -2007 300
rect -2065 221 -2053 255
rect -2019 221 -2007 255
rect -2065 187 -2007 221
rect -2065 153 -2053 187
rect -2019 153 -2007 187
rect -2065 119 -2007 153
rect -2065 85 -2053 119
rect -2019 85 -2007 119
rect -2065 51 -2007 85
rect -2065 17 -2053 51
rect -2019 17 -2007 51
rect -2065 -17 -2007 17
rect -2065 -51 -2053 -17
rect -2019 -51 -2007 -17
rect -2065 -85 -2007 -51
rect -2065 -119 -2053 -85
rect -2019 -119 -2007 -85
rect -2065 -153 -2007 -119
rect -2065 -187 -2053 -153
rect -2019 -187 -2007 -153
rect -2065 -221 -2007 -187
rect -2065 -255 -2053 -221
rect -2019 -255 -2007 -221
rect -2065 -300 -2007 -255
rect -1047 255 -989 300
rect -1047 221 -1035 255
rect -1001 221 -989 255
rect -1047 187 -989 221
rect -1047 153 -1035 187
rect -1001 153 -989 187
rect -1047 119 -989 153
rect -1047 85 -1035 119
rect -1001 85 -989 119
rect -1047 51 -989 85
rect -1047 17 -1035 51
rect -1001 17 -989 51
rect -1047 -17 -989 17
rect -1047 -51 -1035 -17
rect -1001 -51 -989 -17
rect -1047 -85 -989 -51
rect -1047 -119 -1035 -85
rect -1001 -119 -989 -85
rect -1047 -153 -989 -119
rect -1047 -187 -1035 -153
rect -1001 -187 -989 -153
rect -1047 -221 -989 -187
rect -1047 -255 -1035 -221
rect -1001 -255 -989 -221
rect -1047 -300 -989 -255
rect -29 255 29 300
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -300 29 -255
rect 989 255 1047 300
rect 989 221 1001 255
rect 1035 221 1047 255
rect 989 187 1047 221
rect 989 153 1001 187
rect 1035 153 1047 187
rect 989 119 1047 153
rect 989 85 1001 119
rect 1035 85 1047 119
rect 989 51 1047 85
rect 989 17 1001 51
rect 1035 17 1047 51
rect 989 -17 1047 17
rect 989 -51 1001 -17
rect 1035 -51 1047 -17
rect 989 -85 1047 -51
rect 989 -119 1001 -85
rect 1035 -119 1047 -85
rect 989 -153 1047 -119
rect 989 -187 1001 -153
rect 1035 -187 1047 -153
rect 989 -221 1047 -187
rect 989 -255 1001 -221
rect 1035 -255 1047 -221
rect 989 -300 1047 -255
rect 2007 255 2065 300
rect 2007 221 2019 255
rect 2053 221 2065 255
rect 2007 187 2065 221
rect 2007 153 2019 187
rect 2053 153 2065 187
rect 2007 119 2065 153
rect 2007 85 2019 119
rect 2053 85 2065 119
rect 2007 51 2065 85
rect 2007 17 2019 51
rect 2053 17 2065 51
rect 2007 -17 2065 17
rect 2007 -51 2019 -17
rect 2053 -51 2065 -17
rect 2007 -85 2065 -51
rect 2007 -119 2019 -85
rect 2053 -119 2065 -85
rect 2007 -153 2065 -119
rect 2007 -187 2019 -153
rect 2053 -187 2065 -153
rect 2007 -221 2065 -187
rect 2007 -255 2019 -221
rect 2053 -255 2065 -221
rect 2007 -300 2065 -255
rect 3025 255 3083 300
rect 3025 221 3037 255
rect 3071 221 3083 255
rect 3025 187 3083 221
rect 3025 153 3037 187
rect 3071 153 3083 187
rect 3025 119 3083 153
rect 3025 85 3037 119
rect 3071 85 3083 119
rect 3025 51 3083 85
rect 3025 17 3037 51
rect 3071 17 3083 51
rect 3025 -17 3083 17
rect 3025 -51 3037 -17
rect 3071 -51 3083 -17
rect 3025 -85 3083 -51
rect 3025 -119 3037 -85
rect 3071 -119 3083 -85
rect 3025 -153 3083 -119
rect 3025 -187 3037 -153
rect 3071 -187 3083 -153
rect 3025 -221 3083 -187
rect 3025 -255 3037 -221
rect 3071 -255 3083 -221
rect 3025 -300 3083 -255
rect 4043 255 4101 300
rect 4043 221 4055 255
rect 4089 221 4101 255
rect 4043 187 4101 221
rect 4043 153 4055 187
rect 4089 153 4101 187
rect 4043 119 4101 153
rect 4043 85 4055 119
rect 4089 85 4101 119
rect 4043 51 4101 85
rect 4043 17 4055 51
rect 4089 17 4101 51
rect 4043 -17 4101 17
rect 4043 -51 4055 -17
rect 4089 -51 4101 -17
rect 4043 -85 4101 -51
rect 4043 -119 4055 -85
rect 4089 -119 4101 -85
rect 4043 -153 4101 -119
rect 4043 -187 4055 -153
rect 4089 -187 4101 -153
rect 4043 -221 4101 -187
rect 4043 -255 4055 -221
rect 4089 -255 4101 -221
rect 4043 -300 4101 -255
rect 5061 255 5119 300
rect 5061 221 5073 255
rect 5107 221 5119 255
rect 5061 187 5119 221
rect 5061 153 5073 187
rect 5107 153 5119 187
rect 5061 119 5119 153
rect 5061 85 5073 119
rect 5107 85 5119 119
rect 5061 51 5119 85
rect 5061 17 5073 51
rect 5107 17 5119 51
rect 5061 -17 5119 17
rect 5061 -51 5073 -17
rect 5107 -51 5119 -17
rect 5061 -85 5119 -51
rect 5061 -119 5073 -85
rect 5107 -119 5119 -85
rect 5061 -153 5119 -119
rect 5061 -187 5073 -153
rect 5107 -187 5119 -153
rect 5061 -221 5119 -187
rect 5061 -255 5073 -221
rect 5107 -255 5119 -221
rect 5061 -300 5119 -255
rect 6079 255 6137 300
rect 6079 221 6091 255
rect 6125 221 6137 255
rect 6079 187 6137 221
rect 6079 153 6091 187
rect 6125 153 6137 187
rect 6079 119 6137 153
rect 6079 85 6091 119
rect 6125 85 6137 119
rect 6079 51 6137 85
rect 6079 17 6091 51
rect 6125 17 6137 51
rect 6079 -17 6137 17
rect 6079 -51 6091 -17
rect 6125 -51 6137 -17
rect 6079 -85 6137 -51
rect 6079 -119 6091 -85
rect 6125 -119 6137 -85
rect 6079 -153 6137 -119
rect 6079 -187 6091 -153
rect 6125 -187 6137 -153
rect 6079 -221 6137 -187
rect 6079 -255 6091 -221
rect 6125 -255 6137 -221
rect 6079 -300 6137 -255
rect 7097 255 7155 300
rect 7097 221 7109 255
rect 7143 221 7155 255
rect 7097 187 7155 221
rect 7097 153 7109 187
rect 7143 153 7155 187
rect 7097 119 7155 153
rect 7097 85 7109 119
rect 7143 85 7155 119
rect 7097 51 7155 85
rect 7097 17 7109 51
rect 7143 17 7155 51
rect 7097 -17 7155 17
rect 7097 -51 7109 -17
rect 7143 -51 7155 -17
rect 7097 -85 7155 -51
rect 7097 -119 7109 -85
rect 7143 -119 7155 -85
rect 7097 -153 7155 -119
rect 7097 -187 7109 -153
rect 7143 -187 7155 -153
rect 7097 -221 7155 -187
rect 7097 -255 7109 -221
rect 7143 -255 7155 -221
rect 7097 -300 7155 -255
rect 8115 255 8173 300
rect 8115 221 8127 255
rect 8161 221 8173 255
rect 8115 187 8173 221
rect 8115 153 8127 187
rect 8161 153 8173 187
rect 8115 119 8173 153
rect 8115 85 8127 119
rect 8161 85 8173 119
rect 8115 51 8173 85
rect 8115 17 8127 51
rect 8161 17 8173 51
rect 8115 -17 8173 17
rect 8115 -51 8127 -17
rect 8161 -51 8173 -17
rect 8115 -85 8173 -51
rect 8115 -119 8127 -85
rect 8161 -119 8173 -85
rect 8115 -153 8173 -119
rect 8115 -187 8127 -153
rect 8161 -187 8173 -153
rect 8115 -221 8173 -187
rect 8115 -255 8127 -221
rect 8161 -255 8173 -221
rect 8115 -300 8173 -255
rect 9133 255 9191 300
rect 9133 221 9145 255
rect 9179 221 9191 255
rect 9133 187 9191 221
rect 9133 153 9145 187
rect 9179 153 9191 187
rect 9133 119 9191 153
rect 9133 85 9145 119
rect 9179 85 9191 119
rect 9133 51 9191 85
rect 9133 17 9145 51
rect 9179 17 9191 51
rect 9133 -17 9191 17
rect 9133 -51 9145 -17
rect 9179 -51 9191 -17
rect 9133 -85 9191 -51
rect 9133 -119 9145 -85
rect 9179 -119 9191 -85
rect 9133 -153 9191 -119
rect 9133 -187 9145 -153
rect 9179 -187 9191 -153
rect 9133 -221 9191 -187
rect 9133 -255 9145 -221
rect 9179 -255 9191 -221
rect 9133 -300 9191 -255
rect 10151 255 10209 300
rect 10151 221 10163 255
rect 10197 221 10209 255
rect 10151 187 10209 221
rect 10151 153 10163 187
rect 10197 153 10209 187
rect 10151 119 10209 153
rect 10151 85 10163 119
rect 10197 85 10209 119
rect 10151 51 10209 85
rect 10151 17 10163 51
rect 10197 17 10209 51
rect 10151 -17 10209 17
rect 10151 -51 10163 -17
rect 10197 -51 10209 -17
rect 10151 -85 10209 -51
rect 10151 -119 10163 -85
rect 10197 -119 10209 -85
rect 10151 -153 10209 -119
rect 10151 -187 10163 -153
rect 10197 -187 10209 -153
rect 10151 -221 10209 -187
rect 10151 -255 10163 -221
rect 10197 -255 10209 -221
rect 10151 -300 10209 -255
<< ndiffc >>
rect -10197 221 -10163 255
rect -10197 153 -10163 187
rect -10197 85 -10163 119
rect -10197 17 -10163 51
rect -10197 -51 -10163 -17
rect -10197 -119 -10163 -85
rect -10197 -187 -10163 -153
rect -10197 -255 -10163 -221
rect -9179 221 -9145 255
rect -9179 153 -9145 187
rect -9179 85 -9145 119
rect -9179 17 -9145 51
rect -9179 -51 -9145 -17
rect -9179 -119 -9145 -85
rect -9179 -187 -9145 -153
rect -9179 -255 -9145 -221
rect -8161 221 -8127 255
rect -8161 153 -8127 187
rect -8161 85 -8127 119
rect -8161 17 -8127 51
rect -8161 -51 -8127 -17
rect -8161 -119 -8127 -85
rect -8161 -187 -8127 -153
rect -8161 -255 -8127 -221
rect -7143 221 -7109 255
rect -7143 153 -7109 187
rect -7143 85 -7109 119
rect -7143 17 -7109 51
rect -7143 -51 -7109 -17
rect -7143 -119 -7109 -85
rect -7143 -187 -7109 -153
rect -7143 -255 -7109 -221
rect -6125 221 -6091 255
rect -6125 153 -6091 187
rect -6125 85 -6091 119
rect -6125 17 -6091 51
rect -6125 -51 -6091 -17
rect -6125 -119 -6091 -85
rect -6125 -187 -6091 -153
rect -6125 -255 -6091 -221
rect -5107 221 -5073 255
rect -5107 153 -5073 187
rect -5107 85 -5073 119
rect -5107 17 -5073 51
rect -5107 -51 -5073 -17
rect -5107 -119 -5073 -85
rect -5107 -187 -5073 -153
rect -5107 -255 -5073 -221
rect -4089 221 -4055 255
rect -4089 153 -4055 187
rect -4089 85 -4055 119
rect -4089 17 -4055 51
rect -4089 -51 -4055 -17
rect -4089 -119 -4055 -85
rect -4089 -187 -4055 -153
rect -4089 -255 -4055 -221
rect -3071 221 -3037 255
rect -3071 153 -3037 187
rect -3071 85 -3037 119
rect -3071 17 -3037 51
rect -3071 -51 -3037 -17
rect -3071 -119 -3037 -85
rect -3071 -187 -3037 -153
rect -3071 -255 -3037 -221
rect -2053 221 -2019 255
rect -2053 153 -2019 187
rect -2053 85 -2019 119
rect -2053 17 -2019 51
rect -2053 -51 -2019 -17
rect -2053 -119 -2019 -85
rect -2053 -187 -2019 -153
rect -2053 -255 -2019 -221
rect -1035 221 -1001 255
rect -1035 153 -1001 187
rect -1035 85 -1001 119
rect -1035 17 -1001 51
rect -1035 -51 -1001 -17
rect -1035 -119 -1001 -85
rect -1035 -187 -1001 -153
rect -1035 -255 -1001 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 1001 221 1035 255
rect 1001 153 1035 187
rect 1001 85 1035 119
rect 1001 17 1035 51
rect 1001 -51 1035 -17
rect 1001 -119 1035 -85
rect 1001 -187 1035 -153
rect 1001 -255 1035 -221
rect 2019 221 2053 255
rect 2019 153 2053 187
rect 2019 85 2053 119
rect 2019 17 2053 51
rect 2019 -51 2053 -17
rect 2019 -119 2053 -85
rect 2019 -187 2053 -153
rect 2019 -255 2053 -221
rect 3037 221 3071 255
rect 3037 153 3071 187
rect 3037 85 3071 119
rect 3037 17 3071 51
rect 3037 -51 3071 -17
rect 3037 -119 3071 -85
rect 3037 -187 3071 -153
rect 3037 -255 3071 -221
rect 4055 221 4089 255
rect 4055 153 4089 187
rect 4055 85 4089 119
rect 4055 17 4089 51
rect 4055 -51 4089 -17
rect 4055 -119 4089 -85
rect 4055 -187 4089 -153
rect 4055 -255 4089 -221
rect 5073 221 5107 255
rect 5073 153 5107 187
rect 5073 85 5107 119
rect 5073 17 5107 51
rect 5073 -51 5107 -17
rect 5073 -119 5107 -85
rect 5073 -187 5107 -153
rect 5073 -255 5107 -221
rect 6091 221 6125 255
rect 6091 153 6125 187
rect 6091 85 6125 119
rect 6091 17 6125 51
rect 6091 -51 6125 -17
rect 6091 -119 6125 -85
rect 6091 -187 6125 -153
rect 6091 -255 6125 -221
rect 7109 221 7143 255
rect 7109 153 7143 187
rect 7109 85 7143 119
rect 7109 17 7143 51
rect 7109 -51 7143 -17
rect 7109 -119 7143 -85
rect 7109 -187 7143 -153
rect 7109 -255 7143 -221
rect 8127 221 8161 255
rect 8127 153 8161 187
rect 8127 85 8161 119
rect 8127 17 8161 51
rect 8127 -51 8161 -17
rect 8127 -119 8161 -85
rect 8127 -187 8161 -153
rect 8127 -255 8161 -221
rect 9145 221 9179 255
rect 9145 153 9179 187
rect 9145 85 9179 119
rect 9145 17 9179 51
rect 9145 -51 9179 -17
rect 9145 -119 9179 -85
rect 9145 -187 9179 -153
rect 9145 -255 9179 -221
rect 10163 221 10197 255
rect 10163 153 10197 187
rect 10163 85 10197 119
rect 10163 17 10197 51
rect 10163 -51 10197 -17
rect 10163 -119 10197 -85
rect 10163 -187 10197 -153
rect 10163 -255 10197 -221
<< poly >>
rect -9965 372 -9377 388
rect -9965 355 -9926 372
rect -10151 338 -9926 355
rect -9892 338 -9858 372
rect -9824 338 -9790 372
rect -9756 338 -9722 372
rect -9688 338 -9654 372
rect -9620 338 -9586 372
rect -9552 338 -9518 372
rect -9484 338 -9450 372
rect -9416 355 -9377 372
rect -8947 372 -8359 388
rect -8947 355 -8908 372
rect -9416 338 -9191 355
rect -10151 300 -9191 338
rect -9133 338 -8908 355
rect -8874 338 -8840 372
rect -8806 338 -8772 372
rect -8738 338 -8704 372
rect -8670 338 -8636 372
rect -8602 338 -8568 372
rect -8534 338 -8500 372
rect -8466 338 -8432 372
rect -8398 355 -8359 372
rect -7929 372 -7341 388
rect -7929 355 -7890 372
rect -8398 338 -8173 355
rect -9133 300 -8173 338
rect -8115 338 -7890 355
rect -7856 338 -7822 372
rect -7788 338 -7754 372
rect -7720 338 -7686 372
rect -7652 338 -7618 372
rect -7584 338 -7550 372
rect -7516 338 -7482 372
rect -7448 338 -7414 372
rect -7380 355 -7341 372
rect -6911 372 -6323 388
rect -6911 355 -6872 372
rect -7380 338 -7155 355
rect -8115 300 -7155 338
rect -7097 338 -6872 355
rect -6838 338 -6804 372
rect -6770 338 -6736 372
rect -6702 338 -6668 372
rect -6634 338 -6600 372
rect -6566 338 -6532 372
rect -6498 338 -6464 372
rect -6430 338 -6396 372
rect -6362 355 -6323 372
rect -5893 372 -5305 388
rect -5893 355 -5854 372
rect -6362 338 -6137 355
rect -7097 300 -6137 338
rect -6079 338 -5854 355
rect -5820 338 -5786 372
rect -5752 338 -5718 372
rect -5684 338 -5650 372
rect -5616 338 -5582 372
rect -5548 338 -5514 372
rect -5480 338 -5446 372
rect -5412 338 -5378 372
rect -5344 355 -5305 372
rect -4875 372 -4287 388
rect -4875 355 -4836 372
rect -5344 338 -5119 355
rect -6079 300 -5119 338
rect -5061 338 -4836 355
rect -4802 338 -4768 372
rect -4734 338 -4700 372
rect -4666 338 -4632 372
rect -4598 338 -4564 372
rect -4530 338 -4496 372
rect -4462 338 -4428 372
rect -4394 338 -4360 372
rect -4326 355 -4287 372
rect -3857 372 -3269 388
rect -3857 355 -3818 372
rect -4326 338 -4101 355
rect -5061 300 -4101 338
rect -4043 338 -3818 355
rect -3784 338 -3750 372
rect -3716 338 -3682 372
rect -3648 338 -3614 372
rect -3580 338 -3546 372
rect -3512 338 -3478 372
rect -3444 338 -3410 372
rect -3376 338 -3342 372
rect -3308 355 -3269 372
rect -2839 372 -2251 388
rect -2839 355 -2800 372
rect -3308 338 -3083 355
rect -4043 300 -3083 338
rect -3025 338 -2800 355
rect -2766 338 -2732 372
rect -2698 338 -2664 372
rect -2630 338 -2596 372
rect -2562 338 -2528 372
rect -2494 338 -2460 372
rect -2426 338 -2392 372
rect -2358 338 -2324 372
rect -2290 355 -2251 372
rect -1821 372 -1233 388
rect -1821 355 -1782 372
rect -2290 338 -2065 355
rect -3025 300 -2065 338
rect -2007 338 -1782 355
rect -1748 338 -1714 372
rect -1680 338 -1646 372
rect -1612 338 -1578 372
rect -1544 338 -1510 372
rect -1476 338 -1442 372
rect -1408 338 -1374 372
rect -1340 338 -1306 372
rect -1272 355 -1233 372
rect -803 372 -215 388
rect -803 355 -764 372
rect -1272 338 -1047 355
rect -2007 300 -1047 338
rect -989 338 -764 355
rect -730 338 -696 372
rect -662 338 -628 372
rect -594 338 -560 372
rect -526 338 -492 372
rect -458 338 -424 372
rect -390 338 -356 372
rect -322 338 -288 372
rect -254 355 -215 372
rect 215 372 803 388
rect 215 355 254 372
rect -254 338 -29 355
rect -989 300 -29 338
rect 29 338 254 355
rect 288 338 322 372
rect 356 338 390 372
rect 424 338 458 372
rect 492 338 526 372
rect 560 338 594 372
rect 628 338 662 372
rect 696 338 730 372
rect 764 355 803 372
rect 1233 372 1821 388
rect 1233 355 1272 372
rect 764 338 989 355
rect 29 300 989 338
rect 1047 338 1272 355
rect 1306 338 1340 372
rect 1374 338 1408 372
rect 1442 338 1476 372
rect 1510 338 1544 372
rect 1578 338 1612 372
rect 1646 338 1680 372
rect 1714 338 1748 372
rect 1782 355 1821 372
rect 2251 372 2839 388
rect 2251 355 2290 372
rect 1782 338 2007 355
rect 1047 300 2007 338
rect 2065 338 2290 355
rect 2324 338 2358 372
rect 2392 338 2426 372
rect 2460 338 2494 372
rect 2528 338 2562 372
rect 2596 338 2630 372
rect 2664 338 2698 372
rect 2732 338 2766 372
rect 2800 355 2839 372
rect 3269 372 3857 388
rect 3269 355 3308 372
rect 2800 338 3025 355
rect 2065 300 3025 338
rect 3083 338 3308 355
rect 3342 338 3376 372
rect 3410 338 3444 372
rect 3478 338 3512 372
rect 3546 338 3580 372
rect 3614 338 3648 372
rect 3682 338 3716 372
rect 3750 338 3784 372
rect 3818 355 3857 372
rect 4287 372 4875 388
rect 4287 355 4326 372
rect 3818 338 4043 355
rect 3083 300 4043 338
rect 4101 338 4326 355
rect 4360 338 4394 372
rect 4428 338 4462 372
rect 4496 338 4530 372
rect 4564 338 4598 372
rect 4632 338 4666 372
rect 4700 338 4734 372
rect 4768 338 4802 372
rect 4836 355 4875 372
rect 5305 372 5893 388
rect 5305 355 5344 372
rect 4836 338 5061 355
rect 4101 300 5061 338
rect 5119 338 5344 355
rect 5378 338 5412 372
rect 5446 338 5480 372
rect 5514 338 5548 372
rect 5582 338 5616 372
rect 5650 338 5684 372
rect 5718 338 5752 372
rect 5786 338 5820 372
rect 5854 355 5893 372
rect 6323 372 6911 388
rect 6323 355 6362 372
rect 5854 338 6079 355
rect 5119 300 6079 338
rect 6137 338 6362 355
rect 6396 338 6430 372
rect 6464 338 6498 372
rect 6532 338 6566 372
rect 6600 338 6634 372
rect 6668 338 6702 372
rect 6736 338 6770 372
rect 6804 338 6838 372
rect 6872 355 6911 372
rect 7341 372 7929 388
rect 7341 355 7380 372
rect 6872 338 7097 355
rect 6137 300 7097 338
rect 7155 338 7380 355
rect 7414 338 7448 372
rect 7482 338 7516 372
rect 7550 338 7584 372
rect 7618 338 7652 372
rect 7686 338 7720 372
rect 7754 338 7788 372
rect 7822 338 7856 372
rect 7890 355 7929 372
rect 8359 372 8947 388
rect 8359 355 8398 372
rect 7890 338 8115 355
rect 7155 300 8115 338
rect 8173 338 8398 355
rect 8432 338 8466 372
rect 8500 338 8534 372
rect 8568 338 8602 372
rect 8636 338 8670 372
rect 8704 338 8738 372
rect 8772 338 8806 372
rect 8840 338 8874 372
rect 8908 355 8947 372
rect 9377 372 9965 388
rect 9377 355 9416 372
rect 8908 338 9133 355
rect 8173 300 9133 338
rect 9191 338 9416 355
rect 9450 338 9484 372
rect 9518 338 9552 372
rect 9586 338 9620 372
rect 9654 338 9688 372
rect 9722 338 9756 372
rect 9790 338 9824 372
rect 9858 338 9892 372
rect 9926 355 9965 372
rect 9926 338 10151 355
rect 9191 300 10151 338
rect -10151 -338 -9191 -300
rect -10151 -355 -9926 -338
rect -9965 -372 -9926 -355
rect -9892 -372 -9858 -338
rect -9824 -372 -9790 -338
rect -9756 -372 -9722 -338
rect -9688 -372 -9654 -338
rect -9620 -372 -9586 -338
rect -9552 -372 -9518 -338
rect -9484 -372 -9450 -338
rect -9416 -355 -9191 -338
rect -9133 -338 -8173 -300
rect -9133 -355 -8908 -338
rect -9416 -372 -9377 -355
rect -9965 -388 -9377 -372
rect -8947 -372 -8908 -355
rect -8874 -372 -8840 -338
rect -8806 -372 -8772 -338
rect -8738 -372 -8704 -338
rect -8670 -372 -8636 -338
rect -8602 -372 -8568 -338
rect -8534 -372 -8500 -338
rect -8466 -372 -8432 -338
rect -8398 -355 -8173 -338
rect -8115 -338 -7155 -300
rect -8115 -355 -7890 -338
rect -8398 -372 -8359 -355
rect -8947 -388 -8359 -372
rect -7929 -372 -7890 -355
rect -7856 -372 -7822 -338
rect -7788 -372 -7754 -338
rect -7720 -372 -7686 -338
rect -7652 -372 -7618 -338
rect -7584 -372 -7550 -338
rect -7516 -372 -7482 -338
rect -7448 -372 -7414 -338
rect -7380 -355 -7155 -338
rect -7097 -338 -6137 -300
rect -7097 -355 -6872 -338
rect -7380 -372 -7341 -355
rect -7929 -388 -7341 -372
rect -6911 -372 -6872 -355
rect -6838 -372 -6804 -338
rect -6770 -372 -6736 -338
rect -6702 -372 -6668 -338
rect -6634 -372 -6600 -338
rect -6566 -372 -6532 -338
rect -6498 -372 -6464 -338
rect -6430 -372 -6396 -338
rect -6362 -355 -6137 -338
rect -6079 -338 -5119 -300
rect -6079 -355 -5854 -338
rect -6362 -372 -6323 -355
rect -6911 -388 -6323 -372
rect -5893 -372 -5854 -355
rect -5820 -372 -5786 -338
rect -5752 -372 -5718 -338
rect -5684 -372 -5650 -338
rect -5616 -372 -5582 -338
rect -5548 -372 -5514 -338
rect -5480 -372 -5446 -338
rect -5412 -372 -5378 -338
rect -5344 -355 -5119 -338
rect -5061 -338 -4101 -300
rect -5061 -355 -4836 -338
rect -5344 -372 -5305 -355
rect -5893 -388 -5305 -372
rect -4875 -372 -4836 -355
rect -4802 -372 -4768 -338
rect -4734 -372 -4700 -338
rect -4666 -372 -4632 -338
rect -4598 -372 -4564 -338
rect -4530 -372 -4496 -338
rect -4462 -372 -4428 -338
rect -4394 -372 -4360 -338
rect -4326 -355 -4101 -338
rect -4043 -338 -3083 -300
rect -4043 -355 -3818 -338
rect -4326 -372 -4287 -355
rect -4875 -388 -4287 -372
rect -3857 -372 -3818 -355
rect -3784 -372 -3750 -338
rect -3716 -372 -3682 -338
rect -3648 -372 -3614 -338
rect -3580 -372 -3546 -338
rect -3512 -372 -3478 -338
rect -3444 -372 -3410 -338
rect -3376 -372 -3342 -338
rect -3308 -355 -3083 -338
rect -3025 -338 -2065 -300
rect -3025 -355 -2800 -338
rect -3308 -372 -3269 -355
rect -3857 -388 -3269 -372
rect -2839 -372 -2800 -355
rect -2766 -372 -2732 -338
rect -2698 -372 -2664 -338
rect -2630 -372 -2596 -338
rect -2562 -372 -2528 -338
rect -2494 -372 -2460 -338
rect -2426 -372 -2392 -338
rect -2358 -372 -2324 -338
rect -2290 -355 -2065 -338
rect -2007 -338 -1047 -300
rect -2007 -355 -1782 -338
rect -2290 -372 -2251 -355
rect -2839 -388 -2251 -372
rect -1821 -372 -1782 -355
rect -1748 -372 -1714 -338
rect -1680 -372 -1646 -338
rect -1612 -372 -1578 -338
rect -1544 -372 -1510 -338
rect -1476 -372 -1442 -338
rect -1408 -372 -1374 -338
rect -1340 -372 -1306 -338
rect -1272 -355 -1047 -338
rect -989 -338 -29 -300
rect -989 -355 -764 -338
rect -1272 -372 -1233 -355
rect -1821 -388 -1233 -372
rect -803 -372 -764 -355
rect -730 -372 -696 -338
rect -662 -372 -628 -338
rect -594 -372 -560 -338
rect -526 -372 -492 -338
rect -458 -372 -424 -338
rect -390 -372 -356 -338
rect -322 -372 -288 -338
rect -254 -355 -29 -338
rect 29 -338 989 -300
rect 29 -355 254 -338
rect -254 -372 -215 -355
rect -803 -388 -215 -372
rect 215 -372 254 -355
rect 288 -372 322 -338
rect 356 -372 390 -338
rect 424 -372 458 -338
rect 492 -372 526 -338
rect 560 -372 594 -338
rect 628 -372 662 -338
rect 696 -372 730 -338
rect 764 -355 989 -338
rect 1047 -338 2007 -300
rect 1047 -355 1272 -338
rect 764 -372 803 -355
rect 215 -388 803 -372
rect 1233 -372 1272 -355
rect 1306 -372 1340 -338
rect 1374 -372 1408 -338
rect 1442 -372 1476 -338
rect 1510 -372 1544 -338
rect 1578 -372 1612 -338
rect 1646 -372 1680 -338
rect 1714 -372 1748 -338
rect 1782 -355 2007 -338
rect 2065 -338 3025 -300
rect 2065 -355 2290 -338
rect 1782 -372 1821 -355
rect 1233 -388 1821 -372
rect 2251 -372 2290 -355
rect 2324 -372 2358 -338
rect 2392 -372 2426 -338
rect 2460 -372 2494 -338
rect 2528 -372 2562 -338
rect 2596 -372 2630 -338
rect 2664 -372 2698 -338
rect 2732 -372 2766 -338
rect 2800 -355 3025 -338
rect 3083 -338 4043 -300
rect 3083 -355 3308 -338
rect 2800 -372 2839 -355
rect 2251 -388 2839 -372
rect 3269 -372 3308 -355
rect 3342 -372 3376 -338
rect 3410 -372 3444 -338
rect 3478 -372 3512 -338
rect 3546 -372 3580 -338
rect 3614 -372 3648 -338
rect 3682 -372 3716 -338
rect 3750 -372 3784 -338
rect 3818 -355 4043 -338
rect 4101 -338 5061 -300
rect 4101 -355 4326 -338
rect 3818 -372 3857 -355
rect 3269 -388 3857 -372
rect 4287 -372 4326 -355
rect 4360 -372 4394 -338
rect 4428 -372 4462 -338
rect 4496 -372 4530 -338
rect 4564 -372 4598 -338
rect 4632 -372 4666 -338
rect 4700 -372 4734 -338
rect 4768 -372 4802 -338
rect 4836 -355 5061 -338
rect 5119 -338 6079 -300
rect 5119 -355 5344 -338
rect 4836 -372 4875 -355
rect 4287 -388 4875 -372
rect 5305 -372 5344 -355
rect 5378 -372 5412 -338
rect 5446 -372 5480 -338
rect 5514 -372 5548 -338
rect 5582 -372 5616 -338
rect 5650 -372 5684 -338
rect 5718 -372 5752 -338
rect 5786 -372 5820 -338
rect 5854 -355 6079 -338
rect 6137 -338 7097 -300
rect 6137 -355 6362 -338
rect 5854 -372 5893 -355
rect 5305 -388 5893 -372
rect 6323 -372 6362 -355
rect 6396 -372 6430 -338
rect 6464 -372 6498 -338
rect 6532 -372 6566 -338
rect 6600 -372 6634 -338
rect 6668 -372 6702 -338
rect 6736 -372 6770 -338
rect 6804 -372 6838 -338
rect 6872 -355 7097 -338
rect 7155 -338 8115 -300
rect 7155 -355 7380 -338
rect 6872 -372 6911 -355
rect 6323 -388 6911 -372
rect 7341 -372 7380 -355
rect 7414 -372 7448 -338
rect 7482 -372 7516 -338
rect 7550 -372 7584 -338
rect 7618 -372 7652 -338
rect 7686 -372 7720 -338
rect 7754 -372 7788 -338
rect 7822 -372 7856 -338
rect 7890 -355 8115 -338
rect 8173 -338 9133 -300
rect 8173 -355 8398 -338
rect 7890 -372 7929 -355
rect 7341 -388 7929 -372
rect 8359 -372 8398 -355
rect 8432 -372 8466 -338
rect 8500 -372 8534 -338
rect 8568 -372 8602 -338
rect 8636 -372 8670 -338
rect 8704 -372 8738 -338
rect 8772 -372 8806 -338
rect 8840 -372 8874 -338
rect 8908 -355 9133 -338
rect 9191 -338 10151 -300
rect 9191 -355 9416 -338
rect 8908 -372 8947 -355
rect 8359 -388 8947 -372
rect 9377 -372 9416 -355
rect 9450 -372 9484 -338
rect 9518 -372 9552 -338
rect 9586 -372 9620 -338
rect 9654 -372 9688 -338
rect 9722 -372 9756 -338
rect 9790 -372 9824 -338
rect 9858 -372 9892 -338
rect 9926 -355 10151 -338
rect 9926 -372 9965 -355
rect 9377 -388 9965 -372
<< polycont >>
rect -9926 338 -9892 372
rect -9858 338 -9824 372
rect -9790 338 -9756 372
rect -9722 338 -9688 372
rect -9654 338 -9620 372
rect -9586 338 -9552 372
rect -9518 338 -9484 372
rect -9450 338 -9416 372
rect -8908 338 -8874 372
rect -8840 338 -8806 372
rect -8772 338 -8738 372
rect -8704 338 -8670 372
rect -8636 338 -8602 372
rect -8568 338 -8534 372
rect -8500 338 -8466 372
rect -8432 338 -8398 372
rect -7890 338 -7856 372
rect -7822 338 -7788 372
rect -7754 338 -7720 372
rect -7686 338 -7652 372
rect -7618 338 -7584 372
rect -7550 338 -7516 372
rect -7482 338 -7448 372
rect -7414 338 -7380 372
rect -6872 338 -6838 372
rect -6804 338 -6770 372
rect -6736 338 -6702 372
rect -6668 338 -6634 372
rect -6600 338 -6566 372
rect -6532 338 -6498 372
rect -6464 338 -6430 372
rect -6396 338 -6362 372
rect -5854 338 -5820 372
rect -5786 338 -5752 372
rect -5718 338 -5684 372
rect -5650 338 -5616 372
rect -5582 338 -5548 372
rect -5514 338 -5480 372
rect -5446 338 -5412 372
rect -5378 338 -5344 372
rect -4836 338 -4802 372
rect -4768 338 -4734 372
rect -4700 338 -4666 372
rect -4632 338 -4598 372
rect -4564 338 -4530 372
rect -4496 338 -4462 372
rect -4428 338 -4394 372
rect -4360 338 -4326 372
rect -3818 338 -3784 372
rect -3750 338 -3716 372
rect -3682 338 -3648 372
rect -3614 338 -3580 372
rect -3546 338 -3512 372
rect -3478 338 -3444 372
rect -3410 338 -3376 372
rect -3342 338 -3308 372
rect -2800 338 -2766 372
rect -2732 338 -2698 372
rect -2664 338 -2630 372
rect -2596 338 -2562 372
rect -2528 338 -2494 372
rect -2460 338 -2426 372
rect -2392 338 -2358 372
rect -2324 338 -2290 372
rect -1782 338 -1748 372
rect -1714 338 -1680 372
rect -1646 338 -1612 372
rect -1578 338 -1544 372
rect -1510 338 -1476 372
rect -1442 338 -1408 372
rect -1374 338 -1340 372
rect -1306 338 -1272 372
rect -764 338 -730 372
rect -696 338 -662 372
rect -628 338 -594 372
rect -560 338 -526 372
rect -492 338 -458 372
rect -424 338 -390 372
rect -356 338 -322 372
rect -288 338 -254 372
rect 254 338 288 372
rect 322 338 356 372
rect 390 338 424 372
rect 458 338 492 372
rect 526 338 560 372
rect 594 338 628 372
rect 662 338 696 372
rect 730 338 764 372
rect 1272 338 1306 372
rect 1340 338 1374 372
rect 1408 338 1442 372
rect 1476 338 1510 372
rect 1544 338 1578 372
rect 1612 338 1646 372
rect 1680 338 1714 372
rect 1748 338 1782 372
rect 2290 338 2324 372
rect 2358 338 2392 372
rect 2426 338 2460 372
rect 2494 338 2528 372
rect 2562 338 2596 372
rect 2630 338 2664 372
rect 2698 338 2732 372
rect 2766 338 2800 372
rect 3308 338 3342 372
rect 3376 338 3410 372
rect 3444 338 3478 372
rect 3512 338 3546 372
rect 3580 338 3614 372
rect 3648 338 3682 372
rect 3716 338 3750 372
rect 3784 338 3818 372
rect 4326 338 4360 372
rect 4394 338 4428 372
rect 4462 338 4496 372
rect 4530 338 4564 372
rect 4598 338 4632 372
rect 4666 338 4700 372
rect 4734 338 4768 372
rect 4802 338 4836 372
rect 5344 338 5378 372
rect 5412 338 5446 372
rect 5480 338 5514 372
rect 5548 338 5582 372
rect 5616 338 5650 372
rect 5684 338 5718 372
rect 5752 338 5786 372
rect 5820 338 5854 372
rect 6362 338 6396 372
rect 6430 338 6464 372
rect 6498 338 6532 372
rect 6566 338 6600 372
rect 6634 338 6668 372
rect 6702 338 6736 372
rect 6770 338 6804 372
rect 6838 338 6872 372
rect 7380 338 7414 372
rect 7448 338 7482 372
rect 7516 338 7550 372
rect 7584 338 7618 372
rect 7652 338 7686 372
rect 7720 338 7754 372
rect 7788 338 7822 372
rect 7856 338 7890 372
rect 8398 338 8432 372
rect 8466 338 8500 372
rect 8534 338 8568 372
rect 8602 338 8636 372
rect 8670 338 8704 372
rect 8738 338 8772 372
rect 8806 338 8840 372
rect 8874 338 8908 372
rect 9416 338 9450 372
rect 9484 338 9518 372
rect 9552 338 9586 372
rect 9620 338 9654 372
rect 9688 338 9722 372
rect 9756 338 9790 372
rect 9824 338 9858 372
rect 9892 338 9926 372
rect -9926 -372 -9892 -338
rect -9858 -372 -9824 -338
rect -9790 -372 -9756 -338
rect -9722 -372 -9688 -338
rect -9654 -372 -9620 -338
rect -9586 -372 -9552 -338
rect -9518 -372 -9484 -338
rect -9450 -372 -9416 -338
rect -8908 -372 -8874 -338
rect -8840 -372 -8806 -338
rect -8772 -372 -8738 -338
rect -8704 -372 -8670 -338
rect -8636 -372 -8602 -338
rect -8568 -372 -8534 -338
rect -8500 -372 -8466 -338
rect -8432 -372 -8398 -338
rect -7890 -372 -7856 -338
rect -7822 -372 -7788 -338
rect -7754 -372 -7720 -338
rect -7686 -372 -7652 -338
rect -7618 -372 -7584 -338
rect -7550 -372 -7516 -338
rect -7482 -372 -7448 -338
rect -7414 -372 -7380 -338
rect -6872 -372 -6838 -338
rect -6804 -372 -6770 -338
rect -6736 -372 -6702 -338
rect -6668 -372 -6634 -338
rect -6600 -372 -6566 -338
rect -6532 -372 -6498 -338
rect -6464 -372 -6430 -338
rect -6396 -372 -6362 -338
rect -5854 -372 -5820 -338
rect -5786 -372 -5752 -338
rect -5718 -372 -5684 -338
rect -5650 -372 -5616 -338
rect -5582 -372 -5548 -338
rect -5514 -372 -5480 -338
rect -5446 -372 -5412 -338
rect -5378 -372 -5344 -338
rect -4836 -372 -4802 -338
rect -4768 -372 -4734 -338
rect -4700 -372 -4666 -338
rect -4632 -372 -4598 -338
rect -4564 -372 -4530 -338
rect -4496 -372 -4462 -338
rect -4428 -372 -4394 -338
rect -4360 -372 -4326 -338
rect -3818 -372 -3784 -338
rect -3750 -372 -3716 -338
rect -3682 -372 -3648 -338
rect -3614 -372 -3580 -338
rect -3546 -372 -3512 -338
rect -3478 -372 -3444 -338
rect -3410 -372 -3376 -338
rect -3342 -372 -3308 -338
rect -2800 -372 -2766 -338
rect -2732 -372 -2698 -338
rect -2664 -372 -2630 -338
rect -2596 -372 -2562 -338
rect -2528 -372 -2494 -338
rect -2460 -372 -2426 -338
rect -2392 -372 -2358 -338
rect -2324 -372 -2290 -338
rect -1782 -372 -1748 -338
rect -1714 -372 -1680 -338
rect -1646 -372 -1612 -338
rect -1578 -372 -1544 -338
rect -1510 -372 -1476 -338
rect -1442 -372 -1408 -338
rect -1374 -372 -1340 -338
rect -1306 -372 -1272 -338
rect -764 -372 -730 -338
rect -696 -372 -662 -338
rect -628 -372 -594 -338
rect -560 -372 -526 -338
rect -492 -372 -458 -338
rect -424 -372 -390 -338
rect -356 -372 -322 -338
rect -288 -372 -254 -338
rect 254 -372 288 -338
rect 322 -372 356 -338
rect 390 -372 424 -338
rect 458 -372 492 -338
rect 526 -372 560 -338
rect 594 -372 628 -338
rect 662 -372 696 -338
rect 730 -372 764 -338
rect 1272 -372 1306 -338
rect 1340 -372 1374 -338
rect 1408 -372 1442 -338
rect 1476 -372 1510 -338
rect 1544 -372 1578 -338
rect 1612 -372 1646 -338
rect 1680 -372 1714 -338
rect 1748 -372 1782 -338
rect 2290 -372 2324 -338
rect 2358 -372 2392 -338
rect 2426 -372 2460 -338
rect 2494 -372 2528 -338
rect 2562 -372 2596 -338
rect 2630 -372 2664 -338
rect 2698 -372 2732 -338
rect 2766 -372 2800 -338
rect 3308 -372 3342 -338
rect 3376 -372 3410 -338
rect 3444 -372 3478 -338
rect 3512 -372 3546 -338
rect 3580 -372 3614 -338
rect 3648 -372 3682 -338
rect 3716 -372 3750 -338
rect 3784 -372 3818 -338
rect 4326 -372 4360 -338
rect 4394 -372 4428 -338
rect 4462 -372 4496 -338
rect 4530 -372 4564 -338
rect 4598 -372 4632 -338
rect 4666 -372 4700 -338
rect 4734 -372 4768 -338
rect 4802 -372 4836 -338
rect 5344 -372 5378 -338
rect 5412 -372 5446 -338
rect 5480 -372 5514 -338
rect 5548 -372 5582 -338
rect 5616 -372 5650 -338
rect 5684 -372 5718 -338
rect 5752 -372 5786 -338
rect 5820 -372 5854 -338
rect 6362 -372 6396 -338
rect 6430 -372 6464 -338
rect 6498 -372 6532 -338
rect 6566 -372 6600 -338
rect 6634 -372 6668 -338
rect 6702 -372 6736 -338
rect 6770 -372 6804 -338
rect 6838 -372 6872 -338
rect 7380 -372 7414 -338
rect 7448 -372 7482 -338
rect 7516 -372 7550 -338
rect 7584 -372 7618 -338
rect 7652 -372 7686 -338
rect 7720 -372 7754 -338
rect 7788 -372 7822 -338
rect 7856 -372 7890 -338
rect 8398 -372 8432 -338
rect 8466 -372 8500 -338
rect 8534 -372 8568 -338
rect 8602 -372 8636 -338
rect 8670 -372 8704 -338
rect 8738 -372 8772 -338
rect 8806 -372 8840 -338
rect 8874 -372 8908 -338
rect 9416 -372 9450 -338
rect 9484 -372 9518 -338
rect 9552 -372 9586 -338
rect 9620 -372 9654 -338
rect 9688 -372 9722 -338
rect 9756 -372 9790 -338
rect 9824 -372 9858 -338
rect 9892 -372 9926 -338
<< locali >>
rect -9965 338 -9926 372
rect -9892 338 -9868 372
rect -9824 338 -9796 372
rect -9756 338 -9724 372
rect -9688 338 -9654 372
rect -9618 338 -9586 372
rect -9546 338 -9518 372
rect -9474 338 -9450 372
rect -9416 338 -9377 372
rect -8947 338 -8908 372
rect -8874 338 -8850 372
rect -8806 338 -8778 372
rect -8738 338 -8706 372
rect -8670 338 -8636 372
rect -8600 338 -8568 372
rect -8528 338 -8500 372
rect -8456 338 -8432 372
rect -8398 338 -8359 372
rect -7929 338 -7890 372
rect -7856 338 -7832 372
rect -7788 338 -7760 372
rect -7720 338 -7688 372
rect -7652 338 -7618 372
rect -7582 338 -7550 372
rect -7510 338 -7482 372
rect -7438 338 -7414 372
rect -7380 338 -7341 372
rect -6911 338 -6872 372
rect -6838 338 -6814 372
rect -6770 338 -6742 372
rect -6702 338 -6670 372
rect -6634 338 -6600 372
rect -6564 338 -6532 372
rect -6492 338 -6464 372
rect -6420 338 -6396 372
rect -6362 338 -6323 372
rect -5893 338 -5854 372
rect -5820 338 -5796 372
rect -5752 338 -5724 372
rect -5684 338 -5652 372
rect -5616 338 -5582 372
rect -5546 338 -5514 372
rect -5474 338 -5446 372
rect -5402 338 -5378 372
rect -5344 338 -5305 372
rect -4875 338 -4836 372
rect -4802 338 -4778 372
rect -4734 338 -4706 372
rect -4666 338 -4634 372
rect -4598 338 -4564 372
rect -4528 338 -4496 372
rect -4456 338 -4428 372
rect -4384 338 -4360 372
rect -4326 338 -4287 372
rect -3857 338 -3818 372
rect -3784 338 -3760 372
rect -3716 338 -3688 372
rect -3648 338 -3616 372
rect -3580 338 -3546 372
rect -3510 338 -3478 372
rect -3438 338 -3410 372
rect -3366 338 -3342 372
rect -3308 338 -3269 372
rect -2839 338 -2800 372
rect -2766 338 -2742 372
rect -2698 338 -2670 372
rect -2630 338 -2598 372
rect -2562 338 -2528 372
rect -2492 338 -2460 372
rect -2420 338 -2392 372
rect -2348 338 -2324 372
rect -2290 338 -2251 372
rect -1821 338 -1782 372
rect -1748 338 -1724 372
rect -1680 338 -1652 372
rect -1612 338 -1580 372
rect -1544 338 -1510 372
rect -1474 338 -1442 372
rect -1402 338 -1374 372
rect -1330 338 -1306 372
rect -1272 338 -1233 372
rect -803 338 -764 372
rect -730 338 -706 372
rect -662 338 -634 372
rect -594 338 -562 372
rect -526 338 -492 372
rect -456 338 -424 372
rect -384 338 -356 372
rect -312 338 -288 372
rect -254 338 -215 372
rect 215 338 254 372
rect 288 338 312 372
rect 356 338 384 372
rect 424 338 456 372
rect 492 338 526 372
rect 562 338 594 372
rect 634 338 662 372
rect 706 338 730 372
rect 764 338 803 372
rect 1233 338 1272 372
rect 1306 338 1330 372
rect 1374 338 1402 372
rect 1442 338 1474 372
rect 1510 338 1544 372
rect 1580 338 1612 372
rect 1652 338 1680 372
rect 1724 338 1748 372
rect 1782 338 1821 372
rect 2251 338 2290 372
rect 2324 338 2348 372
rect 2392 338 2420 372
rect 2460 338 2492 372
rect 2528 338 2562 372
rect 2598 338 2630 372
rect 2670 338 2698 372
rect 2742 338 2766 372
rect 2800 338 2839 372
rect 3269 338 3308 372
rect 3342 338 3366 372
rect 3410 338 3438 372
rect 3478 338 3510 372
rect 3546 338 3580 372
rect 3616 338 3648 372
rect 3688 338 3716 372
rect 3760 338 3784 372
rect 3818 338 3857 372
rect 4287 338 4326 372
rect 4360 338 4384 372
rect 4428 338 4456 372
rect 4496 338 4528 372
rect 4564 338 4598 372
rect 4634 338 4666 372
rect 4706 338 4734 372
rect 4778 338 4802 372
rect 4836 338 4875 372
rect 5305 338 5344 372
rect 5378 338 5402 372
rect 5446 338 5474 372
rect 5514 338 5546 372
rect 5582 338 5616 372
rect 5652 338 5684 372
rect 5724 338 5752 372
rect 5796 338 5820 372
rect 5854 338 5893 372
rect 6323 338 6362 372
rect 6396 338 6420 372
rect 6464 338 6492 372
rect 6532 338 6564 372
rect 6600 338 6634 372
rect 6670 338 6702 372
rect 6742 338 6770 372
rect 6814 338 6838 372
rect 6872 338 6911 372
rect 7341 338 7380 372
rect 7414 338 7438 372
rect 7482 338 7510 372
rect 7550 338 7582 372
rect 7618 338 7652 372
rect 7688 338 7720 372
rect 7760 338 7788 372
rect 7832 338 7856 372
rect 7890 338 7929 372
rect 8359 338 8398 372
rect 8432 338 8456 372
rect 8500 338 8528 372
rect 8568 338 8600 372
rect 8636 338 8670 372
rect 8706 338 8738 372
rect 8778 338 8806 372
rect 8850 338 8874 372
rect 8908 338 8947 372
rect 9377 338 9416 372
rect 9450 338 9474 372
rect 9518 338 9546 372
rect 9586 338 9618 372
rect 9654 338 9688 372
rect 9724 338 9756 372
rect 9796 338 9824 372
rect 9868 338 9892 372
rect 9926 338 9965 372
rect -10197 269 -10163 304
rect -10197 197 -10163 221
rect -10197 125 -10163 153
rect -10197 53 -10163 85
rect -10197 -17 -10163 17
rect -10197 -85 -10163 -53
rect -10197 -153 -10163 -125
rect -10197 -221 -10163 -197
rect -10197 -304 -10163 -269
rect -9179 269 -9145 304
rect -9179 197 -9145 221
rect -9179 125 -9145 153
rect -9179 53 -9145 85
rect -9179 -17 -9145 17
rect -9179 -85 -9145 -53
rect -9179 -153 -9145 -125
rect -9179 -221 -9145 -197
rect -9179 -304 -9145 -269
rect -8161 269 -8127 304
rect -8161 197 -8127 221
rect -8161 125 -8127 153
rect -8161 53 -8127 85
rect -8161 -17 -8127 17
rect -8161 -85 -8127 -53
rect -8161 -153 -8127 -125
rect -8161 -221 -8127 -197
rect -8161 -304 -8127 -269
rect -7143 269 -7109 304
rect -7143 197 -7109 221
rect -7143 125 -7109 153
rect -7143 53 -7109 85
rect -7143 -17 -7109 17
rect -7143 -85 -7109 -53
rect -7143 -153 -7109 -125
rect -7143 -221 -7109 -197
rect -7143 -304 -7109 -269
rect -6125 269 -6091 304
rect -6125 197 -6091 221
rect -6125 125 -6091 153
rect -6125 53 -6091 85
rect -6125 -17 -6091 17
rect -6125 -85 -6091 -53
rect -6125 -153 -6091 -125
rect -6125 -221 -6091 -197
rect -6125 -304 -6091 -269
rect -5107 269 -5073 304
rect -5107 197 -5073 221
rect -5107 125 -5073 153
rect -5107 53 -5073 85
rect -5107 -17 -5073 17
rect -5107 -85 -5073 -53
rect -5107 -153 -5073 -125
rect -5107 -221 -5073 -197
rect -5107 -304 -5073 -269
rect -4089 269 -4055 304
rect -4089 197 -4055 221
rect -4089 125 -4055 153
rect -4089 53 -4055 85
rect -4089 -17 -4055 17
rect -4089 -85 -4055 -53
rect -4089 -153 -4055 -125
rect -4089 -221 -4055 -197
rect -4089 -304 -4055 -269
rect -3071 269 -3037 304
rect -3071 197 -3037 221
rect -3071 125 -3037 153
rect -3071 53 -3037 85
rect -3071 -17 -3037 17
rect -3071 -85 -3037 -53
rect -3071 -153 -3037 -125
rect -3071 -221 -3037 -197
rect -3071 -304 -3037 -269
rect -2053 269 -2019 304
rect -2053 197 -2019 221
rect -2053 125 -2019 153
rect -2053 53 -2019 85
rect -2053 -17 -2019 17
rect -2053 -85 -2019 -53
rect -2053 -153 -2019 -125
rect -2053 -221 -2019 -197
rect -2053 -304 -2019 -269
rect -1035 269 -1001 304
rect -1035 197 -1001 221
rect -1035 125 -1001 153
rect -1035 53 -1001 85
rect -1035 -17 -1001 17
rect -1035 -85 -1001 -53
rect -1035 -153 -1001 -125
rect -1035 -221 -1001 -197
rect -1035 -304 -1001 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 1001 269 1035 304
rect 1001 197 1035 221
rect 1001 125 1035 153
rect 1001 53 1035 85
rect 1001 -17 1035 17
rect 1001 -85 1035 -53
rect 1001 -153 1035 -125
rect 1001 -221 1035 -197
rect 1001 -304 1035 -269
rect 2019 269 2053 304
rect 2019 197 2053 221
rect 2019 125 2053 153
rect 2019 53 2053 85
rect 2019 -17 2053 17
rect 2019 -85 2053 -53
rect 2019 -153 2053 -125
rect 2019 -221 2053 -197
rect 2019 -304 2053 -269
rect 3037 269 3071 304
rect 3037 197 3071 221
rect 3037 125 3071 153
rect 3037 53 3071 85
rect 3037 -17 3071 17
rect 3037 -85 3071 -53
rect 3037 -153 3071 -125
rect 3037 -221 3071 -197
rect 3037 -304 3071 -269
rect 4055 269 4089 304
rect 4055 197 4089 221
rect 4055 125 4089 153
rect 4055 53 4089 85
rect 4055 -17 4089 17
rect 4055 -85 4089 -53
rect 4055 -153 4089 -125
rect 4055 -221 4089 -197
rect 4055 -304 4089 -269
rect 5073 269 5107 304
rect 5073 197 5107 221
rect 5073 125 5107 153
rect 5073 53 5107 85
rect 5073 -17 5107 17
rect 5073 -85 5107 -53
rect 5073 -153 5107 -125
rect 5073 -221 5107 -197
rect 5073 -304 5107 -269
rect 6091 269 6125 304
rect 6091 197 6125 221
rect 6091 125 6125 153
rect 6091 53 6125 85
rect 6091 -17 6125 17
rect 6091 -85 6125 -53
rect 6091 -153 6125 -125
rect 6091 -221 6125 -197
rect 6091 -304 6125 -269
rect 7109 269 7143 304
rect 7109 197 7143 221
rect 7109 125 7143 153
rect 7109 53 7143 85
rect 7109 -17 7143 17
rect 7109 -85 7143 -53
rect 7109 -153 7143 -125
rect 7109 -221 7143 -197
rect 7109 -304 7143 -269
rect 8127 269 8161 304
rect 8127 197 8161 221
rect 8127 125 8161 153
rect 8127 53 8161 85
rect 8127 -17 8161 17
rect 8127 -85 8161 -53
rect 8127 -153 8161 -125
rect 8127 -221 8161 -197
rect 8127 -304 8161 -269
rect 9145 269 9179 304
rect 9145 197 9179 221
rect 9145 125 9179 153
rect 9145 53 9179 85
rect 9145 -17 9179 17
rect 9145 -85 9179 -53
rect 9145 -153 9179 -125
rect 9145 -221 9179 -197
rect 9145 -304 9179 -269
rect 10163 269 10197 304
rect 10163 197 10197 221
rect 10163 125 10197 153
rect 10163 53 10197 85
rect 10163 -17 10197 17
rect 10163 -85 10197 -53
rect 10163 -153 10197 -125
rect 10163 -221 10197 -197
rect 10163 -304 10197 -269
rect -9965 -372 -9926 -338
rect -9892 -372 -9868 -338
rect -9824 -372 -9796 -338
rect -9756 -372 -9724 -338
rect -9688 -372 -9654 -338
rect -9618 -372 -9586 -338
rect -9546 -372 -9518 -338
rect -9474 -372 -9450 -338
rect -9416 -372 -9377 -338
rect -8947 -372 -8908 -338
rect -8874 -372 -8850 -338
rect -8806 -372 -8778 -338
rect -8738 -372 -8706 -338
rect -8670 -372 -8636 -338
rect -8600 -372 -8568 -338
rect -8528 -372 -8500 -338
rect -8456 -372 -8432 -338
rect -8398 -372 -8359 -338
rect -7929 -372 -7890 -338
rect -7856 -372 -7832 -338
rect -7788 -372 -7760 -338
rect -7720 -372 -7688 -338
rect -7652 -372 -7618 -338
rect -7582 -372 -7550 -338
rect -7510 -372 -7482 -338
rect -7438 -372 -7414 -338
rect -7380 -372 -7341 -338
rect -6911 -372 -6872 -338
rect -6838 -372 -6814 -338
rect -6770 -372 -6742 -338
rect -6702 -372 -6670 -338
rect -6634 -372 -6600 -338
rect -6564 -372 -6532 -338
rect -6492 -372 -6464 -338
rect -6420 -372 -6396 -338
rect -6362 -372 -6323 -338
rect -5893 -372 -5854 -338
rect -5820 -372 -5796 -338
rect -5752 -372 -5724 -338
rect -5684 -372 -5652 -338
rect -5616 -372 -5582 -338
rect -5546 -372 -5514 -338
rect -5474 -372 -5446 -338
rect -5402 -372 -5378 -338
rect -5344 -372 -5305 -338
rect -4875 -372 -4836 -338
rect -4802 -372 -4778 -338
rect -4734 -372 -4706 -338
rect -4666 -372 -4634 -338
rect -4598 -372 -4564 -338
rect -4528 -372 -4496 -338
rect -4456 -372 -4428 -338
rect -4384 -372 -4360 -338
rect -4326 -372 -4287 -338
rect -3857 -372 -3818 -338
rect -3784 -372 -3760 -338
rect -3716 -372 -3688 -338
rect -3648 -372 -3616 -338
rect -3580 -372 -3546 -338
rect -3510 -372 -3478 -338
rect -3438 -372 -3410 -338
rect -3366 -372 -3342 -338
rect -3308 -372 -3269 -338
rect -2839 -372 -2800 -338
rect -2766 -372 -2742 -338
rect -2698 -372 -2670 -338
rect -2630 -372 -2598 -338
rect -2562 -372 -2528 -338
rect -2492 -372 -2460 -338
rect -2420 -372 -2392 -338
rect -2348 -372 -2324 -338
rect -2290 -372 -2251 -338
rect -1821 -372 -1782 -338
rect -1748 -372 -1724 -338
rect -1680 -372 -1652 -338
rect -1612 -372 -1580 -338
rect -1544 -372 -1510 -338
rect -1474 -372 -1442 -338
rect -1402 -372 -1374 -338
rect -1330 -372 -1306 -338
rect -1272 -372 -1233 -338
rect -803 -372 -764 -338
rect -730 -372 -706 -338
rect -662 -372 -634 -338
rect -594 -372 -562 -338
rect -526 -372 -492 -338
rect -456 -372 -424 -338
rect -384 -372 -356 -338
rect -312 -372 -288 -338
rect -254 -372 -215 -338
rect 215 -372 254 -338
rect 288 -372 312 -338
rect 356 -372 384 -338
rect 424 -372 456 -338
rect 492 -372 526 -338
rect 562 -372 594 -338
rect 634 -372 662 -338
rect 706 -372 730 -338
rect 764 -372 803 -338
rect 1233 -372 1272 -338
rect 1306 -372 1330 -338
rect 1374 -372 1402 -338
rect 1442 -372 1474 -338
rect 1510 -372 1544 -338
rect 1580 -372 1612 -338
rect 1652 -372 1680 -338
rect 1724 -372 1748 -338
rect 1782 -372 1821 -338
rect 2251 -372 2290 -338
rect 2324 -372 2348 -338
rect 2392 -372 2420 -338
rect 2460 -372 2492 -338
rect 2528 -372 2562 -338
rect 2598 -372 2630 -338
rect 2670 -372 2698 -338
rect 2742 -372 2766 -338
rect 2800 -372 2839 -338
rect 3269 -372 3308 -338
rect 3342 -372 3366 -338
rect 3410 -372 3438 -338
rect 3478 -372 3510 -338
rect 3546 -372 3580 -338
rect 3616 -372 3648 -338
rect 3688 -372 3716 -338
rect 3760 -372 3784 -338
rect 3818 -372 3857 -338
rect 4287 -372 4326 -338
rect 4360 -372 4384 -338
rect 4428 -372 4456 -338
rect 4496 -372 4528 -338
rect 4564 -372 4598 -338
rect 4634 -372 4666 -338
rect 4706 -372 4734 -338
rect 4778 -372 4802 -338
rect 4836 -372 4875 -338
rect 5305 -372 5344 -338
rect 5378 -372 5402 -338
rect 5446 -372 5474 -338
rect 5514 -372 5546 -338
rect 5582 -372 5616 -338
rect 5652 -372 5684 -338
rect 5724 -372 5752 -338
rect 5796 -372 5820 -338
rect 5854 -372 5893 -338
rect 6323 -372 6362 -338
rect 6396 -372 6420 -338
rect 6464 -372 6492 -338
rect 6532 -372 6564 -338
rect 6600 -372 6634 -338
rect 6670 -372 6702 -338
rect 6742 -372 6770 -338
rect 6814 -372 6838 -338
rect 6872 -372 6911 -338
rect 7341 -372 7380 -338
rect 7414 -372 7438 -338
rect 7482 -372 7510 -338
rect 7550 -372 7582 -338
rect 7618 -372 7652 -338
rect 7688 -372 7720 -338
rect 7760 -372 7788 -338
rect 7832 -372 7856 -338
rect 7890 -372 7929 -338
rect 8359 -372 8398 -338
rect 8432 -372 8456 -338
rect 8500 -372 8528 -338
rect 8568 -372 8600 -338
rect 8636 -372 8670 -338
rect 8706 -372 8738 -338
rect 8778 -372 8806 -338
rect 8850 -372 8874 -338
rect 8908 -372 8947 -338
rect 9377 -372 9416 -338
rect 9450 -372 9474 -338
rect 9518 -372 9546 -338
rect 9586 -372 9618 -338
rect 9654 -372 9688 -338
rect 9724 -372 9756 -338
rect 9796 -372 9824 -338
rect 9868 -372 9892 -338
rect 9926 -372 9965 -338
<< viali >>
rect -9868 338 -9858 372
rect -9858 338 -9834 372
rect -9796 338 -9790 372
rect -9790 338 -9762 372
rect -9724 338 -9722 372
rect -9722 338 -9690 372
rect -9652 338 -9620 372
rect -9620 338 -9618 372
rect -9580 338 -9552 372
rect -9552 338 -9546 372
rect -9508 338 -9484 372
rect -9484 338 -9474 372
rect -8850 338 -8840 372
rect -8840 338 -8816 372
rect -8778 338 -8772 372
rect -8772 338 -8744 372
rect -8706 338 -8704 372
rect -8704 338 -8672 372
rect -8634 338 -8602 372
rect -8602 338 -8600 372
rect -8562 338 -8534 372
rect -8534 338 -8528 372
rect -8490 338 -8466 372
rect -8466 338 -8456 372
rect -7832 338 -7822 372
rect -7822 338 -7798 372
rect -7760 338 -7754 372
rect -7754 338 -7726 372
rect -7688 338 -7686 372
rect -7686 338 -7654 372
rect -7616 338 -7584 372
rect -7584 338 -7582 372
rect -7544 338 -7516 372
rect -7516 338 -7510 372
rect -7472 338 -7448 372
rect -7448 338 -7438 372
rect -6814 338 -6804 372
rect -6804 338 -6780 372
rect -6742 338 -6736 372
rect -6736 338 -6708 372
rect -6670 338 -6668 372
rect -6668 338 -6636 372
rect -6598 338 -6566 372
rect -6566 338 -6564 372
rect -6526 338 -6498 372
rect -6498 338 -6492 372
rect -6454 338 -6430 372
rect -6430 338 -6420 372
rect -5796 338 -5786 372
rect -5786 338 -5762 372
rect -5724 338 -5718 372
rect -5718 338 -5690 372
rect -5652 338 -5650 372
rect -5650 338 -5618 372
rect -5580 338 -5548 372
rect -5548 338 -5546 372
rect -5508 338 -5480 372
rect -5480 338 -5474 372
rect -5436 338 -5412 372
rect -5412 338 -5402 372
rect -4778 338 -4768 372
rect -4768 338 -4744 372
rect -4706 338 -4700 372
rect -4700 338 -4672 372
rect -4634 338 -4632 372
rect -4632 338 -4600 372
rect -4562 338 -4530 372
rect -4530 338 -4528 372
rect -4490 338 -4462 372
rect -4462 338 -4456 372
rect -4418 338 -4394 372
rect -4394 338 -4384 372
rect -3760 338 -3750 372
rect -3750 338 -3726 372
rect -3688 338 -3682 372
rect -3682 338 -3654 372
rect -3616 338 -3614 372
rect -3614 338 -3582 372
rect -3544 338 -3512 372
rect -3512 338 -3510 372
rect -3472 338 -3444 372
rect -3444 338 -3438 372
rect -3400 338 -3376 372
rect -3376 338 -3366 372
rect -2742 338 -2732 372
rect -2732 338 -2708 372
rect -2670 338 -2664 372
rect -2664 338 -2636 372
rect -2598 338 -2596 372
rect -2596 338 -2564 372
rect -2526 338 -2494 372
rect -2494 338 -2492 372
rect -2454 338 -2426 372
rect -2426 338 -2420 372
rect -2382 338 -2358 372
rect -2358 338 -2348 372
rect -1724 338 -1714 372
rect -1714 338 -1690 372
rect -1652 338 -1646 372
rect -1646 338 -1618 372
rect -1580 338 -1578 372
rect -1578 338 -1546 372
rect -1508 338 -1476 372
rect -1476 338 -1474 372
rect -1436 338 -1408 372
rect -1408 338 -1402 372
rect -1364 338 -1340 372
rect -1340 338 -1330 372
rect -706 338 -696 372
rect -696 338 -672 372
rect -634 338 -628 372
rect -628 338 -600 372
rect -562 338 -560 372
rect -560 338 -528 372
rect -490 338 -458 372
rect -458 338 -456 372
rect -418 338 -390 372
rect -390 338 -384 372
rect -346 338 -322 372
rect -322 338 -312 372
rect 312 338 322 372
rect 322 338 346 372
rect 384 338 390 372
rect 390 338 418 372
rect 456 338 458 372
rect 458 338 490 372
rect 528 338 560 372
rect 560 338 562 372
rect 600 338 628 372
rect 628 338 634 372
rect 672 338 696 372
rect 696 338 706 372
rect 1330 338 1340 372
rect 1340 338 1364 372
rect 1402 338 1408 372
rect 1408 338 1436 372
rect 1474 338 1476 372
rect 1476 338 1508 372
rect 1546 338 1578 372
rect 1578 338 1580 372
rect 1618 338 1646 372
rect 1646 338 1652 372
rect 1690 338 1714 372
rect 1714 338 1724 372
rect 2348 338 2358 372
rect 2358 338 2382 372
rect 2420 338 2426 372
rect 2426 338 2454 372
rect 2492 338 2494 372
rect 2494 338 2526 372
rect 2564 338 2596 372
rect 2596 338 2598 372
rect 2636 338 2664 372
rect 2664 338 2670 372
rect 2708 338 2732 372
rect 2732 338 2742 372
rect 3366 338 3376 372
rect 3376 338 3400 372
rect 3438 338 3444 372
rect 3444 338 3472 372
rect 3510 338 3512 372
rect 3512 338 3544 372
rect 3582 338 3614 372
rect 3614 338 3616 372
rect 3654 338 3682 372
rect 3682 338 3688 372
rect 3726 338 3750 372
rect 3750 338 3760 372
rect 4384 338 4394 372
rect 4394 338 4418 372
rect 4456 338 4462 372
rect 4462 338 4490 372
rect 4528 338 4530 372
rect 4530 338 4562 372
rect 4600 338 4632 372
rect 4632 338 4634 372
rect 4672 338 4700 372
rect 4700 338 4706 372
rect 4744 338 4768 372
rect 4768 338 4778 372
rect 5402 338 5412 372
rect 5412 338 5436 372
rect 5474 338 5480 372
rect 5480 338 5508 372
rect 5546 338 5548 372
rect 5548 338 5580 372
rect 5618 338 5650 372
rect 5650 338 5652 372
rect 5690 338 5718 372
rect 5718 338 5724 372
rect 5762 338 5786 372
rect 5786 338 5796 372
rect 6420 338 6430 372
rect 6430 338 6454 372
rect 6492 338 6498 372
rect 6498 338 6526 372
rect 6564 338 6566 372
rect 6566 338 6598 372
rect 6636 338 6668 372
rect 6668 338 6670 372
rect 6708 338 6736 372
rect 6736 338 6742 372
rect 6780 338 6804 372
rect 6804 338 6814 372
rect 7438 338 7448 372
rect 7448 338 7472 372
rect 7510 338 7516 372
rect 7516 338 7544 372
rect 7582 338 7584 372
rect 7584 338 7616 372
rect 7654 338 7686 372
rect 7686 338 7688 372
rect 7726 338 7754 372
rect 7754 338 7760 372
rect 7798 338 7822 372
rect 7822 338 7832 372
rect 8456 338 8466 372
rect 8466 338 8490 372
rect 8528 338 8534 372
rect 8534 338 8562 372
rect 8600 338 8602 372
rect 8602 338 8634 372
rect 8672 338 8704 372
rect 8704 338 8706 372
rect 8744 338 8772 372
rect 8772 338 8778 372
rect 8816 338 8840 372
rect 8840 338 8850 372
rect 9474 338 9484 372
rect 9484 338 9508 372
rect 9546 338 9552 372
rect 9552 338 9580 372
rect 9618 338 9620 372
rect 9620 338 9652 372
rect 9690 338 9722 372
rect 9722 338 9724 372
rect 9762 338 9790 372
rect 9790 338 9796 372
rect 9834 338 9858 372
rect 9858 338 9868 372
rect -10197 255 -10163 269
rect -10197 235 -10163 255
rect -10197 187 -10163 197
rect -10197 163 -10163 187
rect -10197 119 -10163 125
rect -10197 91 -10163 119
rect -10197 51 -10163 53
rect -10197 19 -10163 51
rect -10197 -51 -10163 -19
rect -10197 -53 -10163 -51
rect -10197 -119 -10163 -91
rect -10197 -125 -10163 -119
rect -10197 -187 -10163 -163
rect -10197 -197 -10163 -187
rect -10197 -255 -10163 -235
rect -10197 -269 -10163 -255
rect -9179 255 -9145 269
rect -9179 235 -9145 255
rect -9179 187 -9145 197
rect -9179 163 -9145 187
rect -9179 119 -9145 125
rect -9179 91 -9145 119
rect -9179 51 -9145 53
rect -9179 19 -9145 51
rect -9179 -51 -9145 -19
rect -9179 -53 -9145 -51
rect -9179 -119 -9145 -91
rect -9179 -125 -9145 -119
rect -9179 -187 -9145 -163
rect -9179 -197 -9145 -187
rect -9179 -255 -9145 -235
rect -9179 -269 -9145 -255
rect -8161 255 -8127 269
rect -8161 235 -8127 255
rect -8161 187 -8127 197
rect -8161 163 -8127 187
rect -8161 119 -8127 125
rect -8161 91 -8127 119
rect -8161 51 -8127 53
rect -8161 19 -8127 51
rect -8161 -51 -8127 -19
rect -8161 -53 -8127 -51
rect -8161 -119 -8127 -91
rect -8161 -125 -8127 -119
rect -8161 -187 -8127 -163
rect -8161 -197 -8127 -187
rect -8161 -255 -8127 -235
rect -8161 -269 -8127 -255
rect -7143 255 -7109 269
rect -7143 235 -7109 255
rect -7143 187 -7109 197
rect -7143 163 -7109 187
rect -7143 119 -7109 125
rect -7143 91 -7109 119
rect -7143 51 -7109 53
rect -7143 19 -7109 51
rect -7143 -51 -7109 -19
rect -7143 -53 -7109 -51
rect -7143 -119 -7109 -91
rect -7143 -125 -7109 -119
rect -7143 -187 -7109 -163
rect -7143 -197 -7109 -187
rect -7143 -255 -7109 -235
rect -7143 -269 -7109 -255
rect -6125 255 -6091 269
rect -6125 235 -6091 255
rect -6125 187 -6091 197
rect -6125 163 -6091 187
rect -6125 119 -6091 125
rect -6125 91 -6091 119
rect -6125 51 -6091 53
rect -6125 19 -6091 51
rect -6125 -51 -6091 -19
rect -6125 -53 -6091 -51
rect -6125 -119 -6091 -91
rect -6125 -125 -6091 -119
rect -6125 -187 -6091 -163
rect -6125 -197 -6091 -187
rect -6125 -255 -6091 -235
rect -6125 -269 -6091 -255
rect -5107 255 -5073 269
rect -5107 235 -5073 255
rect -5107 187 -5073 197
rect -5107 163 -5073 187
rect -5107 119 -5073 125
rect -5107 91 -5073 119
rect -5107 51 -5073 53
rect -5107 19 -5073 51
rect -5107 -51 -5073 -19
rect -5107 -53 -5073 -51
rect -5107 -119 -5073 -91
rect -5107 -125 -5073 -119
rect -5107 -187 -5073 -163
rect -5107 -197 -5073 -187
rect -5107 -255 -5073 -235
rect -5107 -269 -5073 -255
rect -4089 255 -4055 269
rect -4089 235 -4055 255
rect -4089 187 -4055 197
rect -4089 163 -4055 187
rect -4089 119 -4055 125
rect -4089 91 -4055 119
rect -4089 51 -4055 53
rect -4089 19 -4055 51
rect -4089 -51 -4055 -19
rect -4089 -53 -4055 -51
rect -4089 -119 -4055 -91
rect -4089 -125 -4055 -119
rect -4089 -187 -4055 -163
rect -4089 -197 -4055 -187
rect -4089 -255 -4055 -235
rect -4089 -269 -4055 -255
rect -3071 255 -3037 269
rect -3071 235 -3037 255
rect -3071 187 -3037 197
rect -3071 163 -3037 187
rect -3071 119 -3037 125
rect -3071 91 -3037 119
rect -3071 51 -3037 53
rect -3071 19 -3037 51
rect -3071 -51 -3037 -19
rect -3071 -53 -3037 -51
rect -3071 -119 -3037 -91
rect -3071 -125 -3037 -119
rect -3071 -187 -3037 -163
rect -3071 -197 -3037 -187
rect -3071 -255 -3037 -235
rect -3071 -269 -3037 -255
rect -2053 255 -2019 269
rect -2053 235 -2019 255
rect -2053 187 -2019 197
rect -2053 163 -2019 187
rect -2053 119 -2019 125
rect -2053 91 -2019 119
rect -2053 51 -2019 53
rect -2053 19 -2019 51
rect -2053 -51 -2019 -19
rect -2053 -53 -2019 -51
rect -2053 -119 -2019 -91
rect -2053 -125 -2019 -119
rect -2053 -187 -2019 -163
rect -2053 -197 -2019 -187
rect -2053 -255 -2019 -235
rect -2053 -269 -2019 -255
rect -1035 255 -1001 269
rect -1035 235 -1001 255
rect -1035 187 -1001 197
rect -1035 163 -1001 187
rect -1035 119 -1001 125
rect -1035 91 -1001 119
rect -1035 51 -1001 53
rect -1035 19 -1001 51
rect -1035 -51 -1001 -19
rect -1035 -53 -1001 -51
rect -1035 -119 -1001 -91
rect -1035 -125 -1001 -119
rect -1035 -187 -1001 -163
rect -1035 -197 -1001 -187
rect -1035 -255 -1001 -235
rect -1035 -269 -1001 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 1001 255 1035 269
rect 1001 235 1035 255
rect 1001 187 1035 197
rect 1001 163 1035 187
rect 1001 119 1035 125
rect 1001 91 1035 119
rect 1001 51 1035 53
rect 1001 19 1035 51
rect 1001 -51 1035 -19
rect 1001 -53 1035 -51
rect 1001 -119 1035 -91
rect 1001 -125 1035 -119
rect 1001 -187 1035 -163
rect 1001 -197 1035 -187
rect 1001 -255 1035 -235
rect 1001 -269 1035 -255
rect 2019 255 2053 269
rect 2019 235 2053 255
rect 2019 187 2053 197
rect 2019 163 2053 187
rect 2019 119 2053 125
rect 2019 91 2053 119
rect 2019 51 2053 53
rect 2019 19 2053 51
rect 2019 -51 2053 -19
rect 2019 -53 2053 -51
rect 2019 -119 2053 -91
rect 2019 -125 2053 -119
rect 2019 -187 2053 -163
rect 2019 -197 2053 -187
rect 2019 -255 2053 -235
rect 2019 -269 2053 -255
rect 3037 255 3071 269
rect 3037 235 3071 255
rect 3037 187 3071 197
rect 3037 163 3071 187
rect 3037 119 3071 125
rect 3037 91 3071 119
rect 3037 51 3071 53
rect 3037 19 3071 51
rect 3037 -51 3071 -19
rect 3037 -53 3071 -51
rect 3037 -119 3071 -91
rect 3037 -125 3071 -119
rect 3037 -187 3071 -163
rect 3037 -197 3071 -187
rect 3037 -255 3071 -235
rect 3037 -269 3071 -255
rect 4055 255 4089 269
rect 4055 235 4089 255
rect 4055 187 4089 197
rect 4055 163 4089 187
rect 4055 119 4089 125
rect 4055 91 4089 119
rect 4055 51 4089 53
rect 4055 19 4089 51
rect 4055 -51 4089 -19
rect 4055 -53 4089 -51
rect 4055 -119 4089 -91
rect 4055 -125 4089 -119
rect 4055 -187 4089 -163
rect 4055 -197 4089 -187
rect 4055 -255 4089 -235
rect 4055 -269 4089 -255
rect 5073 255 5107 269
rect 5073 235 5107 255
rect 5073 187 5107 197
rect 5073 163 5107 187
rect 5073 119 5107 125
rect 5073 91 5107 119
rect 5073 51 5107 53
rect 5073 19 5107 51
rect 5073 -51 5107 -19
rect 5073 -53 5107 -51
rect 5073 -119 5107 -91
rect 5073 -125 5107 -119
rect 5073 -187 5107 -163
rect 5073 -197 5107 -187
rect 5073 -255 5107 -235
rect 5073 -269 5107 -255
rect 6091 255 6125 269
rect 6091 235 6125 255
rect 6091 187 6125 197
rect 6091 163 6125 187
rect 6091 119 6125 125
rect 6091 91 6125 119
rect 6091 51 6125 53
rect 6091 19 6125 51
rect 6091 -51 6125 -19
rect 6091 -53 6125 -51
rect 6091 -119 6125 -91
rect 6091 -125 6125 -119
rect 6091 -187 6125 -163
rect 6091 -197 6125 -187
rect 6091 -255 6125 -235
rect 6091 -269 6125 -255
rect 7109 255 7143 269
rect 7109 235 7143 255
rect 7109 187 7143 197
rect 7109 163 7143 187
rect 7109 119 7143 125
rect 7109 91 7143 119
rect 7109 51 7143 53
rect 7109 19 7143 51
rect 7109 -51 7143 -19
rect 7109 -53 7143 -51
rect 7109 -119 7143 -91
rect 7109 -125 7143 -119
rect 7109 -187 7143 -163
rect 7109 -197 7143 -187
rect 7109 -255 7143 -235
rect 7109 -269 7143 -255
rect 8127 255 8161 269
rect 8127 235 8161 255
rect 8127 187 8161 197
rect 8127 163 8161 187
rect 8127 119 8161 125
rect 8127 91 8161 119
rect 8127 51 8161 53
rect 8127 19 8161 51
rect 8127 -51 8161 -19
rect 8127 -53 8161 -51
rect 8127 -119 8161 -91
rect 8127 -125 8161 -119
rect 8127 -187 8161 -163
rect 8127 -197 8161 -187
rect 8127 -255 8161 -235
rect 8127 -269 8161 -255
rect 9145 255 9179 269
rect 9145 235 9179 255
rect 9145 187 9179 197
rect 9145 163 9179 187
rect 9145 119 9179 125
rect 9145 91 9179 119
rect 9145 51 9179 53
rect 9145 19 9179 51
rect 9145 -51 9179 -19
rect 9145 -53 9179 -51
rect 9145 -119 9179 -91
rect 9145 -125 9179 -119
rect 9145 -187 9179 -163
rect 9145 -197 9179 -187
rect 9145 -255 9179 -235
rect 9145 -269 9179 -255
rect 10163 255 10197 269
rect 10163 235 10197 255
rect 10163 187 10197 197
rect 10163 163 10197 187
rect 10163 119 10197 125
rect 10163 91 10197 119
rect 10163 51 10197 53
rect 10163 19 10197 51
rect 10163 -51 10197 -19
rect 10163 -53 10197 -51
rect 10163 -119 10197 -91
rect 10163 -125 10197 -119
rect 10163 -187 10197 -163
rect 10163 -197 10197 -187
rect 10163 -255 10197 -235
rect 10163 -269 10197 -255
rect -9868 -372 -9858 -338
rect -9858 -372 -9834 -338
rect -9796 -372 -9790 -338
rect -9790 -372 -9762 -338
rect -9724 -372 -9722 -338
rect -9722 -372 -9690 -338
rect -9652 -372 -9620 -338
rect -9620 -372 -9618 -338
rect -9580 -372 -9552 -338
rect -9552 -372 -9546 -338
rect -9508 -372 -9484 -338
rect -9484 -372 -9474 -338
rect -8850 -372 -8840 -338
rect -8840 -372 -8816 -338
rect -8778 -372 -8772 -338
rect -8772 -372 -8744 -338
rect -8706 -372 -8704 -338
rect -8704 -372 -8672 -338
rect -8634 -372 -8602 -338
rect -8602 -372 -8600 -338
rect -8562 -372 -8534 -338
rect -8534 -372 -8528 -338
rect -8490 -372 -8466 -338
rect -8466 -372 -8456 -338
rect -7832 -372 -7822 -338
rect -7822 -372 -7798 -338
rect -7760 -372 -7754 -338
rect -7754 -372 -7726 -338
rect -7688 -372 -7686 -338
rect -7686 -372 -7654 -338
rect -7616 -372 -7584 -338
rect -7584 -372 -7582 -338
rect -7544 -372 -7516 -338
rect -7516 -372 -7510 -338
rect -7472 -372 -7448 -338
rect -7448 -372 -7438 -338
rect -6814 -372 -6804 -338
rect -6804 -372 -6780 -338
rect -6742 -372 -6736 -338
rect -6736 -372 -6708 -338
rect -6670 -372 -6668 -338
rect -6668 -372 -6636 -338
rect -6598 -372 -6566 -338
rect -6566 -372 -6564 -338
rect -6526 -372 -6498 -338
rect -6498 -372 -6492 -338
rect -6454 -372 -6430 -338
rect -6430 -372 -6420 -338
rect -5796 -372 -5786 -338
rect -5786 -372 -5762 -338
rect -5724 -372 -5718 -338
rect -5718 -372 -5690 -338
rect -5652 -372 -5650 -338
rect -5650 -372 -5618 -338
rect -5580 -372 -5548 -338
rect -5548 -372 -5546 -338
rect -5508 -372 -5480 -338
rect -5480 -372 -5474 -338
rect -5436 -372 -5412 -338
rect -5412 -372 -5402 -338
rect -4778 -372 -4768 -338
rect -4768 -372 -4744 -338
rect -4706 -372 -4700 -338
rect -4700 -372 -4672 -338
rect -4634 -372 -4632 -338
rect -4632 -372 -4600 -338
rect -4562 -372 -4530 -338
rect -4530 -372 -4528 -338
rect -4490 -372 -4462 -338
rect -4462 -372 -4456 -338
rect -4418 -372 -4394 -338
rect -4394 -372 -4384 -338
rect -3760 -372 -3750 -338
rect -3750 -372 -3726 -338
rect -3688 -372 -3682 -338
rect -3682 -372 -3654 -338
rect -3616 -372 -3614 -338
rect -3614 -372 -3582 -338
rect -3544 -372 -3512 -338
rect -3512 -372 -3510 -338
rect -3472 -372 -3444 -338
rect -3444 -372 -3438 -338
rect -3400 -372 -3376 -338
rect -3376 -372 -3366 -338
rect -2742 -372 -2732 -338
rect -2732 -372 -2708 -338
rect -2670 -372 -2664 -338
rect -2664 -372 -2636 -338
rect -2598 -372 -2596 -338
rect -2596 -372 -2564 -338
rect -2526 -372 -2494 -338
rect -2494 -372 -2492 -338
rect -2454 -372 -2426 -338
rect -2426 -372 -2420 -338
rect -2382 -372 -2358 -338
rect -2358 -372 -2348 -338
rect -1724 -372 -1714 -338
rect -1714 -372 -1690 -338
rect -1652 -372 -1646 -338
rect -1646 -372 -1618 -338
rect -1580 -372 -1578 -338
rect -1578 -372 -1546 -338
rect -1508 -372 -1476 -338
rect -1476 -372 -1474 -338
rect -1436 -372 -1408 -338
rect -1408 -372 -1402 -338
rect -1364 -372 -1340 -338
rect -1340 -372 -1330 -338
rect -706 -372 -696 -338
rect -696 -372 -672 -338
rect -634 -372 -628 -338
rect -628 -372 -600 -338
rect -562 -372 -560 -338
rect -560 -372 -528 -338
rect -490 -372 -458 -338
rect -458 -372 -456 -338
rect -418 -372 -390 -338
rect -390 -372 -384 -338
rect -346 -372 -322 -338
rect -322 -372 -312 -338
rect 312 -372 322 -338
rect 322 -372 346 -338
rect 384 -372 390 -338
rect 390 -372 418 -338
rect 456 -372 458 -338
rect 458 -372 490 -338
rect 528 -372 560 -338
rect 560 -372 562 -338
rect 600 -372 628 -338
rect 628 -372 634 -338
rect 672 -372 696 -338
rect 696 -372 706 -338
rect 1330 -372 1340 -338
rect 1340 -372 1364 -338
rect 1402 -372 1408 -338
rect 1408 -372 1436 -338
rect 1474 -372 1476 -338
rect 1476 -372 1508 -338
rect 1546 -372 1578 -338
rect 1578 -372 1580 -338
rect 1618 -372 1646 -338
rect 1646 -372 1652 -338
rect 1690 -372 1714 -338
rect 1714 -372 1724 -338
rect 2348 -372 2358 -338
rect 2358 -372 2382 -338
rect 2420 -372 2426 -338
rect 2426 -372 2454 -338
rect 2492 -372 2494 -338
rect 2494 -372 2526 -338
rect 2564 -372 2596 -338
rect 2596 -372 2598 -338
rect 2636 -372 2664 -338
rect 2664 -372 2670 -338
rect 2708 -372 2732 -338
rect 2732 -372 2742 -338
rect 3366 -372 3376 -338
rect 3376 -372 3400 -338
rect 3438 -372 3444 -338
rect 3444 -372 3472 -338
rect 3510 -372 3512 -338
rect 3512 -372 3544 -338
rect 3582 -372 3614 -338
rect 3614 -372 3616 -338
rect 3654 -372 3682 -338
rect 3682 -372 3688 -338
rect 3726 -372 3750 -338
rect 3750 -372 3760 -338
rect 4384 -372 4394 -338
rect 4394 -372 4418 -338
rect 4456 -372 4462 -338
rect 4462 -372 4490 -338
rect 4528 -372 4530 -338
rect 4530 -372 4562 -338
rect 4600 -372 4632 -338
rect 4632 -372 4634 -338
rect 4672 -372 4700 -338
rect 4700 -372 4706 -338
rect 4744 -372 4768 -338
rect 4768 -372 4778 -338
rect 5402 -372 5412 -338
rect 5412 -372 5436 -338
rect 5474 -372 5480 -338
rect 5480 -372 5508 -338
rect 5546 -372 5548 -338
rect 5548 -372 5580 -338
rect 5618 -372 5650 -338
rect 5650 -372 5652 -338
rect 5690 -372 5718 -338
rect 5718 -372 5724 -338
rect 5762 -372 5786 -338
rect 5786 -372 5796 -338
rect 6420 -372 6430 -338
rect 6430 -372 6454 -338
rect 6492 -372 6498 -338
rect 6498 -372 6526 -338
rect 6564 -372 6566 -338
rect 6566 -372 6598 -338
rect 6636 -372 6668 -338
rect 6668 -372 6670 -338
rect 6708 -372 6736 -338
rect 6736 -372 6742 -338
rect 6780 -372 6804 -338
rect 6804 -372 6814 -338
rect 7438 -372 7448 -338
rect 7448 -372 7472 -338
rect 7510 -372 7516 -338
rect 7516 -372 7544 -338
rect 7582 -372 7584 -338
rect 7584 -372 7616 -338
rect 7654 -372 7686 -338
rect 7686 -372 7688 -338
rect 7726 -372 7754 -338
rect 7754 -372 7760 -338
rect 7798 -372 7822 -338
rect 7822 -372 7832 -338
rect 8456 -372 8466 -338
rect 8466 -372 8490 -338
rect 8528 -372 8534 -338
rect 8534 -372 8562 -338
rect 8600 -372 8602 -338
rect 8602 -372 8634 -338
rect 8672 -372 8704 -338
rect 8704 -372 8706 -338
rect 8744 -372 8772 -338
rect 8772 -372 8778 -338
rect 8816 -372 8840 -338
rect 8840 -372 8850 -338
rect 9474 -372 9484 -338
rect 9484 -372 9508 -338
rect 9546 -372 9552 -338
rect 9552 -372 9580 -338
rect 9618 -372 9620 -338
rect 9620 -372 9652 -338
rect 9690 -372 9722 -338
rect 9722 -372 9724 -338
rect 9762 -372 9790 -338
rect 9790 -372 9796 -338
rect 9834 -372 9858 -338
rect 9858 -372 9868 -338
<< metal1 >>
rect -9915 372 -9427 378
rect -9915 338 -9868 372
rect -9834 338 -9796 372
rect -9762 338 -9724 372
rect -9690 338 -9652 372
rect -9618 338 -9580 372
rect -9546 338 -9508 372
rect -9474 338 -9427 372
rect -9915 332 -9427 338
rect -8897 372 -8409 378
rect -8897 338 -8850 372
rect -8816 338 -8778 372
rect -8744 338 -8706 372
rect -8672 338 -8634 372
rect -8600 338 -8562 372
rect -8528 338 -8490 372
rect -8456 338 -8409 372
rect -8897 332 -8409 338
rect -7879 372 -7391 378
rect -7879 338 -7832 372
rect -7798 338 -7760 372
rect -7726 338 -7688 372
rect -7654 338 -7616 372
rect -7582 338 -7544 372
rect -7510 338 -7472 372
rect -7438 338 -7391 372
rect -7879 332 -7391 338
rect -6861 372 -6373 378
rect -6861 338 -6814 372
rect -6780 338 -6742 372
rect -6708 338 -6670 372
rect -6636 338 -6598 372
rect -6564 338 -6526 372
rect -6492 338 -6454 372
rect -6420 338 -6373 372
rect -6861 332 -6373 338
rect -5843 372 -5355 378
rect -5843 338 -5796 372
rect -5762 338 -5724 372
rect -5690 338 -5652 372
rect -5618 338 -5580 372
rect -5546 338 -5508 372
rect -5474 338 -5436 372
rect -5402 338 -5355 372
rect -5843 332 -5355 338
rect -4825 372 -4337 378
rect -4825 338 -4778 372
rect -4744 338 -4706 372
rect -4672 338 -4634 372
rect -4600 338 -4562 372
rect -4528 338 -4490 372
rect -4456 338 -4418 372
rect -4384 338 -4337 372
rect -4825 332 -4337 338
rect -3807 372 -3319 378
rect -3807 338 -3760 372
rect -3726 338 -3688 372
rect -3654 338 -3616 372
rect -3582 338 -3544 372
rect -3510 338 -3472 372
rect -3438 338 -3400 372
rect -3366 338 -3319 372
rect -3807 332 -3319 338
rect -2789 372 -2301 378
rect -2789 338 -2742 372
rect -2708 338 -2670 372
rect -2636 338 -2598 372
rect -2564 338 -2526 372
rect -2492 338 -2454 372
rect -2420 338 -2382 372
rect -2348 338 -2301 372
rect -2789 332 -2301 338
rect -1771 372 -1283 378
rect -1771 338 -1724 372
rect -1690 338 -1652 372
rect -1618 338 -1580 372
rect -1546 338 -1508 372
rect -1474 338 -1436 372
rect -1402 338 -1364 372
rect -1330 338 -1283 372
rect -1771 332 -1283 338
rect -753 372 -265 378
rect -753 338 -706 372
rect -672 338 -634 372
rect -600 338 -562 372
rect -528 338 -490 372
rect -456 338 -418 372
rect -384 338 -346 372
rect -312 338 -265 372
rect -753 332 -265 338
rect 265 372 753 378
rect 265 338 312 372
rect 346 338 384 372
rect 418 338 456 372
rect 490 338 528 372
rect 562 338 600 372
rect 634 338 672 372
rect 706 338 753 372
rect 265 332 753 338
rect 1283 372 1771 378
rect 1283 338 1330 372
rect 1364 338 1402 372
rect 1436 338 1474 372
rect 1508 338 1546 372
rect 1580 338 1618 372
rect 1652 338 1690 372
rect 1724 338 1771 372
rect 1283 332 1771 338
rect 2301 372 2789 378
rect 2301 338 2348 372
rect 2382 338 2420 372
rect 2454 338 2492 372
rect 2526 338 2564 372
rect 2598 338 2636 372
rect 2670 338 2708 372
rect 2742 338 2789 372
rect 2301 332 2789 338
rect 3319 372 3807 378
rect 3319 338 3366 372
rect 3400 338 3438 372
rect 3472 338 3510 372
rect 3544 338 3582 372
rect 3616 338 3654 372
rect 3688 338 3726 372
rect 3760 338 3807 372
rect 3319 332 3807 338
rect 4337 372 4825 378
rect 4337 338 4384 372
rect 4418 338 4456 372
rect 4490 338 4528 372
rect 4562 338 4600 372
rect 4634 338 4672 372
rect 4706 338 4744 372
rect 4778 338 4825 372
rect 4337 332 4825 338
rect 5355 372 5843 378
rect 5355 338 5402 372
rect 5436 338 5474 372
rect 5508 338 5546 372
rect 5580 338 5618 372
rect 5652 338 5690 372
rect 5724 338 5762 372
rect 5796 338 5843 372
rect 5355 332 5843 338
rect 6373 372 6861 378
rect 6373 338 6420 372
rect 6454 338 6492 372
rect 6526 338 6564 372
rect 6598 338 6636 372
rect 6670 338 6708 372
rect 6742 338 6780 372
rect 6814 338 6861 372
rect 6373 332 6861 338
rect 7391 372 7879 378
rect 7391 338 7438 372
rect 7472 338 7510 372
rect 7544 338 7582 372
rect 7616 338 7654 372
rect 7688 338 7726 372
rect 7760 338 7798 372
rect 7832 338 7879 372
rect 7391 332 7879 338
rect 8409 372 8897 378
rect 8409 338 8456 372
rect 8490 338 8528 372
rect 8562 338 8600 372
rect 8634 338 8672 372
rect 8706 338 8744 372
rect 8778 338 8816 372
rect 8850 338 8897 372
rect 8409 332 8897 338
rect 9427 372 9915 378
rect 9427 338 9474 372
rect 9508 338 9546 372
rect 9580 338 9618 372
rect 9652 338 9690 372
rect 9724 338 9762 372
rect 9796 338 9834 372
rect 9868 338 9915 372
rect 9427 332 9915 338
rect -10203 269 -10157 300
rect -10203 235 -10197 269
rect -10163 235 -10157 269
rect -10203 197 -10157 235
rect -10203 163 -10197 197
rect -10163 163 -10157 197
rect -10203 125 -10157 163
rect -10203 91 -10197 125
rect -10163 91 -10157 125
rect -10203 53 -10157 91
rect -10203 19 -10197 53
rect -10163 19 -10157 53
rect -10203 -19 -10157 19
rect -10203 -53 -10197 -19
rect -10163 -53 -10157 -19
rect -10203 -91 -10157 -53
rect -10203 -125 -10197 -91
rect -10163 -125 -10157 -91
rect -10203 -163 -10157 -125
rect -10203 -197 -10197 -163
rect -10163 -197 -10157 -163
rect -10203 -235 -10157 -197
rect -10203 -269 -10197 -235
rect -10163 -269 -10157 -235
rect -10203 -300 -10157 -269
rect -9185 269 -9139 300
rect -9185 235 -9179 269
rect -9145 235 -9139 269
rect -9185 197 -9139 235
rect -9185 163 -9179 197
rect -9145 163 -9139 197
rect -9185 125 -9139 163
rect -9185 91 -9179 125
rect -9145 91 -9139 125
rect -9185 53 -9139 91
rect -9185 19 -9179 53
rect -9145 19 -9139 53
rect -9185 -19 -9139 19
rect -9185 -53 -9179 -19
rect -9145 -53 -9139 -19
rect -9185 -91 -9139 -53
rect -9185 -125 -9179 -91
rect -9145 -125 -9139 -91
rect -9185 -163 -9139 -125
rect -9185 -197 -9179 -163
rect -9145 -197 -9139 -163
rect -9185 -235 -9139 -197
rect -9185 -269 -9179 -235
rect -9145 -269 -9139 -235
rect -9185 -300 -9139 -269
rect -8167 269 -8121 300
rect -8167 235 -8161 269
rect -8127 235 -8121 269
rect -8167 197 -8121 235
rect -8167 163 -8161 197
rect -8127 163 -8121 197
rect -8167 125 -8121 163
rect -8167 91 -8161 125
rect -8127 91 -8121 125
rect -8167 53 -8121 91
rect -8167 19 -8161 53
rect -8127 19 -8121 53
rect -8167 -19 -8121 19
rect -8167 -53 -8161 -19
rect -8127 -53 -8121 -19
rect -8167 -91 -8121 -53
rect -8167 -125 -8161 -91
rect -8127 -125 -8121 -91
rect -8167 -163 -8121 -125
rect -8167 -197 -8161 -163
rect -8127 -197 -8121 -163
rect -8167 -235 -8121 -197
rect -8167 -269 -8161 -235
rect -8127 -269 -8121 -235
rect -8167 -300 -8121 -269
rect -7149 269 -7103 300
rect -7149 235 -7143 269
rect -7109 235 -7103 269
rect -7149 197 -7103 235
rect -7149 163 -7143 197
rect -7109 163 -7103 197
rect -7149 125 -7103 163
rect -7149 91 -7143 125
rect -7109 91 -7103 125
rect -7149 53 -7103 91
rect -7149 19 -7143 53
rect -7109 19 -7103 53
rect -7149 -19 -7103 19
rect -7149 -53 -7143 -19
rect -7109 -53 -7103 -19
rect -7149 -91 -7103 -53
rect -7149 -125 -7143 -91
rect -7109 -125 -7103 -91
rect -7149 -163 -7103 -125
rect -7149 -197 -7143 -163
rect -7109 -197 -7103 -163
rect -7149 -235 -7103 -197
rect -7149 -269 -7143 -235
rect -7109 -269 -7103 -235
rect -7149 -300 -7103 -269
rect -6131 269 -6085 300
rect -6131 235 -6125 269
rect -6091 235 -6085 269
rect -6131 197 -6085 235
rect -6131 163 -6125 197
rect -6091 163 -6085 197
rect -6131 125 -6085 163
rect -6131 91 -6125 125
rect -6091 91 -6085 125
rect -6131 53 -6085 91
rect -6131 19 -6125 53
rect -6091 19 -6085 53
rect -6131 -19 -6085 19
rect -6131 -53 -6125 -19
rect -6091 -53 -6085 -19
rect -6131 -91 -6085 -53
rect -6131 -125 -6125 -91
rect -6091 -125 -6085 -91
rect -6131 -163 -6085 -125
rect -6131 -197 -6125 -163
rect -6091 -197 -6085 -163
rect -6131 -235 -6085 -197
rect -6131 -269 -6125 -235
rect -6091 -269 -6085 -235
rect -6131 -300 -6085 -269
rect -5113 269 -5067 300
rect -5113 235 -5107 269
rect -5073 235 -5067 269
rect -5113 197 -5067 235
rect -5113 163 -5107 197
rect -5073 163 -5067 197
rect -5113 125 -5067 163
rect -5113 91 -5107 125
rect -5073 91 -5067 125
rect -5113 53 -5067 91
rect -5113 19 -5107 53
rect -5073 19 -5067 53
rect -5113 -19 -5067 19
rect -5113 -53 -5107 -19
rect -5073 -53 -5067 -19
rect -5113 -91 -5067 -53
rect -5113 -125 -5107 -91
rect -5073 -125 -5067 -91
rect -5113 -163 -5067 -125
rect -5113 -197 -5107 -163
rect -5073 -197 -5067 -163
rect -5113 -235 -5067 -197
rect -5113 -269 -5107 -235
rect -5073 -269 -5067 -235
rect -5113 -300 -5067 -269
rect -4095 269 -4049 300
rect -4095 235 -4089 269
rect -4055 235 -4049 269
rect -4095 197 -4049 235
rect -4095 163 -4089 197
rect -4055 163 -4049 197
rect -4095 125 -4049 163
rect -4095 91 -4089 125
rect -4055 91 -4049 125
rect -4095 53 -4049 91
rect -4095 19 -4089 53
rect -4055 19 -4049 53
rect -4095 -19 -4049 19
rect -4095 -53 -4089 -19
rect -4055 -53 -4049 -19
rect -4095 -91 -4049 -53
rect -4095 -125 -4089 -91
rect -4055 -125 -4049 -91
rect -4095 -163 -4049 -125
rect -4095 -197 -4089 -163
rect -4055 -197 -4049 -163
rect -4095 -235 -4049 -197
rect -4095 -269 -4089 -235
rect -4055 -269 -4049 -235
rect -4095 -300 -4049 -269
rect -3077 269 -3031 300
rect -3077 235 -3071 269
rect -3037 235 -3031 269
rect -3077 197 -3031 235
rect -3077 163 -3071 197
rect -3037 163 -3031 197
rect -3077 125 -3031 163
rect -3077 91 -3071 125
rect -3037 91 -3031 125
rect -3077 53 -3031 91
rect -3077 19 -3071 53
rect -3037 19 -3031 53
rect -3077 -19 -3031 19
rect -3077 -53 -3071 -19
rect -3037 -53 -3031 -19
rect -3077 -91 -3031 -53
rect -3077 -125 -3071 -91
rect -3037 -125 -3031 -91
rect -3077 -163 -3031 -125
rect -3077 -197 -3071 -163
rect -3037 -197 -3031 -163
rect -3077 -235 -3031 -197
rect -3077 -269 -3071 -235
rect -3037 -269 -3031 -235
rect -3077 -300 -3031 -269
rect -2059 269 -2013 300
rect -2059 235 -2053 269
rect -2019 235 -2013 269
rect -2059 197 -2013 235
rect -2059 163 -2053 197
rect -2019 163 -2013 197
rect -2059 125 -2013 163
rect -2059 91 -2053 125
rect -2019 91 -2013 125
rect -2059 53 -2013 91
rect -2059 19 -2053 53
rect -2019 19 -2013 53
rect -2059 -19 -2013 19
rect -2059 -53 -2053 -19
rect -2019 -53 -2013 -19
rect -2059 -91 -2013 -53
rect -2059 -125 -2053 -91
rect -2019 -125 -2013 -91
rect -2059 -163 -2013 -125
rect -2059 -197 -2053 -163
rect -2019 -197 -2013 -163
rect -2059 -235 -2013 -197
rect -2059 -269 -2053 -235
rect -2019 -269 -2013 -235
rect -2059 -300 -2013 -269
rect -1041 269 -995 300
rect -1041 235 -1035 269
rect -1001 235 -995 269
rect -1041 197 -995 235
rect -1041 163 -1035 197
rect -1001 163 -995 197
rect -1041 125 -995 163
rect -1041 91 -1035 125
rect -1001 91 -995 125
rect -1041 53 -995 91
rect -1041 19 -1035 53
rect -1001 19 -995 53
rect -1041 -19 -995 19
rect -1041 -53 -1035 -19
rect -1001 -53 -995 -19
rect -1041 -91 -995 -53
rect -1041 -125 -1035 -91
rect -1001 -125 -995 -91
rect -1041 -163 -995 -125
rect -1041 -197 -1035 -163
rect -1001 -197 -995 -163
rect -1041 -235 -995 -197
rect -1041 -269 -1035 -235
rect -1001 -269 -995 -235
rect -1041 -300 -995 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 995 269 1041 300
rect 995 235 1001 269
rect 1035 235 1041 269
rect 995 197 1041 235
rect 995 163 1001 197
rect 1035 163 1041 197
rect 995 125 1041 163
rect 995 91 1001 125
rect 1035 91 1041 125
rect 995 53 1041 91
rect 995 19 1001 53
rect 1035 19 1041 53
rect 995 -19 1041 19
rect 995 -53 1001 -19
rect 1035 -53 1041 -19
rect 995 -91 1041 -53
rect 995 -125 1001 -91
rect 1035 -125 1041 -91
rect 995 -163 1041 -125
rect 995 -197 1001 -163
rect 1035 -197 1041 -163
rect 995 -235 1041 -197
rect 995 -269 1001 -235
rect 1035 -269 1041 -235
rect 995 -300 1041 -269
rect 2013 269 2059 300
rect 2013 235 2019 269
rect 2053 235 2059 269
rect 2013 197 2059 235
rect 2013 163 2019 197
rect 2053 163 2059 197
rect 2013 125 2059 163
rect 2013 91 2019 125
rect 2053 91 2059 125
rect 2013 53 2059 91
rect 2013 19 2019 53
rect 2053 19 2059 53
rect 2013 -19 2059 19
rect 2013 -53 2019 -19
rect 2053 -53 2059 -19
rect 2013 -91 2059 -53
rect 2013 -125 2019 -91
rect 2053 -125 2059 -91
rect 2013 -163 2059 -125
rect 2013 -197 2019 -163
rect 2053 -197 2059 -163
rect 2013 -235 2059 -197
rect 2013 -269 2019 -235
rect 2053 -269 2059 -235
rect 2013 -300 2059 -269
rect 3031 269 3077 300
rect 3031 235 3037 269
rect 3071 235 3077 269
rect 3031 197 3077 235
rect 3031 163 3037 197
rect 3071 163 3077 197
rect 3031 125 3077 163
rect 3031 91 3037 125
rect 3071 91 3077 125
rect 3031 53 3077 91
rect 3031 19 3037 53
rect 3071 19 3077 53
rect 3031 -19 3077 19
rect 3031 -53 3037 -19
rect 3071 -53 3077 -19
rect 3031 -91 3077 -53
rect 3031 -125 3037 -91
rect 3071 -125 3077 -91
rect 3031 -163 3077 -125
rect 3031 -197 3037 -163
rect 3071 -197 3077 -163
rect 3031 -235 3077 -197
rect 3031 -269 3037 -235
rect 3071 -269 3077 -235
rect 3031 -300 3077 -269
rect 4049 269 4095 300
rect 4049 235 4055 269
rect 4089 235 4095 269
rect 4049 197 4095 235
rect 4049 163 4055 197
rect 4089 163 4095 197
rect 4049 125 4095 163
rect 4049 91 4055 125
rect 4089 91 4095 125
rect 4049 53 4095 91
rect 4049 19 4055 53
rect 4089 19 4095 53
rect 4049 -19 4095 19
rect 4049 -53 4055 -19
rect 4089 -53 4095 -19
rect 4049 -91 4095 -53
rect 4049 -125 4055 -91
rect 4089 -125 4095 -91
rect 4049 -163 4095 -125
rect 4049 -197 4055 -163
rect 4089 -197 4095 -163
rect 4049 -235 4095 -197
rect 4049 -269 4055 -235
rect 4089 -269 4095 -235
rect 4049 -300 4095 -269
rect 5067 269 5113 300
rect 5067 235 5073 269
rect 5107 235 5113 269
rect 5067 197 5113 235
rect 5067 163 5073 197
rect 5107 163 5113 197
rect 5067 125 5113 163
rect 5067 91 5073 125
rect 5107 91 5113 125
rect 5067 53 5113 91
rect 5067 19 5073 53
rect 5107 19 5113 53
rect 5067 -19 5113 19
rect 5067 -53 5073 -19
rect 5107 -53 5113 -19
rect 5067 -91 5113 -53
rect 5067 -125 5073 -91
rect 5107 -125 5113 -91
rect 5067 -163 5113 -125
rect 5067 -197 5073 -163
rect 5107 -197 5113 -163
rect 5067 -235 5113 -197
rect 5067 -269 5073 -235
rect 5107 -269 5113 -235
rect 5067 -300 5113 -269
rect 6085 269 6131 300
rect 6085 235 6091 269
rect 6125 235 6131 269
rect 6085 197 6131 235
rect 6085 163 6091 197
rect 6125 163 6131 197
rect 6085 125 6131 163
rect 6085 91 6091 125
rect 6125 91 6131 125
rect 6085 53 6131 91
rect 6085 19 6091 53
rect 6125 19 6131 53
rect 6085 -19 6131 19
rect 6085 -53 6091 -19
rect 6125 -53 6131 -19
rect 6085 -91 6131 -53
rect 6085 -125 6091 -91
rect 6125 -125 6131 -91
rect 6085 -163 6131 -125
rect 6085 -197 6091 -163
rect 6125 -197 6131 -163
rect 6085 -235 6131 -197
rect 6085 -269 6091 -235
rect 6125 -269 6131 -235
rect 6085 -300 6131 -269
rect 7103 269 7149 300
rect 7103 235 7109 269
rect 7143 235 7149 269
rect 7103 197 7149 235
rect 7103 163 7109 197
rect 7143 163 7149 197
rect 7103 125 7149 163
rect 7103 91 7109 125
rect 7143 91 7149 125
rect 7103 53 7149 91
rect 7103 19 7109 53
rect 7143 19 7149 53
rect 7103 -19 7149 19
rect 7103 -53 7109 -19
rect 7143 -53 7149 -19
rect 7103 -91 7149 -53
rect 7103 -125 7109 -91
rect 7143 -125 7149 -91
rect 7103 -163 7149 -125
rect 7103 -197 7109 -163
rect 7143 -197 7149 -163
rect 7103 -235 7149 -197
rect 7103 -269 7109 -235
rect 7143 -269 7149 -235
rect 7103 -300 7149 -269
rect 8121 269 8167 300
rect 8121 235 8127 269
rect 8161 235 8167 269
rect 8121 197 8167 235
rect 8121 163 8127 197
rect 8161 163 8167 197
rect 8121 125 8167 163
rect 8121 91 8127 125
rect 8161 91 8167 125
rect 8121 53 8167 91
rect 8121 19 8127 53
rect 8161 19 8167 53
rect 8121 -19 8167 19
rect 8121 -53 8127 -19
rect 8161 -53 8167 -19
rect 8121 -91 8167 -53
rect 8121 -125 8127 -91
rect 8161 -125 8167 -91
rect 8121 -163 8167 -125
rect 8121 -197 8127 -163
rect 8161 -197 8167 -163
rect 8121 -235 8167 -197
rect 8121 -269 8127 -235
rect 8161 -269 8167 -235
rect 8121 -300 8167 -269
rect 9139 269 9185 300
rect 9139 235 9145 269
rect 9179 235 9185 269
rect 9139 197 9185 235
rect 9139 163 9145 197
rect 9179 163 9185 197
rect 9139 125 9185 163
rect 9139 91 9145 125
rect 9179 91 9185 125
rect 9139 53 9185 91
rect 9139 19 9145 53
rect 9179 19 9185 53
rect 9139 -19 9185 19
rect 9139 -53 9145 -19
rect 9179 -53 9185 -19
rect 9139 -91 9185 -53
rect 9139 -125 9145 -91
rect 9179 -125 9185 -91
rect 9139 -163 9185 -125
rect 9139 -197 9145 -163
rect 9179 -197 9185 -163
rect 9139 -235 9185 -197
rect 9139 -269 9145 -235
rect 9179 -269 9185 -235
rect 9139 -300 9185 -269
rect 10157 269 10203 300
rect 10157 235 10163 269
rect 10197 235 10203 269
rect 10157 197 10203 235
rect 10157 163 10163 197
rect 10197 163 10203 197
rect 10157 125 10203 163
rect 10157 91 10163 125
rect 10197 91 10203 125
rect 10157 53 10203 91
rect 10157 19 10163 53
rect 10197 19 10203 53
rect 10157 -19 10203 19
rect 10157 -53 10163 -19
rect 10197 -53 10203 -19
rect 10157 -91 10203 -53
rect 10157 -125 10163 -91
rect 10197 -125 10203 -91
rect 10157 -163 10203 -125
rect 10157 -197 10163 -163
rect 10197 -197 10203 -163
rect 10157 -235 10203 -197
rect 10157 -269 10163 -235
rect 10197 -269 10203 -235
rect 10157 -300 10203 -269
rect -9915 -338 -9427 -332
rect -9915 -372 -9868 -338
rect -9834 -372 -9796 -338
rect -9762 -372 -9724 -338
rect -9690 -372 -9652 -338
rect -9618 -372 -9580 -338
rect -9546 -372 -9508 -338
rect -9474 -372 -9427 -338
rect -9915 -378 -9427 -372
rect -8897 -338 -8409 -332
rect -8897 -372 -8850 -338
rect -8816 -372 -8778 -338
rect -8744 -372 -8706 -338
rect -8672 -372 -8634 -338
rect -8600 -372 -8562 -338
rect -8528 -372 -8490 -338
rect -8456 -372 -8409 -338
rect -8897 -378 -8409 -372
rect -7879 -338 -7391 -332
rect -7879 -372 -7832 -338
rect -7798 -372 -7760 -338
rect -7726 -372 -7688 -338
rect -7654 -372 -7616 -338
rect -7582 -372 -7544 -338
rect -7510 -372 -7472 -338
rect -7438 -372 -7391 -338
rect -7879 -378 -7391 -372
rect -6861 -338 -6373 -332
rect -6861 -372 -6814 -338
rect -6780 -372 -6742 -338
rect -6708 -372 -6670 -338
rect -6636 -372 -6598 -338
rect -6564 -372 -6526 -338
rect -6492 -372 -6454 -338
rect -6420 -372 -6373 -338
rect -6861 -378 -6373 -372
rect -5843 -338 -5355 -332
rect -5843 -372 -5796 -338
rect -5762 -372 -5724 -338
rect -5690 -372 -5652 -338
rect -5618 -372 -5580 -338
rect -5546 -372 -5508 -338
rect -5474 -372 -5436 -338
rect -5402 -372 -5355 -338
rect -5843 -378 -5355 -372
rect -4825 -338 -4337 -332
rect -4825 -372 -4778 -338
rect -4744 -372 -4706 -338
rect -4672 -372 -4634 -338
rect -4600 -372 -4562 -338
rect -4528 -372 -4490 -338
rect -4456 -372 -4418 -338
rect -4384 -372 -4337 -338
rect -4825 -378 -4337 -372
rect -3807 -338 -3319 -332
rect -3807 -372 -3760 -338
rect -3726 -372 -3688 -338
rect -3654 -372 -3616 -338
rect -3582 -372 -3544 -338
rect -3510 -372 -3472 -338
rect -3438 -372 -3400 -338
rect -3366 -372 -3319 -338
rect -3807 -378 -3319 -372
rect -2789 -338 -2301 -332
rect -2789 -372 -2742 -338
rect -2708 -372 -2670 -338
rect -2636 -372 -2598 -338
rect -2564 -372 -2526 -338
rect -2492 -372 -2454 -338
rect -2420 -372 -2382 -338
rect -2348 -372 -2301 -338
rect -2789 -378 -2301 -372
rect -1771 -338 -1283 -332
rect -1771 -372 -1724 -338
rect -1690 -372 -1652 -338
rect -1618 -372 -1580 -338
rect -1546 -372 -1508 -338
rect -1474 -372 -1436 -338
rect -1402 -372 -1364 -338
rect -1330 -372 -1283 -338
rect -1771 -378 -1283 -372
rect -753 -338 -265 -332
rect -753 -372 -706 -338
rect -672 -372 -634 -338
rect -600 -372 -562 -338
rect -528 -372 -490 -338
rect -456 -372 -418 -338
rect -384 -372 -346 -338
rect -312 -372 -265 -338
rect -753 -378 -265 -372
rect 265 -338 753 -332
rect 265 -372 312 -338
rect 346 -372 384 -338
rect 418 -372 456 -338
rect 490 -372 528 -338
rect 562 -372 600 -338
rect 634 -372 672 -338
rect 706 -372 753 -338
rect 265 -378 753 -372
rect 1283 -338 1771 -332
rect 1283 -372 1330 -338
rect 1364 -372 1402 -338
rect 1436 -372 1474 -338
rect 1508 -372 1546 -338
rect 1580 -372 1618 -338
rect 1652 -372 1690 -338
rect 1724 -372 1771 -338
rect 1283 -378 1771 -372
rect 2301 -338 2789 -332
rect 2301 -372 2348 -338
rect 2382 -372 2420 -338
rect 2454 -372 2492 -338
rect 2526 -372 2564 -338
rect 2598 -372 2636 -338
rect 2670 -372 2708 -338
rect 2742 -372 2789 -338
rect 2301 -378 2789 -372
rect 3319 -338 3807 -332
rect 3319 -372 3366 -338
rect 3400 -372 3438 -338
rect 3472 -372 3510 -338
rect 3544 -372 3582 -338
rect 3616 -372 3654 -338
rect 3688 -372 3726 -338
rect 3760 -372 3807 -338
rect 3319 -378 3807 -372
rect 4337 -338 4825 -332
rect 4337 -372 4384 -338
rect 4418 -372 4456 -338
rect 4490 -372 4528 -338
rect 4562 -372 4600 -338
rect 4634 -372 4672 -338
rect 4706 -372 4744 -338
rect 4778 -372 4825 -338
rect 4337 -378 4825 -372
rect 5355 -338 5843 -332
rect 5355 -372 5402 -338
rect 5436 -372 5474 -338
rect 5508 -372 5546 -338
rect 5580 -372 5618 -338
rect 5652 -372 5690 -338
rect 5724 -372 5762 -338
rect 5796 -372 5843 -338
rect 5355 -378 5843 -372
rect 6373 -338 6861 -332
rect 6373 -372 6420 -338
rect 6454 -372 6492 -338
rect 6526 -372 6564 -338
rect 6598 -372 6636 -338
rect 6670 -372 6708 -338
rect 6742 -372 6780 -338
rect 6814 -372 6861 -338
rect 6373 -378 6861 -372
rect 7391 -338 7879 -332
rect 7391 -372 7438 -338
rect 7472 -372 7510 -338
rect 7544 -372 7582 -338
rect 7616 -372 7654 -338
rect 7688 -372 7726 -338
rect 7760 -372 7798 -338
rect 7832 -372 7879 -338
rect 7391 -378 7879 -372
rect 8409 -338 8897 -332
rect 8409 -372 8456 -338
rect 8490 -372 8528 -338
rect 8562 -372 8600 -338
rect 8634 -372 8672 -338
rect 8706 -372 8744 -338
rect 8778 -372 8816 -338
rect 8850 -372 8897 -338
rect 8409 -378 8897 -372
rect 9427 -338 9915 -332
rect 9427 -372 9474 -338
rect 9508 -372 9546 -338
rect 9580 -372 9618 -338
rect 9652 -372 9690 -338
rect 9724 -372 9762 -338
rect 9796 -372 9834 -338
rect 9868 -372 9915 -338
rect 9427 -378 9915 -372
<< end >>
