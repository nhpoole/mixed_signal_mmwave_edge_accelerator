.subckt dff_stdcell D CLK Q QB VDD VSS
*.ipin D
*.ipin CLK
*.opin Q
*.opin QB
*.ipin VDD
*.ipin VSS
x12 CLK D VSS VSS VDD VDD Q QB sky130_fd_sc_hd__dfxbp_1
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfxbp/sky130_fd_sc_hd__dfxbp_1.spice

**** end user architecture code
**.ends
** flattened .save nodes
.ends
