magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1374 -3060 4100 5000
<< nwell >>
rect 402 846 2798 3698
rect 10 522 2798 846
<< pwell >>
rect 412 196 2788 348
rect 412 -1596 564 196
rect 2636 -1596 2788 196
rect 412 -1748 2788 -1596
<< psubdiff >>
rect 438 289 2762 322
rect 438 255 631 289
rect 665 255 699 289
rect 733 255 767 289
rect 801 255 835 289
rect 869 255 903 289
rect 937 255 971 289
rect 1005 255 1039 289
rect 1073 255 1107 289
rect 1141 255 1175 289
rect 1209 255 1243 289
rect 1277 255 1311 289
rect 1345 255 1379 289
rect 1413 255 1447 289
rect 1481 255 1515 289
rect 1549 255 1583 289
rect 1617 255 1651 289
rect 1685 255 1719 289
rect 1753 255 1787 289
rect 1821 255 1855 289
rect 1889 255 1923 289
rect 1957 255 1991 289
rect 2025 255 2059 289
rect 2093 255 2127 289
rect 2161 255 2195 289
rect 2229 255 2263 289
rect 2297 255 2331 289
rect 2365 255 2399 289
rect 2433 255 2467 289
rect 2501 255 2535 289
rect 2569 255 2762 289
rect 438 222 2762 255
rect 438 133 538 222
rect 438 99 471 133
rect 505 99 538 133
rect 438 65 538 99
rect 438 31 471 65
rect 505 31 538 65
rect 438 -3 538 31
rect 438 -37 471 -3
rect 505 -37 538 -3
rect 438 -71 538 -37
rect 438 -105 471 -71
rect 505 -105 538 -71
rect 438 -139 538 -105
rect 438 -173 471 -139
rect 505 -173 538 -139
rect 438 -207 538 -173
rect 438 -241 471 -207
rect 505 -241 538 -207
rect 438 -275 538 -241
rect 438 -309 471 -275
rect 505 -309 538 -275
rect 438 -343 538 -309
rect 438 -377 471 -343
rect 505 -377 538 -343
rect 438 -411 538 -377
rect 438 -445 471 -411
rect 505 -445 538 -411
rect 438 -479 538 -445
rect 438 -513 471 -479
rect 505 -513 538 -479
rect 438 -547 538 -513
rect 438 -581 471 -547
rect 505 -581 538 -547
rect 438 -615 538 -581
rect 438 -649 471 -615
rect 505 -649 538 -615
rect 438 -683 538 -649
rect 438 -717 471 -683
rect 505 -717 538 -683
rect 438 -751 538 -717
rect 438 -785 471 -751
rect 505 -785 538 -751
rect 438 -819 538 -785
rect 438 -853 471 -819
rect 505 -853 538 -819
rect 438 -887 538 -853
rect 438 -921 471 -887
rect 505 -921 538 -887
rect 438 -955 538 -921
rect 438 -989 471 -955
rect 505 -989 538 -955
rect 438 -1023 538 -989
rect 438 -1057 471 -1023
rect 505 -1057 538 -1023
rect 438 -1091 538 -1057
rect 438 -1125 471 -1091
rect 505 -1125 538 -1091
rect 438 -1159 538 -1125
rect 438 -1193 471 -1159
rect 505 -1193 538 -1159
rect 438 -1227 538 -1193
rect 438 -1261 471 -1227
rect 505 -1261 538 -1227
rect 438 -1295 538 -1261
rect 438 -1329 471 -1295
rect 505 -1329 538 -1295
rect 438 -1363 538 -1329
rect 438 -1397 471 -1363
rect 505 -1397 538 -1363
rect 438 -1431 538 -1397
rect 438 -1465 471 -1431
rect 505 -1465 538 -1431
rect 438 -1499 538 -1465
rect 438 -1533 471 -1499
rect 505 -1533 538 -1499
rect 438 -1622 538 -1533
rect 2662 133 2762 222
rect 2662 99 2695 133
rect 2729 99 2762 133
rect 2662 65 2762 99
rect 2662 31 2695 65
rect 2729 31 2762 65
rect 2662 -3 2762 31
rect 2662 -37 2695 -3
rect 2729 -37 2762 -3
rect 2662 -71 2762 -37
rect 2662 -105 2695 -71
rect 2729 -105 2762 -71
rect 2662 -139 2762 -105
rect 2662 -173 2695 -139
rect 2729 -173 2762 -139
rect 2662 -207 2762 -173
rect 2662 -241 2695 -207
rect 2729 -241 2762 -207
rect 2662 -275 2762 -241
rect 2662 -309 2695 -275
rect 2729 -309 2762 -275
rect 2662 -343 2762 -309
rect 2662 -377 2695 -343
rect 2729 -377 2762 -343
rect 2662 -411 2762 -377
rect 2662 -445 2695 -411
rect 2729 -445 2762 -411
rect 2662 -479 2762 -445
rect 2662 -513 2695 -479
rect 2729 -513 2762 -479
rect 2662 -547 2762 -513
rect 2662 -581 2695 -547
rect 2729 -581 2762 -547
rect 2662 -615 2762 -581
rect 2662 -649 2695 -615
rect 2729 -649 2762 -615
rect 2662 -683 2762 -649
rect 2662 -717 2695 -683
rect 2729 -717 2762 -683
rect 2662 -751 2762 -717
rect 2662 -785 2695 -751
rect 2729 -785 2762 -751
rect 2662 -819 2762 -785
rect 2662 -853 2695 -819
rect 2729 -853 2762 -819
rect 2662 -887 2762 -853
rect 2662 -921 2695 -887
rect 2729 -921 2762 -887
rect 2662 -955 2762 -921
rect 2662 -989 2695 -955
rect 2729 -989 2762 -955
rect 2662 -1023 2762 -989
rect 2662 -1057 2695 -1023
rect 2729 -1057 2762 -1023
rect 2662 -1091 2762 -1057
rect 2662 -1125 2695 -1091
rect 2729 -1125 2762 -1091
rect 2662 -1159 2762 -1125
rect 2662 -1193 2695 -1159
rect 2729 -1193 2762 -1159
rect 2662 -1227 2762 -1193
rect 2662 -1261 2695 -1227
rect 2729 -1261 2762 -1227
rect 2662 -1295 2762 -1261
rect 2662 -1329 2695 -1295
rect 2729 -1329 2762 -1295
rect 2662 -1363 2762 -1329
rect 2662 -1397 2695 -1363
rect 2729 -1397 2762 -1363
rect 2662 -1431 2762 -1397
rect 2662 -1465 2695 -1431
rect 2729 -1465 2762 -1431
rect 2662 -1499 2762 -1465
rect 2662 -1533 2695 -1499
rect 2729 -1533 2762 -1499
rect 2662 -1622 2762 -1533
rect 438 -1655 2762 -1622
rect 438 -1689 631 -1655
rect 665 -1689 699 -1655
rect 733 -1689 767 -1655
rect 801 -1689 835 -1655
rect 869 -1689 903 -1655
rect 937 -1689 971 -1655
rect 1005 -1689 1039 -1655
rect 1073 -1689 1107 -1655
rect 1141 -1689 1175 -1655
rect 1209 -1689 1243 -1655
rect 1277 -1689 1311 -1655
rect 1345 -1689 1379 -1655
rect 1413 -1689 1447 -1655
rect 1481 -1689 1515 -1655
rect 1549 -1689 1583 -1655
rect 1617 -1689 1651 -1655
rect 1685 -1689 1719 -1655
rect 1753 -1689 1787 -1655
rect 1821 -1689 1855 -1655
rect 1889 -1689 1923 -1655
rect 1957 -1689 1991 -1655
rect 2025 -1689 2059 -1655
rect 2093 -1689 2127 -1655
rect 2161 -1689 2195 -1655
rect 2229 -1689 2263 -1655
rect 2297 -1689 2331 -1655
rect 2365 -1689 2399 -1655
rect 2433 -1689 2467 -1655
rect 2501 -1689 2535 -1655
rect 2569 -1689 2762 -1655
rect 438 -1722 2762 -1689
<< nsubdiff >>
rect 438 3629 2762 3662
rect 438 3595 631 3629
rect 665 3595 699 3629
rect 733 3595 767 3629
rect 801 3595 835 3629
rect 869 3595 903 3629
rect 937 3595 971 3629
rect 1005 3595 1039 3629
rect 1073 3595 1107 3629
rect 1141 3595 1175 3629
rect 1209 3595 1243 3629
rect 1277 3595 1311 3629
rect 1345 3595 1379 3629
rect 1413 3595 1447 3629
rect 1481 3595 1515 3629
rect 1549 3595 1583 3629
rect 1617 3595 1651 3629
rect 1685 3595 1719 3629
rect 1753 3595 1787 3629
rect 1821 3595 1855 3629
rect 1889 3595 1923 3629
rect 1957 3595 1991 3629
rect 2025 3595 2059 3629
rect 2093 3595 2127 3629
rect 2161 3595 2195 3629
rect 2229 3595 2263 3629
rect 2297 3595 2331 3629
rect 2365 3595 2399 3629
rect 2433 3595 2467 3629
rect 2501 3595 2535 3629
rect 2569 3595 2762 3629
rect 438 3562 2762 3595
rect 438 3487 538 3562
rect 438 3453 471 3487
rect 505 3453 538 3487
rect 438 3419 538 3453
rect 438 3385 471 3419
rect 505 3385 538 3419
rect 438 3351 538 3385
rect 438 3317 471 3351
rect 505 3317 538 3351
rect 438 3283 538 3317
rect 438 3249 471 3283
rect 505 3249 538 3283
rect 438 3215 538 3249
rect 438 3181 471 3215
rect 505 3181 538 3215
rect 438 3147 538 3181
rect 438 3113 471 3147
rect 505 3113 538 3147
rect 438 3079 538 3113
rect 438 3045 471 3079
rect 505 3045 538 3079
rect 438 3011 538 3045
rect 438 2977 471 3011
rect 505 2977 538 3011
rect 438 2943 538 2977
rect 438 2909 471 2943
rect 505 2909 538 2943
rect 438 2875 538 2909
rect 438 2841 471 2875
rect 505 2841 538 2875
rect 438 2807 538 2841
rect 438 2773 471 2807
rect 505 2773 538 2807
rect 438 2739 538 2773
rect 438 2705 471 2739
rect 505 2705 538 2739
rect 438 2671 538 2705
rect 438 2637 471 2671
rect 505 2637 538 2671
rect 438 2603 538 2637
rect 438 2569 471 2603
rect 505 2569 538 2603
rect 438 2535 538 2569
rect 438 2501 471 2535
rect 505 2501 538 2535
rect 438 2467 538 2501
rect 438 2433 471 2467
rect 505 2433 538 2467
rect 438 2399 538 2433
rect 438 2365 471 2399
rect 505 2365 538 2399
rect 438 2331 538 2365
rect 438 2297 471 2331
rect 505 2297 538 2331
rect 438 2263 538 2297
rect 438 2229 471 2263
rect 505 2229 538 2263
rect 438 2195 538 2229
rect 438 2161 471 2195
rect 505 2161 538 2195
rect 438 2127 538 2161
rect 438 2093 471 2127
rect 505 2093 538 2127
rect 438 2059 538 2093
rect 438 2025 471 2059
rect 505 2025 538 2059
rect 438 1991 538 2025
rect 438 1957 471 1991
rect 505 1957 538 1991
rect 438 1923 538 1957
rect 438 1889 471 1923
rect 505 1889 538 1923
rect 438 1855 538 1889
rect 438 1821 471 1855
rect 505 1821 538 1855
rect 438 1787 538 1821
rect 438 1753 471 1787
rect 505 1753 538 1787
rect 438 1719 538 1753
rect 438 1685 471 1719
rect 505 1685 538 1719
rect 438 1651 538 1685
rect 438 1617 471 1651
rect 505 1617 538 1651
rect 438 1583 538 1617
rect 438 1549 471 1583
rect 505 1549 538 1583
rect 438 1515 538 1549
rect 438 1481 471 1515
rect 505 1481 538 1515
rect 438 1447 538 1481
rect 438 1413 471 1447
rect 505 1413 538 1447
rect 438 1379 538 1413
rect 438 1345 471 1379
rect 505 1345 538 1379
rect 438 1311 538 1345
rect 438 1277 471 1311
rect 505 1277 538 1311
rect 438 1243 538 1277
rect 438 1209 471 1243
rect 505 1209 538 1243
rect 438 1175 538 1209
rect 438 1141 471 1175
rect 505 1141 538 1175
rect 438 1107 538 1141
rect 438 1073 471 1107
rect 505 1073 538 1107
rect 438 1039 538 1073
rect 438 1005 471 1039
rect 505 1005 538 1039
rect 438 971 538 1005
rect 438 937 471 971
rect 505 937 538 971
rect 438 903 538 937
rect 438 869 471 903
rect 505 869 538 903
rect 438 835 538 869
rect 438 801 471 835
rect 505 801 538 835
rect 438 767 538 801
rect 438 733 471 767
rect 505 733 538 767
rect 438 658 538 733
rect 2662 3487 2762 3562
rect 2662 3453 2695 3487
rect 2729 3453 2762 3487
rect 2662 3419 2762 3453
rect 2662 3385 2695 3419
rect 2729 3385 2762 3419
rect 2662 3351 2762 3385
rect 2662 3317 2695 3351
rect 2729 3317 2762 3351
rect 2662 3283 2762 3317
rect 2662 3249 2695 3283
rect 2729 3249 2762 3283
rect 2662 3215 2762 3249
rect 2662 3181 2695 3215
rect 2729 3181 2762 3215
rect 2662 3147 2762 3181
rect 2662 3113 2695 3147
rect 2729 3113 2762 3147
rect 2662 3079 2762 3113
rect 2662 3045 2695 3079
rect 2729 3045 2762 3079
rect 2662 3011 2762 3045
rect 2662 2977 2695 3011
rect 2729 2977 2762 3011
rect 2662 2943 2762 2977
rect 2662 2909 2695 2943
rect 2729 2909 2762 2943
rect 2662 2875 2762 2909
rect 2662 2841 2695 2875
rect 2729 2841 2762 2875
rect 2662 2807 2762 2841
rect 2662 2773 2695 2807
rect 2729 2773 2762 2807
rect 2662 2739 2762 2773
rect 2662 2705 2695 2739
rect 2729 2705 2762 2739
rect 2662 2671 2762 2705
rect 2662 2637 2695 2671
rect 2729 2637 2762 2671
rect 2662 2603 2762 2637
rect 2662 2569 2695 2603
rect 2729 2569 2762 2603
rect 2662 2535 2762 2569
rect 2662 2501 2695 2535
rect 2729 2501 2762 2535
rect 2662 2467 2762 2501
rect 2662 2433 2695 2467
rect 2729 2433 2762 2467
rect 2662 2399 2762 2433
rect 2662 2365 2695 2399
rect 2729 2365 2762 2399
rect 2662 2331 2762 2365
rect 2662 2297 2695 2331
rect 2729 2297 2762 2331
rect 2662 2263 2762 2297
rect 2662 2229 2695 2263
rect 2729 2229 2762 2263
rect 2662 2195 2762 2229
rect 2662 2161 2695 2195
rect 2729 2161 2762 2195
rect 2662 2127 2762 2161
rect 2662 2093 2695 2127
rect 2729 2093 2762 2127
rect 2662 2059 2762 2093
rect 2662 2025 2695 2059
rect 2729 2025 2762 2059
rect 2662 1991 2762 2025
rect 2662 1957 2695 1991
rect 2729 1957 2762 1991
rect 2662 1923 2762 1957
rect 2662 1889 2695 1923
rect 2729 1889 2762 1923
rect 2662 1855 2762 1889
rect 2662 1821 2695 1855
rect 2729 1821 2762 1855
rect 2662 1787 2762 1821
rect 2662 1753 2695 1787
rect 2729 1753 2762 1787
rect 2662 1719 2762 1753
rect 2662 1685 2695 1719
rect 2729 1685 2762 1719
rect 2662 1651 2762 1685
rect 2662 1617 2695 1651
rect 2729 1617 2762 1651
rect 2662 1583 2762 1617
rect 2662 1549 2695 1583
rect 2729 1549 2762 1583
rect 2662 1515 2762 1549
rect 2662 1481 2695 1515
rect 2729 1481 2762 1515
rect 2662 1447 2762 1481
rect 2662 1413 2695 1447
rect 2729 1413 2762 1447
rect 2662 1379 2762 1413
rect 2662 1345 2695 1379
rect 2729 1345 2762 1379
rect 2662 1311 2762 1345
rect 2662 1277 2695 1311
rect 2729 1277 2762 1311
rect 2662 1243 2762 1277
rect 2662 1209 2695 1243
rect 2729 1209 2762 1243
rect 2662 1175 2762 1209
rect 2662 1141 2695 1175
rect 2729 1141 2762 1175
rect 2662 1107 2762 1141
rect 2662 1073 2695 1107
rect 2729 1073 2762 1107
rect 2662 1039 2762 1073
rect 2662 1005 2695 1039
rect 2729 1005 2762 1039
rect 2662 971 2762 1005
rect 2662 937 2695 971
rect 2729 937 2762 971
rect 2662 903 2762 937
rect 2662 869 2695 903
rect 2729 869 2762 903
rect 2662 835 2762 869
rect 2662 801 2695 835
rect 2729 801 2762 835
rect 2662 767 2762 801
rect 2662 733 2695 767
rect 2729 733 2762 767
rect 2662 658 2762 733
rect 438 625 2762 658
rect 438 591 631 625
rect 665 591 699 625
rect 733 591 767 625
rect 801 591 835 625
rect 869 591 903 625
rect 937 591 971 625
rect 1005 591 1039 625
rect 1073 591 1107 625
rect 1141 591 1175 625
rect 1209 591 1243 625
rect 1277 591 1311 625
rect 1345 591 1379 625
rect 1413 591 1447 625
rect 1481 591 1515 625
rect 1549 591 1583 625
rect 1617 591 1651 625
rect 1685 591 1719 625
rect 1753 591 1787 625
rect 1821 591 1855 625
rect 1889 591 1923 625
rect 1957 591 1991 625
rect 2025 591 2059 625
rect 2093 591 2127 625
rect 2161 591 2195 625
rect 2229 591 2263 625
rect 2297 591 2331 625
rect 2365 591 2399 625
rect 2433 591 2467 625
rect 2501 591 2535 625
rect 2569 591 2762 625
rect 438 558 2762 591
<< psubdiffcont >>
rect 631 255 665 289
rect 699 255 733 289
rect 767 255 801 289
rect 835 255 869 289
rect 903 255 937 289
rect 971 255 1005 289
rect 1039 255 1073 289
rect 1107 255 1141 289
rect 1175 255 1209 289
rect 1243 255 1277 289
rect 1311 255 1345 289
rect 1379 255 1413 289
rect 1447 255 1481 289
rect 1515 255 1549 289
rect 1583 255 1617 289
rect 1651 255 1685 289
rect 1719 255 1753 289
rect 1787 255 1821 289
rect 1855 255 1889 289
rect 1923 255 1957 289
rect 1991 255 2025 289
rect 2059 255 2093 289
rect 2127 255 2161 289
rect 2195 255 2229 289
rect 2263 255 2297 289
rect 2331 255 2365 289
rect 2399 255 2433 289
rect 2467 255 2501 289
rect 2535 255 2569 289
rect 471 99 505 133
rect 471 31 505 65
rect 471 -37 505 -3
rect 471 -105 505 -71
rect 471 -173 505 -139
rect 471 -241 505 -207
rect 471 -309 505 -275
rect 471 -377 505 -343
rect 471 -445 505 -411
rect 471 -513 505 -479
rect 471 -581 505 -547
rect 471 -649 505 -615
rect 471 -717 505 -683
rect 471 -785 505 -751
rect 471 -853 505 -819
rect 471 -921 505 -887
rect 471 -989 505 -955
rect 471 -1057 505 -1023
rect 471 -1125 505 -1091
rect 471 -1193 505 -1159
rect 471 -1261 505 -1227
rect 471 -1329 505 -1295
rect 471 -1397 505 -1363
rect 471 -1465 505 -1431
rect 471 -1533 505 -1499
rect 2695 99 2729 133
rect 2695 31 2729 65
rect 2695 -37 2729 -3
rect 2695 -105 2729 -71
rect 2695 -173 2729 -139
rect 2695 -241 2729 -207
rect 2695 -309 2729 -275
rect 2695 -377 2729 -343
rect 2695 -445 2729 -411
rect 2695 -513 2729 -479
rect 2695 -581 2729 -547
rect 2695 -649 2729 -615
rect 2695 -717 2729 -683
rect 2695 -785 2729 -751
rect 2695 -853 2729 -819
rect 2695 -921 2729 -887
rect 2695 -989 2729 -955
rect 2695 -1057 2729 -1023
rect 2695 -1125 2729 -1091
rect 2695 -1193 2729 -1159
rect 2695 -1261 2729 -1227
rect 2695 -1329 2729 -1295
rect 2695 -1397 2729 -1363
rect 2695 -1465 2729 -1431
rect 2695 -1533 2729 -1499
rect 631 -1689 665 -1655
rect 699 -1689 733 -1655
rect 767 -1689 801 -1655
rect 835 -1689 869 -1655
rect 903 -1689 937 -1655
rect 971 -1689 1005 -1655
rect 1039 -1689 1073 -1655
rect 1107 -1689 1141 -1655
rect 1175 -1689 1209 -1655
rect 1243 -1689 1277 -1655
rect 1311 -1689 1345 -1655
rect 1379 -1689 1413 -1655
rect 1447 -1689 1481 -1655
rect 1515 -1689 1549 -1655
rect 1583 -1689 1617 -1655
rect 1651 -1689 1685 -1655
rect 1719 -1689 1753 -1655
rect 1787 -1689 1821 -1655
rect 1855 -1689 1889 -1655
rect 1923 -1689 1957 -1655
rect 1991 -1689 2025 -1655
rect 2059 -1689 2093 -1655
rect 2127 -1689 2161 -1655
rect 2195 -1689 2229 -1655
rect 2263 -1689 2297 -1655
rect 2331 -1689 2365 -1655
rect 2399 -1689 2433 -1655
rect 2467 -1689 2501 -1655
rect 2535 -1689 2569 -1655
<< nsubdiffcont >>
rect 631 3595 665 3629
rect 699 3595 733 3629
rect 767 3595 801 3629
rect 835 3595 869 3629
rect 903 3595 937 3629
rect 971 3595 1005 3629
rect 1039 3595 1073 3629
rect 1107 3595 1141 3629
rect 1175 3595 1209 3629
rect 1243 3595 1277 3629
rect 1311 3595 1345 3629
rect 1379 3595 1413 3629
rect 1447 3595 1481 3629
rect 1515 3595 1549 3629
rect 1583 3595 1617 3629
rect 1651 3595 1685 3629
rect 1719 3595 1753 3629
rect 1787 3595 1821 3629
rect 1855 3595 1889 3629
rect 1923 3595 1957 3629
rect 1991 3595 2025 3629
rect 2059 3595 2093 3629
rect 2127 3595 2161 3629
rect 2195 3595 2229 3629
rect 2263 3595 2297 3629
rect 2331 3595 2365 3629
rect 2399 3595 2433 3629
rect 2467 3595 2501 3629
rect 2535 3595 2569 3629
rect 471 3453 505 3487
rect 471 3385 505 3419
rect 471 3317 505 3351
rect 471 3249 505 3283
rect 471 3181 505 3215
rect 471 3113 505 3147
rect 471 3045 505 3079
rect 471 2977 505 3011
rect 471 2909 505 2943
rect 471 2841 505 2875
rect 471 2773 505 2807
rect 471 2705 505 2739
rect 471 2637 505 2671
rect 471 2569 505 2603
rect 471 2501 505 2535
rect 471 2433 505 2467
rect 471 2365 505 2399
rect 471 2297 505 2331
rect 471 2229 505 2263
rect 471 2161 505 2195
rect 471 2093 505 2127
rect 471 2025 505 2059
rect 471 1957 505 1991
rect 471 1889 505 1923
rect 471 1821 505 1855
rect 471 1753 505 1787
rect 471 1685 505 1719
rect 471 1617 505 1651
rect 471 1549 505 1583
rect 471 1481 505 1515
rect 471 1413 505 1447
rect 471 1345 505 1379
rect 471 1277 505 1311
rect 471 1209 505 1243
rect 471 1141 505 1175
rect 471 1073 505 1107
rect 471 1005 505 1039
rect 471 937 505 971
rect 471 869 505 903
rect 471 801 505 835
rect 471 733 505 767
rect 2695 3453 2729 3487
rect 2695 3385 2729 3419
rect 2695 3317 2729 3351
rect 2695 3249 2729 3283
rect 2695 3181 2729 3215
rect 2695 3113 2729 3147
rect 2695 3045 2729 3079
rect 2695 2977 2729 3011
rect 2695 2909 2729 2943
rect 2695 2841 2729 2875
rect 2695 2773 2729 2807
rect 2695 2705 2729 2739
rect 2695 2637 2729 2671
rect 2695 2569 2729 2603
rect 2695 2501 2729 2535
rect 2695 2433 2729 2467
rect 2695 2365 2729 2399
rect 2695 2297 2729 2331
rect 2695 2229 2729 2263
rect 2695 2161 2729 2195
rect 2695 2093 2729 2127
rect 2695 2025 2729 2059
rect 2695 1957 2729 1991
rect 2695 1889 2729 1923
rect 2695 1821 2729 1855
rect 2695 1753 2729 1787
rect 2695 1685 2729 1719
rect 2695 1617 2729 1651
rect 2695 1549 2729 1583
rect 2695 1481 2729 1515
rect 2695 1413 2729 1447
rect 2695 1345 2729 1379
rect 2695 1277 2729 1311
rect 2695 1209 2729 1243
rect 2695 1141 2729 1175
rect 2695 1073 2729 1107
rect 2695 1005 2729 1039
rect 2695 937 2729 971
rect 2695 869 2729 903
rect 2695 801 2729 835
rect 2695 733 2729 767
rect 631 591 665 625
rect 699 591 733 625
rect 767 591 801 625
rect 835 591 869 625
rect 903 591 937 625
rect 971 591 1005 625
rect 1039 591 1073 625
rect 1107 591 1141 625
rect 1175 591 1209 625
rect 1243 591 1277 625
rect 1311 591 1345 625
rect 1379 591 1413 625
rect 1447 591 1481 625
rect 1515 591 1549 625
rect 1583 591 1617 625
rect 1651 591 1685 625
rect 1719 591 1753 625
rect 1787 591 1821 625
rect 1855 591 1889 625
rect 1923 591 1957 625
rect 1991 591 2025 625
rect 2059 591 2093 625
rect 2127 591 2161 625
rect 2195 591 2229 625
rect 2263 591 2297 625
rect 2331 591 2365 625
rect 2399 591 2433 625
rect 2467 591 2501 625
rect 2535 591 2569 625
<< locali >>
rect 438 3629 2762 3662
rect 438 3595 539 3629
rect 573 3595 611 3629
rect 665 3595 683 3629
rect 733 3595 755 3629
rect 801 3595 827 3629
rect 869 3595 899 3629
rect 937 3595 971 3629
rect 1005 3595 1039 3629
rect 1077 3595 1107 3629
rect 1149 3595 1175 3629
rect 1221 3595 1243 3629
rect 1293 3595 1311 3629
rect 1365 3595 1379 3629
rect 1437 3595 1447 3629
rect 1509 3595 1515 3629
rect 1581 3595 1583 3629
rect 1617 3595 1619 3629
rect 1685 3595 1691 3629
rect 1753 3595 1763 3629
rect 1821 3595 1835 3629
rect 1889 3595 1907 3629
rect 1957 3595 1979 3629
rect 2025 3595 2051 3629
rect 2093 3595 2123 3629
rect 2161 3595 2195 3629
rect 2229 3595 2263 3629
rect 2301 3595 2331 3629
rect 2373 3595 2399 3629
rect 2445 3595 2467 3629
rect 2517 3595 2535 3629
rect 2589 3595 2627 3629
rect 2661 3595 2762 3629
rect 438 3562 2762 3595
rect 438 3487 538 3562
rect 438 3453 471 3487
rect 505 3453 538 3487
rect 438 3419 538 3453
rect 438 3353 471 3419
rect 505 3353 538 3419
rect 438 3351 538 3353
rect 438 3317 471 3351
rect 505 3317 538 3351
rect 438 3315 538 3317
rect 438 3249 471 3315
rect 505 3249 538 3315
rect 438 3243 538 3249
rect 438 3181 471 3243
rect 505 3181 538 3243
rect 438 3171 538 3181
rect 438 3113 471 3171
rect 505 3113 538 3171
rect 438 3099 538 3113
rect 438 3045 471 3099
rect 505 3045 538 3099
rect 438 3027 538 3045
rect 438 2977 471 3027
rect 505 2977 538 3027
rect 438 2955 538 2977
rect 438 2909 471 2955
rect 505 2909 538 2955
rect 438 2883 538 2909
rect 438 2841 471 2883
rect 505 2841 538 2883
rect 438 2811 538 2841
rect 438 2773 471 2811
rect 505 2773 538 2811
rect 438 2739 538 2773
rect 438 2705 471 2739
rect 505 2705 538 2739
rect 438 2671 538 2705
rect 438 2633 471 2671
rect 505 2633 538 2671
rect 438 2603 538 2633
rect 438 2561 471 2603
rect 505 2561 538 2603
rect 438 2535 538 2561
rect 438 2489 471 2535
rect 505 2489 538 2535
rect 438 2467 538 2489
rect 438 2417 471 2467
rect 505 2417 538 2467
rect 438 2399 538 2417
rect 438 2345 471 2399
rect 505 2345 538 2399
rect 438 2331 538 2345
rect 438 2273 471 2331
rect 505 2273 538 2331
rect 438 2263 538 2273
rect 438 2201 471 2263
rect 505 2201 538 2263
rect 438 2195 538 2201
rect 438 2129 471 2195
rect 505 2129 538 2195
rect 438 2127 538 2129
rect 438 2093 471 2127
rect 505 2093 538 2127
rect 438 2091 538 2093
rect 438 2025 471 2091
rect 505 2025 538 2091
rect 438 2019 538 2025
rect 438 1957 471 2019
rect 505 1957 538 2019
rect 438 1947 538 1957
rect 438 1889 471 1947
rect 505 1889 538 1947
rect 438 1875 538 1889
rect 438 1821 471 1875
rect 505 1821 538 1875
rect 438 1803 538 1821
rect 438 1753 471 1803
rect 505 1753 538 1803
rect 438 1731 538 1753
rect 438 1685 471 1731
rect 505 1685 538 1731
rect 438 1659 538 1685
rect 438 1617 471 1659
rect 505 1617 538 1659
rect 438 1587 538 1617
rect 438 1549 471 1587
rect 505 1549 538 1587
rect 438 1515 538 1549
rect 438 1481 471 1515
rect 505 1481 538 1515
rect 438 1447 538 1481
rect 438 1409 471 1447
rect 505 1409 538 1447
rect 438 1379 538 1409
rect 438 1337 471 1379
rect 505 1337 538 1379
rect 438 1311 538 1337
rect 438 1265 471 1311
rect 505 1265 538 1311
rect 438 1243 538 1265
rect 438 1193 471 1243
rect 505 1193 538 1243
rect 438 1175 538 1193
rect 438 1121 471 1175
rect 505 1121 538 1175
rect 438 1107 538 1121
rect 438 1049 471 1107
rect 505 1049 538 1107
rect 438 1039 538 1049
rect 438 977 471 1039
rect 505 977 538 1039
rect 438 971 538 977
rect 438 905 471 971
rect 505 905 538 971
rect 438 903 538 905
rect 438 869 471 903
rect 505 869 538 903
rect 438 867 538 869
rect 438 801 471 867
rect 505 801 538 867
rect 438 767 538 801
rect 438 733 471 767
rect 505 733 538 767
rect 438 658 538 733
rect 2662 3487 2762 3562
rect 2662 3453 2695 3487
rect 2729 3453 2762 3487
rect 2662 3419 2762 3453
rect 2662 3353 2695 3419
rect 2729 3353 2762 3419
rect 2662 3351 2762 3353
rect 2662 3317 2695 3351
rect 2729 3317 2762 3351
rect 2662 3315 2762 3317
rect 2662 3249 2695 3315
rect 2729 3249 2762 3315
rect 2662 3243 2762 3249
rect 2662 3181 2695 3243
rect 2729 3181 2762 3243
rect 2662 3171 2762 3181
rect 2662 3113 2695 3171
rect 2729 3113 2762 3171
rect 2662 3099 2762 3113
rect 2662 3045 2695 3099
rect 2729 3045 2762 3099
rect 2662 3027 2762 3045
rect 2662 2977 2695 3027
rect 2729 2977 2762 3027
rect 2662 2955 2762 2977
rect 2662 2909 2695 2955
rect 2729 2909 2762 2955
rect 2662 2883 2762 2909
rect 2662 2841 2695 2883
rect 2729 2841 2762 2883
rect 2662 2811 2762 2841
rect 2662 2773 2695 2811
rect 2729 2773 2762 2811
rect 2662 2739 2762 2773
rect 2662 2705 2695 2739
rect 2729 2705 2762 2739
rect 2662 2671 2762 2705
rect 2662 2633 2695 2671
rect 2729 2633 2762 2671
rect 2662 2603 2762 2633
rect 2662 2561 2695 2603
rect 2729 2561 2762 2603
rect 2662 2535 2762 2561
rect 2662 2489 2695 2535
rect 2729 2489 2762 2535
rect 2662 2467 2762 2489
rect 2662 2417 2695 2467
rect 2729 2417 2762 2467
rect 2662 2399 2762 2417
rect 2662 2345 2695 2399
rect 2729 2345 2762 2399
rect 2662 2331 2762 2345
rect 2662 2273 2695 2331
rect 2729 2273 2762 2331
rect 2662 2263 2762 2273
rect 2662 2201 2695 2263
rect 2729 2201 2762 2263
rect 2662 2195 2762 2201
rect 2662 2129 2695 2195
rect 2729 2129 2762 2195
rect 2662 2127 2762 2129
rect 2662 2093 2695 2127
rect 2729 2093 2762 2127
rect 2662 2091 2762 2093
rect 2662 2025 2695 2091
rect 2729 2025 2762 2091
rect 2662 2019 2762 2025
rect 2662 1957 2695 2019
rect 2729 1957 2762 2019
rect 2662 1947 2762 1957
rect 2662 1889 2695 1947
rect 2729 1889 2762 1947
rect 2662 1875 2762 1889
rect 2662 1821 2695 1875
rect 2729 1821 2762 1875
rect 2662 1803 2762 1821
rect 2662 1753 2695 1803
rect 2729 1753 2762 1803
rect 2662 1731 2762 1753
rect 2662 1685 2695 1731
rect 2729 1685 2762 1731
rect 2662 1659 2762 1685
rect 2662 1617 2695 1659
rect 2729 1617 2762 1659
rect 2662 1587 2762 1617
rect 2662 1549 2695 1587
rect 2729 1549 2762 1587
rect 2662 1515 2762 1549
rect 2662 1481 2695 1515
rect 2729 1481 2762 1515
rect 2662 1447 2762 1481
rect 2662 1409 2695 1447
rect 2729 1409 2762 1447
rect 2662 1379 2762 1409
rect 2662 1337 2695 1379
rect 2729 1337 2762 1379
rect 2662 1311 2762 1337
rect 2662 1265 2695 1311
rect 2729 1265 2762 1311
rect 2662 1243 2762 1265
rect 2662 1193 2695 1243
rect 2729 1193 2762 1243
rect 2662 1175 2762 1193
rect 2662 1121 2695 1175
rect 2729 1121 2762 1175
rect 2662 1107 2762 1121
rect 2662 1049 2695 1107
rect 2729 1049 2762 1107
rect 2662 1039 2762 1049
rect 2662 977 2695 1039
rect 2729 977 2762 1039
rect 2662 971 2762 977
rect 2662 905 2695 971
rect 2729 905 2762 971
rect 2662 903 2762 905
rect 2662 869 2695 903
rect 2729 869 2762 903
rect 2662 867 2762 869
rect 2662 801 2695 867
rect 2729 801 2762 867
rect 2662 767 2762 801
rect 2662 733 2695 767
rect 2729 733 2762 767
rect 2662 658 2762 733
rect 438 625 2762 658
rect 438 591 539 625
rect 573 591 611 625
rect 665 591 683 625
rect 733 591 755 625
rect 801 591 827 625
rect 869 591 899 625
rect 937 591 971 625
rect 1005 591 1039 625
rect 1077 591 1107 625
rect 1149 591 1175 625
rect 1221 591 1243 625
rect 1293 591 1311 625
rect 1365 591 1379 625
rect 1437 591 1447 625
rect 1509 591 1515 625
rect 1581 591 1583 625
rect 1617 591 1619 625
rect 1685 591 1691 625
rect 1753 591 1763 625
rect 1821 591 1835 625
rect 1889 591 1907 625
rect 1957 591 1979 625
rect 2025 591 2051 625
rect 2093 591 2123 625
rect 2161 591 2195 625
rect 2229 591 2263 625
rect 2301 591 2331 625
rect 2373 591 2399 625
rect 2445 591 2467 625
rect 2517 591 2535 625
rect 2589 591 2627 625
rect 2661 591 2762 625
rect 438 558 2762 591
rect 118 519 166 526
rect 118 485 125 519
rect 159 485 166 519
rect 118 478 166 485
rect 220 461 268 468
rect 220 427 227 461
rect 261 427 268 461
rect 220 420 268 427
rect 438 289 2762 322
rect 438 255 539 289
rect 573 255 611 289
rect 665 255 683 289
rect 733 255 755 289
rect 801 255 827 289
rect 869 255 899 289
rect 937 255 971 289
rect 1005 255 1039 289
rect 1077 255 1107 289
rect 1149 255 1175 289
rect 1221 255 1243 289
rect 1293 255 1311 289
rect 1365 255 1379 289
rect 1437 255 1447 289
rect 1509 255 1515 289
rect 1581 255 1583 289
rect 1617 255 1619 289
rect 1685 255 1691 289
rect 1753 255 1763 289
rect 1821 255 1835 289
rect 1889 255 1907 289
rect 1957 255 1979 289
rect 2025 255 2051 289
rect 2093 255 2123 289
rect 2161 255 2195 289
rect 2229 255 2263 289
rect 2301 255 2331 289
rect 2373 255 2399 289
rect 2445 255 2467 289
rect 2517 255 2535 289
rect 2589 255 2627 289
rect 2661 255 2762 289
rect 438 222 2762 255
rect 438 133 538 222
rect 438 75 471 133
rect 505 75 538 133
rect 438 65 538 75
rect 438 3 471 65
rect 505 3 538 65
rect 438 -3 538 3
rect 438 -69 471 -3
rect 505 -69 538 -3
rect 438 -71 538 -69
rect 438 -105 471 -71
rect 505 -105 538 -71
rect 438 -107 538 -105
rect 438 -173 471 -107
rect 505 -173 538 -107
rect 438 -179 538 -173
rect 438 -241 471 -179
rect 505 -241 538 -179
rect 438 -251 538 -241
rect 438 -309 471 -251
rect 505 -309 538 -251
rect 438 -323 538 -309
rect 438 -377 471 -323
rect 505 -377 538 -323
rect 438 -395 538 -377
rect 438 -445 471 -395
rect 505 -445 538 -395
rect 438 -467 538 -445
rect 438 -513 471 -467
rect 505 -513 538 -467
rect 438 -539 538 -513
rect 438 -581 471 -539
rect 505 -581 538 -539
rect 438 -611 538 -581
rect 438 -649 471 -611
rect 505 -649 538 -611
rect 438 -683 538 -649
rect 438 -717 471 -683
rect 505 -717 538 -683
rect 438 -751 538 -717
rect 438 -789 471 -751
rect 505 -789 538 -751
rect 438 -819 538 -789
rect 438 -861 471 -819
rect 505 -861 538 -819
rect 438 -887 538 -861
rect 438 -933 471 -887
rect 505 -933 538 -887
rect 438 -955 538 -933
rect 438 -1005 471 -955
rect 505 -1005 538 -955
rect 438 -1023 538 -1005
rect 438 -1077 471 -1023
rect 505 -1077 538 -1023
rect 438 -1091 538 -1077
rect 438 -1149 471 -1091
rect 505 -1149 538 -1091
rect 438 -1159 538 -1149
rect 438 -1221 471 -1159
rect 505 -1221 538 -1159
rect 438 -1227 538 -1221
rect 438 -1293 471 -1227
rect 505 -1293 538 -1227
rect 438 -1295 538 -1293
rect 438 -1329 471 -1295
rect 505 -1329 538 -1295
rect 438 -1331 538 -1329
rect 438 -1397 471 -1331
rect 505 -1397 538 -1331
rect 438 -1403 538 -1397
rect 438 -1465 471 -1403
rect 505 -1465 538 -1403
rect 438 -1475 538 -1465
rect 438 -1533 471 -1475
rect 505 -1533 538 -1475
rect 438 -1622 538 -1533
rect 2662 133 2762 222
rect 2662 75 2695 133
rect 2729 75 2762 133
rect 2662 65 2762 75
rect 2662 3 2695 65
rect 2729 3 2762 65
rect 2662 -3 2762 3
rect 2662 -69 2695 -3
rect 2729 -69 2762 -3
rect 2662 -71 2762 -69
rect 2662 -105 2695 -71
rect 2729 -105 2762 -71
rect 2662 -107 2762 -105
rect 2662 -173 2695 -107
rect 2729 -173 2762 -107
rect 2662 -179 2762 -173
rect 2662 -241 2695 -179
rect 2729 -241 2762 -179
rect 2662 -251 2762 -241
rect 2662 -309 2695 -251
rect 2729 -309 2762 -251
rect 2662 -323 2762 -309
rect 2662 -377 2695 -323
rect 2729 -377 2762 -323
rect 2662 -395 2762 -377
rect 2662 -445 2695 -395
rect 2729 -445 2762 -395
rect 2662 -467 2762 -445
rect 2662 -513 2695 -467
rect 2729 -513 2762 -467
rect 2662 -539 2762 -513
rect 2662 -581 2695 -539
rect 2729 -581 2762 -539
rect 2662 -611 2762 -581
rect 2662 -649 2695 -611
rect 2729 -649 2762 -611
rect 2662 -683 2762 -649
rect 2662 -717 2695 -683
rect 2729 -717 2762 -683
rect 2662 -751 2762 -717
rect 2662 -789 2695 -751
rect 2729 -789 2762 -751
rect 2662 -819 2762 -789
rect 2662 -861 2695 -819
rect 2729 -861 2762 -819
rect 2662 -887 2762 -861
rect 2662 -933 2695 -887
rect 2729 -933 2762 -887
rect 2662 -955 2762 -933
rect 2662 -1005 2695 -955
rect 2729 -1005 2762 -955
rect 2662 -1023 2762 -1005
rect 2662 -1077 2695 -1023
rect 2729 -1077 2762 -1023
rect 2662 -1091 2762 -1077
rect 2662 -1149 2695 -1091
rect 2729 -1149 2762 -1091
rect 2662 -1159 2762 -1149
rect 2662 -1221 2695 -1159
rect 2729 -1221 2762 -1159
rect 2662 -1227 2762 -1221
rect 2662 -1293 2695 -1227
rect 2729 -1293 2762 -1227
rect 2662 -1295 2762 -1293
rect 2662 -1329 2695 -1295
rect 2729 -1329 2762 -1295
rect 2662 -1331 2762 -1329
rect 2662 -1397 2695 -1331
rect 2729 -1397 2762 -1331
rect 2662 -1403 2762 -1397
rect 2662 -1465 2695 -1403
rect 2729 -1465 2762 -1403
rect 2662 -1475 2762 -1465
rect 2662 -1533 2695 -1475
rect 2729 -1533 2762 -1475
rect 2662 -1622 2762 -1533
rect 438 -1655 2762 -1622
rect 438 -1689 539 -1655
rect 573 -1689 611 -1655
rect 665 -1689 683 -1655
rect 733 -1689 755 -1655
rect 801 -1689 827 -1655
rect 869 -1689 899 -1655
rect 937 -1689 971 -1655
rect 1005 -1689 1039 -1655
rect 1077 -1689 1107 -1655
rect 1149 -1689 1175 -1655
rect 1221 -1689 1243 -1655
rect 1293 -1689 1311 -1655
rect 1365 -1689 1379 -1655
rect 1437 -1689 1447 -1655
rect 1509 -1689 1515 -1655
rect 1581 -1689 1583 -1655
rect 1617 -1689 1619 -1655
rect 1685 -1689 1691 -1655
rect 1753 -1689 1763 -1655
rect 1821 -1689 1835 -1655
rect 1889 -1689 1907 -1655
rect 1957 -1689 1979 -1655
rect 2025 -1689 2051 -1655
rect 2093 -1689 2123 -1655
rect 2161 -1689 2195 -1655
rect 2229 -1689 2263 -1655
rect 2301 -1689 2331 -1655
rect 2373 -1689 2399 -1655
rect 2445 -1689 2467 -1655
rect 2517 -1689 2535 -1655
rect 2589 -1689 2627 -1655
rect 2661 -1689 2762 -1655
rect 438 -1722 2762 -1689
<< viali >>
rect 539 3595 573 3629
rect 611 3595 631 3629
rect 631 3595 645 3629
rect 683 3595 699 3629
rect 699 3595 717 3629
rect 755 3595 767 3629
rect 767 3595 789 3629
rect 827 3595 835 3629
rect 835 3595 861 3629
rect 899 3595 903 3629
rect 903 3595 933 3629
rect 971 3595 1005 3629
rect 1043 3595 1073 3629
rect 1073 3595 1077 3629
rect 1115 3595 1141 3629
rect 1141 3595 1149 3629
rect 1187 3595 1209 3629
rect 1209 3595 1221 3629
rect 1259 3595 1277 3629
rect 1277 3595 1293 3629
rect 1331 3595 1345 3629
rect 1345 3595 1365 3629
rect 1403 3595 1413 3629
rect 1413 3595 1437 3629
rect 1475 3595 1481 3629
rect 1481 3595 1509 3629
rect 1547 3595 1549 3629
rect 1549 3595 1581 3629
rect 1619 3595 1651 3629
rect 1651 3595 1653 3629
rect 1691 3595 1719 3629
rect 1719 3595 1725 3629
rect 1763 3595 1787 3629
rect 1787 3595 1797 3629
rect 1835 3595 1855 3629
rect 1855 3595 1869 3629
rect 1907 3595 1923 3629
rect 1923 3595 1941 3629
rect 1979 3595 1991 3629
rect 1991 3595 2013 3629
rect 2051 3595 2059 3629
rect 2059 3595 2085 3629
rect 2123 3595 2127 3629
rect 2127 3595 2157 3629
rect 2195 3595 2229 3629
rect 2267 3595 2297 3629
rect 2297 3595 2301 3629
rect 2339 3595 2365 3629
rect 2365 3595 2373 3629
rect 2411 3595 2433 3629
rect 2433 3595 2445 3629
rect 2483 3595 2501 3629
rect 2501 3595 2517 3629
rect 2555 3595 2569 3629
rect 2569 3595 2589 3629
rect 2627 3595 2661 3629
rect 471 3385 505 3387
rect 471 3353 505 3385
rect 471 3283 505 3315
rect 471 3281 505 3283
rect 471 3215 505 3243
rect 471 3209 505 3215
rect 471 3147 505 3171
rect 471 3137 505 3147
rect 471 3079 505 3099
rect 471 3065 505 3079
rect 471 3011 505 3027
rect 471 2993 505 3011
rect 471 2943 505 2955
rect 471 2921 505 2943
rect 471 2875 505 2883
rect 471 2849 505 2875
rect 471 2807 505 2811
rect 471 2777 505 2807
rect 471 2705 505 2739
rect 471 2637 505 2667
rect 471 2633 505 2637
rect 471 2569 505 2595
rect 471 2561 505 2569
rect 471 2501 505 2523
rect 471 2489 505 2501
rect 471 2433 505 2451
rect 471 2417 505 2433
rect 471 2365 505 2379
rect 471 2345 505 2365
rect 471 2297 505 2307
rect 471 2273 505 2297
rect 471 2229 505 2235
rect 471 2201 505 2229
rect 471 2161 505 2163
rect 471 2129 505 2161
rect 471 2059 505 2091
rect 471 2057 505 2059
rect 471 1991 505 2019
rect 471 1985 505 1991
rect 471 1923 505 1947
rect 471 1913 505 1923
rect 471 1855 505 1875
rect 471 1841 505 1855
rect 471 1787 505 1803
rect 471 1769 505 1787
rect 471 1719 505 1731
rect 471 1697 505 1719
rect 471 1651 505 1659
rect 471 1625 505 1651
rect 471 1583 505 1587
rect 471 1553 505 1583
rect 471 1481 505 1515
rect 471 1413 505 1443
rect 471 1409 505 1413
rect 471 1345 505 1371
rect 471 1337 505 1345
rect 471 1277 505 1299
rect 471 1265 505 1277
rect 471 1209 505 1227
rect 471 1193 505 1209
rect 471 1141 505 1155
rect 471 1121 505 1141
rect 471 1073 505 1083
rect 471 1049 505 1073
rect 471 1005 505 1011
rect 471 977 505 1005
rect 471 937 505 939
rect 471 905 505 937
rect 471 835 505 867
rect 471 833 505 835
rect 2695 3385 2729 3387
rect 2695 3353 2729 3385
rect 2695 3283 2729 3315
rect 2695 3281 2729 3283
rect 2695 3215 2729 3243
rect 2695 3209 2729 3215
rect 2695 3147 2729 3171
rect 2695 3137 2729 3147
rect 2695 3079 2729 3099
rect 2695 3065 2729 3079
rect 2695 3011 2729 3027
rect 2695 2993 2729 3011
rect 2695 2943 2729 2955
rect 2695 2921 2729 2943
rect 2695 2875 2729 2883
rect 2695 2849 2729 2875
rect 2695 2807 2729 2811
rect 2695 2777 2729 2807
rect 2695 2705 2729 2739
rect 2695 2637 2729 2667
rect 2695 2633 2729 2637
rect 2695 2569 2729 2595
rect 2695 2561 2729 2569
rect 2695 2501 2729 2523
rect 2695 2489 2729 2501
rect 2695 2433 2729 2451
rect 2695 2417 2729 2433
rect 2695 2365 2729 2379
rect 2695 2345 2729 2365
rect 2695 2297 2729 2307
rect 2695 2273 2729 2297
rect 2695 2229 2729 2235
rect 2695 2201 2729 2229
rect 2695 2161 2729 2163
rect 2695 2129 2729 2161
rect 2695 2059 2729 2091
rect 2695 2057 2729 2059
rect 2695 1991 2729 2019
rect 2695 1985 2729 1991
rect 2695 1923 2729 1947
rect 2695 1913 2729 1923
rect 2695 1855 2729 1875
rect 2695 1841 2729 1855
rect 2695 1787 2729 1803
rect 2695 1769 2729 1787
rect 2695 1719 2729 1731
rect 2695 1697 2729 1719
rect 2695 1651 2729 1659
rect 2695 1625 2729 1651
rect 2695 1583 2729 1587
rect 2695 1553 2729 1583
rect 2695 1481 2729 1515
rect 2695 1413 2729 1443
rect 2695 1409 2729 1413
rect 2695 1345 2729 1371
rect 2695 1337 2729 1345
rect 2695 1277 2729 1299
rect 2695 1265 2729 1277
rect 2695 1209 2729 1227
rect 2695 1193 2729 1209
rect 2695 1141 2729 1155
rect 2695 1121 2729 1141
rect 2695 1073 2729 1083
rect 2695 1049 2729 1073
rect 2695 1005 2729 1011
rect 2695 977 2729 1005
rect 2695 937 2729 939
rect 2695 905 2729 937
rect 2695 835 2729 867
rect 2695 833 2729 835
rect 539 591 573 625
rect 611 591 631 625
rect 631 591 645 625
rect 683 591 699 625
rect 699 591 717 625
rect 755 591 767 625
rect 767 591 789 625
rect 827 591 835 625
rect 835 591 861 625
rect 899 591 903 625
rect 903 591 933 625
rect 971 591 1005 625
rect 1043 591 1073 625
rect 1073 591 1077 625
rect 1115 591 1141 625
rect 1141 591 1149 625
rect 1187 591 1209 625
rect 1209 591 1221 625
rect 1259 591 1277 625
rect 1277 591 1293 625
rect 1331 591 1345 625
rect 1345 591 1365 625
rect 1403 591 1413 625
rect 1413 591 1437 625
rect 1475 591 1481 625
rect 1481 591 1509 625
rect 1547 591 1549 625
rect 1549 591 1581 625
rect 1619 591 1651 625
rect 1651 591 1653 625
rect 1691 591 1719 625
rect 1719 591 1725 625
rect 1763 591 1787 625
rect 1787 591 1797 625
rect 1835 591 1855 625
rect 1855 591 1869 625
rect 1907 591 1923 625
rect 1923 591 1941 625
rect 1979 591 1991 625
rect 1991 591 2013 625
rect 2051 591 2059 625
rect 2059 591 2085 625
rect 2123 591 2127 625
rect 2127 591 2157 625
rect 2195 591 2229 625
rect 2267 591 2297 625
rect 2297 591 2301 625
rect 2339 591 2365 625
rect 2365 591 2373 625
rect 2411 591 2433 625
rect 2433 591 2445 625
rect 2483 591 2501 625
rect 2501 591 2517 625
rect 2555 591 2569 625
rect 2569 591 2589 625
rect 2627 591 2661 625
rect 125 485 159 519
rect 227 427 261 461
rect 539 255 573 289
rect 611 255 631 289
rect 631 255 645 289
rect 683 255 699 289
rect 699 255 717 289
rect 755 255 767 289
rect 767 255 789 289
rect 827 255 835 289
rect 835 255 861 289
rect 899 255 903 289
rect 903 255 933 289
rect 971 255 1005 289
rect 1043 255 1073 289
rect 1073 255 1077 289
rect 1115 255 1141 289
rect 1141 255 1149 289
rect 1187 255 1209 289
rect 1209 255 1221 289
rect 1259 255 1277 289
rect 1277 255 1293 289
rect 1331 255 1345 289
rect 1345 255 1365 289
rect 1403 255 1413 289
rect 1413 255 1437 289
rect 1475 255 1481 289
rect 1481 255 1509 289
rect 1547 255 1549 289
rect 1549 255 1581 289
rect 1619 255 1651 289
rect 1651 255 1653 289
rect 1691 255 1719 289
rect 1719 255 1725 289
rect 1763 255 1787 289
rect 1787 255 1797 289
rect 1835 255 1855 289
rect 1855 255 1869 289
rect 1907 255 1923 289
rect 1923 255 1941 289
rect 1979 255 1991 289
rect 1991 255 2013 289
rect 2051 255 2059 289
rect 2059 255 2085 289
rect 2123 255 2127 289
rect 2127 255 2157 289
rect 2195 255 2229 289
rect 2267 255 2297 289
rect 2297 255 2301 289
rect 2339 255 2365 289
rect 2365 255 2373 289
rect 2411 255 2433 289
rect 2433 255 2445 289
rect 2483 255 2501 289
rect 2501 255 2517 289
rect 2555 255 2569 289
rect 2569 255 2589 289
rect 2627 255 2661 289
rect 471 99 505 109
rect 471 75 505 99
rect 471 31 505 37
rect 471 3 505 31
rect 471 -37 505 -35
rect 471 -69 505 -37
rect 471 -139 505 -107
rect 471 -141 505 -139
rect 471 -207 505 -179
rect 471 -213 505 -207
rect 471 -275 505 -251
rect 471 -285 505 -275
rect 471 -343 505 -323
rect 471 -357 505 -343
rect 471 -411 505 -395
rect 471 -429 505 -411
rect 471 -479 505 -467
rect 471 -501 505 -479
rect 471 -547 505 -539
rect 471 -573 505 -547
rect 471 -615 505 -611
rect 471 -645 505 -615
rect 471 -717 505 -683
rect 471 -785 505 -755
rect 471 -789 505 -785
rect 471 -853 505 -827
rect 471 -861 505 -853
rect 471 -921 505 -899
rect 471 -933 505 -921
rect 471 -989 505 -971
rect 471 -1005 505 -989
rect 471 -1057 505 -1043
rect 471 -1077 505 -1057
rect 471 -1125 505 -1115
rect 471 -1149 505 -1125
rect 471 -1193 505 -1187
rect 471 -1221 505 -1193
rect 471 -1261 505 -1259
rect 471 -1293 505 -1261
rect 471 -1363 505 -1331
rect 471 -1365 505 -1363
rect 471 -1431 505 -1403
rect 471 -1437 505 -1431
rect 471 -1499 505 -1475
rect 471 -1509 505 -1499
rect 2695 99 2729 109
rect 2695 75 2729 99
rect 2695 31 2729 37
rect 2695 3 2729 31
rect 2695 -37 2729 -35
rect 2695 -69 2729 -37
rect 2695 -139 2729 -107
rect 2695 -141 2729 -139
rect 2695 -207 2729 -179
rect 2695 -213 2729 -207
rect 2695 -275 2729 -251
rect 2695 -285 2729 -275
rect 2695 -343 2729 -323
rect 2695 -357 2729 -343
rect 2695 -411 2729 -395
rect 2695 -429 2729 -411
rect 2695 -479 2729 -467
rect 2695 -501 2729 -479
rect 2695 -547 2729 -539
rect 2695 -573 2729 -547
rect 2695 -615 2729 -611
rect 2695 -645 2729 -615
rect 2695 -717 2729 -683
rect 2695 -785 2729 -755
rect 2695 -789 2729 -785
rect 2695 -853 2729 -827
rect 2695 -861 2729 -853
rect 2695 -921 2729 -899
rect 2695 -933 2729 -921
rect 2695 -989 2729 -971
rect 2695 -1005 2729 -989
rect 2695 -1057 2729 -1043
rect 2695 -1077 2729 -1057
rect 2695 -1125 2729 -1115
rect 2695 -1149 2729 -1125
rect 2695 -1193 2729 -1187
rect 2695 -1221 2729 -1193
rect 2695 -1261 2729 -1259
rect 2695 -1293 2729 -1261
rect 2695 -1363 2729 -1331
rect 2695 -1365 2729 -1363
rect 2695 -1431 2729 -1403
rect 2695 -1437 2729 -1431
rect 2695 -1499 2729 -1475
rect 2695 -1509 2729 -1499
rect 539 -1689 573 -1655
rect 611 -1689 631 -1655
rect 631 -1689 645 -1655
rect 683 -1689 699 -1655
rect 699 -1689 717 -1655
rect 755 -1689 767 -1655
rect 767 -1689 789 -1655
rect 827 -1689 835 -1655
rect 835 -1689 861 -1655
rect 899 -1689 903 -1655
rect 903 -1689 933 -1655
rect 971 -1689 1005 -1655
rect 1043 -1689 1073 -1655
rect 1073 -1689 1077 -1655
rect 1115 -1689 1141 -1655
rect 1141 -1689 1149 -1655
rect 1187 -1689 1209 -1655
rect 1209 -1689 1221 -1655
rect 1259 -1689 1277 -1655
rect 1277 -1689 1293 -1655
rect 1331 -1689 1345 -1655
rect 1345 -1689 1365 -1655
rect 1403 -1689 1413 -1655
rect 1413 -1689 1437 -1655
rect 1475 -1689 1481 -1655
rect 1481 -1689 1509 -1655
rect 1547 -1689 1549 -1655
rect 1549 -1689 1581 -1655
rect 1619 -1689 1651 -1655
rect 1651 -1689 1653 -1655
rect 1691 -1689 1719 -1655
rect 1719 -1689 1725 -1655
rect 1763 -1689 1787 -1655
rect 1787 -1689 1797 -1655
rect 1835 -1689 1855 -1655
rect 1855 -1689 1869 -1655
rect 1907 -1689 1923 -1655
rect 1923 -1689 1941 -1655
rect 1979 -1689 1991 -1655
rect 1991 -1689 2013 -1655
rect 2051 -1689 2059 -1655
rect 2059 -1689 2085 -1655
rect 2123 -1689 2127 -1655
rect 2127 -1689 2157 -1655
rect 2195 -1689 2229 -1655
rect 2267 -1689 2297 -1655
rect 2297 -1689 2301 -1655
rect 2339 -1689 2365 -1655
rect 2365 -1689 2373 -1655
rect 2411 -1689 2433 -1655
rect 2433 -1689 2445 -1655
rect 2483 -1689 2501 -1655
rect 2501 -1689 2517 -1655
rect 2555 -1689 2569 -1655
rect 2569 -1689 2589 -1655
rect 2627 -1689 2661 -1655
<< metal1 >>
rect 432 3629 2768 3668
rect 432 3595 539 3629
rect 573 3595 611 3629
rect 645 3595 683 3629
rect 717 3595 755 3629
rect 789 3595 827 3629
rect 861 3595 899 3629
rect 933 3595 971 3629
rect 1005 3595 1043 3629
rect 1077 3595 1115 3629
rect 1149 3595 1187 3629
rect 1221 3595 1259 3629
rect 1293 3595 1331 3629
rect 1365 3595 1403 3629
rect 1437 3595 1475 3629
rect 1509 3595 1547 3629
rect 1581 3595 1619 3629
rect 1653 3595 1691 3629
rect 1725 3595 1763 3629
rect 1797 3595 1835 3629
rect 1869 3595 1907 3629
rect 1941 3595 1979 3629
rect 2013 3595 2051 3629
rect 2085 3595 2123 3629
rect 2157 3595 2195 3629
rect 2229 3595 2267 3629
rect 2301 3595 2339 3629
rect 2373 3595 2411 3629
rect 2445 3595 2483 3629
rect 2517 3595 2555 3629
rect 2589 3595 2627 3629
rect 2661 3595 2768 3629
rect 432 3556 2768 3595
rect 432 3528 1154 3556
rect 432 3387 562 3528
rect 432 3353 471 3387
rect 505 3353 562 3387
rect 432 3315 562 3353
rect 432 3281 471 3315
rect 505 3284 562 3315
rect 1126 3284 1154 3528
rect 505 3281 1154 3284
rect 432 3256 1154 3281
rect 2046 3528 2768 3556
rect 2046 3284 2074 3528
rect 2638 3387 2768 3528
rect 2638 3353 2695 3387
rect 2729 3353 2768 3387
rect 2638 3315 2768 3353
rect 2638 3284 2695 3315
rect 2046 3281 2695 3284
rect 2729 3281 2768 3315
rect 2046 3256 2768 3281
rect 432 3243 544 3256
rect 432 3209 471 3243
rect 505 3209 544 3243
rect 432 3171 544 3209
rect 432 3137 471 3171
rect 505 3137 544 3171
rect 432 3099 544 3137
rect 432 3065 471 3099
rect 505 3065 544 3099
rect 2656 3243 2768 3256
rect 2656 3209 2695 3243
rect 2729 3209 2768 3243
rect 2656 3171 2768 3209
rect 2656 3137 2695 3171
rect 2729 3137 2768 3171
rect 2656 3099 2768 3137
rect 432 3027 544 3065
rect 432 2993 471 3027
rect 505 2993 544 3027
rect 432 2955 544 2993
rect 700 3046 2602 3082
rect 700 2994 756 3046
rect 808 2994 820 3046
rect 872 2994 884 3046
rect 936 2994 948 3046
rect 1000 2994 1012 3046
rect 1064 2994 1076 3046
rect 1128 2994 1140 3046
rect 1192 2994 1204 3046
rect 1256 2994 1268 3046
rect 1320 2994 1332 3046
rect 1384 2994 1396 3046
rect 1448 2994 1460 3046
rect 1512 2994 1524 3046
rect 1576 2994 1588 3046
rect 1640 2994 1652 3046
rect 1704 2994 1716 3046
rect 1768 2994 1780 3046
rect 1832 2994 1844 3046
rect 1896 2994 1908 3046
rect 1960 2994 1972 3046
rect 2024 2994 2036 3046
rect 2088 2994 2100 3046
rect 2152 2994 2164 3046
rect 2216 2994 2228 3046
rect 2280 2994 2292 3046
rect 2344 2994 2356 3046
rect 2408 2994 2420 3046
rect 2472 2994 2484 3046
rect 2536 2994 2602 3046
rect 700 2958 2602 2994
rect 2656 3065 2695 3099
rect 2729 3065 2768 3099
rect 2656 3027 2768 3065
rect 2656 2993 2695 3027
rect 2729 2993 2768 3027
rect 432 2921 471 2955
rect 505 2921 544 2955
rect 432 2883 544 2921
rect 432 2849 471 2883
rect 505 2849 544 2883
rect 432 2811 544 2849
rect 432 2777 471 2811
rect 505 2777 544 2811
rect 432 2739 544 2777
rect 432 2705 471 2739
rect 505 2705 544 2739
rect 432 2667 544 2705
rect 432 2633 471 2667
rect 505 2633 544 2667
rect 774 2694 834 2958
rect 904 2694 964 2958
rect 1282 2870 1354 2874
rect 1282 2818 1292 2870
rect 1344 2818 1354 2870
rect 1282 2814 1354 2818
rect 1800 2870 1872 2874
rect 1800 2818 1810 2870
rect 1862 2818 1872 2870
rect 1800 2814 1872 2818
rect 432 2595 544 2633
rect 432 2561 471 2595
rect 505 2561 544 2595
rect 620 2638 692 2642
rect 620 2586 630 2638
rect 682 2586 692 2638
rect 620 2582 692 2586
rect 774 2634 964 2694
rect 432 2523 544 2561
rect 432 2489 471 2523
rect 505 2489 544 2523
rect 432 2451 544 2489
rect 432 2417 471 2451
rect 505 2417 544 2451
rect 432 2379 544 2417
rect 432 2345 471 2379
rect 505 2345 544 2379
rect 432 2307 544 2345
rect 432 2273 471 2307
rect 505 2273 544 2307
rect 432 2235 544 2273
rect 432 2201 471 2235
rect 505 2201 544 2235
rect 432 2163 544 2201
rect 432 2129 471 2163
rect 505 2129 544 2163
rect 432 2091 544 2129
rect 432 2057 471 2091
rect 505 2057 544 2091
rect 432 2019 544 2057
rect 432 1985 471 2019
rect 505 1985 544 2019
rect 432 1947 544 1985
rect 432 1913 471 1947
rect 505 1913 544 1947
rect 432 1875 544 1913
rect 432 1841 471 1875
rect 505 1841 544 1875
rect 432 1803 544 1841
rect 432 1769 471 1803
rect 505 1769 544 1803
rect 432 1731 544 1769
rect 432 1697 471 1731
rect 505 1697 544 1731
rect 432 1659 544 1697
rect 432 1625 471 1659
rect 505 1625 544 1659
rect 432 1587 544 1625
rect 432 1553 471 1587
rect 505 1553 544 1587
rect 432 1515 544 1553
rect 432 1481 471 1515
rect 505 1481 544 1515
rect 432 1443 544 1481
rect 432 1409 471 1443
rect 505 1409 544 1443
rect 432 1371 544 1409
rect 432 1337 471 1371
rect 505 1337 544 1371
rect 432 1299 544 1337
rect 432 1265 471 1299
rect 505 1265 544 1299
rect 432 1227 544 1265
rect 432 1193 471 1227
rect 505 1193 544 1227
rect 432 1155 544 1193
rect 432 1121 471 1155
rect 505 1121 544 1155
rect 432 1083 544 1121
rect 432 1049 471 1083
rect 505 1049 544 1083
rect 432 1011 544 1049
rect 432 977 471 1011
rect 505 977 544 1011
rect 626 2044 686 2582
rect 774 2418 834 2634
rect 904 2506 964 2634
rect 626 1992 630 2044
rect 682 1992 686 2044
rect 626 1068 686 1992
rect 774 1852 834 2118
rect 904 1852 964 2016
rect 774 1792 964 1852
rect 1030 1804 1090 2100
rect 1160 1918 1220 2016
rect 1154 1914 1226 1918
rect 1154 1862 1164 1914
rect 1216 1862 1226 1914
rect 1154 1858 1226 1862
rect 774 1538 834 1792
rect 904 1648 964 1792
rect 1024 1800 1096 1804
rect 1024 1748 1034 1800
rect 1086 1748 1096 1800
rect 1024 1744 1096 1748
rect 626 1064 942 1068
rect 626 1012 880 1064
rect 932 1012 942 1064
rect 626 1008 942 1012
rect 432 939 544 977
rect 1028 956 1088 1260
rect 1288 1252 1348 2814
rect 1538 2758 1610 2762
rect 1538 2706 1548 2758
rect 1600 2706 1610 2758
rect 1538 2702 1610 2706
rect 1410 2638 1482 2642
rect 1410 2586 1420 2638
rect 1472 2586 1482 2638
rect 1410 2582 1482 2586
rect 1416 2506 1476 2582
rect 1544 2418 1604 2702
rect 1666 2638 1738 2642
rect 1666 2586 1676 2638
rect 1728 2586 1738 2638
rect 1666 2582 1738 2586
rect 1672 2504 1732 2582
rect 1806 2390 1866 2814
rect 2194 2682 2254 2958
rect 2322 2682 2382 2958
rect 2656 2955 2768 2993
rect 2656 2921 2695 2955
rect 2729 2921 2768 2955
rect 2656 2883 2768 2921
rect 2656 2849 2695 2883
rect 2729 2849 2768 2883
rect 2656 2811 2768 2849
rect 2656 2777 2695 2811
rect 2729 2777 2768 2811
rect 2468 2758 2540 2762
rect 2468 2706 2478 2758
rect 2530 2706 2540 2758
rect 2468 2702 2540 2706
rect 2656 2739 2768 2777
rect 2656 2705 2695 2739
rect 2729 2705 2768 2739
rect 2194 2622 2382 2682
rect 2194 2508 2254 2622
rect 1412 1914 1484 1918
rect 1412 1862 1422 1914
rect 1474 1862 1484 1914
rect 1412 1858 1484 1862
rect 1670 1914 1742 1918
rect 1670 1862 1680 1914
rect 1732 1862 1742 1914
rect 1670 1858 1742 1862
rect 1418 1650 1478 1858
rect 1542 1800 1614 1804
rect 1542 1748 1552 1800
rect 1604 1748 1614 1800
rect 1542 1744 1614 1748
rect 1548 1558 1608 1744
rect 1676 1654 1736 1858
rect 1800 1546 1860 2132
rect 1934 1918 1994 2016
rect 1928 1914 2000 1918
rect 1928 1862 1938 1914
rect 1990 1862 2000 1914
rect 1928 1858 2000 1862
rect 2064 1804 2124 2124
rect 2322 1860 2382 2622
rect 2058 1800 2130 1804
rect 2058 1748 2068 1800
rect 2120 1748 2130 1800
rect 2058 1744 2130 1748
rect 2190 1800 2382 1860
rect 2190 1650 2250 1800
rect 1160 1068 1220 1158
rect 1154 1064 1226 1068
rect 1154 1012 1164 1064
rect 1216 1012 1226 1064
rect 1154 1008 1226 1012
rect 432 905 471 939
rect 505 905 544 939
rect 432 867 544 905
rect 1022 952 1094 956
rect 1022 900 1032 952
rect 1084 900 1094 952
rect 1022 896 1094 900
rect 432 854 471 867
rect 310 833 471 854
rect 505 833 544 867
rect 310 758 544 833
rect 1544 808 1604 1254
rect 1672 1062 1732 1156
rect 1802 848 1862 1268
rect 1936 1068 1996 1160
rect 1930 1064 2002 1068
rect 1930 1012 1940 1064
rect 1992 1012 2002 1064
rect 1930 1008 2002 1012
rect 2064 956 2124 1292
rect 2188 1070 2248 1152
rect 2322 1070 2382 1800
rect 2188 1010 2382 1070
rect 2058 952 2130 956
rect 2058 900 2068 952
rect 2120 900 2130 952
rect 2058 896 2130 900
rect 1796 844 1868 848
rect 432 664 544 758
rect 1538 804 1610 808
rect 1538 752 1548 804
rect 1600 752 1610 804
rect 1796 792 1806 844
rect 1858 792 1868 844
rect 1796 788 1868 792
rect 1538 748 1610 752
rect 2188 664 2248 1010
rect 2322 664 2382 1010
rect 2474 956 2534 2702
rect 2656 2667 2768 2705
rect 2656 2633 2695 2667
rect 2729 2633 2768 2667
rect 2656 2595 2768 2633
rect 2656 2561 2695 2595
rect 2729 2561 2768 2595
rect 2656 2523 2768 2561
rect 2656 2489 2695 2523
rect 2729 2489 2768 2523
rect 2656 2451 2768 2489
rect 2656 2417 2695 2451
rect 2729 2417 2768 2451
rect 2656 2379 2768 2417
rect 2656 2345 2695 2379
rect 2729 2345 2768 2379
rect 2656 2307 2768 2345
rect 2656 2273 2695 2307
rect 2729 2273 2768 2307
rect 2656 2235 2768 2273
rect 2656 2201 2695 2235
rect 2729 2201 2768 2235
rect 2656 2163 2768 2201
rect 2656 2129 2695 2163
rect 2729 2129 2768 2163
rect 2656 2091 2768 2129
rect 2656 2057 2695 2091
rect 2729 2057 2768 2091
rect 2656 2019 2768 2057
rect 2656 1985 2695 2019
rect 2729 1985 2768 2019
rect 2656 1947 2768 1985
rect 2656 1913 2695 1947
rect 2729 1913 2768 1947
rect 2656 1875 2768 1913
rect 2656 1841 2695 1875
rect 2729 1841 2768 1875
rect 2656 1803 2768 1841
rect 2656 1769 2695 1803
rect 2729 1769 2768 1803
rect 2656 1731 2768 1769
rect 2656 1697 2695 1731
rect 2729 1697 2768 1731
rect 2656 1659 2768 1697
rect 2656 1625 2695 1659
rect 2729 1625 2768 1659
rect 2656 1587 2768 1625
rect 2656 1553 2695 1587
rect 2729 1553 2768 1587
rect 2656 1515 2768 1553
rect 2656 1481 2695 1515
rect 2729 1481 2768 1515
rect 2656 1443 2768 1481
rect 2656 1409 2695 1443
rect 2729 1409 2768 1443
rect 2656 1371 2768 1409
rect 2656 1337 2695 1371
rect 2729 1337 2768 1371
rect 2656 1299 2768 1337
rect 2656 1265 2695 1299
rect 2729 1265 2768 1299
rect 2656 1227 2768 1265
rect 2656 1193 2695 1227
rect 2729 1193 2768 1227
rect 2656 1155 2768 1193
rect 2656 1121 2695 1155
rect 2729 1121 2768 1155
rect 2656 1083 2768 1121
rect 2656 1049 2695 1083
rect 2729 1049 2768 1083
rect 2656 1011 2768 1049
rect 2656 977 2695 1011
rect 2729 977 2768 1011
rect 2468 952 2540 956
rect 2468 900 2478 952
rect 2530 900 2540 952
rect 2468 896 2540 900
rect 2656 939 2768 977
rect 2656 905 2695 939
rect 2729 905 2768 939
rect 2656 867 2768 905
rect 2656 833 2695 867
rect 2729 833 2768 867
rect 2656 664 2768 833
rect 432 625 2768 664
rect 432 591 539 625
rect 573 591 611 625
rect 645 591 683 625
rect 717 591 755 625
rect 789 591 827 625
rect 861 591 899 625
rect 933 591 971 625
rect 1005 591 1043 625
rect 1077 591 1115 625
rect 1149 591 1187 625
rect 1221 591 1259 625
rect 1293 591 1331 625
rect 1365 591 1403 625
rect 1437 591 1475 625
rect 1509 591 1547 625
rect 1581 591 1619 625
rect 1653 591 1691 625
rect 1725 591 1763 625
rect 1797 591 1835 625
rect 1869 591 1907 625
rect 1941 591 1979 625
rect 2013 591 2051 625
rect 2085 591 2123 625
rect 2157 591 2195 625
rect 2229 591 2267 625
rect 2301 591 2339 625
rect 2373 591 2411 625
rect 2445 591 2483 625
rect 2517 591 2555 625
rect 2589 591 2627 625
rect 2661 591 2768 625
rect 432 552 2768 591
rect -108 532 -48 538
rect -108 528 178 532
rect -108 476 -104 528
rect -52 519 178 528
rect -52 485 125 519
rect 159 485 178 519
rect -52 476 178 485
rect -108 472 178 476
rect 214 474 274 480
rect -108 466 -48 472
rect 208 470 280 474
rect 208 418 218 470
rect 270 418 280 470
rect 208 414 280 418
rect 214 408 274 414
rect 432 310 2768 328
rect 314 289 2768 310
rect 314 255 539 289
rect 573 255 611 289
rect 645 255 683 289
rect 717 255 755 289
rect 789 255 827 289
rect 861 255 899 289
rect 933 255 971 289
rect 1005 255 1043 289
rect 1077 255 1115 289
rect 1149 255 1187 289
rect 1221 255 1259 289
rect 1293 255 1331 289
rect 1365 255 1403 289
rect 1437 255 1475 289
rect 1509 255 1547 289
rect 1581 255 1619 289
rect 1653 255 1691 289
rect 1725 255 1763 289
rect 1797 255 1835 289
rect 1869 255 1907 289
rect 1941 255 1979 289
rect 2013 255 2051 289
rect 2085 255 2123 289
rect 2157 255 2195 289
rect 2229 255 2267 289
rect 2301 255 2339 289
rect 2373 255 2411 289
rect 2445 255 2483 289
rect 2517 255 2555 289
rect 2589 255 2627 289
rect 2661 255 2768 289
rect 314 216 2768 255
rect 314 214 544 216
rect 432 109 544 214
rect 432 75 471 109
rect 505 75 544 109
rect 1544 164 1604 174
rect 1544 112 1548 164
rect 1600 112 1604 164
rect 432 37 544 75
rect 1022 98 1094 102
rect 1022 46 1032 98
rect 1084 46 1094 98
rect 1022 42 1094 46
rect 1276 54 1348 58
rect 432 3 471 37
rect 505 3 544 37
rect 432 -35 544 3
rect 432 -69 471 -35
rect 505 -69 544 -35
rect 432 -107 544 -69
rect 432 -141 471 -107
rect 505 -141 544 -107
rect 432 -179 544 -141
rect 432 -213 471 -179
rect 505 -213 544 -179
rect 432 -251 544 -213
rect 432 -285 471 -251
rect 505 -285 544 -251
rect 432 -323 544 -285
rect 1028 -312 1088 42
rect 1276 2 1286 54
rect 1338 2 1348 54
rect 1276 -2 1348 2
rect 1282 -278 1342 -2
rect 1408 -58 1480 -54
rect 1408 -110 1418 -58
rect 1470 -110 1480 -58
rect 1408 -114 1480 -110
rect 1414 -194 1474 -114
rect 1544 -274 1604 112
rect 2656 109 2768 216
rect 2656 75 2695 109
rect 2729 75 2768 109
rect 1796 54 1868 58
rect 1796 2 1806 54
rect 1858 2 1868 54
rect 1796 -2 1868 2
rect 2656 37 2768 75
rect 2656 3 2695 37
rect 2729 3 2768 37
rect 1664 -58 1736 -54
rect 1664 -110 1674 -58
rect 1726 -110 1736 -58
rect 1664 -114 1736 -110
rect 1670 -192 1730 -114
rect 1802 -284 1862 -2
rect 2656 -35 2768 3
rect 2656 -69 2695 -35
rect 2729 -69 2768 -35
rect 2656 -107 2768 -69
rect 2656 -141 2695 -107
rect 2729 -141 2768 -107
rect 2656 -179 2768 -141
rect 2656 -213 2695 -179
rect 2729 -213 2768 -179
rect 2656 -251 2768 -213
rect 2656 -285 2695 -251
rect 2729 -285 2768 -251
rect 432 -357 471 -323
rect 505 -357 544 -323
rect 432 -395 544 -357
rect 432 -429 471 -395
rect 505 -429 544 -395
rect 432 -467 544 -429
rect 432 -501 471 -467
rect 505 -501 544 -467
rect 432 -539 544 -501
rect 432 -573 471 -539
rect 505 -573 544 -539
rect 2656 -323 2768 -285
rect 2656 -357 2695 -323
rect 2729 -357 2768 -323
rect 2656 -395 2768 -357
rect 2656 -429 2695 -395
rect 2729 -429 2768 -395
rect 2656 -467 2768 -429
rect 2656 -501 2695 -467
rect 2729 -501 2768 -467
rect 2656 -539 2768 -501
rect 432 -611 544 -573
rect 432 -645 471 -611
rect 505 -645 544 -611
rect 432 -683 544 -645
rect 432 -717 471 -683
rect 505 -717 544 -683
rect 432 -755 544 -717
rect 432 -789 471 -755
rect 505 -789 544 -755
rect 432 -827 544 -789
rect 432 -861 471 -827
rect 505 -861 544 -827
rect 432 -899 544 -861
rect 432 -933 471 -899
rect 505 -933 544 -899
rect 432 -971 544 -933
rect 432 -1005 471 -971
rect 505 -1005 544 -971
rect 432 -1043 544 -1005
rect 766 -738 826 -564
rect 896 -738 956 -668
rect 766 -798 956 -738
rect 766 -1034 826 -798
rect 896 -1034 956 -798
rect 1022 -864 1082 -582
rect 1156 -750 1216 -666
rect 1930 -750 1990 -666
rect 1150 -754 1222 -750
rect 1150 -806 1160 -754
rect 1212 -806 1222 -754
rect 1150 -810 1222 -806
rect 1924 -754 1996 -750
rect 1924 -806 1934 -754
rect 1986 -806 1996 -754
rect 1924 -810 1996 -806
rect 2058 -864 2118 -564
rect 2186 -744 2246 -668
rect 2314 -744 2374 -572
rect 2186 -804 2374 -744
rect 1016 -868 1088 -864
rect 1016 -920 1026 -868
rect 1078 -920 1088 -868
rect 1016 -924 1088 -920
rect 2052 -868 2124 -864
rect 2052 -920 2062 -868
rect 2114 -920 2124 -868
rect 2052 -924 2124 -920
rect 2186 -1034 2246 -804
rect 2314 -1034 2374 -804
rect 2656 -573 2695 -539
rect 2729 -573 2768 -539
rect 2656 -611 2768 -573
rect 2656 -645 2695 -611
rect 2729 -645 2768 -611
rect 2656 -683 2768 -645
rect 2656 -717 2695 -683
rect 2729 -717 2768 -683
rect 2656 -755 2768 -717
rect 2656 -789 2695 -755
rect 2729 -789 2768 -755
rect 2656 -827 2768 -789
rect 2656 -861 2695 -827
rect 2729 -861 2768 -827
rect 2656 -899 2768 -861
rect 2656 -933 2695 -899
rect 2729 -933 2768 -899
rect 2656 -971 2768 -933
rect 2656 -1005 2695 -971
rect 2729 -1005 2768 -971
rect 432 -1077 471 -1043
rect 505 -1077 544 -1043
rect 432 -1115 544 -1077
rect 432 -1149 471 -1115
rect 505 -1149 544 -1115
rect 432 -1187 544 -1149
rect 656 -1074 2434 -1034
rect 656 -1126 720 -1074
rect 772 -1126 784 -1074
rect 836 -1126 848 -1074
rect 900 -1126 912 -1074
rect 964 -1126 976 -1074
rect 1028 -1126 1040 -1074
rect 1092 -1126 1104 -1074
rect 1156 -1126 1168 -1074
rect 1220 -1126 1232 -1074
rect 1284 -1126 1296 -1074
rect 1348 -1126 1360 -1074
rect 1412 -1126 1424 -1074
rect 1476 -1126 1488 -1074
rect 1540 -1126 1552 -1074
rect 1604 -1126 1616 -1074
rect 1668 -1126 1680 -1074
rect 1732 -1126 1744 -1074
rect 1796 -1126 1808 -1074
rect 1860 -1126 1872 -1074
rect 1924 -1126 1936 -1074
rect 1988 -1126 2000 -1074
rect 2052 -1126 2064 -1074
rect 2116 -1126 2128 -1074
rect 2180 -1126 2192 -1074
rect 2244 -1126 2256 -1074
rect 2308 -1126 2320 -1074
rect 2372 -1126 2434 -1074
rect 656 -1164 2434 -1126
rect 2656 -1043 2768 -1005
rect 2656 -1077 2695 -1043
rect 2729 -1077 2768 -1043
rect 2656 -1115 2768 -1077
rect 2656 -1149 2695 -1115
rect 2729 -1149 2768 -1115
rect 432 -1221 471 -1187
rect 505 -1221 544 -1187
rect 432 -1259 544 -1221
rect 432 -1293 471 -1259
rect 505 -1293 544 -1259
rect 432 -1316 544 -1293
rect 2656 -1187 2768 -1149
rect 2656 -1221 2695 -1187
rect 2729 -1221 2768 -1187
rect 2656 -1259 2768 -1221
rect 2656 -1293 2695 -1259
rect 2729 -1293 2768 -1259
rect 2656 -1316 2768 -1293
rect 432 -1331 1154 -1316
rect 432 -1365 471 -1331
rect 505 -1344 1154 -1331
rect 505 -1365 562 -1344
rect 432 -1403 562 -1365
rect 432 -1437 471 -1403
rect 505 -1437 562 -1403
rect 432 -1475 562 -1437
rect 432 -1509 471 -1475
rect 505 -1509 562 -1475
rect 432 -1588 562 -1509
rect 1126 -1588 1154 -1344
rect 432 -1616 1154 -1588
rect 2046 -1331 2768 -1316
rect 2046 -1344 2695 -1331
rect 2046 -1588 2074 -1344
rect 2638 -1365 2695 -1344
rect 2729 -1365 2768 -1331
rect 2638 -1403 2768 -1365
rect 2638 -1437 2695 -1403
rect 2729 -1437 2768 -1403
rect 2638 -1475 2768 -1437
rect 2638 -1509 2695 -1475
rect 2729 -1509 2768 -1475
rect 2638 -1588 2768 -1509
rect 2046 -1616 2768 -1588
rect 432 -1655 2768 -1616
rect 432 -1689 539 -1655
rect 573 -1689 611 -1655
rect 645 -1689 683 -1655
rect 717 -1689 755 -1655
rect 789 -1689 827 -1655
rect 861 -1689 899 -1655
rect 933 -1689 971 -1655
rect 1005 -1689 1043 -1655
rect 1077 -1689 1115 -1655
rect 1149 -1689 1187 -1655
rect 1221 -1689 1259 -1655
rect 1293 -1689 1331 -1655
rect 1365 -1689 1403 -1655
rect 1437 -1689 1475 -1655
rect 1509 -1689 1547 -1655
rect 1581 -1689 1619 -1655
rect 1653 -1689 1691 -1655
rect 1725 -1689 1763 -1655
rect 1797 -1689 1835 -1655
rect 1869 -1689 1907 -1655
rect 1941 -1689 1979 -1655
rect 2013 -1689 2051 -1655
rect 2085 -1689 2123 -1655
rect 2157 -1689 2195 -1655
rect 2229 -1689 2267 -1655
rect 2301 -1689 2339 -1655
rect 2373 -1689 2411 -1655
rect 2445 -1689 2483 -1655
rect 2517 -1689 2555 -1655
rect 2589 -1689 2627 -1655
rect 2661 -1689 2768 -1655
rect 432 -1728 2768 -1689
<< via1 >>
rect 562 3284 1126 3528
rect 2074 3284 2638 3528
rect 756 2994 808 3046
rect 820 2994 872 3046
rect 884 2994 936 3046
rect 948 2994 1000 3046
rect 1012 2994 1064 3046
rect 1076 2994 1128 3046
rect 1140 2994 1192 3046
rect 1204 2994 1256 3046
rect 1268 2994 1320 3046
rect 1332 2994 1384 3046
rect 1396 2994 1448 3046
rect 1460 2994 1512 3046
rect 1524 2994 1576 3046
rect 1588 2994 1640 3046
rect 1652 2994 1704 3046
rect 1716 2994 1768 3046
rect 1780 2994 1832 3046
rect 1844 2994 1896 3046
rect 1908 2994 1960 3046
rect 1972 2994 2024 3046
rect 2036 2994 2088 3046
rect 2100 2994 2152 3046
rect 2164 2994 2216 3046
rect 2228 2994 2280 3046
rect 2292 2994 2344 3046
rect 2356 2994 2408 3046
rect 2420 2994 2472 3046
rect 2484 2994 2536 3046
rect 1292 2818 1344 2870
rect 1810 2818 1862 2870
rect 630 2586 682 2638
rect 630 1992 682 2044
rect 1164 1862 1216 1914
rect 1034 1748 1086 1800
rect 880 1012 932 1064
rect 1548 2706 1600 2758
rect 1420 2586 1472 2638
rect 1676 2586 1728 2638
rect 2478 2706 2530 2758
rect 1422 1862 1474 1914
rect 1680 1862 1732 1914
rect 1552 1748 1604 1800
rect 1938 1862 1990 1914
rect 2068 1748 2120 1800
rect 1164 1012 1216 1064
rect 1032 900 1084 952
rect 1940 1012 1992 1064
rect 2068 900 2120 952
rect 1548 752 1600 804
rect 1806 792 1858 844
rect 2478 900 2530 952
rect -104 476 -52 528
rect 218 461 270 470
rect 218 427 227 461
rect 227 427 261 461
rect 261 427 270 461
rect 218 418 270 427
rect 1548 112 1600 164
rect 1032 46 1084 98
rect 1286 2 1338 54
rect 1418 -110 1470 -58
rect 1806 2 1858 54
rect 1674 -110 1726 -58
rect 1160 -806 1212 -754
rect 1934 -806 1986 -754
rect 1026 -920 1078 -868
rect 2062 -920 2114 -868
rect 720 -1126 772 -1074
rect 784 -1126 836 -1074
rect 848 -1126 900 -1074
rect 912 -1126 964 -1074
rect 976 -1126 1028 -1074
rect 1040 -1126 1092 -1074
rect 1104 -1126 1156 -1074
rect 1168 -1126 1220 -1074
rect 1232 -1126 1284 -1074
rect 1296 -1126 1348 -1074
rect 1360 -1126 1412 -1074
rect 1424 -1126 1476 -1074
rect 1488 -1126 1540 -1074
rect 1552 -1126 1604 -1074
rect 1616 -1126 1668 -1074
rect 1680 -1126 1732 -1074
rect 1744 -1126 1796 -1074
rect 1808 -1126 1860 -1074
rect 1872 -1126 1924 -1074
rect 1936 -1126 1988 -1074
rect 2000 -1126 2052 -1074
rect 2064 -1126 2116 -1074
rect 2128 -1126 2180 -1074
rect 2192 -1126 2244 -1074
rect 2256 -1126 2308 -1074
rect 2320 -1126 2372 -1074
rect 562 -1588 1126 -1344
rect 2074 -1588 2638 -1344
<< metal2 >>
rect 544 3554 1144 3566
rect 544 3528 576 3554
rect 1112 3528 1144 3554
rect 544 3284 562 3528
rect 1126 3284 1144 3528
rect 544 3258 576 3284
rect 1112 3258 1144 3284
rect 544 3246 1144 3258
rect 2056 3554 2656 3566
rect 2056 3528 2088 3554
rect 2624 3528 2656 3554
rect 2056 3284 2074 3528
rect 2638 3284 2656 3528
rect 2056 3258 2088 3284
rect 2624 3258 2656 3284
rect 2056 3246 2656 3258
rect 700 3048 2602 3082
rect 700 2992 738 3048
rect 794 3046 818 3048
rect 874 3046 898 3048
rect 954 3046 978 3048
rect 1034 3046 1058 3048
rect 1114 3046 1138 3048
rect 1194 3046 1218 3048
rect 1274 3046 1298 3048
rect 1354 3046 1378 3048
rect 1434 3046 1458 3048
rect 1514 3046 1538 3048
rect 1594 3046 1618 3048
rect 1674 3046 1698 3048
rect 1754 3046 1778 3048
rect 1834 3046 1858 3048
rect 1914 3046 1938 3048
rect 1994 3046 2018 3048
rect 2074 3046 2098 3048
rect 2154 3046 2178 3048
rect 2234 3046 2258 3048
rect 2314 3046 2338 3048
rect 2394 3046 2418 3048
rect 2474 3046 2498 3048
rect 808 2994 818 3046
rect 874 2994 884 3046
rect 1128 2994 1138 3046
rect 1194 2994 1204 3046
rect 1448 2994 1458 3046
rect 1514 2994 1524 3046
rect 1768 2994 1778 3046
rect 1834 2994 1844 3046
rect 2088 2994 2098 3046
rect 2154 2994 2164 3046
rect 2408 2994 2418 3046
rect 2474 2994 2484 3046
rect 794 2992 818 2994
rect 874 2992 898 2994
rect 954 2992 978 2994
rect 1034 2992 1058 2994
rect 1114 2992 1138 2994
rect 1194 2992 1218 2994
rect 1274 2992 1298 2994
rect 1354 2992 1378 2994
rect 1434 2992 1458 2994
rect 1514 2992 1538 2994
rect 1594 2992 1618 2994
rect 1674 2992 1698 2994
rect 1754 2992 1778 2994
rect 1834 2992 1858 2994
rect 1914 2992 1938 2994
rect 1994 2992 2018 2994
rect 2074 2992 2098 2994
rect 2154 2992 2178 2994
rect 2234 2992 2258 2994
rect 2314 2992 2338 2994
rect 2394 2992 2418 2994
rect 2474 2992 2498 2994
rect 2554 2992 2602 3048
rect 700 2958 2602 2992
rect 1288 2874 1348 2880
rect 1806 2874 1866 2880
rect 1288 2870 1866 2874
rect 1288 2818 1292 2870
rect 1344 2818 1810 2870
rect 1862 2818 1866 2870
rect 1288 2814 1866 2818
rect 1288 2808 1348 2814
rect 1806 2808 1866 2814
rect 1544 2762 1604 2768
rect 2474 2762 2534 2768
rect 1544 2758 2534 2762
rect 1544 2706 1548 2758
rect 1600 2706 2478 2758
rect 2530 2706 2534 2758
rect 1544 2702 2534 2706
rect 1544 2696 1604 2702
rect 2474 2696 2534 2702
rect 626 2642 686 2648
rect 1416 2642 1476 2648
rect 1672 2642 1732 2648
rect 626 2638 1732 2642
rect 626 2586 630 2638
rect 682 2586 1420 2638
rect 1472 2586 1676 2638
rect 1728 2586 1732 2638
rect 626 2582 1732 2586
rect 626 2576 686 2582
rect 1416 2576 1476 2582
rect 1672 2576 1732 2582
rect -108 2044 692 2048
rect -108 1992 630 2044
rect 682 1992 692 2044
rect -108 1988 692 1992
rect -108 532 -48 1988
rect 1160 1918 1220 1924
rect 1418 1918 1478 1924
rect 1676 1918 1736 1924
rect 1934 1918 1994 1924
rect 628 1914 1994 1918
rect 628 1862 1164 1914
rect 1216 1862 1422 1914
rect 1474 1862 1680 1914
rect 1732 1862 1938 1914
rect 1990 1862 1994 1914
rect 628 1858 1994 1862
rect -114 528 -42 532
rect -114 476 -104 528
rect -52 476 -42 528
rect -114 472 -42 476
rect 628 474 688 1858
rect 1160 1852 1220 1858
rect 1418 1852 1478 1858
rect 1676 1852 1736 1858
rect 1934 1852 1994 1858
rect 1030 1804 1090 1810
rect 1548 1804 1608 1810
rect 2064 1804 2124 1810
rect 1030 1800 2124 1804
rect 1030 1748 1034 1800
rect 1086 1748 1552 1800
rect 1604 1748 2068 1800
rect 2120 1748 2124 1800
rect 1030 1744 2124 1748
rect 1030 1738 1090 1744
rect 1548 1738 1608 1744
rect 2064 1738 2124 1744
rect 208 470 688 474
rect 208 418 218 470
rect 270 418 688 470
rect 208 414 688 418
rect 628 -750 688 414
rect 876 1068 936 1074
rect 1160 1068 1220 1074
rect 1936 1068 1996 1074
rect 876 1064 1996 1068
rect 876 1012 880 1064
rect 932 1012 1164 1064
rect 1216 1012 1940 1064
rect 1992 1012 1996 1064
rect 876 1008 1996 1012
rect 876 -54 936 1008
rect 1160 1002 1220 1008
rect 1936 1002 1996 1008
rect 1028 956 1088 962
rect 2064 956 2124 962
rect 2474 956 2534 962
rect 1028 952 2534 956
rect 1028 900 1032 952
rect 1084 900 2068 952
rect 2120 900 2478 952
rect 2530 900 2534 952
rect 1028 896 2534 900
rect 1028 98 1088 896
rect 2064 890 2124 896
rect 2474 890 2534 896
rect 1802 844 1862 854
rect 1544 804 1604 814
rect 1544 752 1548 804
rect 1600 752 1604 804
rect 1544 168 1604 752
rect 1802 792 1806 844
rect 1858 792 1862 844
rect 1538 164 1610 168
rect 1538 112 1548 164
rect 1600 112 1610 164
rect 1538 108 1610 112
rect 1028 46 1032 98
rect 1084 46 1088 98
rect 1028 36 1088 46
rect 1282 58 1342 64
rect 1802 58 1862 792
rect 1282 54 1862 58
rect 1282 2 1286 54
rect 1338 2 1806 54
rect 1858 2 1862 54
rect 1282 -2 1862 2
rect 1282 -8 1342 -2
rect 1802 -8 1862 -2
rect 1414 -54 1474 -48
rect 1670 -54 1730 -48
rect 876 -58 1730 -54
rect 876 -110 1418 -58
rect 1470 -110 1674 -58
rect 1726 -110 1730 -58
rect 876 -114 1730 -110
rect 1414 -120 1474 -114
rect 1670 -120 1730 -114
rect 1156 -750 1216 -744
rect 1930 -750 1990 -744
rect 628 -754 1990 -750
rect 628 -806 1160 -754
rect 1212 -806 1934 -754
rect 1986 -806 1990 -754
rect 628 -810 1990 -806
rect 1156 -816 1216 -810
rect 1930 -816 1990 -810
rect 1022 -864 1082 -858
rect 2058 -864 2118 -858
rect 1022 -868 2118 -864
rect 1022 -920 1026 -868
rect 1078 -920 2062 -868
rect 2114 -920 2118 -868
rect 1022 -924 2118 -920
rect 1022 -930 1082 -924
rect 2058 -930 2118 -924
rect 656 -1072 2434 -1034
rect 656 -1128 718 -1072
rect 774 -1074 798 -1072
rect 854 -1074 878 -1072
rect 934 -1074 958 -1072
rect 1014 -1074 1038 -1072
rect 1094 -1074 1118 -1072
rect 1174 -1074 1198 -1072
rect 1254 -1074 1278 -1072
rect 1334 -1074 1358 -1072
rect 1414 -1074 1438 -1072
rect 1494 -1074 1518 -1072
rect 1574 -1074 1598 -1072
rect 1654 -1074 1678 -1072
rect 1734 -1074 1758 -1072
rect 1814 -1074 1838 -1072
rect 1894 -1074 1918 -1072
rect 1974 -1074 1998 -1072
rect 2054 -1074 2078 -1072
rect 2134 -1074 2158 -1072
rect 2214 -1074 2238 -1072
rect 2294 -1074 2318 -1072
rect 774 -1126 784 -1074
rect 1028 -1126 1038 -1074
rect 1094 -1126 1104 -1074
rect 1348 -1126 1358 -1074
rect 1414 -1126 1424 -1074
rect 1668 -1126 1678 -1074
rect 1734 -1126 1744 -1074
rect 1988 -1126 1998 -1074
rect 2054 -1126 2064 -1074
rect 2308 -1126 2318 -1074
rect 774 -1128 798 -1126
rect 854 -1128 878 -1126
rect 934 -1128 958 -1126
rect 1014 -1128 1038 -1126
rect 1094 -1128 1118 -1126
rect 1174 -1128 1198 -1126
rect 1254 -1128 1278 -1126
rect 1334 -1128 1358 -1126
rect 1414 -1128 1438 -1126
rect 1494 -1128 1518 -1126
rect 1574 -1128 1598 -1126
rect 1654 -1128 1678 -1126
rect 1734 -1128 1758 -1126
rect 1814 -1128 1838 -1126
rect 1894 -1128 1918 -1126
rect 1974 -1128 1998 -1126
rect 2054 -1128 2078 -1126
rect 2134 -1128 2158 -1126
rect 2214 -1128 2238 -1126
rect 2294 -1128 2318 -1126
rect 2374 -1128 2434 -1072
rect 656 -1164 2434 -1128
rect 544 -1318 1144 -1306
rect 544 -1344 576 -1318
rect 1112 -1344 1144 -1318
rect 544 -1588 562 -1344
rect 1126 -1588 1144 -1344
rect 544 -1614 576 -1588
rect 1112 -1614 1144 -1588
rect 544 -1626 1144 -1614
rect 2056 -1318 2656 -1306
rect 2056 -1344 2088 -1318
rect 2624 -1344 2656 -1318
rect 2056 -1588 2074 -1344
rect 2638 -1588 2656 -1344
rect 2056 -1614 2088 -1588
rect 2624 -1614 2656 -1588
rect 2056 -1626 2656 -1614
<< via2 >>
rect 576 3528 1112 3554
rect 576 3284 1112 3528
rect 576 3258 1112 3284
rect 2088 3528 2624 3554
rect 2088 3284 2624 3528
rect 2088 3258 2624 3284
rect 738 3046 794 3048
rect 818 3046 874 3048
rect 898 3046 954 3048
rect 978 3046 1034 3048
rect 1058 3046 1114 3048
rect 1138 3046 1194 3048
rect 1218 3046 1274 3048
rect 1298 3046 1354 3048
rect 1378 3046 1434 3048
rect 1458 3046 1514 3048
rect 1538 3046 1594 3048
rect 1618 3046 1674 3048
rect 1698 3046 1754 3048
rect 1778 3046 1834 3048
rect 1858 3046 1914 3048
rect 1938 3046 1994 3048
rect 2018 3046 2074 3048
rect 2098 3046 2154 3048
rect 2178 3046 2234 3048
rect 2258 3046 2314 3048
rect 2338 3046 2394 3048
rect 2418 3046 2474 3048
rect 2498 3046 2554 3048
rect 738 2994 756 3046
rect 756 2994 794 3046
rect 818 2994 820 3046
rect 820 2994 872 3046
rect 872 2994 874 3046
rect 898 2994 936 3046
rect 936 2994 948 3046
rect 948 2994 954 3046
rect 978 2994 1000 3046
rect 1000 2994 1012 3046
rect 1012 2994 1034 3046
rect 1058 2994 1064 3046
rect 1064 2994 1076 3046
rect 1076 2994 1114 3046
rect 1138 2994 1140 3046
rect 1140 2994 1192 3046
rect 1192 2994 1194 3046
rect 1218 2994 1256 3046
rect 1256 2994 1268 3046
rect 1268 2994 1274 3046
rect 1298 2994 1320 3046
rect 1320 2994 1332 3046
rect 1332 2994 1354 3046
rect 1378 2994 1384 3046
rect 1384 2994 1396 3046
rect 1396 2994 1434 3046
rect 1458 2994 1460 3046
rect 1460 2994 1512 3046
rect 1512 2994 1514 3046
rect 1538 2994 1576 3046
rect 1576 2994 1588 3046
rect 1588 2994 1594 3046
rect 1618 2994 1640 3046
rect 1640 2994 1652 3046
rect 1652 2994 1674 3046
rect 1698 2994 1704 3046
rect 1704 2994 1716 3046
rect 1716 2994 1754 3046
rect 1778 2994 1780 3046
rect 1780 2994 1832 3046
rect 1832 2994 1834 3046
rect 1858 2994 1896 3046
rect 1896 2994 1908 3046
rect 1908 2994 1914 3046
rect 1938 2994 1960 3046
rect 1960 2994 1972 3046
rect 1972 2994 1994 3046
rect 2018 2994 2024 3046
rect 2024 2994 2036 3046
rect 2036 2994 2074 3046
rect 2098 2994 2100 3046
rect 2100 2994 2152 3046
rect 2152 2994 2154 3046
rect 2178 2994 2216 3046
rect 2216 2994 2228 3046
rect 2228 2994 2234 3046
rect 2258 2994 2280 3046
rect 2280 2994 2292 3046
rect 2292 2994 2314 3046
rect 2338 2994 2344 3046
rect 2344 2994 2356 3046
rect 2356 2994 2394 3046
rect 2418 2994 2420 3046
rect 2420 2994 2472 3046
rect 2472 2994 2474 3046
rect 2498 2994 2536 3046
rect 2536 2994 2554 3046
rect 738 2992 794 2994
rect 818 2992 874 2994
rect 898 2992 954 2994
rect 978 2992 1034 2994
rect 1058 2992 1114 2994
rect 1138 2992 1194 2994
rect 1218 2992 1274 2994
rect 1298 2992 1354 2994
rect 1378 2992 1434 2994
rect 1458 2992 1514 2994
rect 1538 2992 1594 2994
rect 1618 2992 1674 2994
rect 1698 2992 1754 2994
rect 1778 2992 1834 2994
rect 1858 2992 1914 2994
rect 1938 2992 1994 2994
rect 2018 2992 2074 2994
rect 2098 2992 2154 2994
rect 2178 2992 2234 2994
rect 2258 2992 2314 2994
rect 2338 2992 2394 2994
rect 2418 2992 2474 2994
rect 2498 2992 2554 2994
rect 718 -1074 774 -1072
rect 798 -1074 854 -1072
rect 878 -1074 934 -1072
rect 958 -1074 1014 -1072
rect 1038 -1074 1094 -1072
rect 1118 -1074 1174 -1072
rect 1198 -1074 1254 -1072
rect 1278 -1074 1334 -1072
rect 1358 -1074 1414 -1072
rect 1438 -1074 1494 -1072
rect 1518 -1074 1574 -1072
rect 1598 -1074 1654 -1072
rect 1678 -1074 1734 -1072
rect 1758 -1074 1814 -1072
rect 1838 -1074 1894 -1072
rect 1918 -1074 1974 -1072
rect 1998 -1074 2054 -1072
rect 2078 -1074 2134 -1072
rect 2158 -1074 2214 -1072
rect 2238 -1074 2294 -1072
rect 2318 -1074 2374 -1072
rect 718 -1126 720 -1074
rect 720 -1126 772 -1074
rect 772 -1126 774 -1074
rect 798 -1126 836 -1074
rect 836 -1126 848 -1074
rect 848 -1126 854 -1074
rect 878 -1126 900 -1074
rect 900 -1126 912 -1074
rect 912 -1126 934 -1074
rect 958 -1126 964 -1074
rect 964 -1126 976 -1074
rect 976 -1126 1014 -1074
rect 1038 -1126 1040 -1074
rect 1040 -1126 1092 -1074
rect 1092 -1126 1094 -1074
rect 1118 -1126 1156 -1074
rect 1156 -1126 1168 -1074
rect 1168 -1126 1174 -1074
rect 1198 -1126 1220 -1074
rect 1220 -1126 1232 -1074
rect 1232 -1126 1254 -1074
rect 1278 -1126 1284 -1074
rect 1284 -1126 1296 -1074
rect 1296 -1126 1334 -1074
rect 1358 -1126 1360 -1074
rect 1360 -1126 1412 -1074
rect 1412 -1126 1414 -1074
rect 1438 -1126 1476 -1074
rect 1476 -1126 1488 -1074
rect 1488 -1126 1494 -1074
rect 1518 -1126 1540 -1074
rect 1540 -1126 1552 -1074
rect 1552 -1126 1574 -1074
rect 1598 -1126 1604 -1074
rect 1604 -1126 1616 -1074
rect 1616 -1126 1654 -1074
rect 1678 -1126 1680 -1074
rect 1680 -1126 1732 -1074
rect 1732 -1126 1734 -1074
rect 1758 -1126 1796 -1074
rect 1796 -1126 1808 -1074
rect 1808 -1126 1814 -1074
rect 1838 -1126 1860 -1074
rect 1860 -1126 1872 -1074
rect 1872 -1126 1894 -1074
rect 1918 -1126 1924 -1074
rect 1924 -1126 1936 -1074
rect 1936 -1126 1974 -1074
rect 1998 -1126 2000 -1074
rect 2000 -1126 2052 -1074
rect 2052 -1126 2054 -1074
rect 2078 -1126 2116 -1074
rect 2116 -1126 2128 -1074
rect 2128 -1126 2134 -1074
rect 2158 -1126 2180 -1074
rect 2180 -1126 2192 -1074
rect 2192 -1126 2214 -1074
rect 2238 -1126 2244 -1074
rect 2244 -1126 2256 -1074
rect 2256 -1126 2294 -1074
rect 2318 -1126 2320 -1074
rect 2320 -1126 2372 -1074
rect 2372 -1126 2374 -1074
rect 718 -1128 774 -1126
rect 798 -1128 854 -1126
rect 878 -1128 934 -1126
rect 958 -1128 1014 -1126
rect 1038 -1128 1094 -1126
rect 1118 -1128 1174 -1126
rect 1198 -1128 1254 -1126
rect 1278 -1128 1334 -1126
rect 1358 -1128 1414 -1126
rect 1438 -1128 1494 -1126
rect 1518 -1128 1574 -1126
rect 1598 -1128 1654 -1126
rect 1678 -1128 1734 -1126
rect 1758 -1128 1814 -1126
rect 1838 -1128 1894 -1126
rect 1918 -1128 1974 -1126
rect 1998 -1128 2054 -1126
rect 2078 -1128 2134 -1126
rect 2158 -1128 2214 -1126
rect 2238 -1128 2294 -1126
rect 2318 -1128 2374 -1126
rect 576 -1344 1112 -1318
rect 576 -1588 1112 -1344
rect 576 -1614 1112 -1588
rect 2088 -1344 2624 -1318
rect 2088 -1588 2624 -1344
rect 2088 -1614 2624 -1588
<< metal3 >>
rect 534 3554 1154 3561
rect 534 3518 576 3554
rect 1112 3518 1154 3554
rect 534 3294 572 3518
rect 1116 3294 1154 3518
rect 534 3258 576 3294
rect 1112 3258 1154 3294
rect 534 3251 1154 3258
rect 2046 3554 2666 3561
rect 2046 3518 2088 3554
rect 2624 3518 2666 3554
rect 2046 3294 2084 3518
rect 2628 3294 2666 3518
rect 2046 3258 2088 3294
rect 2624 3258 2666 3294
rect 2046 3251 2666 3258
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 798 2988 814 3052
rect 878 2988 894 3052
rect 958 2988 974 3052
rect 1038 2988 1054 3052
rect 1118 2988 1134 3052
rect 1198 2988 1214 3052
rect 1278 2988 1294 3052
rect 1358 2988 1374 3052
rect 1438 2988 1454 3052
rect 1518 2988 1534 3052
rect 1598 2988 1614 3052
rect 1678 2988 1694 3052
rect 1758 2988 1774 3052
rect 1838 2988 1854 3052
rect 1918 2988 1934 3052
rect 1998 2988 2014 3052
rect 2078 2988 2094 3052
rect 2158 2988 2174 3052
rect 2238 2988 2254 3052
rect 2318 2988 2334 3052
rect 2398 2988 2414 3052
rect 2478 2988 2494 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 656 -1068 2434 -1034
rect 656 -1132 714 -1068
rect 778 -1132 794 -1068
rect 858 -1132 874 -1068
rect 938 -1132 954 -1068
rect 1018 -1132 1034 -1068
rect 1098 -1132 1114 -1068
rect 1178 -1132 1194 -1068
rect 1258 -1132 1274 -1068
rect 1338 -1132 1354 -1068
rect 1418 -1132 1434 -1068
rect 1498 -1132 1514 -1068
rect 1578 -1132 1594 -1068
rect 1658 -1132 1674 -1068
rect 1738 -1132 1754 -1068
rect 1818 -1132 1834 -1068
rect 1898 -1132 1914 -1068
rect 1978 -1132 1994 -1068
rect 2058 -1132 2074 -1068
rect 2138 -1132 2154 -1068
rect 2218 -1132 2234 -1068
rect 2298 -1132 2314 -1068
rect 2378 -1132 2434 -1068
rect 656 -1164 2434 -1132
rect 534 -1318 1154 -1311
rect 534 -1354 576 -1318
rect 1112 -1354 1154 -1318
rect 534 -1578 572 -1354
rect 1116 -1578 1154 -1354
rect 534 -1614 576 -1578
rect 1112 -1614 1154 -1578
rect 534 -1621 1154 -1614
rect 2046 -1318 2666 -1311
rect 2046 -1354 2088 -1318
rect 2624 -1354 2666 -1318
rect 2046 -1578 2084 -1354
rect 2628 -1578 2666 -1354
rect 2046 -1614 2088 -1578
rect 2624 -1614 2666 -1578
rect 2046 -1621 2666 -1614
<< via3 >>
rect 572 3294 576 3518
rect 576 3294 1112 3518
rect 1112 3294 1116 3518
rect 2084 3294 2088 3518
rect 2088 3294 2624 3518
rect 2624 3294 2628 3518
rect 734 3048 798 3052
rect 734 2992 738 3048
rect 738 2992 794 3048
rect 794 2992 798 3048
rect 734 2988 798 2992
rect 814 3048 878 3052
rect 814 2992 818 3048
rect 818 2992 874 3048
rect 874 2992 878 3048
rect 814 2988 878 2992
rect 894 3048 958 3052
rect 894 2992 898 3048
rect 898 2992 954 3048
rect 954 2992 958 3048
rect 894 2988 958 2992
rect 974 3048 1038 3052
rect 974 2992 978 3048
rect 978 2992 1034 3048
rect 1034 2992 1038 3048
rect 974 2988 1038 2992
rect 1054 3048 1118 3052
rect 1054 2992 1058 3048
rect 1058 2992 1114 3048
rect 1114 2992 1118 3048
rect 1054 2988 1118 2992
rect 1134 3048 1198 3052
rect 1134 2992 1138 3048
rect 1138 2992 1194 3048
rect 1194 2992 1198 3048
rect 1134 2988 1198 2992
rect 1214 3048 1278 3052
rect 1214 2992 1218 3048
rect 1218 2992 1274 3048
rect 1274 2992 1278 3048
rect 1214 2988 1278 2992
rect 1294 3048 1358 3052
rect 1294 2992 1298 3048
rect 1298 2992 1354 3048
rect 1354 2992 1358 3048
rect 1294 2988 1358 2992
rect 1374 3048 1438 3052
rect 1374 2992 1378 3048
rect 1378 2992 1434 3048
rect 1434 2992 1438 3048
rect 1374 2988 1438 2992
rect 1454 3048 1518 3052
rect 1454 2992 1458 3048
rect 1458 2992 1514 3048
rect 1514 2992 1518 3048
rect 1454 2988 1518 2992
rect 1534 3048 1598 3052
rect 1534 2992 1538 3048
rect 1538 2992 1594 3048
rect 1594 2992 1598 3048
rect 1534 2988 1598 2992
rect 1614 3048 1678 3052
rect 1614 2992 1618 3048
rect 1618 2992 1674 3048
rect 1674 2992 1678 3048
rect 1614 2988 1678 2992
rect 1694 3048 1758 3052
rect 1694 2992 1698 3048
rect 1698 2992 1754 3048
rect 1754 2992 1758 3048
rect 1694 2988 1758 2992
rect 1774 3048 1838 3052
rect 1774 2992 1778 3048
rect 1778 2992 1834 3048
rect 1834 2992 1838 3048
rect 1774 2988 1838 2992
rect 1854 3048 1918 3052
rect 1854 2992 1858 3048
rect 1858 2992 1914 3048
rect 1914 2992 1918 3048
rect 1854 2988 1918 2992
rect 1934 3048 1998 3052
rect 1934 2992 1938 3048
rect 1938 2992 1994 3048
rect 1994 2992 1998 3048
rect 1934 2988 1998 2992
rect 2014 3048 2078 3052
rect 2014 2992 2018 3048
rect 2018 2992 2074 3048
rect 2074 2992 2078 3048
rect 2014 2988 2078 2992
rect 2094 3048 2158 3052
rect 2094 2992 2098 3048
rect 2098 2992 2154 3048
rect 2154 2992 2158 3048
rect 2094 2988 2158 2992
rect 2174 3048 2238 3052
rect 2174 2992 2178 3048
rect 2178 2992 2234 3048
rect 2234 2992 2238 3048
rect 2174 2988 2238 2992
rect 2254 3048 2318 3052
rect 2254 2992 2258 3048
rect 2258 2992 2314 3048
rect 2314 2992 2318 3048
rect 2254 2988 2318 2992
rect 2334 3048 2398 3052
rect 2334 2992 2338 3048
rect 2338 2992 2394 3048
rect 2394 2992 2398 3048
rect 2334 2988 2398 2992
rect 2414 3048 2478 3052
rect 2414 2992 2418 3048
rect 2418 2992 2474 3048
rect 2474 2992 2478 3048
rect 2414 2988 2478 2992
rect 2494 3048 2558 3052
rect 2494 2992 2498 3048
rect 2498 2992 2554 3048
rect 2554 2992 2558 3048
rect 2494 2988 2558 2992
rect 714 -1072 778 -1068
rect 714 -1128 718 -1072
rect 718 -1128 774 -1072
rect 774 -1128 778 -1072
rect 714 -1132 778 -1128
rect 794 -1072 858 -1068
rect 794 -1128 798 -1072
rect 798 -1128 854 -1072
rect 854 -1128 858 -1072
rect 794 -1132 858 -1128
rect 874 -1072 938 -1068
rect 874 -1128 878 -1072
rect 878 -1128 934 -1072
rect 934 -1128 938 -1072
rect 874 -1132 938 -1128
rect 954 -1072 1018 -1068
rect 954 -1128 958 -1072
rect 958 -1128 1014 -1072
rect 1014 -1128 1018 -1072
rect 954 -1132 1018 -1128
rect 1034 -1072 1098 -1068
rect 1034 -1128 1038 -1072
rect 1038 -1128 1094 -1072
rect 1094 -1128 1098 -1072
rect 1034 -1132 1098 -1128
rect 1114 -1072 1178 -1068
rect 1114 -1128 1118 -1072
rect 1118 -1128 1174 -1072
rect 1174 -1128 1178 -1072
rect 1114 -1132 1178 -1128
rect 1194 -1072 1258 -1068
rect 1194 -1128 1198 -1072
rect 1198 -1128 1254 -1072
rect 1254 -1128 1258 -1072
rect 1194 -1132 1258 -1128
rect 1274 -1072 1338 -1068
rect 1274 -1128 1278 -1072
rect 1278 -1128 1334 -1072
rect 1334 -1128 1338 -1072
rect 1274 -1132 1338 -1128
rect 1354 -1072 1418 -1068
rect 1354 -1128 1358 -1072
rect 1358 -1128 1414 -1072
rect 1414 -1128 1418 -1072
rect 1354 -1132 1418 -1128
rect 1434 -1072 1498 -1068
rect 1434 -1128 1438 -1072
rect 1438 -1128 1494 -1072
rect 1494 -1128 1498 -1072
rect 1434 -1132 1498 -1128
rect 1514 -1072 1578 -1068
rect 1514 -1128 1518 -1072
rect 1518 -1128 1574 -1072
rect 1574 -1128 1578 -1072
rect 1514 -1132 1578 -1128
rect 1594 -1072 1658 -1068
rect 1594 -1128 1598 -1072
rect 1598 -1128 1654 -1072
rect 1654 -1128 1658 -1072
rect 1594 -1132 1658 -1128
rect 1674 -1072 1738 -1068
rect 1674 -1128 1678 -1072
rect 1678 -1128 1734 -1072
rect 1734 -1128 1738 -1072
rect 1674 -1132 1738 -1128
rect 1754 -1072 1818 -1068
rect 1754 -1128 1758 -1072
rect 1758 -1128 1814 -1072
rect 1814 -1128 1818 -1072
rect 1754 -1132 1818 -1128
rect 1834 -1072 1898 -1068
rect 1834 -1128 1838 -1072
rect 1838 -1128 1894 -1072
rect 1894 -1128 1898 -1072
rect 1834 -1132 1898 -1128
rect 1914 -1072 1978 -1068
rect 1914 -1128 1918 -1072
rect 1918 -1128 1974 -1072
rect 1974 -1128 1978 -1072
rect 1914 -1132 1978 -1128
rect 1994 -1072 2058 -1068
rect 1994 -1128 1998 -1072
rect 1998 -1128 2054 -1072
rect 2054 -1128 2058 -1072
rect 1994 -1132 2058 -1128
rect 2074 -1072 2138 -1068
rect 2074 -1128 2078 -1072
rect 2078 -1128 2134 -1072
rect 2134 -1128 2138 -1072
rect 2074 -1132 2138 -1128
rect 2154 -1072 2218 -1068
rect 2154 -1128 2158 -1072
rect 2158 -1128 2214 -1072
rect 2214 -1128 2218 -1072
rect 2154 -1132 2218 -1128
rect 2234 -1072 2298 -1068
rect 2234 -1128 2238 -1072
rect 2238 -1128 2294 -1072
rect 2294 -1128 2298 -1072
rect 2234 -1132 2298 -1128
rect 2314 -1072 2378 -1068
rect 2314 -1128 2318 -1072
rect 2318 -1128 2374 -1072
rect 2374 -1128 2378 -1072
rect 2314 -1132 2378 -1128
rect 572 -1578 576 -1354
rect 576 -1578 1112 -1354
rect 1112 -1578 1116 -1354
rect 2084 -1578 2088 -1354
rect 2088 -1578 2624 -1354
rect 2624 -1578 2628 -1354
<< metal4 >>
rect 360 3518 2840 3740
rect 360 3294 572 3518
rect 1116 3294 2084 3518
rect 2628 3294 2840 3518
rect 360 3052 2840 3294
rect 360 2988 734 3052
rect 798 2988 814 3052
rect 878 2988 894 3052
rect 958 2988 974 3052
rect 1038 2988 1054 3052
rect 1118 2988 1134 3052
rect 1198 2988 1214 3052
rect 1278 2988 1294 3052
rect 1358 2988 1374 3052
rect 1438 2988 1454 3052
rect 1518 2988 1534 3052
rect 1598 2988 1614 3052
rect 1678 2988 1694 3052
rect 1758 2988 1774 3052
rect 1838 2988 1854 3052
rect 1918 2988 1934 3052
rect 1998 2988 2014 3052
rect 2078 2988 2094 3052
rect 2158 2988 2174 3052
rect 2238 2988 2254 3052
rect 2318 2988 2334 3052
rect 2398 2988 2414 3052
rect 2478 2988 2494 3052
rect 2558 2988 2840 3052
rect 360 2940 2840 2988
rect 360 -1068 2840 -1000
rect 360 -1132 714 -1068
rect 778 -1132 794 -1068
rect 858 -1132 874 -1068
rect 938 -1132 954 -1068
rect 1018 -1132 1034 -1068
rect 1098 -1132 1114 -1068
rect 1178 -1132 1194 -1068
rect 1258 -1132 1274 -1068
rect 1338 -1132 1354 -1068
rect 1418 -1132 1434 -1068
rect 1498 -1132 1514 -1068
rect 1578 -1132 1594 -1068
rect 1658 -1132 1674 -1068
rect 1738 -1132 1754 -1068
rect 1818 -1132 1834 -1068
rect 1898 -1132 1914 -1068
rect 1978 -1132 1994 -1068
rect 2058 -1132 2074 -1068
rect 2138 -1132 2154 -1068
rect 2218 -1132 2234 -1068
rect 2298 -1132 2314 -1068
rect 2378 -1132 2840 -1068
rect 360 -1354 2840 -1132
rect 360 -1578 572 -1354
rect 1116 -1578 2084 -1354
rect 2628 -1578 2840 -1354
rect 360 -1800 2840 -1578
use sky130_fd_pr__nfet_01v8_V7QVDJ  sky130_fd_pr__nfet_01v8_V7QVDJ_0
timestamp 1626486988
transform 1 0 1571 0 1 -430
box -829 -288 829 288
use sky130_fd_pr__pfet_01v8_hvt_RC2PSP  sky130_fd_pr__pfet_01v8_hvt_RC2PSP_1
timestamp 1626486988
transform 1 0 1576 0 1 1403
box -839 -300 839 300
use sky130_fd_pr__pfet_01v8_hvt_RC2PSP  sky130_fd_pr__pfet_01v8_hvt_RC2PSP_0
timestamp 1626486988
transform 1 0 1576 0 1 2263
box -839 -300 839 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform 1 0 50 0 1 262
box -38 -48 314 592
<< labels >>
flabel metal1 s -26 494 -20 498 1 FreeSans 600 0 0 0 SEL
flabel metal2 s 1570 420 1578 428 1 FreeSans 600 0 0 0 A
flabel metal2 s 1824 440 1832 446 1 FreeSans 600 0 0 0 Y
flabel metal2 s 1048 442 1058 448 1 FreeSans 600 0 0 0 B
flabel metal2 s 434 442 444 452 1 FreeSans 600 0 0 0 SELB
flabel metal4 s 1310 3714 1322 3724 1 FreeSans 600 0 0 0 VDD
flabel metal4 s 1382 -1784 1396 -1776 1 FreeSans 600 0 0 0 VSS
<< properties >>
string FIXED_BBOX 488 -1672 2712 272
<< end >>
