magic
tech sky130A
magscale 1 2
timestamp 1623981199
<< nwell >>
rect -2562 -664 6962 2702
<< pwell >>
rect -2558 -3818 6960 -720
<< nmos >>
rect 3435 -1131 3635 -931
rect 3693 -1131 3893 -931
rect 3951 -1131 4151 -931
rect 4209 -1131 4409 -931
rect 4467 -1131 4667 -931
rect 4725 -1131 4925 -931
rect -1704 -2184 -904 -1984
rect -846 -2184 -46 -1984
rect 12 -2184 812 -1984
rect 870 -2184 1670 -1984
rect 1728 -2184 2528 -1984
rect 2586 -2184 3386 -1984
rect 3444 -2184 4244 -1984
rect 4302 -2184 5102 -1984
rect 5160 -2184 5960 -1984
rect -1704 -2766 -904 -2566
rect -846 -2766 -46 -2566
rect 12 -2766 812 -2566
rect 870 -2766 1670 -2566
rect 1728 -2766 2528 -2566
rect 2586 -2766 3386 -2566
rect 3444 -2766 4244 -2566
rect 4302 -2766 5102 -2566
rect 5160 -2766 5960 -2566
<< scnmos >>
rect -1985 -877 -1955 -793
rect -1901 -877 -1871 -793
rect -1646 -877 -1616 -793
rect -1551 -877 -1521 -805
rect -1455 -877 -1425 -805
rect -1289 -877 -1259 -793
rect -1217 -877 -1187 -793
rect -1085 -877 -1055 -749
rect -986 -877 -956 -805
rect -877 -877 -847 -805
rect -781 -877 -751 -793
rect -632 -877 -602 -793
rect -541 -877 -511 -793
rect -353 -877 -323 -747
rect -165 -877 -135 -793
rect -68 -877 -38 -747
rect 172 -877 202 -747
rect 407 -877 437 -747
rect 491 -877 521 -747
rect 730 -877 760 -747
rect 970 -877 1000 -747
rect 1067 -877 1097 -793
rect 1255 -877 1285 -747
rect 1443 -877 1473 -793
rect 1534 -877 1564 -793
rect 1683 -877 1713 -793
rect 1779 -877 1809 -805
rect 1888 -877 1918 -805
rect 1987 -877 2017 -749
rect 2119 -877 2149 -793
rect 2191 -877 2221 -793
rect 2357 -877 2387 -805
rect 2453 -877 2483 -805
rect 2548 -877 2578 -793
rect 2803 -877 2833 -793
rect 2887 -877 2917 -793
<< pmos >>
rect -2088 1396 -1288 1596
rect -1230 1396 -430 1596
rect -372 1396 428 1596
rect 486 1396 1286 1596
rect 1344 1396 2144 1596
rect 2202 1396 3002 1596
rect 3060 1396 3860 1596
rect 3918 1396 4718 1596
rect 4776 1396 5576 1596
rect 5634 1396 6434 1596
rect -2088 796 -1288 996
rect -1230 796 -430 996
rect -372 796 428 996
rect 486 796 1286 996
rect 1344 796 2144 996
rect 2202 796 3002 996
rect 3060 796 3860 996
rect 3918 796 4718 996
rect 4776 796 5576 996
rect 5634 796 6434 996
rect 3435 -444 3635 -44
rect 3693 -444 3893 -44
rect 3951 -444 4151 -44
rect 4209 -444 4409 -44
rect 4467 -444 4667 -44
rect 4725 -444 4925 -44
<< scpmoshvt >>
rect -1985 -561 -1955 -433
rect -1901 -561 -1871 -433
rect -1634 -511 -1604 -427
rect -1542 -511 -1512 -427
rect -1443 -511 -1413 -427
rect -1303 -511 -1273 -427
rect -1206 -511 -1176 -427
rect -1009 -595 -979 -427
rect -910 -511 -880 -427
rect -824 -511 -794 -427
rect -740 -511 -710 -427
rect -632 -511 -602 -427
rect -548 -511 -518 -427
rect -384 -627 -354 -427
rect -165 -555 -135 -427
rect -68 -627 -38 -427
rect 172 -627 202 -427
rect 407 -627 437 -427
rect 491 -627 521 -427
rect 730 -627 760 -427
rect 970 -627 1000 -427
rect 1067 -555 1097 -427
rect 1286 -627 1316 -427
rect 1450 -511 1480 -427
rect 1534 -511 1564 -427
rect 1642 -511 1672 -427
rect 1726 -511 1756 -427
rect 1812 -511 1842 -427
rect 1911 -595 1941 -427
rect 2108 -511 2138 -427
rect 2205 -511 2235 -427
rect 2345 -511 2375 -427
rect 2444 -511 2474 -427
rect 2536 -511 2566 -427
rect 2803 -561 2833 -433
rect 2887 -561 2917 -433
<< pmoslvt >>
rect 5331 -444 5531 -44
rect 5589 -444 5789 -44
rect 5847 -444 6047 -44
<< nmoslvt >>
rect 5331 -1131 5531 -931
rect 5589 -1131 5789 -931
rect 5847 -1131 6047 -931
<< ndiff >>
rect -2037 -805 -1985 -793
rect -2037 -839 -2029 -805
rect -1995 -839 -1985 -805
rect -2037 -877 -1985 -839
rect -1955 -831 -1901 -793
rect -1955 -865 -1945 -831
rect -1911 -865 -1901 -831
rect -1955 -877 -1901 -865
rect -1871 -805 -1819 -793
rect -1871 -839 -1861 -805
rect -1827 -839 -1819 -805
rect -1871 -877 -1819 -839
rect -1751 -835 -1646 -793
rect -1751 -869 -1739 -835
rect -1705 -869 -1646 -835
rect -1751 -877 -1646 -869
rect -1616 -805 -1566 -793
rect -1135 -793 -1085 -749
rect -1407 -805 -1289 -793
rect -1616 -829 -1551 -805
rect -1616 -863 -1606 -829
rect -1572 -863 -1551 -829
rect -1616 -877 -1551 -863
rect -1521 -829 -1455 -805
rect -1521 -863 -1499 -829
rect -1465 -863 -1455 -829
rect -1521 -877 -1455 -863
rect -1425 -877 -1289 -805
rect -1259 -877 -1217 -793
rect -1187 -831 -1085 -793
rect -1187 -865 -1153 -831
rect -1119 -865 -1085 -831
rect -1187 -877 -1085 -865
rect -1055 -805 -1001 -749
rect -405 -792 -353 -747
rect -831 -805 -781 -793
rect -1055 -835 -986 -805
rect -1055 -869 -1041 -835
rect -1007 -869 -986 -835
rect -1055 -877 -986 -869
rect -956 -831 -877 -805
rect -956 -865 -931 -831
rect -897 -865 -877 -831
rect -956 -877 -877 -865
rect -847 -877 -781 -805
rect -751 -835 -632 -793
rect -751 -869 -719 -835
rect -685 -869 -632 -835
rect -751 -877 -632 -869
rect -602 -877 -541 -793
rect -511 -815 -459 -793
rect -511 -849 -501 -815
rect -467 -849 -459 -815
rect -511 -877 -459 -849
rect -405 -826 -397 -792
rect -363 -826 -353 -792
rect -405 -877 -353 -826
rect -323 -759 -271 -747
rect -323 -793 -313 -759
rect -279 -793 -271 -759
rect -120 -793 -68 -747
rect -323 -827 -271 -793
rect -323 -861 -313 -827
rect -279 -861 -271 -827
rect -323 -877 -271 -861
rect -217 -805 -165 -793
rect -217 -839 -209 -805
rect -175 -839 -165 -805
rect -217 -877 -165 -839
rect -135 -811 -68 -793
rect -135 -845 -112 -811
rect -78 -845 -68 -811
rect -135 -877 -68 -845
rect -38 -781 14 -747
rect -38 -815 -28 -781
rect 6 -815 14 -781
rect -38 -877 14 -815
rect 120 -759 172 -747
rect 120 -793 128 -759
rect 162 -793 172 -759
rect 120 -827 172 -793
rect 120 -861 128 -827
rect 162 -861 172 -827
rect 120 -877 172 -861
rect 202 -759 254 -747
rect 202 -793 212 -759
rect 246 -793 254 -759
rect 202 -827 254 -793
rect 202 -861 212 -827
rect 246 -861 254 -827
rect 202 -877 254 -861
rect 355 -763 407 -747
rect 355 -797 363 -763
rect 397 -797 407 -763
rect 355 -831 407 -797
rect 355 -865 363 -831
rect 397 -865 407 -831
rect 355 -877 407 -865
rect 437 -877 491 -747
rect 521 -763 573 -747
rect 521 -797 531 -763
rect 565 -797 573 -763
rect 521 -831 573 -797
rect 521 -865 531 -831
rect 565 -865 573 -831
rect 521 -877 573 -865
rect 678 -759 730 -747
rect 678 -793 686 -759
rect 720 -793 730 -759
rect 678 -827 730 -793
rect 678 -861 686 -827
rect 720 -861 730 -827
rect 678 -877 730 -861
rect 760 -759 812 -747
rect 760 -793 770 -759
rect 804 -793 812 -759
rect 760 -827 812 -793
rect 760 -861 770 -827
rect 804 -861 812 -827
rect 760 -877 812 -861
rect 918 -781 970 -747
rect 918 -815 926 -781
rect 960 -815 970 -781
rect 918 -877 970 -815
rect 1000 -793 1052 -747
rect 1203 -759 1255 -747
rect 1203 -793 1211 -759
rect 1245 -793 1255 -759
rect 1000 -811 1067 -793
rect 1000 -845 1010 -811
rect 1044 -845 1067 -811
rect 1000 -877 1067 -845
rect 1097 -805 1149 -793
rect 1097 -839 1107 -805
rect 1141 -839 1149 -805
rect 1097 -877 1149 -839
rect 1203 -827 1255 -793
rect 1203 -861 1211 -827
rect 1245 -861 1255 -827
rect 1203 -877 1255 -861
rect 1285 -792 1337 -747
rect 1285 -826 1295 -792
rect 1329 -826 1337 -792
rect 1285 -877 1337 -826
rect 1391 -815 1443 -793
rect 1391 -849 1399 -815
rect 1433 -849 1443 -815
rect 1391 -877 1443 -849
rect 1473 -877 1534 -793
rect 1564 -835 1683 -793
rect 1564 -869 1617 -835
rect 1651 -869 1683 -835
rect 1564 -877 1683 -869
rect 1713 -805 1763 -793
rect 1933 -805 1987 -749
rect 1713 -877 1779 -805
rect 1809 -831 1888 -805
rect 1809 -865 1829 -831
rect 1863 -865 1888 -831
rect 1809 -877 1888 -865
rect 1918 -835 1987 -805
rect 1918 -869 1939 -835
rect 1973 -869 1987 -835
rect 1918 -877 1987 -869
rect 2017 -793 2067 -749
rect 2017 -831 2119 -793
rect 2017 -865 2051 -831
rect 2085 -865 2119 -831
rect 2017 -877 2119 -865
rect 2149 -877 2191 -793
rect 2221 -805 2339 -793
rect 2498 -805 2548 -793
rect 2221 -877 2357 -805
rect 2387 -829 2453 -805
rect 2387 -863 2397 -829
rect 2431 -863 2453 -829
rect 2387 -877 2453 -863
rect 2483 -829 2548 -805
rect 2483 -863 2504 -829
rect 2538 -863 2548 -829
rect 2483 -877 2548 -863
rect 2578 -835 2683 -793
rect 2578 -869 2637 -835
rect 2671 -869 2683 -835
rect 2578 -877 2683 -869
rect 2751 -805 2803 -793
rect 2751 -839 2759 -805
rect 2793 -839 2803 -805
rect 2751 -877 2803 -839
rect 2833 -831 2887 -793
rect 2833 -865 2843 -831
rect 2877 -865 2887 -831
rect 2833 -877 2887 -865
rect 2917 -805 2969 -793
rect 2917 -839 2927 -805
rect 2961 -839 2969 -805
rect 2917 -877 2969 -839
rect 3377 -943 3435 -931
rect 3377 -1119 3389 -943
rect 3423 -1119 3435 -943
rect 3377 -1131 3435 -1119
rect 3635 -943 3693 -931
rect 3635 -1119 3647 -943
rect 3681 -1119 3693 -943
rect 3635 -1131 3693 -1119
rect 3893 -943 3951 -931
rect 3893 -1119 3905 -943
rect 3939 -1119 3951 -943
rect 3893 -1131 3951 -1119
rect 4151 -943 4209 -931
rect 4151 -1119 4163 -943
rect 4197 -1119 4209 -943
rect 4151 -1131 4209 -1119
rect 4409 -943 4467 -931
rect 4409 -1119 4421 -943
rect 4455 -1119 4467 -943
rect 4409 -1131 4467 -1119
rect 4667 -943 4725 -931
rect 4667 -1119 4679 -943
rect 4713 -1119 4725 -943
rect 4667 -1131 4725 -1119
rect 4925 -943 4983 -931
rect 4925 -1119 4937 -943
rect 4971 -1119 4983 -943
rect 4925 -1131 4983 -1119
rect 5273 -943 5331 -931
rect 5273 -1119 5285 -943
rect 5319 -1119 5331 -943
rect 5273 -1131 5331 -1119
rect 5531 -943 5589 -931
rect 5531 -1119 5543 -943
rect 5577 -1119 5589 -943
rect 5531 -1131 5589 -1119
rect 5789 -943 5847 -931
rect 5789 -1119 5801 -943
rect 5835 -1119 5847 -943
rect 5789 -1131 5847 -1119
rect 6047 -943 6105 -931
rect 6047 -1119 6059 -943
rect 6093 -1119 6105 -943
rect 6047 -1131 6105 -1119
rect -1762 -1996 -1704 -1984
rect -1762 -2172 -1750 -1996
rect -1716 -2172 -1704 -1996
rect -1762 -2184 -1704 -2172
rect -904 -1996 -846 -1984
rect -904 -2172 -892 -1996
rect -858 -2172 -846 -1996
rect -904 -2184 -846 -2172
rect -46 -1996 12 -1984
rect -46 -2172 -34 -1996
rect 0 -2172 12 -1996
rect -46 -2184 12 -2172
rect 812 -1996 870 -1984
rect 812 -2172 824 -1996
rect 858 -2172 870 -1996
rect 812 -2184 870 -2172
rect 1670 -1996 1728 -1984
rect 1670 -2172 1682 -1996
rect 1716 -2172 1728 -1996
rect 1670 -2184 1728 -2172
rect 2528 -1996 2586 -1984
rect 2528 -2172 2540 -1996
rect 2574 -2172 2586 -1996
rect 2528 -2184 2586 -2172
rect 3386 -1996 3444 -1984
rect 3386 -2172 3398 -1996
rect 3432 -2172 3444 -1996
rect 3386 -2184 3444 -2172
rect 4244 -1996 4302 -1984
rect 4244 -2172 4256 -1996
rect 4290 -2172 4302 -1996
rect 4244 -2184 4302 -2172
rect 5102 -1996 5160 -1984
rect 5102 -2172 5114 -1996
rect 5148 -2172 5160 -1996
rect 5102 -2184 5160 -2172
rect 5960 -1996 6018 -1984
rect 5960 -2172 5972 -1996
rect 6006 -2172 6018 -1996
rect 5960 -2184 6018 -2172
rect -1762 -2578 -1704 -2566
rect -1762 -2754 -1750 -2578
rect -1716 -2754 -1704 -2578
rect -1762 -2766 -1704 -2754
rect -904 -2578 -846 -2566
rect -904 -2754 -892 -2578
rect -858 -2754 -846 -2578
rect -904 -2766 -846 -2754
rect -46 -2578 12 -2566
rect -46 -2754 -34 -2578
rect 0 -2754 12 -2578
rect -46 -2766 12 -2754
rect 812 -2578 870 -2566
rect 812 -2754 824 -2578
rect 858 -2754 870 -2578
rect 812 -2766 870 -2754
rect 1670 -2578 1728 -2566
rect 1670 -2754 1682 -2578
rect 1716 -2754 1728 -2578
rect 1670 -2766 1728 -2754
rect 2528 -2578 2586 -2566
rect 2528 -2754 2540 -2578
rect 2574 -2754 2586 -2578
rect 2528 -2766 2586 -2754
rect 3386 -2578 3444 -2566
rect 3386 -2754 3398 -2578
rect 3432 -2754 3444 -2578
rect 3386 -2766 3444 -2754
rect 4244 -2578 4302 -2566
rect 4244 -2754 4256 -2578
rect 4290 -2754 4302 -2578
rect 4244 -2766 4302 -2754
rect 5102 -2578 5160 -2566
rect 5102 -2754 5114 -2578
rect 5148 -2754 5160 -2578
rect 5102 -2766 5160 -2754
rect 5960 -2578 6018 -2566
rect 5960 -2754 5972 -2578
rect 6006 -2754 6018 -2578
rect 5960 -2766 6018 -2754
<< pdiff >>
rect -2146 1584 -2088 1596
rect -2146 1408 -2134 1584
rect -2100 1408 -2088 1584
rect -2146 1396 -2088 1408
rect -1288 1584 -1230 1596
rect -1288 1408 -1276 1584
rect -1242 1408 -1230 1584
rect -1288 1396 -1230 1408
rect -430 1584 -372 1596
rect -430 1408 -418 1584
rect -384 1408 -372 1584
rect -430 1396 -372 1408
rect 428 1584 486 1596
rect 428 1408 440 1584
rect 474 1408 486 1584
rect 428 1396 486 1408
rect 1286 1584 1344 1596
rect 1286 1408 1298 1584
rect 1332 1408 1344 1584
rect 1286 1396 1344 1408
rect 2144 1584 2202 1596
rect 2144 1408 2156 1584
rect 2190 1408 2202 1584
rect 2144 1396 2202 1408
rect 3002 1584 3060 1596
rect 3002 1408 3014 1584
rect 3048 1408 3060 1584
rect 3002 1396 3060 1408
rect 3860 1584 3918 1596
rect 3860 1408 3872 1584
rect 3906 1408 3918 1584
rect 3860 1396 3918 1408
rect 4718 1584 4776 1596
rect 4718 1408 4730 1584
rect 4764 1408 4776 1584
rect 4718 1396 4776 1408
rect 5576 1584 5634 1596
rect 5576 1408 5588 1584
rect 5622 1408 5634 1584
rect 5576 1396 5634 1408
rect 6434 1584 6492 1596
rect 6434 1408 6446 1584
rect 6480 1408 6492 1584
rect 6434 1396 6492 1408
rect -2146 984 -2088 996
rect -2146 808 -2134 984
rect -2100 808 -2088 984
rect -2146 796 -2088 808
rect -1288 984 -1230 996
rect -1288 808 -1276 984
rect -1242 808 -1230 984
rect -1288 796 -1230 808
rect -430 984 -372 996
rect -430 808 -418 984
rect -384 808 -372 984
rect -430 796 -372 808
rect 428 984 486 996
rect 428 808 440 984
rect 474 808 486 984
rect 428 796 486 808
rect 1286 984 1344 996
rect 1286 808 1298 984
rect 1332 808 1344 984
rect 1286 796 1344 808
rect 2144 984 2202 996
rect 2144 808 2156 984
rect 2190 808 2202 984
rect 2144 796 2202 808
rect 3002 984 3060 996
rect 3002 808 3014 984
rect 3048 808 3060 984
rect 3002 796 3060 808
rect 3860 984 3918 996
rect 3860 808 3872 984
rect 3906 808 3918 984
rect 3860 796 3918 808
rect 4718 984 4776 996
rect 4718 808 4730 984
rect 4764 808 4776 984
rect 4718 796 4776 808
rect 5576 984 5634 996
rect 5576 808 5588 984
rect 5622 808 5634 984
rect 5576 796 5634 808
rect 6434 984 6492 996
rect 6434 808 6446 984
rect 6480 808 6492 984
rect 6434 796 6492 808
rect -2037 -447 -1985 -433
rect -2037 -481 -2029 -447
rect -1995 -481 -1985 -447
rect -2037 -515 -1985 -481
rect -2037 -549 -2029 -515
rect -1995 -549 -1985 -515
rect -2037 -561 -1985 -549
rect -1955 -463 -1901 -433
rect -1955 -497 -1945 -463
rect -1911 -497 -1901 -463
rect -1955 -561 -1901 -497
rect -1871 -447 -1819 -433
rect -1871 -481 -1861 -447
rect -1827 -481 -1819 -447
rect -1871 -515 -1819 -481
rect -1686 -439 -1634 -427
rect -1686 -473 -1678 -439
rect -1644 -473 -1634 -439
rect -1686 -511 -1634 -473
rect -1604 -447 -1542 -427
rect -1604 -481 -1594 -447
rect -1560 -481 -1542 -447
rect -1604 -511 -1542 -481
rect -1512 -441 -1443 -427
rect -1512 -475 -1501 -441
rect -1467 -475 -1443 -441
rect -1512 -511 -1443 -475
rect -1413 -465 -1303 -427
rect -1413 -499 -1347 -465
rect -1313 -499 -1303 -465
rect -1413 -511 -1303 -499
rect -1273 -449 -1206 -427
rect -1273 -483 -1250 -449
rect -1216 -483 -1206 -449
rect -1273 -511 -1206 -483
rect -1176 -465 -1124 -427
rect -1176 -499 -1166 -465
rect -1132 -499 -1124 -465
rect -1176 -511 -1124 -499
rect -1061 -439 -1009 -427
rect -1061 -473 -1053 -439
rect -1019 -473 -1009 -439
rect -1871 -549 -1861 -515
rect -1827 -549 -1819 -515
rect -1871 -561 -1819 -549
rect -1061 -595 -1009 -473
rect -979 -447 -910 -427
rect -979 -481 -965 -447
rect -931 -481 -910 -447
rect -979 -511 -910 -481
rect -880 -440 -824 -427
rect -880 -474 -868 -440
rect -834 -474 -824 -440
rect -880 -511 -824 -474
rect -794 -511 -740 -427
rect -710 -439 -632 -427
rect -710 -473 -676 -439
rect -642 -473 -632 -439
rect -710 -511 -632 -473
rect -602 -465 -548 -427
rect -602 -499 -592 -465
rect -558 -499 -548 -465
rect -602 -511 -548 -499
rect -518 -439 -384 -427
rect -518 -473 -506 -439
rect -472 -473 -428 -439
rect -394 -473 -384 -439
rect -518 -511 -384 -473
rect -979 -595 -925 -511
rect -434 -627 -384 -511
rect -354 -447 -298 -427
rect -354 -481 -344 -447
rect -310 -481 -298 -447
rect -354 -515 -298 -481
rect -354 -549 -344 -515
rect -310 -549 -298 -515
rect -354 -583 -298 -549
rect -217 -439 -165 -427
rect -217 -473 -209 -439
rect -175 -473 -165 -439
rect -217 -507 -165 -473
rect -217 -541 -209 -507
rect -175 -541 -165 -507
rect -217 -555 -165 -541
rect -135 -439 -68 -427
rect -135 -473 -112 -439
rect -78 -473 -68 -439
rect -135 -507 -68 -473
rect -135 -541 -112 -507
rect -78 -541 -68 -507
rect -135 -555 -68 -541
rect -354 -617 -344 -583
rect -310 -617 -298 -583
rect -354 -627 -298 -617
rect -120 -575 -68 -555
rect -120 -609 -112 -575
rect -78 -609 -68 -575
rect -120 -627 -68 -609
rect -38 -475 14 -427
rect -38 -509 -28 -475
rect 6 -509 14 -475
rect -38 -543 14 -509
rect -38 -577 -28 -543
rect 6 -577 14 -543
rect -38 -627 14 -577
rect 120 -439 172 -427
rect 120 -473 128 -439
rect 162 -473 172 -439
rect 120 -507 172 -473
rect 120 -541 128 -507
rect 162 -541 172 -507
rect 120 -575 172 -541
rect 120 -609 128 -575
rect 162 -609 172 -575
rect 120 -627 172 -609
rect 202 -439 254 -427
rect 202 -473 212 -439
rect 246 -473 254 -439
rect 202 -507 254 -473
rect 202 -541 212 -507
rect 246 -541 254 -507
rect 202 -575 254 -541
rect 202 -609 212 -575
rect 246 -609 254 -575
rect 202 -627 254 -609
rect 355 -439 407 -427
rect 355 -473 363 -439
rect 397 -473 407 -439
rect 355 -507 407 -473
rect 355 -541 363 -507
rect 397 -541 407 -507
rect 355 -575 407 -541
rect 355 -609 363 -575
rect 397 -609 407 -575
rect 355 -627 407 -609
rect 437 -439 491 -427
rect 437 -473 447 -439
rect 481 -473 491 -439
rect 437 -507 491 -473
rect 437 -541 447 -507
rect 481 -541 491 -507
rect 437 -575 491 -541
rect 437 -609 447 -575
rect 481 -609 491 -575
rect 437 -627 491 -609
rect 521 -439 573 -427
rect 521 -473 531 -439
rect 565 -473 573 -439
rect 521 -507 573 -473
rect 521 -541 531 -507
rect 565 -541 573 -507
rect 521 -575 573 -541
rect 521 -609 531 -575
rect 565 -609 573 -575
rect 521 -627 573 -609
rect 678 -439 730 -427
rect 678 -473 686 -439
rect 720 -473 730 -439
rect 678 -507 730 -473
rect 678 -541 686 -507
rect 720 -541 730 -507
rect 678 -575 730 -541
rect 678 -609 686 -575
rect 720 -609 730 -575
rect 678 -627 730 -609
rect 760 -439 812 -427
rect 760 -473 770 -439
rect 804 -473 812 -439
rect 760 -507 812 -473
rect 760 -541 770 -507
rect 804 -541 812 -507
rect 760 -575 812 -541
rect 760 -609 770 -575
rect 804 -609 812 -575
rect 760 -627 812 -609
rect 918 -475 970 -427
rect 918 -509 926 -475
rect 960 -509 970 -475
rect 918 -543 970 -509
rect 918 -577 926 -543
rect 960 -577 970 -543
rect 918 -627 970 -577
rect 1000 -439 1067 -427
rect 1000 -473 1010 -439
rect 1044 -473 1067 -439
rect 1000 -507 1067 -473
rect 1000 -541 1010 -507
rect 1044 -541 1067 -507
rect 1000 -555 1067 -541
rect 1097 -439 1149 -427
rect 1097 -473 1107 -439
rect 1141 -473 1149 -439
rect 1097 -507 1149 -473
rect 1097 -541 1107 -507
rect 1141 -541 1149 -507
rect 1097 -555 1149 -541
rect 1230 -447 1286 -427
rect 1230 -481 1242 -447
rect 1276 -481 1286 -447
rect 1230 -515 1286 -481
rect 1230 -549 1242 -515
rect 1276 -549 1286 -515
rect 1000 -575 1052 -555
rect 1000 -609 1010 -575
rect 1044 -609 1052 -575
rect 1000 -627 1052 -609
rect 1230 -583 1286 -549
rect 1230 -617 1242 -583
rect 1276 -617 1286 -583
rect 1230 -627 1286 -617
rect 1316 -439 1450 -427
rect 1316 -473 1326 -439
rect 1360 -473 1404 -439
rect 1438 -473 1450 -439
rect 1316 -511 1450 -473
rect 1480 -465 1534 -427
rect 1480 -499 1490 -465
rect 1524 -499 1534 -465
rect 1480 -511 1534 -499
rect 1564 -439 1642 -427
rect 1564 -473 1574 -439
rect 1608 -473 1642 -439
rect 1564 -511 1642 -473
rect 1672 -511 1726 -427
rect 1756 -440 1812 -427
rect 1756 -474 1766 -440
rect 1800 -474 1812 -440
rect 1756 -511 1812 -474
rect 1842 -447 1911 -427
rect 1842 -481 1863 -447
rect 1897 -481 1911 -447
rect 1842 -511 1911 -481
rect 1316 -627 1366 -511
rect 1857 -595 1911 -511
rect 1941 -439 1993 -427
rect 1941 -473 1951 -439
rect 1985 -473 1993 -439
rect 1941 -595 1993 -473
rect 2056 -465 2108 -427
rect 2056 -499 2064 -465
rect 2098 -499 2108 -465
rect 2056 -511 2108 -499
rect 2138 -449 2205 -427
rect 2138 -483 2148 -449
rect 2182 -483 2205 -449
rect 2138 -511 2205 -483
rect 2235 -465 2345 -427
rect 2235 -499 2245 -465
rect 2279 -499 2345 -465
rect 2235 -511 2345 -499
rect 2375 -441 2444 -427
rect 2375 -475 2399 -441
rect 2433 -475 2444 -441
rect 2375 -511 2444 -475
rect 2474 -447 2536 -427
rect 2474 -481 2492 -447
rect 2526 -481 2536 -447
rect 2474 -511 2536 -481
rect 2566 -439 2618 -427
rect 2566 -473 2576 -439
rect 2610 -473 2618 -439
rect 2566 -511 2618 -473
rect 2751 -447 2803 -433
rect 2751 -481 2759 -447
rect 2793 -481 2803 -447
rect 2751 -515 2803 -481
rect 2751 -549 2759 -515
rect 2793 -549 2803 -515
rect 2751 -561 2803 -549
rect 2833 -463 2887 -433
rect 2833 -497 2843 -463
rect 2877 -497 2887 -463
rect 2833 -561 2887 -497
rect 2917 -447 2969 -433
rect 2917 -481 2927 -447
rect 2961 -481 2969 -447
rect 2917 -515 2969 -481
rect 2917 -549 2927 -515
rect 2961 -549 2969 -515
rect 2917 -561 2969 -549
rect 3377 -56 3435 -44
rect 3377 -432 3389 -56
rect 3423 -432 3435 -56
rect 3377 -444 3435 -432
rect 3635 -56 3693 -44
rect 3635 -432 3647 -56
rect 3681 -432 3693 -56
rect 3635 -444 3693 -432
rect 3893 -56 3951 -44
rect 3893 -432 3905 -56
rect 3939 -432 3951 -56
rect 3893 -444 3951 -432
rect 4151 -56 4209 -44
rect 4151 -432 4163 -56
rect 4197 -432 4209 -56
rect 4151 -444 4209 -432
rect 4409 -56 4467 -44
rect 4409 -432 4421 -56
rect 4455 -432 4467 -56
rect 4409 -444 4467 -432
rect 4667 -56 4725 -44
rect 4667 -432 4679 -56
rect 4713 -432 4725 -56
rect 4667 -444 4725 -432
rect 4925 -56 4983 -44
rect 4925 -432 4937 -56
rect 4971 -432 4983 -56
rect 4925 -444 4983 -432
rect 5273 -56 5331 -44
rect 5273 -432 5285 -56
rect 5319 -432 5331 -56
rect 5273 -444 5331 -432
rect 5531 -56 5589 -44
rect 5531 -432 5543 -56
rect 5577 -432 5589 -56
rect 5531 -444 5589 -432
rect 5789 -56 5847 -44
rect 5789 -432 5801 -56
rect 5835 -432 5847 -56
rect 5789 -444 5847 -432
rect 6047 -56 6105 -44
rect 6047 -432 6059 -56
rect 6093 -432 6105 -56
rect 6047 -444 6105 -432
<< ndiffc >>
rect -2029 -839 -1995 -805
rect -1945 -865 -1911 -831
rect -1861 -839 -1827 -805
rect -1739 -869 -1705 -835
rect -1606 -863 -1572 -829
rect -1499 -863 -1465 -829
rect -1153 -865 -1119 -831
rect -1041 -869 -1007 -835
rect -931 -865 -897 -831
rect -719 -869 -685 -835
rect -501 -849 -467 -815
rect -397 -826 -363 -792
rect -313 -793 -279 -759
rect -313 -861 -279 -827
rect -209 -839 -175 -805
rect -112 -845 -78 -811
rect -28 -815 6 -781
rect 128 -793 162 -759
rect 128 -861 162 -827
rect 212 -793 246 -759
rect 212 -861 246 -827
rect 363 -797 397 -763
rect 363 -865 397 -831
rect 531 -797 565 -763
rect 531 -865 565 -831
rect 686 -793 720 -759
rect 686 -861 720 -827
rect 770 -793 804 -759
rect 770 -861 804 -827
rect 926 -815 960 -781
rect 1211 -793 1245 -759
rect 1010 -845 1044 -811
rect 1107 -839 1141 -805
rect 1211 -861 1245 -827
rect 1295 -826 1329 -792
rect 1399 -849 1433 -815
rect 1617 -869 1651 -835
rect 1829 -865 1863 -831
rect 1939 -869 1973 -835
rect 2051 -865 2085 -831
rect 2397 -863 2431 -829
rect 2504 -863 2538 -829
rect 2637 -869 2671 -835
rect 2759 -839 2793 -805
rect 2843 -865 2877 -831
rect 2927 -839 2961 -805
rect 3389 -1119 3423 -943
rect 3647 -1119 3681 -943
rect 3905 -1119 3939 -943
rect 4163 -1119 4197 -943
rect 4421 -1119 4455 -943
rect 4679 -1119 4713 -943
rect 4937 -1119 4971 -943
rect 5285 -1119 5319 -943
rect 5543 -1119 5577 -943
rect 5801 -1119 5835 -943
rect 6059 -1119 6093 -943
rect -1750 -2172 -1716 -1996
rect -892 -2172 -858 -1996
rect -34 -2172 0 -1996
rect 824 -2172 858 -1996
rect 1682 -2172 1716 -1996
rect 2540 -2172 2574 -1996
rect 3398 -2172 3432 -1996
rect 4256 -2172 4290 -1996
rect 5114 -2172 5148 -1996
rect 5972 -2172 6006 -1996
rect -1750 -2754 -1716 -2578
rect -892 -2754 -858 -2578
rect -34 -2754 0 -2578
rect 824 -2754 858 -2578
rect 1682 -2754 1716 -2578
rect 2540 -2754 2574 -2578
rect 3398 -2754 3432 -2578
rect 4256 -2754 4290 -2578
rect 5114 -2754 5148 -2578
rect 5972 -2754 6006 -2578
<< pdiffc >>
rect -2134 1408 -2100 1584
rect -1276 1408 -1242 1584
rect -418 1408 -384 1584
rect 440 1408 474 1584
rect 1298 1408 1332 1584
rect 2156 1408 2190 1584
rect 3014 1408 3048 1584
rect 3872 1408 3906 1584
rect 4730 1408 4764 1584
rect 5588 1408 5622 1584
rect 6446 1408 6480 1584
rect -2134 808 -2100 984
rect -1276 808 -1242 984
rect -418 808 -384 984
rect 440 808 474 984
rect 1298 808 1332 984
rect 2156 808 2190 984
rect 3014 808 3048 984
rect 3872 808 3906 984
rect 4730 808 4764 984
rect 5588 808 5622 984
rect 6446 808 6480 984
rect -2029 -481 -1995 -447
rect -2029 -549 -1995 -515
rect -1945 -497 -1911 -463
rect -1861 -481 -1827 -447
rect -1678 -473 -1644 -439
rect -1594 -481 -1560 -447
rect -1501 -475 -1467 -441
rect -1347 -499 -1313 -465
rect -1250 -483 -1216 -449
rect -1166 -499 -1132 -465
rect -1053 -473 -1019 -439
rect -1861 -549 -1827 -515
rect -965 -481 -931 -447
rect -868 -474 -834 -440
rect -676 -473 -642 -439
rect -592 -499 -558 -465
rect -506 -473 -472 -439
rect -428 -473 -394 -439
rect -344 -481 -310 -447
rect -344 -549 -310 -515
rect -209 -473 -175 -439
rect -209 -541 -175 -507
rect -112 -473 -78 -439
rect -112 -541 -78 -507
rect -344 -617 -310 -583
rect -112 -609 -78 -575
rect -28 -509 6 -475
rect -28 -577 6 -543
rect 128 -473 162 -439
rect 128 -541 162 -507
rect 128 -609 162 -575
rect 212 -473 246 -439
rect 212 -541 246 -507
rect 212 -609 246 -575
rect 363 -473 397 -439
rect 363 -541 397 -507
rect 363 -609 397 -575
rect 447 -473 481 -439
rect 447 -541 481 -507
rect 447 -609 481 -575
rect 531 -473 565 -439
rect 531 -541 565 -507
rect 531 -609 565 -575
rect 686 -473 720 -439
rect 686 -541 720 -507
rect 686 -609 720 -575
rect 770 -473 804 -439
rect 770 -541 804 -507
rect 770 -609 804 -575
rect 926 -509 960 -475
rect 926 -577 960 -543
rect 1010 -473 1044 -439
rect 1010 -541 1044 -507
rect 1107 -473 1141 -439
rect 1107 -541 1141 -507
rect 1242 -481 1276 -447
rect 1242 -549 1276 -515
rect 1010 -609 1044 -575
rect 1242 -617 1276 -583
rect 1326 -473 1360 -439
rect 1404 -473 1438 -439
rect 1490 -499 1524 -465
rect 1574 -473 1608 -439
rect 1766 -474 1800 -440
rect 1863 -481 1897 -447
rect 1951 -473 1985 -439
rect 2064 -499 2098 -465
rect 2148 -483 2182 -449
rect 2245 -499 2279 -465
rect 2399 -475 2433 -441
rect 2492 -481 2526 -447
rect 2576 -473 2610 -439
rect 2759 -481 2793 -447
rect 2759 -549 2793 -515
rect 2843 -497 2877 -463
rect 2927 -481 2961 -447
rect 2927 -549 2961 -515
rect 3389 -432 3423 -56
rect 3647 -432 3681 -56
rect 3905 -432 3939 -56
rect 4163 -432 4197 -56
rect 4421 -432 4455 -56
rect 4679 -432 4713 -56
rect 4937 -432 4971 -56
rect 5285 -432 5319 -56
rect 5543 -432 5577 -56
rect 5801 -432 5835 -56
rect 6059 -432 6093 -56
<< psubdiff >>
rect 3275 -791 3371 -757
rect 4989 -791 5085 -757
rect 3275 -853 3309 -791
rect 5051 -853 5085 -791
rect 3275 -1271 3309 -1209
rect 5051 -1271 5085 -1209
rect 3275 -1305 3371 -1271
rect 4989 -1305 5085 -1271
rect 5171 -791 5267 -757
rect 6111 -791 6207 -757
rect 5171 -853 5205 -791
rect 6173 -853 6207 -791
rect 5171 -1271 5205 -1209
rect 6173 -1271 6207 -1209
rect 5171 -1305 5267 -1271
rect 6111 -1305 6207 -1271
rect -2522 -1618 -2360 -1518
rect 6760 -1618 6922 -1518
rect -2522 -1680 -2422 -1618
rect 6822 -1680 6922 -1618
rect -2522 -3682 -2422 -3620
rect 6822 -3682 6922 -3620
rect -2522 -3782 -2360 -3682
rect 6760 -3782 6922 -3682
<< nsubdiff >>
rect -2522 2562 -2360 2662
rect 6760 2562 6922 2662
rect -2522 2500 -2422 2562
rect 6822 2500 6922 2562
rect -2522 458 -2422 520
rect 6822 458 6922 520
rect -2522 358 -2360 458
rect 6760 358 6922 458
rect 3275 105 3371 139
rect 4989 105 5085 139
rect 3275 43 3309 105
rect 5051 43 5085 105
rect 3275 -593 3309 -531
rect 5051 -593 5085 -531
rect 3275 -627 3371 -593
rect 4989 -627 5085 -593
rect 5171 105 5267 139
rect 6111 105 6207 139
rect 5171 43 5205 105
rect 6173 43 6207 105
rect 5171 -593 5205 -531
rect 6173 -593 6207 -531
rect 5171 -627 5267 -593
rect 6111 -627 6207 -593
<< psubdiffcont >>
rect 3371 -791 4989 -757
rect 3275 -1209 3309 -853
rect 5051 -1209 5085 -853
rect 3371 -1305 4989 -1271
rect 5267 -791 6111 -757
rect 5171 -1209 5205 -853
rect 6173 -1209 6207 -853
rect 5267 -1305 6111 -1271
rect -2360 -1618 6760 -1518
rect -2522 -3620 -2422 -1680
rect 6822 -3620 6922 -1680
rect -2360 -3782 6760 -3682
<< nsubdiffcont >>
rect -2360 2562 6760 2662
rect -2522 520 -2422 2500
rect 6822 520 6922 2500
rect -2360 358 6760 458
rect 3371 105 4989 139
rect 3275 -531 3309 43
rect 5051 -531 5085 43
rect 3371 -627 4989 -593
rect 5267 105 6111 139
rect 5171 -531 5205 43
rect 6173 -531 6207 43
rect 5267 -627 6111 -593
<< poly >>
rect -1896 1677 -1480 1693
rect -1896 1660 -1880 1677
rect -2088 1643 -1880 1660
rect -1496 1660 -1480 1677
rect -1038 1677 -622 1693
rect -1038 1660 -1022 1677
rect -1496 1643 -1288 1660
rect -2088 1596 -1288 1643
rect -1230 1643 -1022 1660
rect -638 1660 -622 1677
rect -180 1677 236 1693
rect -180 1660 -164 1677
rect -638 1643 -430 1660
rect -1230 1596 -430 1643
rect -372 1643 -164 1660
rect 220 1660 236 1677
rect 678 1677 1094 1693
rect 678 1660 694 1677
rect 220 1643 428 1660
rect -372 1596 428 1643
rect 486 1643 694 1660
rect 1078 1660 1094 1677
rect 1536 1677 1952 1693
rect 1536 1660 1552 1677
rect 1078 1643 1286 1660
rect 486 1596 1286 1643
rect 1344 1643 1552 1660
rect 1936 1660 1952 1677
rect 2394 1677 2810 1693
rect 2394 1660 2410 1677
rect 1936 1643 2144 1660
rect 1344 1596 2144 1643
rect 2202 1643 2410 1660
rect 2794 1660 2810 1677
rect 3252 1677 3668 1693
rect 3252 1660 3268 1677
rect 2794 1643 3002 1660
rect 2202 1596 3002 1643
rect 3060 1643 3268 1660
rect 3652 1660 3668 1677
rect 4110 1677 4526 1693
rect 4110 1660 4126 1677
rect 3652 1643 3860 1660
rect 3060 1596 3860 1643
rect 3918 1643 4126 1660
rect 4510 1660 4526 1677
rect 4968 1677 5384 1693
rect 4968 1660 4984 1677
rect 4510 1643 4718 1660
rect 3918 1596 4718 1643
rect 4776 1643 4984 1660
rect 5368 1660 5384 1677
rect 5826 1677 6242 1693
rect 5826 1660 5842 1677
rect 5368 1643 5576 1660
rect 4776 1596 5576 1643
rect 5634 1643 5842 1660
rect 6226 1660 6242 1677
rect 6226 1643 6434 1660
rect 5634 1596 6434 1643
rect -2088 1349 -1288 1396
rect -2088 1332 -1880 1349
rect -1896 1315 -1880 1332
rect -1496 1332 -1288 1349
rect -1230 1349 -430 1396
rect -1230 1332 -1022 1349
rect -1496 1315 -1480 1332
rect -1896 1299 -1480 1315
rect -1038 1315 -1022 1332
rect -638 1332 -430 1349
rect -372 1349 428 1396
rect -372 1332 -164 1349
rect -638 1315 -622 1332
rect -1038 1299 -622 1315
rect -180 1315 -164 1332
rect 220 1332 428 1349
rect 486 1349 1286 1396
rect 486 1332 694 1349
rect 220 1315 236 1332
rect -180 1299 236 1315
rect 678 1315 694 1332
rect 1078 1332 1286 1349
rect 1344 1349 2144 1396
rect 1344 1332 1552 1349
rect 1078 1315 1094 1332
rect 678 1299 1094 1315
rect 1536 1315 1552 1332
rect 1936 1332 2144 1349
rect 2202 1349 3002 1396
rect 2202 1332 2410 1349
rect 1936 1315 1952 1332
rect 1536 1299 1952 1315
rect 2394 1315 2410 1332
rect 2794 1332 3002 1349
rect 3060 1349 3860 1396
rect 3060 1332 3268 1349
rect 2794 1315 2810 1332
rect 2394 1299 2810 1315
rect 3252 1315 3268 1332
rect 3652 1332 3860 1349
rect 3918 1349 4718 1396
rect 3918 1332 4126 1349
rect 3652 1315 3668 1332
rect 3252 1299 3668 1315
rect 4110 1315 4126 1332
rect 4510 1332 4718 1349
rect 4776 1349 5576 1396
rect 4776 1332 4984 1349
rect 4510 1315 4526 1332
rect 4110 1299 4526 1315
rect 4968 1315 4984 1332
rect 5368 1332 5576 1349
rect 5634 1349 6434 1396
rect 5634 1332 5842 1349
rect 5368 1315 5384 1332
rect 4968 1299 5384 1315
rect 5826 1315 5842 1332
rect 6226 1332 6434 1349
rect 6226 1315 6242 1332
rect 5826 1299 6242 1315
rect -1896 1077 -1480 1093
rect -1896 1060 -1880 1077
rect -2088 1043 -1880 1060
rect -1496 1060 -1480 1077
rect -1038 1077 -622 1093
rect -1038 1060 -1022 1077
rect -1496 1043 -1288 1060
rect -2088 996 -1288 1043
rect -1230 1043 -1022 1060
rect -638 1060 -622 1077
rect -180 1077 236 1093
rect -180 1060 -164 1077
rect -638 1043 -430 1060
rect -1230 996 -430 1043
rect -372 1043 -164 1060
rect 220 1060 236 1077
rect 678 1077 1094 1093
rect 678 1060 694 1077
rect 220 1043 428 1060
rect -372 996 428 1043
rect 486 1043 694 1060
rect 1078 1060 1094 1077
rect 1536 1077 1952 1093
rect 1536 1060 1552 1077
rect 1078 1043 1286 1060
rect 486 996 1286 1043
rect 1344 1043 1552 1060
rect 1936 1060 1952 1077
rect 2394 1077 2810 1093
rect 2394 1060 2410 1077
rect 1936 1043 2144 1060
rect 1344 996 2144 1043
rect 2202 1043 2410 1060
rect 2794 1060 2810 1077
rect 3252 1077 3668 1093
rect 3252 1060 3268 1077
rect 2794 1043 3002 1060
rect 2202 996 3002 1043
rect 3060 1043 3268 1060
rect 3652 1060 3668 1077
rect 4110 1077 4526 1093
rect 4110 1060 4126 1077
rect 3652 1043 3860 1060
rect 3060 996 3860 1043
rect 3918 1043 4126 1060
rect 4510 1060 4526 1077
rect 4968 1077 5384 1093
rect 4968 1060 4984 1077
rect 4510 1043 4718 1060
rect 3918 996 4718 1043
rect 4776 1043 4984 1060
rect 5368 1060 5384 1077
rect 5826 1077 6242 1093
rect 5826 1060 5842 1077
rect 5368 1043 5576 1060
rect 4776 996 5576 1043
rect 5634 1043 5842 1060
rect 6226 1060 6242 1077
rect 6226 1043 6434 1060
rect 5634 996 6434 1043
rect -2088 749 -1288 796
rect -2088 732 -1880 749
rect -1896 715 -1880 732
rect -1496 732 -1288 749
rect -1230 749 -430 796
rect -1230 732 -1022 749
rect -1496 715 -1480 732
rect -1896 699 -1480 715
rect -1038 715 -1022 732
rect -638 732 -430 749
rect -372 749 428 796
rect -372 732 -164 749
rect -638 715 -622 732
rect -1038 699 -622 715
rect -180 715 -164 732
rect 220 732 428 749
rect 486 749 1286 796
rect 486 732 694 749
rect 220 715 236 732
rect -180 699 236 715
rect 678 715 694 732
rect 1078 732 1286 749
rect 1344 749 2144 796
rect 1344 732 1552 749
rect 1078 715 1094 732
rect 678 699 1094 715
rect 1536 715 1552 732
rect 1936 732 2144 749
rect 2202 749 3002 796
rect 2202 732 2410 749
rect 1936 715 1952 732
rect 1536 699 1952 715
rect 2394 715 2410 732
rect 2794 732 3002 749
rect 3060 749 3860 796
rect 3060 732 3268 749
rect 2794 715 2810 732
rect 2394 699 2810 715
rect 3252 715 3268 732
rect 3652 732 3860 749
rect 3918 749 4718 796
rect 3918 732 4126 749
rect 3652 715 3668 732
rect 3252 699 3668 715
rect 4110 715 4126 732
rect 4510 732 4718 749
rect 4776 749 5576 796
rect 4776 732 4984 749
rect 4510 715 4526 732
rect 4110 699 4526 715
rect 4968 715 4984 732
rect 5368 732 5576 749
rect 5634 749 6434 796
rect 5634 732 5842 749
rect 5368 715 5384 732
rect 4968 699 5384 715
rect 5826 715 5842 732
rect 6226 732 6434 749
rect 6226 715 6242 732
rect 5826 699 6242 715
rect -1985 -433 -1955 -407
rect -1901 -433 -1871 -407
rect -1634 -427 -1604 -401
rect -1542 -427 -1512 -401
rect -1443 -427 -1413 -401
rect -1303 -427 -1273 -401
rect -1206 -427 -1176 -401
rect -1009 -427 -979 -401
rect -910 -427 -880 -401
rect -824 -427 -794 -401
rect -740 -427 -710 -401
rect -632 -427 -602 -401
rect -548 -427 -518 -401
rect -384 -427 -354 -401
rect -165 -427 -135 -401
rect -68 -427 -38 -401
rect 172 -427 202 -401
rect 407 -427 437 -401
rect 491 -427 521 -401
rect 730 -427 760 -401
rect 970 -427 1000 -401
rect 1067 -427 1097 -401
rect 1286 -427 1316 -401
rect 1450 -427 1480 -401
rect 1534 -427 1564 -401
rect 1642 -427 1672 -401
rect 1726 -427 1756 -401
rect 1812 -427 1842 -401
rect 1911 -427 1941 -401
rect 2108 -427 2138 -401
rect 2205 -427 2235 -401
rect 2345 -427 2375 -401
rect 2444 -427 2474 -401
rect 2536 -427 2566 -401
rect -1985 -576 -1955 -561
rect -2018 -606 -1955 -576
rect -2018 -659 -1988 -606
rect -1901 -650 -1871 -561
rect -1634 -598 -1604 -511
rect -1542 -549 -1512 -511
rect -2042 -675 -1988 -659
rect -2042 -709 -2032 -675
rect -1998 -709 -1988 -675
rect -1946 -660 -1871 -650
rect -1946 -694 -1930 -660
rect -1896 -694 -1871 -660
rect -1733 -614 -1604 -598
rect -1558 -559 -1492 -549
rect -1558 -593 -1542 -559
rect -1508 -593 -1492 -559
rect -1558 -603 -1492 -593
rect -1733 -648 -1723 -614
rect -1689 -628 -1604 -614
rect -1689 -648 -1616 -628
rect -1443 -645 -1413 -511
rect -1303 -569 -1273 -511
rect -1303 -585 -1248 -569
rect -1303 -619 -1293 -585
rect -1259 -619 -1248 -585
rect -1303 -635 -1248 -619
rect -1733 -664 -1616 -648
rect -1946 -704 -1871 -694
rect -2042 -725 -1988 -709
rect -2018 -748 -1988 -725
rect -2018 -778 -1955 -748
rect -1985 -793 -1955 -778
rect -1901 -793 -1871 -704
rect -1646 -793 -1616 -664
rect -1551 -675 -1413 -645
rect -1551 -705 -1520 -675
rect -1574 -721 -1520 -705
rect -1574 -755 -1564 -721
rect -1530 -755 -1520 -721
rect -1574 -771 -1520 -755
rect -1478 -727 -1412 -717
rect -1478 -761 -1462 -727
rect -1428 -761 -1412 -727
rect -1478 -771 -1412 -761
rect -1551 -805 -1521 -771
rect -1455 -805 -1425 -771
rect -1289 -793 -1259 -635
rect -1206 -705 -1176 -511
rect -1009 -610 -979 -595
rect -1085 -640 -979 -610
rect -1085 -657 -1055 -640
rect -1121 -673 -1055 -657
rect -1217 -721 -1163 -705
rect -1217 -755 -1207 -721
rect -1173 -755 -1163 -721
rect -1121 -707 -1111 -673
rect -1077 -707 -1055 -673
rect -910 -645 -880 -511
rect -824 -543 -794 -511
rect -838 -559 -784 -543
rect -838 -593 -828 -559
rect -794 -593 -784 -559
rect -838 -609 -784 -593
rect -910 -657 -860 -645
rect -910 -669 -847 -657
rect -910 -675 -823 -669
rect -889 -685 -823 -675
rect -889 -687 -867 -685
rect -1121 -723 -1055 -707
rect -1085 -749 -1055 -723
rect -986 -733 -919 -717
rect -1217 -771 -1163 -755
rect -1217 -793 -1187 -771
rect -986 -767 -963 -733
rect -929 -767 -919 -733
rect -986 -783 -919 -767
rect -877 -719 -867 -687
rect -833 -719 -823 -685
rect -877 -735 -823 -719
rect -740 -695 -710 -511
rect -632 -667 -602 -511
rect -548 -559 -518 -511
rect -560 -575 -506 -559
rect -560 -609 -550 -575
rect -516 -609 -506 -575
rect -560 -625 -506 -609
rect -637 -683 -583 -667
rect -740 -711 -679 -695
rect -740 -731 -723 -711
rect -986 -805 -956 -783
rect -877 -805 -847 -735
rect -781 -745 -723 -731
rect -689 -745 -679 -711
rect -637 -717 -627 -683
rect -593 -717 -583 -683
rect -637 -733 -583 -717
rect -781 -761 -679 -745
rect -781 -793 -751 -761
rect -632 -793 -602 -733
rect -541 -793 -511 -625
rect -165 -591 -135 -555
rect -176 -621 -135 -591
rect -384 -659 -354 -627
rect -176 -659 -146 -621
rect 1067 -591 1097 -555
rect 1067 -621 1108 -591
rect -68 -659 -38 -627
rect 172 -659 202 -627
rect 407 -659 437 -627
rect -455 -675 -146 -659
rect -455 -709 -427 -675
rect -393 -709 -146 -675
rect -455 -725 -146 -709
rect -97 -675 -38 -659
rect -97 -709 -87 -675
rect -53 -709 -38 -675
rect -97 -725 -38 -709
rect 116 -675 202 -659
rect 116 -709 132 -675
rect 166 -709 202 -675
rect 116 -725 202 -709
rect 349 -675 437 -659
rect 349 -709 366 -675
rect 400 -709 437 -675
rect 349 -725 437 -709
rect -353 -747 -323 -725
rect -176 -748 -146 -725
rect -68 -747 -38 -725
rect 172 -747 202 -725
rect 407 -747 437 -725
rect 491 -659 521 -627
rect 730 -659 760 -627
rect 970 -659 1000 -627
rect 1078 -659 1108 -621
rect 1450 -559 1480 -511
rect 1438 -575 1492 -559
rect 1438 -609 1448 -575
rect 1482 -609 1492 -575
rect 1438 -625 1492 -609
rect 1286 -659 1316 -627
rect 491 -675 583 -659
rect 491 -709 534 -675
rect 568 -709 583 -675
rect 491 -725 583 -709
rect 730 -675 816 -659
rect 730 -709 766 -675
rect 800 -709 816 -675
rect 730 -725 816 -709
rect 970 -675 1029 -659
rect 970 -709 985 -675
rect 1019 -709 1029 -675
rect 970 -725 1029 -709
rect 1078 -675 1387 -659
rect 1078 -709 1325 -675
rect 1359 -709 1387 -675
rect 1078 -725 1387 -709
rect 491 -747 521 -725
rect 730 -747 760 -725
rect 970 -747 1000 -725
rect -176 -778 -135 -748
rect -165 -793 -135 -778
rect 1078 -748 1108 -725
rect 1255 -747 1285 -725
rect 1067 -778 1108 -748
rect 1067 -793 1097 -778
rect 1443 -793 1473 -625
rect 1534 -667 1564 -511
rect 1515 -683 1569 -667
rect 1515 -717 1525 -683
rect 1559 -717 1569 -683
rect 1642 -695 1672 -511
rect 1726 -543 1756 -511
rect 1716 -559 1770 -543
rect 1716 -593 1726 -559
rect 1760 -593 1770 -559
rect 1716 -609 1770 -593
rect 1812 -645 1842 -511
rect 2803 -433 2833 -407
rect 2887 -433 2917 -407
rect 1911 -610 1941 -595
rect 1911 -640 2017 -610
rect 1792 -657 1842 -645
rect 1779 -669 1842 -657
rect 1515 -733 1569 -717
rect 1611 -711 1672 -695
rect 1534 -793 1564 -733
rect 1611 -745 1621 -711
rect 1655 -731 1672 -711
rect 1755 -675 1842 -669
rect 1987 -657 2017 -640
rect 1987 -673 2053 -657
rect 1755 -685 1821 -675
rect 1755 -719 1765 -685
rect 1799 -687 1821 -685
rect 1799 -719 1809 -687
rect 1987 -707 2009 -673
rect 2043 -707 2053 -673
rect 2108 -705 2138 -511
rect 2205 -569 2235 -511
rect 2180 -585 2235 -569
rect 2180 -619 2191 -585
rect 2225 -619 2235 -585
rect 2180 -635 2235 -619
rect 1655 -745 1713 -731
rect 1755 -735 1809 -719
rect 1611 -761 1713 -745
rect 1683 -793 1713 -761
rect 1779 -805 1809 -735
rect 1851 -733 1918 -717
rect 1851 -767 1861 -733
rect 1895 -767 1918 -733
rect 1987 -723 2053 -707
rect 2095 -721 2149 -705
rect 1987 -749 2017 -723
rect 1851 -783 1918 -767
rect 1888 -805 1918 -783
rect 2095 -755 2105 -721
rect 2139 -755 2149 -721
rect 2095 -771 2149 -755
rect 2119 -793 2149 -771
rect 2191 -793 2221 -635
rect 2345 -645 2375 -511
rect 2444 -549 2474 -511
rect 2424 -559 2490 -549
rect 2424 -593 2440 -559
rect 2474 -593 2490 -559
rect 2424 -603 2490 -593
rect 2536 -598 2566 -511
rect 3469 37 3601 53
rect 3469 20 3485 37
rect 3435 3 3485 20
rect 3585 20 3601 37
rect 3727 37 3859 53
rect 3727 20 3743 37
rect 3585 3 3635 20
rect 3435 -44 3635 3
rect 3693 3 3743 20
rect 3843 20 3859 37
rect 3985 37 4117 53
rect 3985 20 4001 37
rect 3843 3 3893 20
rect 3693 -44 3893 3
rect 3951 3 4001 20
rect 4101 20 4117 37
rect 4243 37 4375 53
rect 4243 20 4259 37
rect 4101 3 4151 20
rect 3951 -44 4151 3
rect 4209 3 4259 20
rect 4359 20 4375 37
rect 4501 37 4633 53
rect 4501 20 4517 37
rect 4359 3 4409 20
rect 4209 -44 4409 3
rect 4467 3 4517 20
rect 4617 20 4633 37
rect 4759 37 4891 53
rect 4759 20 4775 37
rect 4617 3 4667 20
rect 4467 -44 4667 3
rect 4725 3 4775 20
rect 4875 20 4891 37
rect 4875 3 4925 20
rect 4725 -44 4925 3
rect 3435 -491 3635 -444
rect 3435 -508 3485 -491
rect 2536 -614 2665 -598
rect 2536 -628 2621 -614
rect 2345 -675 2483 -645
rect 2452 -705 2483 -675
rect 2548 -648 2621 -628
rect 2655 -648 2665 -614
rect 2548 -664 2665 -648
rect 2803 -650 2833 -561
rect 2887 -576 2917 -561
rect 2887 -606 2950 -576
rect 2803 -660 2878 -650
rect 2344 -727 2410 -717
rect 2344 -761 2360 -727
rect 2394 -761 2410 -727
rect 2344 -771 2410 -761
rect 2452 -721 2506 -705
rect 2452 -755 2462 -721
rect 2496 -755 2506 -721
rect 2452 -771 2506 -755
rect 2357 -805 2387 -771
rect 2453 -805 2483 -771
rect 2548 -793 2578 -664
rect 2803 -694 2828 -660
rect 2862 -694 2878 -660
rect 2803 -704 2878 -694
rect 2920 -659 2950 -606
rect 3469 -525 3485 -508
rect 3585 -508 3635 -491
rect 3693 -491 3893 -444
rect 3693 -508 3743 -491
rect 3585 -525 3601 -508
rect 3469 -541 3601 -525
rect 3727 -525 3743 -508
rect 3843 -508 3893 -491
rect 3951 -491 4151 -444
rect 3951 -508 4001 -491
rect 3843 -525 3859 -508
rect 3727 -541 3859 -525
rect 3985 -525 4001 -508
rect 4101 -508 4151 -491
rect 4209 -491 4409 -444
rect 4209 -508 4259 -491
rect 4101 -525 4117 -508
rect 3985 -541 4117 -525
rect 4243 -525 4259 -508
rect 4359 -508 4409 -491
rect 4467 -491 4667 -444
rect 4467 -508 4517 -491
rect 4359 -525 4375 -508
rect 4243 -541 4375 -525
rect 4501 -525 4517 -508
rect 4617 -508 4667 -491
rect 4725 -491 4925 -444
rect 4725 -508 4775 -491
rect 4617 -525 4633 -508
rect 4501 -541 4633 -525
rect 4759 -525 4775 -508
rect 4875 -508 4925 -491
rect 4875 -525 4891 -508
rect 4759 -541 4891 -525
rect 5365 37 5497 53
rect 5365 20 5381 37
rect 5331 3 5381 20
rect 5481 20 5497 37
rect 5623 37 5755 53
rect 5623 20 5639 37
rect 5481 3 5531 20
rect 5331 -44 5531 3
rect 5589 3 5639 20
rect 5739 20 5755 37
rect 5881 37 6013 53
rect 5881 20 5897 37
rect 5739 3 5789 20
rect 5589 -44 5789 3
rect 5847 3 5897 20
rect 5997 20 6013 37
rect 5997 3 6047 20
rect 5847 -44 6047 3
rect 5331 -491 5531 -444
rect 5331 -508 5381 -491
rect 5365 -525 5381 -508
rect 5481 -508 5531 -491
rect 5589 -491 5789 -444
rect 5589 -508 5639 -491
rect 5481 -525 5497 -508
rect 5365 -541 5497 -525
rect 5623 -525 5639 -508
rect 5739 -508 5789 -491
rect 5847 -491 6047 -444
rect 5847 -508 5897 -491
rect 5739 -525 5755 -508
rect 5623 -541 5755 -525
rect 5881 -525 5897 -508
rect 5997 -508 6047 -491
rect 5997 -525 6013 -508
rect 5881 -541 6013 -525
rect 2920 -675 2974 -659
rect 2803 -793 2833 -704
rect 2920 -709 2930 -675
rect 2964 -709 2974 -675
rect 2920 -725 2974 -709
rect 2920 -748 2950 -725
rect 2887 -778 2950 -748
rect 2887 -793 2917 -778
rect -1985 -903 -1955 -877
rect -1901 -903 -1871 -877
rect -1646 -903 -1616 -877
rect -1551 -903 -1521 -877
rect -1455 -903 -1425 -877
rect -1289 -903 -1259 -877
rect -1217 -903 -1187 -877
rect -1085 -903 -1055 -877
rect -986 -903 -956 -877
rect -877 -903 -847 -877
rect -781 -903 -751 -877
rect -632 -903 -602 -877
rect -541 -903 -511 -877
rect -353 -903 -323 -877
rect -165 -903 -135 -877
rect -68 -903 -38 -877
rect 172 -903 202 -877
rect 407 -903 437 -877
rect 491 -903 521 -877
rect 730 -903 760 -877
rect 970 -903 1000 -877
rect 1067 -903 1097 -877
rect 1255 -903 1285 -877
rect 1443 -903 1473 -877
rect 1534 -903 1564 -877
rect 1683 -903 1713 -877
rect 1779 -903 1809 -877
rect 1888 -903 1918 -877
rect 1987 -903 2017 -877
rect 2119 -903 2149 -877
rect 2191 -903 2221 -877
rect 2357 -903 2387 -877
rect 2453 -903 2483 -877
rect 2548 -903 2578 -877
rect 2803 -903 2833 -877
rect 2887 -903 2917 -877
rect 3469 -859 3601 -843
rect 3469 -876 3485 -859
rect 3435 -893 3485 -876
rect 3585 -876 3601 -859
rect 3727 -859 3859 -843
rect 3727 -876 3743 -859
rect 3585 -893 3635 -876
rect 3435 -931 3635 -893
rect 3693 -893 3743 -876
rect 3843 -876 3859 -859
rect 3985 -859 4117 -843
rect 3985 -876 4001 -859
rect 3843 -893 3893 -876
rect 3693 -931 3893 -893
rect 3951 -893 4001 -876
rect 4101 -876 4117 -859
rect 4243 -859 4375 -843
rect 4243 -876 4259 -859
rect 4101 -893 4151 -876
rect 3951 -931 4151 -893
rect 4209 -893 4259 -876
rect 4359 -876 4375 -859
rect 4501 -859 4633 -843
rect 4501 -876 4517 -859
rect 4359 -893 4409 -876
rect 4209 -931 4409 -893
rect 4467 -893 4517 -876
rect 4617 -876 4633 -859
rect 4759 -859 4891 -843
rect 4759 -876 4775 -859
rect 4617 -893 4667 -876
rect 4467 -931 4667 -893
rect 4725 -893 4775 -876
rect 4875 -876 4891 -859
rect 4875 -893 4925 -876
rect 4725 -931 4925 -893
rect 3435 -1169 3635 -1131
rect 3435 -1186 3485 -1169
rect 3469 -1203 3485 -1186
rect 3585 -1186 3635 -1169
rect 3693 -1169 3893 -1131
rect 3693 -1186 3743 -1169
rect 3585 -1203 3601 -1186
rect 3469 -1219 3601 -1203
rect 3727 -1203 3743 -1186
rect 3843 -1186 3893 -1169
rect 3951 -1169 4151 -1131
rect 3951 -1186 4001 -1169
rect 3843 -1203 3859 -1186
rect 3727 -1219 3859 -1203
rect 3985 -1203 4001 -1186
rect 4101 -1186 4151 -1169
rect 4209 -1169 4409 -1131
rect 4209 -1186 4259 -1169
rect 4101 -1203 4117 -1186
rect 3985 -1219 4117 -1203
rect 4243 -1203 4259 -1186
rect 4359 -1186 4409 -1169
rect 4467 -1169 4667 -1131
rect 4467 -1186 4517 -1169
rect 4359 -1203 4375 -1186
rect 4243 -1219 4375 -1203
rect 4501 -1203 4517 -1186
rect 4617 -1186 4667 -1169
rect 4725 -1169 4925 -1131
rect 4725 -1186 4775 -1169
rect 4617 -1203 4633 -1186
rect 4501 -1219 4633 -1203
rect 4759 -1203 4775 -1186
rect 4875 -1186 4925 -1169
rect 4875 -1203 4891 -1186
rect 4759 -1219 4891 -1203
rect 5365 -859 5497 -843
rect 5365 -876 5381 -859
rect 5331 -893 5381 -876
rect 5481 -876 5497 -859
rect 5623 -859 5755 -843
rect 5623 -876 5639 -859
rect 5481 -893 5531 -876
rect 5331 -931 5531 -893
rect 5589 -893 5639 -876
rect 5739 -876 5755 -859
rect 5881 -859 6013 -843
rect 5881 -876 5897 -859
rect 5739 -893 5789 -876
rect 5589 -931 5789 -893
rect 5847 -893 5897 -876
rect 5997 -876 6013 -859
rect 5997 -893 6047 -876
rect 5847 -931 6047 -893
rect 5331 -1169 5531 -1131
rect 5331 -1186 5381 -1169
rect 5365 -1203 5381 -1186
rect 5481 -1186 5531 -1169
rect 5589 -1169 5789 -1131
rect 5589 -1186 5639 -1169
rect 5481 -1203 5497 -1186
rect 5365 -1219 5497 -1203
rect 5623 -1203 5639 -1186
rect 5739 -1186 5789 -1169
rect 5847 -1169 6047 -1131
rect 5847 -1186 5897 -1169
rect 5739 -1203 5755 -1186
rect 5623 -1219 5755 -1203
rect 5881 -1203 5897 -1186
rect 5997 -1186 6047 -1169
rect 5997 -1203 6013 -1186
rect 5881 -1219 6013 -1203
rect -1550 -1912 -1058 -1896
rect -1550 -1929 -1534 -1912
rect -1704 -1946 -1534 -1929
rect -1074 -1929 -1058 -1912
rect -692 -1912 -200 -1896
rect -692 -1929 -676 -1912
rect -1074 -1946 -904 -1929
rect -1704 -1984 -904 -1946
rect -846 -1946 -676 -1929
rect -216 -1929 -200 -1912
rect 166 -1912 658 -1896
rect 166 -1929 182 -1912
rect -216 -1946 -46 -1929
rect -846 -1984 -46 -1946
rect 12 -1946 182 -1929
rect 642 -1929 658 -1912
rect 1024 -1912 1516 -1896
rect 1024 -1929 1040 -1912
rect 642 -1946 812 -1929
rect 12 -1984 812 -1946
rect 870 -1946 1040 -1929
rect 1500 -1929 1516 -1912
rect 1882 -1912 2374 -1896
rect 1882 -1929 1898 -1912
rect 1500 -1946 1670 -1929
rect 870 -1984 1670 -1946
rect 1728 -1946 1898 -1929
rect 2358 -1929 2374 -1912
rect 2740 -1912 3232 -1896
rect 2740 -1929 2756 -1912
rect 2358 -1946 2528 -1929
rect 1728 -1984 2528 -1946
rect 2586 -1946 2756 -1929
rect 3216 -1929 3232 -1912
rect 3598 -1912 4090 -1896
rect 3598 -1929 3614 -1912
rect 3216 -1946 3386 -1929
rect 2586 -1984 3386 -1946
rect 3444 -1946 3614 -1929
rect 4074 -1929 4090 -1912
rect 4456 -1912 4948 -1896
rect 4456 -1929 4472 -1912
rect 4074 -1946 4244 -1929
rect 3444 -1984 4244 -1946
rect 4302 -1946 4472 -1929
rect 4932 -1929 4948 -1912
rect 5314 -1912 5806 -1896
rect 5314 -1929 5330 -1912
rect 4932 -1946 5102 -1929
rect 4302 -1984 5102 -1946
rect 5160 -1946 5330 -1929
rect 5790 -1929 5806 -1912
rect 5790 -1946 5960 -1929
rect 5160 -1984 5960 -1946
rect -1704 -2222 -904 -2184
rect -1704 -2239 -1534 -2222
rect -1550 -2256 -1534 -2239
rect -1074 -2239 -904 -2222
rect -846 -2222 -46 -2184
rect -846 -2239 -676 -2222
rect -1074 -2256 -1058 -2239
rect -1550 -2272 -1058 -2256
rect -692 -2256 -676 -2239
rect -216 -2239 -46 -2222
rect 12 -2222 812 -2184
rect 12 -2239 182 -2222
rect -216 -2256 -200 -2239
rect -692 -2272 -200 -2256
rect 166 -2256 182 -2239
rect 642 -2239 812 -2222
rect 870 -2222 1670 -2184
rect 870 -2239 1040 -2222
rect 642 -2256 658 -2239
rect 166 -2272 658 -2256
rect 1024 -2256 1040 -2239
rect 1500 -2239 1670 -2222
rect 1728 -2222 2528 -2184
rect 1728 -2239 1898 -2222
rect 1500 -2256 1516 -2239
rect 1024 -2272 1516 -2256
rect 1882 -2256 1898 -2239
rect 2358 -2239 2528 -2222
rect 2586 -2222 3386 -2184
rect 2586 -2239 2756 -2222
rect 2358 -2256 2374 -2239
rect 1882 -2272 2374 -2256
rect 2740 -2256 2756 -2239
rect 3216 -2239 3386 -2222
rect 3444 -2222 4244 -2184
rect 3444 -2239 3614 -2222
rect 3216 -2256 3232 -2239
rect 2740 -2272 3232 -2256
rect 3598 -2256 3614 -2239
rect 4074 -2239 4244 -2222
rect 4302 -2222 5102 -2184
rect 4302 -2239 4472 -2222
rect 4074 -2256 4090 -2239
rect 3598 -2272 4090 -2256
rect 4456 -2256 4472 -2239
rect 4932 -2239 5102 -2222
rect 5160 -2222 5960 -2184
rect 5160 -2239 5330 -2222
rect 4932 -2256 4948 -2239
rect 4456 -2272 4948 -2256
rect 5314 -2256 5330 -2239
rect 5790 -2239 5960 -2222
rect 5790 -2256 5806 -2239
rect 5314 -2272 5806 -2256
rect -1550 -2494 -1058 -2478
rect -1550 -2511 -1534 -2494
rect -1704 -2528 -1534 -2511
rect -1074 -2511 -1058 -2494
rect -692 -2494 -200 -2478
rect -692 -2511 -676 -2494
rect -1074 -2528 -904 -2511
rect -1704 -2566 -904 -2528
rect -846 -2528 -676 -2511
rect -216 -2511 -200 -2494
rect 166 -2494 658 -2478
rect 166 -2511 182 -2494
rect -216 -2528 -46 -2511
rect -846 -2566 -46 -2528
rect 12 -2528 182 -2511
rect 642 -2511 658 -2494
rect 1024 -2494 1516 -2478
rect 1024 -2511 1040 -2494
rect 642 -2528 812 -2511
rect 12 -2566 812 -2528
rect 870 -2528 1040 -2511
rect 1500 -2511 1516 -2494
rect 1882 -2494 2374 -2478
rect 1882 -2511 1898 -2494
rect 1500 -2528 1670 -2511
rect 870 -2566 1670 -2528
rect 1728 -2528 1898 -2511
rect 2358 -2511 2374 -2494
rect 2740 -2494 3232 -2478
rect 2740 -2511 2756 -2494
rect 2358 -2528 2528 -2511
rect 1728 -2566 2528 -2528
rect 2586 -2528 2756 -2511
rect 3216 -2511 3232 -2494
rect 3598 -2494 4090 -2478
rect 3598 -2511 3614 -2494
rect 3216 -2528 3386 -2511
rect 2586 -2566 3386 -2528
rect 3444 -2528 3614 -2511
rect 4074 -2511 4090 -2494
rect 4456 -2494 4948 -2478
rect 4456 -2511 4472 -2494
rect 4074 -2528 4244 -2511
rect 3444 -2566 4244 -2528
rect 4302 -2528 4472 -2511
rect 4932 -2511 4948 -2494
rect 5314 -2494 5806 -2478
rect 5314 -2511 5330 -2494
rect 4932 -2528 5102 -2511
rect 4302 -2566 5102 -2528
rect 5160 -2528 5330 -2511
rect 5790 -2511 5806 -2494
rect 5790 -2528 5960 -2511
rect 5160 -2566 5960 -2528
rect -1704 -2804 -904 -2766
rect -1704 -2821 -1534 -2804
rect -1550 -2838 -1534 -2821
rect -1074 -2821 -904 -2804
rect -846 -2804 -46 -2766
rect -846 -2821 -676 -2804
rect -1074 -2838 -1058 -2821
rect -1550 -2854 -1058 -2838
rect -692 -2838 -676 -2821
rect -216 -2821 -46 -2804
rect 12 -2804 812 -2766
rect 12 -2821 182 -2804
rect -216 -2838 -200 -2821
rect -692 -2854 -200 -2838
rect 166 -2838 182 -2821
rect 642 -2821 812 -2804
rect 870 -2804 1670 -2766
rect 870 -2821 1040 -2804
rect 642 -2838 658 -2821
rect 166 -2854 658 -2838
rect 1024 -2838 1040 -2821
rect 1500 -2821 1670 -2804
rect 1728 -2804 2528 -2766
rect 1728 -2821 1898 -2804
rect 1500 -2838 1516 -2821
rect 1024 -2854 1516 -2838
rect 1882 -2838 1898 -2821
rect 2358 -2821 2528 -2804
rect 2586 -2804 3386 -2766
rect 2586 -2821 2756 -2804
rect 2358 -2838 2374 -2821
rect 1882 -2854 2374 -2838
rect 2740 -2838 2756 -2821
rect 3216 -2821 3386 -2804
rect 3444 -2804 4244 -2766
rect 3444 -2821 3614 -2804
rect 3216 -2838 3232 -2821
rect 2740 -2854 3232 -2838
rect 3598 -2838 3614 -2821
rect 4074 -2821 4244 -2804
rect 4302 -2804 5102 -2766
rect 4302 -2821 4472 -2804
rect 4074 -2838 4090 -2821
rect 3598 -2854 4090 -2838
rect 4456 -2838 4472 -2821
rect 4932 -2821 5102 -2804
rect 5160 -2804 5960 -2766
rect 5160 -2821 5330 -2804
rect 4932 -2838 4948 -2821
rect 4456 -2854 4948 -2838
rect 5314 -2838 5330 -2821
rect 5790 -2821 5960 -2804
rect 5790 -2838 5806 -2821
rect 5314 -2854 5806 -2838
<< polycont >>
rect -1880 1643 -1496 1677
rect -1022 1643 -638 1677
rect -164 1643 220 1677
rect 694 1643 1078 1677
rect 1552 1643 1936 1677
rect 2410 1643 2794 1677
rect 3268 1643 3652 1677
rect 4126 1643 4510 1677
rect 4984 1643 5368 1677
rect 5842 1643 6226 1677
rect -1880 1315 -1496 1349
rect -1022 1315 -638 1349
rect -164 1315 220 1349
rect 694 1315 1078 1349
rect 1552 1315 1936 1349
rect 2410 1315 2794 1349
rect 3268 1315 3652 1349
rect 4126 1315 4510 1349
rect 4984 1315 5368 1349
rect 5842 1315 6226 1349
rect -1880 1043 -1496 1077
rect -1022 1043 -638 1077
rect -164 1043 220 1077
rect 694 1043 1078 1077
rect 1552 1043 1936 1077
rect 2410 1043 2794 1077
rect 3268 1043 3652 1077
rect 4126 1043 4510 1077
rect 4984 1043 5368 1077
rect 5842 1043 6226 1077
rect -1880 715 -1496 749
rect -1022 715 -638 749
rect -164 715 220 749
rect 694 715 1078 749
rect 1552 715 1936 749
rect 2410 715 2794 749
rect 3268 715 3652 749
rect 4126 715 4510 749
rect 4984 715 5368 749
rect 5842 715 6226 749
rect -2032 -709 -1998 -675
rect -1930 -694 -1896 -660
rect -1542 -593 -1508 -559
rect -1723 -648 -1689 -614
rect -1293 -619 -1259 -585
rect -1564 -755 -1530 -721
rect -1462 -761 -1428 -727
rect -1207 -755 -1173 -721
rect -1111 -707 -1077 -673
rect -828 -593 -794 -559
rect -963 -767 -929 -733
rect -867 -719 -833 -685
rect -550 -609 -516 -575
rect -723 -745 -689 -711
rect -627 -717 -593 -683
rect -427 -709 -393 -675
rect -87 -709 -53 -675
rect 132 -709 166 -675
rect 366 -709 400 -675
rect 1448 -609 1482 -575
rect 534 -709 568 -675
rect 766 -709 800 -675
rect 985 -709 1019 -675
rect 1325 -709 1359 -675
rect 1525 -717 1559 -683
rect 1726 -593 1760 -559
rect 1621 -745 1655 -711
rect 1765 -719 1799 -685
rect 2009 -707 2043 -673
rect 2191 -619 2225 -585
rect 1861 -767 1895 -733
rect 2105 -755 2139 -721
rect 2440 -593 2474 -559
rect 3485 3 3585 37
rect 3743 3 3843 37
rect 4001 3 4101 37
rect 4259 3 4359 37
rect 4517 3 4617 37
rect 4775 3 4875 37
rect 2621 -648 2655 -614
rect 2360 -761 2394 -727
rect 2462 -755 2496 -721
rect 2828 -694 2862 -660
rect 3485 -525 3585 -491
rect 3743 -525 3843 -491
rect 4001 -525 4101 -491
rect 4259 -525 4359 -491
rect 4517 -525 4617 -491
rect 4775 -525 4875 -491
rect 5381 3 5481 37
rect 5639 3 5739 37
rect 5897 3 5997 37
rect 5381 -525 5481 -491
rect 5639 -525 5739 -491
rect 5897 -525 5997 -491
rect 2930 -709 2964 -675
rect 3485 -893 3585 -859
rect 3743 -893 3843 -859
rect 4001 -893 4101 -859
rect 4259 -893 4359 -859
rect 4517 -893 4617 -859
rect 4775 -893 4875 -859
rect 3485 -1203 3585 -1169
rect 3743 -1203 3843 -1169
rect 4001 -1203 4101 -1169
rect 4259 -1203 4359 -1169
rect 4517 -1203 4617 -1169
rect 4775 -1203 4875 -1169
rect 5381 -893 5481 -859
rect 5639 -893 5739 -859
rect 5897 -893 5997 -859
rect 5381 -1203 5481 -1169
rect 5639 -1203 5739 -1169
rect 5897 -1203 5997 -1169
rect -1534 -1946 -1074 -1912
rect -676 -1946 -216 -1912
rect 182 -1946 642 -1912
rect 1040 -1946 1500 -1912
rect 1898 -1946 2358 -1912
rect 2756 -1946 3216 -1912
rect 3614 -1946 4074 -1912
rect 4472 -1946 4932 -1912
rect 5330 -1946 5790 -1912
rect -1534 -2256 -1074 -2222
rect -676 -2256 -216 -2222
rect 182 -2256 642 -2222
rect 1040 -2256 1500 -2222
rect 1898 -2256 2358 -2222
rect 2756 -2256 3216 -2222
rect 3614 -2256 4074 -2222
rect 4472 -2256 4932 -2222
rect 5330 -2256 5790 -2222
rect -1534 -2528 -1074 -2494
rect -676 -2528 -216 -2494
rect 182 -2528 642 -2494
rect 1040 -2528 1500 -2494
rect 1898 -2528 2358 -2494
rect 2756 -2528 3216 -2494
rect 3614 -2528 4074 -2494
rect 4472 -2528 4932 -2494
rect 5330 -2528 5790 -2494
rect -1534 -2838 -1074 -2804
rect -676 -2838 -216 -2804
rect 182 -2838 642 -2804
rect 1040 -2838 1500 -2804
rect 1898 -2838 2358 -2804
rect 2756 -2838 3216 -2804
rect 3614 -2838 4074 -2804
rect 4472 -2838 4932 -2804
rect 5330 -2838 5790 -2804
<< locali >>
rect -2522 2500 -2422 2662
rect 6822 2500 6922 2662
rect -1896 1643 -1880 1677
rect -1496 1643 -1480 1677
rect -1038 1643 -1022 1677
rect -638 1643 -622 1677
rect -180 1643 -164 1677
rect 220 1643 236 1677
rect 678 1643 694 1677
rect 1078 1643 1094 1677
rect 1536 1643 1552 1677
rect 1936 1643 1952 1677
rect 2394 1643 2410 1677
rect 2794 1643 2810 1677
rect 3252 1643 3268 1677
rect 3652 1643 3668 1677
rect 4110 1643 4126 1677
rect 4510 1643 4526 1677
rect 4968 1643 4984 1677
rect 5368 1643 5384 1677
rect 5826 1643 5842 1677
rect 6226 1643 6242 1677
rect -2134 1584 -2100 1600
rect -2134 1392 -2100 1408
rect -1276 1584 -1242 1600
rect -1276 1392 -1242 1408
rect -418 1584 -384 1600
rect -418 1392 -384 1408
rect 440 1584 474 1600
rect 440 1392 474 1408
rect 1298 1584 1332 1600
rect 1298 1392 1332 1408
rect 2156 1584 2190 1600
rect 2156 1392 2190 1408
rect 3014 1584 3048 1600
rect 3014 1392 3048 1408
rect 3872 1584 3906 1600
rect 3872 1392 3906 1408
rect 4730 1584 4764 1600
rect 4730 1392 4764 1408
rect 5588 1584 5622 1600
rect 5588 1392 5622 1408
rect 6446 1584 6480 1600
rect 6446 1392 6480 1408
rect -1896 1315 -1880 1349
rect -1496 1315 -1480 1349
rect -1038 1315 -1022 1349
rect -638 1315 -622 1349
rect -180 1315 -164 1349
rect 220 1315 236 1349
rect 678 1315 694 1349
rect 1078 1315 1094 1349
rect 1536 1315 1552 1349
rect 1936 1315 1952 1349
rect 2394 1315 2410 1349
rect 2794 1315 2810 1349
rect 3252 1315 3268 1349
rect 3652 1315 3668 1349
rect 4110 1315 4126 1349
rect 4510 1315 4526 1349
rect 4968 1315 4984 1349
rect 5368 1315 5384 1349
rect 5826 1315 5842 1349
rect 6226 1315 6242 1349
rect -1896 1043 -1880 1077
rect -1496 1043 -1480 1077
rect -1038 1043 -1022 1077
rect -638 1043 -622 1077
rect -180 1043 -164 1077
rect 220 1043 236 1077
rect 678 1043 694 1077
rect 1078 1043 1094 1077
rect 1536 1043 1552 1077
rect 1936 1043 1952 1077
rect 2394 1043 2410 1077
rect 2794 1043 2810 1077
rect 3252 1043 3268 1077
rect 3652 1043 3668 1077
rect 4110 1043 4126 1077
rect 4510 1043 4526 1077
rect 4968 1043 4984 1077
rect 5368 1043 5384 1077
rect 5826 1043 5842 1077
rect 6226 1043 6242 1077
rect -2134 984 -2100 1000
rect -2134 792 -2100 808
rect -1276 984 -1242 1000
rect -1276 792 -1242 808
rect -418 984 -384 1000
rect -418 792 -384 808
rect 440 984 474 1000
rect 440 792 474 808
rect 1298 984 1332 1000
rect 1298 792 1332 808
rect 2156 984 2190 1000
rect 2156 792 2190 808
rect 3014 984 3048 1000
rect 3014 792 3048 808
rect 3872 984 3906 1000
rect 3872 792 3906 808
rect 4730 984 4764 1000
rect 4730 792 4764 808
rect 5588 984 5622 1000
rect 5588 792 5622 808
rect 6446 984 6480 1000
rect 6446 792 6480 808
rect -1896 715 -1880 749
rect -1496 715 -1480 749
rect -1038 715 -1022 749
rect -638 715 -622 749
rect -180 715 -164 749
rect 220 715 236 749
rect 678 715 694 749
rect 1078 715 1094 749
rect 1536 715 1552 749
rect 1936 715 1952 749
rect 2394 715 2410 749
rect 2794 715 2810 749
rect 3252 715 3268 749
rect 3652 715 3668 749
rect 4110 715 4126 749
rect 4510 715 4526 749
rect 4968 715 4984 749
rect 5368 715 5384 749
rect 5826 715 5842 749
rect 6226 715 6242 749
rect -2522 358 -2422 520
rect 6822 358 6922 520
rect 3275 105 3371 139
rect 4989 105 5085 139
rect 3275 46 3309 105
rect 3308 43 3309 46
rect 5051 44 5085 105
rect 5171 105 5267 139
rect 6111 105 6207 139
rect 5171 44 5205 105
rect 6173 44 6207 105
rect -2064 -397 -2035 -363
rect -2001 -397 -1943 -363
rect -1909 -397 -1851 -363
rect -1817 -397 -1759 -363
rect -1725 -397 -1667 -363
rect -1633 -397 -1575 -363
rect -1541 -397 -1483 -363
rect -1449 -397 -1391 -363
rect -1357 -397 -1299 -363
rect -1265 -397 -1207 -363
rect -1173 -397 -1115 -363
rect -1081 -397 -1023 -363
rect -989 -397 -931 -363
rect -897 -397 -839 -363
rect -805 -397 -747 -363
rect -713 -397 -655 -363
rect -621 -397 -563 -363
rect -529 -397 -471 -363
rect -437 -397 -379 -363
rect -345 -397 -287 -363
rect -253 -397 -195 -363
rect -161 -397 -103 -363
rect -69 -397 -11 -363
rect 23 -397 81 -363
rect 115 -397 173 -363
rect 207 -397 265 -363
rect 299 -397 357 -363
rect 391 -397 449 -363
rect 483 -397 541 -363
rect 575 -397 633 -363
rect 667 -397 725 -363
rect 759 -397 817 -363
rect 851 -397 909 -363
rect 943 -397 1001 -363
rect 1035 -397 1093 -363
rect 1127 -397 1185 -363
rect 1219 -397 1277 -363
rect 1311 -397 1369 -363
rect 1403 -397 1461 -363
rect 1495 -397 1553 -363
rect 1587 -397 1645 -363
rect 1679 -397 1737 -363
rect 1771 -397 1829 -363
rect 1863 -397 1921 -363
rect 1955 -397 2013 -363
rect 2047 -397 2105 -363
rect 2139 -397 2197 -363
rect 2231 -397 2289 -363
rect 2323 -397 2381 -363
rect 2415 -397 2473 -363
rect 2507 -397 2565 -363
rect 2599 -397 2657 -363
rect 2691 -397 2749 -363
rect 2783 -397 2841 -363
rect 2875 -397 2933 -363
rect 2967 -397 2996 -363
rect -2046 -447 -1995 -431
rect -2046 -481 -2029 -447
rect -2046 -515 -1995 -481
rect -1961 -463 -1895 -397
rect -1961 -497 -1945 -463
rect -1911 -497 -1895 -463
rect -1861 -447 -1827 -431
rect -2046 -549 -2029 -515
rect -1861 -515 -1827 -481
rect -1995 -549 -1896 -531
rect -2046 -565 -1896 -549
rect -2046 -666 -1976 -599
rect -2046 -714 -2044 -666
rect -1996 -714 -1976 -666
rect -2046 -729 -1976 -714
rect -1942 -660 -1896 -565
rect -1942 -669 -1930 -660
rect -1908 -703 -1896 -694
rect -1942 -763 -1896 -703
rect -2046 -797 -1896 -763
rect -2046 -805 -1995 -797
rect -2046 -839 -2029 -805
rect -1861 -805 -1827 -567
rect -1793 -442 -1728 -434
rect -1793 -482 -1782 -442
rect -1736 -482 -1728 -442
rect -1793 -591 -1728 -482
rect -1694 -439 -1644 -397
rect -1694 -473 -1678 -439
rect -1694 -489 -1644 -473
rect -1610 -447 -1560 -431
rect -1610 -481 -1594 -447
rect -1610 -497 -1560 -481
rect -1517 -441 -1381 -431
rect -1517 -475 -1501 -441
rect -1467 -475 -1381 -441
rect -1266 -449 -1200 -397
rect -1073 -439 -999 -397
rect -1517 -497 -1381 -475
rect -1610 -523 -1576 -497
rect -1655 -557 -1576 -523
rect -1542 -533 -1449 -531
rect -1781 -614 -1689 -591
rect -1781 -648 -1723 -614
rect -1781 -801 -1689 -648
rect -2046 -855 -1995 -839
rect -1961 -865 -1945 -831
rect -1911 -865 -1895 -831
rect -1655 -829 -1621 -557
rect -1542 -559 -1483 -533
rect -1508 -567 -1483 -559
rect -1508 -593 -1449 -567
rect -1542 -609 -1449 -593
rect -1587 -669 -1517 -647
rect -1587 -703 -1575 -669
rect -1541 -703 -1517 -669
rect -1587 -721 -1517 -703
rect -1587 -755 -1564 -721
rect -1530 -755 -1517 -721
rect -1587 -771 -1517 -755
rect -1483 -727 -1449 -609
rect -1415 -653 -1381 -497
rect -1347 -465 -1313 -449
rect -1266 -483 -1250 -449
rect -1216 -483 -1200 -449
rect -1166 -465 -1132 -449
rect -1347 -517 -1313 -499
rect -1073 -473 -1053 -439
rect -1019 -473 -999 -439
rect -1073 -489 -999 -473
rect -965 -447 -931 -431
rect -1166 -517 -1132 -499
rect -1347 -551 -1132 -517
rect -965 -523 -931 -481
rect -884 -440 -710 -431
rect -884 -474 -868 -440
rect -834 -474 -710 -440
rect -884 -499 -710 -474
rect -676 -439 -626 -397
rect -642 -473 -626 -439
rect -522 -439 -378 -397
rect -676 -489 -626 -473
rect -592 -465 -558 -449
rect -1043 -557 -931 -523
rect -1043 -585 -1009 -557
rect -1309 -619 -1293 -585
rect -1259 -619 -1009 -585
rect -870 -567 -859 -533
rect -825 -559 -778 -533
rect -870 -591 -828 -567
rect -1415 -673 -1077 -653
rect -1415 -687 -1111 -673
rect -1483 -761 -1462 -727
rect -1428 -761 -1412 -727
rect -1483 -771 -1412 -761
rect -1378 -829 -1344 -687
rect -1303 -737 -1207 -721
rect -1269 -771 -1231 -737
rect -1173 -755 -1145 -721
rect -1111 -723 -1077 -707
rect -1197 -771 -1145 -755
rect -1043 -757 -1009 -619
rect -1861 -855 -1827 -839
rect -1961 -907 -1895 -865
rect -1755 -869 -1739 -835
rect -1705 -869 -1689 -835
rect -1655 -863 -1606 -829
rect -1572 -863 -1556 -829
rect -1515 -863 -1499 -829
rect -1465 -863 -1344 -829
rect -1169 -831 -1103 -815
rect -1755 -907 -1689 -869
rect -1169 -865 -1153 -831
rect -1119 -865 -1103 -831
rect -1169 -907 -1103 -865
rect -1061 -835 -1009 -757
rect -971 -593 -828 -591
rect -794 -593 -778 -559
rect -744 -575 -710 -499
rect -522 -473 -506 -439
rect -472 -473 -428 -439
rect -394 -473 -378 -439
rect -344 -447 -263 -431
rect -112 -439 -78 -397
rect -592 -507 -558 -499
rect -310 -481 -263 -447
rect -592 -541 -432 -507
rect -971 -625 -836 -593
rect -744 -609 -550 -575
rect -516 -609 -500 -575
rect -971 -733 -929 -625
rect -744 -627 -710 -609
rect -971 -767 -963 -733
rect -971 -783 -929 -767
rect -895 -669 -825 -659
rect -895 -685 -859 -669
rect -895 -719 -867 -685
rect -833 -719 -825 -703
rect -895 -783 -825 -719
rect -791 -661 -710 -627
rect -791 -817 -757 -661
rect -643 -674 -535 -643
rect -466 -659 -432 -541
rect -344 -515 -263 -481
rect -310 -549 -263 -515
rect -344 -583 -263 -549
rect -310 -617 -263 -583
rect -344 -633 -263 -617
rect -466 -665 -377 -659
rect -609 -683 -535 -674
rect -723 -711 -679 -695
rect -689 -745 -679 -711
rect -643 -717 -627 -708
rect -593 -717 -535 -683
rect -723 -751 -679 -745
rect -583 -737 -535 -717
rect -723 -785 -617 -751
rect -947 -831 -757 -817
rect -1061 -869 -1041 -835
rect -1007 -869 -991 -835
rect -947 -865 -931 -831
rect -897 -865 -757 -831
rect -947 -873 -757 -865
rect -723 -835 -685 -819
rect -723 -869 -719 -835
rect -651 -831 -617 -785
rect -549 -771 -535 -737
rect -583 -797 -535 -771
rect -501 -675 -377 -665
rect -501 -709 -427 -675
rect -393 -709 -377 -675
rect -501 -725 -377 -709
rect -329 -668 -263 -633
rect -329 -716 -320 -668
rect -272 -716 -263 -668
rect -501 -760 -436 -725
rect -329 -759 -263 -716
rect -501 -815 -437 -760
rect -651 -849 -501 -831
rect -467 -849 -437 -815
rect -651 -865 -437 -849
rect -397 -792 -363 -770
rect -723 -907 -685 -869
rect -397 -907 -363 -826
rect -329 -793 -313 -759
rect -279 -793 -263 -759
rect -329 -827 -263 -793
rect -329 -861 -313 -827
rect -279 -861 -263 -827
rect -225 -473 -209 -439
rect -175 -473 -159 -439
rect -225 -507 -159 -473
rect -225 -541 -209 -507
rect -175 -541 -159 -507
rect -225 -659 -159 -541
rect 120 -439 162 -397
rect -112 -507 -78 -473
rect -112 -575 -78 -541
rect -112 -625 -78 -609
rect -28 -475 23 -459
rect 6 -509 23 -475
rect -28 -543 23 -509
rect 6 -577 23 -543
rect -28 -635 23 -577
rect 120 -473 128 -439
rect 120 -507 162 -473
rect 120 -541 128 -507
rect 120 -575 162 -541
rect 120 -609 128 -575
rect 120 -625 162 -609
rect 196 -439 262 -431
rect 196 -470 212 -439
rect 246 -470 262 -439
rect 196 -518 208 -470
rect 256 -518 262 -470
rect 196 -541 212 -518
rect 246 -541 262 -518
rect 196 -575 262 -541
rect 196 -609 212 -575
rect 246 -609 262 -575
rect 196 -627 262 -609
rect 345 -439 397 -397
rect 345 -473 363 -439
rect 345 -507 397 -473
rect 345 -541 363 -507
rect 345 -575 397 -541
rect 345 -609 363 -575
rect 345 -625 397 -609
rect 431 -439 497 -431
rect 431 -473 447 -439
rect 481 -473 497 -439
rect 431 -507 497 -473
rect 431 -541 447 -507
rect 481 -541 497 -507
rect 431 -570 497 -541
rect 431 -612 444 -570
rect 492 -612 497 -570
rect 431 -627 497 -612
rect 531 -439 587 -397
rect 565 -473 587 -439
rect 531 -507 587 -473
rect 565 -541 587 -507
rect 531 -575 587 -541
rect 565 -609 587 -575
rect 531 -625 587 -609
rect 670 -439 736 -431
rect 670 -473 686 -439
rect 720 -473 736 -439
rect 670 -507 736 -473
rect 670 -541 686 -507
rect 720 -541 736 -507
rect 670 -575 736 -541
rect 670 -609 686 -575
rect 720 -609 736 -575
rect 670 -627 736 -609
rect 770 -439 812 -397
rect 804 -473 812 -439
rect 1010 -439 1044 -397
rect 770 -507 812 -473
rect 804 -541 812 -507
rect 770 -575 812 -541
rect 804 -609 812 -575
rect 770 -625 812 -609
rect 909 -475 960 -459
rect 909 -509 926 -475
rect 909 -543 960 -509
rect 909 -577 926 -543
rect -225 -675 -53 -659
rect -225 -709 -87 -675
rect -225 -725 -53 -709
rect -225 -805 -175 -725
rect -19 -765 23 -635
rect 116 -668 182 -661
rect 116 -708 118 -668
rect 116 -709 132 -708
rect 166 -709 182 -668
rect -28 -781 23 -765
rect -225 -839 -209 -805
rect -225 -855 -175 -839
rect -112 -811 -78 -788
rect -329 -869 -263 -861
rect -112 -907 -78 -845
rect 6 -815 23 -781
rect -28 -871 23 -815
rect 116 -759 162 -743
rect 216 -747 262 -627
rect 349 -668 416 -659
rect 349 -709 352 -668
rect 400 -709 416 -668
rect 450 -747 484 -627
rect 518 -668 585 -659
rect 518 -710 526 -668
rect 574 -710 585 -668
rect 518 -713 585 -710
rect 670 -747 716 -627
rect 909 -635 960 -577
rect 1010 -507 1044 -473
rect 1010 -575 1044 -541
rect 1010 -625 1044 -609
rect 1091 -473 1107 -439
rect 1141 -473 1157 -439
rect 1091 -507 1157 -473
rect 1091 -541 1107 -507
rect 1141 -541 1157 -507
rect 750 -668 816 -661
rect 750 -708 764 -668
rect 812 -708 816 -668
rect 750 -709 766 -708
rect 800 -709 816 -708
rect 116 -793 128 -759
rect 116 -827 162 -793
rect 116 -861 128 -827
rect 116 -907 162 -861
rect 196 -759 262 -747
rect 196 -793 212 -759
rect 246 -793 262 -759
rect 196 -827 262 -793
rect 196 -861 212 -827
rect 246 -861 262 -827
rect 196 -873 262 -861
rect 345 -763 484 -747
rect 345 -797 363 -763
rect 397 -797 484 -763
rect 345 -831 484 -797
rect 345 -865 363 -831
rect 397 -865 484 -831
rect 345 -873 484 -865
rect 525 -763 587 -747
rect 525 -797 531 -763
rect 565 -797 587 -763
rect 525 -831 587 -797
rect 525 -865 531 -831
rect 565 -865 587 -831
rect 525 -907 587 -865
rect 670 -759 736 -747
rect 670 -780 686 -759
rect 720 -780 736 -759
rect 670 -828 676 -780
rect 724 -828 736 -780
rect 670 -861 686 -828
rect 720 -861 736 -828
rect 670 -873 736 -861
rect 770 -759 816 -743
rect 804 -793 816 -759
rect 770 -827 816 -793
rect 804 -861 816 -827
rect 770 -907 816 -861
rect 909 -765 951 -635
rect 1091 -659 1157 -541
rect 985 -675 1157 -659
rect 1019 -709 1157 -675
rect 985 -725 1157 -709
rect 909 -781 960 -765
rect 909 -815 926 -781
rect 909 -871 960 -815
rect 1010 -811 1044 -788
rect 1010 -907 1044 -845
rect 1107 -805 1157 -725
rect 1141 -839 1157 -805
rect 1107 -855 1157 -839
rect 1195 -447 1276 -431
rect 1195 -481 1242 -447
rect 1310 -439 1454 -397
rect 1310 -473 1326 -439
rect 1360 -473 1404 -439
rect 1438 -473 1454 -439
rect 1558 -439 1608 -397
rect 1490 -465 1524 -449
rect 1195 -515 1276 -481
rect 1558 -473 1574 -439
rect 1558 -489 1608 -473
rect 1642 -440 1816 -431
rect 1642 -474 1766 -440
rect 1800 -474 1816 -440
rect 1490 -507 1524 -499
rect 1195 -549 1242 -515
rect 1195 -583 1276 -549
rect 1195 -617 1242 -583
rect 1195 -633 1276 -617
rect 1364 -541 1524 -507
rect 1642 -499 1816 -474
rect 1863 -447 1897 -431
rect 1195 -668 1261 -633
rect 1364 -659 1398 -541
rect 1642 -575 1676 -499
rect 1863 -523 1897 -481
rect 1931 -439 2005 -397
rect 1931 -473 1951 -439
rect 1985 -473 2005 -439
rect 2132 -449 2198 -397
rect 2313 -441 2449 -431
rect 1931 -489 2005 -473
rect 2064 -465 2098 -449
rect 2132 -483 2148 -449
rect 2182 -483 2198 -449
rect 2245 -465 2279 -449
rect 2064 -517 2098 -499
rect 2245 -517 2279 -499
rect 1432 -609 1448 -575
rect 1482 -609 1676 -575
rect 1710 -559 1757 -533
rect 1710 -593 1726 -559
rect 1791 -567 1802 -533
rect 1863 -557 1975 -523
rect 2064 -551 2279 -517
rect 2313 -475 2399 -441
rect 2433 -475 2449 -441
rect 2313 -497 2449 -475
rect 2492 -447 2542 -431
rect 2526 -481 2542 -447
rect 2492 -497 2542 -481
rect 2576 -439 2626 -397
rect 2610 -473 2626 -439
rect 2576 -489 2626 -473
rect 2660 -450 2725 -434
rect 1760 -591 1802 -567
rect 1941 -585 1975 -557
rect 1760 -593 1903 -591
rect 1642 -627 1676 -609
rect 1768 -625 1903 -593
rect 1195 -716 1204 -668
rect 1252 -716 1261 -668
rect 1195 -759 1261 -716
rect 1309 -665 1398 -659
rect 1309 -675 1433 -665
rect 1309 -709 1325 -675
rect 1359 -709 1433 -675
rect 1309 -725 1433 -709
rect 1195 -793 1211 -759
rect 1245 -793 1261 -759
rect 1368 -760 1433 -725
rect 1195 -827 1261 -793
rect 1195 -861 1211 -827
rect 1245 -861 1261 -827
rect 1195 -869 1261 -861
rect 1295 -792 1329 -770
rect 1295 -907 1329 -826
rect 1369 -815 1433 -760
rect 1467 -674 1575 -643
rect 1642 -661 1723 -627
rect 1467 -683 1541 -674
rect 1467 -717 1525 -683
rect 1559 -717 1575 -708
rect 1611 -711 1655 -695
rect 1467 -737 1515 -717
rect 1467 -771 1481 -737
rect 1611 -745 1621 -711
rect 1611 -751 1655 -745
rect 1467 -797 1515 -771
rect 1549 -785 1655 -751
rect 1369 -849 1399 -815
rect 1549 -831 1583 -785
rect 1689 -817 1723 -661
rect 1757 -669 1827 -659
rect 1791 -685 1827 -669
rect 1757 -719 1765 -703
rect 1799 -719 1827 -685
rect 1757 -783 1827 -719
rect 1861 -733 1903 -625
rect 1895 -767 1903 -733
rect 1861 -783 1903 -767
rect 1941 -619 2191 -585
rect 2225 -619 2241 -585
rect 1941 -757 1975 -619
rect 2313 -653 2347 -497
rect 2508 -523 2542 -497
rect 2660 -490 2674 -450
rect 2714 -490 2725 -450
rect 2009 -673 2347 -653
rect 2043 -687 2347 -673
rect 2381 -533 2474 -531
rect 2415 -559 2474 -533
rect 2508 -557 2587 -523
rect 2415 -567 2440 -559
rect 2381 -593 2440 -567
rect 2381 -609 2474 -593
rect 2009 -723 2043 -707
rect 2077 -755 2105 -721
rect 2139 -737 2235 -721
rect 1433 -849 1583 -831
rect 1369 -865 1583 -849
rect 1617 -835 1655 -819
rect 1651 -869 1655 -835
rect 1617 -907 1655 -869
rect 1689 -831 1879 -817
rect 1689 -865 1829 -831
rect 1863 -865 1879 -831
rect 1941 -835 1993 -757
rect 2077 -771 2129 -755
rect 2163 -771 2201 -737
rect 1689 -873 1879 -865
rect 1923 -869 1939 -835
rect 1973 -869 1993 -835
rect 2035 -831 2101 -815
rect 2035 -865 2051 -831
rect 2085 -865 2101 -831
rect 2276 -829 2310 -687
rect 2381 -727 2415 -609
rect 2344 -761 2360 -727
rect 2394 -761 2415 -727
rect 2344 -771 2415 -761
rect 2449 -669 2519 -647
rect 2449 -703 2473 -669
rect 2507 -703 2519 -669
rect 2449 -721 2519 -703
rect 2449 -755 2462 -721
rect 2496 -755 2519 -721
rect 2449 -771 2519 -755
rect 2553 -829 2587 -557
rect 2660 -591 2725 -490
rect 2759 -447 2793 -431
rect 2759 -515 2793 -481
rect 2827 -463 2893 -397
rect 2827 -497 2843 -463
rect 2877 -497 2893 -463
rect 2927 -447 2978 -431
rect 2961 -481 2978 -447
rect 2927 -515 2978 -481
rect 2621 -614 2713 -591
rect 2655 -648 2713 -614
rect 2621 -801 2713 -648
rect 2276 -863 2397 -829
rect 2431 -863 2447 -829
rect 2488 -863 2504 -829
rect 2538 -863 2587 -829
rect 2759 -805 2793 -567
rect 2828 -549 2927 -531
rect 2961 -549 2978 -515
rect 3469 3 3485 37
rect 3585 3 3601 37
rect 3727 3 3743 37
rect 3843 3 3859 37
rect 3985 3 4001 37
rect 4101 3 4117 37
rect 4243 3 4259 37
rect 4359 3 4375 37
rect 4501 3 4517 37
rect 4617 3 4633 37
rect 4759 3 4775 37
rect 4875 3 4891 37
rect 3389 -56 3423 -40
rect 3389 -448 3423 -432
rect 3647 -56 3681 -40
rect 3647 -448 3681 -432
rect 3905 -56 3939 -40
rect 3905 -448 3939 -432
rect 4163 -56 4197 -40
rect 4163 -448 4197 -432
rect 4421 -56 4455 -40
rect 4421 -448 4455 -432
rect 4679 -56 4713 -40
rect 4679 -448 4713 -432
rect 4937 -56 4971 -40
rect 4937 -448 4971 -432
rect 3469 -525 3485 -491
rect 3585 -525 3601 -491
rect 3727 -525 3743 -491
rect 3843 -525 3859 -491
rect 3985 -525 4001 -491
rect 4101 -525 4117 -491
rect 4243 -525 4259 -491
rect 4359 -525 4375 -491
rect 4501 -525 4517 -491
rect 4617 -525 4633 -491
rect 4759 -525 4775 -491
rect 4875 -525 4891 -491
rect 5365 3 5381 37
rect 5481 3 5497 37
rect 5623 3 5639 37
rect 5739 3 5755 37
rect 5881 3 5897 37
rect 5997 3 6013 37
rect 5285 -56 5319 -40
rect 5285 -448 5319 -432
rect 5543 -56 5577 -40
rect 5543 -448 5577 -432
rect 5801 -56 5835 -40
rect 5801 -448 5835 -432
rect 6059 -56 6093 -40
rect 6059 -448 6093 -432
rect 5365 -525 5381 -491
rect 5481 -525 5497 -491
rect 5623 -525 5639 -491
rect 5739 -525 5755 -491
rect 5881 -525 5897 -491
rect 5997 -525 6013 -491
rect 2828 -565 2978 -549
rect 2828 -660 2874 -565
rect 3275 -593 3309 -531
rect 5051 -593 5085 -531
rect 2862 -669 2874 -660
rect 2828 -703 2840 -694
rect 2828 -763 2874 -703
rect 2908 -648 2978 -599
rect 3275 -627 3371 -593
rect 4989 -627 5085 -593
rect 5171 -593 5205 -531
rect 6173 -593 6207 -531
rect 5171 -627 5267 -593
rect 6111 -627 6207 -593
rect 2908 -675 2934 -648
rect 2908 -709 2930 -675
rect 2964 -709 2978 -696
rect 2908 -729 2978 -709
rect 2828 -797 2978 -763
rect 2035 -907 2101 -865
rect 2621 -869 2637 -835
rect 2671 -869 2687 -835
rect 2927 -805 2978 -797
rect 2759 -855 2793 -839
rect 2621 -907 2687 -869
rect 2827 -865 2843 -831
rect 2877 -865 2893 -831
rect 2961 -839 2978 -805
rect 2927 -855 2978 -839
rect 3275 -791 3371 -757
rect 4989 -791 5085 -757
rect 3275 -852 3309 -791
rect 3275 -853 3276 -852
rect 2827 -907 2893 -865
rect -2064 -941 -2035 -907
rect -2001 -941 -1943 -907
rect -1909 -941 -1851 -907
rect -1817 -941 -1759 -907
rect -1725 -941 -1667 -907
rect -1633 -941 -1575 -907
rect -1541 -941 -1483 -907
rect -1449 -941 -1391 -907
rect -1357 -941 -1299 -907
rect -1265 -941 -1207 -907
rect -1173 -941 -1115 -907
rect -1081 -941 -1023 -907
rect -989 -941 -931 -907
rect -897 -941 -839 -907
rect -805 -941 -747 -907
rect -713 -941 -655 -907
rect -621 -941 -563 -907
rect -529 -941 -471 -907
rect -437 -941 -379 -907
rect -345 -941 -287 -907
rect -253 -941 -195 -907
rect -161 -941 -103 -907
rect -69 -941 -11 -907
rect 23 -941 81 -907
rect 115 -941 173 -907
rect 207 -941 265 -907
rect 299 -941 357 -907
rect 391 -941 449 -907
rect 483 -941 541 -907
rect 575 -941 633 -907
rect 667 -941 725 -907
rect 759 -941 817 -907
rect 851 -941 909 -907
rect 943 -941 1001 -907
rect 1035 -941 1093 -907
rect 1127 -941 1185 -907
rect 1219 -941 1277 -907
rect 1311 -941 1369 -907
rect 1403 -941 1461 -907
rect 1495 -941 1553 -907
rect 1587 -941 1645 -907
rect 1679 -941 1737 -907
rect 1771 -941 1829 -907
rect 1863 -941 1921 -907
rect 1955 -941 2013 -907
rect 2047 -941 2105 -907
rect 2139 -941 2197 -907
rect 2231 -941 2289 -907
rect 2323 -941 2381 -907
rect 2415 -941 2473 -907
rect 2507 -941 2565 -907
rect 2599 -941 2657 -907
rect 2691 -941 2749 -907
rect 2783 -941 2841 -907
rect 2875 -941 2933 -907
rect 2967 -941 2996 -907
rect 5051 -853 5085 -791
rect 5171 -791 5267 -757
rect 6111 -791 6207 -757
rect 5171 -853 5205 -791
rect 6173 -852 6207 -791
rect 6173 -853 6174 -852
rect 3469 -893 3485 -859
rect 3585 -893 3601 -859
rect 3727 -893 3743 -859
rect 3843 -893 3859 -859
rect 3985 -893 4001 -859
rect 4101 -893 4117 -859
rect 4243 -893 4259 -859
rect 4359 -893 4375 -859
rect 4501 -893 4517 -859
rect 4617 -893 4633 -859
rect 4759 -893 4775 -859
rect 4875 -893 4891 -859
rect 3389 -943 3423 -927
rect 3389 -1135 3423 -1119
rect 3647 -943 3681 -927
rect 3647 -1135 3681 -1119
rect 3905 -943 3939 -927
rect 3905 -1135 3939 -1119
rect 4163 -943 4197 -927
rect 4163 -1135 4197 -1119
rect 4421 -943 4455 -927
rect 4421 -1135 4455 -1119
rect 4679 -943 4713 -927
rect 4679 -1135 4713 -1119
rect 4937 -943 4971 -927
rect 4937 -1135 4971 -1119
rect 3469 -1203 3485 -1169
rect 3585 -1203 3601 -1169
rect 3727 -1203 3743 -1169
rect 3843 -1203 3859 -1169
rect 3985 -1203 4001 -1169
rect 4101 -1203 4117 -1169
rect 4243 -1203 4259 -1169
rect 4359 -1203 4375 -1169
rect 4501 -1203 4517 -1169
rect 4617 -1203 4633 -1169
rect 4759 -1203 4775 -1169
rect 4875 -1203 4891 -1169
rect 5365 -893 5381 -859
rect 5481 -893 5497 -859
rect 5623 -893 5639 -859
rect 5739 -893 5755 -859
rect 5881 -893 5897 -859
rect 5997 -893 6013 -859
rect 5285 -943 5319 -927
rect 5285 -1135 5319 -1119
rect 5543 -943 5577 -927
rect 5543 -1135 5577 -1119
rect 5801 -943 5835 -927
rect 5801 -1135 5835 -1119
rect 6059 -943 6093 -927
rect 6059 -1135 6093 -1119
rect 5365 -1203 5381 -1169
rect 5481 -1203 5497 -1169
rect 5623 -1203 5639 -1169
rect 5739 -1203 5755 -1169
rect 5881 -1203 5897 -1169
rect 5997 -1203 6013 -1169
rect 3275 -1271 3309 -1209
rect 5051 -1271 5085 -1209
rect 3275 -1305 3371 -1271
rect 4989 -1305 5085 -1271
rect 5171 -1271 5205 -1209
rect 6173 -1271 6207 -1209
rect 5171 -1305 5267 -1271
rect 6111 -1305 6207 -1271
rect -2522 -1680 -2422 -1518
rect 6822 -1680 6922 -1518
rect -1550 -1946 -1534 -1912
rect -1074 -1946 -1058 -1912
rect -692 -1946 -676 -1912
rect -216 -1946 -200 -1912
rect 166 -1946 182 -1912
rect 642 -1946 658 -1912
rect 1024 -1946 1040 -1912
rect 1500 -1946 1516 -1912
rect 1882 -1946 1898 -1912
rect 2358 -1946 2374 -1912
rect 2740 -1946 2756 -1912
rect 3216 -1946 3232 -1912
rect 3598 -1946 3614 -1912
rect 4074 -1946 4090 -1912
rect 4456 -1946 4472 -1912
rect 4932 -1946 4948 -1912
rect 5314 -1946 5330 -1912
rect 5790 -1946 5806 -1912
rect -1750 -1996 -1716 -1980
rect -1750 -2188 -1716 -2172
rect -892 -1996 -858 -1980
rect -892 -2188 -858 -2172
rect -34 -1996 0 -1980
rect -34 -2188 0 -2172
rect 824 -1996 858 -1980
rect 824 -2188 858 -2172
rect 1682 -1996 1716 -1980
rect 1682 -2188 1716 -2172
rect 2540 -1996 2574 -1980
rect 2540 -2188 2574 -2172
rect 3398 -1996 3432 -1980
rect 3398 -2188 3432 -2172
rect 4256 -1996 4290 -1980
rect 4256 -2188 4290 -2172
rect 5114 -1996 5148 -1980
rect 5114 -2188 5148 -2172
rect 5972 -1996 6006 -1980
rect 5972 -2188 6006 -2172
rect -1550 -2256 -1534 -2222
rect -1074 -2256 -1058 -2222
rect -692 -2256 -676 -2222
rect -216 -2256 -200 -2222
rect 166 -2256 182 -2222
rect 642 -2256 658 -2222
rect 1024 -2256 1040 -2222
rect 1500 -2256 1516 -2222
rect 1882 -2256 1898 -2222
rect 2358 -2256 2374 -2222
rect 2740 -2256 2756 -2222
rect 3216 -2256 3232 -2222
rect 3598 -2256 3614 -2222
rect 4074 -2256 4090 -2222
rect 4456 -2256 4472 -2222
rect 4932 -2256 4948 -2222
rect 5314 -2256 5330 -2222
rect 5790 -2256 5806 -2222
rect -1550 -2528 -1534 -2494
rect -1074 -2528 -1058 -2494
rect -692 -2528 -676 -2494
rect -216 -2528 -200 -2494
rect 166 -2528 182 -2494
rect 642 -2528 658 -2494
rect 1024 -2528 1040 -2494
rect 1500 -2528 1516 -2494
rect 1882 -2528 1898 -2494
rect 2358 -2528 2374 -2494
rect 2740 -2528 2756 -2494
rect 3216 -2528 3232 -2494
rect 3598 -2528 3614 -2494
rect 4074 -2528 4090 -2494
rect 4456 -2528 4472 -2494
rect 4932 -2528 4948 -2494
rect 5314 -2528 5330 -2494
rect 5790 -2528 5806 -2494
rect -1750 -2578 -1716 -2562
rect -1750 -2770 -1716 -2754
rect -892 -2578 -858 -2562
rect -892 -2770 -858 -2754
rect -34 -2578 0 -2562
rect -34 -2770 0 -2754
rect 824 -2578 858 -2562
rect 824 -2770 858 -2754
rect 1682 -2578 1716 -2562
rect 1682 -2770 1716 -2754
rect 2540 -2578 2574 -2562
rect 2540 -2770 2574 -2754
rect 3398 -2578 3432 -2562
rect 3398 -2770 3432 -2754
rect 4256 -2578 4290 -2562
rect 4256 -2770 4290 -2754
rect 5114 -2578 5148 -2562
rect 5114 -2770 5148 -2754
rect 5972 -2578 6006 -2562
rect 5972 -2770 6006 -2754
rect -1550 -2838 -1534 -2804
rect -1074 -2838 -1058 -2804
rect -692 -2838 -676 -2804
rect -216 -2838 -200 -2804
rect 166 -2838 182 -2804
rect 642 -2838 658 -2804
rect 1024 -2838 1040 -2804
rect 1500 -2838 1516 -2804
rect 1882 -2838 1898 -2804
rect 2358 -2838 2374 -2804
rect 2740 -2838 2756 -2804
rect 3216 -2838 3232 -2804
rect 3598 -2838 3614 -2804
rect 4074 -2838 4090 -2804
rect 4456 -2838 4472 -2804
rect 4932 -2838 4948 -2804
rect 5314 -2838 5330 -2804
rect 5790 -2838 5806 -2804
rect -2522 -3782 -2422 -3620
rect 6822 -3782 6922 -3620
<< viali >>
rect -2422 2562 -2360 2662
rect -2360 2562 6760 2662
rect 6760 2562 6822 2662
rect -2522 563 -2422 2457
rect -1880 1643 -1496 1677
rect -1022 1643 -638 1677
rect -164 1643 220 1677
rect 694 1643 1078 1677
rect 1552 1643 1936 1677
rect 2410 1643 2794 1677
rect 3268 1643 3652 1677
rect 4126 1643 4510 1677
rect 4984 1643 5368 1677
rect 5842 1643 6226 1677
rect -2134 1408 -2100 1584
rect -1276 1408 -1242 1584
rect -418 1408 -384 1584
rect 440 1408 474 1584
rect 1298 1408 1332 1584
rect 2156 1408 2190 1584
rect 3014 1408 3048 1584
rect 3872 1408 3906 1584
rect 4730 1408 4764 1584
rect 5588 1408 5622 1584
rect 6446 1408 6480 1584
rect -1880 1315 -1496 1349
rect -1022 1315 -638 1349
rect -164 1315 220 1349
rect 694 1315 1078 1349
rect 1552 1315 1936 1349
rect 2410 1315 2794 1349
rect 3268 1315 3652 1349
rect 4126 1315 4510 1349
rect 4984 1315 5368 1349
rect 5842 1315 6226 1349
rect -1880 1043 -1496 1077
rect -1022 1043 -638 1077
rect -164 1043 220 1077
rect 694 1043 1078 1077
rect 1552 1043 1936 1077
rect 2410 1043 2794 1077
rect 3268 1043 3652 1077
rect 4126 1043 4510 1077
rect 4984 1043 5368 1077
rect 5842 1043 6226 1077
rect -2134 808 -2100 984
rect -1276 808 -1242 984
rect -418 808 -384 984
rect 440 808 474 984
rect 1298 808 1332 984
rect 2156 808 2190 984
rect 3014 808 3048 984
rect 3872 808 3906 984
rect 4730 808 4764 984
rect 5588 808 5622 984
rect 6446 808 6480 984
rect -1880 715 -1496 749
rect -1022 715 -638 749
rect -164 715 220 749
rect 694 715 1078 749
rect 1552 715 1936 749
rect 2410 715 2794 749
rect 3268 715 3652 749
rect 4126 715 4510 749
rect 4984 715 5368 749
rect 5842 715 6226 749
rect 6822 563 6922 2457
rect -2422 358 -2360 458
rect -2360 358 6760 458
rect 6760 358 6822 458
rect 3274 43 3308 46
rect -2035 -397 -2001 -363
rect -1943 -397 -1909 -363
rect -1851 -397 -1817 -363
rect -1759 -397 -1725 -363
rect -1667 -397 -1633 -363
rect -1575 -397 -1541 -363
rect -1483 -397 -1449 -363
rect -1391 -397 -1357 -363
rect -1299 -397 -1265 -363
rect -1207 -397 -1173 -363
rect -1115 -397 -1081 -363
rect -1023 -397 -989 -363
rect -931 -397 -897 -363
rect -839 -397 -805 -363
rect -747 -397 -713 -363
rect -655 -397 -621 -363
rect -563 -397 -529 -363
rect -471 -397 -437 -363
rect -379 -397 -345 -363
rect -287 -397 -253 -363
rect -195 -397 -161 -363
rect -103 -397 -69 -363
rect -11 -397 23 -363
rect 81 -397 115 -363
rect 173 -397 207 -363
rect 265 -397 299 -363
rect 357 -397 391 -363
rect 449 -397 483 -363
rect 541 -397 575 -363
rect 633 -397 667 -363
rect 725 -397 759 -363
rect 817 -397 851 -363
rect 909 -397 943 -363
rect 1001 -397 1035 -363
rect 1093 -397 1127 -363
rect 1185 -397 1219 -363
rect 1277 -397 1311 -363
rect 1369 -397 1403 -363
rect 1461 -397 1495 -363
rect 1553 -397 1587 -363
rect 1645 -397 1679 -363
rect 1737 -397 1771 -363
rect 1829 -397 1863 -363
rect 1921 -397 1955 -363
rect 2013 -397 2047 -363
rect 2105 -397 2139 -363
rect 2197 -397 2231 -363
rect 2289 -397 2323 -363
rect 2381 -397 2415 -363
rect 2473 -397 2507 -363
rect 2565 -397 2599 -363
rect 2657 -397 2691 -363
rect 2749 -397 2783 -363
rect 2841 -397 2875 -363
rect 2933 -397 2967 -363
rect -2044 -675 -1996 -666
rect -2044 -709 -2032 -675
rect -2032 -709 -1998 -675
rect -1998 -709 -1996 -675
rect -2044 -714 -1996 -709
rect -1942 -694 -1930 -669
rect -1930 -694 -1908 -669
rect -1942 -703 -1908 -694
rect -1861 -549 -1827 -533
rect -1861 -567 -1827 -549
rect -1782 -482 -1736 -442
rect -1483 -567 -1449 -533
rect -1575 -703 -1541 -669
rect -859 -559 -825 -533
rect -859 -567 -828 -559
rect -828 -567 -825 -559
rect -1303 -771 -1269 -737
rect -1231 -755 -1207 -737
rect -1207 -755 -1197 -737
rect -1231 -771 -1197 -755
rect -859 -685 -825 -669
rect -859 -703 -833 -685
rect -833 -703 -825 -685
rect -643 -683 -609 -674
rect -643 -708 -627 -683
rect -627 -708 -609 -683
rect -583 -771 -549 -737
rect -320 -716 -272 -668
rect 208 -473 212 -470
rect 212 -473 246 -470
rect 246 -473 256 -470
rect 208 -507 256 -473
rect 208 -518 212 -507
rect 212 -518 246 -507
rect 246 -518 256 -507
rect 444 -575 492 -570
rect 444 -609 447 -575
rect 447 -609 481 -575
rect 481 -609 492 -575
rect 444 -612 492 -609
rect 118 -675 166 -668
rect 118 -708 132 -675
rect 132 -708 166 -675
rect 352 -675 400 -668
rect 352 -709 366 -675
rect 366 -709 400 -675
rect 352 -710 400 -709
rect 526 -675 574 -668
rect 526 -709 534 -675
rect 534 -709 568 -675
rect 568 -709 574 -675
rect 526 -710 574 -709
rect 764 -675 812 -668
rect 764 -708 766 -675
rect 766 -708 800 -675
rect 800 -708 812 -675
rect 676 -793 686 -780
rect 686 -793 720 -780
rect 720 -793 724 -780
rect 676 -827 724 -793
rect 676 -828 686 -827
rect 686 -828 720 -827
rect 720 -828 724 -827
rect 1757 -559 1791 -533
rect 1757 -567 1760 -559
rect 1760 -567 1791 -559
rect 1204 -716 1252 -668
rect 1541 -683 1575 -674
rect 1541 -708 1559 -683
rect 1559 -708 1575 -683
rect 1481 -771 1515 -737
rect 1757 -685 1791 -669
rect 1757 -703 1765 -685
rect 1765 -703 1791 -685
rect 2674 -490 2714 -450
rect 2381 -567 2415 -533
rect 2129 -755 2139 -737
rect 2139 -755 2163 -737
rect 2129 -771 2163 -755
rect 2201 -771 2235 -737
rect 2473 -703 2507 -669
rect 2759 -549 2793 -533
rect 2759 -567 2793 -549
rect 3274 -530 3275 43
rect 3275 -530 3308 43
rect 5050 43 5086 44
rect 3493 3 3577 37
rect 3751 3 3835 37
rect 4009 3 4093 37
rect 4267 3 4351 37
rect 4525 3 4609 37
rect 4783 3 4867 37
rect 3389 -432 3423 -56
rect 3647 -432 3681 -56
rect 3905 -432 3939 -56
rect 4163 -432 4197 -56
rect 4421 -432 4455 -56
rect 4679 -432 4713 -56
rect 4937 -432 4971 -56
rect 3493 -525 3577 -491
rect 3751 -525 3835 -491
rect 4009 -525 4093 -491
rect 4267 -525 4351 -491
rect 4525 -525 4609 -491
rect 4783 -525 4867 -491
rect 5050 -530 5051 43
rect 5051 -530 5085 43
rect 5085 -530 5086 43
rect 5170 43 5206 44
rect 5170 -530 5171 43
rect 5171 -530 5205 43
rect 5205 -530 5206 43
rect 6172 43 6208 44
rect 5389 3 5473 37
rect 5647 3 5731 37
rect 5905 3 5989 37
rect 5285 -432 5319 -56
rect 5543 -432 5577 -56
rect 5801 -432 5835 -56
rect 6059 -432 6093 -56
rect 5389 -525 5473 -491
rect 5647 -525 5731 -491
rect 5905 -525 5989 -491
rect 6172 -530 6173 43
rect 6173 -530 6207 43
rect 6207 -530 6208 43
rect 2840 -694 2862 -669
rect 2862 -694 2874 -669
rect 2840 -703 2874 -694
rect 2934 -675 2982 -648
rect 2934 -696 2964 -675
rect 2964 -696 2982 -675
rect 3276 -853 3310 -852
rect -2035 -941 -2001 -907
rect -1943 -941 -1909 -907
rect -1851 -941 -1817 -907
rect -1759 -941 -1725 -907
rect -1667 -941 -1633 -907
rect -1575 -941 -1541 -907
rect -1483 -941 -1449 -907
rect -1391 -941 -1357 -907
rect -1299 -941 -1265 -907
rect -1207 -941 -1173 -907
rect -1115 -941 -1081 -907
rect -1023 -941 -989 -907
rect -931 -941 -897 -907
rect -839 -941 -805 -907
rect -747 -941 -713 -907
rect -655 -941 -621 -907
rect -563 -941 -529 -907
rect -471 -941 -437 -907
rect -379 -941 -345 -907
rect -287 -941 -253 -907
rect -195 -941 -161 -907
rect -103 -941 -69 -907
rect -11 -941 23 -907
rect 81 -941 115 -907
rect 173 -941 207 -907
rect 265 -941 299 -907
rect 357 -941 391 -907
rect 449 -941 483 -907
rect 541 -941 575 -907
rect 633 -941 667 -907
rect 725 -941 759 -907
rect 817 -941 851 -907
rect 909 -941 943 -907
rect 1001 -941 1035 -907
rect 1093 -941 1127 -907
rect 1185 -941 1219 -907
rect 1277 -941 1311 -907
rect 1369 -941 1403 -907
rect 1461 -941 1495 -907
rect 1553 -941 1587 -907
rect 1645 -941 1679 -907
rect 1737 -941 1771 -907
rect 1829 -941 1863 -907
rect 1921 -941 1955 -907
rect 2013 -941 2047 -907
rect 2105 -941 2139 -907
rect 2197 -941 2231 -907
rect 2289 -941 2323 -907
rect 2381 -941 2415 -907
rect 2473 -941 2507 -907
rect 2565 -941 2599 -907
rect 2657 -941 2691 -907
rect 2749 -941 2783 -907
rect 2841 -941 2875 -907
rect 2933 -941 2967 -907
rect 3276 -1208 3309 -853
rect 3309 -1208 3310 -853
rect 6174 -853 6208 -852
rect 3493 -893 3577 -859
rect 3751 -893 3835 -859
rect 4009 -893 4093 -859
rect 4267 -893 4351 -859
rect 4525 -893 4609 -859
rect 4783 -893 4867 -859
rect 3389 -1119 3423 -943
rect 3647 -1119 3681 -943
rect 3905 -1119 3939 -943
rect 4163 -1119 4197 -943
rect 4421 -1119 4455 -943
rect 4679 -1119 4713 -943
rect 4937 -1119 4971 -943
rect 3493 -1203 3577 -1169
rect 3751 -1203 3835 -1169
rect 4009 -1203 4093 -1169
rect 4267 -1203 4351 -1169
rect 4525 -1203 4609 -1169
rect 4783 -1203 4867 -1169
rect 5052 -1208 5085 -854
rect 5085 -1208 5086 -854
rect 5172 -1208 5205 -854
rect 5205 -1208 5206 -854
rect 5389 -893 5473 -859
rect 5647 -893 5731 -859
rect 5905 -893 5989 -859
rect 5285 -1119 5319 -943
rect 5543 -1119 5577 -943
rect 5801 -1119 5835 -943
rect 6059 -1119 6093 -943
rect 5389 -1203 5473 -1169
rect 5647 -1203 5731 -1169
rect 5905 -1203 5989 -1169
rect 6174 -1208 6207 -853
rect 6207 -1208 6208 -853
rect -2422 -1618 -2360 -1518
rect -2360 -1618 6760 -1518
rect 6760 -1618 6822 -1518
rect -2522 -3584 -2422 -1716
rect -1496 -1946 -1112 -1912
rect -638 -1946 -254 -1912
rect 220 -1946 604 -1912
rect 1078 -1946 1462 -1912
rect 1936 -1946 2320 -1912
rect 2794 -1946 3178 -1912
rect 3652 -1946 4036 -1912
rect 4510 -1946 4894 -1912
rect 5368 -1946 5752 -1912
rect -1750 -2172 -1716 -1996
rect -892 -2172 -858 -1996
rect -34 -2172 0 -1996
rect 824 -2172 858 -1996
rect 1682 -2172 1716 -1996
rect 2540 -2172 2574 -1996
rect 3398 -2172 3432 -1996
rect 4256 -2172 4290 -1996
rect 5114 -2172 5148 -1996
rect 5972 -2172 6006 -1996
rect -1496 -2256 -1112 -2222
rect -638 -2256 -254 -2222
rect 220 -2256 604 -2222
rect 1078 -2256 1462 -2222
rect 1936 -2256 2320 -2222
rect 2794 -2256 3178 -2222
rect 3652 -2256 4036 -2222
rect 4510 -2256 4894 -2222
rect 5368 -2256 5752 -2222
rect -1496 -2528 -1112 -2494
rect -638 -2528 -254 -2494
rect 220 -2528 604 -2494
rect 1078 -2528 1462 -2494
rect 1936 -2528 2320 -2494
rect 2794 -2528 3178 -2494
rect 3652 -2528 4036 -2494
rect 4510 -2528 4894 -2494
rect 5368 -2528 5752 -2494
rect -1750 -2754 -1716 -2578
rect -892 -2754 -858 -2578
rect -34 -2754 0 -2578
rect 824 -2754 858 -2578
rect 1682 -2754 1716 -2578
rect 2540 -2754 2574 -2578
rect 3398 -2754 3432 -2578
rect 4256 -2754 4290 -2578
rect 5114 -2754 5148 -2578
rect 5972 -2754 6006 -2578
rect -1496 -2838 -1112 -2804
rect -638 -2838 -254 -2804
rect 220 -2838 604 -2804
rect 1078 -2838 1462 -2804
rect 1936 -2838 2320 -2804
rect 2794 -2838 3178 -2804
rect 3652 -2838 4036 -2804
rect 4510 -2838 4894 -2804
rect 5368 -2838 5752 -2804
rect 6822 -3584 6922 -1716
rect -2422 -3782 -2360 -3682
rect -2360 -3782 6760 -3682
rect 6760 -3782 6822 -3682
<< metal1 >>
rect -2528 2662 6928 2668
rect -2528 2562 -2422 2662
rect 6822 2562 6928 2662
rect -2528 2556 6928 2562
rect -2528 2457 -2416 2556
rect -2528 563 -2522 2457
rect -2422 563 -2416 2457
rect -1816 2256 -1806 2556
rect 6206 2256 6216 2556
rect 6816 2457 6928 2556
rect -2340 2140 6730 2174
rect -2340 2030 -2302 2140
rect 6694 2030 6730 2140
rect -2340 1992 6730 2030
rect -2304 1774 -2298 1834
rect -2238 1774 -2232 1834
rect -2146 1806 -2086 1992
rect -1724 1806 -1664 1992
rect -2298 636 -2238 1774
rect -2146 1746 -1664 1806
rect -1296 1774 -1290 1834
rect -1230 1774 -1224 1834
rect -432 1828 -372 1992
rect 1286 1828 1346 1992
rect 3002 1832 3062 1992
rect 4716 1832 4776 1992
rect -2146 1584 -2086 1746
rect -1724 1683 -1664 1746
rect -1892 1677 -1484 1683
rect -1892 1643 -1880 1677
rect -1496 1643 -1484 1677
rect -1892 1637 -1484 1643
rect -2146 1408 -2134 1584
rect -2100 1408 -2086 1584
rect -1290 1584 -1230 1774
rect -432 1768 1346 1828
rect 2134 1768 2140 1828
rect 2200 1768 2206 1828
rect 3002 1772 4776 1832
rect -1034 1677 -626 1683
rect -1034 1643 -1022 1677
rect -638 1643 -626 1677
rect -1034 1637 -626 1643
rect -1290 1536 -1276 1584
rect -2146 1228 -2086 1408
rect -1282 1408 -1276 1536
rect -1242 1536 -1230 1584
rect -432 1584 -372 1768
rect -176 1677 232 1683
rect -176 1643 -164 1677
rect 220 1643 232 1677
rect -176 1637 232 1643
rect 682 1677 1090 1683
rect 682 1643 694 1677
rect 1078 1643 1090 1677
rect 682 1637 1090 1643
rect -1242 1408 -1236 1536
rect -1282 1396 -1236 1408
rect -432 1408 -418 1584
rect -384 1408 -372 1584
rect 434 1584 480 1596
rect 434 1470 440 1584
rect -1892 1349 -1484 1355
rect -1892 1315 -1880 1349
rect -1496 1315 -1484 1349
rect -1892 1309 -1484 1315
rect -1034 1349 -626 1355
rect -1034 1315 -1022 1349
rect -638 1315 -626 1349
rect -1034 1309 -626 1315
rect -1722 1228 -1662 1309
rect -856 1228 -796 1309
rect -2146 1168 -1662 1228
rect -1296 1168 -1290 1228
rect -1230 1168 -1224 1228
rect -862 1168 -856 1228
rect -796 1168 -790 1228
rect -2146 984 -2086 1168
rect -1722 1083 -1662 1168
rect -1892 1077 -1484 1083
rect -1892 1043 -1880 1077
rect -1496 1043 -1484 1077
rect -1892 1037 -1484 1043
rect -2146 808 -2134 984
rect -2100 808 -2086 984
rect -1290 984 -1230 1168
rect -856 1083 -796 1168
rect -1034 1077 -626 1083
rect -1034 1043 -1022 1077
rect -638 1043 -626 1077
rect -1034 1037 -626 1043
rect -1290 942 -1276 984
rect -2146 648 -2086 808
rect -1282 808 -1276 942
rect -1242 942 -1230 984
rect -432 984 -372 1408
rect 426 1408 440 1470
rect 474 1470 480 1584
rect 1286 1584 1346 1768
rect 1540 1677 1948 1683
rect 1540 1643 1552 1677
rect 1936 1643 1948 1677
rect 1540 1637 1948 1643
rect 474 1408 486 1470
rect -176 1349 232 1355
rect -176 1315 -164 1349
rect 220 1315 232 1349
rect -176 1309 232 1315
rect -6 1228 54 1309
rect 426 1228 486 1408
rect 1286 1408 1298 1584
rect 1332 1408 1346 1584
rect 2140 1584 2200 1768
rect 2398 1677 2806 1683
rect 2398 1643 2410 1677
rect 2794 1643 2806 1677
rect 2398 1637 2806 1643
rect 2140 1530 2156 1584
rect 682 1349 1090 1355
rect 682 1315 694 1349
rect 1078 1315 1090 1349
rect 682 1309 1090 1315
rect 856 1228 916 1309
rect -12 1168 -6 1228
rect 54 1168 60 1228
rect 420 1168 426 1228
rect 486 1168 492 1228
rect 850 1168 856 1228
rect 916 1168 922 1228
rect -6 1083 54 1168
rect 856 1083 916 1168
rect -176 1077 232 1083
rect -176 1043 -164 1077
rect 220 1043 232 1077
rect -176 1037 232 1043
rect 682 1077 1090 1083
rect 682 1043 694 1077
rect 1078 1043 1090 1077
rect 682 1037 1090 1043
rect -432 946 -418 984
rect -1242 808 -1236 942
rect -1282 796 -1236 808
rect -424 808 -418 946
rect -384 946 -372 984
rect 434 984 480 996
rect -384 808 -378 946
rect 434 854 440 984
rect -424 796 -378 808
rect 426 808 440 854
rect 474 854 480 984
rect 1286 984 1346 1408
rect 2150 1408 2156 1530
rect 2190 1530 2200 1584
rect 3002 1584 3062 1772
rect 3256 1677 3664 1683
rect 3256 1643 3268 1677
rect 3652 1643 3664 1677
rect 3256 1637 3664 1643
rect 4114 1677 4522 1683
rect 4114 1643 4126 1677
rect 4510 1643 4522 1677
rect 4114 1637 4522 1643
rect 2190 1408 2196 1530
rect 2150 1396 2196 1408
rect 3002 1408 3014 1584
rect 3048 1408 3062 1584
rect 3866 1584 3912 1596
rect 3866 1470 3872 1584
rect 1540 1349 1948 1355
rect 1540 1315 1552 1349
rect 1936 1315 1948 1349
rect 1540 1309 1948 1315
rect 2398 1349 2806 1355
rect 2398 1315 2410 1349
rect 2794 1315 2806 1349
rect 2398 1309 2806 1315
rect 1712 1228 1772 1309
rect 2564 1228 2624 1309
rect 1706 1168 1712 1228
rect 1772 1168 1778 1228
rect 2138 1168 2144 1228
rect 2204 1168 2210 1228
rect 2558 1168 2564 1228
rect 2624 1168 2630 1228
rect 1712 1083 1772 1168
rect 1540 1077 1948 1083
rect 1540 1043 1552 1077
rect 1936 1043 1948 1077
rect 1540 1037 1948 1043
rect 1286 930 1298 984
rect 474 808 486 854
rect -1892 749 -1484 755
rect -1892 715 -1880 749
rect -1496 715 -1484 749
rect -1892 709 -1484 715
rect -1034 749 -626 755
rect -1034 715 -1022 749
rect -638 715 -626 749
rect -1034 709 -626 715
rect -176 749 232 755
rect -176 715 -164 749
rect 220 715 232 749
rect -176 709 232 715
rect -1726 648 -1666 709
rect -2304 576 -2298 636
rect -2238 576 -2232 636
rect -2146 588 -1666 648
rect 426 636 486 808
rect 1292 808 1298 930
rect 1332 930 1346 984
rect 2144 984 2204 1168
rect 2564 1083 2624 1168
rect 2398 1077 2806 1083
rect 2398 1043 2410 1077
rect 2794 1043 2806 1077
rect 2398 1037 2806 1043
rect 2144 938 2156 984
rect 1332 808 1338 930
rect 1292 796 1338 808
rect 2150 808 2156 938
rect 2190 938 2204 984
rect 3002 984 3062 1408
rect 3860 1408 3872 1470
rect 3906 1470 3912 1584
rect 4716 1584 4776 1772
rect 5568 1768 5574 1828
rect 5634 1768 5640 1828
rect 6000 1820 6060 1992
rect 6432 1820 6492 1992
rect 4972 1677 5380 1683
rect 4972 1643 4984 1677
rect 5368 1643 5380 1677
rect 4972 1637 5380 1643
rect 3906 1408 3920 1470
rect 3256 1349 3664 1355
rect 3256 1315 3268 1349
rect 3652 1315 3664 1349
rect 3256 1309 3664 1315
rect 3426 1228 3486 1309
rect 3860 1228 3920 1408
rect 4716 1408 4730 1584
rect 4764 1408 4776 1584
rect 5574 1584 5634 1768
rect 6000 1760 6492 1820
rect 6588 1768 6594 1828
rect 6654 1768 6660 1828
rect 6000 1683 6060 1760
rect 5830 1677 6238 1683
rect 5830 1643 5842 1677
rect 6226 1643 6238 1677
rect 5830 1637 6238 1643
rect 5574 1554 5588 1584
rect 4114 1349 4522 1355
rect 4114 1315 4126 1349
rect 4510 1315 4522 1349
rect 4114 1309 4522 1315
rect 4296 1228 4356 1309
rect 3420 1168 3426 1228
rect 3486 1168 3492 1228
rect 3854 1168 3860 1228
rect 3920 1168 3926 1228
rect 4290 1168 4296 1228
rect 4356 1168 4362 1228
rect 3426 1083 3486 1168
rect 4296 1083 4356 1168
rect 3256 1077 3664 1083
rect 3256 1043 3268 1077
rect 3652 1043 3664 1077
rect 3256 1037 3664 1043
rect 4114 1077 4522 1083
rect 4114 1043 4126 1077
rect 4510 1043 4522 1077
rect 4114 1037 4522 1043
rect 2190 808 2196 938
rect 3002 934 3014 984
rect 2150 796 2196 808
rect 3008 808 3014 934
rect 3048 934 3062 984
rect 3866 984 3912 996
rect 3048 808 3054 934
rect 3866 858 3872 984
rect 3008 796 3054 808
rect 3856 808 3872 858
rect 3906 858 3912 984
rect 4716 984 4776 1408
rect 5582 1408 5588 1554
rect 5622 1554 5634 1584
rect 6432 1584 6492 1760
rect 5622 1408 5628 1554
rect 5582 1396 5628 1408
rect 6432 1408 6446 1584
rect 6480 1408 6492 1584
rect 4972 1349 5380 1355
rect 4972 1315 4984 1349
rect 5368 1315 5380 1349
rect 4972 1309 5380 1315
rect 5830 1349 6238 1355
rect 5830 1315 5842 1349
rect 6226 1315 6238 1349
rect 5830 1309 6238 1315
rect 5136 1228 5196 1309
rect 5130 1168 5136 1228
rect 5196 1168 5202 1228
rect 5570 1168 5576 1228
rect 5636 1168 5642 1228
rect 6000 1226 6060 1309
rect 6432 1226 6492 1408
rect 5136 1083 5196 1168
rect 4972 1077 5380 1083
rect 4972 1043 4984 1077
rect 5368 1043 5380 1077
rect 4972 1037 5380 1043
rect 4716 940 4730 984
rect 3906 808 3916 858
rect 682 749 1090 755
rect 682 715 694 749
rect 1078 715 1090 749
rect 682 709 1090 715
rect 1540 749 1948 755
rect 1540 715 1552 749
rect 1936 715 1948 749
rect 1540 709 1948 715
rect 2398 749 2806 755
rect 2398 715 2410 749
rect 2794 715 2806 749
rect 2398 709 2806 715
rect 3256 749 3664 755
rect 3256 715 3268 749
rect 3652 715 3664 749
rect 3256 709 3664 715
rect 3856 636 3916 808
rect 4724 808 4730 940
rect 4764 940 4776 984
rect 5576 984 5636 1168
rect 6000 1166 6492 1226
rect 6000 1083 6060 1166
rect 5830 1077 6238 1083
rect 5830 1043 5842 1077
rect 6226 1043 6238 1077
rect 5830 1037 6238 1043
rect 4764 808 4770 940
rect 5576 938 5588 984
rect 4724 796 4770 808
rect 5582 808 5588 938
rect 5622 938 5636 984
rect 6432 984 6492 1166
rect 5622 808 5628 938
rect 5582 796 5628 808
rect 6432 808 6446 984
rect 6480 808 6492 984
rect 4114 749 4522 755
rect 4114 715 4126 749
rect 4510 715 4522 749
rect 4114 709 4522 715
rect 4972 749 5380 755
rect 4972 715 4984 749
rect 5368 715 5380 749
rect 4972 709 5380 715
rect 5830 749 6238 755
rect 5830 715 5842 749
rect 6226 715 6238 749
rect 5830 709 6238 715
rect 5996 644 6056 709
rect 6432 644 6492 808
rect -2528 464 -2416 563
rect -2146 464 -2086 588
rect -1726 464 -1666 588
rect 420 576 426 636
rect 486 576 492 636
rect 3850 576 3856 636
rect 3916 576 3922 636
rect 5996 584 6494 644
rect 6594 636 6654 1768
rect 5996 464 6056 584
rect 6432 464 6492 584
rect 6588 576 6594 636
rect 6654 576 6660 636
rect 6816 563 6822 2457
rect 6922 563 6928 2457
rect 6816 464 6928 563
rect -2528 458 6928 464
rect -2528 358 -2422 458
rect 6822 358 6928 458
rect -2528 352 6928 358
rect -2066 -332 -1822 352
rect -1066 -332 -822 352
rect -66 -332 178 352
rect 934 -332 1178 352
rect 1934 -332 2178 352
rect 2750 -332 2994 352
rect 3260 156 3324 352
rect 3376 156 3436 352
rect 3510 156 3570 352
rect 3634 156 3694 352
rect 3260 96 3694 156
rect 3260 46 3324 96
rect -2066 -363 2996 -332
rect -2066 -397 -2035 -363
rect -2001 -397 -1943 -363
rect -1909 -397 -1851 -363
rect -1817 -397 -1759 -363
rect -1725 -397 -1667 -363
rect -1633 -397 -1575 -363
rect -1541 -397 -1483 -363
rect -1449 -397 -1391 -363
rect -1357 -397 -1299 -363
rect -1265 -397 -1207 -363
rect -1173 -397 -1115 -363
rect -1081 -397 -1023 -363
rect -989 -397 -931 -363
rect -897 -397 -839 -363
rect -805 -397 -747 -363
rect -713 -397 -655 -363
rect -621 -397 -563 -363
rect -529 -397 -471 -363
rect -437 -397 -379 -363
rect -345 -397 -287 -363
rect -253 -397 -195 -363
rect -161 -397 -103 -363
rect -69 -397 -11 -363
rect 23 -397 81 -363
rect 115 -397 173 -363
rect 207 -397 265 -363
rect 299 -397 357 -363
rect 391 -397 449 -363
rect 483 -397 541 -363
rect 575 -397 633 -363
rect 667 -397 725 -363
rect 759 -397 817 -363
rect 851 -397 909 -363
rect 943 -397 1001 -363
rect 1035 -397 1093 -363
rect 1127 -397 1185 -363
rect 1219 -397 1277 -363
rect 1311 -397 1369 -363
rect 1403 -397 1461 -363
rect 1495 -397 1553 -363
rect 1587 -397 1645 -363
rect 1679 -397 1737 -363
rect 1771 -397 1829 -363
rect 1863 -397 1921 -363
rect 1955 -397 2013 -363
rect 2047 -397 2105 -363
rect 2139 -397 2197 -363
rect 2231 -397 2289 -363
rect 2323 -397 2381 -363
rect 2415 -397 2473 -363
rect 2507 -397 2565 -363
rect 2599 -397 2657 -363
rect 2691 -397 2749 -363
rect 2783 -397 2841 -363
rect 2875 -397 2933 -363
rect 2967 -397 2996 -363
rect -2066 -428 2996 -397
rect -1794 -442 -1728 -428
rect -1794 -482 -1782 -442
rect -1736 -482 -1728 -442
rect 2660 -450 2726 -428
rect 202 -464 262 -458
rect -1794 -496 -1728 -482
rect 196 -524 202 -464
rect 262 -524 268 -464
rect 2660 -490 2674 -450
rect 2714 -490 2726 -450
rect 2660 -502 2726 -490
rect -1873 -533 -1815 -527
rect -1873 -567 -1861 -533
rect -1827 -536 -1815 -533
rect -1495 -533 -1437 -527
rect -1495 -536 -1483 -533
rect -1827 -564 -1483 -536
rect -1827 -567 -1815 -564
rect -1873 -573 -1815 -567
rect -1495 -567 -1483 -564
rect -1449 -536 -1437 -533
rect -871 -533 -813 -527
rect 202 -530 262 -524
rect -871 -536 -859 -533
rect -1449 -564 -859 -536
rect -1449 -567 -1437 -564
rect -1495 -573 -1437 -567
rect -871 -567 -859 -564
rect -825 -567 -813 -533
rect 1745 -533 1803 -527
rect -871 -573 -813 -567
rect -660 -570 1586 -564
rect -660 -612 444 -570
rect 492 -612 1586 -570
rect 1745 -567 1757 -533
rect 1791 -536 1803 -533
rect 2369 -533 2427 -527
rect 2369 -536 2381 -533
rect 1791 -564 2381 -536
rect 1791 -567 1803 -564
rect 1745 -573 1803 -567
rect 2369 -567 2381 -564
rect 2415 -536 2427 -533
rect 2747 -533 2805 -527
rect 2747 -536 2759 -533
rect 2415 -564 2759 -536
rect 2415 -567 2427 -564
rect 2369 -573 2427 -567
rect 2747 -567 2759 -564
rect 2793 -567 2805 -533
rect 3260 -530 3274 46
rect 3308 -530 3324 46
rect 3376 -56 3436 96
rect 3510 43 3570 96
rect 3481 37 3589 43
rect 3481 3 3493 37
rect 3577 3 3589 37
rect 3481 -3 3589 3
rect 3376 -72 3389 -56
rect 3383 -432 3389 -72
rect 3423 -72 3436 -56
rect 3634 -56 3694 96
rect 4022 156 4082 352
rect 4152 156 4212 352
rect 4280 156 4340 352
rect 4798 164 4858 352
rect 4928 164 4988 352
rect 4022 96 4340 156
rect 4534 98 4540 158
rect 4600 98 4606 158
rect 4022 43 4082 96
rect 3739 37 3847 43
rect 3739 3 3751 37
rect 3835 3 3847 37
rect 3739 -3 3847 3
rect 3997 37 4105 43
rect 3997 3 4009 37
rect 4093 3 4105 37
rect 3997 -3 4105 3
rect 3423 -432 3429 -72
rect 3634 -94 3647 -56
rect 3383 -444 3429 -432
rect 3641 -432 3647 -94
rect 3681 -94 3694 -56
rect 3899 -56 3945 -44
rect 3681 -432 3687 -94
rect 3899 -384 3905 -56
rect 3641 -444 3687 -432
rect 3892 -432 3905 -384
rect 3939 -384 3945 -56
rect 4152 -56 4212 96
rect 4280 43 4340 96
rect 4540 43 4600 98
rect 4662 96 4668 156
rect 4728 96 4734 156
rect 4798 104 4988 164
rect 4255 37 4363 43
rect 4255 3 4267 37
rect 4351 3 4363 37
rect 4255 -3 4363 3
rect 4513 37 4621 43
rect 4513 3 4525 37
rect 4609 3 4621 37
rect 4513 -3 4621 3
rect 4152 -84 4163 -56
rect 3939 -432 3952 -384
rect 3260 -540 3324 -530
rect 3481 -491 3589 -485
rect 3481 -525 3493 -491
rect 3577 -525 3589 -491
rect 3481 -531 3589 -525
rect 3739 -491 3847 -485
rect 3739 -525 3751 -491
rect 3835 -525 3847 -491
rect 3739 -531 3847 -525
rect 2747 -573 2805 -567
rect 3764 -574 3824 -531
rect 3892 -574 3952 -432
rect 4157 -432 4163 -84
rect 4197 -84 4212 -56
rect 4415 -56 4461 -44
rect 4197 -432 4203 -84
rect 4415 -398 4421 -56
rect 4157 -444 4203 -432
rect 4410 -432 4421 -398
rect 4455 -398 4461 -56
rect 4668 -56 4728 96
rect 4798 43 4858 104
rect 4771 37 4879 43
rect 4771 3 4783 37
rect 4867 3 4879 37
rect 4771 -3 4879 3
rect 4668 -96 4679 -56
rect 4455 -432 4470 -398
rect 3997 -491 4105 -485
rect 3997 -525 4009 -491
rect 4093 -525 4105 -491
rect 3997 -531 4105 -525
rect 4255 -491 4363 -485
rect 4255 -525 4267 -491
rect 4351 -525 4363 -491
rect 4255 -531 4363 -525
rect -660 -624 1586 -612
rect -2292 -666 -1984 -660
rect -2292 -714 -2044 -666
rect -1996 -714 -1984 -666
rect -1954 -669 -1896 -663
rect -1954 -703 -1942 -669
rect -1908 -672 -1896 -669
rect -1587 -669 -1529 -663
rect -1587 -672 -1575 -669
rect -1908 -700 -1575 -672
rect -1908 -703 -1896 -700
rect -1954 -709 -1896 -703
rect -1587 -703 -1575 -700
rect -1541 -672 -1529 -669
rect -871 -669 -813 -663
rect -871 -672 -859 -669
rect -1541 -700 -859 -672
rect -1541 -703 -1529 -700
rect -1587 -709 -1529 -703
rect -871 -703 -859 -700
rect -825 -703 -813 -669
rect -871 -709 -813 -703
rect -660 -668 -600 -624
rect 436 -626 496 -624
rect 348 -662 408 -656
rect 840 -662 900 -656
rect -332 -668 348 -662
rect -660 -674 -597 -668
rect -660 -708 -643 -674
rect -609 -708 -597 -674
rect -2292 -720 -1984 -714
rect -660 -731 -597 -708
rect -332 -716 -320 -668
rect -272 -708 118 -668
rect 166 -708 348 -668
rect -272 -716 348 -708
rect -332 -722 348 -716
rect 408 -722 412 -662
rect 514 -668 840 -662
rect 514 -710 526 -668
rect 574 -708 764 -668
rect 812 -708 840 -668
rect 574 -710 840 -708
rect 514 -722 840 -710
rect 900 -668 1264 -662
rect 900 -716 1204 -668
rect 1252 -716 1264 -668
rect 900 -722 1264 -716
rect 1526 -668 1586 -624
rect 3632 -634 3952 -574
rect 2922 -648 3104 -642
rect 1526 -674 1587 -668
rect 1526 -708 1541 -674
rect 1575 -708 1587 -674
rect 348 -728 408 -722
rect 840 -728 900 -722
rect 1526 -731 1587 -708
rect 1745 -669 1803 -663
rect 1745 -703 1757 -669
rect 1791 -672 1803 -669
rect 2461 -669 2519 -663
rect 2461 -672 2473 -669
rect 1791 -700 2473 -672
rect 1791 -703 1803 -700
rect 1745 -709 1803 -703
rect 2461 -703 2473 -700
rect 2507 -672 2519 -669
rect 2828 -669 2886 -663
rect 2828 -672 2840 -669
rect 2507 -700 2840 -672
rect 2507 -703 2519 -700
rect 2461 -709 2519 -703
rect 2828 -703 2840 -700
rect 2874 -703 2886 -669
rect 2922 -696 2934 -648
rect 2982 -696 3104 -648
rect 2922 -702 3104 -696
rect 2828 -709 2886 -703
rect -1315 -737 -1185 -731
rect -1315 -771 -1303 -737
rect -1269 -771 -1231 -737
rect -1197 -740 -1185 -737
rect -660 -737 -537 -731
rect -660 -740 -583 -737
rect -1197 -768 -583 -740
rect -1197 -771 -1185 -768
rect -1315 -777 -1185 -771
rect -595 -771 -583 -768
rect -549 -771 -537 -737
rect 1469 -737 1587 -731
rect -595 -777 -537 -771
rect 670 -774 730 -768
rect 1469 -771 1481 -737
rect 1515 -740 1587 -737
rect 2117 -737 2247 -731
rect 2117 -740 2129 -737
rect 1515 -768 2129 -740
rect 1515 -771 1527 -768
rect 664 -834 670 -774
rect 730 -834 736 -774
rect 1469 -777 1527 -771
rect 2117 -771 2129 -768
rect 2163 -771 2201 -737
rect 2235 -771 2247 -737
rect 2117 -777 2247 -771
rect 670 -840 730 -834
rect 3262 -852 3326 -840
rect -2064 -907 2996 -876
rect -2064 -941 -2035 -907
rect -2001 -941 -1943 -907
rect -1909 -941 -1851 -907
rect -1817 -941 -1759 -907
rect -1725 -941 -1667 -907
rect -1633 -941 -1575 -907
rect -1541 -941 -1483 -907
rect -1449 -941 -1391 -907
rect -1357 -941 -1299 -907
rect -1265 -941 -1207 -907
rect -1173 -941 -1115 -907
rect -1081 -941 -1023 -907
rect -989 -941 -931 -907
rect -897 -941 -839 -907
rect -805 -941 -747 -907
rect -713 -941 -655 -907
rect -621 -941 -563 -907
rect -529 -941 -471 -907
rect -437 -941 -379 -907
rect -345 -941 -287 -907
rect -253 -941 -195 -907
rect -161 -941 -103 -907
rect -69 -941 -11 -907
rect 23 -941 81 -907
rect 115 -941 173 -907
rect 207 -941 265 -907
rect 299 -941 357 -907
rect 391 -941 449 -907
rect 483 -941 541 -907
rect 575 -941 633 -907
rect 667 -941 725 -907
rect 759 -941 817 -907
rect 851 -941 909 -907
rect 943 -941 1001 -907
rect 1035 -941 1093 -907
rect 1127 -941 1185 -907
rect 1219 -941 1277 -907
rect 1311 -941 1369 -907
rect 1403 -941 1461 -907
rect 1495 -941 1553 -907
rect 1587 -941 1645 -907
rect 1679 -941 1737 -907
rect 1771 -941 1829 -907
rect 1863 -941 1921 -907
rect 1955 -941 2013 -907
rect 2047 -941 2105 -907
rect 2139 -941 2197 -907
rect 2231 -941 2289 -907
rect 2323 -941 2381 -907
rect 2415 -941 2473 -907
rect 2507 -941 2565 -907
rect 2599 -941 2657 -907
rect 2691 -941 2749 -907
rect 2783 -941 2841 -907
rect 2875 -941 2933 -907
rect 2967 -941 2996 -907
rect -2064 -942 2996 -941
rect -2066 -972 2996 -942
rect -2066 -1512 -1822 -972
rect -1066 -1512 -822 -972
rect -66 -1512 178 -972
rect 934 -1512 1178 -972
rect 1934 -1512 2178 -972
rect 2752 -1512 2996 -972
rect 3262 -1208 3276 -852
rect 3310 -1208 3326 -852
rect 3481 -859 3589 -853
rect 3481 -893 3493 -859
rect 3577 -893 3589 -859
rect 3481 -899 3589 -893
rect 3383 -943 3429 -931
rect 3383 -1072 3389 -943
rect 3262 -1258 3326 -1208
rect 3376 -1119 3389 -1072
rect 3423 -1072 3429 -943
rect 3632 -943 3692 -634
rect 4410 -744 4470 -432
rect 4673 -432 4679 -96
rect 4713 -96 4728 -56
rect 4928 -56 4988 104
rect 4713 -432 4719 -96
rect 4928 -107 4937 -56
rect 4673 -444 4719 -432
rect 4931 -432 4937 -107
rect 4971 -107 4988 -56
rect 5034 159 5224 352
rect 5274 159 5334 352
rect 5404 159 5464 352
rect 5656 240 5662 300
rect 5722 240 5728 300
rect 5034 99 5464 159
rect 5034 44 5224 99
rect 4971 -432 4977 -107
rect 4931 -444 4977 -432
rect 4513 -491 4621 -485
rect 4513 -525 4525 -491
rect 4609 -525 4621 -491
rect 4513 -531 4621 -525
rect 4771 -491 4879 -485
rect 4771 -525 4783 -491
rect 4867 -525 4879 -491
rect 4771 -531 4879 -525
rect 5034 -530 5050 44
rect 5086 -530 5170 44
rect 5206 -530 5224 44
rect 5274 -56 5334 99
rect 5404 43 5464 99
rect 5526 96 5532 156
rect 5592 96 5598 156
rect 5377 37 5485 43
rect 5377 3 5389 37
rect 5473 3 5485 37
rect 5377 -3 5485 3
rect 5274 -98 5285 -56
rect 5279 -432 5285 -98
rect 5319 -98 5334 -56
rect 5532 -56 5592 96
rect 5662 43 5722 240
rect 5920 164 5980 352
rect 6044 164 6104 352
rect 6158 164 6222 352
rect 5920 104 6222 164
rect 5920 43 5980 104
rect 5635 37 5743 43
rect 5635 3 5647 37
rect 5731 3 5743 37
rect 5635 -3 5743 3
rect 5893 37 6001 43
rect 5893 3 5905 37
rect 5989 3 6001 37
rect 5893 -3 6001 3
rect 5532 -92 5543 -56
rect 5319 -432 5325 -98
rect 5279 -444 5325 -432
rect 5537 -432 5543 -92
rect 5577 -92 5592 -56
rect 5795 -56 5841 -44
rect 5577 -432 5583 -92
rect 5795 -406 5801 -56
rect 5537 -444 5583 -432
rect 5788 -432 5801 -406
rect 5835 -406 5841 -56
rect 6044 -56 6104 104
rect 6044 -84 6059 -56
rect 5835 -432 5848 -406
rect 5034 -544 5224 -530
rect 5377 -491 5485 -485
rect 5377 -525 5389 -491
rect 5473 -525 5485 -491
rect 5377 -531 5485 -525
rect 5635 -491 5743 -485
rect 5635 -525 5647 -491
rect 5731 -525 5743 -491
rect 5635 -531 5743 -525
rect 4410 -804 4598 -744
rect 3739 -859 3847 -853
rect 3739 -893 3751 -859
rect 3835 -893 3847 -859
rect 3739 -899 3847 -893
rect 3997 -859 4105 -853
rect 3997 -893 4009 -859
rect 4093 -893 4105 -859
rect 3997 -899 4105 -893
rect 4255 -859 4363 -853
rect 4255 -893 4267 -859
rect 4351 -893 4363 -859
rect 4255 -899 4363 -893
rect 3632 -982 3647 -943
rect 3423 -1119 3436 -1072
rect 3376 -1258 3436 -1119
rect 3641 -1119 3647 -982
rect 3681 -982 3692 -943
rect 3899 -943 3945 -931
rect 3681 -1119 3687 -982
rect 3899 -1086 3905 -943
rect 3641 -1131 3687 -1119
rect 3892 -1119 3905 -1086
rect 3939 -1086 3945 -943
rect 4157 -943 4203 -931
rect 4157 -1082 4163 -943
rect 3939 -1119 3952 -1086
rect 3481 -1169 3589 -1163
rect 3481 -1203 3493 -1169
rect 3577 -1203 3589 -1169
rect 3481 -1209 3589 -1203
rect 3739 -1169 3847 -1163
rect 3739 -1203 3751 -1169
rect 3835 -1203 3847 -1169
rect 3739 -1209 3847 -1203
rect 3510 -1258 3570 -1209
rect 3262 -1318 3570 -1258
rect 3262 -1512 3326 -1318
rect 3376 -1512 3436 -1318
rect 3510 -1512 3570 -1318
rect 3754 -1394 3814 -1209
rect 3748 -1454 3754 -1394
rect 3814 -1454 3820 -1394
rect 3892 -1396 3952 -1119
rect 4150 -1119 4163 -1082
rect 4197 -1082 4203 -943
rect 4410 -943 4470 -804
rect 4538 -853 4598 -804
rect 4513 -859 4621 -853
rect 4513 -893 4525 -859
rect 4609 -893 4621 -859
rect 4513 -899 4621 -893
rect 4771 -859 4879 -853
rect 4771 -893 4783 -859
rect 4867 -893 4879 -859
rect 4771 -899 4879 -893
rect 5032 -854 5226 -832
rect 4410 -982 4421 -943
rect 4197 -1119 4210 -1082
rect 3997 -1169 4105 -1163
rect 3997 -1203 4009 -1169
rect 4093 -1203 4105 -1169
rect 3997 -1209 4105 -1203
rect 4022 -1260 4082 -1209
rect 4150 -1260 4210 -1119
rect 4415 -1119 4421 -982
rect 4455 -982 4470 -943
rect 4673 -943 4719 -931
rect 4455 -1119 4461 -982
rect 4673 -1080 4679 -943
rect 4415 -1131 4461 -1119
rect 4666 -1119 4679 -1080
rect 4713 -1080 4719 -943
rect 4931 -943 4977 -931
rect 4931 -1080 4937 -943
rect 4713 -1119 4726 -1080
rect 4255 -1169 4363 -1163
rect 4255 -1203 4267 -1169
rect 4351 -1203 4363 -1169
rect 4255 -1209 4363 -1203
rect 4513 -1169 4621 -1163
rect 4513 -1203 4525 -1169
rect 4609 -1203 4621 -1169
rect 4513 -1209 4621 -1203
rect 4280 -1260 4340 -1209
rect 4022 -1320 4340 -1260
rect 3886 -1456 3892 -1396
rect 3952 -1456 3958 -1396
rect 4022 -1512 4082 -1320
rect 4150 -1512 4210 -1320
rect 4280 -1512 4340 -1320
rect 4666 -1272 4726 -1119
rect 4922 -1119 4937 -1080
rect 4971 -1080 4977 -943
rect 4971 -1119 4982 -1080
rect 4771 -1169 4879 -1163
rect 4771 -1203 4783 -1169
rect 4867 -1203 4879 -1169
rect 4771 -1209 4879 -1203
rect 4794 -1272 4854 -1209
rect 4922 -1272 4982 -1119
rect 5032 -1208 5052 -854
rect 5086 -1208 5172 -854
rect 5206 -1208 5226 -854
rect 5377 -859 5485 -853
rect 5377 -893 5389 -859
rect 5473 -893 5485 -859
rect 5377 -899 5485 -893
rect 5635 -859 5743 -853
rect 5635 -893 5647 -859
rect 5731 -893 5743 -859
rect 5635 -899 5743 -893
rect 5279 -943 5325 -931
rect 5279 -1082 5285 -943
rect 5032 -1270 5226 -1208
rect 5274 -1119 5285 -1082
rect 5319 -1082 5325 -943
rect 5537 -943 5583 -931
rect 5319 -1119 5334 -1082
rect 5537 -1088 5543 -943
rect 5274 -1270 5334 -1119
rect 5530 -1119 5543 -1088
rect 5577 -1088 5583 -943
rect 5788 -943 5848 -432
rect 6053 -432 6059 -84
rect 6093 -84 6104 -56
rect 6158 44 6222 104
rect 6093 -432 6099 -84
rect 6053 -444 6099 -432
rect 5893 -491 6001 -485
rect 5893 -525 5905 -491
rect 5989 -525 6001 -491
rect 5893 -531 6001 -525
rect 6158 -530 6172 44
rect 6208 -530 6222 44
rect 6158 -542 6222 -530
rect 6158 -852 6226 -834
rect 5893 -859 6001 -853
rect 5893 -893 5905 -859
rect 5989 -893 6001 -859
rect 5893 -899 6001 -893
rect 5788 -970 5801 -943
rect 5577 -1119 5590 -1088
rect 5377 -1169 5485 -1163
rect 5377 -1203 5389 -1169
rect 5473 -1203 5485 -1169
rect 5377 -1209 5485 -1203
rect 5530 -1182 5590 -1119
rect 5795 -1119 5801 -970
rect 5835 -970 5848 -943
rect 6053 -943 6099 -931
rect 5835 -1119 5841 -970
rect 6053 -1094 6059 -943
rect 5795 -1131 5841 -1119
rect 6048 -1119 6059 -1094
rect 6093 -1094 6099 -943
rect 6093 -1119 6108 -1094
rect 5635 -1169 5743 -1163
rect 5402 -1270 5462 -1209
rect 5530 -1248 5592 -1182
rect 5635 -1203 5647 -1169
rect 5731 -1203 5743 -1169
rect 5635 -1209 5743 -1203
rect 5893 -1169 6001 -1163
rect 5893 -1203 5905 -1169
rect 5989 -1203 6001 -1169
rect 5893 -1209 6001 -1203
rect 5032 -1272 5462 -1270
rect 4666 -1330 5462 -1272
rect 4666 -1332 5226 -1330
rect 5032 -1512 5226 -1332
rect 5532 -1392 5592 -1248
rect 5666 -1274 5726 -1209
rect 5660 -1334 5666 -1274
rect 5726 -1334 5732 -1274
rect 5916 -1276 5976 -1209
rect 6048 -1276 6108 -1119
rect 6158 -1208 6174 -852
rect 6208 -1208 6226 -852
rect 6158 -1276 6226 -1208
rect 5532 -1458 5592 -1452
rect 5916 -1336 6226 -1276
rect 5916 -1512 5976 -1336
rect 6048 -1512 6108 -1336
rect 6158 -1512 6226 -1336
rect -2528 -1518 6928 -1512
rect -2528 -1618 -2422 -1518
rect 6822 -1618 6928 -1518
rect -2528 -1624 6928 -1618
rect -2528 -1716 -2416 -1624
rect 3892 -1674 3952 -1670
rect 5532 -1674 5592 -1668
rect 3892 -1676 5532 -1674
rect -2528 -3584 -2522 -1716
rect -2422 -3584 -2416 -1716
rect 2526 -1736 3892 -1676
rect 3952 -1734 5532 -1676
rect -1764 -1848 -48 -1788
rect 12 -1848 18 -1788
rect 1664 -1848 1670 -1788
rect 1730 -1848 1736 -1788
rect -1764 -1996 -1704 -1848
rect -1340 -1906 -1280 -1848
rect -1508 -1912 -1100 -1906
rect -1508 -1946 -1496 -1912
rect -1112 -1946 -1100 -1912
rect -1508 -1952 -1100 -1946
rect -650 -1912 -242 -1906
rect -650 -1946 -638 -1912
rect -254 -1946 -242 -1912
rect -650 -1952 -242 -1946
rect -1764 -2172 -1750 -1996
rect -1716 -2172 -1704 -1996
rect -898 -1996 -852 -1984
rect -898 -2124 -892 -1996
rect -1764 -2344 -1704 -2172
rect -908 -2172 -892 -2124
rect -858 -2124 -852 -1996
rect -48 -1996 12 -1848
rect 208 -1912 616 -1906
rect 208 -1946 220 -1912
rect 604 -1946 616 -1912
rect 208 -1952 616 -1946
rect 1066 -1912 1474 -1906
rect 1066 -1946 1078 -1912
rect 1462 -1946 1474 -1912
rect 1066 -1952 1474 -1946
rect -48 -2042 -34 -1996
rect -858 -2172 -848 -2124
rect -1508 -2222 -1100 -2216
rect -1508 -2256 -1496 -2222
rect -1112 -2256 -1100 -2222
rect -1508 -2262 -1100 -2256
rect -1348 -2344 -1288 -2262
rect -908 -2340 -848 -2172
rect -40 -2172 -34 -2042
rect 0 -2042 12 -1996
rect 818 -1996 864 -1984
rect 0 -2172 6 -2042
rect 818 -2134 824 -1996
rect -40 -2184 6 -2172
rect 810 -2172 824 -2134
rect 858 -2134 864 -1996
rect 1670 -1996 1730 -1848
rect 1924 -1912 2332 -1906
rect 1924 -1946 1936 -1912
rect 2320 -1946 2332 -1912
rect 1924 -1952 2332 -1946
rect 1670 -2032 1682 -1996
rect 858 -2172 870 -2134
rect -650 -2222 -242 -2216
rect -650 -2256 -638 -2222
rect -254 -2256 -242 -2222
rect -650 -2262 -242 -2256
rect 208 -2222 616 -2216
rect 208 -2256 220 -2222
rect 604 -2256 616 -2222
rect 208 -2262 616 -2256
rect -476 -2340 -416 -2262
rect 378 -2340 438 -2262
rect 810 -2340 870 -2172
rect 1676 -2172 1682 -2032
rect 1716 -2032 1730 -1996
rect 2526 -1996 2586 -1736
rect 3892 -1742 3952 -1736
rect 5532 -1740 5592 -1734
rect 6816 -1716 6928 -1624
rect 2944 -1848 2950 -1788
rect 3010 -1848 3016 -1788
rect 3382 -1848 3388 -1788
rect 3448 -1848 3454 -1788
rect 5092 -1848 5098 -1788
rect 5158 -1848 6018 -1788
rect 2950 -1906 3010 -1848
rect 2782 -1912 3190 -1906
rect 2782 -1946 2794 -1912
rect 3178 -1946 3190 -1912
rect 2782 -1952 3190 -1946
rect 2526 -2026 2540 -1996
rect 1716 -2172 1722 -2032
rect 1676 -2184 1722 -2172
rect 2534 -2172 2540 -2026
rect 2574 -2026 2586 -1996
rect 3388 -1996 3448 -1848
rect 3640 -1912 4048 -1906
rect 3640 -1946 3652 -1912
rect 4036 -1946 4048 -1912
rect 3640 -1952 4048 -1946
rect 4498 -1912 4906 -1906
rect 4498 -1946 4510 -1912
rect 4894 -1946 4906 -1912
rect 4498 -1952 4906 -1946
rect 2574 -2172 2580 -2026
rect 3388 -2036 3398 -1996
rect 2534 -2184 2580 -2172
rect 3392 -2172 3398 -2036
rect 3432 -2036 3448 -1996
rect 4250 -1996 4296 -1984
rect 3432 -2172 3438 -2036
rect 4250 -2122 4256 -1996
rect 3392 -2184 3438 -2172
rect 4244 -2172 4256 -2122
rect 4290 -2122 4296 -1996
rect 5098 -1996 5158 -1848
rect 5518 -1906 5578 -1848
rect 5356 -1912 5764 -1906
rect 5356 -1946 5368 -1912
rect 5752 -1946 5764 -1912
rect 5356 -1952 5764 -1946
rect 5098 -2046 5114 -1996
rect 4290 -2172 4304 -2122
rect 1066 -2222 1474 -2216
rect 1066 -2256 1078 -2222
rect 1462 -2256 1474 -2222
rect 1066 -2262 1474 -2256
rect 1924 -2222 2332 -2216
rect 1924 -2256 1936 -2222
rect 2320 -2256 2332 -2222
rect 1924 -2262 2332 -2256
rect 2782 -2222 3190 -2216
rect 2782 -2256 2794 -2222
rect 3178 -2256 3190 -2222
rect 2782 -2262 3190 -2256
rect 3640 -2222 4048 -2216
rect 3640 -2256 3652 -2222
rect 4036 -2256 4048 -2222
rect 3640 -2262 4048 -2256
rect 1230 -2340 1290 -2262
rect 2094 -2340 2154 -2262
rect 3818 -2340 3878 -2262
rect 4244 -2340 4304 -2172
rect 5108 -2172 5114 -2046
rect 5148 -2046 5158 -1996
rect 5958 -1996 6018 -1848
rect 5148 -2172 5154 -2046
rect 5108 -2184 5154 -2172
rect 5958 -2172 5972 -1996
rect 6006 -2172 6018 -1996
rect 4498 -2222 4906 -2216
rect 4498 -2256 4510 -2222
rect 4894 -2256 4906 -2222
rect 4498 -2262 4906 -2256
rect 5356 -2222 5764 -2216
rect 5356 -2256 5368 -2222
rect 5752 -2256 5764 -2222
rect 5356 -2262 5764 -2256
rect 4666 -2340 4726 -2262
rect 5516 -2336 5576 -2262
rect 5958 -2336 6018 -2172
rect -1764 -2404 -1288 -2344
rect -914 -2400 -908 -2340
rect -848 -2400 -842 -2340
rect -482 -2400 -476 -2340
rect -416 -2400 -410 -2340
rect -58 -2400 -52 -2340
rect 8 -2400 14 -2340
rect 372 -2400 378 -2340
rect 438 -2400 444 -2340
rect 804 -2400 810 -2340
rect 870 -2400 876 -2340
rect 1224 -2400 1230 -2340
rect 1290 -2400 1296 -2340
rect 2088 -2400 2094 -2340
rect 2154 -2400 2160 -2340
rect 2944 -2400 2950 -2340
rect 3010 -2400 3016 -2340
rect 3378 -2400 3384 -2340
rect 3444 -2400 3450 -2340
rect 3812 -2400 3818 -2340
rect 3878 -2400 3884 -2340
rect 4238 -2400 4244 -2340
rect 4304 -2400 4310 -2340
rect 4660 -2400 4666 -2340
rect 4726 -2400 4732 -2340
rect 5094 -2400 5100 -2340
rect 5160 -2400 5166 -2340
rect 5516 -2396 6018 -2336
rect -1764 -2578 -1704 -2404
rect -1348 -2488 -1288 -2404
rect -908 -2406 -848 -2400
rect -476 -2488 -416 -2400
rect -1508 -2494 -1100 -2488
rect -1508 -2528 -1496 -2494
rect -1112 -2528 -1100 -2494
rect -1508 -2534 -1100 -2528
rect -650 -2494 -242 -2488
rect -650 -2528 -638 -2494
rect -254 -2528 -242 -2494
rect -650 -2534 -242 -2528
rect -1764 -2754 -1750 -2578
rect -1716 -2754 -1704 -2578
rect -898 -2578 -852 -2566
rect -898 -2722 -892 -2578
rect -1764 -2892 -1704 -2754
rect -906 -2754 -892 -2722
rect -858 -2722 -852 -2578
rect -52 -2578 8 -2400
rect 378 -2488 438 -2400
rect 2094 -2488 2154 -2400
rect 2950 -2488 3010 -2400
rect 208 -2494 616 -2488
rect 208 -2528 220 -2494
rect 604 -2528 616 -2494
rect 208 -2534 616 -2528
rect 1066 -2494 1474 -2488
rect 1066 -2528 1078 -2494
rect 1462 -2528 1474 -2494
rect 1066 -2534 1474 -2528
rect 1924 -2494 2332 -2488
rect 1924 -2528 1936 -2494
rect 2320 -2528 2332 -2494
rect 1924 -2534 2332 -2528
rect 2782 -2494 3190 -2488
rect 2782 -2528 2794 -2494
rect 3178 -2528 3190 -2494
rect 2782 -2534 3190 -2528
rect -52 -2626 -34 -2578
rect -858 -2754 -846 -2722
rect -1508 -2804 -1100 -2798
rect -1508 -2838 -1496 -2804
rect -1112 -2838 -1100 -2804
rect -1508 -2844 -1100 -2838
rect -1340 -2892 -1280 -2844
rect -906 -2892 -846 -2754
rect -40 -2754 -34 -2626
rect 0 -2626 8 -2578
rect 818 -2578 864 -2566
rect 0 -2754 6 -2626
rect 818 -2700 824 -2578
rect -40 -2766 6 -2754
rect 808 -2754 824 -2700
rect 858 -2700 864 -2578
rect 1676 -2578 1722 -2566
rect 1676 -2696 1682 -2578
rect 858 -2754 868 -2700
rect -650 -2804 -242 -2798
rect -650 -2838 -638 -2804
rect -254 -2838 -242 -2804
rect -650 -2844 -242 -2838
rect 208 -2804 616 -2798
rect 208 -2838 220 -2804
rect 604 -2838 616 -2804
rect 208 -2844 616 -2838
rect -1764 -2952 -846 -2892
rect -1764 -3082 -1704 -2952
rect -1340 -3082 -1280 -2952
rect -906 -3082 -846 -2952
rect 808 -2906 868 -2754
rect 1670 -2754 1682 -2696
rect 1716 -2696 1722 -2578
rect 2534 -2578 2580 -2566
rect 1716 -2754 1730 -2696
rect 2534 -2736 2540 -2578
rect 1066 -2804 1474 -2798
rect 1066 -2838 1078 -2804
rect 1462 -2838 1474 -2804
rect 1066 -2844 1474 -2838
rect 1234 -2906 1294 -2844
rect 1670 -2904 1730 -2754
rect 2526 -2754 2540 -2736
rect 2574 -2736 2580 -2578
rect 3384 -2578 3444 -2400
rect 3818 -2488 3878 -2400
rect 4666 -2488 4726 -2400
rect 3640 -2494 4048 -2488
rect 3640 -2528 3652 -2494
rect 4036 -2528 4048 -2494
rect 3640 -2534 4048 -2528
rect 4498 -2494 4906 -2488
rect 4498 -2528 4510 -2494
rect 4894 -2528 4906 -2494
rect 4498 -2534 4906 -2528
rect 3384 -2636 3398 -2578
rect 2574 -2754 2586 -2736
rect 1924 -2804 2332 -2798
rect 1924 -2838 1936 -2804
rect 2320 -2838 2332 -2804
rect 1924 -2844 2332 -2838
rect 808 -2966 1294 -2906
rect 1664 -2964 1670 -2904
rect 1730 -2964 1736 -2904
rect 808 -3082 868 -2966
rect 1234 -3082 1294 -2966
rect 2526 -3082 2586 -2754
rect 3392 -2754 3398 -2636
rect 3432 -2636 3444 -2578
rect 4250 -2578 4296 -2566
rect 3432 -2754 3438 -2636
rect 4250 -2700 4256 -2578
rect 3392 -2766 3438 -2754
rect 4242 -2754 4256 -2700
rect 4290 -2700 4296 -2578
rect 5100 -2578 5160 -2400
rect 5516 -2488 5576 -2396
rect 5356 -2494 5764 -2488
rect 5356 -2528 5368 -2494
rect 5752 -2528 5764 -2494
rect 5356 -2534 5764 -2528
rect 5100 -2618 5114 -2578
rect 4290 -2754 4302 -2700
rect 2782 -2804 3190 -2798
rect 2782 -2838 2794 -2804
rect 3178 -2838 3190 -2804
rect 2782 -2844 3190 -2838
rect 3640 -2804 4048 -2798
rect 3640 -2838 3652 -2804
rect 4036 -2838 4048 -2804
rect 3640 -2844 4048 -2838
rect 4242 -3082 4302 -2754
rect 5108 -2754 5114 -2618
rect 5148 -2618 5160 -2578
rect 5958 -2578 6018 -2396
rect 5148 -2754 5154 -2618
rect 5108 -2766 5154 -2754
rect 5958 -2754 5972 -2578
rect 6006 -2754 6018 -2578
rect 4498 -2804 4906 -2798
rect 4498 -2838 4510 -2804
rect 4894 -2838 4906 -2804
rect 4498 -2844 4906 -2838
rect 5356 -2804 5764 -2798
rect 5356 -2838 5368 -2804
rect 5752 -2838 5764 -2804
rect 5356 -2844 5764 -2838
rect 5516 -2904 5576 -2844
rect 5958 -2904 6018 -2754
rect 5516 -2964 6018 -2904
rect 5516 -3082 5576 -2964
rect 5958 -3082 6018 -2964
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1782 -3122
rect 6080 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2528 -3676 -2416 -3584
rect -1816 -3676 -1806 -3376
rect 6206 -3676 6216 -3376
rect 6816 -3584 6822 -1716
rect 6922 -3584 6928 -1716
rect 6816 -3676 6928 -3584
rect -2528 -3682 6928 -3676
rect -2528 -3782 -2422 -3682
rect 6822 -3782 6928 -3682
rect -2528 -3788 6928 -3782
<< via1 >>
rect -2416 2256 -1816 2556
rect 6216 2256 6816 2556
rect -2302 2030 6694 2140
rect -2298 1774 -2238 1834
rect -1290 1774 -1230 1834
rect 2140 1768 2200 1828
rect -1290 1168 -1230 1228
rect -856 1168 -796 1228
rect -6 1168 54 1228
rect 426 1168 486 1228
rect 856 1168 916 1228
rect 1712 1168 1772 1228
rect 2144 1168 2204 1228
rect 2564 1168 2624 1228
rect -2298 576 -2238 636
rect 5574 1768 5634 1828
rect 6594 1768 6654 1828
rect 3426 1168 3486 1228
rect 3860 1168 3920 1228
rect 4296 1168 4356 1228
rect 5136 1168 5196 1228
rect 5576 1168 5636 1228
rect 426 576 486 636
rect 3856 576 3916 636
rect 6594 576 6654 636
rect 202 -470 262 -464
rect 202 -518 208 -470
rect 208 -518 256 -470
rect 256 -518 262 -470
rect 202 -524 262 -518
rect 4540 98 4600 158
rect 4668 96 4728 156
rect 348 -668 408 -662
rect 348 -710 352 -668
rect 352 -710 400 -668
rect 400 -710 408 -668
rect 348 -722 408 -710
rect 840 -722 900 -662
rect 670 -780 730 -774
rect 670 -828 676 -780
rect 676 -828 724 -780
rect 724 -828 730 -780
rect 670 -834 730 -828
rect 5662 240 5722 300
rect 5532 96 5592 156
rect 3754 -1454 3814 -1394
rect 3892 -1456 3952 -1396
rect 5666 -1334 5726 -1274
rect 5532 -1452 5592 -1392
rect 3892 -1736 3952 -1676
rect 5532 -1734 5592 -1674
rect -48 -1848 12 -1788
rect 1670 -1848 1730 -1788
rect 2950 -1848 3010 -1788
rect 3388 -1848 3448 -1788
rect 5098 -1848 5158 -1788
rect -908 -2400 -848 -2340
rect -476 -2400 -416 -2340
rect -52 -2400 8 -2340
rect 378 -2400 438 -2340
rect 810 -2400 870 -2340
rect 1230 -2400 1290 -2340
rect 2094 -2400 2154 -2340
rect 2950 -2400 3010 -2340
rect 3384 -2400 3444 -2340
rect 3818 -2400 3878 -2340
rect 4244 -2400 4304 -2340
rect 4666 -2400 4726 -2340
rect 5100 -2400 5160 -2340
rect 1670 -2964 1730 -2904
rect -1782 -3266 6080 -3122
rect -2416 -3676 -1816 -3376
rect 6216 -3676 6816 -3376
<< metal2 >>
rect -2416 2556 -1816 2566
rect -2416 2246 -1816 2256
rect 6216 2556 6816 2566
rect 6216 2246 6816 2256
rect -2340 2140 6730 2174
rect -2340 2030 -2302 2140
rect 6694 2030 6730 2140
rect -2340 1992 6730 2030
rect -2298 1834 -2238 1840
rect -1290 1834 -1230 1840
rect -2238 1774 -1290 1834
rect -2298 1768 -2238 1774
rect -1290 1768 -1230 1774
rect 2140 1828 2200 1834
rect 5574 1828 5634 1834
rect 6594 1828 6654 1834
rect 2200 1768 5574 1828
rect 5634 1768 6594 1828
rect 2140 1762 2200 1768
rect 5574 1762 5634 1768
rect 6594 1762 6654 1768
rect -1290 1228 -1230 1234
rect -856 1228 -796 1234
rect -6 1228 54 1234
rect 426 1228 486 1234
rect 856 1228 916 1234
rect 1712 1228 1772 1234
rect 2144 1228 2204 1234
rect 2564 1228 2624 1234
rect 3426 1228 3486 1234
rect 3860 1228 3920 1234
rect 4296 1228 4356 1234
rect 5136 1228 5196 1234
rect 5576 1228 5636 1234
rect -1230 1168 -856 1228
rect -796 1168 -6 1228
rect 54 1168 426 1228
rect 486 1168 856 1228
rect 916 1168 1712 1228
rect 1772 1168 2144 1228
rect 2204 1168 2564 1228
rect 2624 1168 3426 1228
rect 3486 1168 3860 1228
rect 3920 1168 4296 1228
rect 4356 1168 5136 1228
rect 5196 1168 5576 1228
rect 5636 1168 6776 1228
rect -1290 1162 -1230 1168
rect -856 1162 -796 1168
rect -6 1162 54 1168
rect 426 1162 486 1168
rect 856 1162 916 1168
rect 1712 1162 1772 1168
rect 2144 1162 2204 1168
rect 2564 1162 2624 1168
rect 3426 1162 3486 1168
rect 3860 1162 3920 1168
rect 4296 1162 4356 1168
rect 5136 1162 5196 1168
rect 5576 1162 5636 1168
rect -2298 636 -2238 642
rect 426 636 486 642
rect 3856 636 3916 642
rect 6594 636 6654 642
rect -2238 576 426 636
rect 486 576 3856 636
rect 3916 576 6594 636
rect -2298 570 -2238 576
rect 426 570 486 576
rect 3856 570 3916 576
rect 5662 300 5722 306
rect 202 240 5662 300
rect 202 -464 262 240
rect 5662 234 5722 240
rect 4540 158 4600 164
rect 348 98 4540 158
rect 196 -524 202 -464
rect 262 -524 268 -464
rect 348 -662 408 98
rect 4540 92 4600 98
rect 4668 156 4728 162
rect 5532 156 5592 162
rect 5802 156 5862 576
rect 6594 570 6654 576
rect 4728 96 5532 156
rect 5592 96 5862 156
rect 4668 90 4728 96
rect 5532 90 5592 96
rect 6716 32 6776 1168
rect 6378 -28 6776 32
rect 342 -722 348 -662
rect 408 -722 414 -662
rect 834 -722 840 -662
rect 900 -722 906 -662
rect 664 -834 670 -774
rect 730 -834 736 -774
rect 670 -1394 730 -834
rect 840 -1050 900 -722
rect 840 -1110 3214 -1050
rect 3154 -1274 3214 -1110
rect 5666 -1274 5726 -1268
rect 3154 -1334 5666 -1274
rect 5666 -1340 5726 -1334
rect 3754 -1394 3814 -1388
rect 670 -1454 3754 -1394
rect 3754 -1460 3814 -1454
rect 3892 -1396 3952 -1390
rect 5526 -1452 5532 -1392
rect 5592 -1452 5598 -1392
rect 3892 -1676 3952 -1456
rect 5532 -1674 5592 -1452
rect 3886 -1736 3892 -1676
rect 3952 -1736 3958 -1676
rect 5526 -1734 5532 -1674
rect 5592 -1734 5598 -1674
rect -48 -1788 12 -1782
rect 1670 -1788 1730 -1782
rect 2950 -1788 3010 -1782
rect 3388 -1788 3448 -1782
rect 5098 -1788 5158 -1782
rect 12 -1848 1670 -1788
rect 1730 -1848 2950 -1788
rect 3010 -1848 3388 -1788
rect 3448 -1848 5098 -1788
rect -48 -1854 12 -1848
rect 1670 -1854 1730 -1848
rect 2950 -1854 3010 -1848
rect 3388 -1854 3448 -1848
rect 5098 -1854 5158 -1848
rect -908 -2340 -848 -2334
rect -476 -2340 -416 -2334
rect -52 -2340 8 -2334
rect 378 -2340 438 -2334
rect 810 -2340 870 -2334
rect 1230 -2340 1290 -2334
rect 2094 -2340 2154 -2334
rect 2950 -2340 3010 -2334
rect 3384 -2340 3444 -2334
rect 3818 -2340 3878 -2334
rect 4244 -2340 4304 -2334
rect 4666 -2340 4726 -2334
rect 5100 -2340 5160 -2334
rect -848 -2400 -476 -2340
rect -416 -2400 -52 -2340
rect 8 -2400 378 -2340
rect 438 -2400 810 -2340
rect 870 -2400 1230 -2340
rect 1290 -2400 2094 -2340
rect 2154 -2400 2950 -2340
rect 3010 -2400 3384 -2340
rect 3444 -2400 3818 -2340
rect 3878 -2400 4244 -2340
rect 4304 -2400 4666 -2340
rect 4726 -2400 5100 -2340
rect -908 -2406 -848 -2400
rect -476 -2406 -416 -2400
rect -52 -2406 8 -2400
rect 378 -2406 438 -2400
rect 810 -2406 870 -2400
rect 1230 -2406 1290 -2400
rect 2094 -2406 2154 -2400
rect 2950 -2406 3010 -2400
rect 3384 -2406 3444 -2400
rect 3818 -2406 3878 -2400
rect 4244 -2406 4304 -2400
rect 4666 -2406 4726 -2400
rect 5100 -2406 5160 -2400
rect 1670 -2904 1730 -2898
rect 6378 -2904 6438 -28
rect 1730 -2964 6438 -2904
rect 1670 -2970 1730 -2964
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1782 -3122
rect 6080 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2416 -3376 -1816 -3366
rect -2416 -3686 -1816 -3676
rect 6216 -3376 6816 -3366
rect 6216 -3686 6816 -3676
<< via2 >>
rect -2416 2256 -1816 2556
rect 6216 2256 6816 2556
rect -2302 2030 6694 2140
rect -1782 -3266 6080 -3122
rect -2416 -3676 -1816 -3376
rect 6216 -3676 6816 -3376
<< metal3 >>
rect -2426 2556 -1806 2561
rect -2426 2256 -2416 2556
rect -1816 2256 -1806 2556
rect -2426 2251 -1806 2256
rect 6206 2556 6826 2561
rect 6206 2256 6216 2556
rect 6816 2256 6826 2556
rect 6206 2251 6826 2256
rect -2340 2140 6730 2174
rect -2340 2030 -2302 2140
rect 6694 2030 6730 2140
rect -2340 1992 6730 2030
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1782 -3122
rect 6080 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2426 -3376 -1806 -3371
rect -2426 -3676 -2416 -3376
rect -1816 -3676 -1806 -3376
rect -2426 -3681 -1806 -3676
rect 6206 -3376 6826 -3371
rect 6206 -3676 6216 -3376
rect 6816 -3676 6826 -3376
rect 6206 -3681 6826 -3676
<< via3 >>
rect -2416 2256 -1816 2556
rect 6216 2256 6816 2556
rect -2302 2030 6694 2140
rect -1782 -3266 6080 -3122
rect -2416 -3676 -1816 -3376
rect 6216 -3676 6816 -3376
<< metal4 >>
rect -2600 2556 7000 2740
rect -2600 2256 -2416 2556
rect -1816 2256 6216 2556
rect 6816 2256 7000 2556
rect -2600 2140 7000 2256
rect -2600 2030 -2302 2140
rect 6694 2030 7000 2140
rect -2600 1940 7000 2030
rect -2600 -3122 7000 -3060
rect -2600 -3266 -1782 -3122
rect 6080 -3266 7000 -3122
rect -2600 -3376 7000 -3266
rect -2600 -3676 -2416 -3376
rect -1816 -3676 6216 -3376
rect 6816 -3676 7000 -3376
rect -2600 -3860 7000 -3676
<< labels >>
flabel metal1 2548 -1880 2560 -1874 1 FreeSans 480 0 0 0 vswitchl
flabel metal2 1694 -2378 1704 -2366 1 FreeSans 480 0 0 0 ibiasn
port 6 n
flabel metal1 3656 -862 3666 -854 1 FreeSans 480 0 0 0 vpdiode
flabel metal1 5552 -1226 5564 -1208 1 FreeSans 480 0 0 0 vswitchl
flabel metal2 4962 114 4976 132 1 FreeSans 480 0 0 0 vswitchh
flabel metal2 1104 596 1120 610 1 FreeSans 480 0 0 0 vswitchh
flabel metal1 5812 -840 5822 -830 1 FreeSans 480 0 0 0 vcp
port 5 n
flabel metal1 620 -692 624 -688 1 FreeSans 480 0 0 0 vQB
flabel metal1 294 -700 300 -692 1 FreeSans 480 0 0 0 vQA
flabel metal1 -2200 -692 -2194 -688 1 FreeSans 480 0 0 0 vsig_in
port 4 n
flabel metal1 3070 -680 3078 -676 1 FreeSans 480 0 0 0 vin_div
port 3 n
flabel metal1 300 -592 304 -588 1 FreeSans 480 0 0 0 vRSTN
flabel metal2 944 -1420 952 -1412 1 FreeSans 480 0 0 0 VQBb
flabel metal2 220 -146 228 -138 1 FreeSans 480 0 0 0 vQAb
flabel metal2 1582 1194 1598 1204 1 FreeSans 480 0 0 0 vpbias
flabel metal2 2204 -2944 2214 -2936 1 FreeSans 480 0 0 0 vpbias
flabel metal4 886 2206 898 2222 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel metal4 1252 -3422 1278 -3396 1 FreeSans 480 0 0 0 VSS
port 2 n ground bidirectional
flabel metal1 4436 -580 4442 -570 1 FreeSans 480 0 0 0 vndiode
flabel locali 216 -635 250 -601 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali 216 -703 250 -669 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali 124 -703 158 -669 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/A
flabel nwell 81 -397 115 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell 81 -941 115 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 81 -941 115 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 81 -397 115 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment 52 -924 52 -924 4 sky130_fd_sc_hd__inv_1_1/inv_1
flabel locali 682 -635 716 -601 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 682 -703 716 -669 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 774 -703 808 -669 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 817 -397 851 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 817 -941 851 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 817 -941 851 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 817 -397 851 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 880 -924 880 -924 6 sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali -310 -706 -281 -671 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/Q
flabel locali -8 -703 14 -670 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/Q_N
flabel locali -583 -771 -549 -737 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali -1759 -635 -1725 -601 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/D
flabel locali -2034 -635 -2000 -601 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali -2034 -703 -2000 -669 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali -583 -703 -549 -669 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel metal1 -2035 -941 -2001 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VGND
flabel metal1 -2035 -397 -2001 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VPWR
flabel nwell -2035 -397 -2001 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VPB
flabel pwell -2035 -941 -2001 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VNB
rlabel comment -2064 -924 -2064 -924 4 sky130_fd_sc_hd__dfrbp_1_1/dfrbp_1
rlabel viali -583 -771 -549 -737 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel viali -643 -708 -609 -674 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali -583 -797 -535 -717 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali -643 -717 -535 -643 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 -595 -777 -537 -768 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 -655 -731 -597 -668 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 -655 -740 -537 -731 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 -1315 -740 -1185 -731 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 -1315 -768 -537 -740 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 -1315 -777 -1185 -768 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 1213 -706 1242 -671 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/Q
flabel locali 918 -703 940 -670 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/Q_N
flabel locali 1481 -771 1515 -737 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 2657 -635 2691 -601 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/D
flabel locali 2932 -635 2966 -601 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 2932 -703 2966 -669 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 1481 -703 1515 -669 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel metal1 2933 -941 2967 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VGND
flabel metal1 2933 -397 2967 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VPWR
flabel nwell 2933 -397 2967 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VPB
flabel pwell 2933 -941 2967 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VNB
rlabel comment 2996 -924 2996 -924 6 sky130_fd_sc_hd__dfrbp_1_0/dfrbp_1
rlabel viali 1481 -771 1515 -737 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel viali 1541 -708 1575 -674 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 1467 -797 1515 -717 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 1467 -717 1575 -643 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1469 -777 1527 -768 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1529 -731 1587 -668 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1469 -740 1587 -731 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 2117 -740 2247 -731 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1469 -768 2247 -740 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 2117 -777 2247 -768 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 450 -839 484 -805 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 450 -771 484 -737 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 450 -703 484 -669 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 542 -703 576 -669 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/B
flabel locali 358 -703 392 -669 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/A
flabel nwell 542 -397 576 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell 542 -941 576 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 542 -941 576 -907 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 542 -397 576 -363 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment 604 -924 604 -924 6 sky130_fd_sc_hd__nand2_1_0/nand2_1
<< end >>
