magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 17 199 86 323
rect 194 265 261 339
rect 194 199 286 265
rect 399 289 1915 345
rect 194 124 261 199
rect 1865 171 1915 289
rect 1255 123 1915 171
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 357 89 527
rect 123 323 160 493
rect 194 373 261 527
rect 120 199 160 323
rect 17 17 89 165
rect 123 56 160 199
rect 295 299 365 493
rect 399 413 449 493
rect 483 447 549 527
rect 583 413 617 493
rect 651 447 717 527
rect 751 413 785 493
rect 819 447 885 527
rect 919 413 953 493
rect 987 447 1053 527
rect 1087 413 1915 493
rect 399 379 1915 413
rect 320 255 365 299
rect 320 205 1185 255
rect 1235 205 1831 255
rect 320 165 397 205
rect 194 17 261 89
rect 295 51 397 165
rect 431 131 1221 171
rect 431 51 497 131
rect 531 17 597 97
rect 631 55 665 131
rect 699 17 765 97
rect 799 51 833 131
rect 867 17 933 97
rect 967 55 1001 131
rect 1035 17 1101 97
rect 1135 89 1221 131
rect 1135 51 1915 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 109 252 167 261
rect 1304 252 1362 261
rect 109 224 1362 252
rect 109 215 167 224
rect 1304 215 1362 224
<< labels >>
rlabel locali s 17 199 86 323 6 A
port 1 nsew signal input
rlabel locali s 194 265 261 339 6 TE_B
port 2 nsew signal input
rlabel locali s 194 199 286 265 6 TE_B
port 2 nsew signal input
rlabel locali s 194 124 261 199 6 TE_B
port 2 nsew signal input
rlabel locali s 1865 171 1915 289 6 Z
port 3 nsew signal output
rlabel locali s 1255 123 1915 171 6 Z
port 3 nsew signal output
rlabel locali s 399 289 1915 345 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
