magic
tech sky130A
magscale 1 2
timestamp 1624182449
<< nwell >>
rect 11292 15986 35808 30728
rect 52292 15986 76808 30728
rect 36584 12390 38738 14006
<< pwell >>
rect -1408 -888 35908 15228
rect 39592 -888 76908 15228
<< nmos >>
rect 13578 13734 14538 14334
rect 14596 13734 15556 14334
rect 15614 13734 16574 14334
rect 16632 13734 17592 14334
rect 17650 13734 18610 14334
rect 18668 13734 19628 14334
rect 19686 13734 20646 14334
rect 20704 13734 21664 14334
rect 21722 13734 22682 14334
rect 22740 13734 23700 14334
rect 23758 13734 24718 14334
rect 24776 13734 25736 14334
rect 25794 13734 26754 14334
rect 26812 13734 27772 14334
rect 27830 13734 28790 14334
rect 28848 13734 29808 14334
rect 29866 13734 30826 14334
rect 30884 13734 31844 14334
rect 31902 13734 32862 14334
rect 32920 13734 33880 14334
rect 13578 12916 14538 13516
rect 14596 12916 15556 13516
rect 15614 12916 16574 13516
rect 16632 12916 17592 13516
rect 17650 12916 18610 13516
rect 18668 12916 19628 13516
rect 19686 12916 20646 13516
rect 20704 12916 21664 13516
rect 21722 12916 22682 13516
rect 22740 12916 23700 13516
rect 23758 12916 24718 13516
rect 24776 12916 25736 13516
rect 25794 12916 26754 13516
rect 26812 12916 27772 13516
rect 27830 12916 28790 13516
rect 28848 12916 29808 13516
rect 29866 12916 30826 13516
rect 30884 12916 31844 13516
rect 31902 12916 32862 13516
rect 32920 12916 33880 13516
rect 13578 11538 14538 12138
rect 14596 11538 15556 12138
rect 15614 11538 16574 12138
rect 16632 11538 17592 12138
rect 17650 11538 18610 12138
rect 18668 11538 19628 12138
rect 19686 11538 20646 12138
rect 20704 11538 21664 12138
rect 21722 11538 22682 12138
rect 22740 11538 23700 12138
rect 23758 11538 24718 12138
rect 24776 11538 25736 12138
rect 25794 11538 26754 12138
rect 26812 11538 27772 12138
rect 27830 11538 28790 12138
rect 28848 11538 29808 12138
rect 29866 11538 30826 12138
rect 30884 11538 31844 12138
rect 31902 11538 32862 12138
rect 32920 11538 33880 12138
rect 13578 10306 14538 10906
rect 14596 10306 15556 10906
rect 15614 10306 16574 10906
rect 16632 10306 17592 10906
rect 17650 10306 18610 10906
rect 18668 10306 19628 10906
rect 19686 10306 20646 10906
rect 20704 10306 21664 10906
rect 21722 10306 22682 10906
rect 22740 10306 23700 10906
rect 23758 10306 24718 10906
rect 24776 10306 25736 10906
rect 25794 10306 26754 10906
rect 26812 10306 27772 10906
rect 27830 10306 28790 10906
rect 28848 10306 29808 10906
rect 29866 10306 30826 10906
rect 30884 10306 31844 10906
rect 31902 10306 32862 10906
rect 32920 10306 33880 10906
rect 13576 9072 14536 9672
rect 14594 9072 15554 9672
rect 15612 9072 16572 9672
rect 16630 9072 17590 9672
rect 17648 9072 18608 9672
rect 18666 9072 19626 9672
rect 19684 9072 20644 9672
rect 20702 9072 21662 9672
rect 21720 9072 22680 9672
rect 22738 9072 23698 9672
rect 23756 9072 24716 9672
rect 24774 9072 25734 9672
rect 25792 9072 26752 9672
rect 26810 9072 27770 9672
rect 27828 9072 28788 9672
rect 28846 9072 29806 9672
rect 29864 9072 30824 9672
rect 30882 9072 31842 9672
rect 31900 9072 32860 9672
rect 32918 9072 33878 9672
rect 13576 7838 14536 8438
rect 14594 7838 15554 8438
rect 15612 7838 16572 8438
rect 16630 7838 17590 8438
rect 17648 7838 18608 8438
rect 18666 7838 19626 8438
rect 19684 7838 20644 8438
rect 20702 7838 21662 8438
rect 21720 7838 22680 8438
rect 22738 7838 23698 8438
rect 23756 7838 24716 8438
rect 24774 7838 25734 8438
rect 25792 7838 26752 8438
rect 26810 7838 27770 8438
rect 27828 7838 28788 8438
rect 28846 7838 29806 8438
rect 29864 7838 30824 8438
rect 30882 7838 31842 8438
rect 31900 7838 32860 8438
rect 32918 7838 33878 8438
rect 13576 6606 14536 7206
rect 14594 6606 15554 7206
rect 15612 6606 16572 7206
rect 16630 6606 17590 7206
rect 17648 6606 18608 7206
rect 18666 6606 19626 7206
rect 19684 6606 20644 7206
rect 20702 6606 21662 7206
rect 21720 6606 22680 7206
rect 22738 6606 23698 7206
rect 23756 6606 24716 7206
rect 24774 6606 25734 7206
rect 25792 6606 26752 7206
rect 26810 6606 27770 7206
rect 27828 6606 28788 7206
rect 28846 6606 29806 7206
rect 29864 6606 30824 7206
rect 30882 6606 31842 7206
rect 31900 6606 32860 7206
rect 32918 6606 33878 7206
rect 13576 5372 14536 5972
rect 14594 5372 15554 5972
rect 15612 5372 16572 5972
rect 16630 5372 17590 5972
rect 17648 5372 18608 5972
rect 18666 5372 19626 5972
rect 19684 5372 20644 5972
rect 20702 5372 21662 5972
rect 21720 5372 22680 5972
rect 22738 5372 23698 5972
rect 23756 5372 24716 5972
rect 24774 5372 25734 5972
rect 25792 5372 26752 5972
rect 26810 5372 27770 5972
rect 27828 5372 28788 5972
rect 28846 5372 29806 5972
rect 29864 5372 30824 5972
rect 30882 5372 31842 5972
rect 31900 5372 32860 5972
rect 32918 5372 33878 5972
rect 13576 4138 14536 4738
rect 14594 4138 15554 4738
rect 15612 4138 16572 4738
rect 16630 4138 17590 4738
rect 17648 4138 18608 4738
rect 18666 4138 19626 4738
rect 19684 4138 20644 4738
rect 20702 4138 21662 4738
rect 21720 4138 22680 4738
rect 22738 4138 23698 4738
rect 23756 4138 24716 4738
rect 24774 4138 25734 4738
rect 25792 4138 26752 4738
rect 26810 4138 27770 4738
rect 27828 4138 28788 4738
rect 28846 4138 29806 4738
rect 29864 4138 30824 4738
rect 30882 4138 31842 4738
rect 31900 4138 32860 4738
rect 32918 4138 33878 4738
rect 13576 2906 14536 3506
rect 14594 2906 15554 3506
rect 15612 2906 16572 3506
rect 16630 2906 17590 3506
rect 17648 2906 18608 3506
rect 18666 2906 19626 3506
rect 19684 2906 20644 3506
rect 20702 2906 21662 3506
rect 21720 2906 22680 3506
rect 22738 2906 23698 3506
rect 23756 2906 24716 3506
rect 24774 2906 25734 3506
rect 25792 2906 26752 3506
rect 26810 2906 27770 3506
rect 27828 2906 28788 3506
rect 28846 2906 29806 3506
rect 29864 2906 30824 3506
rect 30882 2906 31842 3506
rect 31900 2906 32860 3506
rect 32918 2906 33878 3506
rect 13576 1672 14536 2272
rect 14594 1672 15554 2272
rect 15612 1672 16572 2272
rect 16630 1672 17590 2272
rect 17648 1672 18608 2272
rect 18666 1672 19626 2272
rect 19684 1672 20644 2272
rect 20702 1672 21662 2272
rect 21720 1672 22680 2272
rect 22738 1672 23698 2272
rect 23756 1672 24716 2272
rect 24774 1672 25734 2272
rect 25792 1672 26752 2272
rect 26810 1672 27770 2272
rect 27828 1672 28788 2272
rect 28846 1672 29806 2272
rect 29864 1672 30824 2272
rect 30882 1672 31842 2272
rect 31900 1672 32860 2272
rect 32918 1672 33878 2272
rect 946 630 1906 1230
rect 1964 630 2924 1230
rect 2982 630 3942 1230
rect 4000 630 4960 1230
rect 5018 630 5978 1230
rect 6036 630 6996 1230
rect 7054 630 8014 1230
rect 8072 630 9032 1230
rect 9090 630 10050 1230
rect 10108 630 11068 1230
rect 13576 440 14536 1040
rect 14594 440 15554 1040
rect 15612 440 16572 1040
rect 16630 440 17590 1040
rect 17648 440 18608 1040
rect 18666 440 19626 1040
rect 19684 440 20644 1040
rect 20702 440 21662 1040
rect 21720 440 22680 1040
rect 22738 440 23698 1040
rect 23756 440 24716 1040
rect 24774 440 25734 1040
rect 25792 440 26752 1040
rect 26810 440 27770 1040
rect 27828 440 28788 1040
rect 28846 440 29806 1040
rect 29864 440 30824 1040
rect 30882 440 31842 1040
rect 31900 440 32860 1040
rect 32918 440 33878 1040
rect -1028 72 -998 202
rect 54578 13734 55538 14334
rect 55596 13734 56556 14334
rect 56614 13734 57574 14334
rect 57632 13734 58592 14334
rect 58650 13734 59610 14334
rect 59668 13734 60628 14334
rect 60686 13734 61646 14334
rect 61704 13734 62664 14334
rect 62722 13734 63682 14334
rect 63740 13734 64700 14334
rect 64758 13734 65718 14334
rect 65776 13734 66736 14334
rect 66794 13734 67754 14334
rect 67812 13734 68772 14334
rect 68830 13734 69790 14334
rect 69848 13734 70808 14334
rect 70866 13734 71826 14334
rect 71884 13734 72844 14334
rect 72902 13734 73862 14334
rect 73920 13734 74880 14334
rect 54578 12916 55538 13516
rect 55596 12916 56556 13516
rect 56614 12916 57574 13516
rect 57632 12916 58592 13516
rect 58650 12916 59610 13516
rect 59668 12916 60628 13516
rect 60686 12916 61646 13516
rect 61704 12916 62664 13516
rect 62722 12916 63682 13516
rect 63740 12916 64700 13516
rect 64758 12916 65718 13516
rect 65776 12916 66736 13516
rect 66794 12916 67754 13516
rect 67812 12916 68772 13516
rect 68830 12916 69790 13516
rect 69848 12916 70808 13516
rect 70866 12916 71826 13516
rect 71884 12916 72844 13516
rect 72902 12916 73862 13516
rect 73920 12916 74880 13516
rect 54578 11538 55538 12138
rect 55596 11538 56556 12138
rect 56614 11538 57574 12138
rect 57632 11538 58592 12138
rect 58650 11538 59610 12138
rect 59668 11538 60628 12138
rect 60686 11538 61646 12138
rect 61704 11538 62664 12138
rect 62722 11538 63682 12138
rect 63740 11538 64700 12138
rect 64758 11538 65718 12138
rect 65776 11538 66736 12138
rect 66794 11538 67754 12138
rect 67812 11538 68772 12138
rect 68830 11538 69790 12138
rect 69848 11538 70808 12138
rect 70866 11538 71826 12138
rect 71884 11538 72844 12138
rect 72902 11538 73862 12138
rect 73920 11538 74880 12138
rect 54578 10306 55538 10906
rect 55596 10306 56556 10906
rect 56614 10306 57574 10906
rect 57632 10306 58592 10906
rect 58650 10306 59610 10906
rect 59668 10306 60628 10906
rect 60686 10306 61646 10906
rect 61704 10306 62664 10906
rect 62722 10306 63682 10906
rect 63740 10306 64700 10906
rect 64758 10306 65718 10906
rect 65776 10306 66736 10906
rect 66794 10306 67754 10906
rect 67812 10306 68772 10906
rect 68830 10306 69790 10906
rect 69848 10306 70808 10906
rect 70866 10306 71826 10906
rect 71884 10306 72844 10906
rect 72902 10306 73862 10906
rect 73920 10306 74880 10906
rect 54576 9072 55536 9672
rect 55594 9072 56554 9672
rect 56612 9072 57572 9672
rect 57630 9072 58590 9672
rect 58648 9072 59608 9672
rect 59666 9072 60626 9672
rect 60684 9072 61644 9672
rect 61702 9072 62662 9672
rect 62720 9072 63680 9672
rect 63738 9072 64698 9672
rect 64756 9072 65716 9672
rect 65774 9072 66734 9672
rect 66792 9072 67752 9672
rect 67810 9072 68770 9672
rect 68828 9072 69788 9672
rect 69846 9072 70806 9672
rect 70864 9072 71824 9672
rect 71882 9072 72842 9672
rect 72900 9072 73860 9672
rect 73918 9072 74878 9672
rect 54576 7838 55536 8438
rect 55594 7838 56554 8438
rect 56612 7838 57572 8438
rect 57630 7838 58590 8438
rect 58648 7838 59608 8438
rect 59666 7838 60626 8438
rect 60684 7838 61644 8438
rect 61702 7838 62662 8438
rect 62720 7838 63680 8438
rect 63738 7838 64698 8438
rect 64756 7838 65716 8438
rect 65774 7838 66734 8438
rect 66792 7838 67752 8438
rect 67810 7838 68770 8438
rect 68828 7838 69788 8438
rect 69846 7838 70806 8438
rect 70864 7838 71824 8438
rect 71882 7838 72842 8438
rect 72900 7838 73860 8438
rect 73918 7838 74878 8438
rect 54576 6606 55536 7206
rect 55594 6606 56554 7206
rect 56612 6606 57572 7206
rect 57630 6606 58590 7206
rect 58648 6606 59608 7206
rect 59666 6606 60626 7206
rect 60684 6606 61644 7206
rect 61702 6606 62662 7206
rect 62720 6606 63680 7206
rect 63738 6606 64698 7206
rect 64756 6606 65716 7206
rect 65774 6606 66734 7206
rect 66792 6606 67752 7206
rect 67810 6606 68770 7206
rect 68828 6606 69788 7206
rect 69846 6606 70806 7206
rect 70864 6606 71824 7206
rect 71882 6606 72842 7206
rect 72900 6606 73860 7206
rect 73918 6606 74878 7206
rect 54576 5372 55536 5972
rect 55594 5372 56554 5972
rect 56612 5372 57572 5972
rect 57630 5372 58590 5972
rect 58648 5372 59608 5972
rect 59666 5372 60626 5972
rect 60684 5372 61644 5972
rect 61702 5372 62662 5972
rect 62720 5372 63680 5972
rect 63738 5372 64698 5972
rect 64756 5372 65716 5972
rect 65774 5372 66734 5972
rect 66792 5372 67752 5972
rect 67810 5372 68770 5972
rect 68828 5372 69788 5972
rect 69846 5372 70806 5972
rect 70864 5372 71824 5972
rect 71882 5372 72842 5972
rect 72900 5372 73860 5972
rect 73918 5372 74878 5972
rect 54576 4138 55536 4738
rect 55594 4138 56554 4738
rect 56612 4138 57572 4738
rect 57630 4138 58590 4738
rect 58648 4138 59608 4738
rect 59666 4138 60626 4738
rect 60684 4138 61644 4738
rect 61702 4138 62662 4738
rect 62720 4138 63680 4738
rect 63738 4138 64698 4738
rect 64756 4138 65716 4738
rect 65774 4138 66734 4738
rect 66792 4138 67752 4738
rect 67810 4138 68770 4738
rect 68828 4138 69788 4738
rect 69846 4138 70806 4738
rect 70864 4138 71824 4738
rect 71882 4138 72842 4738
rect 72900 4138 73860 4738
rect 73918 4138 74878 4738
rect 54576 2906 55536 3506
rect 55594 2906 56554 3506
rect 56612 2906 57572 3506
rect 57630 2906 58590 3506
rect 58648 2906 59608 3506
rect 59666 2906 60626 3506
rect 60684 2906 61644 3506
rect 61702 2906 62662 3506
rect 62720 2906 63680 3506
rect 63738 2906 64698 3506
rect 64756 2906 65716 3506
rect 65774 2906 66734 3506
rect 66792 2906 67752 3506
rect 67810 2906 68770 3506
rect 68828 2906 69788 3506
rect 69846 2906 70806 3506
rect 70864 2906 71824 3506
rect 71882 2906 72842 3506
rect 72900 2906 73860 3506
rect 73918 2906 74878 3506
rect 54576 1672 55536 2272
rect 55594 1672 56554 2272
rect 56612 1672 57572 2272
rect 57630 1672 58590 2272
rect 58648 1672 59608 2272
rect 59666 1672 60626 2272
rect 60684 1672 61644 2272
rect 61702 1672 62662 2272
rect 62720 1672 63680 2272
rect 63738 1672 64698 2272
rect 64756 1672 65716 2272
rect 65774 1672 66734 2272
rect 66792 1672 67752 2272
rect 67810 1672 68770 2272
rect 68828 1672 69788 2272
rect 69846 1672 70806 2272
rect 70864 1672 71824 2272
rect 71882 1672 72842 2272
rect 72900 1672 73860 2272
rect 73918 1672 74878 2272
rect 41946 630 42906 1230
rect 42964 630 43924 1230
rect 43982 630 44942 1230
rect 45000 630 45960 1230
rect 46018 630 46978 1230
rect 47036 630 47996 1230
rect 48054 630 49014 1230
rect 49072 630 50032 1230
rect 50090 630 51050 1230
rect 51108 630 52068 1230
rect 54576 440 55536 1040
rect 55594 440 56554 1040
rect 56612 440 57572 1040
rect 57630 440 58590 1040
rect 58648 440 59608 1040
rect 59666 440 60626 1040
rect 60684 440 61644 1040
rect 61702 440 62662 1040
rect 62720 440 63680 1040
rect 63738 440 64698 1040
rect 64756 440 65716 1040
rect 65774 440 66734 1040
rect 66792 440 67752 1040
rect 67810 440 68770 1040
rect 68828 440 69788 1040
rect 69846 440 70806 1040
rect 70864 440 71824 1040
rect 71882 440 72842 1040
rect 72900 440 73860 1040
rect 73918 440 74878 1040
<< pmos >>
rect 18470 20698 19430 21298
rect 19488 20698 20448 21298
rect 20506 20698 21466 21298
rect 21524 20698 22484 21298
rect 22542 20698 23502 21298
rect 23560 20698 24520 21298
rect 24578 20698 25538 21298
rect 25596 20698 26556 21298
rect 26614 20698 27574 21298
rect 27632 20698 28592 21298
rect 28650 20698 29610 21298
rect 29668 20698 30628 21298
rect 30686 20698 31646 21298
rect 31704 20698 32664 21298
rect 32722 20698 33682 21298
rect 18470 19442 19430 20042
rect 19488 19442 20448 20042
rect 20506 19442 21466 20042
rect 21524 19442 22484 20042
rect 22542 19442 23502 20042
rect 23560 19442 24520 20042
rect 24578 19442 25538 20042
rect 25596 19442 26556 20042
rect 26614 19442 27574 20042
rect 27632 19442 28592 20042
rect 28650 19442 29610 20042
rect 29668 19442 30628 20042
rect 30686 19442 31646 20042
rect 31704 19442 32664 20042
rect 32722 19442 33682 20042
rect 18470 18186 19430 18786
rect 19488 18186 20448 18786
rect 20506 18186 21466 18786
rect 21524 18186 22484 18786
rect 22542 18186 23502 18786
rect 23560 18186 24520 18786
rect 24578 18186 25538 18786
rect 25596 18186 26556 18786
rect 26614 18186 27574 18786
rect 27632 18186 28592 18786
rect 28650 18186 29610 18786
rect 29668 18186 30628 18786
rect 30686 18186 31646 18786
rect 31704 18186 32664 18786
rect 32722 18186 33682 18786
rect 18470 16930 19430 17530
rect 19488 16930 20448 17530
rect 20506 16930 21466 17530
rect 21524 16930 22484 17530
rect 22542 16930 23502 17530
rect 23560 16930 24520 17530
rect 24578 16930 25538 17530
rect 25596 16930 26556 17530
rect 26614 16930 27574 17530
rect 27632 16930 28592 17530
rect 28650 16930 29610 17530
rect 29668 16930 30628 17530
rect 30686 16930 31646 17530
rect 31704 16930 32664 17530
rect 32722 16930 33682 17530
rect 59470 20698 60430 21298
rect 60488 20698 61448 21298
rect 61506 20698 62466 21298
rect 62524 20698 63484 21298
rect 63542 20698 64502 21298
rect 64560 20698 65520 21298
rect 65578 20698 66538 21298
rect 66596 20698 67556 21298
rect 67614 20698 68574 21298
rect 68632 20698 69592 21298
rect 69650 20698 70610 21298
rect 70668 20698 71628 21298
rect 71686 20698 72646 21298
rect 72704 20698 73664 21298
rect 73722 20698 74682 21298
rect 59470 19442 60430 20042
rect 60488 19442 61448 20042
rect 61506 19442 62466 20042
rect 62524 19442 63484 20042
rect 63542 19442 64502 20042
rect 64560 19442 65520 20042
rect 65578 19442 66538 20042
rect 66596 19442 67556 20042
rect 67614 19442 68574 20042
rect 68632 19442 69592 20042
rect 69650 19442 70610 20042
rect 70668 19442 71628 20042
rect 71686 19442 72646 20042
rect 72704 19442 73664 20042
rect 73722 19442 74682 20042
rect 59470 18186 60430 18786
rect 60488 18186 61448 18786
rect 61506 18186 62466 18786
rect 62524 18186 63484 18786
rect 63542 18186 64502 18786
rect 64560 18186 65520 18786
rect 65578 18186 66538 18786
rect 66596 18186 67556 18786
rect 67614 18186 68574 18786
rect 68632 18186 69592 18786
rect 69650 18186 70610 18786
rect 70668 18186 71628 18786
rect 71686 18186 72646 18786
rect 72704 18186 73664 18786
rect 73722 18186 74682 18786
rect 59470 16930 60430 17530
rect 60488 16930 61448 17530
rect 61506 16930 62466 17530
rect 62524 16930 63484 17530
rect 63542 16930 64502 17530
rect 64560 16930 65520 17530
rect 65578 16930 66538 17530
rect 66596 16930 67556 17530
rect 67614 16930 68574 17530
rect 68632 16930 69592 17530
rect 69650 16930 70610 17530
rect 70668 16930 71628 17530
rect 71686 16930 72646 17530
rect 72704 16930 73664 17530
rect 73722 16930 74682 17530
rect 36956 12798 37156 12998
rect 37214 12798 37414 12998
rect 37472 12798 37672 12998
rect 37730 12798 37930 12998
rect 37988 12798 38188 12998
rect 38246 12798 38446 12998
<< pmoslvt >>
rect 17484 27244 18444 27844
rect 18502 27244 19462 27844
rect 19520 27244 20480 27844
rect 20538 27244 21498 27844
rect 21556 27244 22516 27844
rect 22574 27244 23534 27844
rect 23592 27244 24552 27844
rect 24610 27244 25570 27844
rect 25628 27244 26588 27844
rect 26646 27244 27606 27844
rect 27664 27244 28624 27844
rect 28682 27244 29642 27844
rect 29700 27244 30660 27844
rect 30718 27244 31678 27844
rect 31736 27244 32696 27844
rect 32754 27244 33714 27844
rect 17484 26108 18444 26708
rect 18502 26108 19462 26708
rect 19520 26108 20480 26708
rect 20538 26108 21498 26708
rect 21556 26108 22516 26708
rect 22574 26108 23534 26708
rect 23592 26108 24552 26708
rect 24610 26108 25570 26708
rect 25628 26108 26588 26708
rect 26646 26108 27606 26708
rect 27664 26108 28624 26708
rect 28682 26108 29642 26708
rect 29700 26108 30660 26708
rect 30718 26108 31678 26708
rect 31736 26108 32696 26708
rect 32754 26108 33714 26708
rect 17484 24972 18444 25572
rect 18502 24972 19462 25572
rect 19520 24972 20480 25572
rect 20538 24972 21498 25572
rect 21556 24972 22516 25572
rect 22574 24972 23534 25572
rect 23592 24972 24552 25572
rect 24610 24972 25570 25572
rect 25628 24972 26588 25572
rect 26646 24972 27606 25572
rect 27664 24972 28624 25572
rect 28682 24972 29642 25572
rect 29700 24972 30660 25572
rect 30718 24972 31678 25572
rect 31736 24972 32696 25572
rect 32754 24972 33714 25572
rect 18678 23334 19638 23934
rect 19696 23334 20656 23934
rect 20714 23334 21674 23934
rect 21732 23334 22692 23934
rect 22750 23334 23710 23934
rect 23768 23334 24728 23934
rect 24786 23334 25746 23934
rect 25804 23334 26764 23934
rect 26822 23334 27782 23934
rect 27840 23334 28800 23934
rect 28858 23334 29818 23934
rect 29876 23334 30836 23934
rect 30894 23334 31854 23934
rect 31912 23334 32872 23934
rect 18678 22302 19638 22902
rect 19696 22302 20656 22902
rect 20714 22302 21674 22902
rect 21732 22302 22692 22902
rect 22750 22302 23710 22902
rect 23768 22302 24728 22902
rect 24786 22302 25746 22902
rect 25804 22302 26764 22902
rect 26822 22302 27782 22902
rect 27840 22302 28800 22902
rect 28858 22302 29818 22902
rect 29876 22302 30836 22902
rect 30894 22302 31854 22902
rect 31912 22302 32872 22902
rect 13166 20594 14126 21194
rect 14184 20594 15144 21194
rect 15202 20594 16162 21194
rect 16220 20594 17180 21194
rect 13166 19562 14126 20162
rect 14184 19562 15144 20162
rect 15202 19562 16162 20162
rect 16220 19562 17180 20162
rect 13166 18530 14126 19130
rect 14184 18530 15144 19130
rect 15202 18530 16162 19130
rect 16220 18530 17180 19130
rect 13166 17498 14126 18098
rect 14184 17498 15144 18098
rect 15202 17498 16162 18098
rect 16220 17498 17180 18098
rect 58484 27244 59444 27844
rect 59502 27244 60462 27844
rect 60520 27244 61480 27844
rect 61538 27244 62498 27844
rect 62556 27244 63516 27844
rect 63574 27244 64534 27844
rect 64592 27244 65552 27844
rect 65610 27244 66570 27844
rect 66628 27244 67588 27844
rect 67646 27244 68606 27844
rect 68664 27244 69624 27844
rect 69682 27244 70642 27844
rect 70700 27244 71660 27844
rect 71718 27244 72678 27844
rect 72736 27244 73696 27844
rect 73754 27244 74714 27844
rect 58484 26108 59444 26708
rect 59502 26108 60462 26708
rect 60520 26108 61480 26708
rect 61538 26108 62498 26708
rect 62556 26108 63516 26708
rect 63574 26108 64534 26708
rect 64592 26108 65552 26708
rect 65610 26108 66570 26708
rect 66628 26108 67588 26708
rect 67646 26108 68606 26708
rect 68664 26108 69624 26708
rect 69682 26108 70642 26708
rect 70700 26108 71660 26708
rect 71718 26108 72678 26708
rect 72736 26108 73696 26708
rect 73754 26108 74714 26708
rect 58484 24972 59444 25572
rect 59502 24972 60462 25572
rect 60520 24972 61480 25572
rect 61538 24972 62498 25572
rect 62556 24972 63516 25572
rect 63574 24972 64534 25572
rect 64592 24972 65552 25572
rect 65610 24972 66570 25572
rect 66628 24972 67588 25572
rect 67646 24972 68606 25572
rect 68664 24972 69624 25572
rect 69682 24972 70642 25572
rect 70700 24972 71660 25572
rect 71718 24972 72678 25572
rect 72736 24972 73696 25572
rect 73754 24972 74714 25572
rect 59678 23334 60638 23934
rect 60696 23334 61656 23934
rect 61714 23334 62674 23934
rect 62732 23334 63692 23934
rect 63750 23334 64710 23934
rect 64768 23334 65728 23934
rect 65786 23334 66746 23934
rect 66804 23334 67764 23934
rect 67822 23334 68782 23934
rect 68840 23334 69800 23934
rect 69858 23334 70818 23934
rect 70876 23334 71836 23934
rect 71894 23334 72854 23934
rect 72912 23334 73872 23934
rect 59678 22302 60638 22902
rect 60696 22302 61656 22902
rect 61714 22302 62674 22902
rect 62732 22302 63692 22902
rect 63750 22302 64710 22902
rect 64768 22302 65728 22902
rect 65786 22302 66746 22902
rect 66804 22302 67764 22902
rect 67822 22302 68782 22902
rect 68840 22302 69800 22902
rect 69858 22302 70818 22902
rect 70876 22302 71836 22902
rect 71894 22302 72854 22902
rect 72912 22302 73872 22902
rect 54166 20594 55126 21194
rect 55184 20594 56144 21194
rect 56202 20594 57162 21194
rect 57220 20594 58180 21194
rect 54166 19562 55126 20162
rect 55184 19562 56144 20162
rect 56202 19562 57162 20162
rect 57220 19562 58180 20162
rect 54166 18530 55126 19130
rect 55184 18530 56144 19130
rect 56202 18530 57162 19130
rect 57220 18530 58180 19130
rect 54166 17498 55126 18098
rect 55184 17498 56144 18098
rect 56202 17498 57162 18098
rect 57220 17498 58180 18098
<< nmoslvt >>
rect 1812 13258 2772 13858
rect 2830 13258 3790 13858
rect 3848 13258 4808 13858
rect 4866 13258 5826 13858
rect 5884 13258 6844 13858
rect 6902 13258 7862 13858
rect 7920 13258 8880 13858
rect 8938 13258 9898 13858
rect 9956 13258 10916 13858
rect 1812 12440 2772 13040
rect 2830 12440 3790 13040
rect 3848 12440 4808 13040
rect 4866 12440 5826 13040
rect 5884 12440 6844 13040
rect 6902 12440 7862 13040
rect 7920 12440 8880 13040
rect 8938 12440 9898 13040
rect 9956 12440 10916 13040
rect 1812 11622 2772 12222
rect 2830 11622 3790 12222
rect 3848 11622 4808 12222
rect 4866 11622 5826 12222
rect 5884 11622 6844 12222
rect 6902 11622 7862 12222
rect 7920 11622 8880 12222
rect 8938 11622 9898 12222
rect 9956 11622 10916 12222
rect 1812 10804 2772 11404
rect 2830 10804 3790 11404
rect 3848 10804 4808 11404
rect 4866 10804 5826 11404
rect 5884 10804 6844 11404
rect 6902 10804 7862 11404
rect 7920 10804 8880 11404
rect 8938 10804 9898 11404
rect 9956 10804 10916 11404
rect 1812 9986 2772 10586
rect 2830 9986 3790 10586
rect 3848 9986 4808 10586
rect 4866 9986 5826 10586
rect 5884 9986 6844 10586
rect 6902 9986 7862 10586
rect 7920 9986 8880 10586
rect 8938 9986 9898 10586
rect 9956 9986 10916 10586
rect 1812 9168 2772 9768
rect 2830 9168 3790 9768
rect 3848 9168 4808 9768
rect 4866 9168 5826 9768
rect 5884 9168 6844 9768
rect 6902 9168 7862 9768
rect 7920 9168 8880 9768
rect 8938 9168 9898 9768
rect 9956 9168 10916 9768
rect 1812 8350 2772 8950
rect 2830 8350 3790 8950
rect 3848 8350 4808 8950
rect 4866 8350 5826 8950
rect 5884 8350 6844 8950
rect 6902 8350 7862 8950
rect 7920 8350 8880 8950
rect 8938 8350 9898 8950
rect 9956 8350 10916 8950
rect 1812 7532 2772 8132
rect 2830 7532 3790 8132
rect 3848 7532 4808 8132
rect 4866 7532 5826 8132
rect 5884 7532 6844 8132
rect 6902 7532 7862 8132
rect 7920 7532 8880 8132
rect 8938 7532 9898 8132
rect 9956 7532 10916 8132
rect 488 5508 1448 6108
rect 1506 5508 2466 6108
rect 2524 5508 3484 6108
rect 3542 5508 4502 6108
rect 4560 5508 5520 6108
rect 5578 5508 6538 6108
rect 6596 5508 7556 6108
rect 7614 5508 8574 6108
rect 8632 5508 9592 6108
rect 9650 5508 10610 6108
rect 10668 5508 11628 6108
rect 488 4396 1448 4996
rect 1506 4396 2466 4996
rect 2524 4396 3484 4996
rect 3542 4396 4502 4996
rect 4560 4396 5520 4996
rect 5578 4396 6538 4996
rect 6596 4396 7556 4996
rect 7614 4396 8574 4996
rect 8632 4396 9592 4996
rect 9650 4396 10610 4996
rect 10668 4396 11628 4996
rect 488 3284 1448 3884
rect 1506 3284 2466 3884
rect 2524 3284 3484 3884
rect 3542 3284 4502 3884
rect 4560 3284 5520 3884
rect 5578 3284 6538 3884
rect 6596 3284 7556 3884
rect 7614 3284 8574 3884
rect 8632 3284 9592 3884
rect 9650 3284 10610 3884
rect 10668 3284 11628 3884
rect 488 2172 1448 2772
rect 1506 2172 2466 2772
rect 2524 2172 3484 2772
rect 3542 2172 4502 2772
rect 4560 2172 5520 2772
rect 5578 2172 6538 2772
rect 6596 2172 7556 2772
rect 7614 2172 8574 2772
rect 8632 2172 9592 2772
rect 9650 2172 10610 2772
rect 10668 2172 11628 2772
rect 42812 13258 43772 13858
rect 43830 13258 44790 13858
rect 44848 13258 45808 13858
rect 45866 13258 46826 13858
rect 46884 13258 47844 13858
rect 47902 13258 48862 13858
rect 48920 13258 49880 13858
rect 49938 13258 50898 13858
rect 50956 13258 51916 13858
rect 42812 12440 43772 13040
rect 43830 12440 44790 13040
rect 44848 12440 45808 13040
rect 45866 12440 46826 13040
rect 46884 12440 47844 13040
rect 47902 12440 48862 13040
rect 48920 12440 49880 13040
rect 49938 12440 50898 13040
rect 50956 12440 51916 13040
rect 42812 11622 43772 12222
rect 43830 11622 44790 12222
rect 44848 11622 45808 12222
rect 45866 11622 46826 12222
rect 46884 11622 47844 12222
rect 47902 11622 48862 12222
rect 48920 11622 49880 12222
rect 49938 11622 50898 12222
rect 50956 11622 51916 12222
rect 42812 10804 43772 11404
rect 43830 10804 44790 11404
rect 44848 10804 45808 11404
rect 45866 10804 46826 11404
rect 46884 10804 47844 11404
rect 47902 10804 48862 11404
rect 48920 10804 49880 11404
rect 49938 10804 50898 11404
rect 50956 10804 51916 11404
rect 42812 9986 43772 10586
rect 43830 9986 44790 10586
rect 44848 9986 45808 10586
rect 45866 9986 46826 10586
rect 46884 9986 47844 10586
rect 47902 9986 48862 10586
rect 48920 9986 49880 10586
rect 49938 9986 50898 10586
rect 50956 9986 51916 10586
rect 42812 9168 43772 9768
rect 43830 9168 44790 9768
rect 44848 9168 45808 9768
rect 45866 9168 46826 9768
rect 46884 9168 47844 9768
rect 47902 9168 48862 9768
rect 48920 9168 49880 9768
rect 49938 9168 50898 9768
rect 50956 9168 51916 9768
rect 42812 8350 43772 8950
rect 43830 8350 44790 8950
rect 44848 8350 45808 8950
rect 45866 8350 46826 8950
rect 46884 8350 47844 8950
rect 47902 8350 48862 8950
rect 48920 8350 49880 8950
rect 49938 8350 50898 8950
rect 50956 8350 51916 8950
rect 42812 7532 43772 8132
rect 43830 7532 44790 8132
rect 44848 7532 45808 8132
rect 45866 7532 46826 8132
rect 46884 7532 47844 8132
rect 47902 7532 48862 8132
rect 48920 7532 49880 8132
rect 49938 7532 50898 8132
rect 50956 7532 51916 8132
rect 41488 5508 42448 6108
rect 42506 5508 43466 6108
rect 43524 5508 44484 6108
rect 44542 5508 45502 6108
rect 45560 5508 46520 6108
rect 46578 5508 47538 6108
rect 47596 5508 48556 6108
rect 48614 5508 49574 6108
rect 49632 5508 50592 6108
rect 50650 5508 51610 6108
rect 51668 5508 52628 6108
rect 41488 4396 42448 4996
rect 42506 4396 43466 4996
rect 43524 4396 44484 4996
rect 44542 4396 45502 4996
rect 45560 4396 46520 4996
rect 46578 4396 47538 4996
rect 47596 4396 48556 4996
rect 48614 4396 49574 4996
rect 49632 4396 50592 4996
rect 50650 4396 51610 4996
rect 51668 4396 52628 4996
rect 41488 3284 42448 3884
rect 42506 3284 43466 3884
rect 43524 3284 44484 3884
rect 44542 3284 45502 3884
rect 45560 3284 46520 3884
rect 46578 3284 47538 3884
rect 47596 3284 48556 3884
rect 48614 3284 49574 3884
rect 49632 3284 50592 3884
rect 50650 3284 51610 3884
rect 51668 3284 52628 3884
rect 41488 2172 42448 2772
rect 42506 2172 43466 2772
rect 43524 2172 44484 2772
rect 44542 2172 45502 2772
rect 45560 2172 46520 2772
rect 46578 2172 47538 2772
rect 47596 2172 48556 2772
rect 48614 2172 49574 2772
rect 49632 2172 50592 2772
rect 50650 2172 51610 2772
rect 51668 2172 52628 2772
<< ndiff >>
rect 13520 14322 13578 14334
rect 1754 13846 1812 13858
rect 1754 13270 1766 13846
rect 1800 13270 1812 13846
rect 1754 13258 1812 13270
rect 2772 13846 2830 13858
rect 2772 13270 2784 13846
rect 2818 13270 2830 13846
rect 2772 13258 2830 13270
rect 3790 13846 3848 13858
rect 3790 13270 3802 13846
rect 3836 13270 3848 13846
rect 3790 13258 3848 13270
rect 4808 13846 4866 13858
rect 4808 13270 4820 13846
rect 4854 13270 4866 13846
rect 4808 13258 4866 13270
rect 5826 13846 5884 13858
rect 5826 13270 5838 13846
rect 5872 13270 5884 13846
rect 5826 13258 5884 13270
rect 6844 13846 6902 13858
rect 6844 13270 6856 13846
rect 6890 13270 6902 13846
rect 6844 13258 6902 13270
rect 7862 13846 7920 13858
rect 7862 13270 7874 13846
rect 7908 13270 7920 13846
rect 7862 13258 7920 13270
rect 8880 13846 8938 13858
rect 8880 13270 8892 13846
rect 8926 13270 8938 13846
rect 8880 13258 8938 13270
rect 9898 13846 9956 13858
rect 9898 13270 9910 13846
rect 9944 13270 9956 13846
rect 9898 13258 9956 13270
rect 10916 13846 10974 13858
rect 10916 13270 10928 13846
rect 10962 13270 10974 13846
rect 13520 13746 13532 14322
rect 13566 13746 13578 14322
rect 13520 13734 13578 13746
rect 14538 14322 14596 14334
rect 14538 13746 14550 14322
rect 14584 13746 14596 14322
rect 14538 13734 14596 13746
rect 15556 14322 15614 14334
rect 15556 13746 15568 14322
rect 15602 13746 15614 14322
rect 15556 13734 15614 13746
rect 16574 14322 16632 14334
rect 16574 13746 16586 14322
rect 16620 13746 16632 14322
rect 16574 13734 16632 13746
rect 17592 14322 17650 14334
rect 17592 13746 17604 14322
rect 17638 13746 17650 14322
rect 17592 13734 17650 13746
rect 18610 14322 18668 14334
rect 18610 13746 18622 14322
rect 18656 13746 18668 14322
rect 18610 13734 18668 13746
rect 19628 14322 19686 14334
rect 19628 13746 19640 14322
rect 19674 13746 19686 14322
rect 19628 13734 19686 13746
rect 20646 14322 20704 14334
rect 20646 13746 20658 14322
rect 20692 13746 20704 14322
rect 20646 13734 20704 13746
rect 21664 14322 21722 14334
rect 21664 13746 21676 14322
rect 21710 13746 21722 14322
rect 21664 13734 21722 13746
rect 22682 14322 22740 14334
rect 22682 13746 22694 14322
rect 22728 13746 22740 14322
rect 22682 13734 22740 13746
rect 23700 14322 23758 14334
rect 23700 13746 23712 14322
rect 23746 13746 23758 14322
rect 23700 13734 23758 13746
rect 24718 14322 24776 14334
rect 24718 13746 24730 14322
rect 24764 13746 24776 14322
rect 24718 13734 24776 13746
rect 25736 14322 25794 14334
rect 25736 13746 25748 14322
rect 25782 13746 25794 14322
rect 25736 13734 25794 13746
rect 26754 14322 26812 14334
rect 26754 13746 26766 14322
rect 26800 13746 26812 14322
rect 26754 13734 26812 13746
rect 27772 14322 27830 14334
rect 27772 13746 27784 14322
rect 27818 13746 27830 14322
rect 27772 13734 27830 13746
rect 28790 14322 28848 14334
rect 28790 13746 28802 14322
rect 28836 13746 28848 14322
rect 28790 13734 28848 13746
rect 29808 14322 29866 14334
rect 29808 13746 29820 14322
rect 29854 13746 29866 14322
rect 29808 13734 29866 13746
rect 30826 14322 30884 14334
rect 30826 13746 30838 14322
rect 30872 13746 30884 14322
rect 30826 13734 30884 13746
rect 31844 14322 31902 14334
rect 31844 13746 31856 14322
rect 31890 13746 31902 14322
rect 31844 13734 31902 13746
rect 32862 14322 32920 14334
rect 32862 13746 32874 14322
rect 32908 13746 32920 14322
rect 32862 13734 32920 13746
rect 33880 14322 33938 14334
rect 33880 13746 33892 14322
rect 33926 13746 33938 14322
rect 33880 13734 33938 13746
rect 10916 13258 10974 13270
rect 13520 13504 13578 13516
rect 1754 13028 1812 13040
rect 1754 12452 1766 13028
rect 1800 12452 1812 13028
rect 1754 12440 1812 12452
rect 2772 13028 2830 13040
rect 2772 12452 2784 13028
rect 2818 12452 2830 13028
rect 2772 12440 2830 12452
rect 3790 13028 3848 13040
rect 3790 12452 3802 13028
rect 3836 12452 3848 13028
rect 3790 12440 3848 12452
rect 4808 13028 4866 13040
rect 4808 12452 4820 13028
rect 4854 12452 4866 13028
rect 4808 12440 4866 12452
rect 5826 13028 5884 13040
rect 5826 12452 5838 13028
rect 5872 12452 5884 13028
rect 5826 12440 5884 12452
rect 6844 13028 6902 13040
rect 6844 12452 6856 13028
rect 6890 12452 6902 13028
rect 6844 12440 6902 12452
rect 7862 13028 7920 13040
rect 7862 12452 7874 13028
rect 7908 12452 7920 13028
rect 7862 12440 7920 12452
rect 8880 13028 8938 13040
rect 8880 12452 8892 13028
rect 8926 12452 8938 13028
rect 8880 12440 8938 12452
rect 9898 13028 9956 13040
rect 9898 12452 9910 13028
rect 9944 12452 9956 13028
rect 9898 12440 9956 12452
rect 10916 13028 10974 13040
rect 10916 12452 10928 13028
rect 10962 12452 10974 13028
rect 13520 12928 13532 13504
rect 13566 12928 13578 13504
rect 13520 12916 13578 12928
rect 14538 13504 14596 13516
rect 14538 12928 14550 13504
rect 14584 12928 14596 13504
rect 14538 12916 14596 12928
rect 15556 13504 15614 13516
rect 15556 12928 15568 13504
rect 15602 12928 15614 13504
rect 15556 12916 15614 12928
rect 16574 13504 16632 13516
rect 16574 12928 16586 13504
rect 16620 12928 16632 13504
rect 16574 12916 16632 12928
rect 17592 13504 17650 13516
rect 17592 12928 17604 13504
rect 17638 12928 17650 13504
rect 17592 12916 17650 12928
rect 18610 13504 18668 13516
rect 18610 12928 18622 13504
rect 18656 12928 18668 13504
rect 18610 12916 18668 12928
rect 19628 13504 19686 13516
rect 19628 12928 19640 13504
rect 19674 12928 19686 13504
rect 19628 12916 19686 12928
rect 20646 13504 20704 13516
rect 20646 12928 20658 13504
rect 20692 12928 20704 13504
rect 20646 12916 20704 12928
rect 21664 13504 21722 13516
rect 21664 12928 21676 13504
rect 21710 12928 21722 13504
rect 21664 12916 21722 12928
rect 22682 13504 22740 13516
rect 22682 12928 22694 13504
rect 22728 12928 22740 13504
rect 22682 12916 22740 12928
rect 23700 13504 23758 13516
rect 23700 12928 23712 13504
rect 23746 12928 23758 13504
rect 23700 12916 23758 12928
rect 24718 13504 24776 13516
rect 24718 12928 24730 13504
rect 24764 12928 24776 13504
rect 24718 12916 24776 12928
rect 25736 13504 25794 13516
rect 25736 12928 25748 13504
rect 25782 12928 25794 13504
rect 25736 12916 25794 12928
rect 26754 13504 26812 13516
rect 26754 12928 26766 13504
rect 26800 12928 26812 13504
rect 26754 12916 26812 12928
rect 27772 13504 27830 13516
rect 27772 12928 27784 13504
rect 27818 12928 27830 13504
rect 27772 12916 27830 12928
rect 28790 13504 28848 13516
rect 28790 12928 28802 13504
rect 28836 12928 28848 13504
rect 28790 12916 28848 12928
rect 29808 13504 29866 13516
rect 29808 12928 29820 13504
rect 29854 12928 29866 13504
rect 29808 12916 29866 12928
rect 30826 13504 30884 13516
rect 30826 12928 30838 13504
rect 30872 12928 30884 13504
rect 30826 12916 30884 12928
rect 31844 13504 31902 13516
rect 31844 12928 31856 13504
rect 31890 12928 31902 13504
rect 31844 12916 31902 12928
rect 32862 13504 32920 13516
rect 32862 12928 32874 13504
rect 32908 12928 32920 13504
rect 32862 12916 32920 12928
rect 33880 13504 33938 13516
rect 33880 12928 33892 13504
rect 33926 12928 33938 13504
rect 33880 12916 33938 12928
rect 10916 12440 10974 12452
rect 1754 12210 1812 12222
rect 1754 11634 1766 12210
rect 1800 11634 1812 12210
rect 1754 11622 1812 11634
rect 2772 12210 2830 12222
rect 2772 11634 2784 12210
rect 2818 11634 2830 12210
rect 2772 11622 2830 11634
rect 3790 12210 3848 12222
rect 3790 11634 3802 12210
rect 3836 11634 3848 12210
rect 3790 11622 3848 11634
rect 4808 12210 4866 12222
rect 4808 11634 4820 12210
rect 4854 11634 4866 12210
rect 4808 11622 4866 11634
rect 5826 12210 5884 12222
rect 5826 11634 5838 12210
rect 5872 11634 5884 12210
rect 5826 11622 5884 11634
rect 6844 12210 6902 12222
rect 6844 11634 6856 12210
rect 6890 11634 6902 12210
rect 6844 11622 6902 11634
rect 7862 12210 7920 12222
rect 7862 11634 7874 12210
rect 7908 11634 7920 12210
rect 7862 11622 7920 11634
rect 8880 12210 8938 12222
rect 8880 11634 8892 12210
rect 8926 11634 8938 12210
rect 8880 11622 8938 11634
rect 9898 12210 9956 12222
rect 9898 11634 9910 12210
rect 9944 11634 9956 12210
rect 9898 11622 9956 11634
rect 10916 12210 10974 12222
rect 10916 11634 10928 12210
rect 10962 11634 10974 12210
rect 10916 11622 10974 11634
rect 13520 12126 13578 12138
rect 13520 11550 13532 12126
rect 13566 11550 13578 12126
rect 13520 11538 13578 11550
rect 14538 12126 14596 12138
rect 14538 11550 14550 12126
rect 14584 11550 14596 12126
rect 14538 11538 14596 11550
rect 15556 12126 15614 12138
rect 15556 11550 15568 12126
rect 15602 11550 15614 12126
rect 15556 11538 15614 11550
rect 16574 12126 16632 12138
rect 16574 11550 16586 12126
rect 16620 11550 16632 12126
rect 16574 11538 16632 11550
rect 17592 12126 17650 12138
rect 17592 11550 17604 12126
rect 17638 11550 17650 12126
rect 17592 11538 17650 11550
rect 18610 12126 18668 12138
rect 18610 11550 18622 12126
rect 18656 11550 18668 12126
rect 18610 11538 18668 11550
rect 19628 12126 19686 12138
rect 19628 11550 19640 12126
rect 19674 11550 19686 12126
rect 19628 11538 19686 11550
rect 20646 12126 20704 12138
rect 20646 11550 20658 12126
rect 20692 11550 20704 12126
rect 20646 11538 20704 11550
rect 21664 12126 21722 12138
rect 21664 11550 21676 12126
rect 21710 11550 21722 12126
rect 21664 11538 21722 11550
rect 22682 12126 22740 12138
rect 22682 11550 22694 12126
rect 22728 11550 22740 12126
rect 22682 11538 22740 11550
rect 23700 12126 23758 12138
rect 23700 11550 23712 12126
rect 23746 11550 23758 12126
rect 23700 11538 23758 11550
rect 24718 12126 24776 12138
rect 24718 11550 24730 12126
rect 24764 11550 24776 12126
rect 24718 11538 24776 11550
rect 25736 12126 25794 12138
rect 25736 11550 25748 12126
rect 25782 11550 25794 12126
rect 25736 11538 25794 11550
rect 26754 12126 26812 12138
rect 26754 11550 26766 12126
rect 26800 11550 26812 12126
rect 26754 11538 26812 11550
rect 27772 12126 27830 12138
rect 27772 11550 27784 12126
rect 27818 11550 27830 12126
rect 27772 11538 27830 11550
rect 28790 12126 28848 12138
rect 28790 11550 28802 12126
rect 28836 11550 28848 12126
rect 28790 11538 28848 11550
rect 29808 12126 29866 12138
rect 29808 11550 29820 12126
rect 29854 11550 29866 12126
rect 29808 11538 29866 11550
rect 30826 12126 30884 12138
rect 30826 11550 30838 12126
rect 30872 11550 30884 12126
rect 30826 11538 30884 11550
rect 31844 12126 31902 12138
rect 31844 11550 31856 12126
rect 31890 11550 31902 12126
rect 31844 11538 31902 11550
rect 32862 12126 32920 12138
rect 32862 11550 32874 12126
rect 32908 11550 32920 12126
rect 32862 11538 32920 11550
rect 33880 12126 33938 12138
rect 33880 11550 33892 12126
rect 33926 11550 33938 12126
rect 33880 11538 33938 11550
rect 1754 11392 1812 11404
rect 1754 10816 1766 11392
rect 1800 10816 1812 11392
rect 1754 10804 1812 10816
rect 2772 11392 2830 11404
rect 2772 10816 2784 11392
rect 2818 10816 2830 11392
rect 2772 10804 2830 10816
rect 3790 11392 3848 11404
rect 3790 10816 3802 11392
rect 3836 10816 3848 11392
rect 3790 10804 3848 10816
rect 4808 11392 4866 11404
rect 4808 10816 4820 11392
rect 4854 10816 4866 11392
rect 4808 10804 4866 10816
rect 5826 11392 5884 11404
rect 5826 10816 5838 11392
rect 5872 10816 5884 11392
rect 5826 10804 5884 10816
rect 6844 11392 6902 11404
rect 6844 10816 6856 11392
rect 6890 10816 6902 11392
rect 6844 10804 6902 10816
rect 7862 11392 7920 11404
rect 7862 10816 7874 11392
rect 7908 10816 7920 11392
rect 7862 10804 7920 10816
rect 8880 11392 8938 11404
rect 8880 10816 8892 11392
rect 8926 10816 8938 11392
rect 8880 10804 8938 10816
rect 9898 11392 9956 11404
rect 9898 10816 9910 11392
rect 9944 10816 9956 11392
rect 9898 10804 9956 10816
rect 10916 11392 10974 11404
rect 10916 10816 10928 11392
rect 10962 10816 10974 11392
rect 10916 10804 10974 10816
rect 13520 10894 13578 10906
rect 1754 10574 1812 10586
rect 1754 9998 1766 10574
rect 1800 9998 1812 10574
rect 1754 9986 1812 9998
rect 2772 10574 2830 10586
rect 2772 9998 2784 10574
rect 2818 9998 2830 10574
rect 2772 9986 2830 9998
rect 3790 10574 3848 10586
rect 3790 9998 3802 10574
rect 3836 9998 3848 10574
rect 3790 9986 3848 9998
rect 4808 10574 4866 10586
rect 4808 9998 4820 10574
rect 4854 9998 4866 10574
rect 4808 9986 4866 9998
rect 5826 10574 5884 10586
rect 5826 9998 5838 10574
rect 5872 9998 5884 10574
rect 5826 9986 5884 9998
rect 6844 10574 6902 10586
rect 6844 9998 6856 10574
rect 6890 9998 6902 10574
rect 6844 9986 6902 9998
rect 7862 10574 7920 10586
rect 7862 9998 7874 10574
rect 7908 9998 7920 10574
rect 7862 9986 7920 9998
rect 8880 10574 8938 10586
rect 8880 9998 8892 10574
rect 8926 9998 8938 10574
rect 8880 9986 8938 9998
rect 9898 10574 9956 10586
rect 9898 9998 9910 10574
rect 9944 9998 9956 10574
rect 9898 9986 9956 9998
rect 10916 10574 10974 10586
rect 10916 9998 10928 10574
rect 10962 9998 10974 10574
rect 13520 10318 13532 10894
rect 13566 10318 13578 10894
rect 13520 10306 13578 10318
rect 14538 10894 14596 10906
rect 14538 10318 14550 10894
rect 14584 10318 14596 10894
rect 14538 10306 14596 10318
rect 15556 10894 15614 10906
rect 15556 10318 15568 10894
rect 15602 10318 15614 10894
rect 15556 10306 15614 10318
rect 16574 10894 16632 10906
rect 16574 10318 16586 10894
rect 16620 10318 16632 10894
rect 16574 10306 16632 10318
rect 17592 10894 17650 10906
rect 17592 10318 17604 10894
rect 17638 10318 17650 10894
rect 17592 10306 17650 10318
rect 18610 10894 18668 10906
rect 18610 10318 18622 10894
rect 18656 10318 18668 10894
rect 18610 10306 18668 10318
rect 19628 10894 19686 10906
rect 19628 10318 19640 10894
rect 19674 10318 19686 10894
rect 19628 10306 19686 10318
rect 20646 10894 20704 10906
rect 20646 10318 20658 10894
rect 20692 10318 20704 10894
rect 20646 10306 20704 10318
rect 21664 10894 21722 10906
rect 21664 10318 21676 10894
rect 21710 10318 21722 10894
rect 21664 10306 21722 10318
rect 22682 10894 22740 10906
rect 22682 10318 22694 10894
rect 22728 10318 22740 10894
rect 22682 10306 22740 10318
rect 23700 10894 23758 10906
rect 23700 10318 23712 10894
rect 23746 10318 23758 10894
rect 23700 10306 23758 10318
rect 24718 10894 24776 10906
rect 24718 10318 24730 10894
rect 24764 10318 24776 10894
rect 24718 10306 24776 10318
rect 25736 10894 25794 10906
rect 25736 10318 25748 10894
rect 25782 10318 25794 10894
rect 25736 10306 25794 10318
rect 26754 10894 26812 10906
rect 26754 10318 26766 10894
rect 26800 10318 26812 10894
rect 26754 10306 26812 10318
rect 27772 10894 27830 10906
rect 27772 10318 27784 10894
rect 27818 10318 27830 10894
rect 27772 10306 27830 10318
rect 28790 10894 28848 10906
rect 28790 10318 28802 10894
rect 28836 10318 28848 10894
rect 28790 10306 28848 10318
rect 29808 10894 29866 10906
rect 29808 10318 29820 10894
rect 29854 10318 29866 10894
rect 29808 10306 29866 10318
rect 30826 10894 30884 10906
rect 30826 10318 30838 10894
rect 30872 10318 30884 10894
rect 30826 10306 30884 10318
rect 31844 10894 31902 10906
rect 31844 10318 31856 10894
rect 31890 10318 31902 10894
rect 31844 10306 31902 10318
rect 32862 10894 32920 10906
rect 32862 10318 32874 10894
rect 32908 10318 32920 10894
rect 32862 10306 32920 10318
rect 33880 10894 33938 10906
rect 33880 10318 33892 10894
rect 33926 10318 33938 10894
rect 33880 10306 33938 10318
rect 10916 9986 10974 9998
rect 1754 9756 1812 9768
rect 1754 9180 1766 9756
rect 1800 9180 1812 9756
rect 1754 9168 1812 9180
rect 2772 9756 2830 9768
rect 2772 9180 2784 9756
rect 2818 9180 2830 9756
rect 2772 9168 2830 9180
rect 3790 9756 3848 9768
rect 3790 9180 3802 9756
rect 3836 9180 3848 9756
rect 3790 9168 3848 9180
rect 4808 9756 4866 9768
rect 4808 9180 4820 9756
rect 4854 9180 4866 9756
rect 4808 9168 4866 9180
rect 5826 9756 5884 9768
rect 5826 9180 5838 9756
rect 5872 9180 5884 9756
rect 5826 9168 5884 9180
rect 6844 9756 6902 9768
rect 6844 9180 6856 9756
rect 6890 9180 6902 9756
rect 6844 9168 6902 9180
rect 7862 9756 7920 9768
rect 7862 9180 7874 9756
rect 7908 9180 7920 9756
rect 7862 9168 7920 9180
rect 8880 9756 8938 9768
rect 8880 9180 8892 9756
rect 8926 9180 8938 9756
rect 8880 9168 8938 9180
rect 9898 9756 9956 9768
rect 9898 9180 9910 9756
rect 9944 9180 9956 9756
rect 9898 9168 9956 9180
rect 10916 9756 10974 9768
rect 10916 9180 10928 9756
rect 10962 9180 10974 9756
rect 10916 9168 10974 9180
rect 13518 9660 13576 9672
rect 13518 9084 13530 9660
rect 13564 9084 13576 9660
rect 13518 9072 13576 9084
rect 14536 9660 14594 9672
rect 14536 9084 14548 9660
rect 14582 9084 14594 9660
rect 14536 9072 14594 9084
rect 15554 9660 15612 9672
rect 15554 9084 15566 9660
rect 15600 9084 15612 9660
rect 15554 9072 15612 9084
rect 16572 9660 16630 9672
rect 16572 9084 16584 9660
rect 16618 9084 16630 9660
rect 16572 9072 16630 9084
rect 17590 9660 17648 9672
rect 17590 9084 17602 9660
rect 17636 9084 17648 9660
rect 17590 9072 17648 9084
rect 18608 9660 18666 9672
rect 18608 9084 18620 9660
rect 18654 9084 18666 9660
rect 18608 9072 18666 9084
rect 19626 9660 19684 9672
rect 19626 9084 19638 9660
rect 19672 9084 19684 9660
rect 19626 9072 19684 9084
rect 20644 9660 20702 9672
rect 20644 9084 20656 9660
rect 20690 9084 20702 9660
rect 20644 9072 20702 9084
rect 21662 9660 21720 9672
rect 21662 9084 21674 9660
rect 21708 9084 21720 9660
rect 21662 9072 21720 9084
rect 22680 9660 22738 9672
rect 22680 9084 22692 9660
rect 22726 9084 22738 9660
rect 22680 9072 22738 9084
rect 23698 9660 23756 9672
rect 23698 9084 23710 9660
rect 23744 9084 23756 9660
rect 23698 9072 23756 9084
rect 24716 9660 24774 9672
rect 24716 9084 24728 9660
rect 24762 9084 24774 9660
rect 24716 9072 24774 9084
rect 25734 9660 25792 9672
rect 25734 9084 25746 9660
rect 25780 9084 25792 9660
rect 25734 9072 25792 9084
rect 26752 9660 26810 9672
rect 26752 9084 26764 9660
rect 26798 9084 26810 9660
rect 26752 9072 26810 9084
rect 27770 9660 27828 9672
rect 27770 9084 27782 9660
rect 27816 9084 27828 9660
rect 27770 9072 27828 9084
rect 28788 9660 28846 9672
rect 28788 9084 28800 9660
rect 28834 9084 28846 9660
rect 28788 9072 28846 9084
rect 29806 9660 29864 9672
rect 29806 9084 29818 9660
rect 29852 9084 29864 9660
rect 29806 9072 29864 9084
rect 30824 9660 30882 9672
rect 30824 9084 30836 9660
rect 30870 9084 30882 9660
rect 30824 9072 30882 9084
rect 31842 9660 31900 9672
rect 31842 9084 31854 9660
rect 31888 9084 31900 9660
rect 31842 9072 31900 9084
rect 32860 9660 32918 9672
rect 32860 9084 32872 9660
rect 32906 9084 32918 9660
rect 32860 9072 32918 9084
rect 33878 9660 33936 9672
rect 33878 9084 33890 9660
rect 33924 9084 33936 9660
rect 33878 9072 33936 9084
rect 1754 8938 1812 8950
rect 1754 8362 1766 8938
rect 1800 8362 1812 8938
rect 1754 8350 1812 8362
rect 2772 8938 2830 8950
rect 2772 8362 2784 8938
rect 2818 8362 2830 8938
rect 2772 8350 2830 8362
rect 3790 8938 3848 8950
rect 3790 8362 3802 8938
rect 3836 8362 3848 8938
rect 3790 8350 3848 8362
rect 4808 8938 4866 8950
rect 4808 8362 4820 8938
rect 4854 8362 4866 8938
rect 4808 8350 4866 8362
rect 5826 8938 5884 8950
rect 5826 8362 5838 8938
rect 5872 8362 5884 8938
rect 5826 8350 5884 8362
rect 6844 8938 6902 8950
rect 6844 8362 6856 8938
rect 6890 8362 6902 8938
rect 6844 8350 6902 8362
rect 7862 8938 7920 8950
rect 7862 8362 7874 8938
rect 7908 8362 7920 8938
rect 7862 8350 7920 8362
rect 8880 8938 8938 8950
rect 8880 8362 8892 8938
rect 8926 8362 8938 8938
rect 8880 8350 8938 8362
rect 9898 8938 9956 8950
rect 9898 8362 9910 8938
rect 9944 8362 9956 8938
rect 9898 8350 9956 8362
rect 10916 8938 10974 8950
rect 10916 8362 10928 8938
rect 10962 8362 10974 8938
rect 10916 8350 10974 8362
rect 13518 8426 13576 8438
rect 1754 8120 1812 8132
rect 1754 7544 1766 8120
rect 1800 7544 1812 8120
rect 1754 7532 1812 7544
rect 2772 8120 2830 8132
rect 2772 7544 2784 8120
rect 2818 7544 2830 8120
rect 2772 7532 2830 7544
rect 3790 8120 3848 8132
rect 3790 7544 3802 8120
rect 3836 7544 3848 8120
rect 3790 7532 3848 7544
rect 4808 8120 4866 8132
rect 4808 7544 4820 8120
rect 4854 7544 4866 8120
rect 4808 7532 4866 7544
rect 5826 8120 5884 8132
rect 5826 7544 5838 8120
rect 5872 7544 5884 8120
rect 5826 7532 5884 7544
rect 6844 8120 6902 8132
rect 6844 7544 6856 8120
rect 6890 7544 6902 8120
rect 6844 7532 6902 7544
rect 7862 8120 7920 8132
rect 7862 7544 7874 8120
rect 7908 7544 7920 8120
rect 7862 7532 7920 7544
rect 8880 8120 8938 8132
rect 8880 7544 8892 8120
rect 8926 7544 8938 8120
rect 8880 7532 8938 7544
rect 9898 8120 9956 8132
rect 9898 7544 9910 8120
rect 9944 7544 9956 8120
rect 9898 7532 9956 7544
rect 10916 8120 10974 8132
rect 10916 7544 10928 8120
rect 10962 7544 10974 8120
rect 13518 7850 13530 8426
rect 13564 7850 13576 8426
rect 13518 7838 13576 7850
rect 14536 8426 14594 8438
rect 14536 7850 14548 8426
rect 14582 7850 14594 8426
rect 14536 7838 14594 7850
rect 15554 8426 15612 8438
rect 15554 7850 15566 8426
rect 15600 7850 15612 8426
rect 15554 7838 15612 7850
rect 16572 8426 16630 8438
rect 16572 7850 16584 8426
rect 16618 7850 16630 8426
rect 16572 7838 16630 7850
rect 17590 8426 17648 8438
rect 17590 7850 17602 8426
rect 17636 7850 17648 8426
rect 17590 7838 17648 7850
rect 18608 8426 18666 8438
rect 18608 7850 18620 8426
rect 18654 7850 18666 8426
rect 18608 7838 18666 7850
rect 19626 8426 19684 8438
rect 19626 7850 19638 8426
rect 19672 7850 19684 8426
rect 19626 7838 19684 7850
rect 20644 8426 20702 8438
rect 20644 7850 20656 8426
rect 20690 7850 20702 8426
rect 20644 7838 20702 7850
rect 21662 8426 21720 8438
rect 21662 7850 21674 8426
rect 21708 7850 21720 8426
rect 21662 7838 21720 7850
rect 22680 8426 22738 8438
rect 22680 7850 22692 8426
rect 22726 7850 22738 8426
rect 22680 7838 22738 7850
rect 23698 8426 23756 8438
rect 23698 7850 23710 8426
rect 23744 7850 23756 8426
rect 23698 7838 23756 7850
rect 24716 8426 24774 8438
rect 24716 7850 24728 8426
rect 24762 7850 24774 8426
rect 24716 7838 24774 7850
rect 25734 8426 25792 8438
rect 25734 7850 25746 8426
rect 25780 7850 25792 8426
rect 25734 7838 25792 7850
rect 26752 8426 26810 8438
rect 26752 7850 26764 8426
rect 26798 7850 26810 8426
rect 26752 7838 26810 7850
rect 27770 8426 27828 8438
rect 27770 7850 27782 8426
rect 27816 7850 27828 8426
rect 27770 7838 27828 7850
rect 28788 8426 28846 8438
rect 28788 7850 28800 8426
rect 28834 7850 28846 8426
rect 28788 7838 28846 7850
rect 29806 8426 29864 8438
rect 29806 7850 29818 8426
rect 29852 7850 29864 8426
rect 29806 7838 29864 7850
rect 30824 8426 30882 8438
rect 30824 7850 30836 8426
rect 30870 7850 30882 8426
rect 30824 7838 30882 7850
rect 31842 8426 31900 8438
rect 31842 7850 31854 8426
rect 31888 7850 31900 8426
rect 31842 7838 31900 7850
rect 32860 8426 32918 8438
rect 32860 7850 32872 8426
rect 32906 7850 32918 8426
rect 32860 7838 32918 7850
rect 33878 8426 33936 8438
rect 33878 7850 33890 8426
rect 33924 7850 33936 8426
rect 33878 7838 33936 7850
rect 10916 7532 10974 7544
rect 13518 7194 13576 7206
rect 13518 6618 13530 7194
rect 13564 6618 13576 7194
rect 13518 6606 13576 6618
rect 14536 7194 14594 7206
rect 14536 6618 14548 7194
rect 14582 6618 14594 7194
rect 14536 6606 14594 6618
rect 15554 7194 15612 7206
rect 15554 6618 15566 7194
rect 15600 6618 15612 7194
rect 15554 6606 15612 6618
rect 16572 7194 16630 7206
rect 16572 6618 16584 7194
rect 16618 6618 16630 7194
rect 16572 6606 16630 6618
rect 17590 7194 17648 7206
rect 17590 6618 17602 7194
rect 17636 6618 17648 7194
rect 17590 6606 17648 6618
rect 18608 7194 18666 7206
rect 18608 6618 18620 7194
rect 18654 6618 18666 7194
rect 18608 6606 18666 6618
rect 19626 7194 19684 7206
rect 19626 6618 19638 7194
rect 19672 6618 19684 7194
rect 19626 6606 19684 6618
rect 20644 7194 20702 7206
rect 20644 6618 20656 7194
rect 20690 6618 20702 7194
rect 20644 6606 20702 6618
rect 21662 7194 21720 7206
rect 21662 6618 21674 7194
rect 21708 6618 21720 7194
rect 21662 6606 21720 6618
rect 22680 7194 22738 7206
rect 22680 6618 22692 7194
rect 22726 6618 22738 7194
rect 22680 6606 22738 6618
rect 23698 7194 23756 7206
rect 23698 6618 23710 7194
rect 23744 6618 23756 7194
rect 23698 6606 23756 6618
rect 24716 7194 24774 7206
rect 24716 6618 24728 7194
rect 24762 6618 24774 7194
rect 24716 6606 24774 6618
rect 25734 7194 25792 7206
rect 25734 6618 25746 7194
rect 25780 6618 25792 7194
rect 25734 6606 25792 6618
rect 26752 7194 26810 7206
rect 26752 6618 26764 7194
rect 26798 6618 26810 7194
rect 26752 6606 26810 6618
rect 27770 7194 27828 7206
rect 27770 6618 27782 7194
rect 27816 6618 27828 7194
rect 27770 6606 27828 6618
rect 28788 7194 28846 7206
rect 28788 6618 28800 7194
rect 28834 6618 28846 7194
rect 28788 6606 28846 6618
rect 29806 7194 29864 7206
rect 29806 6618 29818 7194
rect 29852 6618 29864 7194
rect 29806 6606 29864 6618
rect 30824 7194 30882 7206
rect 30824 6618 30836 7194
rect 30870 6618 30882 7194
rect 30824 6606 30882 6618
rect 31842 7194 31900 7206
rect 31842 6618 31854 7194
rect 31888 6618 31900 7194
rect 31842 6606 31900 6618
rect 32860 7194 32918 7206
rect 32860 6618 32872 7194
rect 32906 6618 32918 7194
rect 32860 6606 32918 6618
rect 33878 7194 33936 7206
rect 33878 6618 33890 7194
rect 33924 6618 33936 7194
rect 33878 6606 33936 6618
rect 430 6096 488 6108
rect 430 5520 442 6096
rect 476 5520 488 6096
rect 430 5508 488 5520
rect 1448 6096 1506 6108
rect 1448 5520 1460 6096
rect 1494 5520 1506 6096
rect 1448 5508 1506 5520
rect 2466 6096 2524 6108
rect 2466 5520 2478 6096
rect 2512 5520 2524 6096
rect 2466 5508 2524 5520
rect 3484 6096 3542 6108
rect 3484 5520 3496 6096
rect 3530 5520 3542 6096
rect 3484 5508 3542 5520
rect 4502 6096 4560 6108
rect 4502 5520 4514 6096
rect 4548 5520 4560 6096
rect 4502 5508 4560 5520
rect 5520 6096 5578 6108
rect 5520 5520 5532 6096
rect 5566 5520 5578 6096
rect 5520 5508 5578 5520
rect 6538 6096 6596 6108
rect 6538 5520 6550 6096
rect 6584 5520 6596 6096
rect 6538 5508 6596 5520
rect 7556 6096 7614 6108
rect 7556 5520 7568 6096
rect 7602 5520 7614 6096
rect 7556 5508 7614 5520
rect 8574 6096 8632 6108
rect 8574 5520 8586 6096
rect 8620 5520 8632 6096
rect 8574 5508 8632 5520
rect 9592 6096 9650 6108
rect 9592 5520 9604 6096
rect 9638 5520 9650 6096
rect 9592 5508 9650 5520
rect 10610 6096 10668 6108
rect 10610 5520 10622 6096
rect 10656 5520 10668 6096
rect 10610 5508 10668 5520
rect 11628 6096 11686 6108
rect 11628 5520 11640 6096
rect 11674 5520 11686 6096
rect 11628 5508 11686 5520
rect 13518 5960 13576 5972
rect 13518 5384 13530 5960
rect 13564 5384 13576 5960
rect 13518 5372 13576 5384
rect 14536 5960 14594 5972
rect 14536 5384 14548 5960
rect 14582 5384 14594 5960
rect 14536 5372 14594 5384
rect 15554 5960 15612 5972
rect 15554 5384 15566 5960
rect 15600 5384 15612 5960
rect 15554 5372 15612 5384
rect 16572 5960 16630 5972
rect 16572 5384 16584 5960
rect 16618 5384 16630 5960
rect 16572 5372 16630 5384
rect 17590 5960 17648 5972
rect 17590 5384 17602 5960
rect 17636 5384 17648 5960
rect 17590 5372 17648 5384
rect 18608 5960 18666 5972
rect 18608 5384 18620 5960
rect 18654 5384 18666 5960
rect 18608 5372 18666 5384
rect 19626 5960 19684 5972
rect 19626 5384 19638 5960
rect 19672 5384 19684 5960
rect 19626 5372 19684 5384
rect 20644 5960 20702 5972
rect 20644 5384 20656 5960
rect 20690 5384 20702 5960
rect 20644 5372 20702 5384
rect 21662 5960 21720 5972
rect 21662 5384 21674 5960
rect 21708 5384 21720 5960
rect 21662 5372 21720 5384
rect 22680 5960 22738 5972
rect 22680 5384 22692 5960
rect 22726 5384 22738 5960
rect 22680 5372 22738 5384
rect 23698 5960 23756 5972
rect 23698 5384 23710 5960
rect 23744 5384 23756 5960
rect 23698 5372 23756 5384
rect 24716 5960 24774 5972
rect 24716 5384 24728 5960
rect 24762 5384 24774 5960
rect 24716 5372 24774 5384
rect 25734 5960 25792 5972
rect 25734 5384 25746 5960
rect 25780 5384 25792 5960
rect 25734 5372 25792 5384
rect 26752 5960 26810 5972
rect 26752 5384 26764 5960
rect 26798 5384 26810 5960
rect 26752 5372 26810 5384
rect 27770 5960 27828 5972
rect 27770 5384 27782 5960
rect 27816 5384 27828 5960
rect 27770 5372 27828 5384
rect 28788 5960 28846 5972
rect 28788 5384 28800 5960
rect 28834 5384 28846 5960
rect 28788 5372 28846 5384
rect 29806 5960 29864 5972
rect 29806 5384 29818 5960
rect 29852 5384 29864 5960
rect 29806 5372 29864 5384
rect 30824 5960 30882 5972
rect 30824 5384 30836 5960
rect 30870 5384 30882 5960
rect 30824 5372 30882 5384
rect 31842 5960 31900 5972
rect 31842 5384 31854 5960
rect 31888 5384 31900 5960
rect 31842 5372 31900 5384
rect 32860 5960 32918 5972
rect 32860 5384 32872 5960
rect 32906 5384 32918 5960
rect 32860 5372 32918 5384
rect 33878 5960 33936 5972
rect 33878 5384 33890 5960
rect 33924 5384 33936 5960
rect 33878 5372 33936 5384
rect 430 4984 488 4996
rect 430 4408 442 4984
rect 476 4408 488 4984
rect 430 4396 488 4408
rect 1448 4984 1506 4996
rect 1448 4408 1460 4984
rect 1494 4408 1506 4984
rect 1448 4396 1506 4408
rect 2466 4984 2524 4996
rect 2466 4408 2478 4984
rect 2512 4408 2524 4984
rect 2466 4396 2524 4408
rect 3484 4984 3542 4996
rect 3484 4408 3496 4984
rect 3530 4408 3542 4984
rect 3484 4396 3542 4408
rect 4502 4984 4560 4996
rect 4502 4408 4514 4984
rect 4548 4408 4560 4984
rect 4502 4396 4560 4408
rect 5520 4984 5578 4996
rect 5520 4408 5532 4984
rect 5566 4408 5578 4984
rect 5520 4396 5578 4408
rect 6538 4984 6596 4996
rect 6538 4408 6550 4984
rect 6584 4408 6596 4984
rect 6538 4396 6596 4408
rect 7556 4984 7614 4996
rect 7556 4408 7568 4984
rect 7602 4408 7614 4984
rect 7556 4396 7614 4408
rect 8574 4984 8632 4996
rect 8574 4408 8586 4984
rect 8620 4408 8632 4984
rect 8574 4396 8632 4408
rect 9592 4984 9650 4996
rect 9592 4408 9604 4984
rect 9638 4408 9650 4984
rect 9592 4396 9650 4408
rect 10610 4984 10668 4996
rect 10610 4408 10622 4984
rect 10656 4408 10668 4984
rect 10610 4396 10668 4408
rect 11628 4984 11686 4996
rect 11628 4408 11640 4984
rect 11674 4408 11686 4984
rect 11628 4396 11686 4408
rect 13518 4726 13576 4738
rect 13518 4150 13530 4726
rect 13564 4150 13576 4726
rect 13518 4138 13576 4150
rect 14536 4726 14594 4738
rect 14536 4150 14548 4726
rect 14582 4150 14594 4726
rect 14536 4138 14594 4150
rect 15554 4726 15612 4738
rect 15554 4150 15566 4726
rect 15600 4150 15612 4726
rect 15554 4138 15612 4150
rect 16572 4726 16630 4738
rect 16572 4150 16584 4726
rect 16618 4150 16630 4726
rect 16572 4138 16630 4150
rect 17590 4726 17648 4738
rect 17590 4150 17602 4726
rect 17636 4150 17648 4726
rect 17590 4138 17648 4150
rect 18608 4726 18666 4738
rect 18608 4150 18620 4726
rect 18654 4150 18666 4726
rect 18608 4138 18666 4150
rect 19626 4726 19684 4738
rect 19626 4150 19638 4726
rect 19672 4150 19684 4726
rect 19626 4138 19684 4150
rect 20644 4726 20702 4738
rect 20644 4150 20656 4726
rect 20690 4150 20702 4726
rect 20644 4138 20702 4150
rect 21662 4726 21720 4738
rect 21662 4150 21674 4726
rect 21708 4150 21720 4726
rect 21662 4138 21720 4150
rect 22680 4726 22738 4738
rect 22680 4150 22692 4726
rect 22726 4150 22738 4726
rect 22680 4138 22738 4150
rect 23698 4726 23756 4738
rect 23698 4150 23710 4726
rect 23744 4150 23756 4726
rect 23698 4138 23756 4150
rect 24716 4726 24774 4738
rect 24716 4150 24728 4726
rect 24762 4150 24774 4726
rect 24716 4138 24774 4150
rect 25734 4726 25792 4738
rect 25734 4150 25746 4726
rect 25780 4150 25792 4726
rect 25734 4138 25792 4150
rect 26752 4726 26810 4738
rect 26752 4150 26764 4726
rect 26798 4150 26810 4726
rect 26752 4138 26810 4150
rect 27770 4726 27828 4738
rect 27770 4150 27782 4726
rect 27816 4150 27828 4726
rect 27770 4138 27828 4150
rect 28788 4726 28846 4738
rect 28788 4150 28800 4726
rect 28834 4150 28846 4726
rect 28788 4138 28846 4150
rect 29806 4726 29864 4738
rect 29806 4150 29818 4726
rect 29852 4150 29864 4726
rect 29806 4138 29864 4150
rect 30824 4726 30882 4738
rect 30824 4150 30836 4726
rect 30870 4150 30882 4726
rect 30824 4138 30882 4150
rect 31842 4726 31900 4738
rect 31842 4150 31854 4726
rect 31888 4150 31900 4726
rect 31842 4138 31900 4150
rect 32860 4726 32918 4738
rect 32860 4150 32872 4726
rect 32906 4150 32918 4726
rect 32860 4138 32918 4150
rect 33878 4726 33936 4738
rect 33878 4150 33890 4726
rect 33924 4150 33936 4726
rect 33878 4138 33936 4150
rect 430 3872 488 3884
rect 430 3296 442 3872
rect 476 3296 488 3872
rect 430 3284 488 3296
rect 1448 3872 1506 3884
rect 1448 3296 1460 3872
rect 1494 3296 1506 3872
rect 1448 3284 1506 3296
rect 2466 3872 2524 3884
rect 2466 3296 2478 3872
rect 2512 3296 2524 3872
rect 2466 3284 2524 3296
rect 3484 3872 3542 3884
rect 3484 3296 3496 3872
rect 3530 3296 3542 3872
rect 3484 3284 3542 3296
rect 4502 3872 4560 3884
rect 4502 3296 4514 3872
rect 4548 3296 4560 3872
rect 4502 3284 4560 3296
rect 5520 3872 5578 3884
rect 5520 3296 5532 3872
rect 5566 3296 5578 3872
rect 5520 3284 5578 3296
rect 6538 3872 6596 3884
rect 6538 3296 6550 3872
rect 6584 3296 6596 3872
rect 6538 3284 6596 3296
rect 7556 3872 7614 3884
rect 7556 3296 7568 3872
rect 7602 3296 7614 3872
rect 7556 3284 7614 3296
rect 8574 3872 8632 3884
rect 8574 3296 8586 3872
rect 8620 3296 8632 3872
rect 8574 3284 8632 3296
rect 9592 3872 9650 3884
rect 9592 3296 9604 3872
rect 9638 3296 9650 3872
rect 9592 3284 9650 3296
rect 10610 3872 10668 3884
rect 10610 3296 10622 3872
rect 10656 3296 10668 3872
rect 10610 3284 10668 3296
rect 11628 3872 11686 3884
rect 11628 3296 11640 3872
rect 11674 3296 11686 3872
rect 11628 3284 11686 3296
rect 13518 3494 13576 3506
rect 13518 2918 13530 3494
rect 13564 2918 13576 3494
rect 13518 2906 13576 2918
rect 14536 3494 14594 3506
rect 14536 2918 14548 3494
rect 14582 2918 14594 3494
rect 14536 2906 14594 2918
rect 15554 3494 15612 3506
rect 15554 2918 15566 3494
rect 15600 2918 15612 3494
rect 15554 2906 15612 2918
rect 16572 3494 16630 3506
rect 16572 2918 16584 3494
rect 16618 2918 16630 3494
rect 16572 2906 16630 2918
rect 17590 3494 17648 3506
rect 17590 2918 17602 3494
rect 17636 2918 17648 3494
rect 17590 2906 17648 2918
rect 18608 3494 18666 3506
rect 18608 2918 18620 3494
rect 18654 2918 18666 3494
rect 18608 2906 18666 2918
rect 19626 3494 19684 3506
rect 19626 2918 19638 3494
rect 19672 2918 19684 3494
rect 19626 2906 19684 2918
rect 20644 3494 20702 3506
rect 20644 2918 20656 3494
rect 20690 2918 20702 3494
rect 20644 2906 20702 2918
rect 21662 3494 21720 3506
rect 21662 2918 21674 3494
rect 21708 2918 21720 3494
rect 21662 2906 21720 2918
rect 22680 3494 22738 3506
rect 22680 2918 22692 3494
rect 22726 2918 22738 3494
rect 22680 2906 22738 2918
rect 23698 3494 23756 3506
rect 23698 2918 23710 3494
rect 23744 2918 23756 3494
rect 23698 2906 23756 2918
rect 24716 3494 24774 3506
rect 24716 2918 24728 3494
rect 24762 2918 24774 3494
rect 24716 2906 24774 2918
rect 25734 3494 25792 3506
rect 25734 2918 25746 3494
rect 25780 2918 25792 3494
rect 25734 2906 25792 2918
rect 26752 3494 26810 3506
rect 26752 2918 26764 3494
rect 26798 2918 26810 3494
rect 26752 2906 26810 2918
rect 27770 3494 27828 3506
rect 27770 2918 27782 3494
rect 27816 2918 27828 3494
rect 27770 2906 27828 2918
rect 28788 3494 28846 3506
rect 28788 2918 28800 3494
rect 28834 2918 28846 3494
rect 28788 2906 28846 2918
rect 29806 3494 29864 3506
rect 29806 2918 29818 3494
rect 29852 2918 29864 3494
rect 29806 2906 29864 2918
rect 30824 3494 30882 3506
rect 30824 2918 30836 3494
rect 30870 2918 30882 3494
rect 30824 2906 30882 2918
rect 31842 3494 31900 3506
rect 31842 2918 31854 3494
rect 31888 2918 31900 3494
rect 31842 2906 31900 2918
rect 32860 3494 32918 3506
rect 32860 2918 32872 3494
rect 32906 2918 32918 3494
rect 32860 2906 32918 2918
rect 33878 3494 33936 3506
rect 33878 2918 33890 3494
rect 33924 2918 33936 3494
rect 33878 2906 33936 2918
rect 430 2760 488 2772
rect 430 2184 442 2760
rect 476 2184 488 2760
rect 430 2172 488 2184
rect 1448 2760 1506 2772
rect 1448 2184 1460 2760
rect 1494 2184 1506 2760
rect 1448 2172 1506 2184
rect 2466 2760 2524 2772
rect 2466 2184 2478 2760
rect 2512 2184 2524 2760
rect 2466 2172 2524 2184
rect 3484 2760 3542 2772
rect 3484 2184 3496 2760
rect 3530 2184 3542 2760
rect 3484 2172 3542 2184
rect 4502 2760 4560 2772
rect 4502 2184 4514 2760
rect 4548 2184 4560 2760
rect 4502 2172 4560 2184
rect 5520 2760 5578 2772
rect 5520 2184 5532 2760
rect 5566 2184 5578 2760
rect 5520 2172 5578 2184
rect 6538 2760 6596 2772
rect 6538 2184 6550 2760
rect 6584 2184 6596 2760
rect 6538 2172 6596 2184
rect 7556 2760 7614 2772
rect 7556 2184 7568 2760
rect 7602 2184 7614 2760
rect 7556 2172 7614 2184
rect 8574 2760 8632 2772
rect 8574 2184 8586 2760
rect 8620 2184 8632 2760
rect 8574 2172 8632 2184
rect 9592 2760 9650 2772
rect 9592 2184 9604 2760
rect 9638 2184 9650 2760
rect 9592 2172 9650 2184
rect 10610 2760 10668 2772
rect 10610 2184 10622 2760
rect 10656 2184 10668 2760
rect 10610 2172 10668 2184
rect 11628 2760 11686 2772
rect 11628 2184 11640 2760
rect 11674 2184 11686 2760
rect 11628 2172 11686 2184
rect 13518 2260 13576 2272
rect 13518 1684 13530 2260
rect 13564 1684 13576 2260
rect 13518 1672 13576 1684
rect 14536 2260 14594 2272
rect 14536 1684 14548 2260
rect 14582 1684 14594 2260
rect 14536 1672 14594 1684
rect 15554 2260 15612 2272
rect 15554 1684 15566 2260
rect 15600 1684 15612 2260
rect 15554 1672 15612 1684
rect 16572 2260 16630 2272
rect 16572 1684 16584 2260
rect 16618 1684 16630 2260
rect 16572 1672 16630 1684
rect 17590 2260 17648 2272
rect 17590 1684 17602 2260
rect 17636 1684 17648 2260
rect 17590 1672 17648 1684
rect 18608 2260 18666 2272
rect 18608 1684 18620 2260
rect 18654 1684 18666 2260
rect 18608 1672 18666 1684
rect 19626 2260 19684 2272
rect 19626 1684 19638 2260
rect 19672 1684 19684 2260
rect 19626 1672 19684 1684
rect 20644 2260 20702 2272
rect 20644 1684 20656 2260
rect 20690 1684 20702 2260
rect 20644 1672 20702 1684
rect 21662 2260 21720 2272
rect 21662 1684 21674 2260
rect 21708 1684 21720 2260
rect 21662 1672 21720 1684
rect 22680 2260 22738 2272
rect 22680 1684 22692 2260
rect 22726 1684 22738 2260
rect 22680 1672 22738 1684
rect 23698 2260 23756 2272
rect 23698 1684 23710 2260
rect 23744 1684 23756 2260
rect 23698 1672 23756 1684
rect 24716 2260 24774 2272
rect 24716 1684 24728 2260
rect 24762 1684 24774 2260
rect 24716 1672 24774 1684
rect 25734 2260 25792 2272
rect 25734 1684 25746 2260
rect 25780 1684 25792 2260
rect 25734 1672 25792 1684
rect 26752 2260 26810 2272
rect 26752 1684 26764 2260
rect 26798 1684 26810 2260
rect 26752 1672 26810 1684
rect 27770 2260 27828 2272
rect 27770 1684 27782 2260
rect 27816 1684 27828 2260
rect 27770 1672 27828 1684
rect 28788 2260 28846 2272
rect 28788 1684 28800 2260
rect 28834 1684 28846 2260
rect 28788 1672 28846 1684
rect 29806 2260 29864 2272
rect 29806 1684 29818 2260
rect 29852 1684 29864 2260
rect 29806 1672 29864 1684
rect 30824 2260 30882 2272
rect 30824 1684 30836 2260
rect 30870 1684 30882 2260
rect 30824 1672 30882 1684
rect 31842 2260 31900 2272
rect 31842 1684 31854 2260
rect 31888 1684 31900 2260
rect 31842 1672 31900 1684
rect 32860 2260 32918 2272
rect 32860 1684 32872 2260
rect 32906 1684 32918 2260
rect 32860 1672 32918 1684
rect 33878 2260 33936 2272
rect 33878 1684 33890 2260
rect 33924 1684 33936 2260
rect 33878 1672 33936 1684
rect 888 1218 946 1230
rect 888 642 900 1218
rect 934 642 946 1218
rect 888 630 946 642
rect 1906 1218 1964 1230
rect 1906 642 1918 1218
rect 1952 642 1964 1218
rect 1906 630 1964 642
rect 2924 1218 2982 1230
rect 2924 642 2936 1218
rect 2970 642 2982 1218
rect 2924 630 2982 642
rect 3942 1218 4000 1230
rect 3942 642 3954 1218
rect 3988 642 4000 1218
rect 3942 630 4000 642
rect 4960 1218 5018 1230
rect 4960 642 4972 1218
rect 5006 642 5018 1218
rect 4960 630 5018 642
rect 5978 1218 6036 1230
rect 5978 642 5990 1218
rect 6024 642 6036 1218
rect 5978 630 6036 642
rect 6996 1218 7054 1230
rect 6996 642 7008 1218
rect 7042 642 7054 1218
rect 6996 630 7054 642
rect 8014 1218 8072 1230
rect 8014 642 8026 1218
rect 8060 642 8072 1218
rect 8014 630 8072 642
rect 9032 1218 9090 1230
rect 9032 642 9044 1218
rect 9078 642 9090 1218
rect 9032 630 9090 642
rect 10050 1218 10108 1230
rect 10050 642 10062 1218
rect 10096 642 10108 1218
rect 10050 630 10108 642
rect 11068 1218 11126 1230
rect 11068 642 11080 1218
rect 11114 642 11126 1218
rect 11068 630 11126 642
rect 13518 1028 13576 1040
rect 13518 452 13530 1028
rect 13564 452 13576 1028
rect 13518 440 13576 452
rect 14536 1028 14594 1040
rect 14536 452 14548 1028
rect 14582 452 14594 1028
rect 14536 440 14594 452
rect 15554 1028 15612 1040
rect 15554 452 15566 1028
rect 15600 452 15612 1028
rect 15554 440 15612 452
rect 16572 1028 16630 1040
rect 16572 452 16584 1028
rect 16618 452 16630 1028
rect 16572 440 16630 452
rect 17590 1028 17648 1040
rect 17590 452 17602 1028
rect 17636 452 17648 1028
rect 17590 440 17648 452
rect 18608 1028 18666 1040
rect 18608 452 18620 1028
rect 18654 452 18666 1028
rect 18608 440 18666 452
rect 19626 1028 19684 1040
rect 19626 452 19638 1028
rect 19672 452 19684 1028
rect 19626 440 19684 452
rect 20644 1028 20702 1040
rect 20644 452 20656 1028
rect 20690 452 20702 1028
rect 20644 440 20702 452
rect 21662 1028 21720 1040
rect 21662 452 21674 1028
rect 21708 452 21720 1028
rect 21662 440 21720 452
rect 22680 1028 22738 1040
rect 22680 452 22692 1028
rect 22726 452 22738 1028
rect 22680 440 22738 452
rect 23698 1028 23756 1040
rect 23698 452 23710 1028
rect 23744 452 23756 1028
rect 23698 440 23756 452
rect 24716 1028 24774 1040
rect 24716 452 24728 1028
rect 24762 452 24774 1028
rect 24716 440 24774 452
rect 25734 1028 25792 1040
rect 25734 452 25746 1028
rect 25780 452 25792 1028
rect 25734 440 25792 452
rect 26752 1028 26810 1040
rect 26752 452 26764 1028
rect 26798 452 26810 1028
rect 26752 440 26810 452
rect 27770 1028 27828 1040
rect 27770 452 27782 1028
rect 27816 452 27828 1028
rect 27770 440 27828 452
rect 28788 1028 28846 1040
rect 28788 452 28800 1028
rect 28834 452 28846 1028
rect 28788 440 28846 452
rect 29806 1028 29864 1040
rect 29806 452 29818 1028
rect 29852 452 29864 1028
rect 29806 440 29864 452
rect 30824 1028 30882 1040
rect 30824 452 30836 1028
rect 30870 452 30882 1028
rect 30824 440 30882 452
rect 31842 1028 31900 1040
rect 31842 452 31854 1028
rect 31888 452 31900 1028
rect 31842 440 31900 452
rect 32860 1028 32918 1040
rect 32860 452 32872 1028
rect 32906 452 32918 1028
rect 32860 440 32918 452
rect 33878 1028 33936 1040
rect 33878 452 33890 1028
rect 33924 452 33936 1028
rect 33878 440 33936 452
rect -1086 190 -1028 202
rect -1086 84 -1074 190
rect -1040 84 -1028 190
rect -1086 72 -1028 84
rect -998 190 -940 202
rect -998 84 -986 190
rect -952 84 -940 190
rect -998 72 -940 84
rect 54520 14322 54578 14334
rect 42754 13846 42812 13858
rect 42754 13270 42766 13846
rect 42800 13270 42812 13846
rect 42754 13258 42812 13270
rect 43772 13846 43830 13858
rect 43772 13270 43784 13846
rect 43818 13270 43830 13846
rect 43772 13258 43830 13270
rect 44790 13846 44848 13858
rect 44790 13270 44802 13846
rect 44836 13270 44848 13846
rect 44790 13258 44848 13270
rect 45808 13846 45866 13858
rect 45808 13270 45820 13846
rect 45854 13270 45866 13846
rect 45808 13258 45866 13270
rect 46826 13846 46884 13858
rect 46826 13270 46838 13846
rect 46872 13270 46884 13846
rect 46826 13258 46884 13270
rect 47844 13846 47902 13858
rect 47844 13270 47856 13846
rect 47890 13270 47902 13846
rect 47844 13258 47902 13270
rect 48862 13846 48920 13858
rect 48862 13270 48874 13846
rect 48908 13270 48920 13846
rect 48862 13258 48920 13270
rect 49880 13846 49938 13858
rect 49880 13270 49892 13846
rect 49926 13270 49938 13846
rect 49880 13258 49938 13270
rect 50898 13846 50956 13858
rect 50898 13270 50910 13846
rect 50944 13270 50956 13846
rect 50898 13258 50956 13270
rect 51916 13846 51974 13858
rect 51916 13270 51928 13846
rect 51962 13270 51974 13846
rect 54520 13746 54532 14322
rect 54566 13746 54578 14322
rect 54520 13734 54578 13746
rect 55538 14322 55596 14334
rect 55538 13746 55550 14322
rect 55584 13746 55596 14322
rect 55538 13734 55596 13746
rect 56556 14322 56614 14334
rect 56556 13746 56568 14322
rect 56602 13746 56614 14322
rect 56556 13734 56614 13746
rect 57574 14322 57632 14334
rect 57574 13746 57586 14322
rect 57620 13746 57632 14322
rect 57574 13734 57632 13746
rect 58592 14322 58650 14334
rect 58592 13746 58604 14322
rect 58638 13746 58650 14322
rect 58592 13734 58650 13746
rect 59610 14322 59668 14334
rect 59610 13746 59622 14322
rect 59656 13746 59668 14322
rect 59610 13734 59668 13746
rect 60628 14322 60686 14334
rect 60628 13746 60640 14322
rect 60674 13746 60686 14322
rect 60628 13734 60686 13746
rect 61646 14322 61704 14334
rect 61646 13746 61658 14322
rect 61692 13746 61704 14322
rect 61646 13734 61704 13746
rect 62664 14322 62722 14334
rect 62664 13746 62676 14322
rect 62710 13746 62722 14322
rect 62664 13734 62722 13746
rect 63682 14322 63740 14334
rect 63682 13746 63694 14322
rect 63728 13746 63740 14322
rect 63682 13734 63740 13746
rect 64700 14322 64758 14334
rect 64700 13746 64712 14322
rect 64746 13746 64758 14322
rect 64700 13734 64758 13746
rect 65718 14322 65776 14334
rect 65718 13746 65730 14322
rect 65764 13746 65776 14322
rect 65718 13734 65776 13746
rect 66736 14322 66794 14334
rect 66736 13746 66748 14322
rect 66782 13746 66794 14322
rect 66736 13734 66794 13746
rect 67754 14322 67812 14334
rect 67754 13746 67766 14322
rect 67800 13746 67812 14322
rect 67754 13734 67812 13746
rect 68772 14322 68830 14334
rect 68772 13746 68784 14322
rect 68818 13746 68830 14322
rect 68772 13734 68830 13746
rect 69790 14322 69848 14334
rect 69790 13746 69802 14322
rect 69836 13746 69848 14322
rect 69790 13734 69848 13746
rect 70808 14322 70866 14334
rect 70808 13746 70820 14322
rect 70854 13746 70866 14322
rect 70808 13734 70866 13746
rect 71826 14322 71884 14334
rect 71826 13746 71838 14322
rect 71872 13746 71884 14322
rect 71826 13734 71884 13746
rect 72844 14322 72902 14334
rect 72844 13746 72856 14322
rect 72890 13746 72902 14322
rect 72844 13734 72902 13746
rect 73862 14322 73920 14334
rect 73862 13746 73874 14322
rect 73908 13746 73920 14322
rect 73862 13734 73920 13746
rect 74880 14322 74938 14334
rect 74880 13746 74892 14322
rect 74926 13746 74938 14322
rect 74880 13734 74938 13746
rect 51916 13258 51974 13270
rect 54520 13504 54578 13516
rect 42754 13028 42812 13040
rect 42754 12452 42766 13028
rect 42800 12452 42812 13028
rect 42754 12440 42812 12452
rect 43772 13028 43830 13040
rect 43772 12452 43784 13028
rect 43818 12452 43830 13028
rect 43772 12440 43830 12452
rect 44790 13028 44848 13040
rect 44790 12452 44802 13028
rect 44836 12452 44848 13028
rect 44790 12440 44848 12452
rect 45808 13028 45866 13040
rect 45808 12452 45820 13028
rect 45854 12452 45866 13028
rect 45808 12440 45866 12452
rect 46826 13028 46884 13040
rect 46826 12452 46838 13028
rect 46872 12452 46884 13028
rect 46826 12440 46884 12452
rect 47844 13028 47902 13040
rect 47844 12452 47856 13028
rect 47890 12452 47902 13028
rect 47844 12440 47902 12452
rect 48862 13028 48920 13040
rect 48862 12452 48874 13028
rect 48908 12452 48920 13028
rect 48862 12440 48920 12452
rect 49880 13028 49938 13040
rect 49880 12452 49892 13028
rect 49926 12452 49938 13028
rect 49880 12440 49938 12452
rect 50898 13028 50956 13040
rect 50898 12452 50910 13028
rect 50944 12452 50956 13028
rect 50898 12440 50956 12452
rect 51916 13028 51974 13040
rect 51916 12452 51928 13028
rect 51962 12452 51974 13028
rect 54520 12928 54532 13504
rect 54566 12928 54578 13504
rect 54520 12916 54578 12928
rect 55538 13504 55596 13516
rect 55538 12928 55550 13504
rect 55584 12928 55596 13504
rect 55538 12916 55596 12928
rect 56556 13504 56614 13516
rect 56556 12928 56568 13504
rect 56602 12928 56614 13504
rect 56556 12916 56614 12928
rect 57574 13504 57632 13516
rect 57574 12928 57586 13504
rect 57620 12928 57632 13504
rect 57574 12916 57632 12928
rect 58592 13504 58650 13516
rect 58592 12928 58604 13504
rect 58638 12928 58650 13504
rect 58592 12916 58650 12928
rect 59610 13504 59668 13516
rect 59610 12928 59622 13504
rect 59656 12928 59668 13504
rect 59610 12916 59668 12928
rect 60628 13504 60686 13516
rect 60628 12928 60640 13504
rect 60674 12928 60686 13504
rect 60628 12916 60686 12928
rect 61646 13504 61704 13516
rect 61646 12928 61658 13504
rect 61692 12928 61704 13504
rect 61646 12916 61704 12928
rect 62664 13504 62722 13516
rect 62664 12928 62676 13504
rect 62710 12928 62722 13504
rect 62664 12916 62722 12928
rect 63682 13504 63740 13516
rect 63682 12928 63694 13504
rect 63728 12928 63740 13504
rect 63682 12916 63740 12928
rect 64700 13504 64758 13516
rect 64700 12928 64712 13504
rect 64746 12928 64758 13504
rect 64700 12916 64758 12928
rect 65718 13504 65776 13516
rect 65718 12928 65730 13504
rect 65764 12928 65776 13504
rect 65718 12916 65776 12928
rect 66736 13504 66794 13516
rect 66736 12928 66748 13504
rect 66782 12928 66794 13504
rect 66736 12916 66794 12928
rect 67754 13504 67812 13516
rect 67754 12928 67766 13504
rect 67800 12928 67812 13504
rect 67754 12916 67812 12928
rect 68772 13504 68830 13516
rect 68772 12928 68784 13504
rect 68818 12928 68830 13504
rect 68772 12916 68830 12928
rect 69790 13504 69848 13516
rect 69790 12928 69802 13504
rect 69836 12928 69848 13504
rect 69790 12916 69848 12928
rect 70808 13504 70866 13516
rect 70808 12928 70820 13504
rect 70854 12928 70866 13504
rect 70808 12916 70866 12928
rect 71826 13504 71884 13516
rect 71826 12928 71838 13504
rect 71872 12928 71884 13504
rect 71826 12916 71884 12928
rect 72844 13504 72902 13516
rect 72844 12928 72856 13504
rect 72890 12928 72902 13504
rect 72844 12916 72902 12928
rect 73862 13504 73920 13516
rect 73862 12928 73874 13504
rect 73908 12928 73920 13504
rect 73862 12916 73920 12928
rect 74880 13504 74938 13516
rect 74880 12928 74892 13504
rect 74926 12928 74938 13504
rect 74880 12916 74938 12928
rect 51916 12440 51974 12452
rect 42754 12210 42812 12222
rect 42754 11634 42766 12210
rect 42800 11634 42812 12210
rect 42754 11622 42812 11634
rect 43772 12210 43830 12222
rect 43772 11634 43784 12210
rect 43818 11634 43830 12210
rect 43772 11622 43830 11634
rect 44790 12210 44848 12222
rect 44790 11634 44802 12210
rect 44836 11634 44848 12210
rect 44790 11622 44848 11634
rect 45808 12210 45866 12222
rect 45808 11634 45820 12210
rect 45854 11634 45866 12210
rect 45808 11622 45866 11634
rect 46826 12210 46884 12222
rect 46826 11634 46838 12210
rect 46872 11634 46884 12210
rect 46826 11622 46884 11634
rect 47844 12210 47902 12222
rect 47844 11634 47856 12210
rect 47890 11634 47902 12210
rect 47844 11622 47902 11634
rect 48862 12210 48920 12222
rect 48862 11634 48874 12210
rect 48908 11634 48920 12210
rect 48862 11622 48920 11634
rect 49880 12210 49938 12222
rect 49880 11634 49892 12210
rect 49926 11634 49938 12210
rect 49880 11622 49938 11634
rect 50898 12210 50956 12222
rect 50898 11634 50910 12210
rect 50944 11634 50956 12210
rect 50898 11622 50956 11634
rect 51916 12210 51974 12222
rect 51916 11634 51928 12210
rect 51962 11634 51974 12210
rect 51916 11622 51974 11634
rect 54520 12126 54578 12138
rect 54520 11550 54532 12126
rect 54566 11550 54578 12126
rect 54520 11538 54578 11550
rect 55538 12126 55596 12138
rect 55538 11550 55550 12126
rect 55584 11550 55596 12126
rect 55538 11538 55596 11550
rect 56556 12126 56614 12138
rect 56556 11550 56568 12126
rect 56602 11550 56614 12126
rect 56556 11538 56614 11550
rect 57574 12126 57632 12138
rect 57574 11550 57586 12126
rect 57620 11550 57632 12126
rect 57574 11538 57632 11550
rect 58592 12126 58650 12138
rect 58592 11550 58604 12126
rect 58638 11550 58650 12126
rect 58592 11538 58650 11550
rect 59610 12126 59668 12138
rect 59610 11550 59622 12126
rect 59656 11550 59668 12126
rect 59610 11538 59668 11550
rect 60628 12126 60686 12138
rect 60628 11550 60640 12126
rect 60674 11550 60686 12126
rect 60628 11538 60686 11550
rect 61646 12126 61704 12138
rect 61646 11550 61658 12126
rect 61692 11550 61704 12126
rect 61646 11538 61704 11550
rect 62664 12126 62722 12138
rect 62664 11550 62676 12126
rect 62710 11550 62722 12126
rect 62664 11538 62722 11550
rect 63682 12126 63740 12138
rect 63682 11550 63694 12126
rect 63728 11550 63740 12126
rect 63682 11538 63740 11550
rect 64700 12126 64758 12138
rect 64700 11550 64712 12126
rect 64746 11550 64758 12126
rect 64700 11538 64758 11550
rect 65718 12126 65776 12138
rect 65718 11550 65730 12126
rect 65764 11550 65776 12126
rect 65718 11538 65776 11550
rect 66736 12126 66794 12138
rect 66736 11550 66748 12126
rect 66782 11550 66794 12126
rect 66736 11538 66794 11550
rect 67754 12126 67812 12138
rect 67754 11550 67766 12126
rect 67800 11550 67812 12126
rect 67754 11538 67812 11550
rect 68772 12126 68830 12138
rect 68772 11550 68784 12126
rect 68818 11550 68830 12126
rect 68772 11538 68830 11550
rect 69790 12126 69848 12138
rect 69790 11550 69802 12126
rect 69836 11550 69848 12126
rect 69790 11538 69848 11550
rect 70808 12126 70866 12138
rect 70808 11550 70820 12126
rect 70854 11550 70866 12126
rect 70808 11538 70866 11550
rect 71826 12126 71884 12138
rect 71826 11550 71838 12126
rect 71872 11550 71884 12126
rect 71826 11538 71884 11550
rect 72844 12126 72902 12138
rect 72844 11550 72856 12126
rect 72890 11550 72902 12126
rect 72844 11538 72902 11550
rect 73862 12126 73920 12138
rect 73862 11550 73874 12126
rect 73908 11550 73920 12126
rect 73862 11538 73920 11550
rect 74880 12126 74938 12138
rect 74880 11550 74892 12126
rect 74926 11550 74938 12126
rect 74880 11538 74938 11550
rect 42754 11392 42812 11404
rect 42754 10816 42766 11392
rect 42800 10816 42812 11392
rect 42754 10804 42812 10816
rect 43772 11392 43830 11404
rect 43772 10816 43784 11392
rect 43818 10816 43830 11392
rect 43772 10804 43830 10816
rect 44790 11392 44848 11404
rect 44790 10816 44802 11392
rect 44836 10816 44848 11392
rect 44790 10804 44848 10816
rect 45808 11392 45866 11404
rect 45808 10816 45820 11392
rect 45854 10816 45866 11392
rect 45808 10804 45866 10816
rect 46826 11392 46884 11404
rect 46826 10816 46838 11392
rect 46872 10816 46884 11392
rect 46826 10804 46884 10816
rect 47844 11392 47902 11404
rect 47844 10816 47856 11392
rect 47890 10816 47902 11392
rect 47844 10804 47902 10816
rect 48862 11392 48920 11404
rect 48862 10816 48874 11392
rect 48908 10816 48920 11392
rect 48862 10804 48920 10816
rect 49880 11392 49938 11404
rect 49880 10816 49892 11392
rect 49926 10816 49938 11392
rect 49880 10804 49938 10816
rect 50898 11392 50956 11404
rect 50898 10816 50910 11392
rect 50944 10816 50956 11392
rect 50898 10804 50956 10816
rect 51916 11392 51974 11404
rect 51916 10816 51928 11392
rect 51962 10816 51974 11392
rect 51916 10804 51974 10816
rect 54520 10894 54578 10906
rect 42754 10574 42812 10586
rect 42754 9998 42766 10574
rect 42800 9998 42812 10574
rect 42754 9986 42812 9998
rect 43772 10574 43830 10586
rect 43772 9998 43784 10574
rect 43818 9998 43830 10574
rect 43772 9986 43830 9998
rect 44790 10574 44848 10586
rect 44790 9998 44802 10574
rect 44836 9998 44848 10574
rect 44790 9986 44848 9998
rect 45808 10574 45866 10586
rect 45808 9998 45820 10574
rect 45854 9998 45866 10574
rect 45808 9986 45866 9998
rect 46826 10574 46884 10586
rect 46826 9998 46838 10574
rect 46872 9998 46884 10574
rect 46826 9986 46884 9998
rect 47844 10574 47902 10586
rect 47844 9998 47856 10574
rect 47890 9998 47902 10574
rect 47844 9986 47902 9998
rect 48862 10574 48920 10586
rect 48862 9998 48874 10574
rect 48908 9998 48920 10574
rect 48862 9986 48920 9998
rect 49880 10574 49938 10586
rect 49880 9998 49892 10574
rect 49926 9998 49938 10574
rect 49880 9986 49938 9998
rect 50898 10574 50956 10586
rect 50898 9998 50910 10574
rect 50944 9998 50956 10574
rect 50898 9986 50956 9998
rect 51916 10574 51974 10586
rect 51916 9998 51928 10574
rect 51962 9998 51974 10574
rect 54520 10318 54532 10894
rect 54566 10318 54578 10894
rect 54520 10306 54578 10318
rect 55538 10894 55596 10906
rect 55538 10318 55550 10894
rect 55584 10318 55596 10894
rect 55538 10306 55596 10318
rect 56556 10894 56614 10906
rect 56556 10318 56568 10894
rect 56602 10318 56614 10894
rect 56556 10306 56614 10318
rect 57574 10894 57632 10906
rect 57574 10318 57586 10894
rect 57620 10318 57632 10894
rect 57574 10306 57632 10318
rect 58592 10894 58650 10906
rect 58592 10318 58604 10894
rect 58638 10318 58650 10894
rect 58592 10306 58650 10318
rect 59610 10894 59668 10906
rect 59610 10318 59622 10894
rect 59656 10318 59668 10894
rect 59610 10306 59668 10318
rect 60628 10894 60686 10906
rect 60628 10318 60640 10894
rect 60674 10318 60686 10894
rect 60628 10306 60686 10318
rect 61646 10894 61704 10906
rect 61646 10318 61658 10894
rect 61692 10318 61704 10894
rect 61646 10306 61704 10318
rect 62664 10894 62722 10906
rect 62664 10318 62676 10894
rect 62710 10318 62722 10894
rect 62664 10306 62722 10318
rect 63682 10894 63740 10906
rect 63682 10318 63694 10894
rect 63728 10318 63740 10894
rect 63682 10306 63740 10318
rect 64700 10894 64758 10906
rect 64700 10318 64712 10894
rect 64746 10318 64758 10894
rect 64700 10306 64758 10318
rect 65718 10894 65776 10906
rect 65718 10318 65730 10894
rect 65764 10318 65776 10894
rect 65718 10306 65776 10318
rect 66736 10894 66794 10906
rect 66736 10318 66748 10894
rect 66782 10318 66794 10894
rect 66736 10306 66794 10318
rect 67754 10894 67812 10906
rect 67754 10318 67766 10894
rect 67800 10318 67812 10894
rect 67754 10306 67812 10318
rect 68772 10894 68830 10906
rect 68772 10318 68784 10894
rect 68818 10318 68830 10894
rect 68772 10306 68830 10318
rect 69790 10894 69848 10906
rect 69790 10318 69802 10894
rect 69836 10318 69848 10894
rect 69790 10306 69848 10318
rect 70808 10894 70866 10906
rect 70808 10318 70820 10894
rect 70854 10318 70866 10894
rect 70808 10306 70866 10318
rect 71826 10894 71884 10906
rect 71826 10318 71838 10894
rect 71872 10318 71884 10894
rect 71826 10306 71884 10318
rect 72844 10894 72902 10906
rect 72844 10318 72856 10894
rect 72890 10318 72902 10894
rect 72844 10306 72902 10318
rect 73862 10894 73920 10906
rect 73862 10318 73874 10894
rect 73908 10318 73920 10894
rect 73862 10306 73920 10318
rect 74880 10894 74938 10906
rect 74880 10318 74892 10894
rect 74926 10318 74938 10894
rect 74880 10306 74938 10318
rect 51916 9986 51974 9998
rect 42754 9756 42812 9768
rect 42754 9180 42766 9756
rect 42800 9180 42812 9756
rect 42754 9168 42812 9180
rect 43772 9756 43830 9768
rect 43772 9180 43784 9756
rect 43818 9180 43830 9756
rect 43772 9168 43830 9180
rect 44790 9756 44848 9768
rect 44790 9180 44802 9756
rect 44836 9180 44848 9756
rect 44790 9168 44848 9180
rect 45808 9756 45866 9768
rect 45808 9180 45820 9756
rect 45854 9180 45866 9756
rect 45808 9168 45866 9180
rect 46826 9756 46884 9768
rect 46826 9180 46838 9756
rect 46872 9180 46884 9756
rect 46826 9168 46884 9180
rect 47844 9756 47902 9768
rect 47844 9180 47856 9756
rect 47890 9180 47902 9756
rect 47844 9168 47902 9180
rect 48862 9756 48920 9768
rect 48862 9180 48874 9756
rect 48908 9180 48920 9756
rect 48862 9168 48920 9180
rect 49880 9756 49938 9768
rect 49880 9180 49892 9756
rect 49926 9180 49938 9756
rect 49880 9168 49938 9180
rect 50898 9756 50956 9768
rect 50898 9180 50910 9756
rect 50944 9180 50956 9756
rect 50898 9168 50956 9180
rect 51916 9756 51974 9768
rect 51916 9180 51928 9756
rect 51962 9180 51974 9756
rect 51916 9168 51974 9180
rect 54518 9660 54576 9672
rect 54518 9084 54530 9660
rect 54564 9084 54576 9660
rect 54518 9072 54576 9084
rect 55536 9660 55594 9672
rect 55536 9084 55548 9660
rect 55582 9084 55594 9660
rect 55536 9072 55594 9084
rect 56554 9660 56612 9672
rect 56554 9084 56566 9660
rect 56600 9084 56612 9660
rect 56554 9072 56612 9084
rect 57572 9660 57630 9672
rect 57572 9084 57584 9660
rect 57618 9084 57630 9660
rect 57572 9072 57630 9084
rect 58590 9660 58648 9672
rect 58590 9084 58602 9660
rect 58636 9084 58648 9660
rect 58590 9072 58648 9084
rect 59608 9660 59666 9672
rect 59608 9084 59620 9660
rect 59654 9084 59666 9660
rect 59608 9072 59666 9084
rect 60626 9660 60684 9672
rect 60626 9084 60638 9660
rect 60672 9084 60684 9660
rect 60626 9072 60684 9084
rect 61644 9660 61702 9672
rect 61644 9084 61656 9660
rect 61690 9084 61702 9660
rect 61644 9072 61702 9084
rect 62662 9660 62720 9672
rect 62662 9084 62674 9660
rect 62708 9084 62720 9660
rect 62662 9072 62720 9084
rect 63680 9660 63738 9672
rect 63680 9084 63692 9660
rect 63726 9084 63738 9660
rect 63680 9072 63738 9084
rect 64698 9660 64756 9672
rect 64698 9084 64710 9660
rect 64744 9084 64756 9660
rect 64698 9072 64756 9084
rect 65716 9660 65774 9672
rect 65716 9084 65728 9660
rect 65762 9084 65774 9660
rect 65716 9072 65774 9084
rect 66734 9660 66792 9672
rect 66734 9084 66746 9660
rect 66780 9084 66792 9660
rect 66734 9072 66792 9084
rect 67752 9660 67810 9672
rect 67752 9084 67764 9660
rect 67798 9084 67810 9660
rect 67752 9072 67810 9084
rect 68770 9660 68828 9672
rect 68770 9084 68782 9660
rect 68816 9084 68828 9660
rect 68770 9072 68828 9084
rect 69788 9660 69846 9672
rect 69788 9084 69800 9660
rect 69834 9084 69846 9660
rect 69788 9072 69846 9084
rect 70806 9660 70864 9672
rect 70806 9084 70818 9660
rect 70852 9084 70864 9660
rect 70806 9072 70864 9084
rect 71824 9660 71882 9672
rect 71824 9084 71836 9660
rect 71870 9084 71882 9660
rect 71824 9072 71882 9084
rect 72842 9660 72900 9672
rect 72842 9084 72854 9660
rect 72888 9084 72900 9660
rect 72842 9072 72900 9084
rect 73860 9660 73918 9672
rect 73860 9084 73872 9660
rect 73906 9084 73918 9660
rect 73860 9072 73918 9084
rect 74878 9660 74936 9672
rect 74878 9084 74890 9660
rect 74924 9084 74936 9660
rect 74878 9072 74936 9084
rect 42754 8938 42812 8950
rect 42754 8362 42766 8938
rect 42800 8362 42812 8938
rect 42754 8350 42812 8362
rect 43772 8938 43830 8950
rect 43772 8362 43784 8938
rect 43818 8362 43830 8938
rect 43772 8350 43830 8362
rect 44790 8938 44848 8950
rect 44790 8362 44802 8938
rect 44836 8362 44848 8938
rect 44790 8350 44848 8362
rect 45808 8938 45866 8950
rect 45808 8362 45820 8938
rect 45854 8362 45866 8938
rect 45808 8350 45866 8362
rect 46826 8938 46884 8950
rect 46826 8362 46838 8938
rect 46872 8362 46884 8938
rect 46826 8350 46884 8362
rect 47844 8938 47902 8950
rect 47844 8362 47856 8938
rect 47890 8362 47902 8938
rect 47844 8350 47902 8362
rect 48862 8938 48920 8950
rect 48862 8362 48874 8938
rect 48908 8362 48920 8938
rect 48862 8350 48920 8362
rect 49880 8938 49938 8950
rect 49880 8362 49892 8938
rect 49926 8362 49938 8938
rect 49880 8350 49938 8362
rect 50898 8938 50956 8950
rect 50898 8362 50910 8938
rect 50944 8362 50956 8938
rect 50898 8350 50956 8362
rect 51916 8938 51974 8950
rect 51916 8362 51928 8938
rect 51962 8362 51974 8938
rect 51916 8350 51974 8362
rect 54518 8426 54576 8438
rect 42754 8120 42812 8132
rect 42754 7544 42766 8120
rect 42800 7544 42812 8120
rect 42754 7532 42812 7544
rect 43772 8120 43830 8132
rect 43772 7544 43784 8120
rect 43818 7544 43830 8120
rect 43772 7532 43830 7544
rect 44790 8120 44848 8132
rect 44790 7544 44802 8120
rect 44836 7544 44848 8120
rect 44790 7532 44848 7544
rect 45808 8120 45866 8132
rect 45808 7544 45820 8120
rect 45854 7544 45866 8120
rect 45808 7532 45866 7544
rect 46826 8120 46884 8132
rect 46826 7544 46838 8120
rect 46872 7544 46884 8120
rect 46826 7532 46884 7544
rect 47844 8120 47902 8132
rect 47844 7544 47856 8120
rect 47890 7544 47902 8120
rect 47844 7532 47902 7544
rect 48862 8120 48920 8132
rect 48862 7544 48874 8120
rect 48908 7544 48920 8120
rect 48862 7532 48920 7544
rect 49880 8120 49938 8132
rect 49880 7544 49892 8120
rect 49926 7544 49938 8120
rect 49880 7532 49938 7544
rect 50898 8120 50956 8132
rect 50898 7544 50910 8120
rect 50944 7544 50956 8120
rect 50898 7532 50956 7544
rect 51916 8120 51974 8132
rect 51916 7544 51928 8120
rect 51962 7544 51974 8120
rect 54518 7850 54530 8426
rect 54564 7850 54576 8426
rect 54518 7838 54576 7850
rect 55536 8426 55594 8438
rect 55536 7850 55548 8426
rect 55582 7850 55594 8426
rect 55536 7838 55594 7850
rect 56554 8426 56612 8438
rect 56554 7850 56566 8426
rect 56600 7850 56612 8426
rect 56554 7838 56612 7850
rect 57572 8426 57630 8438
rect 57572 7850 57584 8426
rect 57618 7850 57630 8426
rect 57572 7838 57630 7850
rect 58590 8426 58648 8438
rect 58590 7850 58602 8426
rect 58636 7850 58648 8426
rect 58590 7838 58648 7850
rect 59608 8426 59666 8438
rect 59608 7850 59620 8426
rect 59654 7850 59666 8426
rect 59608 7838 59666 7850
rect 60626 8426 60684 8438
rect 60626 7850 60638 8426
rect 60672 7850 60684 8426
rect 60626 7838 60684 7850
rect 61644 8426 61702 8438
rect 61644 7850 61656 8426
rect 61690 7850 61702 8426
rect 61644 7838 61702 7850
rect 62662 8426 62720 8438
rect 62662 7850 62674 8426
rect 62708 7850 62720 8426
rect 62662 7838 62720 7850
rect 63680 8426 63738 8438
rect 63680 7850 63692 8426
rect 63726 7850 63738 8426
rect 63680 7838 63738 7850
rect 64698 8426 64756 8438
rect 64698 7850 64710 8426
rect 64744 7850 64756 8426
rect 64698 7838 64756 7850
rect 65716 8426 65774 8438
rect 65716 7850 65728 8426
rect 65762 7850 65774 8426
rect 65716 7838 65774 7850
rect 66734 8426 66792 8438
rect 66734 7850 66746 8426
rect 66780 7850 66792 8426
rect 66734 7838 66792 7850
rect 67752 8426 67810 8438
rect 67752 7850 67764 8426
rect 67798 7850 67810 8426
rect 67752 7838 67810 7850
rect 68770 8426 68828 8438
rect 68770 7850 68782 8426
rect 68816 7850 68828 8426
rect 68770 7838 68828 7850
rect 69788 8426 69846 8438
rect 69788 7850 69800 8426
rect 69834 7850 69846 8426
rect 69788 7838 69846 7850
rect 70806 8426 70864 8438
rect 70806 7850 70818 8426
rect 70852 7850 70864 8426
rect 70806 7838 70864 7850
rect 71824 8426 71882 8438
rect 71824 7850 71836 8426
rect 71870 7850 71882 8426
rect 71824 7838 71882 7850
rect 72842 8426 72900 8438
rect 72842 7850 72854 8426
rect 72888 7850 72900 8426
rect 72842 7838 72900 7850
rect 73860 8426 73918 8438
rect 73860 7850 73872 8426
rect 73906 7850 73918 8426
rect 73860 7838 73918 7850
rect 74878 8426 74936 8438
rect 74878 7850 74890 8426
rect 74924 7850 74936 8426
rect 74878 7838 74936 7850
rect 51916 7532 51974 7544
rect 54518 7194 54576 7206
rect 54518 6618 54530 7194
rect 54564 6618 54576 7194
rect 54518 6606 54576 6618
rect 55536 7194 55594 7206
rect 55536 6618 55548 7194
rect 55582 6618 55594 7194
rect 55536 6606 55594 6618
rect 56554 7194 56612 7206
rect 56554 6618 56566 7194
rect 56600 6618 56612 7194
rect 56554 6606 56612 6618
rect 57572 7194 57630 7206
rect 57572 6618 57584 7194
rect 57618 6618 57630 7194
rect 57572 6606 57630 6618
rect 58590 7194 58648 7206
rect 58590 6618 58602 7194
rect 58636 6618 58648 7194
rect 58590 6606 58648 6618
rect 59608 7194 59666 7206
rect 59608 6618 59620 7194
rect 59654 6618 59666 7194
rect 59608 6606 59666 6618
rect 60626 7194 60684 7206
rect 60626 6618 60638 7194
rect 60672 6618 60684 7194
rect 60626 6606 60684 6618
rect 61644 7194 61702 7206
rect 61644 6618 61656 7194
rect 61690 6618 61702 7194
rect 61644 6606 61702 6618
rect 62662 7194 62720 7206
rect 62662 6618 62674 7194
rect 62708 6618 62720 7194
rect 62662 6606 62720 6618
rect 63680 7194 63738 7206
rect 63680 6618 63692 7194
rect 63726 6618 63738 7194
rect 63680 6606 63738 6618
rect 64698 7194 64756 7206
rect 64698 6618 64710 7194
rect 64744 6618 64756 7194
rect 64698 6606 64756 6618
rect 65716 7194 65774 7206
rect 65716 6618 65728 7194
rect 65762 6618 65774 7194
rect 65716 6606 65774 6618
rect 66734 7194 66792 7206
rect 66734 6618 66746 7194
rect 66780 6618 66792 7194
rect 66734 6606 66792 6618
rect 67752 7194 67810 7206
rect 67752 6618 67764 7194
rect 67798 6618 67810 7194
rect 67752 6606 67810 6618
rect 68770 7194 68828 7206
rect 68770 6618 68782 7194
rect 68816 6618 68828 7194
rect 68770 6606 68828 6618
rect 69788 7194 69846 7206
rect 69788 6618 69800 7194
rect 69834 6618 69846 7194
rect 69788 6606 69846 6618
rect 70806 7194 70864 7206
rect 70806 6618 70818 7194
rect 70852 6618 70864 7194
rect 70806 6606 70864 6618
rect 71824 7194 71882 7206
rect 71824 6618 71836 7194
rect 71870 6618 71882 7194
rect 71824 6606 71882 6618
rect 72842 7194 72900 7206
rect 72842 6618 72854 7194
rect 72888 6618 72900 7194
rect 72842 6606 72900 6618
rect 73860 7194 73918 7206
rect 73860 6618 73872 7194
rect 73906 6618 73918 7194
rect 73860 6606 73918 6618
rect 74878 7194 74936 7206
rect 74878 6618 74890 7194
rect 74924 6618 74936 7194
rect 74878 6606 74936 6618
rect 41430 6096 41488 6108
rect 41430 5520 41442 6096
rect 41476 5520 41488 6096
rect 41430 5508 41488 5520
rect 42448 6096 42506 6108
rect 42448 5520 42460 6096
rect 42494 5520 42506 6096
rect 42448 5508 42506 5520
rect 43466 6096 43524 6108
rect 43466 5520 43478 6096
rect 43512 5520 43524 6096
rect 43466 5508 43524 5520
rect 44484 6096 44542 6108
rect 44484 5520 44496 6096
rect 44530 5520 44542 6096
rect 44484 5508 44542 5520
rect 45502 6096 45560 6108
rect 45502 5520 45514 6096
rect 45548 5520 45560 6096
rect 45502 5508 45560 5520
rect 46520 6096 46578 6108
rect 46520 5520 46532 6096
rect 46566 5520 46578 6096
rect 46520 5508 46578 5520
rect 47538 6096 47596 6108
rect 47538 5520 47550 6096
rect 47584 5520 47596 6096
rect 47538 5508 47596 5520
rect 48556 6096 48614 6108
rect 48556 5520 48568 6096
rect 48602 5520 48614 6096
rect 48556 5508 48614 5520
rect 49574 6096 49632 6108
rect 49574 5520 49586 6096
rect 49620 5520 49632 6096
rect 49574 5508 49632 5520
rect 50592 6096 50650 6108
rect 50592 5520 50604 6096
rect 50638 5520 50650 6096
rect 50592 5508 50650 5520
rect 51610 6096 51668 6108
rect 51610 5520 51622 6096
rect 51656 5520 51668 6096
rect 51610 5508 51668 5520
rect 52628 6096 52686 6108
rect 52628 5520 52640 6096
rect 52674 5520 52686 6096
rect 52628 5508 52686 5520
rect 54518 5960 54576 5972
rect 54518 5384 54530 5960
rect 54564 5384 54576 5960
rect 54518 5372 54576 5384
rect 55536 5960 55594 5972
rect 55536 5384 55548 5960
rect 55582 5384 55594 5960
rect 55536 5372 55594 5384
rect 56554 5960 56612 5972
rect 56554 5384 56566 5960
rect 56600 5384 56612 5960
rect 56554 5372 56612 5384
rect 57572 5960 57630 5972
rect 57572 5384 57584 5960
rect 57618 5384 57630 5960
rect 57572 5372 57630 5384
rect 58590 5960 58648 5972
rect 58590 5384 58602 5960
rect 58636 5384 58648 5960
rect 58590 5372 58648 5384
rect 59608 5960 59666 5972
rect 59608 5384 59620 5960
rect 59654 5384 59666 5960
rect 59608 5372 59666 5384
rect 60626 5960 60684 5972
rect 60626 5384 60638 5960
rect 60672 5384 60684 5960
rect 60626 5372 60684 5384
rect 61644 5960 61702 5972
rect 61644 5384 61656 5960
rect 61690 5384 61702 5960
rect 61644 5372 61702 5384
rect 62662 5960 62720 5972
rect 62662 5384 62674 5960
rect 62708 5384 62720 5960
rect 62662 5372 62720 5384
rect 63680 5960 63738 5972
rect 63680 5384 63692 5960
rect 63726 5384 63738 5960
rect 63680 5372 63738 5384
rect 64698 5960 64756 5972
rect 64698 5384 64710 5960
rect 64744 5384 64756 5960
rect 64698 5372 64756 5384
rect 65716 5960 65774 5972
rect 65716 5384 65728 5960
rect 65762 5384 65774 5960
rect 65716 5372 65774 5384
rect 66734 5960 66792 5972
rect 66734 5384 66746 5960
rect 66780 5384 66792 5960
rect 66734 5372 66792 5384
rect 67752 5960 67810 5972
rect 67752 5384 67764 5960
rect 67798 5384 67810 5960
rect 67752 5372 67810 5384
rect 68770 5960 68828 5972
rect 68770 5384 68782 5960
rect 68816 5384 68828 5960
rect 68770 5372 68828 5384
rect 69788 5960 69846 5972
rect 69788 5384 69800 5960
rect 69834 5384 69846 5960
rect 69788 5372 69846 5384
rect 70806 5960 70864 5972
rect 70806 5384 70818 5960
rect 70852 5384 70864 5960
rect 70806 5372 70864 5384
rect 71824 5960 71882 5972
rect 71824 5384 71836 5960
rect 71870 5384 71882 5960
rect 71824 5372 71882 5384
rect 72842 5960 72900 5972
rect 72842 5384 72854 5960
rect 72888 5384 72900 5960
rect 72842 5372 72900 5384
rect 73860 5960 73918 5972
rect 73860 5384 73872 5960
rect 73906 5384 73918 5960
rect 73860 5372 73918 5384
rect 74878 5960 74936 5972
rect 74878 5384 74890 5960
rect 74924 5384 74936 5960
rect 74878 5372 74936 5384
rect 41430 4984 41488 4996
rect 41430 4408 41442 4984
rect 41476 4408 41488 4984
rect 41430 4396 41488 4408
rect 42448 4984 42506 4996
rect 42448 4408 42460 4984
rect 42494 4408 42506 4984
rect 42448 4396 42506 4408
rect 43466 4984 43524 4996
rect 43466 4408 43478 4984
rect 43512 4408 43524 4984
rect 43466 4396 43524 4408
rect 44484 4984 44542 4996
rect 44484 4408 44496 4984
rect 44530 4408 44542 4984
rect 44484 4396 44542 4408
rect 45502 4984 45560 4996
rect 45502 4408 45514 4984
rect 45548 4408 45560 4984
rect 45502 4396 45560 4408
rect 46520 4984 46578 4996
rect 46520 4408 46532 4984
rect 46566 4408 46578 4984
rect 46520 4396 46578 4408
rect 47538 4984 47596 4996
rect 47538 4408 47550 4984
rect 47584 4408 47596 4984
rect 47538 4396 47596 4408
rect 48556 4984 48614 4996
rect 48556 4408 48568 4984
rect 48602 4408 48614 4984
rect 48556 4396 48614 4408
rect 49574 4984 49632 4996
rect 49574 4408 49586 4984
rect 49620 4408 49632 4984
rect 49574 4396 49632 4408
rect 50592 4984 50650 4996
rect 50592 4408 50604 4984
rect 50638 4408 50650 4984
rect 50592 4396 50650 4408
rect 51610 4984 51668 4996
rect 51610 4408 51622 4984
rect 51656 4408 51668 4984
rect 51610 4396 51668 4408
rect 52628 4984 52686 4996
rect 52628 4408 52640 4984
rect 52674 4408 52686 4984
rect 52628 4396 52686 4408
rect 54518 4726 54576 4738
rect 54518 4150 54530 4726
rect 54564 4150 54576 4726
rect 54518 4138 54576 4150
rect 55536 4726 55594 4738
rect 55536 4150 55548 4726
rect 55582 4150 55594 4726
rect 55536 4138 55594 4150
rect 56554 4726 56612 4738
rect 56554 4150 56566 4726
rect 56600 4150 56612 4726
rect 56554 4138 56612 4150
rect 57572 4726 57630 4738
rect 57572 4150 57584 4726
rect 57618 4150 57630 4726
rect 57572 4138 57630 4150
rect 58590 4726 58648 4738
rect 58590 4150 58602 4726
rect 58636 4150 58648 4726
rect 58590 4138 58648 4150
rect 59608 4726 59666 4738
rect 59608 4150 59620 4726
rect 59654 4150 59666 4726
rect 59608 4138 59666 4150
rect 60626 4726 60684 4738
rect 60626 4150 60638 4726
rect 60672 4150 60684 4726
rect 60626 4138 60684 4150
rect 61644 4726 61702 4738
rect 61644 4150 61656 4726
rect 61690 4150 61702 4726
rect 61644 4138 61702 4150
rect 62662 4726 62720 4738
rect 62662 4150 62674 4726
rect 62708 4150 62720 4726
rect 62662 4138 62720 4150
rect 63680 4726 63738 4738
rect 63680 4150 63692 4726
rect 63726 4150 63738 4726
rect 63680 4138 63738 4150
rect 64698 4726 64756 4738
rect 64698 4150 64710 4726
rect 64744 4150 64756 4726
rect 64698 4138 64756 4150
rect 65716 4726 65774 4738
rect 65716 4150 65728 4726
rect 65762 4150 65774 4726
rect 65716 4138 65774 4150
rect 66734 4726 66792 4738
rect 66734 4150 66746 4726
rect 66780 4150 66792 4726
rect 66734 4138 66792 4150
rect 67752 4726 67810 4738
rect 67752 4150 67764 4726
rect 67798 4150 67810 4726
rect 67752 4138 67810 4150
rect 68770 4726 68828 4738
rect 68770 4150 68782 4726
rect 68816 4150 68828 4726
rect 68770 4138 68828 4150
rect 69788 4726 69846 4738
rect 69788 4150 69800 4726
rect 69834 4150 69846 4726
rect 69788 4138 69846 4150
rect 70806 4726 70864 4738
rect 70806 4150 70818 4726
rect 70852 4150 70864 4726
rect 70806 4138 70864 4150
rect 71824 4726 71882 4738
rect 71824 4150 71836 4726
rect 71870 4150 71882 4726
rect 71824 4138 71882 4150
rect 72842 4726 72900 4738
rect 72842 4150 72854 4726
rect 72888 4150 72900 4726
rect 72842 4138 72900 4150
rect 73860 4726 73918 4738
rect 73860 4150 73872 4726
rect 73906 4150 73918 4726
rect 73860 4138 73918 4150
rect 74878 4726 74936 4738
rect 74878 4150 74890 4726
rect 74924 4150 74936 4726
rect 74878 4138 74936 4150
rect 41430 3872 41488 3884
rect 41430 3296 41442 3872
rect 41476 3296 41488 3872
rect 41430 3284 41488 3296
rect 42448 3872 42506 3884
rect 42448 3296 42460 3872
rect 42494 3296 42506 3872
rect 42448 3284 42506 3296
rect 43466 3872 43524 3884
rect 43466 3296 43478 3872
rect 43512 3296 43524 3872
rect 43466 3284 43524 3296
rect 44484 3872 44542 3884
rect 44484 3296 44496 3872
rect 44530 3296 44542 3872
rect 44484 3284 44542 3296
rect 45502 3872 45560 3884
rect 45502 3296 45514 3872
rect 45548 3296 45560 3872
rect 45502 3284 45560 3296
rect 46520 3872 46578 3884
rect 46520 3296 46532 3872
rect 46566 3296 46578 3872
rect 46520 3284 46578 3296
rect 47538 3872 47596 3884
rect 47538 3296 47550 3872
rect 47584 3296 47596 3872
rect 47538 3284 47596 3296
rect 48556 3872 48614 3884
rect 48556 3296 48568 3872
rect 48602 3296 48614 3872
rect 48556 3284 48614 3296
rect 49574 3872 49632 3884
rect 49574 3296 49586 3872
rect 49620 3296 49632 3872
rect 49574 3284 49632 3296
rect 50592 3872 50650 3884
rect 50592 3296 50604 3872
rect 50638 3296 50650 3872
rect 50592 3284 50650 3296
rect 51610 3872 51668 3884
rect 51610 3296 51622 3872
rect 51656 3296 51668 3872
rect 51610 3284 51668 3296
rect 52628 3872 52686 3884
rect 52628 3296 52640 3872
rect 52674 3296 52686 3872
rect 52628 3284 52686 3296
rect 54518 3494 54576 3506
rect 54518 2918 54530 3494
rect 54564 2918 54576 3494
rect 54518 2906 54576 2918
rect 55536 3494 55594 3506
rect 55536 2918 55548 3494
rect 55582 2918 55594 3494
rect 55536 2906 55594 2918
rect 56554 3494 56612 3506
rect 56554 2918 56566 3494
rect 56600 2918 56612 3494
rect 56554 2906 56612 2918
rect 57572 3494 57630 3506
rect 57572 2918 57584 3494
rect 57618 2918 57630 3494
rect 57572 2906 57630 2918
rect 58590 3494 58648 3506
rect 58590 2918 58602 3494
rect 58636 2918 58648 3494
rect 58590 2906 58648 2918
rect 59608 3494 59666 3506
rect 59608 2918 59620 3494
rect 59654 2918 59666 3494
rect 59608 2906 59666 2918
rect 60626 3494 60684 3506
rect 60626 2918 60638 3494
rect 60672 2918 60684 3494
rect 60626 2906 60684 2918
rect 61644 3494 61702 3506
rect 61644 2918 61656 3494
rect 61690 2918 61702 3494
rect 61644 2906 61702 2918
rect 62662 3494 62720 3506
rect 62662 2918 62674 3494
rect 62708 2918 62720 3494
rect 62662 2906 62720 2918
rect 63680 3494 63738 3506
rect 63680 2918 63692 3494
rect 63726 2918 63738 3494
rect 63680 2906 63738 2918
rect 64698 3494 64756 3506
rect 64698 2918 64710 3494
rect 64744 2918 64756 3494
rect 64698 2906 64756 2918
rect 65716 3494 65774 3506
rect 65716 2918 65728 3494
rect 65762 2918 65774 3494
rect 65716 2906 65774 2918
rect 66734 3494 66792 3506
rect 66734 2918 66746 3494
rect 66780 2918 66792 3494
rect 66734 2906 66792 2918
rect 67752 3494 67810 3506
rect 67752 2918 67764 3494
rect 67798 2918 67810 3494
rect 67752 2906 67810 2918
rect 68770 3494 68828 3506
rect 68770 2918 68782 3494
rect 68816 2918 68828 3494
rect 68770 2906 68828 2918
rect 69788 3494 69846 3506
rect 69788 2918 69800 3494
rect 69834 2918 69846 3494
rect 69788 2906 69846 2918
rect 70806 3494 70864 3506
rect 70806 2918 70818 3494
rect 70852 2918 70864 3494
rect 70806 2906 70864 2918
rect 71824 3494 71882 3506
rect 71824 2918 71836 3494
rect 71870 2918 71882 3494
rect 71824 2906 71882 2918
rect 72842 3494 72900 3506
rect 72842 2918 72854 3494
rect 72888 2918 72900 3494
rect 72842 2906 72900 2918
rect 73860 3494 73918 3506
rect 73860 2918 73872 3494
rect 73906 2918 73918 3494
rect 73860 2906 73918 2918
rect 74878 3494 74936 3506
rect 74878 2918 74890 3494
rect 74924 2918 74936 3494
rect 74878 2906 74936 2918
rect 41430 2760 41488 2772
rect 41430 2184 41442 2760
rect 41476 2184 41488 2760
rect 41430 2172 41488 2184
rect 42448 2760 42506 2772
rect 42448 2184 42460 2760
rect 42494 2184 42506 2760
rect 42448 2172 42506 2184
rect 43466 2760 43524 2772
rect 43466 2184 43478 2760
rect 43512 2184 43524 2760
rect 43466 2172 43524 2184
rect 44484 2760 44542 2772
rect 44484 2184 44496 2760
rect 44530 2184 44542 2760
rect 44484 2172 44542 2184
rect 45502 2760 45560 2772
rect 45502 2184 45514 2760
rect 45548 2184 45560 2760
rect 45502 2172 45560 2184
rect 46520 2760 46578 2772
rect 46520 2184 46532 2760
rect 46566 2184 46578 2760
rect 46520 2172 46578 2184
rect 47538 2760 47596 2772
rect 47538 2184 47550 2760
rect 47584 2184 47596 2760
rect 47538 2172 47596 2184
rect 48556 2760 48614 2772
rect 48556 2184 48568 2760
rect 48602 2184 48614 2760
rect 48556 2172 48614 2184
rect 49574 2760 49632 2772
rect 49574 2184 49586 2760
rect 49620 2184 49632 2760
rect 49574 2172 49632 2184
rect 50592 2760 50650 2772
rect 50592 2184 50604 2760
rect 50638 2184 50650 2760
rect 50592 2172 50650 2184
rect 51610 2760 51668 2772
rect 51610 2184 51622 2760
rect 51656 2184 51668 2760
rect 51610 2172 51668 2184
rect 52628 2760 52686 2772
rect 52628 2184 52640 2760
rect 52674 2184 52686 2760
rect 52628 2172 52686 2184
rect 54518 2260 54576 2272
rect 54518 1684 54530 2260
rect 54564 1684 54576 2260
rect 54518 1672 54576 1684
rect 55536 2260 55594 2272
rect 55536 1684 55548 2260
rect 55582 1684 55594 2260
rect 55536 1672 55594 1684
rect 56554 2260 56612 2272
rect 56554 1684 56566 2260
rect 56600 1684 56612 2260
rect 56554 1672 56612 1684
rect 57572 2260 57630 2272
rect 57572 1684 57584 2260
rect 57618 1684 57630 2260
rect 57572 1672 57630 1684
rect 58590 2260 58648 2272
rect 58590 1684 58602 2260
rect 58636 1684 58648 2260
rect 58590 1672 58648 1684
rect 59608 2260 59666 2272
rect 59608 1684 59620 2260
rect 59654 1684 59666 2260
rect 59608 1672 59666 1684
rect 60626 2260 60684 2272
rect 60626 1684 60638 2260
rect 60672 1684 60684 2260
rect 60626 1672 60684 1684
rect 61644 2260 61702 2272
rect 61644 1684 61656 2260
rect 61690 1684 61702 2260
rect 61644 1672 61702 1684
rect 62662 2260 62720 2272
rect 62662 1684 62674 2260
rect 62708 1684 62720 2260
rect 62662 1672 62720 1684
rect 63680 2260 63738 2272
rect 63680 1684 63692 2260
rect 63726 1684 63738 2260
rect 63680 1672 63738 1684
rect 64698 2260 64756 2272
rect 64698 1684 64710 2260
rect 64744 1684 64756 2260
rect 64698 1672 64756 1684
rect 65716 2260 65774 2272
rect 65716 1684 65728 2260
rect 65762 1684 65774 2260
rect 65716 1672 65774 1684
rect 66734 2260 66792 2272
rect 66734 1684 66746 2260
rect 66780 1684 66792 2260
rect 66734 1672 66792 1684
rect 67752 2260 67810 2272
rect 67752 1684 67764 2260
rect 67798 1684 67810 2260
rect 67752 1672 67810 1684
rect 68770 2260 68828 2272
rect 68770 1684 68782 2260
rect 68816 1684 68828 2260
rect 68770 1672 68828 1684
rect 69788 2260 69846 2272
rect 69788 1684 69800 2260
rect 69834 1684 69846 2260
rect 69788 1672 69846 1684
rect 70806 2260 70864 2272
rect 70806 1684 70818 2260
rect 70852 1684 70864 2260
rect 70806 1672 70864 1684
rect 71824 2260 71882 2272
rect 71824 1684 71836 2260
rect 71870 1684 71882 2260
rect 71824 1672 71882 1684
rect 72842 2260 72900 2272
rect 72842 1684 72854 2260
rect 72888 1684 72900 2260
rect 72842 1672 72900 1684
rect 73860 2260 73918 2272
rect 73860 1684 73872 2260
rect 73906 1684 73918 2260
rect 73860 1672 73918 1684
rect 74878 2260 74936 2272
rect 74878 1684 74890 2260
rect 74924 1684 74936 2260
rect 74878 1672 74936 1684
rect 41888 1218 41946 1230
rect 41888 642 41900 1218
rect 41934 642 41946 1218
rect 41888 630 41946 642
rect 42906 1218 42964 1230
rect 42906 642 42918 1218
rect 42952 642 42964 1218
rect 42906 630 42964 642
rect 43924 1218 43982 1230
rect 43924 642 43936 1218
rect 43970 642 43982 1218
rect 43924 630 43982 642
rect 44942 1218 45000 1230
rect 44942 642 44954 1218
rect 44988 642 45000 1218
rect 44942 630 45000 642
rect 45960 1218 46018 1230
rect 45960 642 45972 1218
rect 46006 642 46018 1218
rect 45960 630 46018 642
rect 46978 1218 47036 1230
rect 46978 642 46990 1218
rect 47024 642 47036 1218
rect 46978 630 47036 642
rect 47996 1218 48054 1230
rect 47996 642 48008 1218
rect 48042 642 48054 1218
rect 47996 630 48054 642
rect 49014 1218 49072 1230
rect 49014 642 49026 1218
rect 49060 642 49072 1218
rect 49014 630 49072 642
rect 50032 1218 50090 1230
rect 50032 642 50044 1218
rect 50078 642 50090 1218
rect 50032 630 50090 642
rect 51050 1218 51108 1230
rect 51050 642 51062 1218
rect 51096 642 51108 1218
rect 51050 630 51108 642
rect 52068 1218 52126 1230
rect 52068 642 52080 1218
rect 52114 642 52126 1218
rect 52068 630 52126 642
rect 54518 1028 54576 1040
rect 54518 452 54530 1028
rect 54564 452 54576 1028
rect 54518 440 54576 452
rect 55536 1028 55594 1040
rect 55536 452 55548 1028
rect 55582 452 55594 1028
rect 55536 440 55594 452
rect 56554 1028 56612 1040
rect 56554 452 56566 1028
rect 56600 452 56612 1028
rect 56554 440 56612 452
rect 57572 1028 57630 1040
rect 57572 452 57584 1028
rect 57618 452 57630 1028
rect 57572 440 57630 452
rect 58590 1028 58648 1040
rect 58590 452 58602 1028
rect 58636 452 58648 1028
rect 58590 440 58648 452
rect 59608 1028 59666 1040
rect 59608 452 59620 1028
rect 59654 452 59666 1028
rect 59608 440 59666 452
rect 60626 1028 60684 1040
rect 60626 452 60638 1028
rect 60672 452 60684 1028
rect 60626 440 60684 452
rect 61644 1028 61702 1040
rect 61644 452 61656 1028
rect 61690 452 61702 1028
rect 61644 440 61702 452
rect 62662 1028 62720 1040
rect 62662 452 62674 1028
rect 62708 452 62720 1028
rect 62662 440 62720 452
rect 63680 1028 63738 1040
rect 63680 452 63692 1028
rect 63726 452 63738 1028
rect 63680 440 63738 452
rect 64698 1028 64756 1040
rect 64698 452 64710 1028
rect 64744 452 64756 1028
rect 64698 440 64756 452
rect 65716 1028 65774 1040
rect 65716 452 65728 1028
rect 65762 452 65774 1028
rect 65716 440 65774 452
rect 66734 1028 66792 1040
rect 66734 452 66746 1028
rect 66780 452 66792 1028
rect 66734 440 66792 452
rect 67752 1028 67810 1040
rect 67752 452 67764 1028
rect 67798 452 67810 1028
rect 67752 440 67810 452
rect 68770 1028 68828 1040
rect 68770 452 68782 1028
rect 68816 452 68828 1028
rect 68770 440 68828 452
rect 69788 1028 69846 1040
rect 69788 452 69800 1028
rect 69834 452 69846 1028
rect 69788 440 69846 452
rect 70806 1028 70864 1040
rect 70806 452 70818 1028
rect 70852 452 70864 1028
rect 70806 440 70864 452
rect 71824 1028 71882 1040
rect 71824 452 71836 1028
rect 71870 452 71882 1028
rect 71824 440 71882 452
rect 72842 1028 72900 1040
rect 72842 452 72854 1028
rect 72888 452 72900 1028
rect 72842 440 72900 452
rect 73860 1028 73918 1040
rect 73860 452 73872 1028
rect 73906 452 73918 1028
rect 73860 440 73918 452
rect 74878 1028 74936 1040
rect 74878 452 74890 1028
rect 74924 452 74936 1028
rect 74878 440 74936 452
<< pdiff >>
rect 17426 27832 17484 27844
rect 17426 27256 17438 27832
rect 17472 27256 17484 27832
rect 17426 27244 17484 27256
rect 18444 27832 18502 27844
rect 18444 27256 18456 27832
rect 18490 27256 18502 27832
rect 18444 27244 18502 27256
rect 19462 27832 19520 27844
rect 19462 27256 19474 27832
rect 19508 27256 19520 27832
rect 19462 27244 19520 27256
rect 20480 27832 20538 27844
rect 20480 27256 20492 27832
rect 20526 27256 20538 27832
rect 20480 27244 20538 27256
rect 21498 27832 21556 27844
rect 21498 27256 21510 27832
rect 21544 27256 21556 27832
rect 21498 27244 21556 27256
rect 22516 27832 22574 27844
rect 22516 27256 22528 27832
rect 22562 27256 22574 27832
rect 22516 27244 22574 27256
rect 23534 27832 23592 27844
rect 23534 27256 23546 27832
rect 23580 27256 23592 27832
rect 23534 27244 23592 27256
rect 24552 27832 24610 27844
rect 24552 27256 24564 27832
rect 24598 27256 24610 27832
rect 24552 27244 24610 27256
rect 25570 27832 25628 27844
rect 25570 27256 25582 27832
rect 25616 27256 25628 27832
rect 25570 27244 25628 27256
rect 26588 27832 26646 27844
rect 26588 27256 26600 27832
rect 26634 27256 26646 27832
rect 26588 27244 26646 27256
rect 27606 27832 27664 27844
rect 27606 27256 27618 27832
rect 27652 27256 27664 27832
rect 27606 27244 27664 27256
rect 28624 27832 28682 27844
rect 28624 27256 28636 27832
rect 28670 27256 28682 27832
rect 28624 27244 28682 27256
rect 29642 27832 29700 27844
rect 29642 27256 29654 27832
rect 29688 27256 29700 27832
rect 29642 27244 29700 27256
rect 30660 27832 30718 27844
rect 30660 27256 30672 27832
rect 30706 27256 30718 27832
rect 30660 27244 30718 27256
rect 31678 27832 31736 27844
rect 31678 27256 31690 27832
rect 31724 27256 31736 27832
rect 31678 27244 31736 27256
rect 32696 27832 32754 27844
rect 32696 27256 32708 27832
rect 32742 27256 32754 27832
rect 32696 27244 32754 27256
rect 33714 27832 33772 27844
rect 33714 27256 33726 27832
rect 33760 27256 33772 27832
rect 33714 27244 33772 27256
rect 17426 26696 17484 26708
rect 17426 26120 17438 26696
rect 17472 26120 17484 26696
rect 17426 26108 17484 26120
rect 18444 26696 18502 26708
rect 18444 26120 18456 26696
rect 18490 26120 18502 26696
rect 18444 26108 18502 26120
rect 19462 26696 19520 26708
rect 19462 26120 19474 26696
rect 19508 26120 19520 26696
rect 19462 26108 19520 26120
rect 20480 26696 20538 26708
rect 20480 26120 20492 26696
rect 20526 26120 20538 26696
rect 20480 26108 20538 26120
rect 21498 26696 21556 26708
rect 21498 26120 21510 26696
rect 21544 26120 21556 26696
rect 21498 26108 21556 26120
rect 22516 26696 22574 26708
rect 22516 26120 22528 26696
rect 22562 26120 22574 26696
rect 22516 26108 22574 26120
rect 23534 26696 23592 26708
rect 23534 26120 23546 26696
rect 23580 26120 23592 26696
rect 23534 26108 23592 26120
rect 24552 26696 24610 26708
rect 24552 26120 24564 26696
rect 24598 26120 24610 26696
rect 24552 26108 24610 26120
rect 25570 26696 25628 26708
rect 25570 26120 25582 26696
rect 25616 26120 25628 26696
rect 25570 26108 25628 26120
rect 26588 26696 26646 26708
rect 26588 26120 26600 26696
rect 26634 26120 26646 26696
rect 26588 26108 26646 26120
rect 27606 26696 27664 26708
rect 27606 26120 27618 26696
rect 27652 26120 27664 26696
rect 27606 26108 27664 26120
rect 28624 26696 28682 26708
rect 28624 26120 28636 26696
rect 28670 26120 28682 26696
rect 28624 26108 28682 26120
rect 29642 26696 29700 26708
rect 29642 26120 29654 26696
rect 29688 26120 29700 26696
rect 29642 26108 29700 26120
rect 30660 26696 30718 26708
rect 30660 26120 30672 26696
rect 30706 26120 30718 26696
rect 30660 26108 30718 26120
rect 31678 26696 31736 26708
rect 31678 26120 31690 26696
rect 31724 26120 31736 26696
rect 31678 26108 31736 26120
rect 32696 26696 32754 26708
rect 32696 26120 32708 26696
rect 32742 26120 32754 26696
rect 32696 26108 32754 26120
rect 33714 26696 33772 26708
rect 33714 26120 33726 26696
rect 33760 26120 33772 26696
rect 33714 26108 33772 26120
rect 17426 25560 17484 25572
rect 17426 24984 17438 25560
rect 17472 24984 17484 25560
rect 17426 24972 17484 24984
rect 18444 25560 18502 25572
rect 18444 24984 18456 25560
rect 18490 24984 18502 25560
rect 18444 24972 18502 24984
rect 19462 25560 19520 25572
rect 19462 24984 19474 25560
rect 19508 24984 19520 25560
rect 19462 24972 19520 24984
rect 20480 25560 20538 25572
rect 20480 24984 20492 25560
rect 20526 24984 20538 25560
rect 20480 24972 20538 24984
rect 21498 25560 21556 25572
rect 21498 24984 21510 25560
rect 21544 24984 21556 25560
rect 21498 24972 21556 24984
rect 22516 25560 22574 25572
rect 22516 24984 22528 25560
rect 22562 24984 22574 25560
rect 22516 24972 22574 24984
rect 23534 25560 23592 25572
rect 23534 24984 23546 25560
rect 23580 24984 23592 25560
rect 23534 24972 23592 24984
rect 24552 25560 24610 25572
rect 24552 24984 24564 25560
rect 24598 24984 24610 25560
rect 24552 24972 24610 24984
rect 25570 25560 25628 25572
rect 25570 24984 25582 25560
rect 25616 24984 25628 25560
rect 25570 24972 25628 24984
rect 26588 25560 26646 25572
rect 26588 24984 26600 25560
rect 26634 24984 26646 25560
rect 26588 24972 26646 24984
rect 27606 25560 27664 25572
rect 27606 24984 27618 25560
rect 27652 24984 27664 25560
rect 27606 24972 27664 24984
rect 28624 25560 28682 25572
rect 28624 24984 28636 25560
rect 28670 24984 28682 25560
rect 28624 24972 28682 24984
rect 29642 25560 29700 25572
rect 29642 24984 29654 25560
rect 29688 24984 29700 25560
rect 29642 24972 29700 24984
rect 30660 25560 30718 25572
rect 30660 24984 30672 25560
rect 30706 24984 30718 25560
rect 30660 24972 30718 24984
rect 31678 25560 31736 25572
rect 31678 24984 31690 25560
rect 31724 24984 31736 25560
rect 31678 24972 31736 24984
rect 32696 25560 32754 25572
rect 32696 24984 32708 25560
rect 32742 24984 32754 25560
rect 32696 24972 32754 24984
rect 33714 25560 33772 25572
rect 33714 24984 33726 25560
rect 33760 24984 33772 25560
rect 33714 24972 33772 24984
rect 18620 23922 18678 23934
rect 18620 23346 18632 23922
rect 18666 23346 18678 23922
rect 18620 23334 18678 23346
rect 19638 23922 19696 23934
rect 19638 23346 19650 23922
rect 19684 23346 19696 23922
rect 19638 23334 19696 23346
rect 20656 23922 20714 23934
rect 20656 23346 20668 23922
rect 20702 23346 20714 23922
rect 20656 23334 20714 23346
rect 21674 23922 21732 23934
rect 21674 23346 21686 23922
rect 21720 23346 21732 23922
rect 21674 23334 21732 23346
rect 22692 23922 22750 23934
rect 22692 23346 22704 23922
rect 22738 23346 22750 23922
rect 22692 23334 22750 23346
rect 23710 23922 23768 23934
rect 23710 23346 23722 23922
rect 23756 23346 23768 23922
rect 23710 23334 23768 23346
rect 24728 23922 24786 23934
rect 24728 23346 24740 23922
rect 24774 23346 24786 23922
rect 24728 23334 24786 23346
rect 25746 23922 25804 23934
rect 25746 23346 25758 23922
rect 25792 23346 25804 23922
rect 25746 23334 25804 23346
rect 26764 23922 26822 23934
rect 26764 23346 26776 23922
rect 26810 23346 26822 23922
rect 26764 23334 26822 23346
rect 27782 23922 27840 23934
rect 27782 23346 27794 23922
rect 27828 23346 27840 23922
rect 27782 23334 27840 23346
rect 28800 23922 28858 23934
rect 28800 23346 28812 23922
rect 28846 23346 28858 23922
rect 28800 23334 28858 23346
rect 29818 23922 29876 23934
rect 29818 23346 29830 23922
rect 29864 23346 29876 23922
rect 29818 23334 29876 23346
rect 30836 23922 30894 23934
rect 30836 23346 30848 23922
rect 30882 23346 30894 23922
rect 30836 23334 30894 23346
rect 31854 23922 31912 23934
rect 31854 23346 31866 23922
rect 31900 23346 31912 23922
rect 31854 23334 31912 23346
rect 32872 23922 32930 23934
rect 32872 23346 32884 23922
rect 32918 23346 32930 23922
rect 32872 23334 32930 23346
rect 18620 22890 18678 22902
rect 18620 22314 18632 22890
rect 18666 22314 18678 22890
rect 18620 22302 18678 22314
rect 19638 22890 19696 22902
rect 19638 22314 19650 22890
rect 19684 22314 19696 22890
rect 19638 22302 19696 22314
rect 20656 22890 20714 22902
rect 20656 22314 20668 22890
rect 20702 22314 20714 22890
rect 20656 22302 20714 22314
rect 21674 22890 21732 22902
rect 21674 22314 21686 22890
rect 21720 22314 21732 22890
rect 21674 22302 21732 22314
rect 22692 22890 22750 22902
rect 22692 22314 22704 22890
rect 22738 22314 22750 22890
rect 22692 22302 22750 22314
rect 23710 22890 23768 22902
rect 23710 22314 23722 22890
rect 23756 22314 23768 22890
rect 23710 22302 23768 22314
rect 24728 22890 24786 22902
rect 24728 22314 24740 22890
rect 24774 22314 24786 22890
rect 24728 22302 24786 22314
rect 25746 22890 25804 22902
rect 25746 22314 25758 22890
rect 25792 22314 25804 22890
rect 25746 22302 25804 22314
rect 26764 22890 26822 22902
rect 26764 22314 26776 22890
rect 26810 22314 26822 22890
rect 26764 22302 26822 22314
rect 27782 22890 27840 22902
rect 27782 22314 27794 22890
rect 27828 22314 27840 22890
rect 27782 22302 27840 22314
rect 28800 22890 28858 22902
rect 28800 22314 28812 22890
rect 28846 22314 28858 22890
rect 28800 22302 28858 22314
rect 29818 22890 29876 22902
rect 29818 22314 29830 22890
rect 29864 22314 29876 22890
rect 29818 22302 29876 22314
rect 30836 22890 30894 22902
rect 30836 22314 30848 22890
rect 30882 22314 30894 22890
rect 30836 22302 30894 22314
rect 31854 22890 31912 22902
rect 31854 22314 31866 22890
rect 31900 22314 31912 22890
rect 31854 22302 31912 22314
rect 32872 22890 32930 22902
rect 32872 22314 32884 22890
rect 32918 22314 32930 22890
rect 32872 22302 32930 22314
rect 18412 21286 18470 21298
rect 13108 21182 13166 21194
rect 13108 20606 13120 21182
rect 13154 20606 13166 21182
rect 13108 20594 13166 20606
rect 14126 21182 14184 21194
rect 14126 20606 14138 21182
rect 14172 20606 14184 21182
rect 14126 20594 14184 20606
rect 15144 21182 15202 21194
rect 15144 20606 15156 21182
rect 15190 20606 15202 21182
rect 15144 20594 15202 20606
rect 16162 21182 16220 21194
rect 16162 20606 16174 21182
rect 16208 20606 16220 21182
rect 16162 20594 16220 20606
rect 17180 21182 17238 21194
rect 17180 20606 17192 21182
rect 17226 20606 17238 21182
rect 18412 20710 18424 21286
rect 18458 20710 18470 21286
rect 18412 20698 18470 20710
rect 19430 21286 19488 21298
rect 19430 20710 19442 21286
rect 19476 20710 19488 21286
rect 19430 20698 19488 20710
rect 20448 21286 20506 21298
rect 20448 20710 20460 21286
rect 20494 20710 20506 21286
rect 20448 20698 20506 20710
rect 21466 21286 21524 21298
rect 21466 20710 21478 21286
rect 21512 20710 21524 21286
rect 21466 20698 21524 20710
rect 22484 21286 22542 21298
rect 22484 20710 22496 21286
rect 22530 20710 22542 21286
rect 22484 20698 22542 20710
rect 23502 21286 23560 21298
rect 23502 20710 23514 21286
rect 23548 20710 23560 21286
rect 23502 20698 23560 20710
rect 24520 21286 24578 21298
rect 24520 20710 24532 21286
rect 24566 20710 24578 21286
rect 24520 20698 24578 20710
rect 25538 21286 25596 21298
rect 25538 20710 25550 21286
rect 25584 20710 25596 21286
rect 25538 20698 25596 20710
rect 26556 21286 26614 21298
rect 26556 20710 26568 21286
rect 26602 20710 26614 21286
rect 26556 20698 26614 20710
rect 27574 21286 27632 21298
rect 27574 20710 27586 21286
rect 27620 20710 27632 21286
rect 27574 20698 27632 20710
rect 28592 21286 28650 21298
rect 28592 20710 28604 21286
rect 28638 20710 28650 21286
rect 28592 20698 28650 20710
rect 29610 21286 29668 21298
rect 29610 20710 29622 21286
rect 29656 20710 29668 21286
rect 29610 20698 29668 20710
rect 30628 21286 30686 21298
rect 30628 20710 30640 21286
rect 30674 20710 30686 21286
rect 30628 20698 30686 20710
rect 31646 21286 31704 21298
rect 31646 20710 31658 21286
rect 31692 20710 31704 21286
rect 31646 20698 31704 20710
rect 32664 21286 32722 21298
rect 32664 20710 32676 21286
rect 32710 20710 32722 21286
rect 32664 20698 32722 20710
rect 33682 21286 33740 21298
rect 33682 20710 33694 21286
rect 33728 20710 33740 21286
rect 33682 20698 33740 20710
rect 17180 20594 17238 20606
rect 13108 20150 13166 20162
rect 13108 19574 13120 20150
rect 13154 19574 13166 20150
rect 13108 19562 13166 19574
rect 14126 20150 14184 20162
rect 14126 19574 14138 20150
rect 14172 19574 14184 20150
rect 14126 19562 14184 19574
rect 15144 20150 15202 20162
rect 15144 19574 15156 20150
rect 15190 19574 15202 20150
rect 15144 19562 15202 19574
rect 16162 20150 16220 20162
rect 16162 19574 16174 20150
rect 16208 19574 16220 20150
rect 16162 19562 16220 19574
rect 17180 20150 17238 20162
rect 17180 19574 17192 20150
rect 17226 19574 17238 20150
rect 17180 19562 17238 19574
rect 18412 20030 18470 20042
rect 18412 19454 18424 20030
rect 18458 19454 18470 20030
rect 18412 19442 18470 19454
rect 19430 20030 19488 20042
rect 19430 19454 19442 20030
rect 19476 19454 19488 20030
rect 19430 19442 19488 19454
rect 20448 20030 20506 20042
rect 20448 19454 20460 20030
rect 20494 19454 20506 20030
rect 20448 19442 20506 19454
rect 21466 20030 21524 20042
rect 21466 19454 21478 20030
rect 21512 19454 21524 20030
rect 21466 19442 21524 19454
rect 22484 20030 22542 20042
rect 22484 19454 22496 20030
rect 22530 19454 22542 20030
rect 22484 19442 22542 19454
rect 23502 20030 23560 20042
rect 23502 19454 23514 20030
rect 23548 19454 23560 20030
rect 23502 19442 23560 19454
rect 24520 20030 24578 20042
rect 24520 19454 24532 20030
rect 24566 19454 24578 20030
rect 24520 19442 24578 19454
rect 25538 20030 25596 20042
rect 25538 19454 25550 20030
rect 25584 19454 25596 20030
rect 25538 19442 25596 19454
rect 26556 20030 26614 20042
rect 26556 19454 26568 20030
rect 26602 19454 26614 20030
rect 26556 19442 26614 19454
rect 27574 20030 27632 20042
rect 27574 19454 27586 20030
rect 27620 19454 27632 20030
rect 27574 19442 27632 19454
rect 28592 20030 28650 20042
rect 28592 19454 28604 20030
rect 28638 19454 28650 20030
rect 28592 19442 28650 19454
rect 29610 20030 29668 20042
rect 29610 19454 29622 20030
rect 29656 19454 29668 20030
rect 29610 19442 29668 19454
rect 30628 20030 30686 20042
rect 30628 19454 30640 20030
rect 30674 19454 30686 20030
rect 30628 19442 30686 19454
rect 31646 20030 31704 20042
rect 31646 19454 31658 20030
rect 31692 19454 31704 20030
rect 31646 19442 31704 19454
rect 32664 20030 32722 20042
rect 32664 19454 32676 20030
rect 32710 19454 32722 20030
rect 32664 19442 32722 19454
rect 33682 20030 33740 20042
rect 33682 19454 33694 20030
rect 33728 19454 33740 20030
rect 33682 19442 33740 19454
rect 13108 19118 13166 19130
rect 13108 18542 13120 19118
rect 13154 18542 13166 19118
rect 13108 18530 13166 18542
rect 14126 19118 14184 19130
rect 14126 18542 14138 19118
rect 14172 18542 14184 19118
rect 14126 18530 14184 18542
rect 15144 19118 15202 19130
rect 15144 18542 15156 19118
rect 15190 18542 15202 19118
rect 15144 18530 15202 18542
rect 16162 19118 16220 19130
rect 16162 18542 16174 19118
rect 16208 18542 16220 19118
rect 16162 18530 16220 18542
rect 17180 19118 17238 19130
rect 17180 18542 17192 19118
rect 17226 18542 17238 19118
rect 17180 18530 17238 18542
rect 18412 18774 18470 18786
rect 18412 18198 18424 18774
rect 18458 18198 18470 18774
rect 18412 18186 18470 18198
rect 19430 18774 19488 18786
rect 19430 18198 19442 18774
rect 19476 18198 19488 18774
rect 19430 18186 19488 18198
rect 20448 18774 20506 18786
rect 20448 18198 20460 18774
rect 20494 18198 20506 18774
rect 20448 18186 20506 18198
rect 21466 18774 21524 18786
rect 21466 18198 21478 18774
rect 21512 18198 21524 18774
rect 21466 18186 21524 18198
rect 22484 18774 22542 18786
rect 22484 18198 22496 18774
rect 22530 18198 22542 18774
rect 22484 18186 22542 18198
rect 23502 18774 23560 18786
rect 23502 18198 23514 18774
rect 23548 18198 23560 18774
rect 23502 18186 23560 18198
rect 24520 18774 24578 18786
rect 24520 18198 24532 18774
rect 24566 18198 24578 18774
rect 24520 18186 24578 18198
rect 25538 18774 25596 18786
rect 25538 18198 25550 18774
rect 25584 18198 25596 18774
rect 25538 18186 25596 18198
rect 26556 18774 26614 18786
rect 26556 18198 26568 18774
rect 26602 18198 26614 18774
rect 26556 18186 26614 18198
rect 27574 18774 27632 18786
rect 27574 18198 27586 18774
rect 27620 18198 27632 18774
rect 27574 18186 27632 18198
rect 28592 18774 28650 18786
rect 28592 18198 28604 18774
rect 28638 18198 28650 18774
rect 28592 18186 28650 18198
rect 29610 18774 29668 18786
rect 29610 18198 29622 18774
rect 29656 18198 29668 18774
rect 29610 18186 29668 18198
rect 30628 18774 30686 18786
rect 30628 18198 30640 18774
rect 30674 18198 30686 18774
rect 30628 18186 30686 18198
rect 31646 18774 31704 18786
rect 31646 18198 31658 18774
rect 31692 18198 31704 18774
rect 31646 18186 31704 18198
rect 32664 18774 32722 18786
rect 32664 18198 32676 18774
rect 32710 18198 32722 18774
rect 32664 18186 32722 18198
rect 33682 18774 33740 18786
rect 33682 18198 33694 18774
rect 33728 18198 33740 18774
rect 33682 18186 33740 18198
rect 13108 18086 13166 18098
rect 13108 17510 13120 18086
rect 13154 17510 13166 18086
rect 13108 17498 13166 17510
rect 14126 18086 14184 18098
rect 14126 17510 14138 18086
rect 14172 17510 14184 18086
rect 14126 17498 14184 17510
rect 15144 18086 15202 18098
rect 15144 17510 15156 18086
rect 15190 17510 15202 18086
rect 15144 17498 15202 17510
rect 16162 18086 16220 18098
rect 16162 17510 16174 18086
rect 16208 17510 16220 18086
rect 16162 17498 16220 17510
rect 17180 18086 17238 18098
rect 17180 17510 17192 18086
rect 17226 17510 17238 18086
rect 17180 17498 17238 17510
rect 18412 17518 18470 17530
rect 18412 16942 18424 17518
rect 18458 16942 18470 17518
rect 18412 16930 18470 16942
rect 19430 17518 19488 17530
rect 19430 16942 19442 17518
rect 19476 16942 19488 17518
rect 19430 16930 19488 16942
rect 20448 17518 20506 17530
rect 20448 16942 20460 17518
rect 20494 16942 20506 17518
rect 20448 16930 20506 16942
rect 21466 17518 21524 17530
rect 21466 16942 21478 17518
rect 21512 16942 21524 17518
rect 21466 16930 21524 16942
rect 22484 17518 22542 17530
rect 22484 16942 22496 17518
rect 22530 16942 22542 17518
rect 22484 16930 22542 16942
rect 23502 17518 23560 17530
rect 23502 16942 23514 17518
rect 23548 16942 23560 17518
rect 23502 16930 23560 16942
rect 24520 17518 24578 17530
rect 24520 16942 24532 17518
rect 24566 16942 24578 17518
rect 24520 16930 24578 16942
rect 25538 17518 25596 17530
rect 25538 16942 25550 17518
rect 25584 16942 25596 17518
rect 25538 16930 25596 16942
rect 26556 17518 26614 17530
rect 26556 16942 26568 17518
rect 26602 16942 26614 17518
rect 26556 16930 26614 16942
rect 27574 17518 27632 17530
rect 27574 16942 27586 17518
rect 27620 16942 27632 17518
rect 27574 16930 27632 16942
rect 28592 17518 28650 17530
rect 28592 16942 28604 17518
rect 28638 16942 28650 17518
rect 28592 16930 28650 16942
rect 29610 17518 29668 17530
rect 29610 16942 29622 17518
rect 29656 16942 29668 17518
rect 29610 16930 29668 16942
rect 30628 17518 30686 17530
rect 30628 16942 30640 17518
rect 30674 16942 30686 17518
rect 30628 16930 30686 16942
rect 31646 17518 31704 17530
rect 31646 16942 31658 17518
rect 31692 16942 31704 17518
rect 31646 16930 31704 16942
rect 32664 17518 32722 17530
rect 32664 16942 32676 17518
rect 32710 16942 32722 17518
rect 32664 16930 32722 16942
rect 33682 17518 33740 17530
rect 33682 16942 33694 17518
rect 33728 16942 33740 17518
rect 33682 16930 33740 16942
rect 58426 27832 58484 27844
rect 58426 27256 58438 27832
rect 58472 27256 58484 27832
rect 58426 27244 58484 27256
rect 59444 27832 59502 27844
rect 59444 27256 59456 27832
rect 59490 27256 59502 27832
rect 59444 27244 59502 27256
rect 60462 27832 60520 27844
rect 60462 27256 60474 27832
rect 60508 27256 60520 27832
rect 60462 27244 60520 27256
rect 61480 27832 61538 27844
rect 61480 27256 61492 27832
rect 61526 27256 61538 27832
rect 61480 27244 61538 27256
rect 62498 27832 62556 27844
rect 62498 27256 62510 27832
rect 62544 27256 62556 27832
rect 62498 27244 62556 27256
rect 63516 27832 63574 27844
rect 63516 27256 63528 27832
rect 63562 27256 63574 27832
rect 63516 27244 63574 27256
rect 64534 27832 64592 27844
rect 64534 27256 64546 27832
rect 64580 27256 64592 27832
rect 64534 27244 64592 27256
rect 65552 27832 65610 27844
rect 65552 27256 65564 27832
rect 65598 27256 65610 27832
rect 65552 27244 65610 27256
rect 66570 27832 66628 27844
rect 66570 27256 66582 27832
rect 66616 27256 66628 27832
rect 66570 27244 66628 27256
rect 67588 27832 67646 27844
rect 67588 27256 67600 27832
rect 67634 27256 67646 27832
rect 67588 27244 67646 27256
rect 68606 27832 68664 27844
rect 68606 27256 68618 27832
rect 68652 27256 68664 27832
rect 68606 27244 68664 27256
rect 69624 27832 69682 27844
rect 69624 27256 69636 27832
rect 69670 27256 69682 27832
rect 69624 27244 69682 27256
rect 70642 27832 70700 27844
rect 70642 27256 70654 27832
rect 70688 27256 70700 27832
rect 70642 27244 70700 27256
rect 71660 27832 71718 27844
rect 71660 27256 71672 27832
rect 71706 27256 71718 27832
rect 71660 27244 71718 27256
rect 72678 27832 72736 27844
rect 72678 27256 72690 27832
rect 72724 27256 72736 27832
rect 72678 27244 72736 27256
rect 73696 27832 73754 27844
rect 73696 27256 73708 27832
rect 73742 27256 73754 27832
rect 73696 27244 73754 27256
rect 74714 27832 74772 27844
rect 74714 27256 74726 27832
rect 74760 27256 74772 27832
rect 74714 27244 74772 27256
rect 58426 26696 58484 26708
rect 58426 26120 58438 26696
rect 58472 26120 58484 26696
rect 58426 26108 58484 26120
rect 59444 26696 59502 26708
rect 59444 26120 59456 26696
rect 59490 26120 59502 26696
rect 59444 26108 59502 26120
rect 60462 26696 60520 26708
rect 60462 26120 60474 26696
rect 60508 26120 60520 26696
rect 60462 26108 60520 26120
rect 61480 26696 61538 26708
rect 61480 26120 61492 26696
rect 61526 26120 61538 26696
rect 61480 26108 61538 26120
rect 62498 26696 62556 26708
rect 62498 26120 62510 26696
rect 62544 26120 62556 26696
rect 62498 26108 62556 26120
rect 63516 26696 63574 26708
rect 63516 26120 63528 26696
rect 63562 26120 63574 26696
rect 63516 26108 63574 26120
rect 64534 26696 64592 26708
rect 64534 26120 64546 26696
rect 64580 26120 64592 26696
rect 64534 26108 64592 26120
rect 65552 26696 65610 26708
rect 65552 26120 65564 26696
rect 65598 26120 65610 26696
rect 65552 26108 65610 26120
rect 66570 26696 66628 26708
rect 66570 26120 66582 26696
rect 66616 26120 66628 26696
rect 66570 26108 66628 26120
rect 67588 26696 67646 26708
rect 67588 26120 67600 26696
rect 67634 26120 67646 26696
rect 67588 26108 67646 26120
rect 68606 26696 68664 26708
rect 68606 26120 68618 26696
rect 68652 26120 68664 26696
rect 68606 26108 68664 26120
rect 69624 26696 69682 26708
rect 69624 26120 69636 26696
rect 69670 26120 69682 26696
rect 69624 26108 69682 26120
rect 70642 26696 70700 26708
rect 70642 26120 70654 26696
rect 70688 26120 70700 26696
rect 70642 26108 70700 26120
rect 71660 26696 71718 26708
rect 71660 26120 71672 26696
rect 71706 26120 71718 26696
rect 71660 26108 71718 26120
rect 72678 26696 72736 26708
rect 72678 26120 72690 26696
rect 72724 26120 72736 26696
rect 72678 26108 72736 26120
rect 73696 26696 73754 26708
rect 73696 26120 73708 26696
rect 73742 26120 73754 26696
rect 73696 26108 73754 26120
rect 74714 26696 74772 26708
rect 74714 26120 74726 26696
rect 74760 26120 74772 26696
rect 74714 26108 74772 26120
rect 58426 25560 58484 25572
rect 58426 24984 58438 25560
rect 58472 24984 58484 25560
rect 58426 24972 58484 24984
rect 59444 25560 59502 25572
rect 59444 24984 59456 25560
rect 59490 24984 59502 25560
rect 59444 24972 59502 24984
rect 60462 25560 60520 25572
rect 60462 24984 60474 25560
rect 60508 24984 60520 25560
rect 60462 24972 60520 24984
rect 61480 25560 61538 25572
rect 61480 24984 61492 25560
rect 61526 24984 61538 25560
rect 61480 24972 61538 24984
rect 62498 25560 62556 25572
rect 62498 24984 62510 25560
rect 62544 24984 62556 25560
rect 62498 24972 62556 24984
rect 63516 25560 63574 25572
rect 63516 24984 63528 25560
rect 63562 24984 63574 25560
rect 63516 24972 63574 24984
rect 64534 25560 64592 25572
rect 64534 24984 64546 25560
rect 64580 24984 64592 25560
rect 64534 24972 64592 24984
rect 65552 25560 65610 25572
rect 65552 24984 65564 25560
rect 65598 24984 65610 25560
rect 65552 24972 65610 24984
rect 66570 25560 66628 25572
rect 66570 24984 66582 25560
rect 66616 24984 66628 25560
rect 66570 24972 66628 24984
rect 67588 25560 67646 25572
rect 67588 24984 67600 25560
rect 67634 24984 67646 25560
rect 67588 24972 67646 24984
rect 68606 25560 68664 25572
rect 68606 24984 68618 25560
rect 68652 24984 68664 25560
rect 68606 24972 68664 24984
rect 69624 25560 69682 25572
rect 69624 24984 69636 25560
rect 69670 24984 69682 25560
rect 69624 24972 69682 24984
rect 70642 25560 70700 25572
rect 70642 24984 70654 25560
rect 70688 24984 70700 25560
rect 70642 24972 70700 24984
rect 71660 25560 71718 25572
rect 71660 24984 71672 25560
rect 71706 24984 71718 25560
rect 71660 24972 71718 24984
rect 72678 25560 72736 25572
rect 72678 24984 72690 25560
rect 72724 24984 72736 25560
rect 72678 24972 72736 24984
rect 73696 25560 73754 25572
rect 73696 24984 73708 25560
rect 73742 24984 73754 25560
rect 73696 24972 73754 24984
rect 74714 25560 74772 25572
rect 74714 24984 74726 25560
rect 74760 24984 74772 25560
rect 74714 24972 74772 24984
rect 59620 23922 59678 23934
rect 59620 23346 59632 23922
rect 59666 23346 59678 23922
rect 59620 23334 59678 23346
rect 60638 23922 60696 23934
rect 60638 23346 60650 23922
rect 60684 23346 60696 23922
rect 60638 23334 60696 23346
rect 61656 23922 61714 23934
rect 61656 23346 61668 23922
rect 61702 23346 61714 23922
rect 61656 23334 61714 23346
rect 62674 23922 62732 23934
rect 62674 23346 62686 23922
rect 62720 23346 62732 23922
rect 62674 23334 62732 23346
rect 63692 23922 63750 23934
rect 63692 23346 63704 23922
rect 63738 23346 63750 23922
rect 63692 23334 63750 23346
rect 64710 23922 64768 23934
rect 64710 23346 64722 23922
rect 64756 23346 64768 23922
rect 64710 23334 64768 23346
rect 65728 23922 65786 23934
rect 65728 23346 65740 23922
rect 65774 23346 65786 23922
rect 65728 23334 65786 23346
rect 66746 23922 66804 23934
rect 66746 23346 66758 23922
rect 66792 23346 66804 23922
rect 66746 23334 66804 23346
rect 67764 23922 67822 23934
rect 67764 23346 67776 23922
rect 67810 23346 67822 23922
rect 67764 23334 67822 23346
rect 68782 23922 68840 23934
rect 68782 23346 68794 23922
rect 68828 23346 68840 23922
rect 68782 23334 68840 23346
rect 69800 23922 69858 23934
rect 69800 23346 69812 23922
rect 69846 23346 69858 23922
rect 69800 23334 69858 23346
rect 70818 23922 70876 23934
rect 70818 23346 70830 23922
rect 70864 23346 70876 23922
rect 70818 23334 70876 23346
rect 71836 23922 71894 23934
rect 71836 23346 71848 23922
rect 71882 23346 71894 23922
rect 71836 23334 71894 23346
rect 72854 23922 72912 23934
rect 72854 23346 72866 23922
rect 72900 23346 72912 23922
rect 72854 23334 72912 23346
rect 73872 23922 73930 23934
rect 73872 23346 73884 23922
rect 73918 23346 73930 23922
rect 73872 23334 73930 23346
rect 59620 22890 59678 22902
rect 59620 22314 59632 22890
rect 59666 22314 59678 22890
rect 59620 22302 59678 22314
rect 60638 22890 60696 22902
rect 60638 22314 60650 22890
rect 60684 22314 60696 22890
rect 60638 22302 60696 22314
rect 61656 22890 61714 22902
rect 61656 22314 61668 22890
rect 61702 22314 61714 22890
rect 61656 22302 61714 22314
rect 62674 22890 62732 22902
rect 62674 22314 62686 22890
rect 62720 22314 62732 22890
rect 62674 22302 62732 22314
rect 63692 22890 63750 22902
rect 63692 22314 63704 22890
rect 63738 22314 63750 22890
rect 63692 22302 63750 22314
rect 64710 22890 64768 22902
rect 64710 22314 64722 22890
rect 64756 22314 64768 22890
rect 64710 22302 64768 22314
rect 65728 22890 65786 22902
rect 65728 22314 65740 22890
rect 65774 22314 65786 22890
rect 65728 22302 65786 22314
rect 66746 22890 66804 22902
rect 66746 22314 66758 22890
rect 66792 22314 66804 22890
rect 66746 22302 66804 22314
rect 67764 22890 67822 22902
rect 67764 22314 67776 22890
rect 67810 22314 67822 22890
rect 67764 22302 67822 22314
rect 68782 22890 68840 22902
rect 68782 22314 68794 22890
rect 68828 22314 68840 22890
rect 68782 22302 68840 22314
rect 69800 22890 69858 22902
rect 69800 22314 69812 22890
rect 69846 22314 69858 22890
rect 69800 22302 69858 22314
rect 70818 22890 70876 22902
rect 70818 22314 70830 22890
rect 70864 22314 70876 22890
rect 70818 22302 70876 22314
rect 71836 22890 71894 22902
rect 71836 22314 71848 22890
rect 71882 22314 71894 22890
rect 71836 22302 71894 22314
rect 72854 22890 72912 22902
rect 72854 22314 72866 22890
rect 72900 22314 72912 22890
rect 72854 22302 72912 22314
rect 73872 22890 73930 22902
rect 73872 22314 73884 22890
rect 73918 22314 73930 22890
rect 73872 22302 73930 22314
rect 59412 21286 59470 21298
rect 54108 21182 54166 21194
rect 54108 20606 54120 21182
rect 54154 20606 54166 21182
rect 54108 20594 54166 20606
rect 55126 21182 55184 21194
rect 55126 20606 55138 21182
rect 55172 20606 55184 21182
rect 55126 20594 55184 20606
rect 56144 21182 56202 21194
rect 56144 20606 56156 21182
rect 56190 20606 56202 21182
rect 56144 20594 56202 20606
rect 57162 21182 57220 21194
rect 57162 20606 57174 21182
rect 57208 20606 57220 21182
rect 57162 20594 57220 20606
rect 58180 21182 58238 21194
rect 58180 20606 58192 21182
rect 58226 20606 58238 21182
rect 59412 20710 59424 21286
rect 59458 20710 59470 21286
rect 59412 20698 59470 20710
rect 60430 21286 60488 21298
rect 60430 20710 60442 21286
rect 60476 20710 60488 21286
rect 60430 20698 60488 20710
rect 61448 21286 61506 21298
rect 61448 20710 61460 21286
rect 61494 20710 61506 21286
rect 61448 20698 61506 20710
rect 62466 21286 62524 21298
rect 62466 20710 62478 21286
rect 62512 20710 62524 21286
rect 62466 20698 62524 20710
rect 63484 21286 63542 21298
rect 63484 20710 63496 21286
rect 63530 20710 63542 21286
rect 63484 20698 63542 20710
rect 64502 21286 64560 21298
rect 64502 20710 64514 21286
rect 64548 20710 64560 21286
rect 64502 20698 64560 20710
rect 65520 21286 65578 21298
rect 65520 20710 65532 21286
rect 65566 20710 65578 21286
rect 65520 20698 65578 20710
rect 66538 21286 66596 21298
rect 66538 20710 66550 21286
rect 66584 20710 66596 21286
rect 66538 20698 66596 20710
rect 67556 21286 67614 21298
rect 67556 20710 67568 21286
rect 67602 20710 67614 21286
rect 67556 20698 67614 20710
rect 68574 21286 68632 21298
rect 68574 20710 68586 21286
rect 68620 20710 68632 21286
rect 68574 20698 68632 20710
rect 69592 21286 69650 21298
rect 69592 20710 69604 21286
rect 69638 20710 69650 21286
rect 69592 20698 69650 20710
rect 70610 21286 70668 21298
rect 70610 20710 70622 21286
rect 70656 20710 70668 21286
rect 70610 20698 70668 20710
rect 71628 21286 71686 21298
rect 71628 20710 71640 21286
rect 71674 20710 71686 21286
rect 71628 20698 71686 20710
rect 72646 21286 72704 21298
rect 72646 20710 72658 21286
rect 72692 20710 72704 21286
rect 72646 20698 72704 20710
rect 73664 21286 73722 21298
rect 73664 20710 73676 21286
rect 73710 20710 73722 21286
rect 73664 20698 73722 20710
rect 74682 21286 74740 21298
rect 74682 20710 74694 21286
rect 74728 20710 74740 21286
rect 74682 20698 74740 20710
rect 58180 20594 58238 20606
rect 54108 20150 54166 20162
rect 54108 19574 54120 20150
rect 54154 19574 54166 20150
rect 54108 19562 54166 19574
rect 55126 20150 55184 20162
rect 55126 19574 55138 20150
rect 55172 19574 55184 20150
rect 55126 19562 55184 19574
rect 56144 20150 56202 20162
rect 56144 19574 56156 20150
rect 56190 19574 56202 20150
rect 56144 19562 56202 19574
rect 57162 20150 57220 20162
rect 57162 19574 57174 20150
rect 57208 19574 57220 20150
rect 57162 19562 57220 19574
rect 58180 20150 58238 20162
rect 58180 19574 58192 20150
rect 58226 19574 58238 20150
rect 58180 19562 58238 19574
rect 59412 20030 59470 20042
rect 59412 19454 59424 20030
rect 59458 19454 59470 20030
rect 59412 19442 59470 19454
rect 60430 20030 60488 20042
rect 60430 19454 60442 20030
rect 60476 19454 60488 20030
rect 60430 19442 60488 19454
rect 61448 20030 61506 20042
rect 61448 19454 61460 20030
rect 61494 19454 61506 20030
rect 61448 19442 61506 19454
rect 62466 20030 62524 20042
rect 62466 19454 62478 20030
rect 62512 19454 62524 20030
rect 62466 19442 62524 19454
rect 63484 20030 63542 20042
rect 63484 19454 63496 20030
rect 63530 19454 63542 20030
rect 63484 19442 63542 19454
rect 64502 20030 64560 20042
rect 64502 19454 64514 20030
rect 64548 19454 64560 20030
rect 64502 19442 64560 19454
rect 65520 20030 65578 20042
rect 65520 19454 65532 20030
rect 65566 19454 65578 20030
rect 65520 19442 65578 19454
rect 66538 20030 66596 20042
rect 66538 19454 66550 20030
rect 66584 19454 66596 20030
rect 66538 19442 66596 19454
rect 67556 20030 67614 20042
rect 67556 19454 67568 20030
rect 67602 19454 67614 20030
rect 67556 19442 67614 19454
rect 68574 20030 68632 20042
rect 68574 19454 68586 20030
rect 68620 19454 68632 20030
rect 68574 19442 68632 19454
rect 69592 20030 69650 20042
rect 69592 19454 69604 20030
rect 69638 19454 69650 20030
rect 69592 19442 69650 19454
rect 70610 20030 70668 20042
rect 70610 19454 70622 20030
rect 70656 19454 70668 20030
rect 70610 19442 70668 19454
rect 71628 20030 71686 20042
rect 71628 19454 71640 20030
rect 71674 19454 71686 20030
rect 71628 19442 71686 19454
rect 72646 20030 72704 20042
rect 72646 19454 72658 20030
rect 72692 19454 72704 20030
rect 72646 19442 72704 19454
rect 73664 20030 73722 20042
rect 73664 19454 73676 20030
rect 73710 19454 73722 20030
rect 73664 19442 73722 19454
rect 74682 20030 74740 20042
rect 74682 19454 74694 20030
rect 74728 19454 74740 20030
rect 74682 19442 74740 19454
rect 54108 19118 54166 19130
rect 54108 18542 54120 19118
rect 54154 18542 54166 19118
rect 54108 18530 54166 18542
rect 55126 19118 55184 19130
rect 55126 18542 55138 19118
rect 55172 18542 55184 19118
rect 55126 18530 55184 18542
rect 56144 19118 56202 19130
rect 56144 18542 56156 19118
rect 56190 18542 56202 19118
rect 56144 18530 56202 18542
rect 57162 19118 57220 19130
rect 57162 18542 57174 19118
rect 57208 18542 57220 19118
rect 57162 18530 57220 18542
rect 58180 19118 58238 19130
rect 58180 18542 58192 19118
rect 58226 18542 58238 19118
rect 58180 18530 58238 18542
rect 59412 18774 59470 18786
rect 59412 18198 59424 18774
rect 59458 18198 59470 18774
rect 59412 18186 59470 18198
rect 60430 18774 60488 18786
rect 60430 18198 60442 18774
rect 60476 18198 60488 18774
rect 60430 18186 60488 18198
rect 61448 18774 61506 18786
rect 61448 18198 61460 18774
rect 61494 18198 61506 18774
rect 61448 18186 61506 18198
rect 62466 18774 62524 18786
rect 62466 18198 62478 18774
rect 62512 18198 62524 18774
rect 62466 18186 62524 18198
rect 63484 18774 63542 18786
rect 63484 18198 63496 18774
rect 63530 18198 63542 18774
rect 63484 18186 63542 18198
rect 64502 18774 64560 18786
rect 64502 18198 64514 18774
rect 64548 18198 64560 18774
rect 64502 18186 64560 18198
rect 65520 18774 65578 18786
rect 65520 18198 65532 18774
rect 65566 18198 65578 18774
rect 65520 18186 65578 18198
rect 66538 18774 66596 18786
rect 66538 18198 66550 18774
rect 66584 18198 66596 18774
rect 66538 18186 66596 18198
rect 67556 18774 67614 18786
rect 67556 18198 67568 18774
rect 67602 18198 67614 18774
rect 67556 18186 67614 18198
rect 68574 18774 68632 18786
rect 68574 18198 68586 18774
rect 68620 18198 68632 18774
rect 68574 18186 68632 18198
rect 69592 18774 69650 18786
rect 69592 18198 69604 18774
rect 69638 18198 69650 18774
rect 69592 18186 69650 18198
rect 70610 18774 70668 18786
rect 70610 18198 70622 18774
rect 70656 18198 70668 18774
rect 70610 18186 70668 18198
rect 71628 18774 71686 18786
rect 71628 18198 71640 18774
rect 71674 18198 71686 18774
rect 71628 18186 71686 18198
rect 72646 18774 72704 18786
rect 72646 18198 72658 18774
rect 72692 18198 72704 18774
rect 72646 18186 72704 18198
rect 73664 18774 73722 18786
rect 73664 18198 73676 18774
rect 73710 18198 73722 18774
rect 73664 18186 73722 18198
rect 74682 18774 74740 18786
rect 74682 18198 74694 18774
rect 74728 18198 74740 18774
rect 74682 18186 74740 18198
rect 54108 18086 54166 18098
rect 54108 17510 54120 18086
rect 54154 17510 54166 18086
rect 54108 17498 54166 17510
rect 55126 18086 55184 18098
rect 55126 17510 55138 18086
rect 55172 17510 55184 18086
rect 55126 17498 55184 17510
rect 56144 18086 56202 18098
rect 56144 17510 56156 18086
rect 56190 17510 56202 18086
rect 56144 17498 56202 17510
rect 57162 18086 57220 18098
rect 57162 17510 57174 18086
rect 57208 17510 57220 18086
rect 57162 17498 57220 17510
rect 58180 18086 58238 18098
rect 58180 17510 58192 18086
rect 58226 17510 58238 18086
rect 58180 17498 58238 17510
rect 59412 17518 59470 17530
rect 59412 16942 59424 17518
rect 59458 16942 59470 17518
rect 59412 16930 59470 16942
rect 60430 17518 60488 17530
rect 60430 16942 60442 17518
rect 60476 16942 60488 17518
rect 60430 16930 60488 16942
rect 61448 17518 61506 17530
rect 61448 16942 61460 17518
rect 61494 16942 61506 17518
rect 61448 16930 61506 16942
rect 62466 17518 62524 17530
rect 62466 16942 62478 17518
rect 62512 16942 62524 17518
rect 62466 16930 62524 16942
rect 63484 17518 63542 17530
rect 63484 16942 63496 17518
rect 63530 16942 63542 17518
rect 63484 16930 63542 16942
rect 64502 17518 64560 17530
rect 64502 16942 64514 17518
rect 64548 16942 64560 17518
rect 64502 16930 64560 16942
rect 65520 17518 65578 17530
rect 65520 16942 65532 17518
rect 65566 16942 65578 17518
rect 65520 16930 65578 16942
rect 66538 17518 66596 17530
rect 66538 16942 66550 17518
rect 66584 16942 66596 17518
rect 66538 16930 66596 16942
rect 67556 17518 67614 17530
rect 67556 16942 67568 17518
rect 67602 16942 67614 17518
rect 67556 16930 67614 16942
rect 68574 17518 68632 17530
rect 68574 16942 68586 17518
rect 68620 16942 68632 17518
rect 68574 16930 68632 16942
rect 69592 17518 69650 17530
rect 69592 16942 69604 17518
rect 69638 16942 69650 17518
rect 69592 16930 69650 16942
rect 70610 17518 70668 17530
rect 70610 16942 70622 17518
rect 70656 16942 70668 17518
rect 70610 16930 70668 16942
rect 71628 17518 71686 17530
rect 71628 16942 71640 17518
rect 71674 16942 71686 17518
rect 71628 16930 71686 16942
rect 72646 17518 72704 17530
rect 72646 16942 72658 17518
rect 72692 16942 72704 17518
rect 72646 16930 72704 16942
rect 73664 17518 73722 17530
rect 73664 16942 73676 17518
rect 73710 16942 73722 17518
rect 73664 16930 73722 16942
rect 74682 17518 74740 17530
rect 74682 16942 74694 17518
rect 74728 16942 74740 17518
rect 74682 16930 74740 16942
rect 36898 12986 36956 12998
rect 36898 12810 36910 12986
rect 36944 12810 36956 12986
rect 36898 12798 36956 12810
rect 37156 12986 37214 12998
rect 37156 12810 37168 12986
rect 37202 12810 37214 12986
rect 37156 12798 37214 12810
rect 37414 12986 37472 12998
rect 37414 12810 37426 12986
rect 37460 12810 37472 12986
rect 37414 12798 37472 12810
rect 37672 12986 37730 12998
rect 37672 12810 37684 12986
rect 37718 12810 37730 12986
rect 37672 12798 37730 12810
rect 37930 12986 37988 12998
rect 37930 12810 37942 12986
rect 37976 12810 37988 12986
rect 37930 12798 37988 12810
rect 38188 12986 38246 12998
rect 38188 12810 38200 12986
rect 38234 12810 38246 12986
rect 38188 12798 38246 12810
rect 38446 12986 38504 12998
rect 38446 12810 38458 12986
rect 38492 12810 38504 12986
rect 38446 12798 38504 12810
<< ndiffc >>
rect 1766 13270 1800 13846
rect 2784 13270 2818 13846
rect 3802 13270 3836 13846
rect 4820 13270 4854 13846
rect 5838 13270 5872 13846
rect 6856 13270 6890 13846
rect 7874 13270 7908 13846
rect 8892 13270 8926 13846
rect 9910 13270 9944 13846
rect 10928 13270 10962 13846
rect 13532 13746 13566 14322
rect 14550 13746 14584 14322
rect 15568 13746 15602 14322
rect 16586 13746 16620 14322
rect 17604 13746 17638 14322
rect 18622 13746 18656 14322
rect 19640 13746 19674 14322
rect 20658 13746 20692 14322
rect 21676 13746 21710 14322
rect 22694 13746 22728 14322
rect 23712 13746 23746 14322
rect 24730 13746 24764 14322
rect 25748 13746 25782 14322
rect 26766 13746 26800 14322
rect 27784 13746 27818 14322
rect 28802 13746 28836 14322
rect 29820 13746 29854 14322
rect 30838 13746 30872 14322
rect 31856 13746 31890 14322
rect 32874 13746 32908 14322
rect 33892 13746 33926 14322
rect 1766 12452 1800 13028
rect 2784 12452 2818 13028
rect 3802 12452 3836 13028
rect 4820 12452 4854 13028
rect 5838 12452 5872 13028
rect 6856 12452 6890 13028
rect 7874 12452 7908 13028
rect 8892 12452 8926 13028
rect 9910 12452 9944 13028
rect 10928 12452 10962 13028
rect 13532 12928 13566 13504
rect 14550 12928 14584 13504
rect 15568 12928 15602 13504
rect 16586 12928 16620 13504
rect 17604 12928 17638 13504
rect 18622 12928 18656 13504
rect 19640 12928 19674 13504
rect 20658 12928 20692 13504
rect 21676 12928 21710 13504
rect 22694 12928 22728 13504
rect 23712 12928 23746 13504
rect 24730 12928 24764 13504
rect 25748 12928 25782 13504
rect 26766 12928 26800 13504
rect 27784 12928 27818 13504
rect 28802 12928 28836 13504
rect 29820 12928 29854 13504
rect 30838 12928 30872 13504
rect 31856 12928 31890 13504
rect 32874 12928 32908 13504
rect 33892 12928 33926 13504
rect 1766 11634 1800 12210
rect 2784 11634 2818 12210
rect 3802 11634 3836 12210
rect 4820 11634 4854 12210
rect 5838 11634 5872 12210
rect 6856 11634 6890 12210
rect 7874 11634 7908 12210
rect 8892 11634 8926 12210
rect 9910 11634 9944 12210
rect 10928 11634 10962 12210
rect 13532 11550 13566 12126
rect 14550 11550 14584 12126
rect 15568 11550 15602 12126
rect 16586 11550 16620 12126
rect 17604 11550 17638 12126
rect 18622 11550 18656 12126
rect 19640 11550 19674 12126
rect 20658 11550 20692 12126
rect 21676 11550 21710 12126
rect 22694 11550 22728 12126
rect 23712 11550 23746 12126
rect 24730 11550 24764 12126
rect 25748 11550 25782 12126
rect 26766 11550 26800 12126
rect 27784 11550 27818 12126
rect 28802 11550 28836 12126
rect 29820 11550 29854 12126
rect 30838 11550 30872 12126
rect 31856 11550 31890 12126
rect 32874 11550 32908 12126
rect 33892 11550 33926 12126
rect 1766 10816 1800 11392
rect 2784 10816 2818 11392
rect 3802 10816 3836 11392
rect 4820 10816 4854 11392
rect 5838 10816 5872 11392
rect 6856 10816 6890 11392
rect 7874 10816 7908 11392
rect 8892 10816 8926 11392
rect 9910 10816 9944 11392
rect 10928 10816 10962 11392
rect 1766 9998 1800 10574
rect 2784 9998 2818 10574
rect 3802 9998 3836 10574
rect 4820 9998 4854 10574
rect 5838 9998 5872 10574
rect 6856 9998 6890 10574
rect 7874 9998 7908 10574
rect 8892 9998 8926 10574
rect 9910 9998 9944 10574
rect 10928 9998 10962 10574
rect 13532 10318 13566 10894
rect 14550 10318 14584 10894
rect 15568 10318 15602 10894
rect 16586 10318 16620 10894
rect 17604 10318 17638 10894
rect 18622 10318 18656 10894
rect 19640 10318 19674 10894
rect 20658 10318 20692 10894
rect 21676 10318 21710 10894
rect 22694 10318 22728 10894
rect 23712 10318 23746 10894
rect 24730 10318 24764 10894
rect 25748 10318 25782 10894
rect 26766 10318 26800 10894
rect 27784 10318 27818 10894
rect 28802 10318 28836 10894
rect 29820 10318 29854 10894
rect 30838 10318 30872 10894
rect 31856 10318 31890 10894
rect 32874 10318 32908 10894
rect 33892 10318 33926 10894
rect 1766 9180 1800 9756
rect 2784 9180 2818 9756
rect 3802 9180 3836 9756
rect 4820 9180 4854 9756
rect 5838 9180 5872 9756
rect 6856 9180 6890 9756
rect 7874 9180 7908 9756
rect 8892 9180 8926 9756
rect 9910 9180 9944 9756
rect 10928 9180 10962 9756
rect 13530 9084 13564 9660
rect 14548 9084 14582 9660
rect 15566 9084 15600 9660
rect 16584 9084 16618 9660
rect 17602 9084 17636 9660
rect 18620 9084 18654 9660
rect 19638 9084 19672 9660
rect 20656 9084 20690 9660
rect 21674 9084 21708 9660
rect 22692 9084 22726 9660
rect 23710 9084 23744 9660
rect 24728 9084 24762 9660
rect 25746 9084 25780 9660
rect 26764 9084 26798 9660
rect 27782 9084 27816 9660
rect 28800 9084 28834 9660
rect 29818 9084 29852 9660
rect 30836 9084 30870 9660
rect 31854 9084 31888 9660
rect 32872 9084 32906 9660
rect 33890 9084 33924 9660
rect 1766 8362 1800 8938
rect 2784 8362 2818 8938
rect 3802 8362 3836 8938
rect 4820 8362 4854 8938
rect 5838 8362 5872 8938
rect 6856 8362 6890 8938
rect 7874 8362 7908 8938
rect 8892 8362 8926 8938
rect 9910 8362 9944 8938
rect 10928 8362 10962 8938
rect 1766 7544 1800 8120
rect 2784 7544 2818 8120
rect 3802 7544 3836 8120
rect 4820 7544 4854 8120
rect 5838 7544 5872 8120
rect 6856 7544 6890 8120
rect 7874 7544 7908 8120
rect 8892 7544 8926 8120
rect 9910 7544 9944 8120
rect 10928 7544 10962 8120
rect 13530 7850 13564 8426
rect 14548 7850 14582 8426
rect 15566 7850 15600 8426
rect 16584 7850 16618 8426
rect 17602 7850 17636 8426
rect 18620 7850 18654 8426
rect 19638 7850 19672 8426
rect 20656 7850 20690 8426
rect 21674 7850 21708 8426
rect 22692 7850 22726 8426
rect 23710 7850 23744 8426
rect 24728 7850 24762 8426
rect 25746 7850 25780 8426
rect 26764 7850 26798 8426
rect 27782 7850 27816 8426
rect 28800 7850 28834 8426
rect 29818 7850 29852 8426
rect 30836 7850 30870 8426
rect 31854 7850 31888 8426
rect 32872 7850 32906 8426
rect 33890 7850 33924 8426
rect 13530 6618 13564 7194
rect 14548 6618 14582 7194
rect 15566 6618 15600 7194
rect 16584 6618 16618 7194
rect 17602 6618 17636 7194
rect 18620 6618 18654 7194
rect 19638 6618 19672 7194
rect 20656 6618 20690 7194
rect 21674 6618 21708 7194
rect 22692 6618 22726 7194
rect 23710 6618 23744 7194
rect 24728 6618 24762 7194
rect 25746 6618 25780 7194
rect 26764 6618 26798 7194
rect 27782 6618 27816 7194
rect 28800 6618 28834 7194
rect 29818 6618 29852 7194
rect 30836 6618 30870 7194
rect 31854 6618 31888 7194
rect 32872 6618 32906 7194
rect 33890 6618 33924 7194
rect 442 5520 476 6096
rect 1460 5520 1494 6096
rect 2478 5520 2512 6096
rect 3496 5520 3530 6096
rect 4514 5520 4548 6096
rect 5532 5520 5566 6096
rect 6550 5520 6584 6096
rect 7568 5520 7602 6096
rect 8586 5520 8620 6096
rect 9604 5520 9638 6096
rect 10622 5520 10656 6096
rect 11640 5520 11674 6096
rect 13530 5384 13564 5960
rect 14548 5384 14582 5960
rect 15566 5384 15600 5960
rect 16584 5384 16618 5960
rect 17602 5384 17636 5960
rect 18620 5384 18654 5960
rect 19638 5384 19672 5960
rect 20656 5384 20690 5960
rect 21674 5384 21708 5960
rect 22692 5384 22726 5960
rect 23710 5384 23744 5960
rect 24728 5384 24762 5960
rect 25746 5384 25780 5960
rect 26764 5384 26798 5960
rect 27782 5384 27816 5960
rect 28800 5384 28834 5960
rect 29818 5384 29852 5960
rect 30836 5384 30870 5960
rect 31854 5384 31888 5960
rect 32872 5384 32906 5960
rect 33890 5384 33924 5960
rect 442 4408 476 4984
rect 1460 4408 1494 4984
rect 2478 4408 2512 4984
rect 3496 4408 3530 4984
rect 4514 4408 4548 4984
rect 5532 4408 5566 4984
rect 6550 4408 6584 4984
rect 7568 4408 7602 4984
rect 8586 4408 8620 4984
rect 9604 4408 9638 4984
rect 10622 4408 10656 4984
rect 11640 4408 11674 4984
rect 13530 4150 13564 4726
rect 14548 4150 14582 4726
rect 15566 4150 15600 4726
rect 16584 4150 16618 4726
rect 17602 4150 17636 4726
rect 18620 4150 18654 4726
rect 19638 4150 19672 4726
rect 20656 4150 20690 4726
rect 21674 4150 21708 4726
rect 22692 4150 22726 4726
rect 23710 4150 23744 4726
rect 24728 4150 24762 4726
rect 25746 4150 25780 4726
rect 26764 4150 26798 4726
rect 27782 4150 27816 4726
rect 28800 4150 28834 4726
rect 29818 4150 29852 4726
rect 30836 4150 30870 4726
rect 31854 4150 31888 4726
rect 32872 4150 32906 4726
rect 33890 4150 33924 4726
rect 442 3296 476 3872
rect 1460 3296 1494 3872
rect 2478 3296 2512 3872
rect 3496 3296 3530 3872
rect 4514 3296 4548 3872
rect 5532 3296 5566 3872
rect 6550 3296 6584 3872
rect 7568 3296 7602 3872
rect 8586 3296 8620 3872
rect 9604 3296 9638 3872
rect 10622 3296 10656 3872
rect 11640 3296 11674 3872
rect 13530 2918 13564 3494
rect 14548 2918 14582 3494
rect 15566 2918 15600 3494
rect 16584 2918 16618 3494
rect 17602 2918 17636 3494
rect 18620 2918 18654 3494
rect 19638 2918 19672 3494
rect 20656 2918 20690 3494
rect 21674 2918 21708 3494
rect 22692 2918 22726 3494
rect 23710 2918 23744 3494
rect 24728 2918 24762 3494
rect 25746 2918 25780 3494
rect 26764 2918 26798 3494
rect 27782 2918 27816 3494
rect 28800 2918 28834 3494
rect 29818 2918 29852 3494
rect 30836 2918 30870 3494
rect 31854 2918 31888 3494
rect 32872 2918 32906 3494
rect 33890 2918 33924 3494
rect 442 2184 476 2760
rect 1460 2184 1494 2760
rect 2478 2184 2512 2760
rect 3496 2184 3530 2760
rect 4514 2184 4548 2760
rect 5532 2184 5566 2760
rect 6550 2184 6584 2760
rect 7568 2184 7602 2760
rect 8586 2184 8620 2760
rect 9604 2184 9638 2760
rect 10622 2184 10656 2760
rect 11640 2184 11674 2760
rect 13530 1684 13564 2260
rect 14548 1684 14582 2260
rect 15566 1684 15600 2260
rect 16584 1684 16618 2260
rect 17602 1684 17636 2260
rect 18620 1684 18654 2260
rect 19638 1684 19672 2260
rect 20656 1684 20690 2260
rect 21674 1684 21708 2260
rect 22692 1684 22726 2260
rect 23710 1684 23744 2260
rect 24728 1684 24762 2260
rect 25746 1684 25780 2260
rect 26764 1684 26798 2260
rect 27782 1684 27816 2260
rect 28800 1684 28834 2260
rect 29818 1684 29852 2260
rect 30836 1684 30870 2260
rect 31854 1684 31888 2260
rect 32872 1684 32906 2260
rect 33890 1684 33924 2260
rect 900 642 934 1218
rect 1918 642 1952 1218
rect 2936 642 2970 1218
rect 3954 642 3988 1218
rect 4972 642 5006 1218
rect 5990 642 6024 1218
rect 7008 642 7042 1218
rect 8026 642 8060 1218
rect 9044 642 9078 1218
rect 10062 642 10096 1218
rect 11080 642 11114 1218
rect 13530 452 13564 1028
rect 14548 452 14582 1028
rect 15566 452 15600 1028
rect 16584 452 16618 1028
rect 17602 452 17636 1028
rect 18620 452 18654 1028
rect 19638 452 19672 1028
rect 20656 452 20690 1028
rect 21674 452 21708 1028
rect 22692 452 22726 1028
rect 23710 452 23744 1028
rect 24728 452 24762 1028
rect 25746 452 25780 1028
rect 26764 452 26798 1028
rect 27782 452 27816 1028
rect 28800 452 28834 1028
rect 29818 452 29852 1028
rect 30836 452 30870 1028
rect 31854 452 31888 1028
rect 32872 452 32906 1028
rect 33890 452 33924 1028
rect -1074 84 -1040 190
rect -986 84 -952 190
rect 42766 13270 42800 13846
rect 43784 13270 43818 13846
rect 44802 13270 44836 13846
rect 45820 13270 45854 13846
rect 46838 13270 46872 13846
rect 47856 13270 47890 13846
rect 48874 13270 48908 13846
rect 49892 13270 49926 13846
rect 50910 13270 50944 13846
rect 51928 13270 51962 13846
rect 54532 13746 54566 14322
rect 55550 13746 55584 14322
rect 56568 13746 56602 14322
rect 57586 13746 57620 14322
rect 58604 13746 58638 14322
rect 59622 13746 59656 14322
rect 60640 13746 60674 14322
rect 61658 13746 61692 14322
rect 62676 13746 62710 14322
rect 63694 13746 63728 14322
rect 64712 13746 64746 14322
rect 65730 13746 65764 14322
rect 66748 13746 66782 14322
rect 67766 13746 67800 14322
rect 68784 13746 68818 14322
rect 69802 13746 69836 14322
rect 70820 13746 70854 14322
rect 71838 13746 71872 14322
rect 72856 13746 72890 14322
rect 73874 13746 73908 14322
rect 74892 13746 74926 14322
rect 42766 12452 42800 13028
rect 43784 12452 43818 13028
rect 44802 12452 44836 13028
rect 45820 12452 45854 13028
rect 46838 12452 46872 13028
rect 47856 12452 47890 13028
rect 48874 12452 48908 13028
rect 49892 12452 49926 13028
rect 50910 12452 50944 13028
rect 51928 12452 51962 13028
rect 54532 12928 54566 13504
rect 55550 12928 55584 13504
rect 56568 12928 56602 13504
rect 57586 12928 57620 13504
rect 58604 12928 58638 13504
rect 59622 12928 59656 13504
rect 60640 12928 60674 13504
rect 61658 12928 61692 13504
rect 62676 12928 62710 13504
rect 63694 12928 63728 13504
rect 64712 12928 64746 13504
rect 65730 12928 65764 13504
rect 66748 12928 66782 13504
rect 67766 12928 67800 13504
rect 68784 12928 68818 13504
rect 69802 12928 69836 13504
rect 70820 12928 70854 13504
rect 71838 12928 71872 13504
rect 72856 12928 72890 13504
rect 73874 12928 73908 13504
rect 74892 12928 74926 13504
rect 42766 11634 42800 12210
rect 43784 11634 43818 12210
rect 44802 11634 44836 12210
rect 45820 11634 45854 12210
rect 46838 11634 46872 12210
rect 47856 11634 47890 12210
rect 48874 11634 48908 12210
rect 49892 11634 49926 12210
rect 50910 11634 50944 12210
rect 51928 11634 51962 12210
rect 54532 11550 54566 12126
rect 55550 11550 55584 12126
rect 56568 11550 56602 12126
rect 57586 11550 57620 12126
rect 58604 11550 58638 12126
rect 59622 11550 59656 12126
rect 60640 11550 60674 12126
rect 61658 11550 61692 12126
rect 62676 11550 62710 12126
rect 63694 11550 63728 12126
rect 64712 11550 64746 12126
rect 65730 11550 65764 12126
rect 66748 11550 66782 12126
rect 67766 11550 67800 12126
rect 68784 11550 68818 12126
rect 69802 11550 69836 12126
rect 70820 11550 70854 12126
rect 71838 11550 71872 12126
rect 72856 11550 72890 12126
rect 73874 11550 73908 12126
rect 74892 11550 74926 12126
rect 42766 10816 42800 11392
rect 43784 10816 43818 11392
rect 44802 10816 44836 11392
rect 45820 10816 45854 11392
rect 46838 10816 46872 11392
rect 47856 10816 47890 11392
rect 48874 10816 48908 11392
rect 49892 10816 49926 11392
rect 50910 10816 50944 11392
rect 51928 10816 51962 11392
rect 42766 9998 42800 10574
rect 43784 9998 43818 10574
rect 44802 9998 44836 10574
rect 45820 9998 45854 10574
rect 46838 9998 46872 10574
rect 47856 9998 47890 10574
rect 48874 9998 48908 10574
rect 49892 9998 49926 10574
rect 50910 9998 50944 10574
rect 51928 9998 51962 10574
rect 54532 10318 54566 10894
rect 55550 10318 55584 10894
rect 56568 10318 56602 10894
rect 57586 10318 57620 10894
rect 58604 10318 58638 10894
rect 59622 10318 59656 10894
rect 60640 10318 60674 10894
rect 61658 10318 61692 10894
rect 62676 10318 62710 10894
rect 63694 10318 63728 10894
rect 64712 10318 64746 10894
rect 65730 10318 65764 10894
rect 66748 10318 66782 10894
rect 67766 10318 67800 10894
rect 68784 10318 68818 10894
rect 69802 10318 69836 10894
rect 70820 10318 70854 10894
rect 71838 10318 71872 10894
rect 72856 10318 72890 10894
rect 73874 10318 73908 10894
rect 74892 10318 74926 10894
rect 42766 9180 42800 9756
rect 43784 9180 43818 9756
rect 44802 9180 44836 9756
rect 45820 9180 45854 9756
rect 46838 9180 46872 9756
rect 47856 9180 47890 9756
rect 48874 9180 48908 9756
rect 49892 9180 49926 9756
rect 50910 9180 50944 9756
rect 51928 9180 51962 9756
rect 54530 9084 54564 9660
rect 55548 9084 55582 9660
rect 56566 9084 56600 9660
rect 57584 9084 57618 9660
rect 58602 9084 58636 9660
rect 59620 9084 59654 9660
rect 60638 9084 60672 9660
rect 61656 9084 61690 9660
rect 62674 9084 62708 9660
rect 63692 9084 63726 9660
rect 64710 9084 64744 9660
rect 65728 9084 65762 9660
rect 66746 9084 66780 9660
rect 67764 9084 67798 9660
rect 68782 9084 68816 9660
rect 69800 9084 69834 9660
rect 70818 9084 70852 9660
rect 71836 9084 71870 9660
rect 72854 9084 72888 9660
rect 73872 9084 73906 9660
rect 74890 9084 74924 9660
rect 42766 8362 42800 8938
rect 43784 8362 43818 8938
rect 44802 8362 44836 8938
rect 45820 8362 45854 8938
rect 46838 8362 46872 8938
rect 47856 8362 47890 8938
rect 48874 8362 48908 8938
rect 49892 8362 49926 8938
rect 50910 8362 50944 8938
rect 51928 8362 51962 8938
rect 42766 7544 42800 8120
rect 43784 7544 43818 8120
rect 44802 7544 44836 8120
rect 45820 7544 45854 8120
rect 46838 7544 46872 8120
rect 47856 7544 47890 8120
rect 48874 7544 48908 8120
rect 49892 7544 49926 8120
rect 50910 7544 50944 8120
rect 51928 7544 51962 8120
rect 54530 7850 54564 8426
rect 55548 7850 55582 8426
rect 56566 7850 56600 8426
rect 57584 7850 57618 8426
rect 58602 7850 58636 8426
rect 59620 7850 59654 8426
rect 60638 7850 60672 8426
rect 61656 7850 61690 8426
rect 62674 7850 62708 8426
rect 63692 7850 63726 8426
rect 64710 7850 64744 8426
rect 65728 7850 65762 8426
rect 66746 7850 66780 8426
rect 67764 7850 67798 8426
rect 68782 7850 68816 8426
rect 69800 7850 69834 8426
rect 70818 7850 70852 8426
rect 71836 7850 71870 8426
rect 72854 7850 72888 8426
rect 73872 7850 73906 8426
rect 74890 7850 74924 8426
rect 54530 6618 54564 7194
rect 55548 6618 55582 7194
rect 56566 6618 56600 7194
rect 57584 6618 57618 7194
rect 58602 6618 58636 7194
rect 59620 6618 59654 7194
rect 60638 6618 60672 7194
rect 61656 6618 61690 7194
rect 62674 6618 62708 7194
rect 63692 6618 63726 7194
rect 64710 6618 64744 7194
rect 65728 6618 65762 7194
rect 66746 6618 66780 7194
rect 67764 6618 67798 7194
rect 68782 6618 68816 7194
rect 69800 6618 69834 7194
rect 70818 6618 70852 7194
rect 71836 6618 71870 7194
rect 72854 6618 72888 7194
rect 73872 6618 73906 7194
rect 74890 6618 74924 7194
rect 41442 5520 41476 6096
rect 42460 5520 42494 6096
rect 43478 5520 43512 6096
rect 44496 5520 44530 6096
rect 45514 5520 45548 6096
rect 46532 5520 46566 6096
rect 47550 5520 47584 6096
rect 48568 5520 48602 6096
rect 49586 5520 49620 6096
rect 50604 5520 50638 6096
rect 51622 5520 51656 6096
rect 52640 5520 52674 6096
rect 54530 5384 54564 5960
rect 55548 5384 55582 5960
rect 56566 5384 56600 5960
rect 57584 5384 57618 5960
rect 58602 5384 58636 5960
rect 59620 5384 59654 5960
rect 60638 5384 60672 5960
rect 61656 5384 61690 5960
rect 62674 5384 62708 5960
rect 63692 5384 63726 5960
rect 64710 5384 64744 5960
rect 65728 5384 65762 5960
rect 66746 5384 66780 5960
rect 67764 5384 67798 5960
rect 68782 5384 68816 5960
rect 69800 5384 69834 5960
rect 70818 5384 70852 5960
rect 71836 5384 71870 5960
rect 72854 5384 72888 5960
rect 73872 5384 73906 5960
rect 74890 5384 74924 5960
rect 41442 4408 41476 4984
rect 42460 4408 42494 4984
rect 43478 4408 43512 4984
rect 44496 4408 44530 4984
rect 45514 4408 45548 4984
rect 46532 4408 46566 4984
rect 47550 4408 47584 4984
rect 48568 4408 48602 4984
rect 49586 4408 49620 4984
rect 50604 4408 50638 4984
rect 51622 4408 51656 4984
rect 52640 4408 52674 4984
rect 54530 4150 54564 4726
rect 55548 4150 55582 4726
rect 56566 4150 56600 4726
rect 57584 4150 57618 4726
rect 58602 4150 58636 4726
rect 59620 4150 59654 4726
rect 60638 4150 60672 4726
rect 61656 4150 61690 4726
rect 62674 4150 62708 4726
rect 63692 4150 63726 4726
rect 64710 4150 64744 4726
rect 65728 4150 65762 4726
rect 66746 4150 66780 4726
rect 67764 4150 67798 4726
rect 68782 4150 68816 4726
rect 69800 4150 69834 4726
rect 70818 4150 70852 4726
rect 71836 4150 71870 4726
rect 72854 4150 72888 4726
rect 73872 4150 73906 4726
rect 74890 4150 74924 4726
rect 41442 3296 41476 3872
rect 42460 3296 42494 3872
rect 43478 3296 43512 3872
rect 44496 3296 44530 3872
rect 45514 3296 45548 3872
rect 46532 3296 46566 3872
rect 47550 3296 47584 3872
rect 48568 3296 48602 3872
rect 49586 3296 49620 3872
rect 50604 3296 50638 3872
rect 51622 3296 51656 3872
rect 52640 3296 52674 3872
rect 54530 2918 54564 3494
rect 55548 2918 55582 3494
rect 56566 2918 56600 3494
rect 57584 2918 57618 3494
rect 58602 2918 58636 3494
rect 59620 2918 59654 3494
rect 60638 2918 60672 3494
rect 61656 2918 61690 3494
rect 62674 2918 62708 3494
rect 63692 2918 63726 3494
rect 64710 2918 64744 3494
rect 65728 2918 65762 3494
rect 66746 2918 66780 3494
rect 67764 2918 67798 3494
rect 68782 2918 68816 3494
rect 69800 2918 69834 3494
rect 70818 2918 70852 3494
rect 71836 2918 71870 3494
rect 72854 2918 72888 3494
rect 73872 2918 73906 3494
rect 74890 2918 74924 3494
rect 41442 2184 41476 2760
rect 42460 2184 42494 2760
rect 43478 2184 43512 2760
rect 44496 2184 44530 2760
rect 45514 2184 45548 2760
rect 46532 2184 46566 2760
rect 47550 2184 47584 2760
rect 48568 2184 48602 2760
rect 49586 2184 49620 2760
rect 50604 2184 50638 2760
rect 51622 2184 51656 2760
rect 52640 2184 52674 2760
rect 54530 1684 54564 2260
rect 55548 1684 55582 2260
rect 56566 1684 56600 2260
rect 57584 1684 57618 2260
rect 58602 1684 58636 2260
rect 59620 1684 59654 2260
rect 60638 1684 60672 2260
rect 61656 1684 61690 2260
rect 62674 1684 62708 2260
rect 63692 1684 63726 2260
rect 64710 1684 64744 2260
rect 65728 1684 65762 2260
rect 66746 1684 66780 2260
rect 67764 1684 67798 2260
rect 68782 1684 68816 2260
rect 69800 1684 69834 2260
rect 70818 1684 70852 2260
rect 71836 1684 71870 2260
rect 72854 1684 72888 2260
rect 73872 1684 73906 2260
rect 74890 1684 74924 2260
rect 41900 642 41934 1218
rect 42918 642 42952 1218
rect 43936 642 43970 1218
rect 44954 642 44988 1218
rect 45972 642 46006 1218
rect 46990 642 47024 1218
rect 48008 642 48042 1218
rect 49026 642 49060 1218
rect 50044 642 50078 1218
rect 51062 642 51096 1218
rect 52080 642 52114 1218
rect 54530 452 54564 1028
rect 55548 452 55582 1028
rect 56566 452 56600 1028
rect 57584 452 57618 1028
rect 58602 452 58636 1028
rect 59620 452 59654 1028
rect 60638 452 60672 1028
rect 61656 452 61690 1028
rect 62674 452 62708 1028
rect 63692 452 63726 1028
rect 64710 452 64744 1028
rect 65728 452 65762 1028
rect 66746 452 66780 1028
rect 67764 452 67798 1028
rect 68782 452 68816 1028
rect 69800 452 69834 1028
rect 70818 452 70852 1028
rect 71836 452 71870 1028
rect 72854 452 72888 1028
rect 73872 452 73906 1028
rect 74890 452 74924 1028
<< pdiffc >>
rect 17438 27256 17472 27832
rect 18456 27256 18490 27832
rect 19474 27256 19508 27832
rect 20492 27256 20526 27832
rect 21510 27256 21544 27832
rect 22528 27256 22562 27832
rect 23546 27256 23580 27832
rect 24564 27256 24598 27832
rect 25582 27256 25616 27832
rect 26600 27256 26634 27832
rect 27618 27256 27652 27832
rect 28636 27256 28670 27832
rect 29654 27256 29688 27832
rect 30672 27256 30706 27832
rect 31690 27256 31724 27832
rect 32708 27256 32742 27832
rect 33726 27256 33760 27832
rect 17438 26120 17472 26696
rect 18456 26120 18490 26696
rect 19474 26120 19508 26696
rect 20492 26120 20526 26696
rect 21510 26120 21544 26696
rect 22528 26120 22562 26696
rect 23546 26120 23580 26696
rect 24564 26120 24598 26696
rect 25582 26120 25616 26696
rect 26600 26120 26634 26696
rect 27618 26120 27652 26696
rect 28636 26120 28670 26696
rect 29654 26120 29688 26696
rect 30672 26120 30706 26696
rect 31690 26120 31724 26696
rect 32708 26120 32742 26696
rect 33726 26120 33760 26696
rect 17438 24984 17472 25560
rect 18456 24984 18490 25560
rect 19474 24984 19508 25560
rect 20492 24984 20526 25560
rect 21510 24984 21544 25560
rect 22528 24984 22562 25560
rect 23546 24984 23580 25560
rect 24564 24984 24598 25560
rect 25582 24984 25616 25560
rect 26600 24984 26634 25560
rect 27618 24984 27652 25560
rect 28636 24984 28670 25560
rect 29654 24984 29688 25560
rect 30672 24984 30706 25560
rect 31690 24984 31724 25560
rect 32708 24984 32742 25560
rect 33726 24984 33760 25560
rect 18632 23346 18666 23922
rect 19650 23346 19684 23922
rect 20668 23346 20702 23922
rect 21686 23346 21720 23922
rect 22704 23346 22738 23922
rect 23722 23346 23756 23922
rect 24740 23346 24774 23922
rect 25758 23346 25792 23922
rect 26776 23346 26810 23922
rect 27794 23346 27828 23922
rect 28812 23346 28846 23922
rect 29830 23346 29864 23922
rect 30848 23346 30882 23922
rect 31866 23346 31900 23922
rect 32884 23346 32918 23922
rect 18632 22314 18666 22890
rect 19650 22314 19684 22890
rect 20668 22314 20702 22890
rect 21686 22314 21720 22890
rect 22704 22314 22738 22890
rect 23722 22314 23756 22890
rect 24740 22314 24774 22890
rect 25758 22314 25792 22890
rect 26776 22314 26810 22890
rect 27794 22314 27828 22890
rect 28812 22314 28846 22890
rect 29830 22314 29864 22890
rect 30848 22314 30882 22890
rect 31866 22314 31900 22890
rect 32884 22314 32918 22890
rect 13120 20606 13154 21182
rect 14138 20606 14172 21182
rect 15156 20606 15190 21182
rect 16174 20606 16208 21182
rect 17192 20606 17226 21182
rect 18424 20710 18458 21286
rect 19442 20710 19476 21286
rect 20460 20710 20494 21286
rect 21478 20710 21512 21286
rect 22496 20710 22530 21286
rect 23514 20710 23548 21286
rect 24532 20710 24566 21286
rect 25550 20710 25584 21286
rect 26568 20710 26602 21286
rect 27586 20710 27620 21286
rect 28604 20710 28638 21286
rect 29622 20710 29656 21286
rect 30640 20710 30674 21286
rect 31658 20710 31692 21286
rect 32676 20710 32710 21286
rect 33694 20710 33728 21286
rect 13120 19574 13154 20150
rect 14138 19574 14172 20150
rect 15156 19574 15190 20150
rect 16174 19574 16208 20150
rect 17192 19574 17226 20150
rect 18424 19454 18458 20030
rect 19442 19454 19476 20030
rect 20460 19454 20494 20030
rect 21478 19454 21512 20030
rect 22496 19454 22530 20030
rect 23514 19454 23548 20030
rect 24532 19454 24566 20030
rect 25550 19454 25584 20030
rect 26568 19454 26602 20030
rect 27586 19454 27620 20030
rect 28604 19454 28638 20030
rect 29622 19454 29656 20030
rect 30640 19454 30674 20030
rect 31658 19454 31692 20030
rect 32676 19454 32710 20030
rect 33694 19454 33728 20030
rect 13120 18542 13154 19118
rect 14138 18542 14172 19118
rect 15156 18542 15190 19118
rect 16174 18542 16208 19118
rect 17192 18542 17226 19118
rect 18424 18198 18458 18774
rect 19442 18198 19476 18774
rect 20460 18198 20494 18774
rect 21478 18198 21512 18774
rect 22496 18198 22530 18774
rect 23514 18198 23548 18774
rect 24532 18198 24566 18774
rect 25550 18198 25584 18774
rect 26568 18198 26602 18774
rect 27586 18198 27620 18774
rect 28604 18198 28638 18774
rect 29622 18198 29656 18774
rect 30640 18198 30674 18774
rect 31658 18198 31692 18774
rect 32676 18198 32710 18774
rect 33694 18198 33728 18774
rect 13120 17510 13154 18086
rect 14138 17510 14172 18086
rect 15156 17510 15190 18086
rect 16174 17510 16208 18086
rect 17192 17510 17226 18086
rect 18424 16942 18458 17518
rect 19442 16942 19476 17518
rect 20460 16942 20494 17518
rect 21478 16942 21512 17518
rect 22496 16942 22530 17518
rect 23514 16942 23548 17518
rect 24532 16942 24566 17518
rect 25550 16942 25584 17518
rect 26568 16942 26602 17518
rect 27586 16942 27620 17518
rect 28604 16942 28638 17518
rect 29622 16942 29656 17518
rect 30640 16942 30674 17518
rect 31658 16942 31692 17518
rect 32676 16942 32710 17518
rect 33694 16942 33728 17518
rect 58438 27256 58472 27832
rect 59456 27256 59490 27832
rect 60474 27256 60508 27832
rect 61492 27256 61526 27832
rect 62510 27256 62544 27832
rect 63528 27256 63562 27832
rect 64546 27256 64580 27832
rect 65564 27256 65598 27832
rect 66582 27256 66616 27832
rect 67600 27256 67634 27832
rect 68618 27256 68652 27832
rect 69636 27256 69670 27832
rect 70654 27256 70688 27832
rect 71672 27256 71706 27832
rect 72690 27256 72724 27832
rect 73708 27256 73742 27832
rect 74726 27256 74760 27832
rect 58438 26120 58472 26696
rect 59456 26120 59490 26696
rect 60474 26120 60508 26696
rect 61492 26120 61526 26696
rect 62510 26120 62544 26696
rect 63528 26120 63562 26696
rect 64546 26120 64580 26696
rect 65564 26120 65598 26696
rect 66582 26120 66616 26696
rect 67600 26120 67634 26696
rect 68618 26120 68652 26696
rect 69636 26120 69670 26696
rect 70654 26120 70688 26696
rect 71672 26120 71706 26696
rect 72690 26120 72724 26696
rect 73708 26120 73742 26696
rect 74726 26120 74760 26696
rect 58438 24984 58472 25560
rect 59456 24984 59490 25560
rect 60474 24984 60508 25560
rect 61492 24984 61526 25560
rect 62510 24984 62544 25560
rect 63528 24984 63562 25560
rect 64546 24984 64580 25560
rect 65564 24984 65598 25560
rect 66582 24984 66616 25560
rect 67600 24984 67634 25560
rect 68618 24984 68652 25560
rect 69636 24984 69670 25560
rect 70654 24984 70688 25560
rect 71672 24984 71706 25560
rect 72690 24984 72724 25560
rect 73708 24984 73742 25560
rect 74726 24984 74760 25560
rect 59632 23346 59666 23922
rect 60650 23346 60684 23922
rect 61668 23346 61702 23922
rect 62686 23346 62720 23922
rect 63704 23346 63738 23922
rect 64722 23346 64756 23922
rect 65740 23346 65774 23922
rect 66758 23346 66792 23922
rect 67776 23346 67810 23922
rect 68794 23346 68828 23922
rect 69812 23346 69846 23922
rect 70830 23346 70864 23922
rect 71848 23346 71882 23922
rect 72866 23346 72900 23922
rect 73884 23346 73918 23922
rect 59632 22314 59666 22890
rect 60650 22314 60684 22890
rect 61668 22314 61702 22890
rect 62686 22314 62720 22890
rect 63704 22314 63738 22890
rect 64722 22314 64756 22890
rect 65740 22314 65774 22890
rect 66758 22314 66792 22890
rect 67776 22314 67810 22890
rect 68794 22314 68828 22890
rect 69812 22314 69846 22890
rect 70830 22314 70864 22890
rect 71848 22314 71882 22890
rect 72866 22314 72900 22890
rect 73884 22314 73918 22890
rect 54120 20606 54154 21182
rect 55138 20606 55172 21182
rect 56156 20606 56190 21182
rect 57174 20606 57208 21182
rect 58192 20606 58226 21182
rect 59424 20710 59458 21286
rect 60442 20710 60476 21286
rect 61460 20710 61494 21286
rect 62478 20710 62512 21286
rect 63496 20710 63530 21286
rect 64514 20710 64548 21286
rect 65532 20710 65566 21286
rect 66550 20710 66584 21286
rect 67568 20710 67602 21286
rect 68586 20710 68620 21286
rect 69604 20710 69638 21286
rect 70622 20710 70656 21286
rect 71640 20710 71674 21286
rect 72658 20710 72692 21286
rect 73676 20710 73710 21286
rect 74694 20710 74728 21286
rect 54120 19574 54154 20150
rect 55138 19574 55172 20150
rect 56156 19574 56190 20150
rect 57174 19574 57208 20150
rect 58192 19574 58226 20150
rect 59424 19454 59458 20030
rect 60442 19454 60476 20030
rect 61460 19454 61494 20030
rect 62478 19454 62512 20030
rect 63496 19454 63530 20030
rect 64514 19454 64548 20030
rect 65532 19454 65566 20030
rect 66550 19454 66584 20030
rect 67568 19454 67602 20030
rect 68586 19454 68620 20030
rect 69604 19454 69638 20030
rect 70622 19454 70656 20030
rect 71640 19454 71674 20030
rect 72658 19454 72692 20030
rect 73676 19454 73710 20030
rect 74694 19454 74728 20030
rect 54120 18542 54154 19118
rect 55138 18542 55172 19118
rect 56156 18542 56190 19118
rect 57174 18542 57208 19118
rect 58192 18542 58226 19118
rect 59424 18198 59458 18774
rect 60442 18198 60476 18774
rect 61460 18198 61494 18774
rect 62478 18198 62512 18774
rect 63496 18198 63530 18774
rect 64514 18198 64548 18774
rect 65532 18198 65566 18774
rect 66550 18198 66584 18774
rect 67568 18198 67602 18774
rect 68586 18198 68620 18774
rect 69604 18198 69638 18774
rect 70622 18198 70656 18774
rect 71640 18198 71674 18774
rect 72658 18198 72692 18774
rect 73676 18198 73710 18774
rect 74694 18198 74728 18774
rect 54120 17510 54154 18086
rect 55138 17510 55172 18086
rect 56156 17510 56190 18086
rect 57174 17510 57208 18086
rect 58192 17510 58226 18086
rect 59424 16942 59458 17518
rect 60442 16942 60476 17518
rect 61460 16942 61494 17518
rect 62478 16942 62512 17518
rect 63496 16942 63530 17518
rect 64514 16942 64548 17518
rect 65532 16942 65566 17518
rect 66550 16942 66584 17518
rect 67568 16942 67602 17518
rect 68586 16942 68620 17518
rect 69604 16942 69638 17518
rect 70622 16942 70656 17518
rect 71640 16942 71674 17518
rect 72658 16942 72692 17518
rect 73676 16942 73710 17518
rect 74694 16942 74728 17518
rect 36910 12810 36944 12986
rect 37168 12810 37202 12986
rect 37426 12810 37460 12986
rect 37684 12810 37718 12986
rect 37942 12810 37976 12986
rect 38200 12810 38234 12986
rect 38458 12810 38492 12986
<< psubdiff >>
rect -1372 15092 -1210 15192
rect 35710 15092 35872 15192
rect -1372 15030 -1272 15092
rect 35772 15030 35872 15092
rect 14036 14586 14118 14610
rect 14036 14552 14060 14586
rect 14094 14552 14118 14586
rect 14036 14528 14118 14552
rect 15054 14586 15136 14610
rect 15054 14552 15078 14586
rect 15112 14552 15136 14586
rect 15054 14528 15136 14552
rect 16072 14586 16154 14610
rect 16072 14552 16096 14586
rect 16130 14552 16154 14586
rect 16072 14528 16154 14552
rect 17090 14586 17172 14610
rect 17090 14552 17114 14586
rect 17148 14552 17172 14586
rect 17090 14528 17172 14552
rect 18108 14586 18190 14610
rect 18108 14552 18132 14586
rect 18166 14552 18190 14586
rect 18108 14528 18190 14552
rect 19126 14586 19208 14610
rect 19126 14552 19150 14586
rect 19184 14552 19208 14586
rect 19126 14528 19208 14552
rect 20144 14586 20226 14610
rect 20144 14552 20168 14586
rect 20202 14552 20226 14586
rect 20144 14528 20226 14552
rect 21162 14586 21244 14610
rect 21162 14552 21186 14586
rect 21220 14552 21244 14586
rect 21162 14528 21244 14552
rect 22180 14586 22262 14610
rect 22180 14552 22204 14586
rect 22238 14552 22262 14586
rect 22180 14528 22262 14552
rect 23198 14586 23280 14610
rect 23198 14552 23222 14586
rect 23256 14552 23280 14586
rect 23198 14528 23280 14552
rect 24216 14586 24298 14610
rect 24216 14552 24240 14586
rect 24274 14552 24298 14586
rect 24216 14528 24298 14552
rect 25234 14586 25316 14610
rect 25234 14552 25258 14586
rect 25292 14552 25316 14586
rect 25234 14528 25316 14552
rect 26252 14586 26334 14610
rect 26252 14552 26276 14586
rect 26310 14552 26334 14586
rect 26252 14528 26334 14552
rect 27270 14586 27352 14610
rect 27270 14552 27294 14586
rect 27328 14552 27352 14586
rect 27270 14528 27352 14552
rect 28288 14586 28370 14610
rect 28288 14552 28312 14586
rect 28346 14552 28370 14586
rect 28288 14528 28370 14552
rect 29306 14586 29388 14610
rect 29306 14552 29330 14586
rect 29364 14552 29388 14586
rect 29306 14528 29388 14552
rect 30324 14586 30406 14610
rect 30324 14552 30348 14586
rect 30382 14552 30406 14586
rect 30324 14528 30406 14552
rect 31342 14586 31424 14610
rect 31342 14552 31366 14586
rect 31400 14552 31424 14586
rect 31342 14528 31424 14552
rect 32360 14586 32442 14610
rect 32360 14552 32384 14586
rect 32418 14552 32442 14586
rect 32360 14528 32442 14552
rect 33378 14586 33460 14610
rect 33378 14552 33402 14586
rect 33436 14552 33460 14586
rect 33378 14528 33460 14552
rect 1742 13984 1824 14008
rect 1742 13950 1766 13984
rect 1800 13950 1824 13984
rect 1742 13926 1824 13950
rect 2760 13984 2842 14008
rect 2760 13950 2784 13984
rect 2818 13950 2842 13984
rect 2760 13926 2842 13950
rect 3778 13984 3860 14008
rect 3778 13950 3802 13984
rect 3836 13950 3860 13984
rect 3778 13926 3860 13950
rect 4796 13984 4878 14008
rect 4796 13950 4820 13984
rect 4854 13950 4878 13984
rect 4796 13926 4878 13950
rect 5814 13984 5896 14008
rect 5814 13950 5838 13984
rect 5872 13950 5896 13984
rect 5814 13926 5896 13950
rect 6832 13984 6914 14008
rect 6832 13950 6856 13984
rect 6890 13950 6914 13984
rect 6832 13926 6914 13950
rect 7850 13984 7932 14008
rect 7850 13950 7874 13984
rect 7908 13950 7932 13984
rect 7850 13926 7932 13950
rect 8868 13984 8950 14008
rect 8868 13950 8892 13984
rect 8926 13950 8950 13984
rect 8868 13926 8950 13950
rect 9886 13984 9968 14008
rect 9886 13950 9910 13984
rect 9944 13950 9968 13984
rect 9886 13926 9968 13950
rect 10914 13984 10996 14008
rect 10914 13950 10938 13984
rect 10972 13950 10996 13984
rect 10914 13926 10996 13950
rect 1742 13166 1824 13190
rect 1742 13132 1766 13166
rect 1800 13132 1824 13166
rect 1742 13108 1824 13132
rect 2760 13166 2842 13190
rect 2760 13132 2784 13166
rect 2818 13132 2842 13166
rect 2760 13108 2842 13132
rect 3778 13166 3860 13190
rect 3778 13132 3802 13166
rect 3836 13132 3860 13166
rect 3778 13108 3860 13132
rect 4796 13166 4878 13190
rect 4796 13132 4820 13166
rect 4854 13132 4878 13166
rect 4796 13108 4878 13132
rect 5814 13166 5896 13190
rect 5814 13132 5838 13166
rect 5872 13132 5896 13166
rect 5814 13108 5896 13132
rect 6832 13166 6914 13190
rect 6832 13132 6856 13166
rect 6890 13132 6914 13166
rect 6832 13108 6914 13132
rect 7850 13166 7932 13190
rect 7850 13132 7874 13166
rect 7908 13132 7932 13166
rect 7850 13108 7932 13132
rect 8868 13166 8950 13190
rect 8868 13132 8892 13166
rect 8926 13132 8950 13166
rect 8868 13108 8950 13132
rect 9886 13166 9968 13190
rect 9886 13132 9910 13166
rect 9944 13132 9968 13166
rect 9886 13108 9968 13132
rect 10914 13166 10996 13190
rect 10914 13132 10938 13166
rect 10972 13132 10996 13166
rect 10914 13108 10996 13132
rect 14048 12560 14130 12584
rect 14048 12526 14072 12560
rect 14106 12526 14130 12560
rect 14048 12502 14130 12526
rect 15066 12560 15148 12584
rect 15066 12526 15090 12560
rect 15124 12526 15148 12560
rect 15066 12502 15148 12526
rect 16084 12560 16166 12584
rect 16084 12526 16108 12560
rect 16142 12526 16166 12560
rect 16084 12502 16166 12526
rect 17102 12560 17184 12584
rect 17102 12526 17126 12560
rect 17160 12526 17184 12560
rect 17102 12502 17184 12526
rect 18120 12560 18202 12584
rect 18120 12526 18144 12560
rect 18178 12526 18202 12560
rect 18120 12502 18202 12526
rect 19138 12560 19220 12584
rect 19138 12526 19162 12560
rect 19196 12526 19220 12560
rect 19138 12502 19220 12526
rect 20156 12560 20238 12584
rect 20156 12526 20180 12560
rect 20214 12526 20238 12560
rect 20156 12502 20238 12526
rect 21174 12560 21256 12584
rect 21174 12526 21198 12560
rect 21232 12526 21256 12560
rect 21174 12502 21256 12526
rect 22192 12560 22274 12584
rect 22192 12526 22216 12560
rect 22250 12526 22274 12560
rect 22192 12502 22274 12526
rect 23210 12560 23292 12584
rect 23210 12526 23234 12560
rect 23268 12526 23292 12560
rect 23210 12502 23292 12526
rect 24228 12560 24310 12584
rect 24228 12526 24252 12560
rect 24286 12526 24310 12560
rect 24228 12502 24310 12526
rect 25246 12560 25328 12584
rect 25246 12526 25270 12560
rect 25304 12526 25328 12560
rect 25246 12502 25328 12526
rect 26264 12560 26346 12584
rect 26264 12526 26288 12560
rect 26322 12526 26346 12560
rect 26264 12502 26346 12526
rect 27282 12560 27364 12584
rect 27282 12526 27306 12560
rect 27340 12526 27364 12560
rect 27282 12502 27364 12526
rect 28300 12560 28382 12584
rect 28300 12526 28324 12560
rect 28358 12526 28382 12560
rect 28300 12502 28382 12526
rect 29318 12560 29400 12584
rect 29318 12526 29342 12560
rect 29376 12526 29400 12560
rect 29318 12502 29400 12526
rect 30336 12560 30418 12584
rect 30336 12526 30360 12560
rect 30394 12526 30418 12560
rect 30336 12502 30418 12526
rect 31354 12560 31436 12584
rect 31354 12526 31378 12560
rect 31412 12526 31436 12560
rect 31354 12502 31436 12526
rect 32372 12560 32454 12584
rect 32372 12526 32396 12560
rect 32430 12526 32454 12560
rect 32372 12502 32454 12526
rect 33390 12560 33472 12584
rect 33390 12526 33414 12560
rect 33448 12526 33472 12560
rect 33390 12502 33472 12526
rect 1742 12348 1824 12372
rect 1742 12314 1766 12348
rect 1800 12314 1824 12348
rect 1742 12290 1824 12314
rect 2760 12348 2842 12372
rect 2760 12314 2784 12348
rect 2818 12314 2842 12348
rect 2760 12290 2842 12314
rect 3778 12348 3860 12372
rect 3778 12314 3802 12348
rect 3836 12314 3860 12348
rect 3778 12290 3860 12314
rect 4796 12348 4878 12372
rect 4796 12314 4820 12348
rect 4854 12314 4878 12348
rect 4796 12290 4878 12314
rect 5814 12348 5896 12372
rect 5814 12314 5838 12348
rect 5872 12314 5896 12348
rect 5814 12290 5896 12314
rect 6832 12348 6914 12372
rect 6832 12314 6856 12348
rect 6890 12314 6914 12348
rect 6832 12290 6914 12314
rect 7850 12348 7932 12372
rect 7850 12314 7874 12348
rect 7908 12314 7932 12348
rect 7850 12290 7932 12314
rect 8868 12348 8950 12372
rect 8868 12314 8892 12348
rect 8926 12314 8950 12348
rect 8868 12290 8950 12314
rect 9886 12348 9968 12372
rect 9886 12314 9910 12348
rect 9944 12314 9968 12348
rect 9886 12290 9968 12314
rect 10914 12348 10996 12372
rect 10914 12314 10938 12348
rect 10972 12314 10996 12348
rect 10914 12290 10996 12314
rect 1742 11530 1824 11554
rect 1742 11496 1766 11530
rect 1800 11496 1824 11530
rect 1742 11472 1824 11496
rect 2760 11530 2842 11554
rect 2760 11496 2784 11530
rect 2818 11496 2842 11530
rect 2760 11472 2842 11496
rect 3778 11530 3860 11554
rect 3778 11496 3802 11530
rect 3836 11496 3860 11530
rect 3778 11472 3860 11496
rect 4796 11530 4878 11554
rect 4796 11496 4820 11530
rect 4854 11496 4878 11530
rect 4796 11472 4878 11496
rect 5814 11530 5896 11554
rect 5814 11496 5838 11530
rect 5872 11496 5896 11530
rect 5814 11472 5896 11496
rect 6832 11530 6914 11554
rect 6832 11496 6856 11530
rect 6890 11496 6914 11530
rect 6832 11472 6914 11496
rect 7850 11530 7932 11554
rect 7850 11496 7874 11530
rect 7908 11496 7932 11530
rect 7850 11472 7932 11496
rect 8868 11530 8950 11554
rect 8868 11496 8892 11530
rect 8926 11496 8950 11530
rect 8868 11472 8950 11496
rect 9886 11530 9968 11554
rect 9886 11496 9910 11530
rect 9944 11496 9968 11530
rect 9886 11472 9968 11496
rect 10914 11530 10996 11554
rect 10914 11496 10938 11530
rect 10972 11496 10996 11530
rect 10914 11472 10996 11496
rect 14036 11254 14118 11278
rect 14036 11220 14060 11254
rect 14094 11220 14118 11254
rect 14036 11196 14118 11220
rect 15054 11254 15136 11278
rect 15054 11220 15078 11254
rect 15112 11220 15136 11254
rect 15054 11196 15136 11220
rect 16072 11254 16154 11278
rect 16072 11220 16096 11254
rect 16130 11220 16154 11254
rect 16072 11196 16154 11220
rect 17090 11254 17172 11278
rect 17090 11220 17114 11254
rect 17148 11220 17172 11254
rect 17090 11196 17172 11220
rect 18108 11254 18190 11278
rect 18108 11220 18132 11254
rect 18166 11220 18190 11254
rect 18108 11196 18190 11220
rect 19126 11254 19208 11278
rect 19126 11220 19150 11254
rect 19184 11220 19208 11254
rect 19126 11196 19208 11220
rect 20144 11254 20226 11278
rect 20144 11220 20168 11254
rect 20202 11220 20226 11254
rect 20144 11196 20226 11220
rect 21162 11254 21244 11278
rect 21162 11220 21186 11254
rect 21220 11220 21244 11254
rect 21162 11196 21244 11220
rect 22180 11254 22262 11278
rect 22180 11220 22204 11254
rect 22238 11220 22262 11254
rect 22180 11196 22262 11220
rect 23198 11254 23280 11278
rect 23198 11220 23222 11254
rect 23256 11220 23280 11254
rect 23198 11196 23280 11220
rect 24216 11254 24298 11278
rect 24216 11220 24240 11254
rect 24274 11220 24298 11254
rect 24216 11196 24298 11220
rect 25234 11254 25316 11278
rect 25234 11220 25258 11254
rect 25292 11220 25316 11254
rect 25234 11196 25316 11220
rect 26252 11254 26334 11278
rect 26252 11220 26276 11254
rect 26310 11220 26334 11254
rect 26252 11196 26334 11220
rect 27270 11254 27352 11278
rect 27270 11220 27294 11254
rect 27328 11220 27352 11254
rect 27270 11196 27352 11220
rect 28288 11254 28370 11278
rect 28288 11220 28312 11254
rect 28346 11220 28370 11254
rect 28288 11196 28370 11220
rect 29306 11254 29388 11278
rect 29306 11220 29330 11254
rect 29364 11220 29388 11254
rect 29306 11196 29388 11220
rect 30324 11254 30406 11278
rect 30324 11220 30348 11254
rect 30382 11220 30406 11254
rect 30324 11196 30406 11220
rect 31342 11254 31424 11278
rect 31342 11220 31366 11254
rect 31400 11220 31424 11254
rect 31342 11196 31424 11220
rect 32360 11254 32442 11278
rect 32360 11220 32384 11254
rect 32418 11220 32442 11254
rect 32360 11196 32442 11220
rect 33378 11254 33460 11278
rect 33378 11220 33402 11254
rect 33436 11220 33460 11254
rect 33378 11196 33460 11220
rect 1742 10712 1824 10736
rect 1742 10678 1766 10712
rect 1800 10678 1824 10712
rect 1742 10654 1824 10678
rect 2760 10712 2842 10736
rect 2760 10678 2784 10712
rect 2818 10678 2842 10712
rect 2760 10654 2842 10678
rect 3778 10712 3860 10736
rect 3778 10678 3802 10712
rect 3836 10678 3860 10712
rect 3778 10654 3860 10678
rect 4796 10712 4878 10736
rect 4796 10678 4820 10712
rect 4854 10678 4878 10712
rect 4796 10654 4878 10678
rect 5814 10712 5896 10736
rect 5814 10678 5838 10712
rect 5872 10678 5896 10712
rect 5814 10654 5896 10678
rect 6832 10712 6914 10736
rect 6832 10678 6856 10712
rect 6890 10678 6914 10712
rect 6832 10654 6914 10678
rect 7850 10712 7932 10736
rect 7850 10678 7874 10712
rect 7908 10678 7932 10712
rect 7850 10654 7932 10678
rect 8868 10712 8950 10736
rect 8868 10678 8892 10712
rect 8926 10678 8950 10712
rect 8868 10654 8950 10678
rect 9886 10712 9968 10736
rect 9886 10678 9910 10712
rect 9944 10678 9968 10712
rect 9886 10654 9968 10678
rect 10914 10712 10996 10736
rect 10914 10678 10938 10712
rect 10972 10678 10996 10712
rect 10914 10654 10996 10678
rect 14024 10018 14106 10042
rect 1742 9894 1824 9918
rect 1742 9860 1766 9894
rect 1800 9860 1824 9894
rect 1742 9836 1824 9860
rect 2760 9894 2842 9918
rect 2760 9860 2784 9894
rect 2818 9860 2842 9894
rect 2760 9836 2842 9860
rect 3778 9894 3860 9918
rect 3778 9860 3802 9894
rect 3836 9860 3860 9894
rect 3778 9836 3860 9860
rect 4796 9894 4878 9918
rect 4796 9860 4820 9894
rect 4854 9860 4878 9894
rect 4796 9836 4878 9860
rect 5814 9894 5896 9918
rect 5814 9860 5838 9894
rect 5872 9860 5896 9894
rect 5814 9836 5896 9860
rect 6832 9894 6914 9918
rect 6832 9860 6856 9894
rect 6890 9860 6914 9894
rect 6832 9836 6914 9860
rect 7850 9894 7932 9918
rect 7850 9860 7874 9894
rect 7908 9860 7932 9894
rect 7850 9836 7932 9860
rect 8868 9894 8950 9918
rect 14024 9984 14048 10018
rect 14082 9984 14106 10018
rect 14024 9960 14106 9984
rect 15042 10018 15124 10042
rect 15042 9984 15066 10018
rect 15100 9984 15124 10018
rect 15042 9960 15124 9984
rect 16060 10018 16142 10042
rect 16060 9984 16084 10018
rect 16118 9984 16142 10018
rect 16060 9960 16142 9984
rect 17078 10018 17160 10042
rect 17078 9984 17102 10018
rect 17136 9984 17160 10018
rect 17078 9960 17160 9984
rect 18096 10018 18178 10042
rect 18096 9984 18120 10018
rect 18154 9984 18178 10018
rect 18096 9960 18178 9984
rect 19114 10018 19196 10042
rect 19114 9984 19138 10018
rect 19172 9984 19196 10018
rect 19114 9960 19196 9984
rect 20132 10018 20214 10042
rect 20132 9984 20156 10018
rect 20190 9984 20214 10018
rect 20132 9960 20214 9984
rect 21150 10018 21232 10042
rect 21150 9984 21174 10018
rect 21208 9984 21232 10018
rect 21150 9960 21232 9984
rect 22168 10018 22250 10042
rect 22168 9984 22192 10018
rect 22226 9984 22250 10018
rect 22168 9960 22250 9984
rect 23186 10018 23268 10042
rect 23186 9984 23210 10018
rect 23244 9984 23268 10018
rect 23186 9960 23268 9984
rect 24204 10018 24286 10042
rect 24204 9984 24228 10018
rect 24262 9984 24286 10018
rect 24204 9960 24286 9984
rect 25222 10018 25304 10042
rect 25222 9984 25246 10018
rect 25280 9984 25304 10018
rect 25222 9960 25304 9984
rect 26240 10018 26322 10042
rect 26240 9984 26264 10018
rect 26298 9984 26322 10018
rect 26240 9960 26322 9984
rect 27258 10018 27340 10042
rect 27258 9984 27282 10018
rect 27316 9984 27340 10018
rect 27258 9960 27340 9984
rect 28276 10018 28358 10042
rect 28276 9984 28300 10018
rect 28334 9984 28358 10018
rect 28276 9960 28358 9984
rect 29294 10018 29376 10042
rect 29294 9984 29318 10018
rect 29352 9984 29376 10018
rect 29294 9960 29376 9984
rect 30312 10018 30394 10042
rect 30312 9984 30336 10018
rect 30370 9984 30394 10018
rect 30312 9960 30394 9984
rect 31330 10018 31412 10042
rect 31330 9984 31354 10018
rect 31388 9984 31412 10018
rect 31330 9960 31412 9984
rect 32348 10018 32430 10042
rect 32348 9984 32372 10018
rect 32406 9984 32430 10018
rect 32348 9960 32430 9984
rect 33366 10018 33448 10042
rect 33366 9984 33390 10018
rect 33424 9984 33448 10018
rect 33366 9960 33448 9984
rect 8868 9860 8892 9894
rect 8926 9860 8950 9894
rect 8868 9836 8950 9860
rect 9886 9894 9968 9918
rect 9886 9860 9910 9894
rect 9944 9860 9968 9894
rect 9886 9836 9968 9860
rect 10914 9894 10996 9918
rect 10914 9860 10938 9894
rect 10972 9860 10996 9894
rect 10914 9836 10996 9860
rect 1742 9076 1824 9100
rect 1742 9042 1766 9076
rect 1800 9042 1824 9076
rect 1742 9018 1824 9042
rect 2760 9076 2842 9100
rect 2760 9042 2784 9076
rect 2818 9042 2842 9076
rect 2760 9018 2842 9042
rect 3778 9076 3860 9100
rect 3778 9042 3802 9076
rect 3836 9042 3860 9076
rect 3778 9018 3860 9042
rect 4796 9076 4878 9100
rect 4796 9042 4820 9076
rect 4854 9042 4878 9076
rect 4796 9018 4878 9042
rect 5814 9076 5896 9100
rect 5814 9042 5838 9076
rect 5872 9042 5896 9076
rect 5814 9018 5896 9042
rect 6832 9076 6914 9100
rect 6832 9042 6856 9076
rect 6890 9042 6914 9076
rect 6832 9018 6914 9042
rect 7850 9076 7932 9100
rect 7850 9042 7874 9076
rect 7908 9042 7932 9076
rect 7850 9018 7932 9042
rect 8868 9076 8950 9100
rect 8868 9042 8892 9076
rect 8926 9042 8950 9076
rect 8868 9018 8950 9042
rect 9886 9076 9968 9100
rect 9886 9042 9910 9076
rect 9944 9042 9968 9076
rect 9886 9018 9968 9042
rect 10914 9076 10996 9100
rect 10914 9042 10938 9076
rect 10972 9042 10996 9076
rect 10914 9018 10996 9042
rect 14024 8794 14106 8818
rect 14024 8760 14048 8794
rect 14082 8760 14106 8794
rect 14024 8736 14106 8760
rect 15042 8794 15124 8818
rect 15042 8760 15066 8794
rect 15100 8760 15124 8794
rect 15042 8736 15124 8760
rect 16060 8794 16142 8818
rect 16060 8760 16084 8794
rect 16118 8760 16142 8794
rect 16060 8736 16142 8760
rect 17078 8794 17160 8818
rect 17078 8760 17102 8794
rect 17136 8760 17160 8794
rect 17078 8736 17160 8760
rect 18096 8794 18178 8818
rect 18096 8760 18120 8794
rect 18154 8760 18178 8794
rect 18096 8736 18178 8760
rect 19114 8794 19196 8818
rect 19114 8760 19138 8794
rect 19172 8760 19196 8794
rect 19114 8736 19196 8760
rect 20132 8794 20214 8818
rect 20132 8760 20156 8794
rect 20190 8760 20214 8794
rect 20132 8736 20214 8760
rect 21150 8794 21232 8818
rect 21150 8760 21174 8794
rect 21208 8760 21232 8794
rect 21150 8736 21232 8760
rect 22168 8794 22250 8818
rect 22168 8760 22192 8794
rect 22226 8760 22250 8794
rect 22168 8736 22250 8760
rect 23186 8794 23268 8818
rect 23186 8760 23210 8794
rect 23244 8760 23268 8794
rect 23186 8736 23268 8760
rect 24204 8794 24286 8818
rect 24204 8760 24228 8794
rect 24262 8760 24286 8794
rect 24204 8736 24286 8760
rect 25222 8794 25304 8818
rect 25222 8760 25246 8794
rect 25280 8760 25304 8794
rect 25222 8736 25304 8760
rect 26240 8794 26322 8818
rect 26240 8760 26264 8794
rect 26298 8760 26322 8794
rect 26240 8736 26322 8760
rect 27258 8794 27340 8818
rect 27258 8760 27282 8794
rect 27316 8760 27340 8794
rect 27258 8736 27340 8760
rect 28276 8794 28358 8818
rect 28276 8760 28300 8794
rect 28334 8760 28358 8794
rect 28276 8736 28358 8760
rect 29294 8794 29376 8818
rect 29294 8760 29318 8794
rect 29352 8760 29376 8794
rect 29294 8736 29376 8760
rect 30312 8794 30394 8818
rect 30312 8760 30336 8794
rect 30370 8760 30394 8794
rect 30312 8736 30394 8760
rect 31330 8794 31412 8818
rect 31330 8760 31354 8794
rect 31388 8760 31412 8794
rect 31330 8736 31412 8760
rect 32348 8794 32430 8818
rect 32348 8760 32372 8794
rect 32406 8760 32430 8794
rect 32348 8736 32430 8760
rect 33366 8794 33448 8818
rect 33366 8760 33390 8794
rect 33424 8760 33448 8794
rect 33366 8736 33448 8760
rect 1742 8258 1824 8282
rect 1742 8224 1766 8258
rect 1800 8224 1824 8258
rect 1742 8200 1824 8224
rect 2760 8258 2842 8282
rect 2760 8224 2784 8258
rect 2818 8224 2842 8258
rect 2760 8200 2842 8224
rect 3778 8258 3860 8282
rect 3778 8224 3802 8258
rect 3836 8224 3860 8258
rect 3778 8200 3860 8224
rect 4796 8258 4878 8282
rect 4796 8224 4820 8258
rect 4854 8224 4878 8258
rect 4796 8200 4878 8224
rect 5814 8258 5896 8282
rect 5814 8224 5838 8258
rect 5872 8224 5896 8258
rect 5814 8200 5896 8224
rect 6832 8258 6914 8282
rect 6832 8224 6856 8258
rect 6890 8224 6914 8258
rect 6832 8200 6914 8224
rect 7850 8258 7932 8282
rect 7850 8224 7874 8258
rect 7908 8224 7932 8258
rect 7850 8200 7932 8224
rect 8868 8258 8950 8282
rect 8868 8224 8892 8258
rect 8926 8224 8950 8258
rect 8868 8200 8950 8224
rect 9886 8258 9968 8282
rect 9886 8224 9910 8258
rect 9944 8224 9968 8258
rect 9886 8200 9968 8224
rect 10914 8258 10996 8282
rect 10914 8224 10938 8258
rect 10972 8224 10996 8258
rect 10914 8200 10996 8224
rect 14036 7558 14118 7582
rect 14036 7524 14060 7558
rect 14094 7524 14118 7558
rect 14036 7500 14118 7524
rect 15054 7558 15136 7582
rect 15054 7524 15078 7558
rect 15112 7524 15136 7558
rect 15054 7500 15136 7524
rect 16072 7558 16154 7582
rect 16072 7524 16096 7558
rect 16130 7524 16154 7558
rect 16072 7500 16154 7524
rect 17090 7558 17172 7582
rect 17090 7524 17114 7558
rect 17148 7524 17172 7558
rect 17090 7500 17172 7524
rect 18108 7558 18190 7582
rect 18108 7524 18132 7558
rect 18166 7524 18190 7558
rect 18108 7500 18190 7524
rect 19126 7558 19208 7582
rect 19126 7524 19150 7558
rect 19184 7524 19208 7558
rect 19126 7500 19208 7524
rect 20144 7558 20226 7582
rect 20144 7524 20168 7558
rect 20202 7524 20226 7558
rect 20144 7500 20226 7524
rect 21162 7558 21244 7582
rect 21162 7524 21186 7558
rect 21220 7524 21244 7558
rect 21162 7500 21244 7524
rect 22180 7558 22262 7582
rect 22180 7524 22204 7558
rect 22238 7524 22262 7558
rect 22180 7500 22262 7524
rect 23198 7558 23280 7582
rect 23198 7524 23222 7558
rect 23256 7524 23280 7558
rect 23198 7500 23280 7524
rect 24216 7558 24298 7582
rect 24216 7524 24240 7558
rect 24274 7524 24298 7558
rect 24216 7500 24298 7524
rect 25234 7558 25316 7582
rect 25234 7524 25258 7558
rect 25292 7524 25316 7558
rect 25234 7500 25316 7524
rect 26252 7558 26334 7582
rect 26252 7524 26276 7558
rect 26310 7524 26334 7558
rect 26252 7500 26334 7524
rect 27270 7558 27352 7582
rect 27270 7524 27294 7558
rect 27328 7524 27352 7558
rect 27270 7500 27352 7524
rect 28288 7558 28370 7582
rect 28288 7524 28312 7558
rect 28346 7524 28370 7558
rect 28288 7500 28370 7524
rect 29306 7558 29388 7582
rect 29306 7524 29330 7558
rect 29364 7524 29388 7558
rect 29306 7500 29388 7524
rect 30324 7558 30406 7582
rect 30324 7524 30348 7558
rect 30382 7524 30406 7558
rect 30324 7500 30406 7524
rect 31342 7558 31424 7582
rect 31342 7524 31366 7558
rect 31400 7524 31424 7558
rect 31342 7500 31424 7524
rect 32360 7558 32442 7582
rect 32360 7524 32384 7558
rect 32418 7524 32442 7558
rect 32360 7500 32442 7524
rect 33378 7558 33460 7582
rect 33378 7524 33402 7558
rect 33436 7524 33460 7558
rect 33378 7500 33460 7524
rect 1730 7364 1812 7388
rect 1730 7330 1754 7364
rect 1788 7330 1812 7364
rect 1730 7306 1812 7330
rect 2748 7364 2830 7388
rect 2748 7330 2772 7364
rect 2806 7330 2830 7364
rect 2748 7306 2830 7330
rect 3766 7364 3848 7388
rect 3766 7330 3790 7364
rect 3824 7330 3848 7364
rect 3766 7306 3848 7330
rect 4784 7364 4866 7388
rect 4784 7330 4808 7364
rect 4842 7330 4866 7364
rect 4784 7306 4866 7330
rect 5802 7364 5884 7388
rect 5802 7330 5826 7364
rect 5860 7330 5884 7364
rect 5802 7306 5884 7330
rect 6820 7364 6902 7388
rect 6820 7330 6844 7364
rect 6878 7330 6902 7364
rect 6820 7306 6902 7330
rect 7838 7364 7920 7388
rect 7838 7330 7862 7364
rect 7896 7330 7920 7364
rect 7838 7306 7920 7330
rect 8856 7364 8938 7388
rect 8856 7330 8880 7364
rect 8914 7330 8938 7364
rect 8856 7306 8938 7330
rect 9874 7364 9956 7388
rect 9874 7330 9898 7364
rect 9932 7330 9956 7364
rect 9874 7306 9956 7330
rect 10902 7364 10984 7388
rect 10902 7330 10926 7364
rect 10960 7330 10984 7364
rect 10902 7306 10984 7330
rect 934 6416 1016 6440
rect 934 6382 958 6416
rect 992 6382 1016 6416
rect 934 6358 1016 6382
rect 1952 6416 2034 6440
rect 1952 6382 1976 6416
rect 2010 6382 2034 6416
rect 1952 6358 2034 6382
rect 2970 6416 3052 6440
rect 2970 6382 2994 6416
rect 3028 6382 3052 6416
rect 2970 6358 3052 6382
rect 3988 6416 4070 6440
rect 3988 6382 4012 6416
rect 4046 6382 4070 6416
rect 3988 6358 4070 6382
rect 5006 6416 5088 6440
rect 5006 6382 5030 6416
rect 5064 6382 5088 6416
rect 5006 6358 5088 6382
rect 6024 6416 6106 6440
rect 6024 6382 6048 6416
rect 6082 6382 6106 6416
rect 6024 6358 6106 6382
rect 7042 6416 7124 6440
rect 7042 6382 7066 6416
rect 7100 6382 7124 6416
rect 7042 6358 7124 6382
rect 8060 6416 8142 6440
rect 8060 6382 8084 6416
rect 8118 6382 8142 6416
rect 8060 6358 8142 6382
rect 9078 6416 9160 6440
rect 9078 6382 9102 6416
rect 9136 6382 9160 6416
rect 9078 6358 9160 6382
rect 10096 6416 10178 6440
rect 10096 6382 10120 6416
rect 10154 6382 10178 6416
rect 10096 6358 10178 6382
rect 11114 6416 11196 6440
rect 11114 6382 11138 6416
rect 11172 6382 11196 6416
rect 11114 6358 11196 6382
rect 14036 6310 14118 6334
rect 14036 6276 14060 6310
rect 14094 6276 14118 6310
rect 14036 6252 14118 6276
rect 15054 6310 15136 6334
rect 15054 6276 15078 6310
rect 15112 6276 15136 6310
rect 15054 6252 15136 6276
rect 16072 6310 16154 6334
rect 16072 6276 16096 6310
rect 16130 6276 16154 6310
rect 16072 6252 16154 6276
rect 17090 6310 17172 6334
rect 17090 6276 17114 6310
rect 17148 6276 17172 6310
rect 17090 6252 17172 6276
rect 18108 6310 18190 6334
rect 18108 6276 18132 6310
rect 18166 6276 18190 6310
rect 18108 6252 18190 6276
rect 19126 6310 19208 6334
rect 19126 6276 19150 6310
rect 19184 6276 19208 6310
rect 19126 6252 19208 6276
rect 20144 6310 20226 6334
rect 20144 6276 20168 6310
rect 20202 6276 20226 6310
rect 20144 6252 20226 6276
rect 21162 6310 21244 6334
rect 21162 6276 21186 6310
rect 21220 6276 21244 6310
rect 21162 6252 21244 6276
rect 22180 6310 22262 6334
rect 22180 6276 22204 6310
rect 22238 6276 22262 6310
rect 22180 6252 22262 6276
rect 23198 6310 23280 6334
rect 23198 6276 23222 6310
rect 23256 6276 23280 6310
rect 23198 6252 23280 6276
rect 24216 6310 24298 6334
rect 24216 6276 24240 6310
rect 24274 6276 24298 6310
rect 24216 6252 24298 6276
rect 25234 6310 25316 6334
rect 25234 6276 25258 6310
rect 25292 6276 25316 6310
rect 25234 6252 25316 6276
rect 26252 6310 26334 6334
rect 26252 6276 26276 6310
rect 26310 6276 26334 6310
rect 26252 6252 26334 6276
rect 27270 6310 27352 6334
rect 27270 6276 27294 6310
rect 27328 6276 27352 6310
rect 27270 6252 27352 6276
rect 28288 6310 28370 6334
rect 28288 6276 28312 6310
rect 28346 6276 28370 6310
rect 28288 6252 28370 6276
rect 29306 6310 29388 6334
rect 29306 6276 29330 6310
rect 29364 6276 29388 6310
rect 29306 6252 29388 6276
rect 30324 6310 30406 6334
rect 30324 6276 30348 6310
rect 30382 6276 30406 6310
rect 30324 6252 30406 6276
rect 31342 6310 31424 6334
rect 31342 6276 31366 6310
rect 31400 6276 31424 6310
rect 31342 6252 31424 6276
rect 32360 6310 32442 6334
rect 32360 6276 32384 6310
rect 32418 6276 32442 6310
rect 32360 6252 32442 6276
rect 33378 6310 33460 6334
rect 33378 6276 33402 6310
rect 33436 6276 33460 6310
rect 33378 6252 33460 6276
rect 946 5274 1028 5298
rect 946 5240 970 5274
rect 1004 5240 1028 5274
rect 946 5216 1028 5240
rect 1964 5274 2046 5298
rect 1964 5240 1988 5274
rect 2022 5240 2046 5274
rect 1964 5216 2046 5240
rect 2982 5274 3064 5298
rect 2982 5240 3006 5274
rect 3040 5240 3064 5274
rect 2982 5216 3064 5240
rect 4000 5274 4082 5298
rect 4000 5240 4024 5274
rect 4058 5240 4082 5274
rect 4000 5216 4082 5240
rect 5018 5274 5100 5298
rect 5018 5240 5042 5274
rect 5076 5240 5100 5274
rect 5018 5216 5100 5240
rect 6036 5274 6118 5298
rect 6036 5240 6060 5274
rect 6094 5240 6118 5274
rect 6036 5216 6118 5240
rect 7054 5274 7136 5298
rect 7054 5240 7078 5274
rect 7112 5240 7136 5274
rect 7054 5216 7136 5240
rect 8072 5274 8154 5298
rect 8072 5240 8096 5274
rect 8130 5240 8154 5274
rect 8072 5216 8154 5240
rect 9090 5274 9172 5298
rect 9090 5240 9114 5274
rect 9148 5240 9172 5274
rect 9090 5216 9172 5240
rect 10108 5274 10190 5298
rect 10108 5240 10132 5274
rect 10166 5240 10190 5274
rect 10108 5216 10190 5240
rect 11126 5274 11208 5298
rect 11126 5240 11150 5274
rect 11184 5240 11208 5274
rect 11126 5216 11208 5240
rect 14012 5074 14094 5098
rect 14012 5040 14036 5074
rect 14070 5040 14094 5074
rect 14012 5016 14094 5040
rect 15030 5074 15112 5098
rect 15030 5040 15054 5074
rect 15088 5040 15112 5074
rect 15030 5016 15112 5040
rect 16048 5074 16130 5098
rect 16048 5040 16072 5074
rect 16106 5040 16130 5074
rect 16048 5016 16130 5040
rect 17066 5074 17148 5098
rect 17066 5040 17090 5074
rect 17124 5040 17148 5074
rect 17066 5016 17148 5040
rect 18084 5074 18166 5098
rect 18084 5040 18108 5074
rect 18142 5040 18166 5074
rect 18084 5016 18166 5040
rect 19102 5074 19184 5098
rect 19102 5040 19126 5074
rect 19160 5040 19184 5074
rect 19102 5016 19184 5040
rect 20120 5074 20202 5098
rect 20120 5040 20144 5074
rect 20178 5040 20202 5074
rect 20120 5016 20202 5040
rect 21138 5074 21220 5098
rect 21138 5040 21162 5074
rect 21196 5040 21220 5074
rect 21138 5016 21220 5040
rect 22156 5074 22238 5098
rect 22156 5040 22180 5074
rect 22214 5040 22238 5074
rect 22156 5016 22238 5040
rect 23174 5074 23256 5098
rect 23174 5040 23198 5074
rect 23232 5040 23256 5074
rect 23174 5016 23256 5040
rect 24192 5074 24274 5098
rect 24192 5040 24216 5074
rect 24250 5040 24274 5074
rect 24192 5016 24274 5040
rect 25210 5074 25292 5098
rect 25210 5040 25234 5074
rect 25268 5040 25292 5074
rect 25210 5016 25292 5040
rect 26228 5074 26310 5098
rect 26228 5040 26252 5074
rect 26286 5040 26310 5074
rect 26228 5016 26310 5040
rect 27246 5074 27328 5098
rect 27246 5040 27270 5074
rect 27304 5040 27328 5074
rect 27246 5016 27328 5040
rect 28264 5074 28346 5098
rect 28264 5040 28288 5074
rect 28322 5040 28346 5074
rect 28264 5016 28346 5040
rect 29282 5074 29364 5098
rect 29282 5040 29306 5074
rect 29340 5040 29364 5074
rect 29282 5016 29364 5040
rect 30300 5074 30382 5098
rect 30300 5040 30324 5074
rect 30358 5040 30382 5074
rect 30300 5016 30382 5040
rect 31318 5074 31400 5098
rect 31318 5040 31342 5074
rect 31376 5040 31400 5074
rect 31318 5016 31400 5040
rect 32336 5074 32418 5098
rect 32336 5040 32360 5074
rect 32394 5040 32418 5074
rect 32336 5016 32418 5040
rect 33354 5074 33436 5098
rect 33354 5040 33378 5074
rect 33412 5040 33436 5074
rect 33354 5016 33436 5040
rect 924 4166 1006 4190
rect 924 4132 948 4166
rect 982 4132 1006 4166
rect 924 4108 1006 4132
rect 1942 4166 2024 4190
rect 1942 4132 1966 4166
rect 2000 4132 2024 4166
rect 1942 4108 2024 4132
rect 2960 4166 3042 4190
rect 2960 4132 2984 4166
rect 3018 4132 3042 4166
rect 2960 4108 3042 4132
rect 3978 4166 4060 4190
rect 3978 4132 4002 4166
rect 4036 4132 4060 4166
rect 3978 4108 4060 4132
rect 4996 4166 5078 4190
rect 4996 4132 5020 4166
rect 5054 4132 5078 4166
rect 4996 4108 5078 4132
rect 6014 4166 6096 4190
rect 6014 4132 6038 4166
rect 6072 4132 6096 4166
rect 6014 4108 6096 4132
rect 7032 4166 7114 4190
rect 7032 4132 7056 4166
rect 7090 4132 7114 4166
rect 7032 4108 7114 4132
rect 8050 4166 8132 4190
rect 8050 4132 8074 4166
rect 8108 4132 8132 4166
rect 8050 4108 8132 4132
rect 9068 4166 9150 4190
rect 9068 4132 9092 4166
rect 9126 4132 9150 4166
rect 9068 4108 9150 4132
rect 10086 4166 10168 4190
rect 10086 4132 10110 4166
rect 10144 4132 10168 4166
rect 10086 4108 10168 4132
rect 11104 4166 11186 4190
rect 11104 4132 11128 4166
rect 11162 4132 11186 4166
rect 11104 4108 11186 4132
rect 14024 3850 14106 3874
rect 14024 3816 14048 3850
rect 14082 3816 14106 3850
rect 14024 3792 14106 3816
rect 15042 3850 15124 3874
rect 15042 3816 15066 3850
rect 15100 3816 15124 3850
rect 15042 3792 15124 3816
rect 16060 3850 16142 3874
rect 16060 3816 16084 3850
rect 16118 3816 16142 3850
rect 16060 3792 16142 3816
rect 17078 3850 17160 3874
rect 17078 3816 17102 3850
rect 17136 3816 17160 3850
rect 17078 3792 17160 3816
rect 18096 3850 18178 3874
rect 18096 3816 18120 3850
rect 18154 3816 18178 3850
rect 18096 3792 18178 3816
rect 19114 3850 19196 3874
rect 19114 3816 19138 3850
rect 19172 3816 19196 3850
rect 19114 3792 19196 3816
rect 20132 3850 20214 3874
rect 20132 3816 20156 3850
rect 20190 3816 20214 3850
rect 20132 3792 20214 3816
rect 21150 3850 21232 3874
rect 21150 3816 21174 3850
rect 21208 3816 21232 3850
rect 21150 3792 21232 3816
rect 22168 3850 22250 3874
rect 22168 3816 22192 3850
rect 22226 3816 22250 3850
rect 22168 3792 22250 3816
rect 23186 3850 23268 3874
rect 23186 3816 23210 3850
rect 23244 3816 23268 3850
rect 23186 3792 23268 3816
rect 24204 3850 24286 3874
rect 24204 3816 24228 3850
rect 24262 3816 24286 3850
rect 24204 3792 24286 3816
rect 25222 3850 25304 3874
rect 25222 3816 25246 3850
rect 25280 3816 25304 3850
rect 25222 3792 25304 3816
rect 26240 3850 26322 3874
rect 26240 3816 26264 3850
rect 26298 3816 26322 3850
rect 26240 3792 26322 3816
rect 27258 3850 27340 3874
rect 27258 3816 27282 3850
rect 27316 3816 27340 3850
rect 27258 3792 27340 3816
rect 28276 3850 28358 3874
rect 28276 3816 28300 3850
rect 28334 3816 28358 3850
rect 28276 3792 28358 3816
rect 29294 3850 29376 3874
rect 29294 3816 29318 3850
rect 29352 3816 29376 3850
rect 29294 3792 29376 3816
rect 30312 3850 30394 3874
rect 30312 3816 30336 3850
rect 30370 3816 30394 3850
rect 30312 3792 30394 3816
rect 31330 3850 31412 3874
rect 31330 3816 31354 3850
rect 31388 3816 31412 3850
rect 31330 3792 31412 3816
rect 32348 3850 32430 3874
rect 32348 3816 32372 3850
rect 32406 3816 32430 3850
rect 32348 3792 32430 3816
rect 33366 3850 33448 3874
rect 33366 3816 33390 3850
rect 33424 3816 33448 3850
rect 33366 3792 33448 3816
rect 924 3060 1006 3084
rect 924 3026 948 3060
rect 982 3026 1006 3060
rect 924 3002 1006 3026
rect 1942 3060 2024 3084
rect 1942 3026 1966 3060
rect 2000 3026 2024 3060
rect 1942 3002 2024 3026
rect 2960 3060 3042 3084
rect 2960 3026 2984 3060
rect 3018 3026 3042 3060
rect 2960 3002 3042 3026
rect 3978 3060 4060 3084
rect 3978 3026 4002 3060
rect 4036 3026 4060 3060
rect 3978 3002 4060 3026
rect 4996 3060 5078 3084
rect 4996 3026 5020 3060
rect 5054 3026 5078 3060
rect 4996 3002 5078 3026
rect 6014 3060 6096 3084
rect 6014 3026 6038 3060
rect 6072 3026 6096 3060
rect 6014 3002 6096 3026
rect 7032 3060 7114 3084
rect 7032 3026 7056 3060
rect 7090 3026 7114 3060
rect 7032 3002 7114 3026
rect 8050 3060 8132 3084
rect 8050 3026 8074 3060
rect 8108 3026 8132 3060
rect 8050 3002 8132 3026
rect 9068 3060 9150 3084
rect 9068 3026 9092 3060
rect 9126 3026 9150 3060
rect 9068 3002 9150 3026
rect 10086 3060 10168 3084
rect 10086 3026 10110 3060
rect 10144 3026 10168 3060
rect 10086 3002 10168 3026
rect 11104 3060 11186 3084
rect 11104 3026 11128 3060
rect 11162 3026 11186 3060
rect 11104 3002 11186 3026
rect 14024 2614 14106 2638
rect 14024 2580 14048 2614
rect 14082 2580 14106 2614
rect 14024 2556 14106 2580
rect 15042 2614 15124 2638
rect 15042 2580 15066 2614
rect 15100 2580 15124 2614
rect 15042 2556 15124 2580
rect 16060 2614 16142 2638
rect 16060 2580 16084 2614
rect 16118 2580 16142 2614
rect 16060 2556 16142 2580
rect 17078 2614 17160 2638
rect 17078 2580 17102 2614
rect 17136 2580 17160 2614
rect 17078 2556 17160 2580
rect 18096 2614 18178 2638
rect 18096 2580 18120 2614
rect 18154 2580 18178 2614
rect 18096 2556 18178 2580
rect 19114 2614 19196 2638
rect 19114 2580 19138 2614
rect 19172 2580 19196 2614
rect 19114 2556 19196 2580
rect 20132 2614 20214 2638
rect 20132 2580 20156 2614
rect 20190 2580 20214 2614
rect 20132 2556 20214 2580
rect 21150 2614 21232 2638
rect 21150 2580 21174 2614
rect 21208 2580 21232 2614
rect 21150 2556 21232 2580
rect 22168 2614 22250 2638
rect 22168 2580 22192 2614
rect 22226 2580 22250 2614
rect 22168 2556 22250 2580
rect 23186 2614 23268 2638
rect 23186 2580 23210 2614
rect 23244 2580 23268 2614
rect 23186 2556 23268 2580
rect 24204 2614 24286 2638
rect 24204 2580 24228 2614
rect 24262 2580 24286 2614
rect 24204 2556 24286 2580
rect 25222 2614 25304 2638
rect 25222 2580 25246 2614
rect 25280 2580 25304 2614
rect 25222 2556 25304 2580
rect 26240 2614 26322 2638
rect 26240 2580 26264 2614
rect 26298 2580 26322 2614
rect 26240 2556 26322 2580
rect 27258 2614 27340 2638
rect 27258 2580 27282 2614
rect 27316 2580 27340 2614
rect 27258 2556 27340 2580
rect 28276 2614 28358 2638
rect 28276 2580 28300 2614
rect 28334 2580 28358 2614
rect 28276 2556 28358 2580
rect 29294 2614 29376 2638
rect 29294 2580 29318 2614
rect 29352 2580 29376 2614
rect 29294 2556 29376 2580
rect 30312 2614 30394 2638
rect 30312 2580 30336 2614
rect 30370 2580 30394 2614
rect 30312 2556 30394 2580
rect 31330 2614 31412 2638
rect 31330 2580 31354 2614
rect 31388 2580 31412 2614
rect 31330 2556 31412 2580
rect 32348 2614 32430 2638
rect 32348 2580 32372 2614
rect 32406 2580 32430 2614
rect 32348 2556 32430 2580
rect 33366 2614 33448 2638
rect 33366 2580 33390 2614
rect 33424 2580 33448 2614
rect 33366 2556 33448 2580
rect 924 1718 1006 1742
rect 924 1684 948 1718
rect 982 1684 1006 1718
rect 924 1660 1006 1684
rect 1942 1718 2024 1742
rect 1942 1684 1966 1718
rect 2000 1684 2024 1718
rect 1942 1660 2024 1684
rect 2960 1718 3042 1742
rect 2960 1684 2984 1718
rect 3018 1684 3042 1718
rect 2960 1660 3042 1684
rect 3978 1718 4060 1742
rect 3978 1684 4002 1718
rect 4036 1684 4060 1718
rect 3978 1660 4060 1684
rect 4996 1718 5078 1742
rect 4996 1684 5020 1718
rect 5054 1684 5078 1718
rect 4996 1660 5078 1684
rect 6014 1718 6096 1742
rect 6014 1684 6038 1718
rect 6072 1684 6096 1718
rect 6014 1660 6096 1684
rect 7032 1718 7114 1742
rect 7032 1684 7056 1718
rect 7090 1684 7114 1718
rect 7032 1660 7114 1684
rect 8050 1718 8132 1742
rect 8050 1684 8074 1718
rect 8108 1684 8132 1718
rect 8050 1660 8132 1684
rect 9068 1718 9150 1742
rect 9068 1684 9092 1718
rect 9126 1684 9150 1718
rect 9068 1660 9150 1684
rect 10086 1718 10168 1742
rect 10086 1684 10110 1718
rect 10144 1684 10168 1718
rect 10086 1660 10168 1684
rect 11104 1718 11186 1742
rect 11104 1684 11128 1718
rect 11162 1684 11186 1718
rect 11104 1660 11186 1684
rect 14036 1368 14118 1392
rect 14036 1334 14060 1368
rect 14094 1334 14118 1368
rect 14036 1310 14118 1334
rect 15054 1368 15136 1392
rect 15054 1334 15078 1368
rect 15112 1334 15136 1368
rect 15054 1310 15136 1334
rect 16072 1368 16154 1392
rect 16072 1334 16096 1368
rect 16130 1334 16154 1368
rect 16072 1310 16154 1334
rect 17090 1368 17172 1392
rect 17090 1334 17114 1368
rect 17148 1334 17172 1368
rect 17090 1310 17172 1334
rect 18108 1368 18190 1392
rect 18108 1334 18132 1368
rect 18166 1334 18190 1368
rect 18108 1310 18190 1334
rect 19126 1368 19208 1392
rect 19126 1334 19150 1368
rect 19184 1334 19208 1368
rect 19126 1310 19208 1334
rect 20144 1368 20226 1392
rect 20144 1334 20168 1368
rect 20202 1334 20226 1368
rect 20144 1310 20226 1334
rect 21162 1368 21244 1392
rect 21162 1334 21186 1368
rect 21220 1334 21244 1368
rect 21162 1310 21244 1334
rect 22180 1368 22262 1392
rect 22180 1334 22204 1368
rect 22238 1334 22262 1368
rect 22180 1310 22262 1334
rect 23198 1368 23280 1392
rect 23198 1334 23222 1368
rect 23256 1334 23280 1368
rect 23198 1310 23280 1334
rect 24216 1368 24298 1392
rect 24216 1334 24240 1368
rect 24274 1334 24298 1368
rect 24216 1310 24298 1334
rect 25234 1368 25316 1392
rect 25234 1334 25258 1368
rect 25292 1334 25316 1368
rect 25234 1310 25316 1334
rect 26252 1368 26334 1392
rect 26252 1334 26276 1368
rect 26310 1334 26334 1368
rect 26252 1310 26334 1334
rect 27270 1368 27352 1392
rect 27270 1334 27294 1368
rect 27328 1334 27352 1368
rect 27270 1310 27352 1334
rect 28288 1368 28370 1392
rect 28288 1334 28312 1368
rect 28346 1334 28370 1368
rect 28288 1310 28370 1334
rect 29306 1368 29388 1392
rect 29306 1334 29330 1368
rect 29364 1334 29388 1368
rect 29306 1310 29388 1334
rect 30324 1368 30406 1392
rect 30324 1334 30348 1368
rect 30382 1334 30406 1368
rect 30324 1310 30406 1334
rect 31342 1368 31424 1392
rect 31342 1334 31366 1368
rect 31400 1334 31424 1368
rect 31342 1310 31424 1334
rect 32360 1368 32442 1392
rect 32360 1334 32384 1368
rect 32418 1334 32442 1368
rect 32360 1310 32442 1334
rect 33378 1368 33460 1392
rect 33378 1334 33402 1368
rect 33436 1334 33460 1368
rect 33378 1310 33460 1334
rect -1188 362 -1092 396
rect -934 362 -838 396
rect -1188 223 -1154 362
rect -872 223 -838 362
rect -1188 -102 -1154 51
rect 734 272 816 296
rect 734 238 758 272
rect 792 238 816 272
rect 734 214 816 238
rect 1752 272 1834 296
rect 1752 238 1776 272
rect 1810 238 1834 272
rect 1752 214 1834 238
rect 2770 272 2852 296
rect 2770 238 2794 272
rect 2828 238 2852 272
rect 2770 214 2852 238
rect 3788 272 3870 296
rect 3788 238 3812 272
rect 3846 238 3870 272
rect 3788 214 3870 238
rect 4806 272 4888 296
rect 4806 238 4830 272
rect 4864 238 4888 272
rect 4806 214 4888 238
rect 5824 272 5906 296
rect 5824 238 5848 272
rect 5882 238 5906 272
rect 5824 214 5906 238
rect 6842 272 6924 296
rect 6842 238 6866 272
rect 6900 238 6924 272
rect 6842 214 6924 238
rect 7860 272 7942 296
rect 7860 238 7884 272
rect 7918 238 7942 272
rect 7860 214 7942 238
rect 8878 272 8960 296
rect 8878 238 8902 272
rect 8936 238 8960 272
rect 8878 214 8960 238
rect 9896 272 9978 296
rect 9896 238 9920 272
rect 9954 238 9978 272
rect 9896 214 9978 238
rect 10914 272 10996 296
rect 10914 238 10938 272
rect 10972 238 10996 272
rect 10914 214 10996 238
rect 14024 190 14106 214
rect 14024 156 14048 190
rect 14082 156 14106 190
rect 14024 132 14106 156
rect 15042 190 15124 214
rect 15042 156 15066 190
rect 15100 156 15124 190
rect 15042 132 15124 156
rect 16060 190 16142 214
rect 16060 156 16084 190
rect 16118 156 16142 190
rect 16060 132 16142 156
rect 17078 190 17160 214
rect 17078 156 17102 190
rect 17136 156 17160 190
rect 17078 132 17160 156
rect 18096 190 18178 214
rect 18096 156 18120 190
rect 18154 156 18178 190
rect 18096 132 18178 156
rect 19114 190 19196 214
rect 19114 156 19138 190
rect 19172 156 19196 190
rect 19114 132 19196 156
rect 20132 190 20214 214
rect 20132 156 20156 190
rect 20190 156 20214 190
rect 20132 132 20214 156
rect 21150 190 21232 214
rect 21150 156 21174 190
rect 21208 156 21232 190
rect 21150 132 21232 156
rect 22168 190 22250 214
rect 22168 156 22192 190
rect 22226 156 22250 190
rect 22168 132 22250 156
rect 23186 190 23268 214
rect 23186 156 23210 190
rect 23244 156 23268 190
rect 23186 132 23268 156
rect 24204 190 24286 214
rect 24204 156 24228 190
rect 24262 156 24286 190
rect 24204 132 24286 156
rect 25222 190 25304 214
rect 25222 156 25246 190
rect 25280 156 25304 190
rect 25222 132 25304 156
rect 26240 190 26322 214
rect 26240 156 26264 190
rect 26298 156 26322 190
rect 26240 132 26322 156
rect 27258 190 27340 214
rect 27258 156 27282 190
rect 27316 156 27340 190
rect 27258 132 27340 156
rect 28276 190 28358 214
rect 28276 156 28300 190
rect 28334 156 28358 190
rect 28276 132 28358 156
rect 29294 190 29376 214
rect 29294 156 29318 190
rect 29352 156 29376 190
rect 29294 132 29376 156
rect 30312 190 30394 214
rect 30312 156 30336 190
rect 30370 156 30394 190
rect 30312 132 30394 156
rect 31330 190 31412 214
rect 31330 156 31354 190
rect 31388 156 31412 190
rect 31330 132 31412 156
rect 32348 190 32430 214
rect 32348 156 32372 190
rect 32406 156 32430 190
rect 32348 132 32430 156
rect 33366 190 33448 214
rect 33366 156 33390 190
rect 33424 156 33448 190
rect 33366 132 33448 156
rect -872 -102 -838 51
rect -1188 -136 -1092 -102
rect -934 -136 -838 -102
rect -1372 -752 -1272 -690
rect 39628 15092 39790 15192
rect 76710 15092 76872 15192
rect 39628 15030 39728 15092
rect 35772 -752 35872 -690
rect -1372 -852 -1210 -752
rect 35710 -852 35872 -752
rect 76772 15030 76872 15092
rect 55036 14586 55118 14610
rect 55036 14552 55060 14586
rect 55094 14552 55118 14586
rect 55036 14528 55118 14552
rect 56054 14586 56136 14610
rect 56054 14552 56078 14586
rect 56112 14552 56136 14586
rect 56054 14528 56136 14552
rect 57072 14586 57154 14610
rect 57072 14552 57096 14586
rect 57130 14552 57154 14586
rect 57072 14528 57154 14552
rect 58090 14586 58172 14610
rect 58090 14552 58114 14586
rect 58148 14552 58172 14586
rect 58090 14528 58172 14552
rect 59108 14586 59190 14610
rect 59108 14552 59132 14586
rect 59166 14552 59190 14586
rect 59108 14528 59190 14552
rect 60126 14586 60208 14610
rect 60126 14552 60150 14586
rect 60184 14552 60208 14586
rect 60126 14528 60208 14552
rect 61144 14586 61226 14610
rect 61144 14552 61168 14586
rect 61202 14552 61226 14586
rect 61144 14528 61226 14552
rect 62162 14586 62244 14610
rect 62162 14552 62186 14586
rect 62220 14552 62244 14586
rect 62162 14528 62244 14552
rect 63180 14586 63262 14610
rect 63180 14552 63204 14586
rect 63238 14552 63262 14586
rect 63180 14528 63262 14552
rect 64198 14586 64280 14610
rect 64198 14552 64222 14586
rect 64256 14552 64280 14586
rect 64198 14528 64280 14552
rect 65216 14586 65298 14610
rect 65216 14552 65240 14586
rect 65274 14552 65298 14586
rect 65216 14528 65298 14552
rect 66234 14586 66316 14610
rect 66234 14552 66258 14586
rect 66292 14552 66316 14586
rect 66234 14528 66316 14552
rect 67252 14586 67334 14610
rect 67252 14552 67276 14586
rect 67310 14552 67334 14586
rect 67252 14528 67334 14552
rect 68270 14586 68352 14610
rect 68270 14552 68294 14586
rect 68328 14552 68352 14586
rect 68270 14528 68352 14552
rect 69288 14586 69370 14610
rect 69288 14552 69312 14586
rect 69346 14552 69370 14586
rect 69288 14528 69370 14552
rect 70306 14586 70388 14610
rect 70306 14552 70330 14586
rect 70364 14552 70388 14586
rect 70306 14528 70388 14552
rect 71324 14586 71406 14610
rect 71324 14552 71348 14586
rect 71382 14552 71406 14586
rect 71324 14528 71406 14552
rect 72342 14586 72424 14610
rect 72342 14552 72366 14586
rect 72400 14552 72424 14586
rect 72342 14528 72424 14552
rect 73360 14586 73442 14610
rect 73360 14552 73384 14586
rect 73418 14552 73442 14586
rect 73360 14528 73442 14552
rect 74378 14586 74460 14610
rect 74378 14552 74402 14586
rect 74436 14552 74460 14586
rect 74378 14528 74460 14552
rect 42742 13984 42824 14008
rect 42742 13950 42766 13984
rect 42800 13950 42824 13984
rect 42742 13926 42824 13950
rect 43760 13984 43842 14008
rect 43760 13950 43784 13984
rect 43818 13950 43842 13984
rect 43760 13926 43842 13950
rect 44778 13984 44860 14008
rect 44778 13950 44802 13984
rect 44836 13950 44860 13984
rect 44778 13926 44860 13950
rect 45796 13984 45878 14008
rect 45796 13950 45820 13984
rect 45854 13950 45878 13984
rect 45796 13926 45878 13950
rect 46814 13984 46896 14008
rect 46814 13950 46838 13984
rect 46872 13950 46896 13984
rect 46814 13926 46896 13950
rect 47832 13984 47914 14008
rect 47832 13950 47856 13984
rect 47890 13950 47914 13984
rect 47832 13926 47914 13950
rect 48850 13984 48932 14008
rect 48850 13950 48874 13984
rect 48908 13950 48932 13984
rect 48850 13926 48932 13950
rect 49868 13984 49950 14008
rect 49868 13950 49892 13984
rect 49926 13950 49950 13984
rect 49868 13926 49950 13950
rect 50886 13984 50968 14008
rect 50886 13950 50910 13984
rect 50944 13950 50968 13984
rect 50886 13926 50968 13950
rect 51914 13984 51996 14008
rect 51914 13950 51938 13984
rect 51972 13950 51996 13984
rect 51914 13926 51996 13950
rect 42742 13166 42824 13190
rect 42742 13132 42766 13166
rect 42800 13132 42824 13166
rect 42742 13108 42824 13132
rect 43760 13166 43842 13190
rect 43760 13132 43784 13166
rect 43818 13132 43842 13166
rect 43760 13108 43842 13132
rect 44778 13166 44860 13190
rect 44778 13132 44802 13166
rect 44836 13132 44860 13166
rect 44778 13108 44860 13132
rect 45796 13166 45878 13190
rect 45796 13132 45820 13166
rect 45854 13132 45878 13166
rect 45796 13108 45878 13132
rect 46814 13166 46896 13190
rect 46814 13132 46838 13166
rect 46872 13132 46896 13166
rect 46814 13108 46896 13132
rect 47832 13166 47914 13190
rect 47832 13132 47856 13166
rect 47890 13132 47914 13166
rect 47832 13108 47914 13132
rect 48850 13166 48932 13190
rect 48850 13132 48874 13166
rect 48908 13132 48932 13166
rect 48850 13108 48932 13132
rect 49868 13166 49950 13190
rect 49868 13132 49892 13166
rect 49926 13132 49950 13166
rect 49868 13108 49950 13132
rect 50886 13166 50968 13190
rect 50886 13132 50910 13166
rect 50944 13132 50968 13166
rect 50886 13108 50968 13132
rect 51914 13166 51996 13190
rect 51914 13132 51938 13166
rect 51972 13132 51996 13166
rect 51914 13108 51996 13132
rect 55048 12560 55130 12584
rect 55048 12526 55072 12560
rect 55106 12526 55130 12560
rect 55048 12502 55130 12526
rect 56066 12560 56148 12584
rect 56066 12526 56090 12560
rect 56124 12526 56148 12560
rect 56066 12502 56148 12526
rect 57084 12560 57166 12584
rect 57084 12526 57108 12560
rect 57142 12526 57166 12560
rect 57084 12502 57166 12526
rect 58102 12560 58184 12584
rect 58102 12526 58126 12560
rect 58160 12526 58184 12560
rect 58102 12502 58184 12526
rect 59120 12560 59202 12584
rect 59120 12526 59144 12560
rect 59178 12526 59202 12560
rect 59120 12502 59202 12526
rect 60138 12560 60220 12584
rect 60138 12526 60162 12560
rect 60196 12526 60220 12560
rect 60138 12502 60220 12526
rect 61156 12560 61238 12584
rect 61156 12526 61180 12560
rect 61214 12526 61238 12560
rect 61156 12502 61238 12526
rect 62174 12560 62256 12584
rect 62174 12526 62198 12560
rect 62232 12526 62256 12560
rect 62174 12502 62256 12526
rect 63192 12560 63274 12584
rect 63192 12526 63216 12560
rect 63250 12526 63274 12560
rect 63192 12502 63274 12526
rect 64210 12560 64292 12584
rect 64210 12526 64234 12560
rect 64268 12526 64292 12560
rect 64210 12502 64292 12526
rect 65228 12560 65310 12584
rect 65228 12526 65252 12560
rect 65286 12526 65310 12560
rect 65228 12502 65310 12526
rect 66246 12560 66328 12584
rect 66246 12526 66270 12560
rect 66304 12526 66328 12560
rect 66246 12502 66328 12526
rect 67264 12560 67346 12584
rect 67264 12526 67288 12560
rect 67322 12526 67346 12560
rect 67264 12502 67346 12526
rect 68282 12560 68364 12584
rect 68282 12526 68306 12560
rect 68340 12526 68364 12560
rect 68282 12502 68364 12526
rect 69300 12560 69382 12584
rect 69300 12526 69324 12560
rect 69358 12526 69382 12560
rect 69300 12502 69382 12526
rect 70318 12560 70400 12584
rect 70318 12526 70342 12560
rect 70376 12526 70400 12560
rect 70318 12502 70400 12526
rect 71336 12560 71418 12584
rect 71336 12526 71360 12560
rect 71394 12526 71418 12560
rect 71336 12502 71418 12526
rect 72354 12560 72436 12584
rect 72354 12526 72378 12560
rect 72412 12526 72436 12560
rect 72354 12502 72436 12526
rect 73372 12560 73454 12584
rect 73372 12526 73396 12560
rect 73430 12526 73454 12560
rect 73372 12502 73454 12526
rect 74390 12560 74472 12584
rect 74390 12526 74414 12560
rect 74448 12526 74472 12560
rect 74390 12502 74472 12526
rect 42742 12348 42824 12372
rect 42742 12314 42766 12348
rect 42800 12314 42824 12348
rect 42742 12290 42824 12314
rect 43760 12348 43842 12372
rect 43760 12314 43784 12348
rect 43818 12314 43842 12348
rect 43760 12290 43842 12314
rect 44778 12348 44860 12372
rect 44778 12314 44802 12348
rect 44836 12314 44860 12348
rect 44778 12290 44860 12314
rect 45796 12348 45878 12372
rect 45796 12314 45820 12348
rect 45854 12314 45878 12348
rect 45796 12290 45878 12314
rect 46814 12348 46896 12372
rect 46814 12314 46838 12348
rect 46872 12314 46896 12348
rect 46814 12290 46896 12314
rect 47832 12348 47914 12372
rect 47832 12314 47856 12348
rect 47890 12314 47914 12348
rect 47832 12290 47914 12314
rect 48850 12348 48932 12372
rect 48850 12314 48874 12348
rect 48908 12314 48932 12348
rect 48850 12290 48932 12314
rect 49868 12348 49950 12372
rect 49868 12314 49892 12348
rect 49926 12314 49950 12348
rect 49868 12290 49950 12314
rect 50886 12348 50968 12372
rect 50886 12314 50910 12348
rect 50944 12314 50968 12348
rect 50886 12290 50968 12314
rect 51914 12348 51996 12372
rect 51914 12314 51938 12348
rect 51972 12314 51996 12348
rect 51914 12290 51996 12314
rect 42742 11530 42824 11554
rect 42742 11496 42766 11530
rect 42800 11496 42824 11530
rect 42742 11472 42824 11496
rect 43760 11530 43842 11554
rect 43760 11496 43784 11530
rect 43818 11496 43842 11530
rect 43760 11472 43842 11496
rect 44778 11530 44860 11554
rect 44778 11496 44802 11530
rect 44836 11496 44860 11530
rect 44778 11472 44860 11496
rect 45796 11530 45878 11554
rect 45796 11496 45820 11530
rect 45854 11496 45878 11530
rect 45796 11472 45878 11496
rect 46814 11530 46896 11554
rect 46814 11496 46838 11530
rect 46872 11496 46896 11530
rect 46814 11472 46896 11496
rect 47832 11530 47914 11554
rect 47832 11496 47856 11530
rect 47890 11496 47914 11530
rect 47832 11472 47914 11496
rect 48850 11530 48932 11554
rect 48850 11496 48874 11530
rect 48908 11496 48932 11530
rect 48850 11472 48932 11496
rect 49868 11530 49950 11554
rect 49868 11496 49892 11530
rect 49926 11496 49950 11530
rect 49868 11472 49950 11496
rect 50886 11530 50968 11554
rect 50886 11496 50910 11530
rect 50944 11496 50968 11530
rect 50886 11472 50968 11496
rect 51914 11530 51996 11554
rect 51914 11496 51938 11530
rect 51972 11496 51996 11530
rect 51914 11472 51996 11496
rect 55036 11254 55118 11278
rect 55036 11220 55060 11254
rect 55094 11220 55118 11254
rect 55036 11196 55118 11220
rect 56054 11254 56136 11278
rect 56054 11220 56078 11254
rect 56112 11220 56136 11254
rect 56054 11196 56136 11220
rect 57072 11254 57154 11278
rect 57072 11220 57096 11254
rect 57130 11220 57154 11254
rect 57072 11196 57154 11220
rect 58090 11254 58172 11278
rect 58090 11220 58114 11254
rect 58148 11220 58172 11254
rect 58090 11196 58172 11220
rect 59108 11254 59190 11278
rect 59108 11220 59132 11254
rect 59166 11220 59190 11254
rect 59108 11196 59190 11220
rect 60126 11254 60208 11278
rect 60126 11220 60150 11254
rect 60184 11220 60208 11254
rect 60126 11196 60208 11220
rect 61144 11254 61226 11278
rect 61144 11220 61168 11254
rect 61202 11220 61226 11254
rect 61144 11196 61226 11220
rect 62162 11254 62244 11278
rect 62162 11220 62186 11254
rect 62220 11220 62244 11254
rect 62162 11196 62244 11220
rect 63180 11254 63262 11278
rect 63180 11220 63204 11254
rect 63238 11220 63262 11254
rect 63180 11196 63262 11220
rect 64198 11254 64280 11278
rect 64198 11220 64222 11254
rect 64256 11220 64280 11254
rect 64198 11196 64280 11220
rect 65216 11254 65298 11278
rect 65216 11220 65240 11254
rect 65274 11220 65298 11254
rect 65216 11196 65298 11220
rect 66234 11254 66316 11278
rect 66234 11220 66258 11254
rect 66292 11220 66316 11254
rect 66234 11196 66316 11220
rect 67252 11254 67334 11278
rect 67252 11220 67276 11254
rect 67310 11220 67334 11254
rect 67252 11196 67334 11220
rect 68270 11254 68352 11278
rect 68270 11220 68294 11254
rect 68328 11220 68352 11254
rect 68270 11196 68352 11220
rect 69288 11254 69370 11278
rect 69288 11220 69312 11254
rect 69346 11220 69370 11254
rect 69288 11196 69370 11220
rect 70306 11254 70388 11278
rect 70306 11220 70330 11254
rect 70364 11220 70388 11254
rect 70306 11196 70388 11220
rect 71324 11254 71406 11278
rect 71324 11220 71348 11254
rect 71382 11220 71406 11254
rect 71324 11196 71406 11220
rect 72342 11254 72424 11278
rect 72342 11220 72366 11254
rect 72400 11220 72424 11254
rect 72342 11196 72424 11220
rect 73360 11254 73442 11278
rect 73360 11220 73384 11254
rect 73418 11220 73442 11254
rect 73360 11196 73442 11220
rect 74378 11254 74460 11278
rect 74378 11220 74402 11254
rect 74436 11220 74460 11254
rect 74378 11196 74460 11220
rect 42742 10712 42824 10736
rect 42742 10678 42766 10712
rect 42800 10678 42824 10712
rect 42742 10654 42824 10678
rect 43760 10712 43842 10736
rect 43760 10678 43784 10712
rect 43818 10678 43842 10712
rect 43760 10654 43842 10678
rect 44778 10712 44860 10736
rect 44778 10678 44802 10712
rect 44836 10678 44860 10712
rect 44778 10654 44860 10678
rect 45796 10712 45878 10736
rect 45796 10678 45820 10712
rect 45854 10678 45878 10712
rect 45796 10654 45878 10678
rect 46814 10712 46896 10736
rect 46814 10678 46838 10712
rect 46872 10678 46896 10712
rect 46814 10654 46896 10678
rect 47832 10712 47914 10736
rect 47832 10678 47856 10712
rect 47890 10678 47914 10712
rect 47832 10654 47914 10678
rect 48850 10712 48932 10736
rect 48850 10678 48874 10712
rect 48908 10678 48932 10712
rect 48850 10654 48932 10678
rect 49868 10712 49950 10736
rect 49868 10678 49892 10712
rect 49926 10678 49950 10712
rect 49868 10654 49950 10678
rect 50886 10712 50968 10736
rect 50886 10678 50910 10712
rect 50944 10678 50968 10712
rect 50886 10654 50968 10678
rect 51914 10712 51996 10736
rect 51914 10678 51938 10712
rect 51972 10678 51996 10712
rect 51914 10654 51996 10678
rect 55024 10018 55106 10042
rect 42742 9894 42824 9918
rect 42742 9860 42766 9894
rect 42800 9860 42824 9894
rect 42742 9836 42824 9860
rect 43760 9894 43842 9918
rect 43760 9860 43784 9894
rect 43818 9860 43842 9894
rect 43760 9836 43842 9860
rect 44778 9894 44860 9918
rect 44778 9860 44802 9894
rect 44836 9860 44860 9894
rect 44778 9836 44860 9860
rect 45796 9894 45878 9918
rect 45796 9860 45820 9894
rect 45854 9860 45878 9894
rect 45796 9836 45878 9860
rect 46814 9894 46896 9918
rect 46814 9860 46838 9894
rect 46872 9860 46896 9894
rect 46814 9836 46896 9860
rect 47832 9894 47914 9918
rect 47832 9860 47856 9894
rect 47890 9860 47914 9894
rect 47832 9836 47914 9860
rect 48850 9894 48932 9918
rect 48850 9860 48874 9894
rect 48908 9860 48932 9894
rect 48850 9836 48932 9860
rect 49868 9894 49950 9918
rect 55024 9984 55048 10018
rect 55082 9984 55106 10018
rect 55024 9960 55106 9984
rect 56042 10018 56124 10042
rect 56042 9984 56066 10018
rect 56100 9984 56124 10018
rect 56042 9960 56124 9984
rect 57060 10018 57142 10042
rect 57060 9984 57084 10018
rect 57118 9984 57142 10018
rect 57060 9960 57142 9984
rect 58078 10018 58160 10042
rect 58078 9984 58102 10018
rect 58136 9984 58160 10018
rect 58078 9960 58160 9984
rect 59096 10018 59178 10042
rect 59096 9984 59120 10018
rect 59154 9984 59178 10018
rect 59096 9960 59178 9984
rect 60114 10018 60196 10042
rect 60114 9984 60138 10018
rect 60172 9984 60196 10018
rect 60114 9960 60196 9984
rect 61132 10018 61214 10042
rect 61132 9984 61156 10018
rect 61190 9984 61214 10018
rect 61132 9960 61214 9984
rect 62150 10018 62232 10042
rect 62150 9984 62174 10018
rect 62208 9984 62232 10018
rect 62150 9960 62232 9984
rect 63168 10018 63250 10042
rect 63168 9984 63192 10018
rect 63226 9984 63250 10018
rect 63168 9960 63250 9984
rect 64186 10018 64268 10042
rect 64186 9984 64210 10018
rect 64244 9984 64268 10018
rect 64186 9960 64268 9984
rect 65204 10018 65286 10042
rect 65204 9984 65228 10018
rect 65262 9984 65286 10018
rect 65204 9960 65286 9984
rect 66222 10018 66304 10042
rect 66222 9984 66246 10018
rect 66280 9984 66304 10018
rect 66222 9960 66304 9984
rect 67240 10018 67322 10042
rect 67240 9984 67264 10018
rect 67298 9984 67322 10018
rect 67240 9960 67322 9984
rect 68258 10018 68340 10042
rect 68258 9984 68282 10018
rect 68316 9984 68340 10018
rect 68258 9960 68340 9984
rect 69276 10018 69358 10042
rect 69276 9984 69300 10018
rect 69334 9984 69358 10018
rect 69276 9960 69358 9984
rect 70294 10018 70376 10042
rect 70294 9984 70318 10018
rect 70352 9984 70376 10018
rect 70294 9960 70376 9984
rect 71312 10018 71394 10042
rect 71312 9984 71336 10018
rect 71370 9984 71394 10018
rect 71312 9960 71394 9984
rect 72330 10018 72412 10042
rect 72330 9984 72354 10018
rect 72388 9984 72412 10018
rect 72330 9960 72412 9984
rect 73348 10018 73430 10042
rect 73348 9984 73372 10018
rect 73406 9984 73430 10018
rect 73348 9960 73430 9984
rect 74366 10018 74448 10042
rect 74366 9984 74390 10018
rect 74424 9984 74448 10018
rect 74366 9960 74448 9984
rect 49868 9860 49892 9894
rect 49926 9860 49950 9894
rect 49868 9836 49950 9860
rect 50886 9894 50968 9918
rect 50886 9860 50910 9894
rect 50944 9860 50968 9894
rect 50886 9836 50968 9860
rect 51914 9894 51996 9918
rect 51914 9860 51938 9894
rect 51972 9860 51996 9894
rect 51914 9836 51996 9860
rect 42742 9076 42824 9100
rect 42742 9042 42766 9076
rect 42800 9042 42824 9076
rect 42742 9018 42824 9042
rect 43760 9076 43842 9100
rect 43760 9042 43784 9076
rect 43818 9042 43842 9076
rect 43760 9018 43842 9042
rect 44778 9076 44860 9100
rect 44778 9042 44802 9076
rect 44836 9042 44860 9076
rect 44778 9018 44860 9042
rect 45796 9076 45878 9100
rect 45796 9042 45820 9076
rect 45854 9042 45878 9076
rect 45796 9018 45878 9042
rect 46814 9076 46896 9100
rect 46814 9042 46838 9076
rect 46872 9042 46896 9076
rect 46814 9018 46896 9042
rect 47832 9076 47914 9100
rect 47832 9042 47856 9076
rect 47890 9042 47914 9076
rect 47832 9018 47914 9042
rect 48850 9076 48932 9100
rect 48850 9042 48874 9076
rect 48908 9042 48932 9076
rect 48850 9018 48932 9042
rect 49868 9076 49950 9100
rect 49868 9042 49892 9076
rect 49926 9042 49950 9076
rect 49868 9018 49950 9042
rect 50886 9076 50968 9100
rect 50886 9042 50910 9076
rect 50944 9042 50968 9076
rect 50886 9018 50968 9042
rect 51914 9076 51996 9100
rect 51914 9042 51938 9076
rect 51972 9042 51996 9076
rect 51914 9018 51996 9042
rect 55024 8794 55106 8818
rect 55024 8760 55048 8794
rect 55082 8760 55106 8794
rect 55024 8736 55106 8760
rect 56042 8794 56124 8818
rect 56042 8760 56066 8794
rect 56100 8760 56124 8794
rect 56042 8736 56124 8760
rect 57060 8794 57142 8818
rect 57060 8760 57084 8794
rect 57118 8760 57142 8794
rect 57060 8736 57142 8760
rect 58078 8794 58160 8818
rect 58078 8760 58102 8794
rect 58136 8760 58160 8794
rect 58078 8736 58160 8760
rect 59096 8794 59178 8818
rect 59096 8760 59120 8794
rect 59154 8760 59178 8794
rect 59096 8736 59178 8760
rect 60114 8794 60196 8818
rect 60114 8760 60138 8794
rect 60172 8760 60196 8794
rect 60114 8736 60196 8760
rect 61132 8794 61214 8818
rect 61132 8760 61156 8794
rect 61190 8760 61214 8794
rect 61132 8736 61214 8760
rect 62150 8794 62232 8818
rect 62150 8760 62174 8794
rect 62208 8760 62232 8794
rect 62150 8736 62232 8760
rect 63168 8794 63250 8818
rect 63168 8760 63192 8794
rect 63226 8760 63250 8794
rect 63168 8736 63250 8760
rect 64186 8794 64268 8818
rect 64186 8760 64210 8794
rect 64244 8760 64268 8794
rect 64186 8736 64268 8760
rect 65204 8794 65286 8818
rect 65204 8760 65228 8794
rect 65262 8760 65286 8794
rect 65204 8736 65286 8760
rect 66222 8794 66304 8818
rect 66222 8760 66246 8794
rect 66280 8760 66304 8794
rect 66222 8736 66304 8760
rect 67240 8794 67322 8818
rect 67240 8760 67264 8794
rect 67298 8760 67322 8794
rect 67240 8736 67322 8760
rect 68258 8794 68340 8818
rect 68258 8760 68282 8794
rect 68316 8760 68340 8794
rect 68258 8736 68340 8760
rect 69276 8794 69358 8818
rect 69276 8760 69300 8794
rect 69334 8760 69358 8794
rect 69276 8736 69358 8760
rect 70294 8794 70376 8818
rect 70294 8760 70318 8794
rect 70352 8760 70376 8794
rect 70294 8736 70376 8760
rect 71312 8794 71394 8818
rect 71312 8760 71336 8794
rect 71370 8760 71394 8794
rect 71312 8736 71394 8760
rect 72330 8794 72412 8818
rect 72330 8760 72354 8794
rect 72388 8760 72412 8794
rect 72330 8736 72412 8760
rect 73348 8794 73430 8818
rect 73348 8760 73372 8794
rect 73406 8760 73430 8794
rect 73348 8736 73430 8760
rect 74366 8794 74448 8818
rect 74366 8760 74390 8794
rect 74424 8760 74448 8794
rect 74366 8736 74448 8760
rect 42742 8258 42824 8282
rect 42742 8224 42766 8258
rect 42800 8224 42824 8258
rect 42742 8200 42824 8224
rect 43760 8258 43842 8282
rect 43760 8224 43784 8258
rect 43818 8224 43842 8258
rect 43760 8200 43842 8224
rect 44778 8258 44860 8282
rect 44778 8224 44802 8258
rect 44836 8224 44860 8258
rect 44778 8200 44860 8224
rect 45796 8258 45878 8282
rect 45796 8224 45820 8258
rect 45854 8224 45878 8258
rect 45796 8200 45878 8224
rect 46814 8258 46896 8282
rect 46814 8224 46838 8258
rect 46872 8224 46896 8258
rect 46814 8200 46896 8224
rect 47832 8258 47914 8282
rect 47832 8224 47856 8258
rect 47890 8224 47914 8258
rect 47832 8200 47914 8224
rect 48850 8258 48932 8282
rect 48850 8224 48874 8258
rect 48908 8224 48932 8258
rect 48850 8200 48932 8224
rect 49868 8258 49950 8282
rect 49868 8224 49892 8258
rect 49926 8224 49950 8258
rect 49868 8200 49950 8224
rect 50886 8258 50968 8282
rect 50886 8224 50910 8258
rect 50944 8224 50968 8258
rect 50886 8200 50968 8224
rect 51914 8258 51996 8282
rect 51914 8224 51938 8258
rect 51972 8224 51996 8258
rect 51914 8200 51996 8224
rect 55036 7558 55118 7582
rect 55036 7524 55060 7558
rect 55094 7524 55118 7558
rect 55036 7500 55118 7524
rect 56054 7558 56136 7582
rect 56054 7524 56078 7558
rect 56112 7524 56136 7558
rect 56054 7500 56136 7524
rect 57072 7558 57154 7582
rect 57072 7524 57096 7558
rect 57130 7524 57154 7558
rect 57072 7500 57154 7524
rect 58090 7558 58172 7582
rect 58090 7524 58114 7558
rect 58148 7524 58172 7558
rect 58090 7500 58172 7524
rect 59108 7558 59190 7582
rect 59108 7524 59132 7558
rect 59166 7524 59190 7558
rect 59108 7500 59190 7524
rect 60126 7558 60208 7582
rect 60126 7524 60150 7558
rect 60184 7524 60208 7558
rect 60126 7500 60208 7524
rect 61144 7558 61226 7582
rect 61144 7524 61168 7558
rect 61202 7524 61226 7558
rect 61144 7500 61226 7524
rect 62162 7558 62244 7582
rect 62162 7524 62186 7558
rect 62220 7524 62244 7558
rect 62162 7500 62244 7524
rect 63180 7558 63262 7582
rect 63180 7524 63204 7558
rect 63238 7524 63262 7558
rect 63180 7500 63262 7524
rect 64198 7558 64280 7582
rect 64198 7524 64222 7558
rect 64256 7524 64280 7558
rect 64198 7500 64280 7524
rect 65216 7558 65298 7582
rect 65216 7524 65240 7558
rect 65274 7524 65298 7558
rect 65216 7500 65298 7524
rect 66234 7558 66316 7582
rect 66234 7524 66258 7558
rect 66292 7524 66316 7558
rect 66234 7500 66316 7524
rect 67252 7558 67334 7582
rect 67252 7524 67276 7558
rect 67310 7524 67334 7558
rect 67252 7500 67334 7524
rect 68270 7558 68352 7582
rect 68270 7524 68294 7558
rect 68328 7524 68352 7558
rect 68270 7500 68352 7524
rect 69288 7558 69370 7582
rect 69288 7524 69312 7558
rect 69346 7524 69370 7558
rect 69288 7500 69370 7524
rect 70306 7558 70388 7582
rect 70306 7524 70330 7558
rect 70364 7524 70388 7558
rect 70306 7500 70388 7524
rect 71324 7558 71406 7582
rect 71324 7524 71348 7558
rect 71382 7524 71406 7558
rect 71324 7500 71406 7524
rect 72342 7558 72424 7582
rect 72342 7524 72366 7558
rect 72400 7524 72424 7558
rect 72342 7500 72424 7524
rect 73360 7558 73442 7582
rect 73360 7524 73384 7558
rect 73418 7524 73442 7558
rect 73360 7500 73442 7524
rect 74378 7558 74460 7582
rect 74378 7524 74402 7558
rect 74436 7524 74460 7558
rect 74378 7500 74460 7524
rect 42730 7364 42812 7388
rect 42730 7330 42754 7364
rect 42788 7330 42812 7364
rect 42730 7306 42812 7330
rect 43748 7364 43830 7388
rect 43748 7330 43772 7364
rect 43806 7330 43830 7364
rect 43748 7306 43830 7330
rect 44766 7364 44848 7388
rect 44766 7330 44790 7364
rect 44824 7330 44848 7364
rect 44766 7306 44848 7330
rect 45784 7364 45866 7388
rect 45784 7330 45808 7364
rect 45842 7330 45866 7364
rect 45784 7306 45866 7330
rect 46802 7364 46884 7388
rect 46802 7330 46826 7364
rect 46860 7330 46884 7364
rect 46802 7306 46884 7330
rect 47820 7364 47902 7388
rect 47820 7330 47844 7364
rect 47878 7330 47902 7364
rect 47820 7306 47902 7330
rect 48838 7364 48920 7388
rect 48838 7330 48862 7364
rect 48896 7330 48920 7364
rect 48838 7306 48920 7330
rect 49856 7364 49938 7388
rect 49856 7330 49880 7364
rect 49914 7330 49938 7364
rect 49856 7306 49938 7330
rect 50874 7364 50956 7388
rect 50874 7330 50898 7364
rect 50932 7330 50956 7364
rect 50874 7306 50956 7330
rect 51902 7364 51984 7388
rect 51902 7330 51926 7364
rect 51960 7330 51984 7364
rect 51902 7306 51984 7330
rect 41934 6416 42016 6440
rect 41934 6382 41958 6416
rect 41992 6382 42016 6416
rect 41934 6358 42016 6382
rect 42952 6416 43034 6440
rect 42952 6382 42976 6416
rect 43010 6382 43034 6416
rect 42952 6358 43034 6382
rect 43970 6416 44052 6440
rect 43970 6382 43994 6416
rect 44028 6382 44052 6416
rect 43970 6358 44052 6382
rect 44988 6416 45070 6440
rect 44988 6382 45012 6416
rect 45046 6382 45070 6416
rect 44988 6358 45070 6382
rect 46006 6416 46088 6440
rect 46006 6382 46030 6416
rect 46064 6382 46088 6416
rect 46006 6358 46088 6382
rect 47024 6416 47106 6440
rect 47024 6382 47048 6416
rect 47082 6382 47106 6416
rect 47024 6358 47106 6382
rect 48042 6416 48124 6440
rect 48042 6382 48066 6416
rect 48100 6382 48124 6416
rect 48042 6358 48124 6382
rect 49060 6416 49142 6440
rect 49060 6382 49084 6416
rect 49118 6382 49142 6416
rect 49060 6358 49142 6382
rect 50078 6416 50160 6440
rect 50078 6382 50102 6416
rect 50136 6382 50160 6416
rect 50078 6358 50160 6382
rect 51096 6416 51178 6440
rect 51096 6382 51120 6416
rect 51154 6382 51178 6416
rect 51096 6358 51178 6382
rect 52114 6416 52196 6440
rect 52114 6382 52138 6416
rect 52172 6382 52196 6416
rect 52114 6358 52196 6382
rect 55036 6310 55118 6334
rect 55036 6276 55060 6310
rect 55094 6276 55118 6310
rect 55036 6252 55118 6276
rect 56054 6310 56136 6334
rect 56054 6276 56078 6310
rect 56112 6276 56136 6310
rect 56054 6252 56136 6276
rect 57072 6310 57154 6334
rect 57072 6276 57096 6310
rect 57130 6276 57154 6310
rect 57072 6252 57154 6276
rect 58090 6310 58172 6334
rect 58090 6276 58114 6310
rect 58148 6276 58172 6310
rect 58090 6252 58172 6276
rect 59108 6310 59190 6334
rect 59108 6276 59132 6310
rect 59166 6276 59190 6310
rect 59108 6252 59190 6276
rect 60126 6310 60208 6334
rect 60126 6276 60150 6310
rect 60184 6276 60208 6310
rect 60126 6252 60208 6276
rect 61144 6310 61226 6334
rect 61144 6276 61168 6310
rect 61202 6276 61226 6310
rect 61144 6252 61226 6276
rect 62162 6310 62244 6334
rect 62162 6276 62186 6310
rect 62220 6276 62244 6310
rect 62162 6252 62244 6276
rect 63180 6310 63262 6334
rect 63180 6276 63204 6310
rect 63238 6276 63262 6310
rect 63180 6252 63262 6276
rect 64198 6310 64280 6334
rect 64198 6276 64222 6310
rect 64256 6276 64280 6310
rect 64198 6252 64280 6276
rect 65216 6310 65298 6334
rect 65216 6276 65240 6310
rect 65274 6276 65298 6310
rect 65216 6252 65298 6276
rect 66234 6310 66316 6334
rect 66234 6276 66258 6310
rect 66292 6276 66316 6310
rect 66234 6252 66316 6276
rect 67252 6310 67334 6334
rect 67252 6276 67276 6310
rect 67310 6276 67334 6310
rect 67252 6252 67334 6276
rect 68270 6310 68352 6334
rect 68270 6276 68294 6310
rect 68328 6276 68352 6310
rect 68270 6252 68352 6276
rect 69288 6310 69370 6334
rect 69288 6276 69312 6310
rect 69346 6276 69370 6310
rect 69288 6252 69370 6276
rect 70306 6310 70388 6334
rect 70306 6276 70330 6310
rect 70364 6276 70388 6310
rect 70306 6252 70388 6276
rect 71324 6310 71406 6334
rect 71324 6276 71348 6310
rect 71382 6276 71406 6310
rect 71324 6252 71406 6276
rect 72342 6310 72424 6334
rect 72342 6276 72366 6310
rect 72400 6276 72424 6310
rect 72342 6252 72424 6276
rect 73360 6310 73442 6334
rect 73360 6276 73384 6310
rect 73418 6276 73442 6310
rect 73360 6252 73442 6276
rect 74378 6310 74460 6334
rect 74378 6276 74402 6310
rect 74436 6276 74460 6310
rect 74378 6252 74460 6276
rect 41946 5274 42028 5298
rect 41946 5240 41970 5274
rect 42004 5240 42028 5274
rect 41946 5216 42028 5240
rect 42964 5274 43046 5298
rect 42964 5240 42988 5274
rect 43022 5240 43046 5274
rect 42964 5216 43046 5240
rect 43982 5274 44064 5298
rect 43982 5240 44006 5274
rect 44040 5240 44064 5274
rect 43982 5216 44064 5240
rect 45000 5274 45082 5298
rect 45000 5240 45024 5274
rect 45058 5240 45082 5274
rect 45000 5216 45082 5240
rect 46018 5274 46100 5298
rect 46018 5240 46042 5274
rect 46076 5240 46100 5274
rect 46018 5216 46100 5240
rect 47036 5274 47118 5298
rect 47036 5240 47060 5274
rect 47094 5240 47118 5274
rect 47036 5216 47118 5240
rect 48054 5274 48136 5298
rect 48054 5240 48078 5274
rect 48112 5240 48136 5274
rect 48054 5216 48136 5240
rect 49072 5274 49154 5298
rect 49072 5240 49096 5274
rect 49130 5240 49154 5274
rect 49072 5216 49154 5240
rect 50090 5274 50172 5298
rect 50090 5240 50114 5274
rect 50148 5240 50172 5274
rect 50090 5216 50172 5240
rect 51108 5274 51190 5298
rect 51108 5240 51132 5274
rect 51166 5240 51190 5274
rect 51108 5216 51190 5240
rect 52126 5274 52208 5298
rect 52126 5240 52150 5274
rect 52184 5240 52208 5274
rect 52126 5216 52208 5240
rect 55012 5074 55094 5098
rect 55012 5040 55036 5074
rect 55070 5040 55094 5074
rect 55012 5016 55094 5040
rect 56030 5074 56112 5098
rect 56030 5040 56054 5074
rect 56088 5040 56112 5074
rect 56030 5016 56112 5040
rect 57048 5074 57130 5098
rect 57048 5040 57072 5074
rect 57106 5040 57130 5074
rect 57048 5016 57130 5040
rect 58066 5074 58148 5098
rect 58066 5040 58090 5074
rect 58124 5040 58148 5074
rect 58066 5016 58148 5040
rect 59084 5074 59166 5098
rect 59084 5040 59108 5074
rect 59142 5040 59166 5074
rect 59084 5016 59166 5040
rect 60102 5074 60184 5098
rect 60102 5040 60126 5074
rect 60160 5040 60184 5074
rect 60102 5016 60184 5040
rect 61120 5074 61202 5098
rect 61120 5040 61144 5074
rect 61178 5040 61202 5074
rect 61120 5016 61202 5040
rect 62138 5074 62220 5098
rect 62138 5040 62162 5074
rect 62196 5040 62220 5074
rect 62138 5016 62220 5040
rect 63156 5074 63238 5098
rect 63156 5040 63180 5074
rect 63214 5040 63238 5074
rect 63156 5016 63238 5040
rect 64174 5074 64256 5098
rect 64174 5040 64198 5074
rect 64232 5040 64256 5074
rect 64174 5016 64256 5040
rect 65192 5074 65274 5098
rect 65192 5040 65216 5074
rect 65250 5040 65274 5074
rect 65192 5016 65274 5040
rect 66210 5074 66292 5098
rect 66210 5040 66234 5074
rect 66268 5040 66292 5074
rect 66210 5016 66292 5040
rect 67228 5074 67310 5098
rect 67228 5040 67252 5074
rect 67286 5040 67310 5074
rect 67228 5016 67310 5040
rect 68246 5074 68328 5098
rect 68246 5040 68270 5074
rect 68304 5040 68328 5074
rect 68246 5016 68328 5040
rect 69264 5074 69346 5098
rect 69264 5040 69288 5074
rect 69322 5040 69346 5074
rect 69264 5016 69346 5040
rect 70282 5074 70364 5098
rect 70282 5040 70306 5074
rect 70340 5040 70364 5074
rect 70282 5016 70364 5040
rect 71300 5074 71382 5098
rect 71300 5040 71324 5074
rect 71358 5040 71382 5074
rect 71300 5016 71382 5040
rect 72318 5074 72400 5098
rect 72318 5040 72342 5074
rect 72376 5040 72400 5074
rect 72318 5016 72400 5040
rect 73336 5074 73418 5098
rect 73336 5040 73360 5074
rect 73394 5040 73418 5074
rect 73336 5016 73418 5040
rect 74354 5074 74436 5098
rect 74354 5040 74378 5074
rect 74412 5040 74436 5074
rect 74354 5016 74436 5040
rect 41924 4166 42006 4190
rect 41924 4132 41948 4166
rect 41982 4132 42006 4166
rect 41924 4108 42006 4132
rect 42942 4166 43024 4190
rect 42942 4132 42966 4166
rect 43000 4132 43024 4166
rect 42942 4108 43024 4132
rect 43960 4166 44042 4190
rect 43960 4132 43984 4166
rect 44018 4132 44042 4166
rect 43960 4108 44042 4132
rect 44978 4166 45060 4190
rect 44978 4132 45002 4166
rect 45036 4132 45060 4166
rect 44978 4108 45060 4132
rect 45996 4166 46078 4190
rect 45996 4132 46020 4166
rect 46054 4132 46078 4166
rect 45996 4108 46078 4132
rect 47014 4166 47096 4190
rect 47014 4132 47038 4166
rect 47072 4132 47096 4166
rect 47014 4108 47096 4132
rect 48032 4166 48114 4190
rect 48032 4132 48056 4166
rect 48090 4132 48114 4166
rect 48032 4108 48114 4132
rect 49050 4166 49132 4190
rect 49050 4132 49074 4166
rect 49108 4132 49132 4166
rect 49050 4108 49132 4132
rect 50068 4166 50150 4190
rect 50068 4132 50092 4166
rect 50126 4132 50150 4166
rect 50068 4108 50150 4132
rect 51086 4166 51168 4190
rect 51086 4132 51110 4166
rect 51144 4132 51168 4166
rect 51086 4108 51168 4132
rect 52104 4166 52186 4190
rect 52104 4132 52128 4166
rect 52162 4132 52186 4166
rect 52104 4108 52186 4132
rect 55024 3850 55106 3874
rect 55024 3816 55048 3850
rect 55082 3816 55106 3850
rect 55024 3792 55106 3816
rect 56042 3850 56124 3874
rect 56042 3816 56066 3850
rect 56100 3816 56124 3850
rect 56042 3792 56124 3816
rect 57060 3850 57142 3874
rect 57060 3816 57084 3850
rect 57118 3816 57142 3850
rect 57060 3792 57142 3816
rect 58078 3850 58160 3874
rect 58078 3816 58102 3850
rect 58136 3816 58160 3850
rect 58078 3792 58160 3816
rect 59096 3850 59178 3874
rect 59096 3816 59120 3850
rect 59154 3816 59178 3850
rect 59096 3792 59178 3816
rect 60114 3850 60196 3874
rect 60114 3816 60138 3850
rect 60172 3816 60196 3850
rect 60114 3792 60196 3816
rect 61132 3850 61214 3874
rect 61132 3816 61156 3850
rect 61190 3816 61214 3850
rect 61132 3792 61214 3816
rect 62150 3850 62232 3874
rect 62150 3816 62174 3850
rect 62208 3816 62232 3850
rect 62150 3792 62232 3816
rect 63168 3850 63250 3874
rect 63168 3816 63192 3850
rect 63226 3816 63250 3850
rect 63168 3792 63250 3816
rect 64186 3850 64268 3874
rect 64186 3816 64210 3850
rect 64244 3816 64268 3850
rect 64186 3792 64268 3816
rect 65204 3850 65286 3874
rect 65204 3816 65228 3850
rect 65262 3816 65286 3850
rect 65204 3792 65286 3816
rect 66222 3850 66304 3874
rect 66222 3816 66246 3850
rect 66280 3816 66304 3850
rect 66222 3792 66304 3816
rect 67240 3850 67322 3874
rect 67240 3816 67264 3850
rect 67298 3816 67322 3850
rect 67240 3792 67322 3816
rect 68258 3850 68340 3874
rect 68258 3816 68282 3850
rect 68316 3816 68340 3850
rect 68258 3792 68340 3816
rect 69276 3850 69358 3874
rect 69276 3816 69300 3850
rect 69334 3816 69358 3850
rect 69276 3792 69358 3816
rect 70294 3850 70376 3874
rect 70294 3816 70318 3850
rect 70352 3816 70376 3850
rect 70294 3792 70376 3816
rect 71312 3850 71394 3874
rect 71312 3816 71336 3850
rect 71370 3816 71394 3850
rect 71312 3792 71394 3816
rect 72330 3850 72412 3874
rect 72330 3816 72354 3850
rect 72388 3816 72412 3850
rect 72330 3792 72412 3816
rect 73348 3850 73430 3874
rect 73348 3816 73372 3850
rect 73406 3816 73430 3850
rect 73348 3792 73430 3816
rect 74366 3850 74448 3874
rect 74366 3816 74390 3850
rect 74424 3816 74448 3850
rect 74366 3792 74448 3816
rect 41924 3060 42006 3084
rect 41924 3026 41948 3060
rect 41982 3026 42006 3060
rect 41924 3002 42006 3026
rect 42942 3060 43024 3084
rect 42942 3026 42966 3060
rect 43000 3026 43024 3060
rect 42942 3002 43024 3026
rect 43960 3060 44042 3084
rect 43960 3026 43984 3060
rect 44018 3026 44042 3060
rect 43960 3002 44042 3026
rect 44978 3060 45060 3084
rect 44978 3026 45002 3060
rect 45036 3026 45060 3060
rect 44978 3002 45060 3026
rect 45996 3060 46078 3084
rect 45996 3026 46020 3060
rect 46054 3026 46078 3060
rect 45996 3002 46078 3026
rect 47014 3060 47096 3084
rect 47014 3026 47038 3060
rect 47072 3026 47096 3060
rect 47014 3002 47096 3026
rect 48032 3060 48114 3084
rect 48032 3026 48056 3060
rect 48090 3026 48114 3060
rect 48032 3002 48114 3026
rect 49050 3060 49132 3084
rect 49050 3026 49074 3060
rect 49108 3026 49132 3060
rect 49050 3002 49132 3026
rect 50068 3060 50150 3084
rect 50068 3026 50092 3060
rect 50126 3026 50150 3060
rect 50068 3002 50150 3026
rect 51086 3060 51168 3084
rect 51086 3026 51110 3060
rect 51144 3026 51168 3060
rect 51086 3002 51168 3026
rect 52104 3060 52186 3084
rect 52104 3026 52128 3060
rect 52162 3026 52186 3060
rect 52104 3002 52186 3026
rect 55024 2614 55106 2638
rect 55024 2580 55048 2614
rect 55082 2580 55106 2614
rect 55024 2556 55106 2580
rect 56042 2614 56124 2638
rect 56042 2580 56066 2614
rect 56100 2580 56124 2614
rect 56042 2556 56124 2580
rect 57060 2614 57142 2638
rect 57060 2580 57084 2614
rect 57118 2580 57142 2614
rect 57060 2556 57142 2580
rect 58078 2614 58160 2638
rect 58078 2580 58102 2614
rect 58136 2580 58160 2614
rect 58078 2556 58160 2580
rect 59096 2614 59178 2638
rect 59096 2580 59120 2614
rect 59154 2580 59178 2614
rect 59096 2556 59178 2580
rect 60114 2614 60196 2638
rect 60114 2580 60138 2614
rect 60172 2580 60196 2614
rect 60114 2556 60196 2580
rect 61132 2614 61214 2638
rect 61132 2580 61156 2614
rect 61190 2580 61214 2614
rect 61132 2556 61214 2580
rect 62150 2614 62232 2638
rect 62150 2580 62174 2614
rect 62208 2580 62232 2614
rect 62150 2556 62232 2580
rect 63168 2614 63250 2638
rect 63168 2580 63192 2614
rect 63226 2580 63250 2614
rect 63168 2556 63250 2580
rect 64186 2614 64268 2638
rect 64186 2580 64210 2614
rect 64244 2580 64268 2614
rect 64186 2556 64268 2580
rect 65204 2614 65286 2638
rect 65204 2580 65228 2614
rect 65262 2580 65286 2614
rect 65204 2556 65286 2580
rect 66222 2614 66304 2638
rect 66222 2580 66246 2614
rect 66280 2580 66304 2614
rect 66222 2556 66304 2580
rect 67240 2614 67322 2638
rect 67240 2580 67264 2614
rect 67298 2580 67322 2614
rect 67240 2556 67322 2580
rect 68258 2614 68340 2638
rect 68258 2580 68282 2614
rect 68316 2580 68340 2614
rect 68258 2556 68340 2580
rect 69276 2614 69358 2638
rect 69276 2580 69300 2614
rect 69334 2580 69358 2614
rect 69276 2556 69358 2580
rect 70294 2614 70376 2638
rect 70294 2580 70318 2614
rect 70352 2580 70376 2614
rect 70294 2556 70376 2580
rect 71312 2614 71394 2638
rect 71312 2580 71336 2614
rect 71370 2580 71394 2614
rect 71312 2556 71394 2580
rect 72330 2614 72412 2638
rect 72330 2580 72354 2614
rect 72388 2580 72412 2614
rect 72330 2556 72412 2580
rect 73348 2614 73430 2638
rect 73348 2580 73372 2614
rect 73406 2580 73430 2614
rect 73348 2556 73430 2580
rect 74366 2614 74448 2638
rect 74366 2580 74390 2614
rect 74424 2580 74448 2614
rect 74366 2556 74448 2580
rect 41924 1718 42006 1742
rect 41924 1684 41948 1718
rect 41982 1684 42006 1718
rect 41924 1660 42006 1684
rect 42942 1718 43024 1742
rect 42942 1684 42966 1718
rect 43000 1684 43024 1718
rect 42942 1660 43024 1684
rect 43960 1718 44042 1742
rect 43960 1684 43984 1718
rect 44018 1684 44042 1718
rect 43960 1660 44042 1684
rect 44978 1718 45060 1742
rect 44978 1684 45002 1718
rect 45036 1684 45060 1718
rect 44978 1660 45060 1684
rect 45996 1718 46078 1742
rect 45996 1684 46020 1718
rect 46054 1684 46078 1718
rect 45996 1660 46078 1684
rect 47014 1718 47096 1742
rect 47014 1684 47038 1718
rect 47072 1684 47096 1718
rect 47014 1660 47096 1684
rect 48032 1718 48114 1742
rect 48032 1684 48056 1718
rect 48090 1684 48114 1718
rect 48032 1660 48114 1684
rect 49050 1718 49132 1742
rect 49050 1684 49074 1718
rect 49108 1684 49132 1718
rect 49050 1660 49132 1684
rect 50068 1718 50150 1742
rect 50068 1684 50092 1718
rect 50126 1684 50150 1718
rect 50068 1660 50150 1684
rect 51086 1718 51168 1742
rect 51086 1684 51110 1718
rect 51144 1684 51168 1718
rect 51086 1660 51168 1684
rect 52104 1718 52186 1742
rect 52104 1684 52128 1718
rect 52162 1684 52186 1718
rect 52104 1660 52186 1684
rect 55036 1368 55118 1392
rect 55036 1334 55060 1368
rect 55094 1334 55118 1368
rect 55036 1310 55118 1334
rect 56054 1368 56136 1392
rect 56054 1334 56078 1368
rect 56112 1334 56136 1368
rect 56054 1310 56136 1334
rect 57072 1368 57154 1392
rect 57072 1334 57096 1368
rect 57130 1334 57154 1368
rect 57072 1310 57154 1334
rect 58090 1368 58172 1392
rect 58090 1334 58114 1368
rect 58148 1334 58172 1368
rect 58090 1310 58172 1334
rect 59108 1368 59190 1392
rect 59108 1334 59132 1368
rect 59166 1334 59190 1368
rect 59108 1310 59190 1334
rect 60126 1368 60208 1392
rect 60126 1334 60150 1368
rect 60184 1334 60208 1368
rect 60126 1310 60208 1334
rect 61144 1368 61226 1392
rect 61144 1334 61168 1368
rect 61202 1334 61226 1368
rect 61144 1310 61226 1334
rect 62162 1368 62244 1392
rect 62162 1334 62186 1368
rect 62220 1334 62244 1368
rect 62162 1310 62244 1334
rect 63180 1368 63262 1392
rect 63180 1334 63204 1368
rect 63238 1334 63262 1368
rect 63180 1310 63262 1334
rect 64198 1368 64280 1392
rect 64198 1334 64222 1368
rect 64256 1334 64280 1368
rect 64198 1310 64280 1334
rect 65216 1368 65298 1392
rect 65216 1334 65240 1368
rect 65274 1334 65298 1368
rect 65216 1310 65298 1334
rect 66234 1368 66316 1392
rect 66234 1334 66258 1368
rect 66292 1334 66316 1368
rect 66234 1310 66316 1334
rect 67252 1368 67334 1392
rect 67252 1334 67276 1368
rect 67310 1334 67334 1368
rect 67252 1310 67334 1334
rect 68270 1368 68352 1392
rect 68270 1334 68294 1368
rect 68328 1334 68352 1368
rect 68270 1310 68352 1334
rect 69288 1368 69370 1392
rect 69288 1334 69312 1368
rect 69346 1334 69370 1368
rect 69288 1310 69370 1334
rect 70306 1368 70388 1392
rect 70306 1334 70330 1368
rect 70364 1334 70388 1368
rect 70306 1310 70388 1334
rect 71324 1368 71406 1392
rect 71324 1334 71348 1368
rect 71382 1334 71406 1368
rect 71324 1310 71406 1334
rect 72342 1368 72424 1392
rect 72342 1334 72366 1368
rect 72400 1334 72424 1368
rect 72342 1310 72424 1334
rect 73360 1368 73442 1392
rect 73360 1334 73384 1368
rect 73418 1334 73442 1368
rect 73360 1310 73442 1334
rect 74378 1368 74460 1392
rect 74378 1334 74402 1368
rect 74436 1334 74460 1368
rect 74378 1310 74460 1334
rect 41734 272 41816 296
rect 41734 238 41758 272
rect 41792 238 41816 272
rect 41734 214 41816 238
rect 42752 272 42834 296
rect 42752 238 42776 272
rect 42810 238 42834 272
rect 42752 214 42834 238
rect 43770 272 43852 296
rect 43770 238 43794 272
rect 43828 238 43852 272
rect 43770 214 43852 238
rect 44788 272 44870 296
rect 44788 238 44812 272
rect 44846 238 44870 272
rect 44788 214 44870 238
rect 45806 272 45888 296
rect 45806 238 45830 272
rect 45864 238 45888 272
rect 45806 214 45888 238
rect 46824 272 46906 296
rect 46824 238 46848 272
rect 46882 238 46906 272
rect 46824 214 46906 238
rect 47842 272 47924 296
rect 47842 238 47866 272
rect 47900 238 47924 272
rect 47842 214 47924 238
rect 48860 272 48942 296
rect 48860 238 48884 272
rect 48918 238 48942 272
rect 48860 214 48942 238
rect 49878 272 49960 296
rect 49878 238 49902 272
rect 49936 238 49960 272
rect 49878 214 49960 238
rect 50896 272 50978 296
rect 50896 238 50920 272
rect 50954 238 50978 272
rect 50896 214 50978 238
rect 51914 272 51996 296
rect 51914 238 51938 272
rect 51972 238 51996 272
rect 51914 214 51996 238
rect 55024 190 55106 214
rect 55024 156 55048 190
rect 55082 156 55106 190
rect 55024 132 55106 156
rect 56042 190 56124 214
rect 56042 156 56066 190
rect 56100 156 56124 190
rect 56042 132 56124 156
rect 57060 190 57142 214
rect 57060 156 57084 190
rect 57118 156 57142 190
rect 57060 132 57142 156
rect 58078 190 58160 214
rect 58078 156 58102 190
rect 58136 156 58160 190
rect 58078 132 58160 156
rect 59096 190 59178 214
rect 59096 156 59120 190
rect 59154 156 59178 190
rect 59096 132 59178 156
rect 60114 190 60196 214
rect 60114 156 60138 190
rect 60172 156 60196 190
rect 60114 132 60196 156
rect 61132 190 61214 214
rect 61132 156 61156 190
rect 61190 156 61214 190
rect 61132 132 61214 156
rect 62150 190 62232 214
rect 62150 156 62174 190
rect 62208 156 62232 190
rect 62150 132 62232 156
rect 63168 190 63250 214
rect 63168 156 63192 190
rect 63226 156 63250 190
rect 63168 132 63250 156
rect 64186 190 64268 214
rect 64186 156 64210 190
rect 64244 156 64268 190
rect 64186 132 64268 156
rect 65204 190 65286 214
rect 65204 156 65228 190
rect 65262 156 65286 190
rect 65204 132 65286 156
rect 66222 190 66304 214
rect 66222 156 66246 190
rect 66280 156 66304 190
rect 66222 132 66304 156
rect 67240 190 67322 214
rect 67240 156 67264 190
rect 67298 156 67322 190
rect 67240 132 67322 156
rect 68258 190 68340 214
rect 68258 156 68282 190
rect 68316 156 68340 190
rect 68258 132 68340 156
rect 69276 190 69358 214
rect 69276 156 69300 190
rect 69334 156 69358 190
rect 69276 132 69358 156
rect 70294 190 70376 214
rect 70294 156 70318 190
rect 70352 156 70376 190
rect 70294 132 70376 156
rect 71312 190 71394 214
rect 71312 156 71336 190
rect 71370 156 71394 190
rect 71312 132 71394 156
rect 72330 190 72412 214
rect 72330 156 72354 190
rect 72388 156 72412 190
rect 72330 132 72412 156
rect 73348 190 73430 214
rect 73348 156 73372 190
rect 73406 156 73430 190
rect 73348 132 73430 156
rect 74366 190 74448 214
rect 74366 156 74390 190
rect 74424 156 74448 190
rect 74366 132 74448 156
rect 39628 -752 39728 -690
rect 76772 -752 76872 -690
rect 39628 -852 39790 -752
rect 76710 -852 76872 -752
<< nsubdiff >>
rect 11328 30592 11490 30692
rect 35610 30592 35772 30692
rect 11328 30530 11428 30592
rect 35672 30530 35772 30592
rect 17922 28148 18004 28174
rect 17922 28114 17946 28148
rect 17980 28114 18004 28148
rect 17922 28090 18004 28114
rect 18940 28148 19022 28174
rect 18940 28114 18964 28148
rect 18998 28114 19022 28148
rect 18940 28090 19022 28114
rect 19958 28148 20040 28174
rect 19958 28114 19982 28148
rect 20016 28114 20040 28148
rect 19958 28090 20040 28114
rect 20976 28148 21058 28174
rect 20976 28114 21000 28148
rect 21034 28114 21058 28148
rect 20976 28090 21058 28114
rect 21994 28148 22076 28174
rect 21994 28114 22018 28148
rect 22052 28114 22076 28148
rect 21994 28090 22076 28114
rect 23012 28148 23094 28174
rect 23012 28114 23036 28148
rect 23070 28114 23094 28148
rect 23012 28090 23094 28114
rect 24030 28148 24112 28174
rect 24030 28114 24054 28148
rect 24088 28114 24112 28148
rect 24030 28090 24112 28114
rect 25048 28148 25130 28174
rect 25048 28114 25072 28148
rect 25106 28114 25130 28148
rect 25048 28090 25130 28114
rect 26066 28148 26148 28174
rect 26066 28114 26090 28148
rect 26124 28114 26148 28148
rect 26066 28090 26148 28114
rect 27084 28148 27166 28174
rect 27084 28114 27108 28148
rect 27142 28114 27166 28148
rect 27084 28090 27166 28114
rect 28102 28148 28184 28174
rect 28102 28114 28126 28148
rect 28160 28114 28184 28148
rect 28102 28090 28184 28114
rect 29120 28148 29202 28174
rect 29120 28114 29144 28148
rect 29178 28114 29202 28148
rect 29120 28090 29202 28114
rect 30138 28148 30220 28174
rect 30138 28114 30162 28148
rect 30196 28114 30220 28148
rect 30138 28090 30220 28114
rect 31156 28148 31238 28174
rect 31156 28114 31180 28148
rect 31214 28114 31238 28148
rect 31156 28090 31238 28114
rect 32174 28148 32256 28174
rect 32174 28114 32198 28148
rect 32232 28114 32256 28148
rect 32174 28090 32256 28114
rect 33192 28148 33274 28174
rect 33192 28114 33216 28148
rect 33250 28114 33274 28148
rect 33192 28090 33274 28114
rect 17944 26994 18026 27020
rect 17944 26960 17968 26994
rect 18002 26960 18026 26994
rect 17944 26936 18026 26960
rect 18962 26994 19044 27020
rect 18962 26960 18986 26994
rect 19020 26960 19044 26994
rect 18962 26936 19044 26960
rect 19980 26994 20062 27020
rect 19980 26960 20004 26994
rect 20038 26960 20062 26994
rect 19980 26936 20062 26960
rect 20998 26994 21080 27020
rect 20998 26960 21022 26994
rect 21056 26960 21080 26994
rect 20998 26936 21080 26960
rect 22016 26994 22098 27020
rect 22016 26960 22040 26994
rect 22074 26960 22098 26994
rect 22016 26936 22098 26960
rect 23034 26994 23116 27020
rect 23034 26960 23058 26994
rect 23092 26960 23116 26994
rect 23034 26936 23116 26960
rect 24052 26994 24134 27020
rect 24052 26960 24076 26994
rect 24110 26960 24134 26994
rect 24052 26936 24134 26960
rect 25070 26994 25152 27020
rect 25070 26960 25094 26994
rect 25128 26960 25152 26994
rect 25070 26936 25152 26960
rect 26088 26994 26170 27020
rect 26088 26960 26112 26994
rect 26146 26960 26170 26994
rect 26088 26936 26170 26960
rect 27106 26994 27188 27020
rect 27106 26960 27130 26994
rect 27164 26960 27188 26994
rect 27106 26936 27188 26960
rect 28124 26994 28206 27020
rect 28124 26960 28148 26994
rect 28182 26960 28206 26994
rect 28124 26936 28206 26960
rect 29142 26994 29224 27020
rect 29142 26960 29166 26994
rect 29200 26960 29224 26994
rect 29142 26936 29224 26960
rect 30160 26994 30242 27020
rect 30160 26960 30184 26994
rect 30218 26960 30242 26994
rect 30160 26936 30242 26960
rect 31178 26994 31260 27020
rect 31178 26960 31202 26994
rect 31236 26960 31260 26994
rect 31178 26936 31260 26960
rect 32196 26994 32278 27020
rect 32196 26960 32220 26994
rect 32254 26960 32278 26994
rect 32196 26936 32278 26960
rect 33214 26994 33296 27020
rect 33214 26960 33238 26994
rect 33272 26960 33296 26994
rect 33214 26936 33296 26960
rect 17922 25862 18004 25888
rect 17922 25828 17946 25862
rect 17980 25828 18004 25862
rect 17922 25804 18004 25828
rect 18940 25862 19022 25888
rect 18940 25828 18964 25862
rect 18998 25828 19022 25862
rect 18940 25804 19022 25828
rect 19958 25862 20040 25888
rect 19958 25828 19982 25862
rect 20016 25828 20040 25862
rect 19958 25804 20040 25828
rect 20976 25862 21058 25888
rect 20976 25828 21000 25862
rect 21034 25828 21058 25862
rect 20976 25804 21058 25828
rect 21994 25862 22076 25888
rect 21994 25828 22018 25862
rect 22052 25828 22076 25862
rect 21994 25804 22076 25828
rect 23012 25862 23094 25888
rect 23012 25828 23036 25862
rect 23070 25828 23094 25862
rect 23012 25804 23094 25828
rect 24030 25862 24112 25888
rect 24030 25828 24054 25862
rect 24088 25828 24112 25862
rect 24030 25804 24112 25828
rect 25048 25862 25130 25888
rect 25048 25828 25072 25862
rect 25106 25828 25130 25862
rect 25048 25804 25130 25828
rect 26066 25862 26148 25888
rect 26066 25828 26090 25862
rect 26124 25828 26148 25862
rect 26066 25804 26148 25828
rect 27084 25862 27166 25888
rect 27084 25828 27108 25862
rect 27142 25828 27166 25862
rect 27084 25804 27166 25828
rect 28102 25862 28184 25888
rect 28102 25828 28126 25862
rect 28160 25828 28184 25862
rect 28102 25804 28184 25828
rect 29120 25862 29202 25888
rect 29120 25828 29144 25862
rect 29178 25828 29202 25862
rect 29120 25804 29202 25828
rect 30138 25862 30220 25888
rect 30138 25828 30162 25862
rect 30196 25828 30220 25862
rect 30138 25804 30220 25828
rect 31156 25862 31238 25888
rect 31156 25828 31180 25862
rect 31214 25828 31238 25862
rect 31156 25804 31238 25828
rect 32174 25862 32256 25888
rect 32174 25828 32198 25862
rect 32232 25828 32256 25862
rect 32174 25804 32256 25828
rect 33192 25862 33274 25888
rect 33192 25828 33216 25862
rect 33250 25828 33274 25862
rect 33192 25804 33274 25828
rect 17922 24480 18004 24506
rect 17922 24446 17946 24480
rect 17980 24446 18004 24480
rect 17922 24422 18004 24446
rect 18940 24480 19022 24506
rect 18940 24446 18964 24480
rect 18998 24446 19022 24480
rect 18940 24422 19022 24446
rect 19958 24480 20040 24506
rect 19958 24446 19982 24480
rect 20016 24446 20040 24480
rect 19958 24422 20040 24446
rect 20976 24480 21058 24506
rect 20976 24446 21000 24480
rect 21034 24446 21058 24480
rect 20976 24422 21058 24446
rect 21994 24480 22076 24506
rect 21994 24446 22018 24480
rect 22052 24446 22076 24480
rect 21994 24422 22076 24446
rect 23012 24480 23094 24506
rect 23012 24446 23036 24480
rect 23070 24446 23094 24480
rect 23012 24422 23094 24446
rect 24030 24480 24112 24506
rect 24030 24446 24054 24480
rect 24088 24446 24112 24480
rect 24030 24422 24112 24446
rect 25048 24480 25130 24506
rect 25048 24446 25072 24480
rect 25106 24446 25130 24480
rect 25048 24422 25130 24446
rect 26066 24480 26148 24506
rect 26066 24446 26090 24480
rect 26124 24446 26148 24480
rect 26066 24422 26148 24446
rect 27084 24480 27166 24506
rect 27084 24446 27108 24480
rect 27142 24446 27166 24480
rect 27084 24422 27166 24446
rect 28102 24480 28184 24506
rect 28102 24446 28126 24480
rect 28160 24446 28184 24480
rect 28102 24422 28184 24446
rect 29120 24480 29202 24506
rect 29120 24446 29144 24480
rect 29178 24446 29202 24480
rect 29120 24422 29202 24446
rect 30138 24480 30220 24506
rect 30138 24446 30162 24480
rect 30196 24446 30220 24480
rect 30138 24422 30220 24446
rect 31156 24480 31238 24506
rect 31156 24446 31180 24480
rect 31214 24446 31238 24480
rect 31156 24422 31238 24446
rect 32174 24480 32256 24506
rect 32174 24446 32198 24480
rect 32232 24446 32256 24480
rect 32174 24422 32256 24446
rect 33192 24480 33274 24506
rect 33192 24446 33216 24480
rect 33250 24446 33274 24480
rect 33192 24422 33274 24446
rect 18610 23132 18692 23158
rect 18610 23098 18634 23132
rect 18668 23098 18692 23132
rect 18610 23074 18692 23098
rect 19628 23132 19710 23158
rect 19628 23098 19652 23132
rect 19686 23098 19710 23132
rect 19628 23074 19710 23098
rect 20646 23132 20728 23158
rect 20646 23098 20670 23132
rect 20704 23098 20728 23132
rect 20646 23074 20728 23098
rect 21664 23132 21746 23158
rect 21664 23098 21688 23132
rect 21722 23098 21746 23132
rect 21664 23074 21746 23098
rect 22682 23132 22764 23158
rect 22682 23098 22706 23132
rect 22740 23098 22764 23132
rect 22682 23074 22764 23098
rect 23700 23132 23782 23158
rect 23700 23098 23724 23132
rect 23758 23098 23782 23132
rect 23700 23074 23782 23098
rect 24718 23132 24800 23158
rect 24718 23098 24742 23132
rect 24776 23098 24800 23132
rect 24718 23074 24800 23098
rect 25736 23132 25818 23158
rect 25736 23098 25760 23132
rect 25794 23098 25818 23132
rect 25736 23074 25818 23098
rect 26754 23132 26836 23158
rect 26754 23098 26778 23132
rect 26812 23098 26836 23132
rect 26754 23074 26836 23098
rect 27772 23132 27854 23158
rect 27772 23098 27796 23132
rect 27830 23098 27854 23132
rect 27772 23074 27854 23098
rect 28790 23132 28872 23158
rect 28790 23098 28814 23132
rect 28848 23098 28872 23132
rect 28790 23074 28872 23098
rect 29808 23132 29890 23158
rect 29808 23098 29832 23132
rect 29866 23098 29890 23132
rect 29808 23074 29890 23098
rect 30826 23132 30908 23158
rect 30826 23098 30850 23132
rect 30884 23098 30908 23132
rect 30826 23074 30908 23098
rect 31844 23132 31926 23158
rect 31844 23098 31868 23132
rect 31902 23098 31926 23132
rect 31844 23074 31926 23098
rect 32862 23132 32944 23158
rect 32862 23098 32886 23132
rect 32920 23098 32944 23132
rect 32862 23074 32944 23098
rect 18216 21854 18298 21880
rect 18216 21820 18240 21854
rect 18274 21820 18298 21854
rect 18216 21796 18298 21820
rect 19234 21854 19316 21880
rect 19234 21820 19258 21854
rect 19292 21820 19316 21854
rect 19234 21796 19316 21820
rect 20252 21854 20334 21880
rect 20252 21820 20276 21854
rect 20310 21820 20334 21854
rect 20252 21796 20334 21820
rect 21270 21854 21352 21880
rect 21270 21820 21294 21854
rect 21328 21820 21352 21854
rect 21270 21796 21352 21820
rect 22288 21854 22370 21880
rect 22288 21820 22312 21854
rect 22346 21820 22370 21854
rect 22288 21796 22370 21820
rect 23306 21854 23388 21880
rect 23306 21820 23330 21854
rect 23364 21820 23388 21854
rect 23306 21796 23388 21820
rect 24324 21854 24406 21880
rect 24324 21820 24348 21854
rect 24382 21820 24406 21854
rect 24324 21796 24406 21820
rect 25342 21854 25424 21880
rect 25342 21820 25366 21854
rect 25400 21820 25424 21854
rect 25342 21796 25424 21820
rect 26360 21854 26442 21880
rect 26360 21820 26384 21854
rect 26418 21820 26442 21854
rect 26360 21796 26442 21820
rect 27378 21854 27460 21880
rect 27378 21820 27402 21854
rect 27436 21820 27460 21854
rect 27378 21796 27460 21820
rect 28396 21854 28478 21880
rect 28396 21820 28420 21854
rect 28454 21820 28478 21854
rect 28396 21796 28478 21820
rect 29414 21854 29496 21880
rect 29414 21820 29438 21854
rect 29472 21820 29496 21854
rect 29414 21796 29496 21820
rect 30432 21854 30514 21880
rect 30432 21820 30456 21854
rect 30490 21820 30514 21854
rect 30432 21796 30514 21820
rect 31450 21854 31532 21880
rect 31450 21820 31474 21854
rect 31508 21820 31532 21854
rect 31450 21796 31532 21820
rect 32468 21854 32550 21880
rect 32468 21820 32492 21854
rect 32526 21820 32550 21854
rect 32468 21796 32550 21820
rect 33486 21854 33568 21880
rect 33486 21820 33510 21854
rect 33544 21820 33568 21854
rect 33486 21796 33568 21820
rect 13618 21544 13700 21570
rect 13618 21510 13642 21544
rect 13676 21510 13700 21544
rect 13618 21486 13700 21510
rect 14636 21544 14718 21570
rect 14636 21510 14660 21544
rect 14694 21510 14718 21544
rect 14636 21486 14718 21510
rect 15654 21544 15736 21570
rect 15654 21510 15678 21544
rect 15712 21510 15736 21544
rect 15654 21486 15736 21510
rect 16672 21544 16754 21570
rect 16672 21510 16696 21544
rect 16730 21510 16754 21544
rect 16672 21486 16754 21510
rect 13094 20390 13176 20416
rect 13094 20356 13118 20390
rect 13152 20356 13176 20390
rect 13094 20332 13176 20356
rect 14112 20390 14194 20416
rect 14112 20356 14136 20390
rect 14170 20356 14194 20390
rect 14112 20332 14194 20356
rect 15130 20390 15212 20416
rect 15130 20356 15154 20390
rect 15188 20356 15212 20390
rect 15130 20332 15212 20356
rect 16148 20390 16230 20416
rect 16148 20356 16172 20390
rect 16206 20356 16230 20390
rect 16148 20332 16230 20356
rect 18306 20406 18388 20432
rect 18306 20372 18330 20406
rect 18364 20372 18388 20406
rect 18306 20348 18388 20372
rect 19324 20406 19406 20432
rect 19324 20372 19348 20406
rect 19382 20372 19406 20406
rect 19324 20348 19406 20372
rect 20342 20406 20424 20432
rect 20342 20372 20366 20406
rect 20400 20372 20424 20406
rect 20342 20348 20424 20372
rect 21360 20406 21442 20432
rect 21360 20372 21384 20406
rect 21418 20372 21442 20406
rect 21360 20348 21442 20372
rect 22378 20406 22460 20432
rect 22378 20372 22402 20406
rect 22436 20372 22460 20406
rect 22378 20348 22460 20372
rect 23396 20406 23478 20432
rect 23396 20372 23420 20406
rect 23454 20372 23478 20406
rect 23396 20348 23478 20372
rect 24414 20406 24496 20432
rect 24414 20372 24438 20406
rect 24472 20372 24496 20406
rect 24414 20348 24496 20372
rect 25432 20406 25514 20432
rect 25432 20372 25456 20406
rect 25490 20372 25514 20406
rect 25432 20348 25514 20372
rect 26450 20406 26532 20432
rect 26450 20372 26474 20406
rect 26508 20372 26532 20406
rect 26450 20348 26532 20372
rect 27468 20406 27550 20432
rect 27468 20372 27492 20406
rect 27526 20372 27550 20406
rect 27468 20348 27550 20372
rect 28486 20406 28568 20432
rect 28486 20372 28510 20406
rect 28544 20372 28568 20406
rect 28486 20348 28568 20372
rect 29504 20406 29586 20432
rect 29504 20372 29528 20406
rect 29562 20372 29586 20406
rect 29504 20348 29586 20372
rect 30522 20406 30604 20432
rect 30522 20372 30546 20406
rect 30580 20372 30604 20406
rect 30522 20348 30604 20372
rect 31540 20406 31622 20432
rect 31540 20372 31564 20406
rect 31598 20372 31622 20406
rect 31540 20348 31622 20372
rect 32558 20406 32640 20432
rect 32558 20372 32582 20406
rect 32616 20372 32640 20406
rect 32558 20348 32640 20372
rect 33576 20406 33658 20432
rect 33576 20372 33600 20406
rect 33634 20372 33658 20406
rect 33576 20348 33658 20372
rect 13104 19362 13186 19388
rect 13104 19328 13128 19362
rect 13162 19328 13186 19362
rect 13104 19304 13186 19328
rect 14122 19362 14204 19388
rect 14122 19328 14146 19362
rect 14180 19328 14204 19362
rect 14122 19304 14204 19328
rect 15140 19362 15222 19388
rect 15140 19328 15164 19362
rect 15198 19328 15222 19362
rect 15140 19304 15222 19328
rect 16158 19362 16240 19388
rect 16158 19328 16182 19362
rect 16216 19328 16240 19362
rect 16158 19304 16240 19328
rect 18330 19138 18412 19164
rect 18330 19104 18354 19138
rect 18388 19104 18412 19138
rect 18330 19080 18412 19104
rect 19348 19138 19430 19164
rect 19348 19104 19372 19138
rect 19406 19104 19430 19138
rect 19348 19080 19430 19104
rect 20366 19138 20448 19164
rect 20366 19104 20390 19138
rect 20424 19104 20448 19138
rect 20366 19080 20448 19104
rect 21384 19138 21466 19164
rect 21384 19104 21408 19138
rect 21442 19104 21466 19138
rect 21384 19080 21466 19104
rect 22402 19138 22484 19164
rect 22402 19104 22426 19138
rect 22460 19104 22484 19138
rect 22402 19080 22484 19104
rect 23420 19138 23502 19164
rect 23420 19104 23444 19138
rect 23478 19104 23502 19138
rect 23420 19080 23502 19104
rect 24438 19138 24520 19164
rect 24438 19104 24462 19138
rect 24496 19104 24520 19138
rect 24438 19080 24520 19104
rect 25456 19138 25538 19164
rect 25456 19104 25480 19138
rect 25514 19104 25538 19138
rect 25456 19080 25538 19104
rect 26474 19138 26556 19164
rect 26474 19104 26498 19138
rect 26532 19104 26556 19138
rect 26474 19080 26556 19104
rect 27492 19138 27574 19164
rect 27492 19104 27516 19138
rect 27550 19104 27574 19138
rect 27492 19080 27574 19104
rect 28510 19138 28592 19164
rect 28510 19104 28534 19138
rect 28568 19104 28592 19138
rect 28510 19080 28592 19104
rect 29528 19138 29610 19164
rect 29528 19104 29552 19138
rect 29586 19104 29610 19138
rect 29528 19080 29610 19104
rect 30546 19138 30628 19164
rect 30546 19104 30570 19138
rect 30604 19104 30628 19138
rect 30546 19080 30628 19104
rect 31564 19138 31646 19164
rect 31564 19104 31588 19138
rect 31622 19104 31646 19138
rect 31564 19080 31646 19104
rect 32582 19138 32664 19164
rect 32582 19104 32606 19138
rect 32640 19104 32664 19138
rect 32582 19080 32664 19104
rect 33600 19138 33682 19164
rect 33600 19104 33624 19138
rect 33658 19104 33682 19138
rect 33600 19080 33682 19104
rect 13094 18334 13176 18360
rect 13094 18300 13118 18334
rect 13152 18300 13176 18334
rect 13094 18276 13176 18300
rect 14112 18334 14194 18360
rect 14112 18300 14136 18334
rect 14170 18300 14194 18334
rect 14112 18276 14194 18300
rect 15130 18334 15212 18360
rect 15130 18300 15154 18334
rect 15188 18300 15212 18334
rect 15130 18276 15212 18300
rect 16148 18334 16230 18360
rect 16148 18300 16172 18334
rect 16206 18300 16230 18334
rect 16148 18276 16230 18300
rect 18194 17894 18276 17920
rect 18194 17860 18218 17894
rect 18252 17860 18276 17894
rect 18194 17836 18276 17860
rect 19212 17894 19294 17920
rect 19212 17860 19236 17894
rect 19270 17860 19294 17894
rect 19212 17836 19294 17860
rect 20230 17894 20312 17920
rect 20230 17860 20254 17894
rect 20288 17860 20312 17894
rect 20230 17836 20312 17860
rect 21248 17894 21330 17920
rect 21248 17860 21272 17894
rect 21306 17860 21330 17894
rect 21248 17836 21330 17860
rect 22266 17894 22348 17920
rect 22266 17860 22290 17894
rect 22324 17860 22348 17894
rect 22266 17836 22348 17860
rect 23284 17894 23366 17920
rect 23284 17860 23308 17894
rect 23342 17860 23366 17894
rect 23284 17836 23366 17860
rect 24302 17894 24384 17920
rect 24302 17860 24326 17894
rect 24360 17860 24384 17894
rect 24302 17836 24384 17860
rect 25320 17894 25402 17920
rect 25320 17860 25344 17894
rect 25378 17860 25402 17894
rect 25320 17836 25402 17860
rect 26338 17894 26420 17920
rect 26338 17860 26362 17894
rect 26396 17860 26420 17894
rect 26338 17836 26420 17860
rect 27356 17894 27438 17920
rect 27356 17860 27380 17894
rect 27414 17860 27438 17894
rect 27356 17836 27438 17860
rect 28374 17894 28456 17920
rect 28374 17860 28398 17894
rect 28432 17860 28456 17894
rect 28374 17836 28456 17860
rect 29392 17894 29474 17920
rect 29392 17860 29416 17894
rect 29450 17860 29474 17894
rect 29392 17836 29474 17860
rect 30410 17894 30492 17920
rect 30410 17860 30434 17894
rect 30468 17860 30492 17894
rect 30410 17836 30492 17860
rect 31428 17894 31510 17920
rect 31428 17860 31452 17894
rect 31486 17860 31510 17894
rect 31428 17836 31510 17860
rect 32446 17894 32528 17920
rect 32446 17860 32470 17894
rect 32504 17860 32528 17894
rect 32446 17836 32528 17860
rect 33464 17894 33546 17920
rect 33464 17860 33488 17894
rect 33522 17860 33546 17894
rect 33464 17836 33546 17860
rect 13618 17182 13700 17208
rect 13618 17148 13642 17182
rect 13676 17148 13700 17182
rect 13618 17124 13700 17148
rect 14636 17182 14718 17208
rect 14636 17148 14660 17182
rect 14694 17148 14718 17182
rect 14636 17124 14718 17148
rect 15654 17182 15736 17208
rect 15654 17148 15678 17182
rect 15712 17148 15736 17182
rect 15654 17124 15736 17148
rect 16672 17182 16754 17208
rect 16672 17148 16696 17182
rect 16730 17148 16754 17182
rect 16672 17124 16754 17148
rect 11328 16122 11428 16184
rect 35672 16122 35772 16184
rect 11328 16022 11490 16122
rect 35610 16022 35772 16122
rect 52328 30592 52490 30692
rect 76610 30592 76772 30692
rect 52328 30530 52428 30592
rect 76672 30530 76772 30592
rect 58922 28148 59004 28174
rect 58922 28114 58946 28148
rect 58980 28114 59004 28148
rect 58922 28090 59004 28114
rect 59940 28148 60022 28174
rect 59940 28114 59964 28148
rect 59998 28114 60022 28148
rect 59940 28090 60022 28114
rect 60958 28148 61040 28174
rect 60958 28114 60982 28148
rect 61016 28114 61040 28148
rect 60958 28090 61040 28114
rect 61976 28148 62058 28174
rect 61976 28114 62000 28148
rect 62034 28114 62058 28148
rect 61976 28090 62058 28114
rect 62994 28148 63076 28174
rect 62994 28114 63018 28148
rect 63052 28114 63076 28148
rect 62994 28090 63076 28114
rect 64012 28148 64094 28174
rect 64012 28114 64036 28148
rect 64070 28114 64094 28148
rect 64012 28090 64094 28114
rect 65030 28148 65112 28174
rect 65030 28114 65054 28148
rect 65088 28114 65112 28148
rect 65030 28090 65112 28114
rect 66048 28148 66130 28174
rect 66048 28114 66072 28148
rect 66106 28114 66130 28148
rect 66048 28090 66130 28114
rect 67066 28148 67148 28174
rect 67066 28114 67090 28148
rect 67124 28114 67148 28148
rect 67066 28090 67148 28114
rect 68084 28148 68166 28174
rect 68084 28114 68108 28148
rect 68142 28114 68166 28148
rect 68084 28090 68166 28114
rect 69102 28148 69184 28174
rect 69102 28114 69126 28148
rect 69160 28114 69184 28148
rect 69102 28090 69184 28114
rect 70120 28148 70202 28174
rect 70120 28114 70144 28148
rect 70178 28114 70202 28148
rect 70120 28090 70202 28114
rect 71138 28148 71220 28174
rect 71138 28114 71162 28148
rect 71196 28114 71220 28148
rect 71138 28090 71220 28114
rect 72156 28148 72238 28174
rect 72156 28114 72180 28148
rect 72214 28114 72238 28148
rect 72156 28090 72238 28114
rect 73174 28148 73256 28174
rect 73174 28114 73198 28148
rect 73232 28114 73256 28148
rect 73174 28090 73256 28114
rect 74192 28148 74274 28174
rect 74192 28114 74216 28148
rect 74250 28114 74274 28148
rect 74192 28090 74274 28114
rect 58944 26994 59026 27020
rect 58944 26960 58968 26994
rect 59002 26960 59026 26994
rect 58944 26936 59026 26960
rect 59962 26994 60044 27020
rect 59962 26960 59986 26994
rect 60020 26960 60044 26994
rect 59962 26936 60044 26960
rect 60980 26994 61062 27020
rect 60980 26960 61004 26994
rect 61038 26960 61062 26994
rect 60980 26936 61062 26960
rect 61998 26994 62080 27020
rect 61998 26960 62022 26994
rect 62056 26960 62080 26994
rect 61998 26936 62080 26960
rect 63016 26994 63098 27020
rect 63016 26960 63040 26994
rect 63074 26960 63098 26994
rect 63016 26936 63098 26960
rect 64034 26994 64116 27020
rect 64034 26960 64058 26994
rect 64092 26960 64116 26994
rect 64034 26936 64116 26960
rect 65052 26994 65134 27020
rect 65052 26960 65076 26994
rect 65110 26960 65134 26994
rect 65052 26936 65134 26960
rect 66070 26994 66152 27020
rect 66070 26960 66094 26994
rect 66128 26960 66152 26994
rect 66070 26936 66152 26960
rect 67088 26994 67170 27020
rect 67088 26960 67112 26994
rect 67146 26960 67170 26994
rect 67088 26936 67170 26960
rect 68106 26994 68188 27020
rect 68106 26960 68130 26994
rect 68164 26960 68188 26994
rect 68106 26936 68188 26960
rect 69124 26994 69206 27020
rect 69124 26960 69148 26994
rect 69182 26960 69206 26994
rect 69124 26936 69206 26960
rect 70142 26994 70224 27020
rect 70142 26960 70166 26994
rect 70200 26960 70224 26994
rect 70142 26936 70224 26960
rect 71160 26994 71242 27020
rect 71160 26960 71184 26994
rect 71218 26960 71242 26994
rect 71160 26936 71242 26960
rect 72178 26994 72260 27020
rect 72178 26960 72202 26994
rect 72236 26960 72260 26994
rect 72178 26936 72260 26960
rect 73196 26994 73278 27020
rect 73196 26960 73220 26994
rect 73254 26960 73278 26994
rect 73196 26936 73278 26960
rect 74214 26994 74296 27020
rect 74214 26960 74238 26994
rect 74272 26960 74296 26994
rect 74214 26936 74296 26960
rect 58922 25862 59004 25888
rect 58922 25828 58946 25862
rect 58980 25828 59004 25862
rect 58922 25804 59004 25828
rect 59940 25862 60022 25888
rect 59940 25828 59964 25862
rect 59998 25828 60022 25862
rect 59940 25804 60022 25828
rect 60958 25862 61040 25888
rect 60958 25828 60982 25862
rect 61016 25828 61040 25862
rect 60958 25804 61040 25828
rect 61976 25862 62058 25888
rect 61976 25828 62000 25862
rect 62034 25828 62058 25862
rect 61976 25804 62058 25828
rect 62994 25862 63076 25888
rect 62994 25828 63018 25862
rect 63052 25828 63076 25862
rect 62994 25804 63076 25828
rect 64012 25862 64094 25888
rect 64012 25828 64036 25862
rect 64070 25828 64094 25862
rect 64012 25804 64094 25828
rect 65030 25862 65112 25888
rect 65030 25828 65054 25862
rect 65088 25828 65112 25862
rect 65030 25804 65112 25828
rect 66048 25862 66130 25888
rect 66048 25828 66072 25862
rect 66106 25828 66130 25862
rect 66048 25804 66130 25828
rect 67066 25862 67148 25888
rect 67066 25828 67090 25862
rect 67124 25828 67148 25862
rect 67066 25804 67148 25828
rect 68084 25862 68166 25888
rect 68084 25828 68108 25862
rect 68142 25828 68166 25862
rect 68084 25804 68166 25828
rect 69102 25862 69184 25888
rect 69102 25828 69126 25862
rect 69160 25828 69184 25862
rect 69102 25804 69184 25828
rect 70120 25862 70202 25888
rect 70120 25828 70144 25862
rect 70178 25828 70202 25862
rect 70120 25804 70202 25828
rect 71138 25862 71220 25888
rect 71138 25828 71162 25862
rect 71196 25828 71220 25862
rect 71138 25804 71220 25828
rect 72156 25862 72238 25888
rect 72156 25828 72180 25862
rect 72214 25828 72238 25862
rect 72156 25804 72238 25828
rect 73174 25862 73256 25888
rect 73174 25828 73198 25862
rect 73232 25828 73256 25862
rect 73174 25804 73256 25828
rect 74192 25862 74274 25888
rect 74192 25828 74216 25862
rect 74250 25828 74274 25862
rect 74192 25804 74274 25828
rect 58922 24480 59004 24506
rect 58922 24446 58946 24480
rect 58980 24446 59004 24480
rect 58922 24422 59004 24446
rect 59940 24480 60022 24506
rect 59940 24446 59964 24480
rect 59998 24446 60022 24480
rect 59940 24422 60022 24446
rect 60958 24480 61040 24506
rect 60958 24446 60982 24480
rect 61016 24446 61040 24480
rect 60958 24422 61040 24446
rect 61976 24480 62058 24506
rect 61976 24446 62000 24480
rect 62034 24446 62058 24480
rect 61976 24422 62058 24446
rect 62994 24480 63076 24506
rect 62994 24446 63018 24480
rect 63052 24446 63076 24480
rect 62994 24422 63076 24446
rect 64012 24480 64094 24506
rect 64012 24446 64036 24480
rect 64070 24446 64094 24480
rect 64012 24422 64094 24446
rect 65030 24480 65112 24506
rect 65030 24446 65054 24480
rect 65088 24446 65112 24480
rect 65030 24422 65112 24446
rect 66048 24480 66130 24506
rect 66048 24446 66072 24480
rect 66106 24446 66130 24480
rect 66048 24422 66130 24446
rect 67066 24480 67148 24506
rect 67066 24446 67090 24480
rect 67124 24446 67148 24480
rect 67066 24422 67148 24446
rect 68084 24480 68166 24506
rect 68084 24446 68108 24480
rect 68142 24446 68166 24480
rect 68084 24422 68166 24446
rect 69102 24480 69184 24506
rect 69102 24446 69126 24480
rect 69160 24446 69184 24480
rect 69102 24422 69184 24446
rect 70120 24480 70202 24506
rect 70120 24446 70144 24480
rect 70178 24446 70202 24480
rect 70120 24422 70202 24446
rect 71138 24480 71220 24506
rect 71138 24446 71162 24480
rect 71196 24446 71220 24480
rect 71138 24422 71220 24446
rect 72156 24480 72238 24506
rect 72156 24446 72180 24480
rect 72214 24446 72238 24480
rect 72156 24422 72238 24446
rect 73174 24480 73256 24506
rect 73174 24446 73198 24480
rect 73232 24446 73256 24480
rect 73174 24422 73256 24446
rect 74192 24480 74274 24506
rect 74192 24446 74216 24480
rect 74250 24446 74274 24480
rect 74192 24422 74274 24446
rect 59610 23132 59692 23158
rect 59610 23098 59634 23132
rect 59668 23098 59692 23132
rect 59610 23074 59692 23098
rect 60628 23132 60710 23158
rect 60628 23098 60652 23132
rect 60686 23098 60710 23132
rect 60628 23074 60710 23098
rect 61646 23132 61728 23158
rect 61646 23098 61670 23132
rect 61704 23098 61728 23132
rect 61646 23074 61728 23098
rect 62664 23132 62746 23158
rect 62664 23098 62688 23132
rect 62722 23098 62746 23132
rect 62664 23074 62746 23098
rect 63682 23132 63764 23158
rect 63682 23098 63706 23132
rect 63740 23098 63764 23132
rect 63682 23074 63764 23098
rect 64700 23132 64782 23158
rect 64700 23098 64724 23132
rect 64758 23098 64782 23132
rect 64700 23074 64782 23098
rect 65718 23132 65800 23158
rect 65718 23098 65742 23132
rect 65776 23098 65800 23132
rect 65718 23074 65800 23098
rect 66736 23132 66818 23158
rect 66736 23098 66760 23132
rect 66794 23098 66818 23132
rect 66736 23074 66818 23098
rect 67754 23132 67836 23158
rect 67754 23098 67778 23132
rect 67812 23098 67836 23132
rect 67754 23074 67836 23098
rect 68772 23132 68854 23158
rect 68772 23098 68796 23132
rect 68830 23098 68854 23132
rect 68772 23074 68854 23098
rect 69790 23132 69872 23158
rect 69790 23098 69814 23132
rect 69848 23098 69872 23132
rect 69790 23074 69872 23098
rect 70808 23132 70890 23158
rect 70808 23098 70832 23132
rect 70866 23098 70890 23132
rect 70808 23074 70890 23098
rect 71826 23132 71908 23158
rect 71826 23098 71850 23132
rect 71884 23098 71908 23132
rect 71826 23074 71908 23098
rect 72844 23132 72926 23158
rect 72844 23098 72868 23132
rect 72902 23098 72926 23132
rect 72844 23074 72926 23098
rect 73862 23132 73944 23158
rect 73862 23098 73886 23132
rect 73920 23098 73944 23132
rect 73862 23074 73944 23098
rect 59216 21854 59298 21880
rect 59216 21820 59240 21854
rect 59274 21820 59298 21854
rect 59216 21796 59298 21820
rect 60234 21854 60316 21880
rect 60234 21820 60258 21854
rect 60292 21820 60316 21854
rect 60234 21796 60316 21820
rect 61252 21854 61334 21880
rect 61252 21820 61276 21854
rect 61310 21820 61334 21854
rect 61252 21796 61334 21820
rect 62270 21854 62352 21880
rect 62270 21820 62294 21854
rect 62328 21820 62352 21854
rect 62270 21796 62352 21820
rect 63288 21854 63370 21880
rect 63288 21820 63312 21854
rect 63346 21820 63370 21854
rect 63288 21796 63370 21820
rect 64306 21854 64388 21880
rect 64306 21820 64330 21854
rect 64364 21820 64388 21854
rect 64306 21796 64388 21820
rect 65324 21854 65406 21880
rect 65324 21820 65348 21854
rect 65382 21820 65406 21854
rect 65324 21796 65406 21820
rect 66342 21854 66424 21880
rect 66342 21820 66366 21854
rect 66400 21820 66424 21854
rect 66342 21796 66424 21820
rect 67360 21854 67442 21880
rect 67360 21820 67384 21854
rect 67418 21820 67442 21854
rect 67360 21796 67442 21820
rect 68378 21854 68460 21880
rect 68378 21820 68402 21854
rect 68436 21820 68460 21854
rect 68378 21796 68460 21820
rect 69396 21854 69478 21880
rect 69396 21820 69420 21854
rect 69454 21820 69478 21854
rect 69396 21796 69478 21820
rect 70414 21854 70496 21880
rect 70414 21820 70438 21854
rect 70472 21820 70496 21854
rect 70414 21796 70496 21820
rect 71432 21854 71514 21880
rect 71432 21820 71456 21854
rect 71490 21820 71514 21854
rect 71432 21796 71514 21820
rect 72450 21854 72532 21880
rect 72450 21820 72474 21854
rect 72508 21820 72532 21854
rect 72450 21796 72532 21820
rect 73468 21854 73550 21880
rect 73468 21820 73492 21854
rect 73526 21820 73550 21854
rect 73468 21796 73550 21820
rect 74486 21854 74568 21880
rect 74486 21820 74510 21854
rect 74544 21820 74568 21854
rect 74486 21796 74568 21820
rect 54618 21544 54700 21570
rect 54618 21510 54642 21544
rect 54676 21510 54700 21544
rect 54618 21486 54700 21510
rect 55636 21544 55718 21570
rect 55636 21510 55660 21544
rect 55694 21510 55718 21544
rect 55636 21486 55718 21510
rect 56654 21544 56736 21570
rect 56654 21510 56678 21544
rect 56712 21510 56736 21544
rect 56654 21486 56736 21510
rect 57672 21544 57754 21570
rect 57672 21510 57696 21544
rect 57730 21510 57754 21544
rect 57672 21486 57754 21510
rect 54094 20390 54176 20416
rect 54094 20356 54118 20390
rect 54152 20356 54176 20390
rect 54094 20332 54176 20356
rect 55112 20390 55194 20416
rect 55112 20356 55136 20390
rect 55170 20356 55194 20390
rect 55112 20332 55194 20356
rect 56130 20390 56212 20416
rect 56130 20356 56154 20390
rect 56188 20356 56212 20390
rect 56130 20332 56212 20356
rect 57148 20390 57230 20416
rect 57148 20356 57172 20390
rect 57206 20356 57230 20390
rect 57148 20332 57230 20356
rect 59306 20406 59388 20432
rect 59306 20372 59330 20406
rect 59364 20372 59388 20406
rect 59306 20348 59388 20372
rect 60324 20406 60406 20432
rect 60324 20372 60348 20406
rect 60382 20372 60406 20406
rect 60324 20348 60406 20372
rect 61342 20406 61424 20432
rect 61342 20372 61366 20406
rect 61400 20372 61424 20406
rect 61342 20348 61424 20372
rect 62360 20406 62442 20432
rect 62360 20372 62384 20406
rect 62418 20372 62442 20406
rect 62360 20348 62442 20372
rect 63378 20406 63460 20432
rect 63378 20372 63402 20406
rect 63436 20372 63460 20406
rect 63378 20348 63460 20372
rect 64396 20406 64478 20432
rect 64396 20372 64420 20406
rect 64454 20372 64478 20406
rect 64396 20348 64478 20372
rect 65414 20406 65496 20432
rect 65414 20372 65438 20406
rect 65472 20372 65496 20406
rect 65414 20348 65496 20372
rect 66432 20406 66514 20432
rect 66432 20372 66456 20406
rect 66490 20372 66514 20406
rect 66432 20348 66514 20372
rect 67450 20406 67532 20432
rect 67450 20372 67474 20406
rect 67508 20372 67532 20406
rect 67450 20348 67532 20372
rect 68468 20406 68550 20432
rect 68468 20372 68492 20406
rect 68526 20372 68550 20406
rect 68468 20348 68550 20372
rect 69486 20406 69568 20432
rect 69486 20372 69510 20406
rect 69544 20372 69568 20406
rect 69486 20348 69568 20372
rect 70504 20406 70586 20432
rect 70504 20372 70528 20406
rect 70562 20372 70586 20406
rect 70504 20348 70586 20372
rect 71522 20406 71604 20432
rect 71522 20372 71546 20406
rect 71580 20372 71604 20406
rect 71522 20348 71604 20372
rect 72540 20406 72622 20432
rect 72540 20372 72564 20406
rect 72598 20372 72622 20406
rect 72540 20348 72622 20372
rect 73558 20406 73640 20432
rect 73558 20372 73582 20406
rect 73616 20372 73640 20406
rect 73558 20348 73640 20372
rect 74576 20406 74658 20432
rect 74576 20372 74600 20406
rect 74634 20372 74658 20406
rect 74576 20348 74658 20372
rect 54104 19362 54186 19388
rect 54104 19328 54128 19362
rect 54162 19328 54186 19362
rect 54104 19304 54186 19328
rect 55122 19362 55204 19388
rect 55122 19328 55146 19362
rect 55180 19328 55204 19362
rect 55122 19304 55204 19328
rect 56140 19362 56222 19388
rect 56140 19328 56164 19362
rect 56198 19328 56222 19362
rect 56140 19304 56222 19328
rect 57158 19362 57240 19388
rect 57158 19328 57182 19362
rect 57216 19328 57240 19362
rect 57158 19304 57240 19328
rect 59330 19138 59412 19164
rect 59330 19104 59354 19138
rect 59388 19104 59412 19138
rect 59330 19080 59412 19104
rect 60348 19138 60430 19164
rect 60348 19104 60372 19138
rect 60406 19104 60430 19138
rect 60348 19080 60430 19104
rect 61366 19138 61448 19164
rect 61366 19104 61390 19138
rect 61424 19104 61448 19138
rect 61366 19080 61448 19104
rect 62384 19138 62466 19164
rect 62384 19104 62408 19138
rect 62442 19104 62466 19138
rect 62384 19080 62466 19104
rect 63402 19138 63484 19164
rect 63402 19104 63426 19138
rect 63460 19104 63484 19138
rect 63402 19080 63484 19104
rect 64420 19138 64502 19164
rect 64420 19104 64444 19138
rect 64478 19104 64502 19138
rect 64420 19080 64502 19104
rect 65438 19138 65520 19164
rect 65438 19104 65462 19138
rect 65496 19104 65520 19138
rect 65438 19080 65520 19104
rect 66456 19138 66538 19164
rect 66456 19104 66480 19138
rect 66514 19104 66538 19138
rect 66456 19080 66538 19104
rect 67474 19138 67556 19164
rect 67474 19104 67498 19138
rect 67532 19104 67556 19138
rect 67474 19080 67556 19104
rect 68492 19138 68574 19164
rect 68492 19104 68516 19138
rect 68550 19104 68574 19138
rect 68492 19080 68574 19104
rect 69510 19138 69592 19164
rect 69510 19104 69534 19138
rect 69568 19104 69592 19138
rect 69510 19080 69592 19104
rect 70528 19138 70610 19164
rect 70528 19104 70552 19138
rect 70586 19104 70610 19138
rect 70528 19080 70610 19104
rect 71546 19138 71628 19164
rect 71546 19104 71570 19138
rect 71604 19104 71628 19138
rect 71546 19080 71628 19104
rect 72564 19138 72646 19164
rect 72564 19104 72588 19138
rect 72622 19104 72646 19138
rect 72564 19080 72646 19104
rect 73582 19138 73664 19164
rect 73582 19104 73606 19138
rect 73640 19104 73664 19138
rect 73582 19080 73664 19104
rect 74600 19138 74682 19164
rect 74600 19104 74624 19138
rect 74658 19104 74682 19138
rect 74600 19080 74682 19104
rect 54094 18334 54176 18360
rect 54094 18300 54118 18334
rect 54152 18300 54176 18334
rect 54094 18276 54176 18300
rect 55112 18334 55194 18360
rect 55112 18300 55136 18334
rect 55170 18300 55194 18334
rect 55112 18276 55194 18300
rect 56130 18334 56212 18360
rect 56130 18300 56154 18334
rect 56188 18300 56212 18334
rect 56130 18276 56212 18300
rect 57148 18334 57230 18360
rect 57148 18300 57172 18334
rect 57206 18300 57230 18334
rect 57148 18276 57230 18300
rect 59194 17894 59276 17920
rect 59194 17860 59218 17894
rect 59252 17860 59276 17894
rect 59194 17836 59276 17860
rect 60212 17894 60294 17920
rect 60212 17860 60236 17894
rect 60270 17860 60294 17894
rect 60212 17836 60294 17860
rect 61230 17894 61312 17920
rect 61230 17860 61254 17894
rect 61288 17860 61312 17894
rect 61230 17836 61312 17860
rect 62248 17894 62330 17920
rect 62248 17860 62272 17894
rect 62306 17860 62330 17894
rect 62248 17836 62330 17860
rect 63266 17894 63348 17920
rect 63266 17860 63290 17894
rect 63324 17860 63348 17894
rect 63266 17836 63348 17860
rect 64284 17894 64366 17920
rect 64284 17860 64308 17894
rect 64342 17860 64366 17894
rect 64284 17836 64366 17860
rect 65302 17894 65384 17920
rect 65302 17860 65326 17894
rect 65360 17860 65384 17894
rect 65302 17836 65384 17860
rect 66320 17894 66402 17920
rect 66320 17860 66344 17894
rect 66378 17860 66402 17894
rect 66320 17836 66402 17860
rect 67338 17894 67420 17920
rect 67338 17860 67362 17894
rect 67396 17860 67420 17894
rect 67338 17836 67420 17860
rect 68356 17894 68438 17920
rect 68356 17860 68380 17894
rect 68414 17860 68438 17894
rect 68356 17836 68438 17860
rect 69374 17894 69456 17920
rect 69374 17860 69398 17894
rect 69432 17860 69456 17894
rect 69374 17836 69456 17860
rect 70392 17894 70474 17920
rect 70392 17860 70416 17894
rect 70450 17860 70474 17894
rect 70392 17836 70474 17860
rect 71410 17894 71492 17920
rect 71410 17860 71434 17894
rect 71468 17860 71492 17894
rect 71410 17836 71492 17860
rect 72428 17894 72510 17920
rect 72428 17860 72452 17894
rect 72486 17860 72510 17894
rect 72428 17836 72510 17860
rect 73446 17894 73528 17920
rect 73446 17860 73470 17894
rect 73504 17860 73528 17894
rect 73446 17836 73528 17860
rect 74464 17894 74546 17920
rect 74464 17860 74488 17894
rect 74522 17860 74546 17894
rect 74464 17836 74546 17860
rect 54618 17182 54700 17208
rect 54618 17148 54642 17182
rect 54676 17148 54700 17182
rect 54618 17124 54700 17148
rect 55636 17182 55718 17208
rect 55636 17148 55660 17182
rect 55694 17148 55718 17182
rect 55636 17124 55718 17148
rect 56654 17182 56736 17208
rect 56654 17148 56678 17182
rect 56712 17148 56736 17182
rect 56654 17124 56736 17148
rect 57672 17182 57754 17208
rect 57672 17148 57696 17182
rect 57730 17148 57754 17182
rect 57672 17124 57754 17148
rect 52328 16122 52428 16184
rect 76672 16122 76772 16184
rect 52328 16022 52490 16122
rect 76610 16022 76772 16122
rect 36718 13870 36880 13970
rect 38520 13870 38682 13970
rect 36718 13808 36818 13870
rect 38582 13808 38682 13870
rect 36718 12526 36818 12588
rect 38582 12526 38682 12588
rect 36718 12426 36880 12526
rect 38520 12426 38682 12526
<< psubdiffcont >>
rect -1210 15092 35710 15192
rect -1372 -690 -1272 15030
rect 14060 14552 14094 14586
rect 15078 14552 15112 14586
rect 16096 14552 16130 14586
rect 17114 14552 17148 14586
rect 18132 14552 18166 14586
rect 19150 14552 19184 14586
rect 20168 14552 20202 14586
rect 21186 14552 21220 14586
rect 22204 14552 22238 14586
rect 23222 14552 23256 14586
rect 24240 14552 24274 14586
rect 25258 14552 25292 14586
rect 26276 14552 26310 14586
rect 27294 14552 27328 14586
rect 28312 14552 28346 14586
rect 29330 14552 29364 14586
rect 30348 14552 30382 14586
rect 31366 14552 31400 14586
rect 32384 14552 32418 14586
rect 33402 14552 33436 14586
rect 1766 13950 1800 13984
rect 2784 13950 2818 13984
rect 3802 13950 3836 13984
rect 4820 13950 4854 13984
rect 5838 13950 5872 13984
rect 6856 13950 6890 13984
rect 7874 13950 7908 13984
rect 8892 13950 8926 13984
rect 9910 13950 9944 13984
rect 10938 13950 10972 13984
rect 1766 13132 1800 13166
rect 2784 13132 2818 13166
rect 3802 13132 3836 13166
rect 4820 13132 4854 13166
rect 5838 13132 5872 13166
rect 6856 13132 6890 13166
rect 7874 13132 7908 13166
rect 8892 13132 8926 13166
rect 9910 13132 9944 13166
rect 10938 13132 10972 13166
rect 14072 12526 14106 12560
rect 15090 12526 15124 12560
rect 16108 12526 16142 12560
rect 17126 12526 17160 12560
rect 18144 12526 18178 12560
rect 19162 12526 19196 12560
rect 20180 12526 20214 12560
rect 21198 12526 21232 12560
rect 22216 12526 22250 12560
rect 23234 12526 23268 12560
rect 24252 12526 24286 12560
rect 25270 12526 25304 12560
rect 26288 12526 26322 12560
rect 27306 12526 27340 12560
rect 28324 12526 28358 12560
rect 29342 12526 29376 12560
rect 30360 12526 30394 12560
rect 31378 12526 31412 12560
rect 32396 12526 32430 12560
rect 33414 12526 33448 12560
rect 1766 12314 1800 12348
rect 2784 12314 2818 12348
rect 3802 12314 3836 12348
rect 4820 12314 4854 12348
rect 5838 12314 5872 12348
rect 6856 12314 6890 12348
rect 7874 12314 7908 12348
rect 8892 12314 8926 12348
rect 9910 12314 9944 12348
rect 10938 12314 10972 12348
rect 1766 11496 1800 11530
rect 2784 11496 2818 11530
rect 3802 11496 3836 11530
rect 4820 11496 4854 11530
rect 5838 11496 5872 11530
rect 6856 11496 6890 11530
rect 7874 11496 7908 11530
rect 8892 11496 8926 11530
rect 9910 11496 9944 11530
rect 10938 11496 10972 11530
rect 14060 11220 14094 11254
rect 15078 11220 15112 11254
rect 16096 11220 16130 11254
rect 17114 11220 17148 11254
rect 18132 11220 18166 11254
rect 19150 11220 19184 11254
rect 20168 11220 20202 11254
rect 21186 11220 21220 11254
rect 22204 11220 22238 11254
rect 23222 11220 23256 11254
rect 24240 11220 24274 11254
rect 25258 11220 25292 11254
rect 26276 11220 26310 11254
rect 27294 11220 27328 11254
rect 28312 11220 28346 11254
rect 29330 11220 29364 11254
rect 30348 11220 30382 11254
rect 31366 11220 31400 11254
rect 32384 11220 32418 11254
rect 33402 11220 33436 11254
rect 1766 10678 1800 10712
rect 2784 10678 2818 10712
rect 3802 10678 3836 10712
rect 4820 10678 4854 10712
rect 5838 10678 5872 10712
rect 6856 10678 6890 10712
rect 7874 10678 7908 10712
rect 8892 10678 8926 10712
rect 9910 10678 9944 10712
rect 10938 10678 10972 10712
rect 1766 9860 1800 9894
rect 2784 9860 2818 9894
rect 3802 9860 3836 9894
rect 4820 9860 4854 9894
rect 5838 9860 5872 9894
rect 6856 9860 6890 9894
rect 7874 9860 7908 9894
rect 14048 9984 14082 10018
rect 15066 9984 15100 10018
rect 16084 9984 16118 10018
rect 17102 9984 17136 10018
rect 18120 9984 18154 10018
rect 19138 9984 19172 10018
rect 20156 9984 20190 10018
rect 21174 9984 21208 10018
rect 22192 9984 22226 10018
rect 23210 9984 23244 10018
rect 24228 9984 24262 10018
rect 25246 9984 25280 10018
rect 26264 9984 26298 10018
rect 27282 9984 27316 10018
rect 28300 9984 28334 10018
rect 29318 9984 29352 10018
rect 30336 9984 30370 10018
rect 31354 9984 31388 10018
rect 32372 9984 32406 10018
rect 33390 9984 33424 10018
rect 8892 9860 8926 9894
rect 9910 9860 9944 9894
rect 10938 9860 10972 9894
rect 1766 9042 1800 9076
rect 2784 9042 2818 9076
rect 3802 9042 3836 9076
rect 4820 9042 4854 9076
rect 5838 9042 5872 9076
rect 6856 9042 6890 9076
rect 7874 9042 7908 9076
rect 8892 9042 8926 9076
rect 9910 9042 9944 9076
rect 10938 9042 10972 9076
rect 14048 8760 14082 8794
rect 15066 8760 15100 8794
rect 16084 8760 16118 8794
rect 17102 8760 17136 8794
rect 18120 8760 18154 8794
rect 19138 8760 19172 8794
rect 20156 8760 20190 8794
rect 21174 8760 21208 8794
rect 22192 8760 22226 8794
rect 23210 8760 23244 8794
rect 24228 8760 24262 8794
rect 25246 8760 25280 8794
rect 26264 8760 26298 8794
rect 27282 8760 27316 8794
rect 28300 8760 28334 8794
rect 29318 8760 29352 8794
rect 30336 8760 30370 8794
rect 31354 8760 31388 8794
rect 32372 8760 32406 8794
rect 33390 8760 33424 8794
rect 1766 8224 1800 8258
rect 2784 8224 2818 8258
rect 3802 8224 3836 8258
rect 4820 8224 4854 8258
rect 5838 8224 5872 8258
rect 6856 8224 6890 8258
rect 7874 8224 7908 8258
rect 8892 8224 8926 8258
rect 9910 8224 9944 8258
rect 10938 8224 10972 8258
rect 14060 7524 14094 7558
rect 15078 7524 15112 7558
rect 16096 7524 16130 7558
rect 17114 7524 17148 7558
rect 18132 7524 18166 7558
rect 19150 7524 19184 7558
rect 20168 7524 20202 7558
rect 21186 7524 21220 7558
rect 22204 7524 22238 7558
rect 23222 7524 23256 7558
rect 24240 7524 24274 7558
rect 25258 7524 25292 7558
rect 26276 7524 26310 7558
rect 27294 7524 27328 7558
rect 28312 7524 28346 7558
rect 29330 7524 29364 7558
rect 30348 7524 30382 7558
rect 31366 7524 31400 7558
rect 32384 7524 32418 7558
rect 33402 7524 33436 7558
rect 1754 7330 1788 7364
rect 2772 7330 2806 7364
rect 3790 7330 3824 7364
rect 4808 7330 4842 7364
rect 5826 7330 5860 7364
rect 6844 7330 6878 7364
rect 7862 7330 7896 7364
rect 8880 7330 8914 7364
rect 9898 7330 9932 7364
rect 10926 7330 10960 7364
rect 958 6382 992 6416
rect 1976 6382 2010 6416
rect 2994 6382 3028 6416
rect 4012 6382 4046 6416
rect 5030 6382 5064 6416
rect 6048 6382 6082 6416
rect 7066 6382 7100 6416
rect 8084 6382 8118 6416
rect 9102 6382 9136 6416
rect 10120 6382 10154 6416
rect 11138 6382 11172 6416
rect 14060 6276 14094 6310
rect 15078 6276 15112 6310
rect 16096 6276 16130 6310
rect 17114 6276 17148 6310
rect 18132 6276 18166 6310
rect 19150 6276 19184 6310
rect 20168 6276 20202 6310
rect 21186 6276 21220 6310
rect 22204 6276 22238 6310
rect 23222 6276 23256 6310
rect 24240 6276 24274 6310
rect 25258 6276 25292 6310
rect 26276 6276 26310 6310
rect 27294 6276 27328 6310
rect 28312 6276 28346 6310
rect 29330 6276 29364 6310
rect 30348 6276 30382 6310
rect 31366 6276 31400 6310
rect 32384 6276 32418 6310
rect 33402 6276 33436 6310
rect 970 5240 1004 5274
rect 1988 5240 2022 5274
rect 3006 5240 3040 5274
rect 4024 5240 4058 5274
rect 5042 5240 5076 5274
rect 6060 5240 6094 5274
rect 7078 5240 7112 5274
rect 8096 5240 8130 5274
rect 9114 5240 9148 5274
rect 10132 5240 10166 5274
rect 11150 5240 11184 5274
rect 14036 5040 14070 5074
rect 15054 5040 15088 5074
rect 16072 5040 16106 5074
rect 17090 5040 17124 5074
rect 18108 5040 18142 5074
rect 19126 5040 19160 5074
rect 20144 5040 20178 5074
rect 21162 5040 21196 5074
rect 22180 5040 22214 5074
rect 23198 5040 23232 5074
rect 24216 5040 24250 5074
rect 25234 5040 25268 5074
rect 26252 5040 26286 5074
rect 27270 5040 27304 5074
rect 28288 5040 28322 5074
rect 29306 5040 29340 5074
rect 30324 5040 30358 5074
rect 31342 5040 31376 5074
rect 32360 5040 32394 5074
rect 33378 5040 33412 5074
rect 948 4132 982 4166
rect 1966 4132 2000 4166
rect 2984 4132 3018 4166
rect 4002 4132 4036 4166
rect 5020 4132 5054 4166
rect 6038 4132 6072 4166
rect 7056 4132 7090 4166
rect 8074 4132 8108 4166
rect 9092 4132 9126 4166
rect 10110 4132 10144 4166
rect 11128 4132 11162 4166
rect 14048 3816 14082 3850
rect 15066 3816 15100 3850
rect 16084 3816 16118 3850
rect 17102 3816 17136 3850
rect 18120 3816 18154 3850
rect 19138 3816 19172 3850
rect 20156 3816 20190 3850
rect 21174 3816 21208 3850
rect 22192 3816 22226 3850
rect 23210 3816 23244 3850
rect 24228 3816 24262 3850
rect 25246 3816 25280 3850
rect 26264 3816 26298 3850
rect 27282 3816 27316 3850
rect 28300 3816 28334 3850
rect 29318 3816 29352 3850
rect 30336 3816 30370 3850
rect 31354 3816 31388 3850
rect 32372 3816 32406 3850
rect 33390 3816 33424 3850
rect 948 3026 982 3060
rect 1966 3026 2000 3060
rect 2984 3026 3018 3060
rect 4002 3026 4036 3060
rect 5020 3026 5054 3060
rect 6038 3026 6072 3060
rect 7056 3026 7090 3060
rect 8074 3026 8108 3060
rect 9092 3026 9126 3060
rect 10110 3026 10144 3060
rect 11128 3026 11162 3060
rect 14048 2580 14082 2614
rect 15066 2580 15100 2614
rect 16084 2580 16118 2614
rect 17102 2580 17136 2614
rect 18120 2580 18154 2614
rect 19138 2580 19172 2614
rect 20156 2580 20190 2614
rect 21174 2580 21208 2614
rect 22192 2580 22226 2614
rect 23210 2580 23244 2614
rect 24228 2580 24262 2614
rect 25246 2580 25280 2614
rect 26264 2580 26298 2614
rect 27282 2580 27316 2614
rect 28300 2580 28334 2614
rect 29318 2580 29352 2614
rect 30336 2580 30370 2614
rect 31354 2580 31388 2614
rect 32372 2580 32406 2614
rect 33390 2580 33424 2614
rect 948 1684 982 1718
rect 1966 1684 2000 1718
rect 2984 1684 3018 1718
rect 4002 1684 4036 1718
rect 5020 1684 5054 1718
rect 6038 1684 6072 1718
rect 7056 1684 7090 1718
rect 8074 1684 8108 1718
rect 9092 1684 9126 1718
rect 10110 1684 10144 1718
rect 11128 1684 11162 1718
rect 14060 1334 14094 1368
rect 15078 1334 15112 1368
rect 16096 1334 16130 1368
rect 17114 1334 17148 1368
rect 18132 1334 18166 1368
rect 19150 1334 19184 1368
rect 20168 1334 20202 1368
rect 21186 1334 21220 1368
rect 22204 1334 22238 1368
rect 23222 1334 23256 1368
rect 24240 1334 24274 1368
rect 25258 1334 25292 1368
rect 26276 1334 26310 1368
rect 27294 1334 27328 1368
rect 28312 1334 28346 1368
rect 29330 1334 29364 1368
rect 30348 1334 30382 1368
rect 31366 1334 31400 1368
rect 32384 1334 32418 1368
rect 33402 1334 33436 1368
rect -1092 362 -934 396
rect -1188 51 -1154 223
rect -872 51 -838 223
rect 758 238 792 272
rect 1776 238 1810 272
rect 2794 238 2828 272
rect 3812 238 3846 272
rect 4830 238 4864 272
rect 5848 238 5882 272
rect 6866 238 6900 272
rect 7884 238 7918 272
rect 8902 238 8936 272
rect 9920 238 9954 272
rect 10938 238 10972 272
rect 14048 156 14082 190
rect 15066 156 15100 190
rect 16084 156 16118 190
rect 17102 156 17136 190
rect 18120 156 18154 190
rect 19138 156 19172 190
rect 20156 156 20190 190
rect 21174 156 21208 190
rect 22192 156 22226 190
rect 23210 156 23244 190
rect 24228 156 24262 190
rect 25246 156 25280 190
rect 26264 156 26298 190
rect 27282 156 27316 190
rect 28300 156 28334 190
rect 29318 156 29352 190
rect 30336 156 30370 190
rect 31354 156 31388 190
rect 32372 156 32406 190
rect 33390 156 33424 190
rect -1092 -136 -934 -102
rect 35772 -690 35872 15030
rect 39790 15092 76710 15192
rect -1210 -852 35710 -752
rect 39628 -690 39728 15030
rect 55060 14552 55094 14586
rect 56078 14552 56112 14586
rect 57096 14552 57130 14586
rect 58114 14552 58148 14586
rect 59132 14552 59166 14586
rect 60150 14552 60184 14586
rect 61168 14552 61202 14586
rect 62186 14552 62220 14586
rect 63204 14552 63238 14586
rect 64222 14552 64256 14586
rect 65240 14552 65274 14586
rect 66258 14552 66292 14586
rect 67276 14552 67310 14586
rect 68294 14552 68328 14586
rect 69312 14552 69346 14586
rect 70330 14552 70364 14586
rect 71348 14552 71382 14586
rect 72366 14552 72400 14586
rect 73384 14552 73418 14586
rect 74402 14552 74436 14586
rect 42766 13950 42800 13984
rect 43784 13950 43818 13984
rect 44802 13950 44836 13984
rect 45820 13950 45854 13984
rect 46838 13950 46872 13984
rect 47856 13950 47890 13984
rect 48874 13950 48908 13984
rect 49892 13950 49926 13984
rect 50910 13950 50944 13984
rect 51938 13950 51972 13984
rect 42766 13132 42800 13166
rect 43784 13132 43818 13166
rect 44802 13132 44836 13166
rect 45820 13132 45854 13166
rect 46838 13132 46872 13166
rect 47856 13132 47890 13166
rect 48874 13132 48908 13166
rect 49892 13132 49926 13166
rect 50910 13132 50944 13166
rect 51938 13132 51972 13166
rect 55072 12526 55106 12560
rect 56090 12526 56124 12560
rect 57108 12526 57142 12560
rect 58126 12526 58160 12560
rect 59144 12526 59178 12560
rect 60162 12526 60196 12560
rect 61180 12526 61214 12560
rect 62198 12526 62232 12560
rect 63216 12526 63250 12560
rect 64234 12526 64268 12560
rect 65252 12526 65286 12560
rect 66270 12526 66304 12560
rect 67288 12526 67322 12560
rect 68306 12526 68340 12560
rect 69324 12526 69358 12560
rect 70342 12526 70376 12560
rect 71360 12526 71394 12560
rect 72378 12526 72412 12560
rect 73396 12526 73430 12560
rect 74414 12526 74448 12560
rect 42766 12314 42800 12348
rect 43784 12314 43818 12348
rect 44802 12314 44836 12348
rect 45820 12314 45854 12348
rect 46838 12314 46872 12348
rect 47856 12314 47890 12348
rect 48874 12314 48908 12348
rect 49892 12314 49926 12348
rect 50910 12314 50944 12348
rect 51938 12314 51972 12348
rect 42766 11496 42800 11530
rect 43784 11496 43818 11530
rect 44802 11496 44836 11530
rect 45820 11496 45854 11530
rect 46838 11496 46872 11530
rect 47856 11496 47890 11530
rect 48874 11496 48908 11530
rect 49892 11496 49926 11530
rect 50910 11496 50944 11530
rect 51938 11496 51972 11530
rect 55060 11220 55094 11254
rect 56078 11220 56112 11254
rect 57096 11220 57130 11254
rect 58114 11220 58148 11254
rect 59132 11220 59166 11254
rect 60150 11220 60184 11254
rect 61168 11220 61202 11254
rect 62186 11220 62220 11254
rect 63204 11220 63238 11254
rect 64222 11220 64256 11254
rect 65240 11220 65274 11254
rect 66258 11220 66292 11254
rect 67276 11220 67310 11254
rect 68294 11220 68328 11254
rect 69312 11220 69346 11254
rect 70330 11220 70364 11254
rect 71348 11220 71382 11254
rect 72366 11220 72400 11254
rect 73384 11220 73418 11254
rect 74402 11220 74436 11254
rect 42766 10678 42800 10712
rect 43784 10678 43818 10712
rect 44802 10678 44836 10712
rect 45820 10678 45854 10712
rect 46838 10678 46872 10712
rect 47856 10678 47890 10712
rect 48874 10678 48908 10712
rect 49892 10678 49926 10712
rect 50910 10678 50944 10712
rect 51938 10678 51972 10712
rect 42766 9860 42800 9894
rect 43784 9860 43818 9894
rect 44802 9860 44836 9894
rect 45820 9860 45854 9894
rect 46838 9860 46872 9894
rect 47856 9860 47890 9894
rect 48874 9860 48908 9894
rect 55048 9984 55082 10018
rect 56066 9984 56100 10018
rect 57084 9984 57118 10018
rect 58102 9984 58136 10018
rect 59120 9984 59154 10018
rect 60138 9984 60172 10018
rect 61156 9984 61190 10018
rect 62174 9984 62208 10018
rect 63192 9984 63226 10018
rect 64210 9984 64244 10018
rect 65228 9984 65262 10018
rect 66246 9984 66280 10018
rect 67264 9984 67298 10018
rect 68282 9984 68316 10018
rect 69300 9984 69334 10018
rect 70318 9984 70352 10018
rect 71336 9984 71370 10018
rect 72354 9984 72388 10018
rect 73372 9984 73406 10018
rect 74390 9984 74424 10018
rect 49892 9860 49926 9894
rect 50910 9860 50944 9894
rect 51938 9860 51972 9894
rect 42766 9042 42800 9076
rect 43784 9042 43818 9076
rect 44802 9042 44836 9076
rect 45820 9042 45854 9076
rect 46838 9042 46872 9076
rect 47856 9042 47890 9076
rect 48874 9042 48908 9076
rect 49892 9042 49926 9076
rect 50910 9042 50944 9076
rect 51938 9042 51972 9076
rect 55048 8760 55082 8794
rect 56066 8760 56100 8794
rect 57084 8760 57118 8794
rect 58102 8760 58136 8794
rect 59120 8760 59154 8794
rect 60138 8760 60172 8794
rect 61156 8760 61190 8794
rect 62174 8760 62208 8794
rect 63192 8760 63226 8794
rect 64210 8760 64244 8794
rect 65228 8760 65262 8794
rect 66246 8760 66280 8794
rect 67264 8760 67298 8794
rect 68282 8760 68316 8794
rect 69300 8760 69334 8794
rect 70318 8760 70352 8794
rect 71336 8760 71370 8794
rect 72354 8760 72388 8794
rect 73372 8760 73406 8794
rect 74390 8760 74424 8794
rect 42766 8224 42800 8258
rect 43784 8224 43818 8258
rect 44802 8224 44836 8258
rect 45820 8224 45854 8258
rect 46838 8224 46872 8258
rect 47856 8224 47890 8258
rect 48874 8224 48908 8258
rect 49892 8224 49926 8258
rect 50910 8224 50944 8258
rect 51938 8224 51972 8258
rect 55060 7524 55094 7558
rect 56078 7524 56112 7558
rect 57096 7524 57130 7558
rect 58114 7524 58148 7558
rect 59132 7524 59166 7558
rect 60150 7524 60184 7558
rect 61168 7524 61202 7558
rect 62186 7524 62220 7558
rect 63204 7524 63238 7558
rect 64222 7524 64256 7558
rect 65240 7524 65274 7558
rect 66258 7524 66292 7558
rect 67276 7524 67310 7558
rect 68294 7524 68328 7558
rect 69312 7524 69346 7558
rect 70330 7524 70364 7558
rect 71348 7524 71382 7558
rect 72366 7524 72400 7558
rect 73384 7524 73418 7558
rect 74402 7524 74436 7558
rect 42754 7330 42788 7364
rect 43772 7330 43806 7364
rect 44790 7330 44824 7364
rect 45808 7330 45842 7364
rect 46826 7330 46860 7364
rect 47844 7330 47878 7364
rect 48862 7330 48896 7364
rect 49880 7330 49914 7364
rect 50898 7330 50932 7364
rect 51926 7330 51960 7364
rect 41958 6382 41992 6416
rect 42976 6382 43010 6416
rect 43994 6382 44028 6416
rect 45012 6382 45046 6416
rect 46030 6382 46064 6416
rect 47048 6382 47082 6416
rect 48066 6382 48100 6416
rect 49084 6382 49118 6416
rect 50102 6382 50136 6416
rect 51120 6382 51154 6416
rect 52138 6382 52172 6416
rect 55060 6276 55094 6310
rect 56078 6276 56112 6310
rect 57096 6276 57130 6310
rect 58114 6276 58148 6310
rect 59132 6276 59166 6310
rect 60150 6276 60184 6310
rect 61168 6276 61202 6310
rect 62186 6276 62220 6310
rect 63204 6276 63238 6310
rect 64222 6276 64256 6310
rect 65240 6276 65274 6310
rect 66258 6276 66292 6310
rect 67276 6276 67310 6310
rect 68294 6276 68328 6310
rect 69312 6276 69346 6310
rect 70330 6276 70364 6310
rect 71348 6276 71382 6310
rect 72366 6276 72400 6310
rect 73384 6276 73418 6310
rect 74402 6276 74436 6310
rect 41970 5240 42004 5274
rect 42988 5240 43022 5274
rect 44006 5240 44040 5274
rect 45024 5240 45058 5274
rect 46042 5240 46076 5274
rect 47060 5240 47094 5274
rect 48078 5240 48112 5274
rect 49096 5240 49130 5274
rect 50114 5240 50148 5274
rect 51132 5240 51166 5274
rect 52150 5240 52184 5274
rect 55036 5040 55070 5074
rect 56054 5040 56088 5074
rect 57072 5040 57106 5074
rect 58090 5040 58124 5074
rect 59108 5040 59142 5074
rect 60126 5040 60160 5074
rect 61144 5040 61178 5074
rect 62162 5040 62196 5074
rect 63180 5040 63214 5074
rect 64198 5040 64232 5074
rect 65216 5040 65250 5074
rect 66234 5040 66268 5074
rect 67252 5040 67286 5074
rect 68270 5040 68304 5074
rect 69288 5040 69322 5074
rect 70306 5040 70340 5074
rect 71324 5040 71358 5074
rect 72342 5040 72376 5074
rect 73360 5040 73394 5074
rect 74378 5040 74412 5074
rect 41948 4132 41982 4166
rect 42966 4132 43000 4166
rect 43984 4132 44018 4166
rect 45002 4132 45036 4166
rect 46020 4132 46054 4166
rect 47038 4132 47072 4166
rect 48056 4132 48090 4166
rect 49074 4132 49108 4166
rect 50092 4132 50126 4166
rect 51110 4132 51144 4166
rect 52128 4132 52162 4166
rect 55048 3816 55082 3850
rect 56066 3816 56100 3850
rect 57084 3816 57118 3850
rect 58102 3816 58136 3850
rect 59120 3816 59154 3850
rect 60138 3816 60172 3850
rect 61156 3816 61190 3850
rect 62174 3816 62208 3850
rect 63192 3816 63226 3850
rect 64210 3816 64244 3850
rect 65228 3816 65262 3850
rect 66246 3816 66280 3850
rect 67264 3816 67298 3850
rect 68282 3816 68316 3850
rect 69300 3816 69334 3850
rect 70318 3816 70352 3850
rect 71336 3816 71370 3850
rect 72354 3816 72388 3850
rect 73372 3816 73406 3850
rect 74390 3816 74424 3850
rect 41948 3026 41982 3060
rect 42966 3026 43000 3060
rect 43984 3026 44018 3060
rect 45002 3026 45036 3060
rect 46020 3026 46054 3060
rect 47038 3026 47072 3060
rect 48056 3026 48090 3060
rect 49074 3026 49108 3060
rect 50092 3026 50126 3060
rect 51110 3026 51144 3060
rect 52128 3026 52162 3060
rect 55048 2580 55082 2614
rect 56066 2580 56100 2614
rect 57084 2580 57118 2614
rect 58102 2580 58136 2614
rect 59120 2580 59154 2614
rect 60138 2580 60172 2614
rect 61156 2580 61190 2614
rect 62174 2580 62208 2614
rect 63192 2580 63226 2614
rect 64210 2580 64244 2614
rect 65228 2580 65262 2614
rect 66246 2580 66280 2614
rect 67264 2580 67298 2614
rect 68282 2580 68316 2614
rect 69300 2580 69334 2614
rect 70318 2580 70352 2614
rect 71336 2580 71370 2614
rect 72354 2580 72388 2614
rect 73372 2580 73406 2614
rect 74390 2580 74424 2614
rect 41948 1684 41982 1718
rect 42966 1684 43000 1718
rect 43984 1684 44018 1718
rect 45002 1684 45036 1718
rect 46020 1684 46054 1718
rect 47038 1684 47072 1718
rect 48056 1684 48090 1718
rect 49074 1684 49108 1718
rect 50092 1684 50126 1718
rect 51110 1684 51144 1718
rect 52128 1684 52162 1718
rect 55060 1334 55094 1368
rect 56078 1334 56112 1368
rect 57096 1334 57130 1368
rect 58114 1334 58148 1368
rect 59132 1334 59166 1368
rect 60150 1334 60184 1368
rect 61168 1334 61202 1368
rect 62186 1334 62220 1368
rect 63204 1334 63238 1368
rect 64222 1334 64256 1368
rect 65240 1334 65274 1368
rect 66258 1334 66292 1368
rect 67276 1334 67310 1368
rect 68294 1334 68328 1368
rect 69312 1334 69346 1368
rect 70330 1334 70364 1368
rect 71348 1334 71382 1368
rect 72366 1334 72400 1368
rect 73384 1334 73418 1368
rect 74402 1334 74436 1368
rect 41758 238 41792 272
rect 42776 238 42810 272
rect 43794 238 43828 272
rect 44812 238 44846 272
rect 45830 238 45864 272
rect 46848 238 46882 272
rect 47866 238 47900 272
rect 48884 238 48918 272
rect 49902 238 49936 272
rect 50920 238 50954 272
rect 51938 238 51972 272
rect 55048 156 55082 190
rect 56066 156 56100 190
rect 57084 156 57118 190
rect 58102 156 58136 190
rect 59120 156 59154 190
rect 60138 156 60172 190
rect 61156 156 61190 190
rect 62174 156 62208 190
rect 63192 156 63226 190
rect 64210 156 64244 190
rect 65228 156 65262 190
rect 66246 156 66280 190
rect 67264 156 67298 190
rect 68282 156 68316 190
rect 69300 156 69334 190
rect 70318 156 70352 190
rect 71336 156 71370 190
rect 72354 156 72388 190
rect 73372 156 73406 190
rect 74390 156 74424 190
rect 76772 -690 76872 15030
rect 39790 -852 76710 -752
<< nsubdiffcont >>
rect 11490 30592 35610 30692
rect 11328 16184 11428 30530
rect 17946 28114 17980 28148
rect 18964 28114 18998 28148
rect 19982 28114 20016 28148
rect 21000 28114 21034 28148
rect 22018 28114 22052 28148
rect 23036 28114 23070 28148
rect 24054 28114 24088 28148
rect 25072 28114 25106 28148
rect 26090 28114 26124 28148
rect 27108 28114 27142 28148
rect 28126 28114 28160 28148
rect 29144 28114 29178 28148
rect 30162 28114 30196 28148
rect 31180 28114 31214 28148
rect 32198 28114 32232 28148
rect 33216 28114 33250 28148
rect 17968 26960 18002 26994
rect 18986 26960 19020 26994
rect 20004 26960 20038 26994
rect 21022 26960 21056 26994
rect 22040 26960 22074 26994
rect 23058 26960 23092 26994
rect 24076 26960 24110 26994
rect 25094 26960 25128 26994
rect 26112 26960 26146 26994
rect 27130 26960 27164 26994
rect 28148 26960 28182 26994
rect 29166 26960 29200 26994
rect 30184 26960 30218 26994
rect 31202 26960 31236 26994
rect 32220 26960 32254 26994
rect 33238 26960 33272 26994
rect 17946 25828 17980 25862
rect 18964 25828 18998 25862
rect 19982 25828 20016 25862
rect 21000 25828 21034 25862
rect 22018 25828 22052 25862
rect 23036 25828 23070 25862
rect 24054 25828 24088 25862
rect 25072 25828 25106 25862
rect 26090 25828 26124 25862
rect 27108 25828 27142 25862
rect 28126 25828 28160 25862
rect 29144 25828 29178 25862
rect 30162 25828 30196 25862
rect 31180 25828 31214 25862
rect 32198 25828 32232 25862
rect 33216 25828 33250 25862
rect 17946 24446 17980 24480
rect 18964 24446 18998 24480
rect 19982 24446 20016 24480
rect 21000 24446 21034 24480
rect 22018 24446 22052 24480
rect 23036 24446 23070 24480
rect 24054 24446 24088 24480
rect 25072 24446 25106 24480
rect 26090 24446 26124 24480
rect 27108 24446 27142 24480
rect 28126 24446 28160 24480
rect 29144 24446 29178 24480
rect 30162 24446 30196 24480
rect 31180 24446 31214 24480
rect 32198 24446 32232 24480
rect 33216 24446 33250 24480
rect 18634 23098 18668 23132
rect 19652 23098 19686 23132
rect 20670 23098 20704 23132
rect 21688 23098 21722 23132
rect 22706 23098 22740 23132
rect 23724 23098 23758 23132
rect 24742 23098 24776 23132
rect 25760 23098 25794 23132
rect 26778 23098 26812 23132
rect 27796 23098 27830 23132
rect 28814 23098 28848 23132
rect 29832 23098 29866 23132
rect 30850 23098 30884 23132
rect 31868 23098 31902 23132
rect 32886 23098 32920 23132
rect 18240 21820 18274 21854
rect 19258 21820 19292 21854
rect 20276 21820 20310 21854
rect 21294 21820 21328 21854
rect 22312 21820 22346 21854
rect 23330 21820 23364 21854
rect 24348 21820 24382 21854
rect 25366 21820 25400 21854
rect 26384 21820 26418 21854
rect 27402 21820 27436 21854
rect 28420 21820 28454 21854
rect 29438 21820 29472 21854
rect 30456 21820 30490 21854
rect 31474 21820 31508 21854
rect 32492 21820 32526 21854
rect 33510 21820 33544 21854
rect 13642 21510 13676 21544
rect 14660 21510 14694 21544
rect 15678 21510 15712 21544
rect 16696 21510 16730 21544
rect 13118 20356 13152 20390
rect 14136 20356 14170 20390
rect 15154 20356 15188 20390
rect 16172 20356 16206 20390
rect 18330 20372 18364 20406
rect 19348 20372 19382 20406
rect 20366 20372 20400 20406
rect 21384 20372 21418 20406
rect 22402 20372 22436 20406
rect 23420 20372 23454 20406
rect 24438 20372 24472 20406
rect 25456 20372 25490 20406
rect 26474 20372 26508 20406
rect 27492 20372 27526 20406
rect 28510 20372 28544 20406
rect 29528 20372 29562 20406
rect 30546 20372 30580 20406
rect 31564 20372 31598 20406
rect 32582 20372 32616 20406
rect 33600 20372 33634 20406
rect 13128 19328 13162 19362
rect 14146 19328 14180 19362
rect 15164 19328 15198 19362
rect 16182 19328 16216 19362
rect 18354 19104 18388 19138
rect 19372 19104 19406 19138
rect 20390 19104 20424 19138
rect 21408 19104 21442 19138
rect 22426 19104 22460 19138
rect 23444 19104 23478 19138
rect 24462 19104 24496 19138
rect 25480 19104 25514 19138
rect 26498 19104 26532 19138
rect 27516 19104 27550 19138
rect 28534 19104 28568 19138
rect 29552 19104 29586 19138
rect 30570 19104 30604 19138
rect 31588 19104 31622 19138
rect 32606 19104 32640 19138
rect 33624 19104 33658 19138
rect 13118 18300 13152 18334
rect 14136 18300 14170 18334
rect 15154 18300 15188 18334
rect 16172 18300 16206 18334
rect 18218 17860 18252 17894
rect 19236 17860 19270 17894
rect 20254 17860 20288 17894
rect 21272 17860 21306 17894
rect 22290 17860 22324 17894
rect 23308 17860 23342 17894
rect 24326 17860 24360 17894
rect 25344 17860 25378 17894
rect 26362 17860 26396 17894
rect 27380 17860 27414 17894
rect 28398 17860 28432 17894
rect 29416 17860 29450 17894
rect 30434 17860 30468 17894
rect 31452 17860 31486 17894
rect 32470 17860 32504 17894
rect 33488 17860 33522 17894
rect 13642 17148 13676 17182
rect 14660 17148 14694 17182
rect 15678 17148 15712 17182
rect 16696 17148 16730 17182
rect 35672 16184 35772 30530
rect 11490 16022 35610 16122
rect 52490 30592 76610 30692
rect 52328 16184 52428 30530
rect 58946 28114 58980 28148
rect 59964 28114 59998 28148
rect 60982 28114 61016 28148
rect 62000 28114 62034 28148
rect 63018 28114 63052 28148
rect 64036 28114 64070 28148
rect 65054 28114 65088 28148
rect 66072 28114 66106 28148
rect 67090 28114 67124 28148
rect 68108 28114 68142 28148
rect 69126 28114 69160 28148
rect 70144 28114 70178 28148
rect 71162 28114 71196 28148
rect 72180 28114 72214 28148
rect 73198 28114 73232 28148
rect 74216 28114 74250 28148
rect 58968 26960 59002 26994
rect 59986 26960 60020 26994
rect 61004 26960 61038 26994
rect 62022 26960 62056 26994
rect 63040 26960 63074 26994
rect 64058 26960 64092 26994
rect 65076 26960 65110 26994
rect 66094 26960 66128 26994
rect 67112 26960 67146 26994
rect 68130 26960 68164 26994
rect 69148 26960 69182 26994
rect 70166 26960 70200 26994
rect 71184 26960 71218 26994
rect 72202 26960 72236 26994
rect 73220 26960 73254 26994
rect 74238 26960 74272 26994
rect 58946 25828 58980 25862
rect 59964 25828 59998 25862
rect 60982 25828 61016 25862
rect 62000 25828 62034 25862
rect 63018 25828 63052 25862
rect 64036 25828 64070 25862
rect 65054 25828 65088 25862
rect 66072 25828 66106 25862
rect 67090 25828 67124 25862
rect 68108 25828 68142 25862
rect 69126 25828 69160 25862
rect 70144 25828 70178 25862
rect 71162 25828 71196 25862
rect 72180 25828 72214 25862
rect 73198 25828 73232 25862
rect 74216 25828 74250 25862
rect 58946 24446 58980 24480
rect 59964 24446 59998 24480
rect 60982 24446 61016 24480
rect 62000 24446 62034 24480
rect 63018 24446 63052 24480
rect 64036 24446 64070 24480
rect 65054 24446 65088 24480
rect 66072 24446 66106 24480
rect 67090 24446 67124 24480
rect 68108 24446 68142 24480
rect 69126 24446 69160 24480
rect 70144 24446 70178 24480
rect 71162 24446 71196 24480
rect 72180 24446 72214 24480
rect 73198 24446 73232 24480
rect 74216 24446 74250 24480
rect 59634 23098 59668 23132
rect 60652 23098 60686 23132
rect 61670 23098 61704 23132
rect 62688 23098 62722 23132
rect 63706 23098 63740 23132
rect 64724 23098 64758 23132
rect 65742 23098 65776 23132
rect 66760 23098 66794 23132
rect 67778 23098 67812 23132
rect 68796 23098 68830 23132
rect 69814 23098 69848 23132
rect 70832 23098 70866 23132
rect 71850 23098 71884 23132
rect 72868 23098 72902 23132
rect 73886 23098 73920 23132
rect 59240 21820 59274 21854
rect 60258 21820 60292 21854
rect 61276 21820 61310 21854
rect 62294 21820 62328 21854
rect 63312 21820 63346 21854
rect 64330 21820 64364 21854
rect 65348 21820 65382 21854
rect 66366 21820 66400 21854
rect 67384 21820 67418 21854
rect 68402 21820 68436 21854
rect 69420 21820 69454 21854
rect 70438 21820 70472 21854
rect 71456 21820 71490 21854
rect 72474 21820 72508 21854
rect 73492 21820 73526 21854
rect 74510 21820 74544 21854
rect 54642 21510 54676 21544
rect 55660 21510 55694 21544
rect 56678 21510 56712 21544
rect 57696 21510 57730 21544
rect 54118 20356 54152 20390
rect 55136 20356 55170 20390
rect 56154 20356 56188 20390
rect 57172 20356 57206 20390
rect 59330 20372 59364 20406
rect 60348 20372 60382 20406
rect 61366 20372 61400 20406
rect 62384 20372 62418 20406
rect 63402 20372 63436 20406
rect 64420 20372 64454 20406
rect 65438 20372 65472 20406
rect 66456 20372 66490 20406
rect 67474 20372 67508 20406
rect 68492 20372 68526 20406
rect 69510 20372 69544 20406
rect 70528 20372 70562 20406
rect 71546 20372 71580 20406
rect 72564 20372 72598 20406
rect 73582 20372 73616 20406
rect 74600 20372 74634 20406
rect 54128 19328 54162 19362
rect 55146 19328 55180 19362
rect 56164 19328 56198 19362
rect 57182 19328 57216 19362
rect 59354 19104 59388 19138
rect 60372 19104 60406 19138
rect 61390 19104 61424 19138
rect 62408 19104 62442 19138
rect 63426 19104 63460 19138
rect 64444 19104 64478 19138
rect 65462 19104 65496 19138
rect 66480 19104 66514 19138
rect 67498 19104 67532 19138
rect 68516 19104 68550 19138
rect 69534 19104 69568 19138
rect 70552 19104 70586 19138
rect 71570 19104 71604 19138
rect 72588 19104 72622 19138
rect 73606 19104 73640 19138
rect 74624 19104 74658 19138
rect 54118 18300 54152 18334
rect 55136 18300 55170 18334
rect 56154 18300 56188 18334
rect 57172 18300 57206 18334
rect 59218 17860 59252 17894
rect 60236 17860 60270 17894
rect 61254 17860 61288 17894
rect 62272 17860 62306 17894
rect 63290 17860 63324 17894
rect 64308 17860 64342 17894
rect 65326 17860 65360 17894
rect 66344 17860 66378 17894
rect 67362 17860 67396 17894
rect 68380 17860 68414 17894
rect 69398 17860 69432 17894
rect 70416 17860 70450 17894
rect 71434 17860 71468 17894
rect 72452 17860 72486 17894
rect 73470 17860 73504 17894
rect 74488 17860 74522 17894
rect 54642 17148 54676 17182
rect 55660 17148 55694 17182
rect 56678 17148 56712 17182
rect 57696 17148 57730 17182
rect 76672 16184 76772 30530
rect 52490 16022 76610 16122
rect 36880 13870 38520 13970
rect 36718 12588 36818 13808
rect 38582 12588 38682 13808
rect 36880 12426 38520 12526
<< poly >>
rect 17670 27925 18258 27941
rect 17670 27908 17686 27925
rect 17484 27891 17686 27908
rect 18242 27908 18258 27925
rect 18688 27925 19276 27941
rect 18688 27908 18704 27925
rect 18242 27891 18444 27908
rect 17484 27844 18444 27891
rect 18502 27891 18704 27908
rect 19260 27908 19276 27925
rect 19706 27925 20294 27941
rect 19706 27908 19722 27925
rect 19260 27891 19462 27908
rect 18502 27844 19462 27891
rect 19520 27891 19722 27908
rect 20278 27908 20294 27925
rect 20724 27925 21312 27941
rect 20724 27908 20740 27925
rect 20278 27891 20480 27908
rect 19520 27844 20480 27891
rect 20538 27891 20740 27908
rect 21296 27908 21312 27925
rect 21742 27925 22330 27941
rect 21742 27908 21758 27925
rect 21296 27891 21498 27908
rect 20538 27844 21498 27891
rect 21556 27891 21758 27908
rect 22314 27908 22330 27925
rect 22760 27925 23348 27941
rect 22760 27908 22776 27925
rect 22314 27891 22516 27908
rect 21556 27844 22516 27891
rect 22574 27891 22776 27908
rect 23332 27908 23348 27925
rect 23778 27925 24366 27941
rect 23778 27908 23794 27925
rect 23332 27891 23534 27908
rect 22574 27844 23534 27891
rect 23592 27891 23794 27908
rect 24350 27908 24366 27925
rect 24796 27925 25384 27941
rect 24796 27908 24812 27925
rect 24350 27891 24552 27908
rect 23592 27844 24552 27891
rect 24610 27891 24812 27908
rect 25368 27908 25384 27925
rect 25814 27925 26402 27941
rect 25814 27908 25830 27925
rect 25368 27891 25570 27908
rect 24610 27844 25570 27891
rect 25628 27891 25830 27908
rect 26386 27908 26402 27925
rect 26832 27925 27420 27941
rect 26832 27908 26848 27925
rect 26386 27891 26588 27908
rect 25628 27844 26588 27891
rect 26646 27891 26848 27908
rect 27404 27908 27420 27925
rect 27850 27925 28438 27941
rect 27850 27908 27866 27925
rect 27404 27891 27606 27908
rect 26646 27844 27606 27891
rect 27664 27891 27866 27908
rect 28422 27908 28438 27925
rect 28868 27925 29456 27941
rect 28868 27908 28884 27925
rect 28422 27891 28624 27908
rect 27664 27844 28624 27891
rect 28682 27891 28884 27908
rect 29440 27908 29456 27925
rect 29886 27925 30474 27941
rect 29886 27908 29902 27925
rect 29440 27891 29642 27908
rect 28682 27844 29642 27891
rect 29700 27891 29902 27908
rect 30458 27908 30474 27925
rect 30904 27925 31492 27941
rect 30904 27908 30920 27925
rect 30458 27891 30660 27908
rect 29700 27844 30660 27891
rect 30718 27891 30920 27908
rect 31476 27908 31492 27925
rect 31922 27925 32510 27941
rect 31922 27908 31938 27925
rect 31476 27891 31678 27908
rect 30718 27844 31678 27891
rect 31736 27891 31938 27908
rect 32494 27908 32510 27925
rect 32940 27925 33528 27941
rect 32940 27908 32956 27925
rect 32494 27891 32696 27908
rect 31736 27844 32696 27891
rect 32754 27891 32956 27908
rect 33512 27908 33528 27925
rect 33512 27891 33714 27908
rect 32754 27844 33714 27891
rect 17484 27197 18444 27244
rect 17484 27180 17686 27197
rect 17670 27163 17686 27180
rect 18242 27180 18444 27197
rect 18502 27197 19462 27244
rect 18502 27180 18704 27197
rect 18242 27163 18258 27180
rect 17670 27147 18258 27163
rect 18688 27163 18704 27180
rect 19260 27180 19462 27197
rect 19520 27197 20480 27244
rect 19520 27180 19722 27197
rect 19260 27163 19276 27180
rect 18688 27147 19276 27163
rect 19706 27163 19722 27180
rect 20278 27180 20480 27197
rect 20538 27197 21498 27244
rect 20538 27180 20740 27197
rect 20278 27163 20294 27180
rect 19706 27147 20294 27163
rect 20724 27163 20740 27180
rect 21296 27180 21498 27197
rect 21556 27197 22516 27244
rect 21556 27180 21758 27197
rect 21296 27163 21312 27180
rect 20724 27147 21312 27163
rect 21742 27163 21758 27180
rect 22314 27180 22516 27197
rect 22574 27197 23534 27244
rect 22574 27180 22776 27197
rect 22314 27163 22330 27180
rect 21742 27147 22330 27163
rect 22760 27163 22776 27180
rect 23332 27180 23534 27197
rect 23592 27197 24552 27244
rect 23592 27180 23794 27197
rect 23332 27163 23348 27180
rect 22760 27147 23348 27163
rect 23778 27163 23794 27180
rect 24350 27180 24552 27197
rect 24610 27197 25570 27244
rect 24610 27180 24812 27197
rect 24350 27163 24366 27180
rect 23778 27147 24366 27163
rect 24796 27163 24812 27180
rect 25368 27180 25570 27197
rect 25628 27197 26588 27244
rect 25628 27180 25830 27197
rect 25368 27163 25384 27180
rect 24796 27147 25384 27163
rect 25814 27163 25830 27180
rect 26386 27180 26588 27197
rect 26646 27197 27606 27244
rect 26646 27180 26848 27197
rect 26386 27163 26402 27180
rect 25814 27147 26402 27163
rect 26832 27163 26848 27180
rect 27404 27180 27606 27197
rect 27664 27197 28624 27244
rect 27664 27180 27866 27197
rect 27404 27163 27420 27180
rect 26832 27147 27420 27163
rect 27850 27163 27866 27180
rect 28422 27180 28624 27197
rect 28682 27197 29642 27244
rect 28682 27180 28884 27197
rect 28422 27163 28438 27180
rect 27850 27147 28438 27163
rect 28868 27163 28884 27180
rect 29440 27180 29642 27197
rect 29700 27197 30660 27244
rect 29700 27180 29902 27197
rect 29440 27163 29456 27180
rect 28868 27147 29456 27163
rect 29886 27163 29902 27180
rect 30458 27180 30660 27197
rect 30718 27197 31678 27244
rect 30718 27180 30920 27197
rect 30458 27163 30474 27180
rect 29886 27147 30474 27163
rect 30904 27163 30920 27180
rect 31476 27180 31678 27197
rect 31736 27197 32696 27244
rect 31736 27180 31938 27197
rect 31476 27163 31492 27180
rect 30904 27147 31492 27163
rect 31922 27163 31938 27180
rect 32494 27180 32696 27197
rect 32754 27197 33714 27244
rect 32754 27180 32956 27197
rect 32494 27163 32510 27180
rect 31922 27147 32510 27163
rect 32940 27163 32956 27180
rect 33512 27180 33714 27197
rect 33512 27163 33528 27180
rect 32940 27147 33528 27163
rect 17670 26789 18258 26805
rect 17670 26772 17686 26789
rect 17484 26755 17686 26772
rect 18242 26772 18258 26789
rect 18688 26789 19276 26805
rect 18688 26772 18704 26789
rect 18242 26755 18444 26772
rect 17484 26708 18444 26755
rect 18502 26755 18704 26772
rect 19260 26772 19276 26789
rect 19706 26789 20294 26805
rect 19706 26772 19722 26789
rect 19260 26755 19462 26772
rect 18502 26708 19462 26755
rect 19520 26755 19722 26772
rect 20278 26772 20294 26789
rect 20724 26789 21312 26805
rect 20724 26772 20740 26789
rect 20278 26755 20480 26772
rect 19520 26708 20480 26755
rect 20538 26755 20740 26772
rect 21296 26772 21312 26789
rect 21742 26789 22330 26805
rect 21742 26772 21758 26789
rect 21296 26755 21498 26772
rect 20538 26708 21498 26755
rect 21556 26755 21758 26772
rect 22314 26772 22330 26789
rect 22760 26789 23348 26805
rect 22760 26772 22776 26789
rect 22314 26755 22516 26772
rect 21556 26708 22516 26755
rect 22574 26755 22776 26772
rect 23332 26772 23348 26789
rect 23778 26789 24366 26805
rect 23778 26772 23794 26789
rect 23332 26755 23534 26772
rect 22574 26708 23534 26755
rect 23592 26755 23794 26772
rect 24350 26772 24366 26789
rect 24796 26789 25384 26805
rect 24796 26772 24812 26789
rect 24350 26755 24552 26772
rect 23592 26708 24552 26755
rect 24610 26755 24812 26772
rect 25368 26772 25384 26789
rect 25814 26789 26402 26805
rect 25814 26772 25830 26789
rect 25368 26755 25570 26772
rect 24610 26708 25570 26755
rect 25628 26755 25830 26772
rect 26386 26772 26402 26789
rect 26832 26789 27420 26805
rect 26832 26772 26848 26789
rect 26386 26755 26588 26772
rect 25628 26708 26588 26755
rect 26646 26755 26848 26772
rect 27404 26772 27420 26789
rect 27850 26789 28438 26805
rect 27850 26772 27866 26789
rect 27404 26755 27606 26772
rect 26646 26708 27606 26755
rect 27664 26755 27866 26772
rect 28422 26772 28438 26789
rect 28868 26789 29456 26805
rect 28868 26772 28884 26789
rect 28422 26755 28624 26772
rect 27664 26708 28624 26755
rect 28682 26755 28884 26772
rect 29440 26772 29456 26789
rect 29886 26789 30474 26805
rect 29886 26772 29902 26789
rect 29440 26755 29642 26772
rect 28682 26708 29642 26755
rect 29700 26755 29902 26772
rect 30458 26772 30474 26789
rect 30904 26789 31492 26805
rect 30904 26772 30920 26789
rect 30458 26755 30660 26772
rect 29700 26708 30660 26755
rect 30718 26755 30920 26772
rect 31476 26772 31492 26789
rect 31922 26789 32510 26805
rect 31922 26772 31938 26789
rect 31476 26755 31678 26772
rect 30718 26708 31678 26755
rect 31736 26755 31938 26772
rect 32494 26772 32510 26789
rect 32940 26789 33528 26805
rect 32940 26772 32956 26789
rect 32494 26755 32696 26772
rect 31736 26708 32696 26755
rect 32754 26755 32956 26772
rect 33512 26772 33528 26789
rect 33512 26755 33714 26772
rect 32754 26708 33714 26755
rect 17484 26061 18444 26108
rect 17484 26044 17686 26061
rect 17670 26027 17686 26044
rect 18242 26044 18444 26061
rect 18502 26061 19462 26108
rect 18502 26044 18704 26061
rect 18242 26027 18258 26044
rect 17670 26011 18258 26027
rect 18688 26027 18704 26044
rect 19260 26044 19462 26061
rect 19520 26061 20480 26108
rect 19520 26044 19722 26061
rect 19260 26027 19276 26044
rect 18688 26011 19276 26027
rect 19706 26027 19722 26044
rect 20278 26044 20480 26061
rect 20538 26061 21498 26108
rect 20538 26044 20740 26061
rect 20278 26027 20294 26044
rect 19706 26011 20294 26027
rect 20724 26027 20740 26044
rect 21296 26044 21498 26061
rect 21556 26061 22516 26108
rect 21556 26044 21758 26061
rect 21296 26027 21312 26044
rect 20724 26011 21312 26027
rect 21742 26027 21758 26044
rect 22314 26044 22516 26061
rect 22574 26061 23534 26108
rect 22574 26044 22776 26061
rect 22314 26027 22330 26044
rect 21742 26011 22330 26027
rect 22760 26027 22776 26044
rect 23332 26044 23534 26061
rect 23592 26061 24552 26108
rect 23592 26044 23794 26061
rect 23332 26027 23348 26044
rect 22760 26011 23348 26027
rect 23778 26027 23794 26044
rect 24350 26044 24552 26061
rect 24610 26061 25570 26108
rect 24610 26044 24812 26061
rect 24350 26027 24366 26044
rect 23778 26011 24366 26027
rect 24796 26027 24812 26044
rect 25368 26044 25570 26061
rect 25628 26061 26588 26108
rect 25628 26044 25830 26061
rect 25368 26027 25384 26044
rect 24796 26011 25384 26027
rect 25814 26027 25830 26044
rect 26386 26044 26588 26061
rect 26646 26061 27606 26108
rect 26646 26044 26848 26061
rect 26386 26027 26402 26044
rect 25814 26011 26402 26027
rect 26832 26027 26848 26044
rect 27404 26044 27606 26061
rect 27664 26061 28624 26108
rect 27664 26044 27866 26061
rect 27404 26027 27420 26044
rect 26832 26011 27420 26027
rect 27850 26027 27866 26044
rect 28422 26044 28624 26061
rect 28682 26061 29642 26108
rect 28682 26044 28884 26061
rect 28422 26027 28438 26044
rect 27850 26011 28438 26027
rect 28868 26027 28884 26044
rect 29440 26044 29642 26061
rect 29700 26061 30660 26108
rect 29700 26044 29902 26061
rect 29440 26027 29456 26044
rect 28868 26011 29456 26027
rect 29886 26027 29902 26044
rect 30458 26044 30660 26061
rect 30718 26061 31678 26108
rect 30718 26044 30920 26061
rect 30458 26027 30474 26044
rect 29886 26011 30474 26027
rect 30904 26027 30920 26044
rect 31476 26044 31678 26061
rect 31736 26061 32696 26108
rect 31736 26044 31938 26061
rect 31476 26027 31492 26044
rect 30904 26011 31492 26027
rect 31922 26027 31938 26044
rect 32494 26044 32696 26061
rect 32754 26061 33714 26108
rect 32754 26044 32956 26061
rect 32494 26027 32510 26044
rect 31922 26011 32510 26027
rect 32940 26027 32956 26044
rect 33512 26044 33714 26061
rect 33512 26027 33528 26044
rect 32940 26011 33528 26027
rect 17670 25653 18258 25669
rect 17670 25636 17686 25653
rect 17484 25619 17686 25636
rect 18242 25636 18258 25653
rect 18688 25653 19276 25669
rect 18688 25636 18704 25653
rect 18242 25619 18444 25636
rect 17484 25572 18444 25619
rect 18502 25619 18704 25636
rect 19260 25636 19276 25653
rect 19706 25653 20294 25669
rect 19706 25636 19722 25653
rect 19260 25619 19462 25636
rect 18502 25572 19462 25619
rect 19520 25619 19722 25636
rect 20278 25636 20294 25653
rect 20724 25653 21312 25669
rect 20724 25636 20740 25653
rect 20278 25619 20480 25636
rect 19520 25572 20480 25619
rect 20538 25619 20740 25636
rect 21296 25636 21312 25653
rect 21742 25653 22330 25669
rect 21742 25636 21758 25653
rect 21296 25619 21498 25636
rect 20538 25572 21498 25619
rect 21556 25619 21758 25636
rect 22314 25636 22330 25653
rect 22760 25653 23348 25669
rect 22760 25636 22776 25653
rect 22314 25619 22516 25636
rect 21556 25572 22516 25619
rect 22574 25619 22776 25636
rect 23332 25636 23348 25653
rect 23778 25653 24366 25669
rect 23778 25636 23794 25653
rect 23332 25619 23534 25636
rect 22574 25572 23534 25619
rect 23592 25619 23794 25636
rect 24350 25636 24366 25653
rect 24796 25653 25384 25669
rect 24796 25636 24812 25653
rect 24350 25619 24552 25636
rect 23592 25572 24552 25619
rect 24610 25619 24812 25636
rect 25368 25636 25384 25653
rect 25814 25653 26402 25669
rect 25814 25636 25830 25653
rect 25368 25619 25570 25636
rect 24610 25572 25570 25619
rect 25628 25619 25830 25636
rect 26386 25636 26402 25653
rect 26832 25653 27420 25669
rect 26832 25636 26848 25653
rect 26386 25619 26588 25636
rect 25628 25572 26588 25619
rect 26646 25619 26848 25636
rect 27404 25636 27420 25653
rect 27850 25653 28438 25669
rect 27850 25636 27866 25653
rect 27404 25619 27606 25636
rect 26646 25572 27606 25619
rect 27664 25619 27866 25636
rect 28422 25636 28438 25653
rect 28868 25653 29456 25669
rect 28868 25636 28884 25653
rect 28422 25619 28624 25636
rect 27664 25572 28624 25619
rect 28682 25619 28884 25636
rect 29440 25636 29456 25653
rect 29886 25653 30474 25669
rect 29886 25636 29902 25653
rect 29440 25619 29642 25636
rect 28682 25572 29642 25619
rect 29700 25619 29902 25636
rect 30458 25636 30474 25653
rect 30904 25653 31492 25669
rect 30904 25636 30920 25653
rect 30458 25619 30660 25636
rect 29700 25572 30660 25619
rect 30718 25619 30920 25636
rect 31476 25636 31492 25653
rect 31922 25653 32510 25669
rect 31922 25636 31938 25653
rect 31476 25619 31678 25636
rect 30718 25572 31678 25619
rect 31736 25619 31938 25636
rect 32494 25636 32510 25653
rect 32940 25653 33528 25669
rect 32940 25636 32956 25653
rect 32494 25619 32696 25636
rect 31736 25572 32696 25619
rect 32754 25619 32956 25636
rect 33512 25636 33528 25653
rect 33512 25619 33714 25636
rect 32754 25572 33714 25619
rect 17484 24925 18444 24972
rect 17484 24908 17686 24925
rect 17670 24891 17686 24908
rect 18242 24908 18444 24925
rect 18502 24925 19462 24972
rect 18502 24908 18704 24925
rect 18242 24891 18258 24908
rect 17670 24875 18258 24891
rect 18688 24891 18704 24908
rect 19260 24908 19462 24925
rect 19520 24925 20480 24972
rect 19520 24908 19722 24925
rect 19260 24891 19276 24908
rect 18688 24875 19276 24891
rect 19706 24891 19722 24908
rect 20278 24908 20480 24925
rect 20538 24925 21498 24972
rect 20538 24908 20740 24925
rect 20278 24891 20294 24908
rect 19706 24875 20294 24891
rect 20724 24891 20740 24908
rect 21296 24908 21498 24925
rect 21556 24925 22516 24972
rect 21556 24908 21758 24925
rect 21296 24891 21312 24908
rect 20724 24875 21312 24891
rect 21742 24891 21758 24908
rect 22314 24908 22516 24925
rect 22574 24925 23534 24972
rect 22574 24908 22776 24925
rect 22314 24891 22330 24908
rect 21742 24875 22330 24891
rect 22760 24891 22776 24908
rect 23332 24908 23534 24925
rect 23592 24925 24552 24972
rect 23592 24908 23794 24925
rect 23332 24891 23348 24908
rect 22760 24875 23348 24891
rect 23778 24891 23794 24908
rect 24350 24908 24552 24925
rect 24610 24925 25570 24972
rect 24610 24908 24812 24925
rect 24350 24891 24366 24908
rect 23778 24875 24366 24891
rect 24796 24891 24812 24908
rect 25368 24908 25570 24925
rect 25628 24925 26588 24972
rect 25628 24908 25830 24925
rect 25368 24891 25384 24908
rect 24796 24875 25384 24891
rect 25814 24891 25830 24908
rect 26386 24908 26588 24925
rect 26646 24925 27606 24972
rect 26646 24908 26848 24925
rect 26386 24891 26402 24908
rect 25814 24875 26402 24891
rect 26832 24891 26848 24908
rect 27404 24908 27606 24925
rect 27664 24925 28624 24972
rect 27664 24908 27866 24925
rect 27404 24891 27420 24908
rect 26832 24875 27420 24891
rect 27850 24891 27866 24908
rect 28422 24908 28624 24925
rect 28682 24925 29642 24972
rect 28682 24908 28884 24925
rect 28422 24891 28438 24908
rect 27850 24875 28438 24891
rect 28868 24891 28884 24908
rect 29440 24908 29642 24925
rect 29700 24925 30660 24972
rect 29700 24908 29902 24925
rect 29440 24891 29456 24908
rect 28868 24875 29456 24891
rect 29886 24891 29902 24908
rect 30458 24908 30660 24925
rect 30718 24925 31678 24972
rect 30718 24908 30920 24925
rect 30458 24891 30474 24908
rect 29886 24875 30474 24891
rect 30904 24891 30920 24908
rect 31476 24908 31678 24925
rect 31736 24925 32696 24972
rect 31736 24908 31938 24925
rect 31476 24891 31492 24908
rect 30904 24875 31492 24891
rect 31922 24891 31938 24908
rect 32494 24908 32696 24925
rect 32754 24925 33714 24972
rect 32754 24908 32956 24925
rect 32494 24891 32510 24908
rect 31922 24875 32510 24891
rect 32940 24891 32956 24908
rect 33512 24908 33714 24925
rect 33512 24891 33528 24908
rect 32940 24875 33528 24891
rect 18864 24015 19452 24031
rect 18864 23998 18880 24015
rect 18678 23981 18880 23998
rect 19436 23998 19452 24015
rect 19882 24015 20470 24031
rect 19882 23998 19898 24015
rect 19436 23981 19638 23998
rect 18678 23934 19638 23981
rect 19696 23981 19898 23998
rect 20454 23998 20470 24015
rect 20900 24015 21488 24031
rect 20900 23998 20916 24015
rect 20454 23981 20656 23998
rect 19696 23934 20656 23981
rect 20714 23981 20916 23998
rect 21472 23998 21488 24015
rect 21918 24015 22506 24031
rect 21918 23998 21934 24015
rect 21472 23981 21674 23998
rect 20714 23934 21674 23981
rect 21732 23981 21934 23998
rect 22490 23998 22506 24015
rect 22936 24015 23524 24031
rect 22936 23998 22952 24015
rect 22490 23981 22692 23998
rect 21732 23934 22692 23981
rect 22750 23981 22952 23998
rect 23508 23998 23524 24015
rect 23954 24015 24542 24031
rect 23954 23998 23970 24015
rect 23508 23981 23710 23998
rect 22750 23934 23710 23981
rect 23768 23981 23970 23998
rect 24526 23998 24542 24015
rect 24972 24015 25560 24031
rect 24972 23998 24988 24015
rect 24526 23981 24728 23998
rect 23768 23934 24728 23981
rect 24786 23981 24988 23998
rect 25544 23998 25560 24015
rect 25990 24015 26578 24031
rect 25990 23998 26006 24015
rect 25544 23981 25746 23998
rect 24786 23934 25746 23981
rect 25804 23981 26006 23998
rect 26562 23998 26578 24015
rect 27008 24015 27596 24031
rect 27008 23998 27024 24015
rect 26562 23981 26764 23998
rect 25804 23934 26764 23981
rect 26822 23981 27024 23998
rect 27580 23998 27596 24015
rect 28026 24015 28614 24031
rect 28026 23998 28042 24015
rect 27580 23981 27782 23998
rect 26822 23934 27782 23981
rect 27840 23981 28042 23998
rect 28598 23998 28614 24015
rect 29044 24015 29632 24031
rect 29044 23998 29060 24015
rect 28598 23981 28800 23998
rect 27840 23934 28800 23981
rect 28858 23981 29060 23998
rect 29616 23998 29632 24015
rect 30062 24015 30650 24031
rect 30062 23998 30078 24015
rect 29616 23981 29818 23998
rect 28858 23934 29818 23981
rect 29876 23981 30078 23998
rect 30634 23998 30650 24015
rect 31080 24015 31668 24031
rect 31080 23998 31096 24015
rect 30634 23981 30836 23998
rect 29876 23934 30836 23981
rect 30894 23981 31096 23998
rect 31652 23998 31668 24015
rect 32098 24015 32686 24031
rect 32098 23998 32114 24015
rect 31652 23981 31854 23998
rect 30894 23934 31854 23981
rect 31912 23981 32114 23998
rect 32670 23998 32686 24015
rect 32670 23981 32872 23998
rect 31912 23934 32872 23981
rect 18678 23287 19638 23334
rect 18678 23270 18880 23287
rect 18864 23253 18880 23270
rect 19436 23270 19638 23287
rect 19696 23287 20656 23334
rect 19696 23270 19898 23287
rect 19436 23253 19452 23270
rect 18864 23237 19452 23253
rect 19882 23253 19898 23270
rect 20454 23270 20656 23287
rect 20714 23287 21674 23334
rect 20714 23270 20916 23287
rect 20454 23253 20470 23270
rect 19882 23237 20470 23253
rect 20900 23253 20916 23270
rect 21472 23270 21674 23287
rect 21732 23287 22692 23334
rect 21732 23270 21934 23287
rect 21472 23253 21488 23270
rect 20900 23237 21488 23253
rect 21918 23253 21934 23270
rect 22490 23270 22692 23287
rect 22750 23287 23710 23334
rect 22750 23270 22952 23287
rect 22490 23253 22506 23270
rect 21918 23237 22506 23253
rect 22936 23253 22952 23270
rect 23508 23270 23710 23287
rect 23768 23287 24728 23334
rect 23768 23270 23970 23287
rect 23508 23253 23524 23270
rect 22936 23237 23524 23253
rect 23954 23253 23970 23270
rect 24526 23270 24728 23287
rect 24786 23287 25746 23334
rect 24786 23270 24988 23287
rect 24526 23253 24542 23270
rect 23954 23237 24542 23253
rect 24972 23253 24988 23270
rect 25544 23270 25746 23287
rect 25804 23287 26764 23334
rect 25804 23270 26006 23287
rect 25544 23253 25560 23270
rect 24972 23237 25560 23253
rect 25990 23253 26006 23270
rect 26562 23270 26764 23287
rect 26822 23287 27782 23334
rect 26822 23270 27024 23287
rect 26562 23253 26578 23270
rect 25990 23237 26578 23253
rect 27008 23253 27024 23270
rect 27580 23270 27782 23287
rect 27840 23287 28800 23334
rect 27840 23270 28042 23287
rect 27580 23253 27596 23270
rect 27008 23237 27596 23253
rect 28026 23253 28042 23270
rect 28598 23270 28800 23287
rect 28858 23287 29818 23334
rect 28858 23270 29060 23287
rect 28598 23253 28614 23270
rect 28026 23237 28614 23253
rect 29044 23253 29060 23270
rect 29616 23270 29818 23287
rect 29876 23287 30836 23334
rect 29876 23270 30078 23287
rect 29616 23253 29632 23270
rect 29044 23237 29632 23253
rect 30062 23253 30078 23270
rect 30634 23270 30836 23287
rect 30894 23287 31854 23334
rect 30894 23270 31096 23287
rect 30634 23253 30650 23270
rect 30062 23237 30650 23253
rect 31080 23253 31096 23270
rect 31652 23270 31854 23287
rect 31912 23287 32872 23334
rect 31912 23270 32114 23287
rect 31652 23253 31668 23270
rect 31080 23237 31668 23253
rect 32098 23253 32114 23270
rect 32670 23270 32872 23287
rect 32670 23253 32686 23270
rect 32098 23237 32686 23253
rect 18864 22983 19452 22999
rect 18864 22966 18880 22983
rect 18678 22949 18880 22966
rect 19436 22966 19452 22983
rect 19882 22983 20470 22999
rect 19882 22966 19898 22983
rect 19436 22949 19638 22966
rect 18678 22902 19638 22949
rect 19696 22949 19898 22966
rect 20454 22966 20470 22983
rect 20900 22983 21488 22999
rect 20900 22966 20916 22983
rect 20454 22949 20656 22966
rect 19696 22902 20656 22949
rect 20714 22949 20916 22966
rect 21472 22966 21488 22983
rect 21918 22983 22506 22999
rect 21918 22966 21934 22983
rect 21472 22949 21674 22966
rect 20714 22902 21674 22949
rect 21732 22949 21934 22966
rect 22490 22966 22506 22983
rect 22936 22983 23524 22999
rect 22936 22966 22952 22983
rect 22490 22949 22692 22966
rect 21732 22902 22692 22949
rect 22750 22949 22952 22966
rect 23508 22966 23524 22983
rect 23954 22983 24542 22999
rect 23954 22966 23970 22983
rect 23508 22949 23710 22966
rect 22750 22902 23710 22949
rect 23768 22949 23970 22966
rect 24526 22966 24542 22983
rect 24972 22983 25560 22999
rect 24972 22966 24988 22983
rect 24526 22949 24728 22966
rect 23768 22902 24728 22949
rect 24786 22949 24988 22966
rect 25544 22966 25560 22983
rect 25990 22983 26578 22999
rect 25990 22966 26006 22983
rect 25544 22949 25746 22966
rect 24786 22902 25746 22949
rect 25804 22949 26006 22966
rect 26562 22966 26578 22983
rect 27008 22983 27596 22999
rect 27008 22966 27024 22983
rect 26562 22949 26764 22966
rect 25804 22902 26764 22949
rect 26822 22949 27024 22966
rect 27580 22966 27596 22983
rect 28026 22983 28614 22999
rect 28026 22966 28042 22983
rect 27580 22949 27782 22966
rect 26822 22902 27782 22949
rect 27840 22949 28042 22966
rect 28598 22966 28614 22983
rect 29044 22983 29632 22999
rect 29044 22966 29060 22983
rect 28598 22949 28800 22966
rect 27840 22902 28800 22949
rect 28858 22949 29060 22966
rect 29616 22966 29632 22983
rect 30062 22983 30650 22999
rect 30062 22966 30078 22983
rect 29616 22949 29818 22966
rect 28858 22902 29818 22949
rect 29876 22949 30078 22966
rect 30634 22966 30650 22983
rect 31080 22983 31668 22999
rect 31080 22966 31096 22983
rect 30634 22949 30836 22966
rect 29876 22902 30836 22949
rect 30894 22949 31096 22966
rect 31652 22966 31668 22983
rect 32098 22983 32686 22999
rect 32098 22966 32114 22983
rect 31652 22949 31854 22966
rect 30894 22902 31854 22949
rect 31912 22949 32114 22966
rect 32670 22966 32686 22983
rect 32670 22949 32872 22966
rect 31912 22902 32872 22949
rect 18678 22255 19638 22302
rect 18678 22238 18880 22255
rect 18864 22221 18880 22238
rect 19436 22238 19638 22255
rect 19696 22255 20656 22302
rect 19696 22238 19898 22255
rect 19436 22221 19452 22238
rect 18864 22205 19452 22221
rect 19882 22221 19898 22238
rect 20454 22238 20656 22255
rect 20714 22255 21674 22302
rect 20714 22238 20916 22255
rect 20454 22221 20470 22238
rect 19882 22205 20470 22221
rect 20900 22221 20916 22238
rect 21472 22238 21674 22255
rect 21732 22255 22692 22302
rect 21732 22238 21934 22255
rect 21472 22221 21488 22238
rect 20900 22205 21488 22221
rect 21918 22221 21934 22238
rect 22490 22238 22692 22255
rect 22750 22255 23710 22302
rect 22750 22238 22952 22255
rect 22490 22221 22506 22238
rect 21918 22205 22506 22221
rect 22936 22221 22952 22238
rect 23508 22238 23710 22255
rect 23768 22255 24728 22302
rect 23768 22238 23970 22255
rect 23508 22221 23524 22238
rect 22936 22205 23524 22221
rect 23954 22221 23970 22238
rect 24526 22238 24728 22255
rect 24786 22255 25746 22302
rect 24786 22238 24988 22255
rect 24526 22221 24542 22238
rect 23954 22205 24542 22221
rect 24972 22221 24988 22238
rect 25544 22238 25746 22255
rect 25804 22255 26764 22302
rect 25804 22238 26006 22255
rect 25544 22221 25560 22238
rect 24972 22205 25560 22221
rect 25990 22221 26006 22238
rect 26562 22238 26764 22255
rect 26822 22255 27782 22302
rect 26822 22238 27024 22255
rect 26562 22221 26578 22238
rect 25990 22205 26578 22221
rect 27008 22221 27024 22238
rect 27580 22238 27782 22255
rect 27840 22255 28800 22302
rect 27840 22238 28042 22255
rect 27580 22221 27596 22238
rect 27008 22205 27596 22221
rect 28026 22221 28042 22238
rect 28598 22238 28800 22255
rect 28858 22255 29818 22302
rect 28858 22238 29060 22255
rect 28598 22221 28614 22238
rect 28026 22205 28614 22221
rect 29044 22221 29060 22238
rect 29616 22238 29818 22255
rect 29876 22255 30836 22302
rect 29876 22238 30078 22255
rect 29616 22221 29632 22238
rect 29044 22205 29632 22221
rect 30062 22221 30078 22238
rect 30634 22238 30836 22255
rect 30894 22255 31854 22302
rect 30894 22238 31096 22255
rect 30634 22221 30650 22238
rect 30062 22205 30650 22221
rect 31080 22221 31096 22238
rect 31652 22238 31854 22255
rect 31912 22255 32872 22302
rect 31912 22238 32114 22255
rect 31652 22221 31668 22238
rect 31080 22205 31668 22221
rect 32098 22221 32114 22238
rect 32670 22238 32872 22255
rect 32670 22221 32686 22238
rect 32098 22205 32686 22221
rect 18656 21379 19244 21395
rect 18656 21362 18672 21379
rect 18470 21345 18672 21362
rect 19228 21362 19244 21379
rect 19674 21379 20262 21395
rect 19674 21362 19690 21379
rect 19228 21345 19430 21362
rect 18470 21298 19430 21345
rect 19488 21345 19690 21362
rect 20246 21362 20262 21379
rect 20692 21379 21280 21395
rect 20692 21362 20708 21379
rect 20246 21345 20448 21362
rect 19488 21298 20448 21345
rect 20506 21345 20708 21362
rect 21264 21362 21280 21379
rect 21710 21379 22298 21395
rect 21710 21362 21726 21379
rect 21264 21345 21466 21362
rect 20506 21298 21466 21345
rect 21524 21345 21726 21362
rect 22282 21362 22298 21379
rect 22728 21379 23316 21395
rect 22728 21362 22744 21379
rect 22282 21345 22484 21362
rect 21524 21298 22484 21345
rect 22542 21345 22744 21362
rect 23300 21362 23316 21379
rect 23746 21379 24334 21395
rect 23746 21362 23762 21379
rect 23300 21345 23502 21362
rect 22542 21298 23502 21345
rect 23560 21345 23762 21362
rect 24318 21362 24334 21379
rect 24764 21379 25352 21395
rect 24764 21362 24780 21379
rect 24318 21345 24520 21362
rect 23560 21298 24520 21345
rect 24578 21345 24780 21362
rect 25336 21362 25352 21379
rect 25782 21379 26370 21395
rect 25782 21362 25798 21379
rect 25336 21345 25538 21362
rect 24578 21298 25538 21345
rect 25596 21345 25798 21362
rect 26354 21362 26370 21379
rect 26800 21379 27388 21395
rect 26800 21362 26816 21379
rect 26354 21345 26556 21362
rect 25596 21298 26556 21345
rect 26614 21345 26816 21362
rect 27372 21362 27388 21379
rect 27818 21379 28406 21395
rect 27818 21362 27834 21379
rect 27372 21345 27574 21362
rect 26614 21298 27574 21345
rect 27632 21345 27834 21362
rect 28390 21362 28406 21379
rect 28836 21379 29424 21395
rect 28836 21362 28852 21379
rect 28390 21345 28592 21362
rect 27632 21298 28592 21345
rect 28650 21345 28852 21362
rect 29408 21362 29424 21379
rect 29854 21379 30442 21395
rect 29854 21362 29870 21379
rect 29408 21345 29610 21362
rect 28650 21298 29610 21345
rect 29668 21345 29870 21362
rect 30426 21362 30442 21379
rect 30872 21379 31460 21395
rect 30872 21362 30888 21379
rect 30426 21345 30628 21362
rect 29668 21298 30628 21345
rect 30686 21345 30888 21362
rect 31444 21362 31460 21379
rect 31890 21379 32478 21395
rect 31890 21362 31906 21379
rect 31444 21345 31646 21362
rect 30686 21298 31646 21345
rect 31704 21345 31906 21362
rect 32462 21362 32478 21379
rect 32908 21379 33496 21395
rect 32908 21362 32924 21379
rect 32462 21345 32664 21362
rect 31704 21298 32664 21345
rect 32722 21345 32924 21362
rect 33480 21362 33496 21379
rect 33480 21345 33682 21362
rect 32722 21298 33682 21345
rect 13352 21275 13940 21291
rect 13352 21258 13368 21275
rect 13166 21241 13368 21258
rect 13924 21258 13940 21275
rect 14370 21275 14958 21291
rect 14370 21258 14386 21275
rect 13924 21241 14126 21258
rect 13166 21194 14126 21241
rect 14184 21241 14386 21258
rect 14942 21258 14958 21275
rect 15388 21275 15976 21291
rect 15388 21258 15404 21275
rect 14942 21241 15144 21258
rect 14184 21194 15144 21241
rect 15202 21241 15404 21258
rect 15960 21258 15976 21275
rect 16406 21275 16994 21291
rect 16406 21258 16422 21275
rect 15960 21241 16162 21258
rect 15202 21194 16162 21241
rect 16220 21241 16422 21258
rect 16978 21258 16994 21275
rect 16978 21241 17180 21258
rect 16220 21194 17180 21241
rect 18470 20651 19430 20698
rect 18470 20634 18672 20651
rect 18656 20617 18672 20634
rect 19228 20634 19430 20651
rect 19488 20651 20448 20698
rect 19488 20634 19690 20651
rect 19228 20617 19244 20634
rect 18656 20601 19244 20617
rect 19674 20617 19690 20634
rect 20246 20634 20448 20651
rect 20506 20651 21466 20698
rect 20506 20634 20708 20651
rect 20246 20617 20262 20634
rect 19674 20601 20262 20617
rect 20692 20617 20708 20634
rect 21264 20634 21466 20651
rect 21524 20651 22484 20698
rect 21524 20634 21726 20651
rect 21264 20617 21280 20634
rect 20692 20601 21280 20617
rect 21710 20617 21726 20634
rect 22282 20634 22484 20651
rect 22542 20651 23502 20698
rect 22542 20634 22744 20651
rect 22282 20617 22298 20634
rect 21710 20601 22298 20617
rect 22728 20617 22744 20634
rect 23300 20634 23502 20651
rect 23560 20651 24520 20698
rect 23560 20634 23762 20651
rect 23300 20617 23316 20634
rect 22728 20601 23316 20617
rect 23746 20617 23762 20634
rect 24318 20634 24520 20651
rect 24578 20651 25538 20698
rect 24578 20634 24780 20651
rect 24318 20617 24334 20634
rect 23746 20601 24334 20617
rect 24764 20617 24780 20634
rect 25336 20634 25538 20651
rect 25596 20651 26556 20698
rect 25596 20634 25798 20651
rect 25336 20617 25352 20634
rect 24764 20601 25352 20617
rect 25782 20617 25798 20634
rect 26354 20634 26556 20651
rect 26614 20651 27574 20698
rect 26614 20634 26816 20651
rect 26354 20617 26370 20634
rect 25782 20601 26370 20617
rect 26800 20617 26816 20634
rect 27372 20634 27574 20651
rect 27632 20651 28592 20698
rect 27632 20634 27834 20651
rect 27372 20617 27388 20634
rect 26800 20601 27388 20617
rect 27818 20617 27834 20634
rect 28390 20634 28592 20651
rect 28650 20651 29610 20698
rect 28650 20634 28852 20651
rect 28390 20617 28406 20634
rect 27818 20601 28406 20617
rect 28836 20617 28852 20634
rect 29408 20634 29610 20651
rect 29668 20651 30628 20698
rect 29668 20634 29870 20651
rect 29408 20617 29424 20634
rect 28836 20601 29424 20617
rect 29854 20617 29870 20634
rect 30426 20634 30628 20651
rect 30686 20651 31646 20698
rect 30686 20634 30888 20651
rect 30426 20617 30442 20634
rect 29854 20601 30442 20617
rect 30872 20617 30888 20634
rect 31444 20634 31646 20651
rect 31704 20651 32664 20698
rect 31704 20634 31906 20651
rect 31444 20617 31460 20634
rect 30872 20601 31460 20617
rect 31890 20617 31906 20634
rect 32462 20634 32664 20651
rect 32722 20651 33682 20698
rect 32722 20634 32924 20651
rect 32462 20617 32478 20634
rect 31890 20601 32478 20617
rect 32908 20617 32924 20634
rect 33480 20634 33682 20651
rect 33480 20617 33496 20634
rect 32908 20601 33496 20617
rect 13166 20547 14126 20594
rect 13166 20530 13368 20547
rect 13352 20513 13368 20530
rect 13924 20530 14126 20547
rect 14184 20547 15144 20594
rect 14184 20530 14386 20547
rect 13924 20513 13940 20530
rect 13352 20497 13940 20513
rect 14370 20513 14386 20530
rect 14942 20530 15144 20547
rect 15202 20547 16162 20594
rect 15202 20530 15404 20547
rect 14942 20513 14958 20530
rect 14370 20497 14958 20513
rect 15388 20513 15404 20530
rect 15960 20530 16162 20547
rect 16220 20547 17180 20594
rect 16220 20530 16422 20547
rect 15960 20513 15976 20530
rect 15388 20497 15976 20513
rect 16406 20513 16422 20530
rect 16978 20530 17180 20547
rect 16978 20513 16994 20530
rect 16406 20497 16994 20513
rect 13352 20243 13940 20259
rect 13352 20226 13368 20243
rect 13166 20209 13368 20226
rect 13924 20226 13940 20243
rect 14370 20243 14958 20259
rect 14370 20226 14386 20243
rect 13924 20209 14126 20226
rect 13166 20162 14126 20209
rect 14184 20209 14386 20226
rect 14942 20226 14958 20243
rect 15388 20243 15976 20259
rect 15388 20226 15404 20243
rect 14942 20209 15144 20226
rect 14184 20162 15144 20209
rect 15202 20209 15404 20226
rect 15960 20226 15976 20243
rect 16406 20243 16994 20259
rect 16406 20226 16422 20243
rect 15960 20209 16162 20226
rect 15202 20162 16162 20209
rect 16220 20209 16422 20226
rect 16978 20226 16994 20243
rect 16978 20209 17180 20226
rect 16220 20162 17180 20209
rect 18656 20123 19244 20139
rect 18656 20106 18672 20123
rect 18470 20089 18672 20106
rect 19228 20106 19244 20123
rect 19674 20123 20262 20139
rect 19674 20106 19690 20123
rect 19228 20089 19430 20106
rect 18470 20042 19430 20089
rect 19488 20089 19690 20106
rect 20246 20106 20262 20123
rect 20692 20123 21280 20139
rect 20692 20106 20708 20123
rect 20246 20089 20448 20106
rect 19488 20042 20448 20089
rect 20506 20089 20708 20106
rect 21264 20106 21280 20123
rect 21710 20123 22298 20139
rect 21710 20106 21726 20123
rect 21264 20089 21466 20106
rect 20506 20042 21466 20089
rect 21524 20089 21726 20106
rect 22282 20106 22298 20123
rect 22728 20123 23316 20139
rect 22728 20106 22744 20123
rect 22282 20089 22484 20106
rect 21524 20042 22484 20089
rect 22542 20089 22744 20106
rect 23300 20106 23316 20123
rect 23746 20123 24334 20139
rect 23746 20106 23762 20123
rect 23300 20089 23502 20106
rect 22542 20042 23502 20089
rect 23560 20089 23762 20106
rect 24318 20106 24334 20123
rect 24764 20123 25352 20139
rect 24764 20106 24780 20123
rect 24318 20089 24520 20106
rect 23560 20042 24520 20089
rect 24578 20089 24780 20106
rect 25336 20106 25352 20123
rect 25782 20123 26370 20139
rect 25782 20106 25798 20123
rect 25336 20089 25538 20106
rect 24578 20042 25538 20089
rect 25596 20089 25798 20106
rect 26354 20106 26370 20123
rect 26800 20123 27388 20139
rect 26800 20106 26816 20123
rect 26354 20089 26556 20106
rect 25596 20042 26556 20089
rect 26614 20089 26816 20106
rect 27372 20106 27388 20123
rect 27818 20123 28406 20139
rect 27818 20106 27834 20123
rect 27372 20089 27574 20106
rect 26614 20042 27574 20089
rect 27632 20089 27834 20106
rect 28390 20106 28406 20123
rect 28836 20123 29424 20139
rect 28836 20106 28852 20123
rect 28390 20089 28592 20106
rect 27632 20042 28592 20089
rect 28650 20089 28852 20106
rect 29408 20106 29424 20123
rect 29854 20123 30442 20139
rect 29854 20106 29870 20123
rect 29408 20089 29610 20106
rect 28650 20042 29610 20089
rect 29668 20089 29870 20106
rect 30426 20106 30442 20123
rect 30872 20123 31460 20139
rect 30872 20106 30888 20123
rect 30426 20089 30628 20106
rect 29668 20042 30628 20089
rect 30686 20089 30888 20106
rect 31444 20106 31460 20123
rect 31890 20123 32478 20139
rect 31890 20106 31906 20123
rect 31444 20089 31646 20106
rect 30686 20042 31646 20089
rect 31704 20089 31906 20106
rect 32462 20106 32478 20123
rect 32908 20123 33496 20139
rect 32908 20106 32924 20123
rect 32462 20089 32664 20106
rect 31704 20042 32664 20089
rect 32722 20089 32924 20106
rect 33480 20106 33496 20123
rect 33480 20089 33682 20106
rect 32722 20042 33682 20089
rect 13166 19515 14126 19562
rect 13166 19498 13368 19515
rect 13352 19481 13368 19498
rect 13924 19498 14126 19515
rect 14184 19515 15144 19562
rect 14184 19498 14386 19515
rect 13924 19481 13940 19498
rect 13352 19465 13940 19481
rect 14370 19481 14386 19498
rect 14942 19498 15144 19515
rect 15202 19515 16162 19562
rect 15202 19498 15404 19515
rect 14942 19481 14958 19498
rect 14370 19465 14958 19481
rect 15388 19481 15404 19498
rect 15960 19498 16162 19515
rect 16220 19515 17180 19562
rect 16220 19498 16422 19515
rect 15960 19481 15976 19498
rect 15388 19465 15976 19481
rect 16406 19481 16422 19498
rect 16978 19498 17180 19515
rect 16978 19481 16994 19498
rect 16406 19465 16994 19481
rect 18470 19395 19430 19442
rect 18470 19378 18672 19395
rect 18656 19361 18672 19378
rect 19228 19378 19430 19395
rect 19488 19395 20448 19442
rect 19488 19378 19690 19395
rect 19228 19361 19244 19378
rect 18656 19345 19244 19361
rect 19674 19361 19690 19378
rect 20246 19378 20448 19395
rect 20506 19395 21466 19442
rect 20506 19378 20708 19395
rect 20246 19361 20262 19378
rect 19674 19345 20262 19361
rect 20692 19361 20708 19378
rect 21264 19378 21466 19395
rect 21524 19395 22484 19442
rect 21524 19378 21726 19395
rect 21264 19361 21280 19378
rect 20692 19345 21280 19361
rect 21710 19361 21726 19378
rect 22282 19378 22484 19395
rect 22542 19395 23502 19442
rect 22542 19378 22744 19395
rect 22282 19361 22298 19378
rect 21710 19345 22298 19361
rect 22728 19361 22744 19378
rect 23300 19378 23502 19395
rect 23560 19395 24520 19442
rect 23560 19378 23762 19395
rect 23300 19361 23316 19378
rect 22728 19345 23316 19361
rect 23746 19361 23762 19378
rect 24318 19378 24520 19395
rect 24578 19395 25538 19442
rect 24578 19378 24780 19395
rect 24318 19361 24334 19378
rect 23746 19345 24334 19361
rect 24764 19361 24780 19378
rect 25336 19378 25538 19395
rect 25596 19395 26556 19442
rect 25596 19378 25798 19395
rect 25336 19361 25352 19378
rect 24764 19345 25352 19361
rect 25782 19361 25798 19378
rect 26354 19378 26556 19395
rect 26614 19395 27574 19442
rect 26614 19378 26816 19395
rect 26354 19361 26370 19378
rect 25782 19345 26370 19361
rect 26800 19361 26816 19378
rect 27372 19378 27574 19395
rect 27632 19395 28592 19442
rect 27632 19378 27834 19395
rect 27372 19361 27388 19378
rect 26800 19345 27388 19361
rect 27818 19361 27834 19378
rect 28390 19378 28592 19395
rect 28650 19395 29610 19442
rect 28650 19378 28852 19395
rect 28390 19361 28406 19378
rect 27818 19345 28406 19361
rect 28836 19361 28852 19378
rect 29408 19378 29610 19395
rect 29668 19395 30628 19442
rect 29668 19378 29870 19395
rect 29408 19361 29424 19378
rect 28836 19345 29424 19361
rect 29854 19361 29870 19378
rect 30426 19378 30628 19395
rect 30686 19395 31646 19442
rect 30686 19378 30888 19395
rect 30426 19361 30442 19378
rect 29854 19345 30442 19361
rect 30872 19361 30888 19378
rect 31444 19378 31646 19395
rect 31704 19395 32664 19442
rect 31704 19378 31906 19395
rect 31444 19361 31460 19378
rect 30872 19345 31460 19361
rect 31890 19361 31906 19378
rect 32462 19378 32664 19395
rect 32722 19395 33682 19442
rect 32722 19378 32924 19395
rect 32462 19361 32478 19378
rect 31890 19345 32478 19361
rect 32908 19361 32924 19378
rect 33480 19378 33682 19395
rect 33480 19361 33496 19378
rect 32908 19345 33496 19361
rect 13352 19211 13940 19227
rect 13352 19194 13368 19211
rect 13166 19177 13368 19194
rect 13924 19194 13940 19211
rect 14370 19211 14958 19227
rect 14370 19194 14386 19211
rect 13924 19177 14126 19194
rect 13166 19130 14126 19177
rect 14184 19177 14386 19194
rect 14942 19194 14958 19211
rect 15388 19211 15976 19227
rect 15388 19194 15404 19211
rect 14942 19177 15144 19194
rect 14184 19130 15144 19177
rect 15202 19177 15404 19194
rect 15960 19194 15976 19211
rect 16406 19211 16994 19227
rect 16406 19194 16422 19211
rect 15960 19177 16162 19194
rect 15202 19130 16162 19177
rect 16220 19177 16422 19194
rect 16978 19194 16994 19211
rect 16978 19177 17180 19194
rect 16220 19130 17180 19177
rect 18656 18867 19244 18883
rect 18656 18850 18672 18867
rect 18470 18833 18672 18850
rect 19228 18850 19244 18867
rect 19674 18867 20262 18883
rect 19674 18850 19690 18867
rect 19228 18833 19430 18850
rect 18470 18786 19430 18833
rect 19488 18833 19690 18850
rect 20246 18850 20262 18867
rect 20692 18867 21280 18883
rect 20692 18850 20708 18867
rect 20246 18833 20448 18850
rect 19488 18786 20448 18833
rect 20506 18833 20708 18850
rect 21264 18850 21280 18867
rect 21710 18867 22298 18883
rect 21710 18850 21726 18867
rect 21264 18833 21466 18850
rect 20506 18786 21466 18833
rect 21524 18833 21726 18850
rect 22282 18850 22298 18867
rect 22728 18867 23316 18883
rect 22728 18850 22744 18867
rect 22282 18833 22484 18850
rect 21524 18786 22484 18833
rect 22542 18833 22744 18850
rect 23300 18850 23316 18867
rect 23746 18867 24334 18883
rect 23746 18850 23762 18867
rect 23300 18833 23502 18850
rect 22542 18786 23502 18833
rect 23560 18833 23762 18850
rect 24318 18850 24334 18867
rect 24764 18867 25352 18883
rect 24764 18850 24780 18867
rect 24318 18833 24520 18850
rect 23560 18786 24520 18833
rect 24578 18833 24780 18850
rect 25336 18850 25352 18867
rect 25782 18867 26370 18883
rect 25782 18850 25798 18867
rect 25336 18833 25538 18850
rect 24578 18786 25538 18833
rect 25596 18833 25798 18850
rect 26354 18850 26370 18867
rect 26800 18867 27388 18883
rect 26800 18850 26816 18867
rect 26354 18833 26556 18850
rect 25596 18786 26556 18833
rect 26614 18833 26816 18850
rect 27372 18850 27388 18867
rect 27818 18867 28406 18883
rect 27818 18850 27834 18867
rect 27372 18833 27574 18850
rect 26614 18786 27574 18833
rect 27632 18833 27834 18850
rect 28390 18850 28406 18867
rect 28836 18867 29424 18883
rect 28836 18850 28852 18867
rect 28390 18833 28592 18850
rect 27632 18786 28592 18833
rect 28650 18833 28852 18850
rect 29408 18850 29424 18867
rect 29854 18867 30442 18883
rect 29854 18850 29870 18867
rect 29408 18833 29610 18850
rect 28650 18786 29610 18833
rect 29668 18833 29870 18850
rect 30426 18850 30442 18867
rect 30872 18867 31460 18883
rect 30872 18850 30888 18867
rect 30426 18833 30628 18850
rect 29668 18786 30628 18833
rect 30686 18833 30888 18850
rect 31444 18850 31460 18867
rect 31890 18867 32478 18883
rect 31890 18850 31906 18867
rect 31444 18833 31646 18850
rect 30686 18786 31646 18833
rect 31704 18833 31906 18850
rect 32462 18850 32478 18867
rect 32908 18867 33496 18883
rect 32908 18850 32924 18867
rect 32462 18833 32664 18850
rect 31704 18786 32664 18833
rect 32722 18833 32924 18850
rect 33480 18850 33496 18867
rect 33480 18833 33682 18850
rect 32722 18786 33682 18833
rect 13166 18483 14126 18530
rect 13166 18466 13368 18483
rect 13352 18449 13368 18466
rect 13924 18466 14126 18483
rect 14184 18483 15144 18530
rect 14184 18466 14386 18483
rect 13924 18449 13940 18466
rect 13352 18433 13940 18449
rect 14370 18449 14386 18466
rect 14942 18466 15144 18483
rect 15202 18483 16162 18530
rect 15202 18466 15404 18483
rect 14942 18449 14958 18466
rect 14370 18433 14958 18449
rect 15388 18449 15404 18466
rect 15960 18466 16162 18483
rect 16220 18483 17180 18530
rect 16220 18466 16422 18483
rect 15960 18449 15976 18466
rect 15388 18433 15976 18449
rect 16406 18449 16422 18466
rect 16978 18466 17180 18483
rect 16978 18449 16994 18466
rect 16406 18433 16994 18449
rect 13352 18179 13940 18195
rect 13352 18162 13368 18179
rect 13166 18145 13368 18162
rect 13924 18162 13940 18179
rect 14370 18179 14958 18195
rect 14370 18162 14386 18179
rect 13924 18145 14126 18162
rect 13166 18098 14126 18145
rect 14184 18145 14386 18162
rect 14942 18162 14958 18179
rect 15388 18179 15976 18195
rect 15388 18162 15404 18179
rect 14942 18145 15144 18162
rect 14184 18098 15144 18145
rect 15202 18145 15404 18162
rect 15960 18162 15976 18179
rect 16406 18179 16994 18195
rect 16406 18162 16422 18179
rect 15960 18145 16162 18162
rect 15202 18098 16162 18145
rect 16220 18145 16422 18162
rect 16978 18162 16994 18179
rect 16978 18145 17180 18162
rect 16220 18098 17180 18145
rect 18470 18139 19430 18186
rect 18470 18122 18672 18139
rect 18656 18105 18672 18122
rect 19228 18122 19430 18139
rect 19488 18139 20448 18186
rect 19488 18122 19690 18139
rect 19228 18105 19244 18122
rect 18656 18089 19244 18105
rect 19674 18105 19690 18122
rect 20246 18122 20448 18139
rect 20506 18139 21466 18186
rect 20506 18122 20708 18139
rect 20246 18105 20262 18122
rect 19674 18089 20262 18105
rect 20692 18105 20708 18122
rect 21264 18122 21466 18139
rect 21524 18139 22484 18186
rect 21524 18122 21726 18139
rect 21264 18105 21280 18122
rect 20692 18089 21280 18105
rect 21710 18105 21726 18122
rect 22282 18122 22484 18139
rect 22542 18139 23502 18186
rect 22542 18122 22744 18139
rect 22282 18105 22298 18122
rect 21710 18089 22298 18105
rect 22728 18105 22744 18122
rect 23300 18122 23502 18139
rect 23560 18139 24520 18186
rect 23560 18122 23762 18139
rect 23300 18105 23316 18122
rect 22728 18089 23316 18105
rect 23746 18105 23762 18122
rect 24318 18122 24520 18139
rect 24578 18139 25538 18186
rect 24578 18122 24780 18139
rect 24318 18105 24334 18122
rect 23746 18089 24334 18105
rect 24764 18105 24780 18122
rect 25336 18122 25538 18139
rect 25596 18139 26556 18186
rect 25596 18122 25798 18139
rect 25336 18105 25352 18122
rect 24764 18089 25352 18105
rect 25782 18105 25798 18122
rect 26354 18122 26556 18139
rect 26614 18139 27574 18186
rect 26614 18122 26816 18139
rect 26354 18105 26370 18122
rect 25782 18089 26370 18105
rect 26800 18105 26816 18122
rect 27372 18122 27574 18139
rect 27632 18139 28592 18186
rect 27632 18122 27834 18139
rect 27372 18105 27388 18122
rect 26800 18089 27388 18105
rect 27818 18105 27834 18122
rect 28390 18122 28592 18139
rect 28650 18139 29610 18186
rect 28650 18122 28852 18139
rect 28390 18105 28406 18122
rect 27818 18089 28406 18105
rect 28836 18105 28852 18122
rect 29408 18122 29610 18139
rect 29668 18139 30628 18186
rect 29668 18122 29870 18139
rect 29408 18105 29424 18122
rect 28836 18089 29424 18105
rect 29854 18105 29870 18122
rect 30426 18122 30628 18139
rect 30686 18139 31646 18186
rect 30686 18122 30888 18139
rect 30426 18105 30442 18122
rect 29854 18089 30442 18105
rect 30872 18105 30888 18122
rect 31444 18122 31646 18139
rect 31704 18139 32664 18186
rect 31704 18122 31906 18139
rect 31444 18105 31460 18122
rect 30872 18089 31460 18105
rect 31890 18105 31906 18122
rect 32462 18122 32664 18139
rect 32722 18139 33682 18186
rect 32722 18122 32924 18139
rect 32462 18105 32478 18122
rect 31890 18089 32478 18105
rect 32908 18105 32924 18122
rect 33480 18122 33682 18139
rect 33480 18105 33496 18122
rect 32908 18089 33496 18105
rect 18656 17611 19244 17627
rect 18656 17594 18672 17611
rect 18470 17577 18672 17594
rect 19228 17594 19244 17611
rect 19674 17611 20262 17627
rect 19674 17594 19690 17611
rect 19228 17577 19430 17594
rect 18470 17530 19430 17577
rect 19488 17577 19690 17594
rect 20246 17594 20262 17611
rect 20692 17611 21280 17627
rect 20692 17594 20708 17611
rect 20246 17577 20448 17594
rect 19488 17530 20448 17577
rect 20506 17577 20708 17594
rect 21264 17594 21280 17611
rect 21710 17611 22298 17627
rect 21710 17594 21726 17611
rect 21264 17577 21466 17594
rect 20506 17530 21466 17577
rect 21524 17577 21726 17594
rect 22282 17594 22298 17611
rect 22728 17611 23316 17627
rect 22728 17594 22744 17611
rect 22282 17577 22484 17594
rect 21524 17530 22484 17577
rect 22542 17577 22744 17594
rect 23300 17594 23316 17611
rect 23746 17611 24334 17627
rect 23746 17594 23762 17611
rect 23300 17577 23502 17594
rect 22542 17530 23502 17577
rect 23560 17577 23762 17594
rect 24318 17594 24334 17611
rect 24764 17611 25352 17627
rect 24764 17594 24780 17611
rect 24318 17577 24520 17594
rect 23560 17530 24520 17577
rect 24578 17577 24780 17594
rect 25336 17594 25352 17611
rect 25782 17611 26370 17627
rect 25782 17594 25798 17611
rect 25336 17577 25538 17594
rect 24578 17530 25538 17577
rect 25596 17577 25798 17594
rect 26354 17594 26370 17611
rect 26800 17611 27388 17627
rect 26800 17594 26816 17611
rect 26354 17577 26556 17594
rect 25596 17530 26556 17577
rect 26614 17577 26816 17594
rect 27372 17594 27388 17611
rect 27818 17611 28406 17627
rect 27818 17594 27834 17611
rect 27372 17577 27574 17594
rect 26614 17530 27574 17577
rect 27632 17577 27834 17594
rect 28390 17594 28406 17611
rect 28836 17611 29424 17627
rect 28836 17594 28852 17611
rect 28390 17577 28592 17594
rect 27632 17530 28592 17577
rect 28650 17577 28852 17594
rect 29408 17594 29424 17611
rect 29854 17611 30442 17627
rect 29854 17594 29870 17611
rect 29408 17577 29610 17594
rect 28650 17530 29610 17577
rect 29668 17577 29870 17594
rect 30426 17594 30442 17611
rect 30872 17611 31460 17627
rect 30872 17594 30888 17611
rect 30426 17577 30628 17594
rect 29668 17530 30628 17577
rect 30686 17577 30888 17594
rect 31444 17594 31460 17611
rect 31890 17611 32478 17627
rect 31890 17594 31906 17611
rect 31444 17577 31646 17594
rect 30686 17530 31646 17577
rect 31704 17577 31906 17594
rect 32462 17594 32478 17611
rect 32908 17611 33496 17627
rect 32908 17594 32924 17611
rect 32462 17577 32664 17594
rect 31704 17530 32664 17577
rect 32722 17577 32924 17594
rect 33480 17594 33496 17611
rect 33480 17577 33682 17594
rect 32722 17530 33682 17577
rect 13166 17451 14126 17498
rect 13166 17434 13368 17451
rect 13352 17417 13368 17434
rect 13924 17434 14126 17451
rect 14184 17451 15144 17498
rect 14184 17434 14386 17451
rect 13924 17417 13940 17434
rect 13352 17401 13940 17417
rect 14370 17417 14386 17434
rect 14942 17434 15144 17451
rect 15202 17451 16162 17498
rect 15202 17434 15404 17451
rect 14942 17417 14958 17434
rect 14370 17401 14958 17417
rect 15388 17417 15404 17434
rect 15960 17434 16162 17451
rect 16220 17451 17180 17498
rect 16220 17434 16422 17451
rect 15960 17417 15976 17434
rect 15388 17401 15976 17417
rect 16406 17417 16422 17434
rect 16978 17434 17180 17451
rect 16978 17417 16994 17434
rect 16406 17401 16994 17417
rect 18470 16883 19430 16930
rect 18470 16866 18672 16883
rect 18656 16849 18672 16866
rect 19228 16866 19430 16883
rect 19488 16883 20448 16930
rect 19488 16866 19690 16883
rect 19228 16849 19244 16866
rect 18656 16833 19244 16849
rect 19674 16849 19690 16866
rect 20246 16866 20448 16883
rect 20506 16883 21466 16930
rect 20506 16866 20708 16883
rect 20246 16849 20262 16866
rect 19674 16833 20262 16849
rect 20692 16849 20708 16866
rect 21264 16866 21466 16883
rect 21524 16883 22484 16930
rect 21524 16866 21726 16883
rect 21264 16849 21280 16866
rect 20692 16833 21280 16849
rect 21710 16849 21726 16866
rect 22282 16866 22484 16883
rect 22542 16883 23502 16930
rect 22542 16866 22744 16883
rect 22282 16849 22298 16866
rect 21710 16833 22298 16849
rect 22728 16849 22744 16866
rect 23300 16866 23502 16883
rect 23560 16883 24520 16930
rect 23560 16866 23762 16883
rect 23300 16849 23316 16866
rect 22728 16833 23316 16849
rect 23746 16849 23762 16866
rect 24318 16866 24520 16883
rect 24578 16883 25538 16930
rect 24578 16866 24780 16883
rect 24318 16849 24334 16866
rect 23746 16833 24334 16849
rect 24764 16849 24780 16866
rect 25336 16866 25538 16883
rect 25596 16883 26556 16930
rect 25596 16866 25798 16883
rect 25336 16849 25352 16866
rect 24764 16833 25352 16849
rect 25782 16849 25798 16866
rect 26354 16866 26556 16883
rect 26614 16883 27574 16930
rect 26614 16866 26816 16883
rect 26354 16849 26370 16866
rect 25782 16833 26370 16849
rect 26800 16849 26816 16866
rect 27372 16866 27574 16883
rect 27632 16883 28592 16930
rect 27632 16866 27834 16883
rect 27372 16849 27388 16866
rect 26800 16833 27388 16849
rect 27818 16849 27834 16866
rect 28390 16866 28592 16883
rect 28650 16883 29610 16930
rect 28650 16866 28852 16883
rect 28390 16849 28406 16866
rect 27818 16833 28406 16849
rect 28836 16849 28852 16866
rect 29408 16866 29610 16883
rect 29668 16883 30628 16930
rect 29668 16866 29870 16883
rect 29408 16849 29424 16866
rect 28836 16833 29424 16849
rect 29854 16849 29870 16866
rect 30426 16866 30628 16883
rect 30686 16883 31646 16930
rect 30686 16866 30888 16883
rect 30426 16849 30442 16866
rect 29854 16833 30442 16849
rect 30872 16849 30888 16866
rect 31444 16866 31646 16883
rect 31704 16883 32664 16930
rect 31704 16866 31906 16883
rect 31444 16849 31460 16866
rect 30872 16833 31460 16849
rect 31890 16849 31906 16866
rect 32462 16866 32664 16883
rect 32722 16883 33682 16930
rect 32722 16866 32924 16883
rect 32462 16849 32478 16866
rect 31890 16833 32478 16849
rect 32908 16849 32924 16866
rect 33480 16866 33682 16883
rect 33480 16849 33496 16866
rect 32908 16833 33496 16849
rect 58670 27925 59258 27941
rect 58670 27908 58686 27925
rect 58484 27891 58686 27908
rect 59242 27908 59258 27925
rect 59688 27925 60276 27941
rect 59688 27908 59704 27925
rect 59242 27891 59444 27908
rect 58484 27844 59444 27891
rect 59502 27891 59704 27908
rect 60260 27908 60276 27925
rect 60706 27925 61294 27941
rect 60706 27908 60722 27925
rect 60260 27891 60462 27908
rect 59502 27844 60462 27891
rect 60520 27891 60722 27908
rect 61278 27908 61294 27925
rect 61724 27925 62312 27941
rect 61724 27908 61740 27925
rect 61278 27891 61480 27908
rect 60520 27844 61480 27891
rect 61538 27891 61740 27908
rect 62296 27908 62312 27925
rect 62742 27925 63330 27941
rect 62742 27908 62758 27925
rect 62296 27891 62498 27908
rect 61538 27844 62498 27891
rect 62556 27891 62758 27908
rect 63314 27908 63330 27925
rect 63760 27925 64348 27941
rect 63760 27908 63776 27925
rect 63314 27891 63516 27908
rect 62556 27844 63516 27891
rect 63574 27891 63776 27908
rect 64332 27908 64348 27925
rect 64778 27925 65366 27941
rect 64778 27908 64794 27925
rect 64332 27891 64534 27908
rect 63574 27844 64534 27891
rect 64592 27891 64794 27908
rect 65350 27908 65366 27925
rect 65796 27925 66384 27941
rect 65796 27908 65812 27925
rect 65350 27891 65552 27908
rect 64592 27844 65552 27891
rect 65610 27891 65812 27908
rect 66368 27908 66384 27925
rect 66814 27925 67402 27941
rect 66814 27908 66830 27925
rect 66368 27891 66570 27908
rect 65610 27844 66570 27891
rect 66628 27891 66830 27908
rect 67386 27908 67402 27925
rect 67832 27925 68420 27941
rect 67832 27908 67848 27925
rect 67386 27891 67588 27908
rect 66628 27844 67588 27891
rect 67646 27891 67848 27908
rect 68404 27908 68420 27925
rect 68850 27925 69438 27941
rect 68850 27908 68866 27925
rect 68404 27891 68606 27908
rect 67646 27844 68606 27891
rect 68664 27891 68866 27908
rect 69422 27908 69438 27925
rect 69868 27925 70456 27941
rect 69868 27908 69884 27925
rect 69422 27891 69624 27908
rect 68664 27844 69624 27891
rect 69682 27891 69884 27908
rect 70440 27908 70456 27925
rect 70886 27925 71474 27941
rect 70886 27908 70902 27925
rect 70440 27891 70642 27908
rect 69682 27844 70642 27891
rect 70700 27891 70902 27908
rect 71458 27908 71474 27925
rect 71904 27925 72492 27941
rect 71904 27908 71920 27925
rect 71458 27891 71660 27908
rect 70700 27844 71660 27891
rect 71718 27891 71920 27908
rect 72476 27908 72492 27925
rect 72922 27925 73510 27941
rect 72922 27908 72938 27925
rect 72476 27891 72678 27908
rect 71718 27844 72678 27891
rect 72736 27891 72938 27908
rect 73494 27908 73510 27925
rect 73940 27925 74528 27941
rect 73940 27908 73956 27925
rect 73494 27891 73696 27908
rect 72736 27844 73696 27891
rect 73754 27891 73956 27908
rect 74512 27908 74528 27925
rect 74512 27891 74714 27908
rect 73754 27844 74714 27891
rect 58484 27197 59444 27244
rect 58484 27180 58686 27197
rect 58670 27163 58686 27180
rect 59242 27180 59444 27197
rect 59502 27197 60462 27244
rect 59502 27180 59704 27197
rect 59242 27163 59258 27180
rect 58670 27147 59258 27163
rect 59688 27163 59704 27180
rect 60260 27180 60462 27197
rect 60520 27197 61480 27244
rect 60520 27180 60722 27197
rect 60260 27163 60276 27180
rect 59688 27147 60276 27163
rect 60706 27163 60722 27180
rect 61278 27180 61480 27197
rect 61538 27197 62498 27244
rect 61538 27180 61740 27197
rect 61278 27163 61294 27180
rect 60706 27147 61294 27163
rect 61724 27163 61740 27180
rect 62296 27180 62498 27197
rect 62556 27197 63516 27244
rect 62556 27180 62758 27197
rect 62296 27163 62312 27180
rect 61724 27147 62312 27163
rect 62742 27163 62758 27180
rect 63314 27180 63516 27197
rect 63574 27197 64534 27244
rect 63574 27180 63776 27197
rect 63314 27163 63330 27180
rect 62742 27147 63330 27163
rect 63760 27163 63776 27180
rect 64332 27180 64534 27197
rect 64592 27197 65552 27244
rect 64592 27180 64794 27197
rect 64332 27163 64348 27180
rect 63760 27147 64348 27163
rect 64778 27163 64794 27180
rect 65350 27180 65552 27197
rect 65610 27197 66570 27244
rect 65610 27180 65812 27197
rect 65350 27163 65366 27180
rect 64778 27147 65366 27163
rect 65796 27163 65812 27180
rect 66368 27180 66570 27197
rect 66628 27197 67588 27244
rect 66628 27180 66830 27197
rect 66368 27163 66384 27180
rect 65796 27147 66384 27163
rect 66814 27163 66830 27180
rect 67386 27180 67588 27197
rect 67646 27197 68606 27244
rect 67646 27180 67848 27197
rect 67386 27163 67402 27180
rect 66814 27147 67402 27163
rect 67832 27163 67848 27180
rect 68404 27180 68606 27197
rect 68664 27197 69624 27244
rect 68664 27180 68866 27197
rect 68404 27163 68420 27180
rect 67832 27147 68420 27163
rect 68850 27163 68866 27180
rect 69422 27180 69624 27197
rect 69682 27197 70642 27244
rect 69682 27180 69884 27197
rect 69422 27163 69438 27180
rect 68850 27147 69438 27163
rect 69868 27163 69884 27180
rect 70440 27180 70642 27197
rect 70700 27197 71660 27244
rect 70700 27180 70902 27197
rect 70440 27163 70456 27180
rect 69868 27147 70456 27163
rect 70886 27163 70902 27180
rect 71458 27180 71660 27197
rect 71718 27197 72678 27244
rect 71718 27180 71920 27197
rect 71458 27163 71474 27180
rect 70886 27147 71474 27163
rect 71904 27163 71920 27180
rect 72476 27180 72678 27197
rect 72736 27197 73696 27244
rect 72736 27180 72938 27197
rect 72476 27163 72492 27180
rect 71904 27147 72492 27163
rect 72922 27163 72938 27180
rect 73494 27180 73696 27197
rect 73754 27197 74714 27244
rect 73754 27180 73956 27197
rect 73494 27163 73510 27180
rect 72922 27147 73510 27163
rect 73940 27163 73956 27180
rect 74512 27180 74714 27197
rect 74512 27163 74528 27180
rect 73940 27147 74528 27163
rect 58670 26789 59258 26805
rect 58670 26772 58686 26789
rect 58484 26755 58686 26772
rect 59242 26772 59258 26789
rect 59688 26789 60276 26805
rect 59688 26772 59704 26789
rect 59242 26755 59444 26772
rect 58484 26708 59444 26755
rect 59502 26755 59704 26772
rect 60260 26772 60276 26789
rect 60706 26789 61294 26805
rect 60706 26772 60722 26789
rect 60260 26755 60462 26772
rect 59502 26708 60462 26755
rect 60520 26755 60722 26772
rect 61278 26772 61294 26789
rect 61724 26789 62312 26805
rect 61724 26772 61740 26789
rect 61278 26755 61480 26772
rect 60520 26708 61480 26755
rect 61538 26755 61740 26772
rect 62296 26772 62312 26789
rect 62742 26789 63330 26805
rect 62742 26772 62758 26789
rect 62296 26755 62498 26772
rect 61538 26708 62498 26755
rect 62556 26755 62758 26772
rect 63314 26772 63330 26789
rect 63760 26789 64348 26805
rect 63760 26772 63776 26789
rect 63314 26755 63516 26772
rect 62556 26708 63516 26755
rect 63574 26755 63776 26772
rect 64332 26772 64348 26789
rect 64778 26789 65366 26805
rect 64778 26772 64794 26789
rect 64332 26755 64534 26772
rect 63574 26708 64534 26755
rect 64592 26755 64794 26772
rect 65350 26772 65366 26789
rect 65796 26789 66384 26805
rect 65796 26772 65812 26789
rect 65350 26755 65552 26772
rect 64592 26708 65552 26755
rect 65610 26755 65812 26772
rect 66368 26772 66384 26789
rect 66814 26789 67402 26805
rect 66814 26772 66830 26789
rect 66368 26755 66570 26772
rect 65610 26708 66570 26755
rect 66628 26755 66830 26772
rect 67386 26772 67402 26789
rect 67832 26789 68420 26805
rect 67832 26772 67848 26789
rect 67386 26755 67588 26772
rect 66628 26708 67588 26755
rect 67646 26755 67848 26772
rect 68404 26772 68420 26789
rect 68850 26789 69438 26805
rect 68850 26772 68866 26789
rect 68404 26755 68606 26772
rect 67646 26708 68606 26755
rect 68664 26755 68866 26772
rect 69422 26772 69438 26789
rect 69868 26789 70456 26805
rect 69868 26772 69884 26789
rect 69422 26755 69624 26772
rect 68664 26708 69624 26755
rect 69682 26755 69884 26772
rect 70440 26772 70456 26789
rect 70886 26789 71474 26805
rect 70886 26772 70902 26789
rect 70440 26755 70642 26772
rect 69682 26708 70642 26755
rect 70700 26755 70902 26772
rect 71458 26772 71474 26789
rect 71904 26789 72492 26805
rect 71904 26772 71920 26789
rect 71458 26755 71660 26772
rect 70700 26708 71660 26755
rect 71718 26755 71920 26772
rect 72476 26772 72492 26789
rect 72922 26789 73510 26805
rect 72922 26772 72938 26789
rect 72476 26755 72678 26772
rect 71718 26708 72678 26755
rect 72736 26755 72938 26772
rect 73494 26772 73510 26789
rect 73940 26789 74528 26805
rect 73940 26772 73956 26789
rect 73494 26755 73696 26772
rect 72736 26708 73696 26755
rect 73754 26755 73956 26772
rect 74512 26772 74528 26789
rect 74512 26755 74714 26772
rect 73754 26708 74714 26755
rect 58484 26061 59444 26108
rect 58484 26044 58686 26061
rect 58670 26027 58686 26044
rect 59242 26044 59444 26061
rect 59502 26061 60462 26108
rect 59502 26044 59704 26061
rect 59242 26027 59258 26044
rect 58670 26011 59258 26027
rect 59688 26027 59704 26044
rect 60260 26044 60462 26061
rect 60520 26061 61480 26108
rect 60520 26044 60722 26061
rect 60260 26027 60276 26044
rect 59688 26011 60276 26027
rect 60706 26027 60722 26044
rect 61278 26044 61480 26061
rect 61538 26061 62498 26108
rect 61538 26044 61740 26061
rect 61278 26027 61294 26044
rect 60706 26011 61294 26027
rect 61724 26027 61740 26044
rect 62296 26044 62498 26061
rect 62556 26061 63516 26108
rect 62556 26044 62758 26061
rect 62296 26027 62312 26044
rect 61724 26011 62312 26027
rect 62742 26027 62758 26044
rect 63314 26044 63516 26061
rect 63574 26061 64534 26108
rect 63574 26044 63776 26061
rect 63314 26027 63330 26044
rect 62742 26011 63330 26027
rect 63760 26027 63776 26044
rect 64332 26044 64534 26061
rect 64592 26061 65552 26108
rect 64592 26044 64794 26061
rect 64332 26027 64348 26044
rect 63760 26011 64348 26027
rect 64778 26027 64794 26044
rect 65350 26044 65552 26061
rect 65610 26061 66570 26108
rect 65610 26044 65812 26061
rect 65350 26027 65366 26044
rect 64778 26011 65366 26027
rect 65796 26027 65812 26044
rect 66368 26044 66570 26061
rect 66628 26061 67588 26108
rect 66628 26044 66830 26061
rect 66368 26027 66384 26044
rect 65796 26011 66384 26027
rect 66814 26027 66830 26044
rect 67386 26044 67588 26061
rect 67646 26061 68606 26108
rect 67646 26044 67848 26061
rect 67386 26027 67402 26044
rect 66814 26011 67402 26027
rect 67832 26027 67848 26044
rect 68404 26044 68606 26061
rect 68664 26061 69624 26108
rect 68664 26044 68866 26061
rect 68404 26027 68420 26044
rect 67832 26011 68420 26027
rect 68850 26027 68866 26044
rect 69422 26044 69624 26061
rect 69682 26061 70642 26108
rect 69682 26044 69884 26061
rect 69422 26027 69438 26044
rect 68850 26011 69438 26027
rect 69868 26027 69884 26044
rect 70440 26044 70642 26061
rect 70700 26061 71660 26108
rect 70700 26044 70902 26061
rect 70440 26027 70456 26044
rect 69868 26011 70456 26027
rect 70886 26027 70902 26044
rect 71458 26044 71660 26061
rect 71718 26061 72678 26108
rect 71718 26044 71920 26061
rect 71458 26027 71474 26044
rect 70886 26011 71474 26027
rect 71904 26027 71920 26044
rect 72476 26044 72678 26061
rect 72736 26061 73696 26108
rect 72736 26044 72938 26061
rect 72476 26027 72492 26044
rect 71904 26011 72492 26027
rect 72922 26027 72938 26044
rect 73494 26044 73696 26061
rect 73754 26061 74714 26108
rect 73754 26044 73956 26061
rect 73494 26027 73510 26044
rect 72922 26011 73510 26027
rect 73940 26027 73956 26044
rect 74512 26044 74714 26061
rect 74512 26027 74528 26044
rect 73940 26011 74528 26027
rect 58670 25653 59258 25669
rect 58670 25636 58686 25653
rect 58484 25619 58686 25636
rect 59242 25636 59258 25653
rect 59688 25653 60276 25669
rect 59688 25636 59704 25653
rect 59242 25619 59444 25636
rect 58484 25572 59444 25619
rect 59502 25619 59704 25636
rect 60260 25636 60276 25653
rect 60706 25653 61294 25669
rect 60706 25636 60722 25653
rect 60260 25619 60462 25636
rect 59502 25572 60462 25619
rect 60520 25619 60722 25636
rect 61278 25636 61294 25653
rect 61724 25653 62312 25669
rect 61724 25636 61740 25653
rect 61278 25619 61480 25636
rect 60520 25572 61480 25619
rect 61538 25619 61740 25636
rect 62296 25636 62312 25653
rect 62742 25653 63330 25669
rect 62742 25636 62758 25653
rect 62296 25619 62498 25636
rect 61538 25572 62498 25619
rect 62556 25619 62758 25636
rect 63314 25636 63330 25653
rect 63760 25653 64348 25669
rect 63760 25636 63776 25653
rect 63314 25619 63516 25636
rect 62556 25572 63516 25619
rect 63574 25619 63776 25636
rect 64332 25636 64348 25653
rect 64778 25653 65366 25669
rect 64778 25636 64794 25653
rect 64332 25619 64534 25636
rect 63574 25572 64534 25619
rect 64592 25619 64794 25636
rect 65350 25636 65366 25653
rect 65796 25653 66384 25669
rect 65796 25636 65812 25653
rect 65350 25619 65552 25636
rect 64592 25572 65552 25619
rect 65610 25619 65812 25636
rect 66368 25636 66384 25653
rect 66814 25653 67402 25669
rect 66814 25636 66830 25653
rect 66368 25619 66570 25636
rect 65610 25572 66570 25619
rect 66628 25619 66830 25636
rect 67386 25636 67402 25653
rect 67832 25653 68420 25669
rect 67832 25636 67848 25653
rect 67386 25619 67588 25636
rect 66628 25572 67588 25619
rect 67646 25619 67848 25636
rect 68404 25636 68420 25653
rect 68850 25653 69438 25669
rect 68850 25636 68866 25653
rect 68404 25619 68606 25636
rect 67646 25572 68606 25619
rect 68664 25619 68866 25636
rect 69422 25636 69438 25653
rect 69868 25653 70456 25669
rect 69868 25636 69884 25653
rect 69422 25619 69624 25636
rect 68664 25572 69624 25619
rect 69682 25619 69884 25636
rect 70440 25636 70456 25653
rect 70886 25653 71474 25669
rect 70886 25636 70902 25653
rect 70440 25619 70642 25636
rect 69682 25572 70642 25619
rect 70700 25619 70902 25636
rect 71458 25636 71474 25653
rect 71904 25653 72492 25669
rect 71904 25636 71920 25653
rect 71458 25619 71660 25636
rect 70700 25572 71660 25619
rect 71718 25619 71920 25636
rect 72476 25636 72492 25653
rect 72922 25653 73510 25669
rect 72922 25636 72938 25653
rect 72476 25619 72678 25636
rect 71718 25572 72678 25619
rect 72736 25619 72938 25636
rect 73494 25636 73510 25653
rect 73940 25653 74528 25669
rect 73940 25636 73956 25653
rect 73494 25619 73696 25636
rect 72736 25572 73696 25619
rect 73754 25619 73956 25636
rect 74512 25636 74528 25653
rect 74512 25619 74714 25636
rect 73754 25572 74714 25619
rect 58484 24925 59444 24972
rect 58484 24908 58686 24925
rect 58670 24891 58686 24908
rect 59242 24908 59444 24925
rect 59502 24925 60462 24972
rect 59502 24908 59704 24925
rect 59242 24891 59258 24908
rect 58670 24875 59258 24891
rect 59688 24891 59704 24908
rect 60260 24908 60462 24925
rect 60520 24925 61480 24972
rect 60520 24908 60722 24925
rect 60260 24891 60276 24908
rect 59688 24875 60276 24891
rect 60706 24891 60722 24908
rect 61278 24908 61480 24925
rect 61538 24925 62498 24972
rect 61538 24908 61740 24925
rect 61278 24891 61294 24908
rect 60706 24875 61294 24891
rect 61724 24891 61740 24908
rect 62296 24908 62498 24925
rect 62556 24925 63516 24972
rect 62556 24908 62758 24925
rect 62296 24891 62312 24908
rect 61724 24875 62312 24891
rect 62742 24891 62758 24908
rect 63314 24908 63516 24925
rect 63574 24925 64534 24972
rect 63574 24908 63776 24925
rect 63314 24891 63330 24908
rect 62742 24875 63330 24891
rect 63760 24891 63776 24908
rect 64332 24908 64534 24925
rect 64592 24925 65552 24972
rect 64592 24908 64794 24925
rect 64332 24891 64348 24908
rect 63760 24875 64348 24891
rect 64778 24891 64794 24908
rect 65350 24908 65552 24925
rect 65610 24925 66570 24972
rect 65610 24908 65812 24925
rect 65350 24891 65366 24908
rect 64778 24875 65366 24891
rect 65796 24891 65812 24908
rect 66368 24908 66570 24925
rect 66628 24925 67588 24972
rect 66628 24908 66830 24925
rect 66368 24891 66384 24908
rect 65796 24875 66384 24891
rect 66814 24891 66830 24908
rect 67386 24908 67588 24925
rect 67646 24925 68606 24972
rect 67646 24908 67848 24925
rect 67386 24891 67402 24908
rect 66814 24875 67402 24891
rect 67832 24891 67848 24908
rect 68404 24908 68606 24925
rect 68664 24925 69624 24972
rect 68664 24908 68866 24925
rect 68404 24891 68420 24908
rect 67832 24875 68420 24891
rect 68850 24891 68866 24908
rect 69422 24908 69624 24925
rect 69682 24925 70642 24972
rect 69682 24908 69884 24925
rect 69422 24891 69438 24908
rect 68850 24875 69438 24891
rect 69868 24891 69884 24908
rect 70440 24908 70642 24925
rect 70700 24925 71660 24972
rect 70700 24908 70902 24925
rect 70440 24891 70456 24908
rect 69868 24875 70456 24891
rect 70886 24891 70902 24908
rect 71458 24908 71660 24925
rect 71718 24925 72678 24972
rect 71718 24908 71920 24925
rect 71458 24891 71474 24908
rect 70886 24875 71474 24891
rect 71904 24891 71920 24908
rect 72476 24908 72678 24925
rect 72736 24925 73696 24972
rect 72736 24908 72938 24925
rect 72476 24891 72492 24908
rect 71904 24875 72492 24891
rect 72922 24891 72938 24908
rect 73494 24908 73696 24925
rect 73754 24925 74714 24972
rect 73754 24908 73956 24925
rect 73494 24891 73510 24908
rect 72922 24875 73510 24891
rect 73940 24891 73956 24908
rect 74512 24908 74714 24925
rect 74512 24891 74528 24908
rect 73940 24875 74528 24891
rect 59864 24015 60452 24031
rect 59864 23998 59880 24015
rect 59678 23981 59880 23998
rect 60436 23998 60452 24015
rect 60882 24015 61470 24031
rect 60882 23998 60898 24015
rect 60436 23981 60638 23998
rect 59678 23934 60638 23981
rect 60696 23981 60898 23998
rect 61454 23998 61470 24015
rect 61900 24015 62488 24031
rect 61900 23998 61916 24015
rect 61454 23981 61656 23998
rect 60696 23934 61656 23981
rect 61714 23981 61916 23998
rect 62472 23998 62488 24015
rect 62918 24015 63506 24031
rect 62918 23998 62934 24015
rect 62472 23981 62674 23998
rect 61714 23934 62674 23981
rect 62732 23981 62934 23998
rect 63490 23998 63506 24015
rect 63936 24015 64524 24031
rect 63936 23998 63952 24015
rect 63490 23981 63692 23998
rect 62732 23934 63692 23981
rect 63750 23981 63952 23998
rect 64508 23998 64524 24015
rect 64954 24015 65542 24031
rect 64954 23998 64970 24015
rect 64508 23981 64710 23998
rect 63750 23934 64710 23981
rect 64768 23981 64970 23998
rect 65526 23998 65542 24015
rect 65972 24015 66560 24031
rect 65972 23998 65988 24015
rect 65526 23981 65728 23998
rect 64768 23934 65728 23981
rect 65786 23981 65988 23998
rect 66544 23998 66560 24015
rect 66990 24015 67578 24031
rect 66990 23998 67006 24015
rect 66544 23981 66746 23998
rect 65786 23934 66746 23981
rect 66804 23981 67006 23998
rect 67562 23998 67578 24015
rect 68008 24015 68596 24031
rect 68008 23998 68024 24015
rect 67562 23981 67764 23998
rect 66804 23934 67764 23981
rect 67822 23981 68024 23998
rect 68580 23998 68596 24015
rect 69026 24015 69614 24031
rect 69026 23998 69042 24015
rect 68580 23981 68782 23998
rect 67822 23934 68782 23981
rect 68840 23981 69042 23998
rect 69598 23998 69614 24015
rect 70044 24015 70632 24031
rect 70044 23998 70060 24015
rect 69598 23981 69800 23998
rect 68840 23934 69800 23981
rect 69858 23981 70060 23998
rect 70616 23998 70632 24015
rect 71062 24015 71650 24031
rect 71062 23998 71078 24015
rect 70616 23981 70818 23998
rect 69858 23934 70818 23981
rect 70876 23981 71078 23998
rect 71634 23998 71650 24015
rect 72080 24015 72668 24031
rect 72080 23998 72096 24015
rect 71634 23981 71836 23998
rect 70876 23934 71836 23981
rect 71894 23981 72096 23998
rect 72652 23998 72668 24015
rect 73098 24015 73686 24031
rect 73098 23998 73114 24015
rect 72652 23981 72854 23998
rect 71894 23934 72854 23981
rect 72912 23981 73114 23998
rect 73670 23998 73686 24015
rect 73670 23981 73872 23998
rect 72912 23934 73872 23981
rect 59678 23287 60638 23334
rect 59678 23270 59880 23287
rect 59864 23253 59880 23270
rect 60436 23270 60638 23287
rect 60696 23287 61656 23334
rect 60696 23270 60898 23287
rect 60436 23253 60452 23270
rect 59864 23237 60452 23253
rect 60882 23253 60898 23270
rect 61454 23270 61656 23287
rect 61714 23287 62674 23334
rect 61714 23270 61916 23287
rect 61454 23253 61470 23270
rect 60882 23237 61470 23253
rect 61900 23253 61916 23270
rect 62472 23270 62674 23287
rect 62732 23287 63692 23334
rect 62732 23270 62934 23287
rect 62472 23253 62488 23270
rect 61900 23237 62488 23253
rect 62918 23253 62934 23270
rect 63490 23270 63692 23287
rect 63750 23287 64710 23334
rect 63750 23270 63952 23287
rect 63490 23253 63506 23270
rect 62918 23237 63506 23253
rect 63936 23253 63952 23270
rect 64508 23270 64710 23287
rect 64768 23287 65728 23334
rect 64768 23270 64970 23287
rect 64508 23253 64524 23270
rect 63936 23237 64524 23253
rect 64954 23253 64970 23270
rect 65526 23270 65728 23287
rect 65786 23287 66746 23334
rect 65786 23270 65988 23287
rect 65526 23253 65542 23270
rect 64954 23237 65542 23253
rect 65972 23253 65988 23270
rect 66544 23270 66746 23287
rect 66804 23287 67764 23334
rect 66804 23270 67006 23287
rect 66544 23253 66560 23270
rect 65972 23237 66560 23253
rect 66990 23253 67006 23270
rect 67562 23270 67764 23287
rect 67822 23287 68782 23334
rect 67822 23270 68024 23287
rect 67562 23253 67578 23270
rect 66990 23237 67578 23253
rect 68008 23253 68024 23270
rect 68580 23270 68782 23287
rect 68840 23287 69800 23334
rect 68840 23270 69042 23287
rect 68580 23253 68596 23270
rect 68008 23237 68596 23253
rect 69026 23253 69042 23270
rect 69598 23270 69800 23287
rect 69858 23287 70818 23334
rect 69858 23270 70060 23287
rect 69598 23253 69614 23270
rect 69026 23237 69614 23253
rect 70044 23253 70060 23270
rect 70616 23270 70818 23287
rect 70876 23287 71836 23334
rect 70876 23270 71078 23287
rect 70616 23253 70632 23270
rect 70044 23237 70632 23253
rect 71062 23253 71078 23270
rect 71634 23270 71836 23287
rect 71894 23287 72854 23334
rect 71894 23270 72096 23287
rect 71634 23253 71650 23270
rect 71062 23237 71650 23253
rect 72080 23253 72096 23270
rect 72652 23270 72854 23287
rect 72912 23287 73872 23334
rect 72912 23270 73114 23287
rect 72652 23253 72668 23270
rect 72080 23237 72668 23253
rect 73098 23253 73114 23270
rect 73670 23270 73872 23287
rect 73670 23253 73686 23270
rect 73098 23237 73686 23253
rect 59864 22983 60452 22999
rect 59864 22966 59880 22983
rect 59678 22949 59880 22966
rect 60436 22966 60452 22983
rect 60882 22983 61470 22999
rect 60882 22966 60898 22983
rect 60436 22949 60638 22966
rect 59678 22902 60638 22949
rect 60696 22949 60898 22966
rect 61454 22966 61470 22983
rect 61900 22983 62488 22999
rect 61900 22966 61916 22983
rect 61454 22949 61656 22966
rect 60696 22902 61656 22949
rect 61714 22949 61916 22966
rect 62472 22966 62488 22983
rect 62918 22983 63506 22999
rect 62918 22966 62934 22983
rect 62472 22949 62674 22966
rect 61714 22902 62674 22949
rect 62732 22949 62934 22966
rect 63490 22966 63506 22983
rect 63936 22983 64524 22999
rect 63936 22966 63952 22983
rect 63490 22949 63692 22966
rect 62732 22902 63692 22949
rect 63750 22949 63952 22966
rect 64508 22966 64524 22983
rect 64954 22983 65542 22999
rect 64954 22966 64970 22983
rect 64508 22949 64710 22966
rect 63750 22902 64710 22949
rect 64768 22949 64970 22966
rect 65526 22966 65542 22983
rect 65972 22983 66560 22999
rect 65972 22966 65988 22983
rect 65526 22949 65728 22966
rect 64768 22902 65728 22949
rect 65786 22949 65988 22966
rect 66544 22966 66560 22983
rect 66990 22983 67578 22999
rect 66990 22966 67006 22983
rect 66544 22949 66746 22966
rect 65786 22902 66746 22949
rect 66804 22949 67006 22966
rect 67562 22966 67578 22983
rect 68008 22983 68596 22999
rect 68008 22966 68024 22983
rect 67562 22949 67764 22966
rect 66804 22902 67764 22949
rect 67822 22949 68024 22966
rect 68580 22966 68596 22983
rect 69026 22983 69614 22999
rect 69026 22966 69042 22983
rect 68580 22949 68782 22966
rect 67822 22902 68782 22949
rect 68840 22949 69042 22966
rect 69598 22966 69614 22983
rect 70044 22983 70632 22999
rect 70044 22966 70060 22983
rect 69598 22949 69800 22966
rect 68840 22902 69800 22949
rect 69858 22949 70060 22966
rect 70616 22966 70632 22983
rect 71062 22983 71650 22999
rect 71062 22966 71078 22983
rect 70616 22949 70818 22966
rect 69858 22902 70818 22949
rect 70876 22949 71078 22966
rect 71634 22966 71650 22983
rect 72080 22983 72668 22999
rect 72080 22966 72096 22983
rect 71634 22949 71836 22966
rect 70876 22902 71836 22949
rect 71894 22949 72096 22966
rect 72652 22966 72668 22983
rect 73098 22983 73686 22999
rect 73098 22966 73114 22983
rect 72652 22949 72854 22966
rect 71894 22902 72854 22949
rect 72912 22949 73114 22966
rect 73670 22966 73686 22983
rect 73670 22949 73872 22966
rect 72912 22902 73872 22949
rect 59678 22255 60638 22302
rect 59678 22238 59880 22255
rect 59864 22221 59880 22238
rect 60436 22238 60638 22255
rect 60696 22255 61656 22302
rect 60696 22238 60898 22255
rect 60436 22221 60452 22238
rect 59864 22205 60452 22221
rect 60882 22221 60898 22238
rect 61454 22238 61656 22255
rect 61714 22255 62674 22302
rect 61714 22238 61916 22255
rect 61454 22221 61470 22238
rect 60882 22205 61470 22221
rect 61900 22221 61916 22238
rect 62472 22238 62674 22255
rect 62732 22255 63692 22302
rect 62732 22238 62934 22255
rect 62472 22221 62488 22238
rect 61900 22205 62488 22221
rect 62918 22221 62934 22238
rect 63490 22238 63692 22255
rect 63750 22255 64710 22302
rect 63750 22238 63952 22255
rect 63490 22221 63506 22238
rect 62918 22205 63506 22221
rect 63936 22221 63952 22238
rect 64508 22238 64710 22255
rect 64768 22255 65728 22302
rect 64768 22238 64970 22255
rect 64508 22221 64524 22238
rect 63936 22205 64524 22221
rect 64954 22221 64970 22238
rect 65526 22238 65728 22255
rect 65786 22255 66746 22302
rect 65786 22238 65988 22255
rect 65526 22221 65542 22238
rect 64954 22205 65542 22221
rect 65972 22221 65988 22238
rect 66544 22238 66746 22255
rect 66804 22255 67764 22302
rect 66804 22238 67006 22255
rect 66544 22221 66560 22238
rect 65972 22205 66560 22221
rect 66990 22221 67006 22238
rect 67562 22238 67764 22255
rect 67822 22255 68782 22302
rect 67822 22238 68024 22255
rect 67562 22221 67578 22238
rect 66990 22205 67578 22221
rect 68008 22221 68024 22238
rect 68580 22238 68782 22255
rect 68840 22255 69800 22302
rect 68840 22238 69042 22255
rect 68580 22221 68596 22238
rect 68008 22205 68596 22221
rect 69026 22221 69042 22238
rect 69598 22238 69800 22255
rect 69858 22255 70818 22302
rect 69858 22238 70060 22255
rect 69598 22221 69614 22238
rect 69026 22205 69614 22221
rect 70044 22221 70060 22238
rect 70616 22238 70818 22255
rect 70876 22255 71836 22302
rect 70876 22238 71078 22255
rect 70616 22221 70632 22238
rect 70044 22205 70632 22221
rect 71062 22221 71078 22238
rect 71634 22238 71836 22255
rect 71894 22255 72854 22302
rect 71894 22238 72096 22255
rect 71634 22221 71650 22238
rect 71062 22205 71650 22221
rect 72080 22221 72096 22238
rect 72652 22238 72854 22255
rect 72912 22255 73872 22302
rect 72912 22238 73114 22255
rect 72652 22221 72668 22238
rect 72080 22205 72668 22221
rect 73098 22221 73114 22238
rect 73670 22238 73872 22255
rect 73670 22221 73686 22238
rect 73098 22205 73686 22221
rect 59656 21379 60244 21395
rect 59656 21362 59672 21379
rect 59470 21345 59672 21362
rect 60228 21362 60244 21379
rect 60674 21379 61262 21395
rect 60674 21362 60690 21379
rect 60228 21345 60430 21362
rect 59470 21298 60430 21345
rect 60488 21345 60690 21362
rect 61246 21362 61262 21379
rect 61692 21379 62280 21395
rect 61692 21362 61708 21379
rect 61246 21345 61448 21362
rect 60488 21298 61448 21345
rect 61506 21345 61708 21362
rect 62264 21362 62280 21379
rect 62710 21379 63298 21395
rect 62710 21362 62726 21379
rect 62264 21345 62466 21362
rect 61506 21298 62466 21345
rect 62524 21345 62726 21362
rect 63282 21362 63298 21379
rect 63728 21379 64316 21395
rect 63728 21362 63744 21379
rect 63282 21345 63484 21362
rect 62524 21298 63484 21345
rect 63542 21345 63744 21362
rect 64300 21362 64316 21379
rect 64746 21379 65334 21395
rect 64746 21362 64762 21379
rect 64300 21345 64502 21362
rect 63542 21298 64502 21345
rect 64560 21345 64762 21362
rect 65318 21362 65334 21379
rect 65764 21379 66352 21395
rect 65764 21362 65780 21379
rect 65318 21345 65520 21362
rect 64560 21298 65520 21345
rect 65578 21345 65780 21362
rect 66336 21362 66352 21379
rect 66782 21379 67370 21395
rect 66782 21362 66798 21379
rect 66336 21345 66538 21362
rect 65578 21298 66538 21345
rect 66596 21345 66798 21362
rect 67354 21362 67370 21379
rect 67800 21379 68388 21395
rect 67800 21362 67816 21379
rect 67354 21345 67556 21362
rect 66596 21298 67556 21345
rect 67614 21345 67816 21362
rect 68372 21362 68388 21379
rect 68818 21379 69406 21395
rect 68818 21362 68834 21379
rect 68372 21345 68574 21362
rect 67614 21298 68574 21345
rect 68632 21345 68834 21362
rect 69390 21362 69406 21379
rect 69836 21379 70424 21395
rect 69836 21362 69852 21379
rect 69390 21345 69592 21362
rect 68632 21298 69592 21345
rect 69650 21345 69852 21362
rect 70408 21362 70424 21379
rect 70854 21379 71442 21395
rect 70854 21362 70870 21379
rect 70408 21345 70610 21362
rect 69650 21298 70610 21345
rect 70668 21345 70870 21362
rect 71426 21362 71442 21379
rect 71872 21379 72460 21395
rect 71872 21362 71888 21379
rect 71426 21345 71628 21362
rect 70668 21298 71628 21345
rect 71686 21345 71888 21362
rect 72444 21362 72460 21379
rect 72890 21379 73478 21395
rect 72890 21362 72906 21379
rect 72444 21345 72646 21362
rect 71686 21298 72646 21345
rect 72704 21345 72906 21362
rect 73462 21362 73478 21379
rect 73908 21379 74496 21395
rect 73908 21362 73924 21379
rect 73462 21345 73664 21362
rect 72704 21298 73664 21345
rect 73722 21345 73924 21362
rect 74480 21362 74496 21379
rect 74480 21345 74682 21362
rect 73722 21298 74682 21345
rect 54352 21275 54940 21291
rect 54352 21258 54368 21275
rect 54166 21241 54368 21258
rect 54924 21258 54940 21275
rect 55370 21275 55958 21291
rect 55370 21258 55386 21275
rect 54924 21241 55126 21258
rect 54166 21194 55126 21241
rect 55184 21241 55386 21258
rect 55942 21258 55958 21275
rect 56388 21275 56976 21291
rect 56388 21258 56404 21275
rect 55942 21241 56144 21258
rect 55184 21194 56144 21241
rect 56202 21241 56404 21258
rect 56960 21258 56976 21275
rect 57406 21275 57994 21291
rect 57406 21258 57422 21275
rect 56960 21241 57162 21258
rect 56202 21194 57162 21241
rect 57220 21241 57422 21258
rect 57978 21258 57994 21275
rect 57978 21241 58180 21258
rect 57220 21194 58180 21241
rect 59470 20651 60430 20698
rect 59470 20634 59672 20651
rect 59656 20617 59672 20634
rect 60228 20634 60430 20651
rect 60488 20651 61448 20698
rect 60488 20634 60690 20651
rect 60228 20617 60244 20634
rect 59656 20601 60244 20617
rect 60674 20617 60690 20634
rect 61246 20634 61448 20651
rect 61506 20651 62466 20698
rect 61506 20634 61708 20651
rect 61246 20617 61262 20634
rect 60674 20601 61262 20617
rect 61692 20617 61708 20634
rect 62264 20634 62466 20651
rect 62524 20651 63484 20698
rect 62524 20634 62726 20651
rect 62264 20617 62280 20634
rect 61692 20601 62280 20617
rect 62710 20617 62726 20634
rect 63282 20634 63484 20651
rect 63542 20651 64502 20698
rect 63542 20634 63744 20651
rect 63282 20617 63298 20634
rect 62710 20601 63298 20617
rect 63728 20617 63744 20634
rect 64300 20634 64502 20651
rect 64560 20651 65520 20698
rect 64560 20634 64762 20651
rect 64300 20617 64316 20634
rect 63728 20601 64316 20617
rect 64746 20617 64762 20634
rect 65318 20634 65520 20651
rect 65578 20651 66538 20698
rect 65578 20634 65780 20651
rect 65318 20617 65334 20634
rect 64746 20601 65334 20617
rect 65764 20617 65780 20634
rect 66336 20634 66538 20651
rect 66596 20651 67556 20698
rect 66596 20634 66798 20651
rect 66336 20617 66352 20634
rect 65764 20601 66352 20617
rect 66782 20617 66798 20634
rect 67354 20634 67556 20651
rect 67614 20651 68574 20698
rect 67614 20634 67816 20651
rect 67354 20617 67370 20634
rect 66782 20601 67370 20617
rect 67800 20617 67816 20634
rect 68372 20634 68574 20651
rect 68632 20651 69592 20698
rect 68632 20634 68834 20651
rect 68372 20617 68388 20634
rect 67800 20601 68388 20617
rect 68818 20617 68834 20634
rect 69390 20634 69592 20651
rect 69650 20651 70610 20698
rect 69650 20634 69852 20651
rect 69390 20617 69406 20634
rect 68818 20601 69406 20617
rect 69836 20617 69852 20634
rect 70408 20634 70610 20651
rect 70668 20651 71628 20698
rect 70668 20634 70870 20651
rect 70408 20617 70424 20634
rect 69836 20601 70424 20617
rect 70854 20617 70870 20634
rect 71426 20634 71628 20651
rect 71686 20651 72646 20698
rect 71686 20634 71888 20651
rect 71426 20617 71442 20634
rect 70854 20601 71442 20617
rect 71872 20617 71888 20634
rect 72444 20634 72646 20651
rect 72704 20651 73664 20698
rect 72704 20634 72906 20651
rect 72444 20617 72460 20634
rect 71872 20601 72460 20617
rect 72890 20617 72906 20634
rect 73462 20634 73664 20651
rect 73722 20651 74682 20698
rect 73722 20634 73924 20651
rect 73462 20617 73478 20634
rect 72890 20601 73478 20617
rect 73908 20617 73924 20634
rect 74480 20634 74682 20651
rect 74480 20617 74496 20634
rect 73908 20601 74496 20617
rect 54166 20547 55126 20594
rect 54166 20530 54368 20547
rect 54352 20513 54368 20530
rect 54924 20530 55126 20547
rect 55184 20547 56144 20594
rect 55184 20530 55386 20547
rect 54924 20513 54940 20530
rect 54352 20497 54940 20513
rect 55370 20513 55386 20530
rect 55942 20530 56144 20547
rect 56202 20547 57162 20594
rect 56202 20530 56404 20547
rect 55942 20513 55958 20530
rect 55370 20497 55958 20513
rect 56388 20513 56404 20530
rect 56960 20530 57162 20547
rect 57220 20547 58180 20594
rect 57220 20530 57422 20547
rect 56960 20513 56976 20530
rect 56388 20497 56976 20513
rect 57406 20513 57422 20530
rect 57978 20530 58180 20547
rect 57978 20513 57994 20530
rect 57406 20497 57994 20513
rect 54352 20243 54940 20259
rect 54352 20226 54368 20243
rect 54166 20209 54368 20226
rect 54924 20226 54940 20243
rect 55370 20243 55958 20259
rect 55370 20226 55386 20243
rect 54924 20209 55126 20226
rect 54166 20162 55126 20209
rect 55184 20209 55386 20226
rect 55942 20226 55958 20243
rect 56388 20243 56976 20259
rect 56388 20226 56404 20243
rect 55942 20209 56144 20226
rect 55184 20162 56144 20209
rect 56202 20209 56404 20226
rect 56960 20226 56976 20243
rect 57406 20243 57994 20259
rect 57406 20226 57422 20243
rect 56960 20209 57162 20226
rect 56202 20162 57162 20209
rect 57220 20209 57422 20226
rect 57978 20226 57994 20243
rect 57978 20209 58180 20226
rect 57220 20162 58180 20209
rect 59656 20123 60244 20139
rect 59656 20106 59672 20123
rect 59470 20089 59672 20106
rect 60228 20106 60244 20123
rect 60674 20123 61262 20139
rect 60674 20106 60690 20123
rect 60228 20089 60430 20106
rect 59470 20042 60430 20089
rect 60488 20089 60690 20106
rect 61246 20106 61262 20123
rect 61692 20123 62280 20139
rect 61692 20106 61708 20123
rect 61246 20089 61448 20106
rect 60488 20042 61448 20089
rect 61506 20089 61708 20106
rect 62264 20106 62280 20123
rect 62710 20123 63298 20139
rect 62710 20106 62726 20123
rect 62264 20089 62466 20106
rect 61506 20042 62466 20089
rect 62524 20089 62726 20106
rect 63282 20106 63298 20123
rect 63728 20123 64316 20139
rect 63728 20106 63744 20123
rect 63282 20089 63484 20106
rect 62524 20042 63484 20089
rect 63542 20089 63744 20106
rect 64300 20106 64316 20123
rect 64746 20123 65334 20139
rect 64746 20106 64762 20123
rect 64300 20089 64502 20106
rect 63542 20042 64502 20089
rect 64560 20089 64762 20106
rect 65318 20106 65334 20123
rect 65764 20123 66352 20139
rect 65764 20106 65780 20123
rect 65318 20089 65520 20106
rect 64560 20042 65520 20089
rect 65578 20089 65780 20106
rect 66336 20106 66352 20123
rect 66782 20123 67370 20139
rect 66782 20106 66798 20123
rect 66336 20089 66538 20106
rect 65578 20042 66538 20089
rect 66596 20089 66798 20106
rect 67354 20106 67370 20123
rect 67800 20123 68388 20139
rect 67800 20106 67816 20123
rect 67354 20089 67556 20106
rect 66596 20042 67556 20089
rect 67614 20089 67816 20106
rect 68372 20106 68388 20123
rect 68818 20123 69406 20139
rect 68818 20106 68834 20123
rect 68372 20089 68574 20106
rect 67614 20042 68574 20089
rect 68632 20089 68834 20106
rect 69390 20106 69406 20123
rect 69836 20123 70424 20139
rect 69836 20106 69852 20123
rect 69390 20089 69592 20106
rect 68632 20042 69592 20089
rect 69650 20089 69852 20106
rect 70408 20106 70424 20123
rect 70854 20123 71442 20139
rect 70854 20106 70870 20123
rect 70408 20089 70610 20106
rect 69650 20042 70610 20089
rect 70668 20089 70870 20106
rect 71426 20106 71442 20123
rect 71872 20123 72460 20139
rect 71872 20106 71888 20123
rect 71426 20089 71628 20106
rect 70668 20042 71628 20089
rect 71686 20089 71888 20106
rect 72444 20106 72460 20123
rect 72890 20123 73478 20139
rect 72890 20106 72906 20123
rect 72444 20089 72646 20106
rect 71686 20042 72646 20089
rect 72704 20089 72906 20106
rect 73462 20106 73478 20123
rect 73908 20123 74496 20139
rect 73908 20106 73924 20123
rect 73462 20089 73664 20106
rect 72704 20042 73664 20089
rect 73722 20089 73924 20106
rect 74480 20106 74496 20123
rect 74480 20089 74682 20106
rect 73722 20042 74682 20089
rect 54166 19515 55126 19562
rect 54166 19498 54368 19515
rect 54352 19481 54368 19498
rect 54924 19498 55126 19515
rect 55184 19515 56144 19562
rect 55184 19498 55386 19515
rect 54924 19481 54940 19498
rect 54352 19465 54940 19481
rect 55370 19481 55386 19498
rect 55942 19498 56144 19515
rect 56202 19515 57162 19562
rect 56202 19498 56404 19515
rect 55942 19481 55958 19498
rect 55370 19465 55958 19481
rect 56388 19481 56404 19498
rect 56960 19498 57162 19515
rect 57220 19515 58180 19562
rect 57220 19498 57422 19515
rect 56960 19481 56976 19498
rect 56388 19465 56976 19481
rect 57406 19481 57422 19498
rect 57978 19498 58180 19515
rect 57978 19481 57994 19498
rect 57406 19465 57994 19481
rect 59470 19395 60430 19442
rect 59470 19378 59672 19395
rect 59656 19361 59672 19378
rect 60228 19378 60430 19395
rect 60488 19395 61448 19442
rect 60488 19378 60690 19395
rect 60228 19361 60244 19378
rect 59656 19345 60244 19361
rect 60674 19361 60690 19378
rect 61246 19378 61448 19395
rect 61506 19395 62466 19442
rect 61506 19378 61708 19395
rect 61246 19361 61262 19378
rect 60674 19345 61262 19361
rect 61692 19361 61708 19378
rect 62264 19378 62466 19395
rect 62524 19395 63484 19442
rect 62524 19378 62726 19395
rect 62264 19361 62280 19378
rect 61692 19345 62280 19361
rect 62710 19361 62726 19378
rect 63282 19378 63484 19395
rect 63542 19395 64502 19442
rect 63542 19378 63744 19395
rect 63282 19361 63298 19378
rect 62710 19345 63298 19361
rect 63728 19361 63744 19378
rect 64300 19378 64502 19395
rect 64560 19395 65520 19442
rect 64560 19378 64762 19395
rect 64300 19361 64316 19378
rect 63728 19345 64316 19361
rect 64746 19361 64762 19378
rect 65318 19378 65520 19395
rect 65578 19395 66538 19442
rect 65578 19378 65780 19395
rect 65318 19361 65334 19378
rect 64746 19345 65334 19361
rect 65764 19361 65780 19378
rect 66336 19378 66538 19395
rect 66596 19395 67556 19442
rect 66596 19378 66798 19395
rect 66336 19361 66352 19378
rect 65764 19345 66352 19361
rect 66782 19361 66798 19378
rect 67354 19378 67556 19395
rect 67614 19395 68574 19442
rect 67614 19378 67816 19395
rect 67354 19361 67370 19378
rect 66782 19345 67370 19361
rect 67800 19361 67816 19378
rect 68372 19378 68574 19395
rect 68632 19395 69592 19442
rect 68632 19378 68834 19395
rect 68372 19361 68388 19378
rect 67800 19345 68388 19361
rect 68818 19361 68834 19378
rect 69390 19378 69592 19395
rect 69650 19395 70610 19442
rect 69650 19378 69852 19395
rect 69390 19361 69406 19378
rect 68818 19345 69406 19361
rect 69836 19361 69852 19378
rect 70408 19378 70610 19395
rect 70668 19395 71628 19442
rect 70668 19378 70870 19395
rect 70408 19361 70424 19378
rect 69836 19345 70424 19361
rect 70854 19361 70870 19378
rect 71426 19378 71628 19395
rect 71686 19395 72646 19442
rect 71686 19378 71888 19395
rect 71426 19361 71442 19378
rect 70854 19345 71442 19361
rect 71872 19361 71888 19378
rect 72444 19378 72646 19395
rect 72704 19395 73664 19442
rect 72704 19378 72906 19395
rect 72444 19361 72460 19378
rect 71872 19345 72460 19361
rect 72890 19361 72906 19378
rect 73462 19378 73664 19395
rect 73722 19395 74682 19442
rect 73722 19378 73924 19395
rect 73462 19361 73478 19378
rect 72890 19345 73478 19361
rect 73908 19361 73924 19378
rect 74480 19378 74682 19395
rect 74480 19361 74496 19378
rect 73908 19345 74496 19361
rect 54352 19211 54940 19227
rect 54352 19194 54368 19211
rect 54166 19177 54368 19194
rect 54924 19194 54940 19211
rect 55370 19211 55958 19227
rect 55370 19194 55386 19211
rect 54924 19177 55126 19194
rect 54166 19130 55126 19177
rect 55184 19177 55386 19194
rect 55942 19194 55958 19211
rect 56388 19211 56976 19227
rect 56388 19194 56404 19211
rect 55942 19177 56144 19194
rect 55184 19130 56144 19177
rect 56202 19177 56404 19194
rect 56960 19194 56976 19211
rect 57406 19211 57994 19227
rect 57406 19194 57422 19211
rect 56960 19177 57162 19194
rect 56202 19130 57162 19177
rect 57220 19177 57422 19194
rect 57978 19194 57994 19211
rect 57978 19177 58180 19194
rect 57220 19130 58180 19177
rect 59656 18867 60244 18883
rect 59656 18850 59672 18867
rect 59470 18833 59672 18850
rect 60228 18850 60244 18867
rect 60674 18867 61262 18883
rect 60674 18850 60690 18867
rect 60228 18833 60430 18850
rect 59470 18786 60430 18833
rect 60488 18833 60690 18850
rect 61246 18850 61262 18867
rect 61692 18867 62280 18883
rect 61692 18850 61708 18867
rect 61246 18833 61448 18850
rect 60488 18786 61448 18833
rect 61506 18833 61708 18850
rect 62264 18850 62280 18867
rect 62710 18867 63298 18883
rect 62710 18850 62726 18867
rect 62264 18833 62466 18850
rect 61506 18786 62466 18833
rect 62524 18833 62726 18850
rect 63282 18850 63298 18867
rect 63728 18867 64316 18883
rect 63728 18850 63744 18867
rect 63282 18833 63484 18850
rect 62524 18786 63484 18833
rect 63542 18833 63744 18850
rect 64300 18850 64316 18867
rect 64746 18867 65334 18883
rect 64746 18850 64762 18867
rect 64300 18833 64502 18850
rect 63542 18786 64502 18833
rect 64560 18833 64762 18850
rect 65318 18850 65334 18867
rect 65764 18867 66352 18883
rect 65764 18850 65780 18867
rect 65318 18833 65520 18850
rect 64560 18786 65520 18833
rect 65578 18833 65780 18850
rect 66336 18850 66352 18867
rect 66782 18867 67370 18883
rect 66782 18850 66798 18867
rect 66336 18833 66538 18850
rect 65578 18786 66538 18833
rect 66596 18833 66798 18850
rect 67354 18850 67370 18867
rect 67800 18867 68388 18883
rect 67800 18850 67816 18867
rect 67354 18833 67556 18850
rect 66596 18786 67556 18833
rect 67614 18833 67816 18850
rect 68372 18850 68388 18867
rect 68818 18867 69406 18883
rect 68818 18850 68834 18867
rect 68372 18833 68574 18850
rect 67614 18786 68574 18833
rect 68632 18833 68834 18850
rect 69390 18850 69406 18867
rect 69836 18867 70424 18883
rect 69836 18850 69852 18867
rect 69390 18833 69592 18850
rect 68632 18786 69592 18833
rect 69650 18833 69852 18850
rect 70408 18850 70424 18867
rect 70854 18867 71442 18883
rect 70854 18850 70870 18867
rect 70408 18833 70610 18850
rect 69650 18786 70610 18833
rect 70668 18833 70870 18850
rect 71426 18850 71442 18867
rect 71872 18867 72460 18883
rect 71872 18850 71888 18867
rect 71426 18833 71628 18850
rect 70668 18786 71628 18833
rect 71686 18833 71888 18850
rect 72444 18850 72460 18867
rect 72890 18867 73478 18883
rect 72890 18850 72906 18867
rect 72444 18833 72646 18850
rect 71686 18786 72646 18833
rect 72704 18833 72906 18850
rect 73462 18850 73478 18867
rect 73908 18867 74496 18883
rect 73908 18850 73924 18867
rect 73462 18833 73664 18850
rect 72704 18786 73664 18833
rect 73722 18833 73924 18850
rect 74480 18850 74496 18867
rect 74480 18833 74682 18850
rect 73722 18786 74682 18833
rect 54166 18483 55126 18530
rect 54166 18466 54368 18483
rect 54352 18449 54368 18466
rect 54924 18466 55126 18483
rect 55184 18483 56144 18530
rect 55184 18466 55386 18483
rect 54924 18449 54940 18466
rect 54352 18433 54940 18449
rect 55370 18449 55386 18466
rect 55942 18466 56144 18483
rect 56202 18483 57162 18530
rect 56202 18466 56404 18483
rect 55942 18449 55958 18466
rect 55370 18433 55958 18449
rect 56388 18449 56404 18466
rect 56960 18466 57162 18483
rect 57220 18483 58180 18530
rect 57220 18466 57422 18483
rect 56960 18449 56976 18466
rect 56388 18433 56976 18449
rect 57406 18449 57422 18466
rect 57978 18466 58180 18483
rect 57978 18449 57994 18466
rect 57406 18433 57994 18449
rect 54352 18179 54940 18195
rect 54352 18162 54368 18179
rect 54166 18145 54368 18162
rect 54924 18162 54940 18179
rect 55370 18179 55958 18195
rect 55370 18162 55386 18179
rect 54924 18145 55126 18162
rect 54166 18098 55126 18145
rect 55184 18145 55386 18162
rect 55942 18162 55958 18179
rect 56388 18179 56976 18195
rect 56388 18162 56404 18179
rect 55942 18145 56144 18162
rect 55184 18098 56144 18145
rect 56202 18145 56404 18162
rect 56960 18162 56976 18179
rect 57406 18179 57994 18195
rect 57406 18162 57422 18179
rect 56960 18145 57162 18162
rect 56202 18098 57162 18145
rect 57220 18145 57422 18162
rect 57978 18162 57994 18179
rect 57978 18145 58180 18162
rect 57220 18098 58180 18145
rect 59470 18139 60430 18186
rect 59470 18122 59672 18139
rect 59656 18105 59672 18122
rect 60228 18122 60430 18139
rect 60488 18139 61448 18186
rect 60488 18122 60690 18139
rect 60228 18105 60244 18122
rect 59656 18089 60244 18105
rect 60674 18105 60690 18122
rect 61246 18122 61448 18139
rect 61506 18139 62466 18186
rect 61506 18122 61708 18139
rect 61246 18105 61262 18122
rect 60674 18089 61262 18105
rect 61692 18105 61708 18122
rect 62264 18122 62466 18139
rect 62524 18139 63484 18186
rect 62524 18122 62726 18139
rect 62264 18105 62280 18122
rect 61692 18089 62280 18105
rect 62710 18105 62726 18122
rect 63282 18122 63484 18139
rect 63542 18139 64502 18186
rect 63542 18122 63744 18139
rect 63282 18105 63298 18122
rect 62710 18089 63298 18105
rect 63728 18105 63744 18122
rect 64300 18122 64502 18139
rect 64560 18139 65520 18186
rect 64560 18122 64762 18139
rect 64300 18105 64316 18122
rect 63728 18089 64316 18105
rect 64746 18105 64762 18122
rect 65318 18122 65520 18139
rect 65578 18139 66538 18186
rect 65578 18122 65780 18139
rect 65318 18105 65334 18122
rect 64746 18089 65334 18105
rect 65764 18105 65780 18122
rect 66336 18122 66538 18139
rect 66596 18139 67556 18186
rect 66596 18122 66798 18139
rect 66336 18105 66352 18122
rect 65764 18089 66352 18105
rect 66782 18105 66798 18122
rect 67354 18122 67556 18139
rect 67614 18139 68574 18186
rect 67614 18122 67816 18139
rect 67354 18105 67370 18122
rect 66782 18089 67370 18105
rect 67800 18105 67816 18122
rect 68372 18122 68574 18139
rect 68632 18139 69592 18186
rect 68632 18122 68834 18139
rect 68372 18105 68388 18122
rect 67800 18089 68388 18105
rect 68818 18105 68834 18122
rect 69390 18122 69592 18139
rect 69650 18139 70610 18186
rect 69650 18122 69852 18139
rect 69390 18105 69406 18122
rect 68818 18089 69406 18105
rect 69836 18105 69852 18122
rect 70408 18122 70610 18139
rect 70668 18139 71628 18186
rect 70668 18122 70870 18139
rect 70408 18105 70424 18122
rect 69836 18089 70424 18105
rect 70854 18105 70870 18122
rect 71426 18122 71628 18139
rect 71686 18139 72646 18186
rect 71686 18122 71888 18139
rect 71426 18105 71442 18122
rect 70854 18089 71442 18105
rect 71872 18105 71888 18122
rect 72444 18122 72646 18139
rect 72704 18139 73664 18186
rect 72704 18122 72906 18139
rect 72444 18105 72460 18122
rect 71872 18089 72460 18105
rect 72890 18105 72906 18122
rect 73462 18122 73664 18139
rect 73722 18139 74682 18186
rect 73722 18122 73924 18139
rect 73462 18105 73478 18122
rect 72890 18089 73478 18105
rect 73908 18105 73924 18122
rect 74480 18122 74682 18139
rect 74480 18105 74496 18122
rect 73908 18089 74496 18105
rect 59656 17611 60244 17627
rect 59656 17594 59672 17611
rect 59470 17577 59672 17594
rect 60228 17594 60244 17611
rect 60674 17611 61262 17627
rect 60674 17594 60690 17611
rect 60228 17577 60430 17594
rect 59470 17530 60430 17577
rect 60488 17577 60690 17594
rect 61246 17594 61262 17611
rect 61692 17611 62280 17627
rect 61692 17594 61708 17611
rect 61246 17577 61448 17594
rect 60488 17530 61448 17577
rect 61506 17577 61708 17594
rect 62264 17594 62280 17611
rect 62710 17611 63298 17627
rect 62710 17594 62726 17611
rect 62264 17577 62466 17594
rect 61506 17530 62466 17577
rect 62524 17577 62726 17594
rect 63282 17594 63298 17611
rect 63728 17611 64316 17627
rect 63728 17594 63744 17611
rect 63282 17577 63484 17594
rect 62524 17530 63484 17577
rect 63542 17577 63744 17594
rect 64300 17594 64316 17611
rect 64746 17611 65334 17627
rect 64746 17594 64762 17611
rect 64300 17577 64502 17594
rect 63542 17530 64502 17577
rect 64560 17577 64762 17594
rect 65318 17594 65334 17611
rect 65764 17611 66352 17627
rect 65764 17594 65780 17611
rect 65318 17577 65520 17594
rect 64560 17530 65520 17577
rect 65578 17577 65780 17594
rect 66336 17594 66352 17611
rect 66782 17611 67370 17627
rect 66782 17594 66798 17611
rect 66336 17577 66538 17594
rect 65578 17530 66538 17577
rect 66596 17577 66798 17594
rect 67354 17594 67370 17611
rect 67800 17611 68388 17627
rect 67800 17594 67816 17611
rect 67354 17577 67556 17594
rect 66596 17530 67556 17577
rect 67614 17577 67816 17594
rect 68372 17594 68388 17611
rect 68818 17611 69406 17627
rect 68818 17594 68834 17611
rect 68372 17577 68574 17594
rect 67614 17530 68574 17577
rect 68632 17577 68834 17594
rect 69390 17594 69406 17611
rect 69836 17611 70424 17627
rect 69836 17594 69852 17611
rect 69390 17577 69592 17594
rect 68632 17530 69592 17577
rect 69650 17577 69852 17594
rect 70408 17594 70424 17611
rect 70854 17611 71442 17627
rect 70854 17594 70870 17611
rect 70408 17577 70610 17594
rect 69650 17530 70610 17577
rect 70668 17577 70870 17594
rect 71426 17594 71442 17611
rect 71872 17611 72460 17627
rect 71872 17594 71888 17611
rect 71426 17577 71628 17594
rect 70668 17530 71628 17577
rect 71686 17577 71888 17594
rect 72444 17594 72460 17611
rect 72890 17611 73478 17627
rect 72890 17594 72906 17611
rect 72444 17577 72646 17594
rect 71686 17530 72646 17577
rect 72704 17577 72906 17594
rect 73462 17594 73478 17611
rect 73908 17611 74496 17627
rect 73908 17594 73924 17611
rect 73462 17577 73664 17594
rect 72704 17530 73664 17577
rect 73722 17577 73924 17594
rect 74480 17594 74496 17611
rect 74480 17577 74682 17594
rect 73722 17530 74682 17577
rect 54166 17451 55126 17498
rect 54166 17434 54368 17451
rect 54352 17417 54368 17434
rect 54924 17434 55126 17451
rect 55184 17451 56144 17498
rect 55184 17434 55386 17451
rect 54924 17417 54940 17434
rect 54352 17401 54940 17417
rect 55370 17417 55386 17434
rect 55942 17434 56144 17451
rect 56202 17451 57162 17498
rect 56202 17434 56404 17451
rect 55942 17417 55958 17434
rect 55370 17401 55958 17417
rect 56388 17417 56404 17434
rect 56960 17434 57162 17451
rect 57220 17451 58180 17498
rect 57220 17434 57422 17451
rect 56960 17417 56976 17434
rect 56388 17401 56976 17417
rect 57406 17417 57422 17434
rect 57978 17434 58180 17451
rect 57978 17417 57994 17434
rect 57406 17401 57994 17417
rect 59470 16883 60430 16930
rect 59470 16866 59672 16883
rect 59656 16849 59672 16866
rect 60228 16866 60430 16883
rect 60488 16883 61448 16930
rect 60488 16866 60690 16883
rect 60228 16849 60244 16866
rect 59656 16833 60244 16849
rect 60674 16849 60690 16866
rect 61246 16866 61448 16883
rect 61506 16883 62466 16930
rect 61506 16866 61708 16883
rect 61246 16849 61262 16866
rect 60674 16833 61262 16849
rect 61692 16849 61708 16866
rect 62264 16866 62466 16883
rect 62524 16883 63484 16930
rect 62524 16866 62726 16883
rect 62264 16849 62280 16866
rect 61692 16833 62280 16849
rect 62710 16849 62726 16866
rect 63282 16866 63484 16883
rect 63542 16883 64502 16930
rect 63542 16866 63744 16883
rect 63282 16849 63298 16866
rect 62710 16833 63298 16849
rect 63728 16849 63744 16866
rect 64300 16866 64502 16883
rect 64560 16883 65520 16930
rect 64560 16866 64762 16883
rect 64300 16849 64316 16866
rect 63728 16833 64316 16849
rect 64746 16849 64762 16866
rect 65318 16866 65520 16883
rect 65578 16883 66538 16930
rect 65578 16866 65780 16883
rect 65318 16849 65334 16866
rect 64746 16833 65334 16849
rect 65764 16849 65780 16866
rect 66336 16866 66538 16883
rect 66596 16883 67556 16930
rect 66596 16866 66798 16883
rect 66336 16849 66352 16866
rect 65764 16833 66352 16849
rect 66782 16849 66798 16866
rect 67354 16866 67556 16883
rect 67614 16883 68574 16930
rect 67614 16866 67816 16883
rect 67354 16849 67370 16866
rect 66782 16833 67370 16849
rect 67800 16849 67816 16866
rect 68372 16866 68574 16883
rect 68632 16883 69592 16930
rect 68632 16866 68834 16883
rect 68372 16849 68388 16866
rect 67800 16833 68388 16849
rect 68818 16849 68834 16866
rect 69390 16866 69592 16883
rect 69650 16883 70610 16930
rect 69650 16866 69852 16883
rect 69390 16849 69406 16866
rect 68818 16833 69406 16849
rect 69836 16849 69852 16866
rect 70408 16866 70610 16883
rect 70668 16883 71628 16930
rect 70668 16866 70870 16883
rect 70408 16849 70424 16866
rect 69836 16833 70424 16849
rect 70854 16849 70870 16866
rect 71426 16866 71628 16883
rect 71686 16883 72646 16930
rect 71686 16866 71888 16883
rect 71426 16849 71442 16866
rect 70854 16833 71442 16849
rect 71872 16849 71888 16866
rect 72444 16866 72646 16883
rect 72704 16883 73664 16930
rect 72704 16866 72906 16883
rect 72444 16849 72460 16866
rect 71872 16833 72460 16849
rect 72890 16849 72906 16866
rect 73462 16866 73664 16883
rect 73722 16883 74682 16930
rect 73722 16866 73924 16883
rect 73462 16849 73478 16866
rect 72890 16833 73478 16849
rect 73908 16849 73924 16866
rect 74480 16866 74682 16883
rect 74480 16849 74496 16866
rect 73908 16833 74496 16849
rect 13764 14406 14352 14422
rect 13764 14389 13780 14406
rect 13578 14372 13780 14389
rect 14336 14389 14352 14406
rect 14782 14406 15370 14422
rect 14782 14389 14798 14406
rect 14336 14372 14538 14389
rect 13578 14334 14538 14372
rect 14596 14372 14798 14389
rect 15354 14389 15370 14406
rect 15800 14406 16388 14422
rect 15800 14389 15816 14406
rect 15354 14372 15556 14389
rect 14596 14334 15556 14372
rect 15614 14372 15816 14389
rect 16372 14389 16388 14406
rect 16818 14406 17406 14422
rect 16818 14389 16834 14406
rect 16372 14372 16574 14389
rect 15614 14334 16574 14372
rect 16632 14372 16834 14389
rect 17390 14389 17406 14406
rect 17836 14406 18424 14422
rect 17836 14389 17852 14406
rect 17390 14372 17592 14389
rect 16632 14334 17592 14372
rect 17650 14372 17852 14389
rect 18408 14389 18424 14406
rect 18854 14406 19442 14422
rect 18854 14389 18870 14406
rect 18408 14372 18610 14389
rect 17650 14334 18610 14372
rect 18668 14372 18870 14389
rect 19426 14389 19442 14406
rect 19872 14406 20460 14422
rect 19872 14389 19888 14406
rect 19426 14372 19628 14389
rect 18668 14334 19628 14372
rect 19686 14372 19888 14389
rect 20444 14389 20460 14406
rect 20890 14406 21478 14422
rect 20890 14389 20906 14406
rect 20444 14372 20646 14389
rect 19686 14334 20646 14372
rect 20704 14372 20906 14389
rect 21462 14389 21478 14406
rect 21908 14406 22496 14422
rect 21908 14389 21924 14406
rect 21462 14372 21664 14389
rect 20704 14334 21664 14372
rect 21722 14372 21924 14389
rect 22480 14389 22496 14406
rect 22926 14406 23514 14422
rect 22926 14389 22942 14406
rect 22480 14372 22682 14389
rect 21722 14334 22682 14372
rect 22740 14372 22942 14389
rect 23498 14389 23514 14406
rect 23944 14406 24532 14422
rect 23944 14389 23960 14406
rect 23498 14372 23700 14389
rect 22740 14334 23700 14372
rect 23758 14372 23960 14389
rect 24516 14389 24532 14406
rect 24962 14406 25550 14422
rect 24962 14389 24978 14406
rect 24516 14372 24718 14389
rect 23758 14334 24718 14372
rect 24776 14372 24978 14389
rect 25534 14389 25550 14406
rect 25980 14406 26568 14422
rect 25980 14389 25996 14406
rect 25534 14372 25736 14389
rect 24776 14334 25736 14372
rect 25794 14372 25996 14389
rect 26552 14389 26568 14406
rect 26998 14406 27586 14422
rect 26998 14389 27014 14406
rect 26552 14372 26754 14389
rect 25794 14334 26754 14372
rect 26812 14372 27014 14389
rect 27570 14389 27586 14406
rect 28016 14406 28604 14422
rect 28016 14389 28032 14406
rect 27570 14372 27772 14389
rect 26812 14334 27772 14372
rect 27830 14372 28032 14389
rect 28588 14389 28604 14406
rect 29034 14406 29622 14422
rect 29034 14389 29050 14406
rect 28588 14372 28790 14389
rect 27830 14334 28790 14372
rect 28848 14372 29050 14389
rect 29606 14389 29622 14406
rect 30052 14406 30640 14422
rect 30052 14389 30068 14406
rect 29606 14372 29808 14389
rect 28848 14334 29808 14372
rect 29866 14372 30068 14389
rect 30624 14389 30640 14406
rect 31070 14406 31658 14422
rect 31070 14389 31086 14406
rect 30624 14372 30826 14389
rect 29866 14334 30826 14372
rect 30884 14372 31086 14389
rect 31642 14389 31658 14406
rect 32088 14406 32676 14422
rect 32088 14389 32104 14406
rect 31642 14372 31844 14389
rect 30884 14334 31844 14372
rect 31902 14372 32104 14389
rect 32660 14389 32676 14406
rect 33106 14406 33694 14422
rect 33106 14389 33122 14406
rect 32660 14372 32862 14389
rect 31902 14334 32862 14372
rect 32920 14372 33122 14389
rect 33678 14389 33694 14406
rect 33678 14372 33880 14389
rect 32920 14334 33880 14372
rect 1998 13930 2586 13946
rect 1998 13913 2014 13930
rect 1812 13896 2014 13913
rect 2570 13913 2586 13930
rect 3016 13930 3604 13946
rect 3016 13913 3032 13930
rect 2570 13896 2772 13913
rect 1812 13858 2772 13896
rect 2830 13896 3032 13913
rect 3588 13913 3604 13930
rect 4034 13930 4622 13946
rect 4034 13913 4050 13930
rect 3588 13896 3790 13913
rect 2830 13858 3790 13896
rect 3848 13896 4050 13913
rect 4606 13913 4622 13930
rect 5052 13930 5640 13946
rect 5052 13913 5068 13930
rect 4606 13896 4808 13913
rect 3848 13858 4808 13896
rect 4866 13896 5068 13913
rect 5624 13913 5640 13930
rect 6070 13930 6658 13946
rect 6070 13913 6086 13930
rect 5624 13896 5826 13913
rect 4866 13858 5826 13896
rect 5884 13896 6086 13913
rect 6642 13913 6658 13930
rect 7088 13930 7676 13946
rect 7088 13913 7104 13930
rect 6642 13896 6844 13913
rect 5884 13858 6844 13896
rect 6902 13896 7104 13913
rect 7660 13913 7676 13930
rect 8106 13930 8694 13946
rect 8106 13913 8122 13930
rect 7660 13896 7862 13913
rect 6902 13858 7862 13896
rect 7920 13896 8122 13913
rect 8678 13913 8694 13930
rect 9124 13930 9712 13946
rect 9124 13913 9140 13930
rect 8678 13896 8880 13913
rect 7920 13858 8880 13896
rect 8938 13896 9140 13913
rect 9696 13913 9712 13930
rect 10142 13930 10730 13946
rect 10142 13913 10158 13930
rect 9696 13896 9898 13913
rect 8938 13858 9898 13896
rect 9956 13896 10158 13913
rect 10714 13913 10730 13930
rect 10714 13896 10916 13913
rect 9956 13858 10916 13896
rect 13578 13696 14538 13734
rect 13578 13679 13780 13696
rect 13764 13662 13780 13679
rect 14336 13679 14538 13696
rect 14596 13696 15556 13734
rect 14596 13679 14798 13696
rect 14336 13662 14352 13679
rect 13764 13646 14352 13662
rect 14782 13662 14798 13679
rect 15354 13679 15556 13696
rect 15614 13696 16574 13734
rect 15614 13679 15816 13696
rect 15354 13662 15370 13679
rect 14782 13646 15370 13662
rect 15800 13662 15816 13679
rect 16372 13679 16574 13696
rect 16632 13696 17592 13734
rect 16632 13679 16834 13696
rect 16372 13662 16388 13679
rect 15800 13646 16388 13662
rect 16818 13662 16834 13679
rect 17390 13679 17592 13696
rect 17650 13696 18610 13734
rect 17650 13679 17852 13696
rect 17390 13662 17406 13679
rect 16818 13646 17406 13662
rect 17836 13662 17852 13679
rect 18408 13679 18610 13696
rect 18668 13696 19628 13734
rect 18668 13679 18870 13696
rect 18408 13662 18424 13679
rect 17836 13646 18424 13662
rect 18854 13662 18870 13679
rect 19426 13679 19628 13696
rect 19686 13696 20646 13734
rect 19686 13679 19888 13696
rect 19426 13662 19442 13679
rect 18854 13646 19442 13662
rect 19872 13662 19888 13679
rect 20444 13679 20646 13696
rect 20704 13696 21664 13734
rect 20704 13679 20906 13696
rect 20444 13662 20460 13679
rect 19872 13646 20460 13662
rect 20890 13662 20906 13679
rect 21462 13679 21664 13696
rect 21722 13696 22682 13734
rect 21722 13679 21924 13696
rect 21462 13662 21478 13679
rect 20890 13646 21478 13662
rect 21908 13662 21924 13679
rect 22480 13679 22682 13696
rect 22740 13696 23700 13734
rect 22740 13679 22942 13696
rect 22480 13662 22496 13679
rect 21908 13646 22496 13662
rect 22926 13662 22942 13679
rect 23498 13679 23700 13696
rect 23758 13696 24718 13734
rect 23758 13679 23960 13696
rect 23498 13662 23514 13679
rect 22926 13646 23514 13662
rect 23944 13662 23960 13679
rect 24516 13679 24718 13696
rect 24776 13696 25736 13734
rect 24776 13679 24978 13696
rect 24516 13662 24532 13679
rect 23944 13646 24532 13662
rect 24962 13662 24978 13679
rect 25534 13679 25736 13696
rect 25794 13696 26754 13734
rect 25794 13679 25996 13696
rect 25534 13662 25550 13679
rect 24962 13646 25550 13662
rect 25980 13662 25996 13679
rect 26552 13679 26754 13696
rect 26812 13696 27772 13734
rect 26812 13679 27014 13696
rect 26552 13662 26568 13679
rect 25980 13646 26568 13662
rect 26998 13662 27014 13679
rect 27570 13679 27772 13696
rect 27830 13696 28790 13734
rect 27830 13679 28032 13696
rect 27570 13662 27586 13679
rect 26998 13646 27586 13662
rect 28016 13662 28032 13679
rect 28588 13679 28790 13696
rect 28848 13696 29808 13734
rect 28848 13679 29050 13696
rect 28588 13662 28604 13679
rect 28016 13646 28604 13662
rect 29034 13662 29050 13679
rect 29606 13679 29808 13696
rect 29866 13696 30826 13734
rect 29866 13679 30068 13696
rect 29606 13662 29622 13679
rect 29034 13646 29622 13662
rect 30052 13662 30068 13679
rect 30624 13679 30826 13696
rect 30884 13696 31844 13734
rect 30884 13679 31086 13696
rect 30624 13662 30640 13679
rect 30052 13646 30640 13662
rect 31070 13662 31086 13679
rect 31642 13679 31844 13696
rect 31902 13696 32862 13734
rect 31902 13679 32104 13696
rect 31642 13662 31658 13679
rect 31070 13646 31658 13662
rect 32088 13662 32104 13679
rect 32660 13679 32862 13696
rect 32920 13696 33880 13734
rect 32920 13679 33122 13696
rect 32660 13662 32676 13679
rect 32088 13646 32676 13662
rect 33106 13662 33122 13679
rect 33678 13679 33880 13696
rect 33678 13662 33694 13679
rect 33106 13646 33694 13662
rect 13764 13588 14352 13604
rect 13764 13571 13780 13588
rect 13578 13554 13780 13571
rect 14336 13571 14352 13588
rect 14782 13588 15370 13604
rect 14782 13571 14798 13588
rect 14336 13554 14538 13571
rect 13578 13516 14538 13554
rect 14596 13554 14798 13571
rect 15354 13571 15370 13588
rect 15800 13588 16388 13604
rect 15800 13571 15816 13588
rect 15354 13554 15556 13571
rect 14596 13516 15556 13554
rect 15614 13554 15816 13571
rect 16372 13571 16388 13588
rect 16818 13588 17406 13604
rect 16818 13571 16834 13588
rect 16372 13554 16574 13571
rect 15614 13516 16574 13554
rect 16632 13554 16834 13571
rect 17390 13571 17406 13588
rect 17836 13588 18424 13604
rect 17836 13571 17852 13588
rect 17390 13554 17592 13571
rect 16632 13516 17592 13554
rect 17650 13554 17852 13571
rect 18408 13571 18424 13588
rect 18854 13588 19442 13604
rect 18854 13571 18870 13588
rect 18408 13554 18610 13571
rect 17650 13516 18610 13554
rect 18668 13554 18870 13571
rect 19426 13571 19442 13588
rect 19872 13588 20460 13604
rect 19872 13571 19888 13588
rect 19426 13554 19628 13571
rect 18668 13516 19628 13554
rect 19686 13554 19888 13571
rect 20444 13571 20460 13588
rect 20890 13588 21478 13604
rect 20890 13571 20906 13588
rect 20444 13554 20646 13571
rect 19686 13516 20646 13554
rect 20704 13554 20906 13571
rect 21462 13571 21478 13588
rect 21908 13588 22496 13604
rect 21908 13571 21924 13588
rect 21462 13554 21664 13571
rect 20704 13516 21664 13554
rect 21722 13554 21924 13571
rect 22480 13571 22496 13588
rect 22926 13588 23514 13604
rect 22926 13571 22942 13588
rect 22480 13554 22682 13571
rect 21722 13516 22682 13554
rect 22740 13554 22942 13571
rect 23498 13571 23514 13588
rect 23944 13588 24532 13604
rect 23944 13571 23960 13588
rect 23498 13554 23700 13571
rect 22740 13516 23700 13554
rect 23758 13554 23960 13571
rect 24516 13571 24532 13588
rect 24962 13588 25550 13604
rect 24962 13571 24978 13588
rect 24516 13554 24718 13571
rect 23758 13516 24718 13554
rect 24776 13554 24978 13571
rect 25534 13571 25550 13588
rect 25980 13588 26568 13604
rect 25980 13571 25996 13588
rect 25534 13554 25736 13571
rect 24776 13516 25736 13554
rect 25794 13554 25996 13571
rect 26552 13571 26568 13588
rect 26998 13588 27586 13604
rect 26998 13571 27014 13588
rect 26552 13554 26754 13571
rect 25794 13516 26754 13554
rect 26812 13554 27014 13571
rect 27570 13571 27586 13588
rect 28016 13588 28604 13604
rect 28016 13571 28032 13588
rect 27570 13554 27772 13571
rect 26812 13516 27772 13554
rect 27830 13554 28032 13571
rect 28588 13571 28604 13588
rect 29034 13588 29622 13604
rect 29034 13571 29050 13588
rect 28588 13554 28790 13571
rect 27830 13516 28790 13554
rect 28848 13554 29050 13571
rect 29606 13571 29622 13588
rect 30052 13588 30640 13604
rect 30052 13571 30068 13588
rect 29606 13554 29808 13571
rect 28848 13516 29808 13554
rect 29866 13554 30068 13571
rect 30624 13571 30640 13588
rect 31070 13588 31658 13604
rect 31070 13571 31086 13588
rect 30624 13554 30826 13571
rect 29866 13516 30826 13554
rect 30884 13554 31086 13571
rect 31642 13571 31658 13588
rect 32088 13588 32676 13604
rect 32088 13571 32104 13588
rect 31642 13554 31844 13571
rect 30884 13516 31844 13554
rect 31902 13554 32104 13571
rect 32660 13571 32676 13588
rect 33106 13588 33694 13604
rect 33106 13571 33122 13588
rect 32660 13554 32862 13571
rect 31902 13516 32862 13554
rect 32920 13554 33122 13571
rect 33678 13571 33694 13588
rect 33678 13554 33880 13571
rect 32920 13516 33880 13554
rect 1812 13220 2772 13258
rect 1812 13203 2014 13220
rect 1998 13186 2014 13203
rect 2570 13203 2772 13220
rect 2830 13220 3790 13258
rect 2830 13203 3032 13220
rect 2570 13186 2586 13203
rect 1998 13170 2586 13186
rect 3016 13186 3032 13203
rect 3588 13203 3790 13220
rect 3848 13220 4808 13258
rect 3848 13203 4050 13220
rect 3588 13186 3604 13203
rect 3016 13170 3604 13186
rect 1998 13112 2586 13128
rect 1998 13095 2014 13112
rect 1812 13078 2014 13095
rect 2570 13095 2586 13112
rect 4034 13186 4050 13203
rect 4606 13203 4808 13220
rect 4866 13220 5826 13258
rect 4866 13203 5068 13220
rect 4606 13186 4622 13203
rect 4034 13170 4622 13186
rect 3016 13112 3604 13128
rect 3016 13095 3032 13112
rect 2570 13078 2772 13095
rect 1812 13040 2772 13078
rect 2830 13078 3032 13095
rect 3588 13095 3604 13112
rect 5052 13186 5068 13203
rect 5624 13203 5826 13220
rect 5884 13220 6844 13258
rect 5884 13203 6086 13220
rect 5624 13186 5640 13203
rect 5052 13170 5640 13186
rect 4034 13112 4622 13128
rect 4034 13095 4050 13112
rect 3588 13078 3790 13095
rect 2830 13040 3790 13078
rect 3848 13078 4050 13095
rect 4606 13095 4622 13112
rect 6070 13186 6086 13203
rect 6642 13203 6844 13220
rect 6902 13220 7862 13258
rect 6902 13203 7104 13220
rect 6642 13186 6658 13203
rect 6070 13170 6658 13186
rect 5052 13112 5640 13128
rect 5052 13095 5068 13112
rect 4606 13078 4808 13095
rect 3848 13040 4808 13078
rect 4866 13078 5068 13095
rect 5624 13095 5640 13112
rect 7088 13186 7104 13203
rect 7660 13203 7862 13220
rect 7920 13220 8880 13258
rect 7920 13203 8122 13220
rect 7660 13186 7676 13203
rect 7088 13170 7676 13186
rect 6070 13112 6658 13128
rect 6070 13095 6086 13112
rect 5624 13078 5826 13095
rect 4866 13040 5826 13078
rect 5884 13078 6086 13095
rect 6642 13095 6658 13112
rect 8106 13186 8122 13203
rect 8678 13203 8880 13220
rect 8938 13220 9898 13258
rect 8938 13203 9140 13220
rect 8678 13186 8694 13203
rect 8106 13170 8694 13186
rect 7088 13112 7676 13128
rect 7088 13095 7104 13112
rect 6642 13078 6844 13095
rect 5884 13040 6844 13078
rect 6902 13078 7104 13095
rect 7660 13095 7676 13112
rect 9124 13186 9140 13203
rect 9696 13203 9898 13220
rect 9956 13220 10916 13258
rect 9956 13203 10158 13220
rect 9696 13186 9712 13203
rect 9124 13170 9712 13186
rect 8106 13112 8694 13128
rect 8106 13095 8122 13112
rect 7660 13078 7862 13095
rect 6902 13040 7862 13078
rect 7920 13078 8122 13095
rect 8678 13095 8694 13112
rect 10142 13186 10158 13203
rect 10714 13203 10916 13220
rect 10714 13186 10730 13203
rect 10142 13170 10730 13186
rect 9124 13112 9712 13128
rect 9124 13095 9140 13112
rect 8678 13078 8880 13095
rect 7920 13040 8880 13078
rect 8938 13078 9140 13095
rect 9696 13095 9712 13112
rect 10142 13112 10730 13128
rect 10142 13095 10158 13112
rect 9696 13078 9898 13095
rect 8938 13040 9898 13078
rect 9956 13078 10158 13095
rect 10714 13095 10730 13112
rect 10714 13078 10916 13095
rect 9956 13040 10916 13078
rect 13578 12878 14538 12916
rect 13578 12861 13780 12878
rect 13764 12844 13780 12861
rect 14336 12861 14538 12878
rect 14596 12878 15556 12916
rect 14596 12861 14798 12878
rect 14336 12844 14352 12861
rect 13764 12828 14352 12844
rect 14782 12844 14798 12861
rect 15354 12861 15556 12878
rect 15614 12878 16574 12916
rect 15614 12861 15816 12878
rect 15354 12844 15370 12861
rect 14782 12828 15370 12844
rect 15800 12844 15816 12861
rect 16372 12861 16574 12878
rect 16632 12878 17592 12916
rect 16632 12861 16834 12878
rect 16372 12844 16388 12861
rect 15800 12828 16388 12844
rect 16818 12844 16834 12861
rect 17390 12861 17592 12878
rect 17650 12878 18610 12916
rect 17650 12861 17852 12878
rect 17390 12844 17406 12861
rect 16818 12828 17406 12844
rect 17836 12844 17852 12861
rect 18408 12861 18610 12878
rect 18668 12878 19628 12916
rect 18668 12861 18870 12878
rect 18408 12844 18424 12861
rect 17836 12828 18424 12844
rect 18854 12844 18870 12861
rect 19426 12861 19628 12878
rect 19686 12878 20646 12916
rect 19686 12861 19888 12878
rect 19426 12844 19442 12861
rect 18854 12828 19442 12844
rect 19872 12844 19888 12861
rect 20444 12861 20646 12878
rect 20704 12878 21664 12916
rect 20704 12861 20906 12878
rect 20444 12844 20460 12861
rect 19872 12828 20460 12844
rect 20890 12844 20906 12861
rect 21462 12861 21664 12878
rect 21722 12878 22682 12916
rect 21722 12861 21924 12878
rect 21462 12844 21478 12861
rect 20890 12828 21478 12844
rect 21908 12844 21924 12861
rect 22480 12861 22682 12878
rect 22740 12878 23700 12916
rect 22740 12861 22942 12878
rect 22480 12844 22496 12861
rect 21908 12828 22496 12844
rect 22926 12844 22942 12861
rect 23498 12861 23700 12878
rect 23758 12878 24718 12916
rect 23758 12861 23960 12878
rect 23498 12844 23514 12861
rect 22926 12828 23514 12844
rect 23944 12844 23960 12861
rect 24516 12861 24718 12878
rect 24776 12878 25736 12916
rect 24776 12861 24978 12878
rect 24516 12844 24532 12861
rect 23944 12828 24532 12844
rect 24962 12844 24978 12861
rect 25534 12861 25736 12878
rect 25794 12878 26754 12916
rect 25794 12861 25996 12878
rect 25534 12844 25550 12861
rect 24962 12828 25550 12844
rect 25980 12844 25996 12861
rect 26552 12861 26754 12878
rect 26812 12878 27772 12916
rect 26812 12861 27014 12878
rect 26552 12844 26568 12861
rect 25980 12828 26568 12844
rect 26998 12844 27014 12861
rect 27570 12861 27772 12878
rect 27830 12878 28790 12916
rect 27830 12861 28032 12878
rect 27570 12844 27586 12861
rect 26998 12828 27586 12844
rect 28016 12844 28032 12861
rect 28588 12861 28790 12878
rect 28848 12878 29808 12916
rect 28848 12861 29050 12878
rect 28588 12844 28604 12861
rect 28016 12828 28604 12844
rect 29034 12844 29050 12861
rect 29606 12861 29808 12878
rect 29866 12878 30826 12916
rect 29866 12861 30068 12878
rect 29606 12844 29622 12861
rect 29034 12828 29622 12844
rect 30052 12844 30068 12861
rect 30624 12861 30826 12878
rect 30884 12878 31844 12916
rect 30884 12861 31086 12878
rect 30624 12844 30640 12861
rect 30052 12828 30640 12844
rect 31070 12844 31086 12861
rect 31642 12861 31844 12878
rect 31902 12878 32862 12916
rect 31902 12861 32104 12878
rect 31642 12844 31658 12861
rect 31070 12828 31658 12844
rect 32088 12844 32104 12861
rect 32660 12861 32862 12878
rect 32920 12878 33880 12916
rect 32920 12861 33122 12878
rect 32660 12844 32676 12861
rect 32088 12828 32676 12844
rect 33106 12844 33122 12861
rect 33678 12861 33880 12878
rect 33678 12844 33694 12861
rect 33106 12828 33694 12844
rect 1812 12402 2772 12440
rect 1812 12385 2014 12402
rect 1998 12368 2014 12385
rect 2570 12385 2772 12402
rect 2830 12402 3790 12440
rect 2830 12385 3032 12402
rect 2570 12368 2586 12385
rect 1998 12352 2586 12368
rect 3016 12368 3032 12385
rect 3588 12385 3790 12402
rect 3848 12402 4808 12440
rect 3848 12385 4050 12402
rect 3588 12368 3604 12385
rect 3016 12352 3604 12368
rect 1998 12294 2586 12310
rect 1998 12277 2014 12294
rect 1812 12260 2014 12277
rect 2570 12277 2586 12294
rect 4034 12368 4050 12385
rect 4606 12385 4808 12402
rect 4866 12402 5826 12440
rect 4866 12385 5068 12402
rect 4606 12368 4622 12385
rect 4034 12352 4622 12368
rect 3016 12294 3604 12310
rect 3016 12277 3032 12294
rect 2570 12260 2772 12277
rect 1812 12222 2772 12260
rect 2830 12260 3032 12277
rect 3588 12277 3604 12294
rect 5052 12368 5068 12385
rect 5624 12385 5826 12402
rect 5884 12402 6844 12440
rect 5884 12385 6086 12402
rect 5624 12368 5640 12385
rect 5052 12352 5640 12368
rect 4034 12294 4622 12310
rect 4034 12277 4050 12294
rect 3588 12260 3790 12277
rect 2830 12222 3790 12260
rect 3848 12260 4050 12277
rect 4606 12277 4622 12294
rect 6070 12368 6086 12385
rect 6642 12385 6844 12402
rect 6902 12402 7862 12440
rect 6902 12385 7104 12402
rect 6642 12368 6658 12385
rect 6070 12352 6658 12368
rect 5052 12294 5640 12310
rect 5052 12277 5068 12294
rect 4606 12260 4808 12277
rect 3848 12222 4808 12260
rect 4866 12260 5068 12277
rect 5624 12277 5640 12294
rect 7088 12368 7104 12385
rect 7660 12385 7862 12402
rect 7920 12402 8880 12440
rect 7920 12385 8122 12402
rect 7660 12368 7676 12385
rect 7088 12352 7676 12368
rect 6070 12294 6658 12310
rect 6070 12277 6086 12294
rect 5624 12260 5826 12277
rect 4866 12222 5826 12260
rect 5884 12260 6086 12277
rect 6642 12277 6658 12294
rect 8106 12368 8122 12385
rect 8678 12385 8880 12402
rect 8938 12402 9898 12440
rect 8938 12385 9140 12402
rect 8678 12368 8694 12385
rect 8106 12352 8694 12368
rect 7088 12294 7676 12310
rect 7088 12277 7104 12294
rect 6642 12260 6844 12277
rect 5884 12222 6844 12260
rect 6902 12260 7104 12277
rect 7660 12277 7676 12294
rect 9124 12368 9140 12385
rect 9696 12385 9898 12402
rect 9956 12402 10916 12440
rect 9956 12385 10158 12402
rect 9696 12368 9712 12385
rect 9124 12352 9712 12368
rect 8106 12294 8694 12310
rect 8106 12277 8122 12294
rect 7660 12260 7862 12277
rect 6902 12222 7862 12260
rect 7920 12260 8122 12277
rect 8678 12277 8694 12294
rect 10142 12368 10158 12385
rect 10714 12385 10916 12402
rect 10714 12368 10730 12385
rect 10142 12352 10730 12368
rect 9124 12294 9712 12310
rect 9124 12277 9140 12294
rect 8678 12260 8880 12277
rect 7920 12222 8880 12260
rect 8938 12260 9140 12277
rect 9696 12277 9712 12294
rect 10142 12294 10730 12310
rect 10142 12277 10158 12294
rect 9696 12260 9898 12277
rect 8938 12222 9898 12260
rect 9956 12260 10158 12277
rect 10714 12277 10730 12294
rect 10714 12260 10916 12277
rect 9956 12222 10916 12260
rect 13764 12210 14352 12226
rect 13764 12193 13780 12210
rect 13578 12176 13780 12193
rect 14336 12193 14352 12210
rect 14782 12210 15370 12226
rect 14782 12193 14798 12210
rect 14336 12176 14538 12193
rect 13578 12138 14538 12176
rect 14596 12176 14798 12193
rect 15354 12193 15370 12210
rect 15800 12210 16388 12226
rect 15800 12193 15816 12210
rect 15354 12176 15556 12193
rect 14596 12138 15556 12176
rect 15614 12176 15816 12193
rect 16372 12193 16388 12210
rect 16818 12210 17406 12226
rect 16818 12193 16834 12210
rect 16372 12176 16574 12193
rect 15614 12138 16574 12176
rect 16632 12176 16834 12193
rect 17390 12193 17406 12210
rect 17836 12210 18424 12226
rect 17836 12193 17852 12210
rect 17390 12176 17592 12193
rect 16632 12138 17592 12176
rect 17650 12176 17852 12193
rect 18408 12193 18424 12210
rect 18854 12210 19442 12226
rect 18854 12193 18870 12210
rect 18408 12176 18610 12193
rect 17650 12138 18610 12176
rect 18668 12176 18870 12193
rect 19426 12193 19442 12210
rect 19872 12210 20460 12226
rect 19872 12193 19888 12210
rect 19426 12176 19628 12193
rect 18668 12138 19628 12176
rect 19686 12176 19888 12193
rect 20444 12193 20460 12210
rect 20890 12210 21478 12226
rect 20890 12193 20906 12210
rect 20444 12176 20646 12193
rect 19686 12138 20646 12176
rect 20704 12176 20906 12193
rect 21462 12193 21478 12210
rect 21908 12210 22496 12226
rect 21908 12193 21924 12210
rect 21462 12176 21664 12193
rect 20704 12138 21664 12176
rect 21722 12176 21924 12193
rect 22480 12193 22496 12210
rect 22926 12210 23514 12226
rect 22926 12193 22942 12210
rect 22480 12176 22682 12193
rect 21722 12138 22682 12176
rect 22740 12176 22942 12193
rect 23498 12193 23514 12210
rect 23944 12210 24532 12226
rect 23944 12193 23960 12210
rect 23498 12176 23700 12193
rect 22740 12138 23700 12176
rect 23758 12176 23960 12193
rect 24516 12193 24532 12210
rect 24962 12210 25550 12226
rect 24962 12193 24978 12210
rect 24516 12176 24718 12193
rect 23758 12138 24718 12176
rect 24776 12176 24978 12193
rect 25534 12193 25550 12210
rect 25980 12210 26568 12226
rect 25980 12193 25996 12210
rect 25534 12176 25736 12193
rect 24776 12138 25736 12176
rect 25794 12176 25996 12193
rect 26552 12193 26568 12210
rect 26998 12210 27586 12226
rect 26998 12193 27014 12210
rect 26552 12176 26754 12193
rect 25794 12138 26754 12176
rect 26812 12176 27014 12193
rect 27570 12193 27586 12210
rect 28016 12210 28604 12226
rect 28016 12193 28032 12210
rect 27570 12176 27772 12193
rect 26812 12138 27772 12176
rect 27830 12176 28032 12193
rect 28588 12193 28604 12210
rect 29034 12210 29622 12226
rect 29034 12193 29050 12210
rect 28588 12176 28790 12193
rect 27830 12138 28790 12176
rect 28848 12176 29050 12193
rect 29606 12193 29622 12210
rect 30052 12210 30640 12226
rect 30052 12193 30068 12210
rect 29606 12176 29808 12193
rect 28848 12138 29808 12176
rect 29866 12176 30068 12193
rect 30624 12193 30640 12210
rect 31070 12210 31658 12226
rect 31070 12193 31086 12210
rect 30624 12176 30826 12193
rect 29866 12138 30826 12176
rect 30884 12176 31086 12193
rect 31642 12193 31658 12210
rect 32088 12210 32676 12226
rect 32088 12193 32104 12210
rect 31642 12176 31844 12193
rect 30884 12138 31844 12176
rect 31902 12176 32104 12193
rect 32660 12193 32676 12210
rect 33106 12210 33694 12226
rect 33106 12193 33122 12210
rect 32660 12176 32862 12193
rect 31902 12138 32862 12176
rect 32920 12176 33122 12193
rect 33678 12193 33694 12210
rect 33678 12176 33880 12193
rect 32920 12138 33880 12176
rect 1812 11584 2772 11622
rect 1812 11567 2014 11584
rect 1998 11550 2014 11567
rect 2570 11567 2772 11584
rect 2830 11584 3790 11622
rect 2830 11567 3032 11584
rect 2570 11550 2586 11567
rect 1998 11534 2586 11550
rect 3016 11550 3032 11567
rect 3588 11567 3790 11584
rect 3848 11584 4808 11622
rect 3848 11567 4050 11584
rect 3588 11550 3604 11567
rect 3016 11534 3604 11550
rect 1998 11476 2586 11492
rect 1998 11459 2014 11476
rect 1812 11442 2014 11459
rect 2570 11459 2586 11476
rect 4034 11550 4050 11567
rect 4606 11567 4808 11584
rect 4866 11584 5826 11622
rect 4866 11567 5068 11584
rect 4606 11550 4622 11567
rect 4034 11534 4622 11550
rect 3016 11476 3604 11492
rect 3016 11459 3032 11476
rect 2570 11442 2772 11459
rect 1812 11404 2772 11442
rect 2830 11442 3032 11459
rect 3588 11459 3604 11476
rect 5052 11550 5068 11567
rect 5624 11567 5826 11584
rect 5884 11584 6844 11622
rect 5884 11567 6086 11584
rect 5624 11550 5640 11567
rect 5052 11534 5640 11550
rect 4034 11476 4622 11492
rect 4034 11459 4050 11476
rect 3588 11442 3790 11459
rect 2830 11404 3790 11442
rect 3848 11442 4050 11459
rect 4606 11459 4622 11476
rect 6070 11550 6086 11567
rect 6642 11567 6844 11584
rect 6902 11584 7862 11622
rect 6902 11567 7104 11584
rect 6642 11550 6658 11567
rect 6070 11534 6658 11550
rect 5052 11476 5640 11492
rect 5052 11459 5068 11476
rect 4606 11442 4808 11459
rect 3848 11404 4808 11442
rect 4866 11442 5068 11459
rect 5624 11459 5640 11476
rect 7088 11550 7104 11567
rect 7660 11567 7862 11584
rect 7920 11584 8880 11622
rect 7920 11567 8122 11584
rect 7660 11550 7676 11567
rect 7088 11534 7676 11550
rect 6070 11476 6658 11492
rect 6070 11459 6086 11476
rect 5624 11442 5826 11459
rect 4866 11404 5826 11442
rect 5884 11442 6086 11459
rect 6642 11459 6658 11476
rect 8106 11550 8122 11567
rect 8678 11567 8880 11584
rect 8938 11584 9898 11622
rect 8938 11567 9140 11584
rect 8678 11550 8694 11567
rect 8106 11534 8694 11550
rect 7088 11476 7676 11492
rect 7088 11459 7104 11476
rect 6642 11442 6844 11459
rect 5884 11404 6844 11442
rect 6902 11442 7104 11459
rect 7660 11459 7676 11476
rect 9124 11550 9140 11567
rect 9696 11567 9898 11584
rect 9956 11584 10916 11622
rect 9956 11567 10158 11584
rect 9696 11550 9712 11567
rect 9124 11534 9712 11550
rect 8106 11476 8694 11492
rect 8106 11459 8122 11476
rect 7660 11442 7862 11459
rect 6902 11404 7862 11442
rect 7920 11442 8122 11459
rect 8678 11459 8694 11476
rect 10142 11550 10158 11567
rect 10714 11567 10916 11584
rect 10714 11550 10730 11567
rect 10142 11534 10730 11550
rect 9124 11476 9712 11492
rect 9124 11459 9140 11476
rect 8678 11442 8880 11459
rect 7920 11404 8880 11442
rect 8938 11442 9140 11459
rect 9696 11459 9712 11476
rect 10142 11476 10730 11492
rect 10142 11459 10158 11476
rect 9696 11442 9898 11459
rect 8938 11404 9898 11442
rect 9956 11442 10158 11459
rect 10714 11459 10730 11476
rect 13578 11500 14538 11538
rect 13578 11483 13780 11500
rect 13764 11466 13780 11483
rect 14336 11483 14538 11500
rect 14596 11500 15556 11538
rect 14596 11483 14798 11500
rect 14336 11466 14352 11483
rect 10714 11442 10916 11459
rect 13764 11450 14352 11466
rect 14782 11466 14798 11483
rect 15354 11483 15556 11500
rect 15614 11500 16574 11538
rect 15614 11483 15816 11500
rect 15354 11466 15370 11483
rect 14782 11450 15370 11466
rect 15800 11466 15816 11483
rect 16372 11483 16574 11500
rect 16632 11500 17592 11538
rect 16632 11483 16834 11500
rect 16372 11466 16388 11483
rect 15800 11450 16388 11466
rect 16818 11466 16834 11483
rect 17390 11483 17592 11500
rect 17650 11500 18610 11538
rect 17650 11483 17852 11500
rect 17390 11466 17406 11483
rect 16818 11450 17406 11466
rect 17836 11466 17852 11483
rect 18408 11483 18610 11500
rect 18668 11500 19628 11538
rect 18668 11483 18870 11500
rect 18408 11466 18424 11483
rect 17836 11450 18424 11466
rect 18854 11466 18870 11483
rect 19426 11483 19628 11500
rect 19686 11500 20646 11538
rect 19686 11483 19888 11500
rect 19426 11466 19442 11483
rect 18854 11450 19442 11466
rect 19872 11466 19888 11483
rect 20444 11483 20646 11500
rect 20704 11500 21664 11538
rect 20704 11483 20906 11500
rect 20444 11466 20460 11483
rect 19872 11450 20460 11466
rect 20890 11466 20906 11483
rect 21462 11483 21664 11500
rect 21722 11500 22682 11538
rect 21722 11483 21924 11500
rect 21462 11466 21478 11483
rect 20890 11450 21478 11466
rect 21908 11466 21924 11483
rect 22480 11483 22682 11500
rect 22740 11500 23700 11538
rect 22740 11483 22942 11500
rect 22480 11466 22496 11483
rect 21908 11450 22496 11466
rect 22926 11466 22942 11483
rect 23498 11483 23700 11500
rect 23758 11500 24718 11538
rect 23758 11483 23960 11500
rect 23498 11466 23514 11483
rect 22926 11450 23514 11466
rect 23944 11466 23960 11483
rect 24516 11483 24718 11500
rect 24776 11500 25736 11538
rect 24776 11483 24978 11500
rect 24516 11466 24532 11483
rect 23944 11450 24532 11466
rect 24962 11466 24978 11483
rect 25534 11483 25736 11500
rect 25794 11500 26754 11538
rect 25794 11483 25996 11500
rect 25534 11466 25550 11483
rect 24962 11450 25550 11466
rect 25980 11466 25996 11483
rect 26552 11483 26754 11500
rect 26812 11500 27772 11538
rect 26812 11483 27014 11500
rect 26552 11466 26568 11483
rect 25980 11450 26568 11466
rect 26998 11466 27014 11483
rect 27570 11483 27772 11500
rect 27830 11500 28790 11538
rect 27830 11483 28032 11500
rect 27570 11466 27586 11483
rect 26998 11450 27586 11466
rect 28016 11466 28032 11483
rect 28588 11483 28790 11500
rect 28848 11500 29808 11538
rect 28848 11483 29050 11500
rect 28588 11466 28604 11483
rect 28016 11450 28604 11466
rect 29034 11466 29050 11483
rect 29606 11483 29808 11500
rect 29866 11500 30826 11538
rect 29866 11483 30068 11500
rect 29606 11466 29622 11483
rect 29034 11450 29622 11466
rect 30052 11466 30068 11483
rect 30624 11483 30826 11500
rect 30884 11500 31844 11538
rect 30884 11483 31086 11500
rect 30624 11466 30640 11483
rect 30052 11450 30640 11466
rect 31070 11466 31086 11483
rect 31642 11483 31844 11500
rect 31902 11500 32862 11538
rect 31902 11483 32104 11500
rect 31642 11466 31658 11483
rect 31070 11450 31658 11466
rect 32088 11466 32104 11483
rect 32660 11483 32862 11500
rect 32920 11500 33880 11538
rect 32920 11483 33122 11500
rect 32660 11466 32676 11483
rect 32088 11450 32676 11466
rect 33106 11466 33122 11483
rect 33678 11483 33880 11500
rect 33678 11466 33694 11483
rect 33106 11450 33694 11466
rect 9956 11404 10916 11442
rect 13764 10978 14352 10994
rect 13764 10961 13780 10978
rect 13578 10944 13780 10961
rect 14336 10961 14352 10978
rect 14782 10978 15370 10994
rect 14782 10961 14798 10978
rect 14336 10944 14538 10961
rect 13578 10906 14538 10944
rect 14596 10944 14798 10961
rect 15354 10961 15370 10978
rect 15800 10978 16388 10994
rect 15800 10961 15816 10978
rect 15354 10944 15556 10961
rect 14596 10906 15556 10944
rect 15614 10944 15816 10961
rect 16372 10961 16388 10978
rect 16818 10978 17406 10994
rect 16818 10961 16834 10978
rect 16372 10944 16574 10961
rect 15614 10906 16574 10944
rect 16632 10944 16834 10961
rect 17390 10961 17406 10978
rect 17836 10978 18424 10994
rect 17836 10961 17852 10978
rect 17390 10944 17592 10961
rect 16632 10906 17592 10944
rect 17650 10944 17852 10961
rect 18408 10961 18424 10978
rect 18854 10978 19442 10994
rect 18854 10961 18870 10978
rect 18408 10944 18610 10961
rect 17650 10906 18610 10944
rect 18668 10944 18870 10961
rect 19426 10961 19442 10978
rect 19872 10978 20460 10994
rect 19872 10961 19888 10978
rect 19426 10944 19628 10961
rect 18668 10906 19628 10944
rect 19686 10944 19888 10961
rect 20444 10961 20460 10978
rect 20890 10978 21478 10994
rect 20890 10961 20906 10978
rect 20444 10944 20646 10961
rect 19686 10906 20646 10944
rect 20704 10944 20906 10961
rect 21462 10961 21478 10978
rect 21908 10978 22496 10994
rect 21908 10961 21924 10978
rect 21462 10944 21664 10961
rect 20704 10906 21664 10944
rect 21722 10944 21924 10961
rect 22480 10961 22496 10978
rect 22926 10978 23514 10994
rect 22926 10961 22942 10978
rect 22480 10944 22682 10961
rect 21722 10906 22682 10944
rect 22740 10944 22942 10961
rect 23498 10961 23514 10978
rect 23944 10978 24532 10994
rect 23944 10961 23960 10978
rect 23498 10944 23700 10961
rect 22740 10906 23700 10944
rect 23758 10944 23960 10961
rect 24516 10961 24532 10978
rect 24962 10978 25550 10994
rect 24962 10961 24978 10978
rect 24516 10944 24718 10961
rect 23758 10906 24718 10944
rect 24776 10944 24978 10961
rect 25534 10961 25550 10978
rect 25980 10978 26568 10994
rect 25980 10961 25996 10978
rect 25534 10944 25736 10961
rect 24776 10906 25736 10944
rect 25794 10944 25996 10961
rect 26552 10961 26568 10978
rect 26998 10978 27586 10994
rect 26998 10961 27014 10978
rect 26552 10944 26754 10961
rect 25794 10906 26754 10944
rect 26812 10944 27014 10961
rect 27570 10961 27586 10978
rect 28016 10978 28604 10994
rect 28016 10961 28032 10978
rect 27570 10944 27772 10961
rect 26812 10906 27772 10944
rect 27830 10944 28032 10961
rect 28588 10961 28604 10978
rect 29034 10978 29622 10994
rect 29034 10961 29050 10978
rect 28588 10944 28790 10961
rect 27830 10906 28790 10944
rect 28848 10944 29050 10961
rect 29606 10961 29622 10978
rect 30052 10978 30640 10994
rect 30052 10961 30068 10978
rect 29606 10944 29808 10961
rect 28848 10906 29808 10944
rect 29866 10944 30068 10961
rect 30624 10961 30640 10978
rect 31070 10978 31658 10994
rect 31070 10961 31086 10978
rect 30624 10944 30826 10961
rect 29866 10906 30826 10944
rect 30884 10944 31086 10961
rect 31642 10961 31658 10978
rect 32088 10978 32676 10994
rect 32088 10961 32104 10978
rect 31642 10944 31844 10961
rect 30884 10906 31844 10944
rect 31902 10944 32104 10961
rect 32660 10961 32676 10978
rect 33106 10978 33694 10994
rect 33106 10961 33122 10978
rect 32660 10944 32862 10961
rect 31902 10906 32862 10944
rect 32920 10944 33122 10961
rect 33678 10961 33694 10978
rect 33678 10944 33880 10961
rect 32920 10906 33880 10944
rect 1812 10766 2772 10804
rect 1812 10749 2014 10766
rect 1998 10732 2014 10749
rect 2570 10749 2772 10766
rect 2830 10766 3790 10804
rect 2830 10749 3032 10766
rect 2570 10732 2586 10749
rect 1998 10716 2586 10732
rect 3016 10732 3032 10749
rect 3588 10749 3790 10766
rect 3848 10766 4808 10804
rect 3848 10749 4050 10766
rect 3588 10732 3604 10749
rect 3016 10716 3604 10732
rect 1998 10658 2586 10674
rect 1998 10641 2014 10658
rect 1812 10624 2014 10641
rect 2570 10641 2586 10658
rect 4034 10732 4050 10749
rect 4606 10749 4808 10766
rect 4866 10766 5826 10804
rect 4866 10749 5068 10766
rect 4606 10732 4622 10749
rect 4034 10716 4622 10732
rect 3016 10658 3604 10674
rect 3016 10641 3032 10658
rect 2570 10624 2772 10641
rect 1812 10586 2772 10624
rect 2830 10624 3032 10641
rect 3588 10641 3604 10658
rect 5052 10732 5068 10749
rect 5624 10749 5826 10766
rect 5884 10766 6844 10804
rect 5884 10749 6086 10766
rect 5624 10732 5640 10749
rect 5052 10716 5640 10732
rect 4034 10658 4622 10674
rect 4034 10641 4050 10658
rect 3588 10624 3790 10641
rect 2830 10586 3790 10624
rect 3848 10624 4050 10641
rect 4606 10641 4622 10658
rect 6070 10732 6086 10749
rect 6642 10749 6844 10766
rect 6902 10766 7862 10804
rect 6902 10749 7104 10766
rect 6642 10732 6658 10749
rect 6070 10716 6658 10732
rect 5052 10658 5640 10674
rect 5052 10641 5068 10658
rect 4606 10624 4808 10641
rect 3848 10586 4808 10624
rect 4866 10624 5068 10641
rect 5624 10641 5640 10658
rect 7088 10732 7104 10749
rect 7660 10749 7862 10766
rect 7920 10766 8880 10804
rect 7920 10749 8122 10766
rect 7660 10732 7676 10749
rect 7088 10716 7676 10732
rect 6070 10658 6658 10674
rect 6070 10641 6086 10658
rect 5624 10624 5826 10641
rect 4866 10586 5826 10624
rect 5884 10624 6086 10641
rect 6642 10641 6658 10658
rect 8106 10732 8122 10749
rect 8678 10749 8880 10766
rect 8938 10766 9898 10804
rect 8938 10749 9140 10766
rect 8678 10732 8694 10749
rect 8106 10716 8694 10732
rect 7088 10658 7676 10674
rect 7088 10641 7104 10658
rect 6642 10624 6844 10641
rect 5884 10586 6844 10624
rect 6902 10624 7104 10641
rect 7660 10641 7676 10658
rect 9124 10732 9140 10749
rect 9696 10749 9898 10766
rect 9956 10766 10916 10804
rect 9956 10749 10158 10766
rect 9696 10732 9712 10749
rect 9124 10716 9712 10732
rect 8106 10658 8694 10674
rect 8106 10641 8122 10658
rect 7660 10624 7862 10641
rect 6902 10586 7862 10624
rect 7920 10624 8122 10641
rect 8678 10641 8694 10658
rect 10142 10732 10158 10749
rect 10714 10749 10916 10766
rect 10714 10732 10730 10749
rect 10142 10716 10730 10732
rect 9124 10658 9712 10674
rect 9124 10641 9140 10658
rect 8678 10624 8880 10641
rect 7920 10586 8880 10624
rect 8938 10624 9140 10641
rect 9696 10641 9712 10658
rect 10142 10658 10730 10674
rect 10142 10641 10158 10658
rect 9696 10624 9898 10641
rect 8938 10586 9898 10624
rect 9956 10624 10158 10641
rect 10714 10641 10730 10658
rect 10714 10624 10916 10641
rect 9956 10586 10916 10624
rect 13578 10268 14538 10306
rect 13578 10251 13780 10268
rect 13764 10234 13780 10251
rect 14336 10251 14538 10268
rect 14596 10268 15556 10306
rect 14596 10251 14798 10268
rect 14336 10234 14352 10251
rect 13764 10218 14352 10234
rect 14782 10234 14798 10251
rect 15354 10251 15556 10268
rect 15614 10268 16574 10306
rect 15614 10251 15816 10268
rect 15354 10234 15370 10251
rect 14782 10218 15370 10234
rect 15800 10234 15816 10251
rect 16372 10251 16574 10268
rect 16632 10268 17592 10306
rect 16632 10251 16834 10268
rect 16372 10234 16388 10251
rect 15800 10218 16388 10234
rect 16818 10234 16834 10251
rect 17390 10251 17592 10268
rect 17650 10268 18610 10306
rect 17650 10251 17852 10268
rect 17390 10234 17406 10251
rect 16818 10218 17406 10234
rect 17836 10234 17852 10251
rect 18408 10251 18610 10268
rect 18668 10268 19628 10306
rect 18668 10251 18870 10268
rect 18408 10234 18424 10251
rect 17836 10218 18424 10234
rect 18854 10234 18870 10251
rect 19426 10251 19628 10268
rect 19686 10268 20646 10306
rect 19686 10251 19888 10268
rect 19426 10234 19442 10251
rect 18854 10218 19442 10234
rect 19872 10234 19888 10251
rect 20444 10251 20646 10268
rect 20704 10268 21664 10306
rect 20704 10251 20906 10268
rect 20444 10234 20460 10251
rect 19872 10218 20460 10234
rect 20890 10234 20906 10251
rect 21462 10251 21664 10268
rect 21722 10268 22682 10306
rect 21722 10251 21924 10268
rect 21462 10234 21478 10251
rect 20890 10218 21478 10234
rect 21908 10234 21924 10251
rect 22480 10251 22682 10268
rect 22740 10268 23700 10306
rect 22740 10251 22942 10268
rect 22480 10234 22496 10251
rect 21908 10218 22496 10234
rect 22926 10234 22942 10251
rect 23498 10251 23700 10268
rect 23758 10268 24718 10306
rect 23758 10251 23960 10268
rect 23498 10234 23514 10251
rect 22926 10218 23514 10234
rect 23944 10234 23960 10251
rect 24516 10251 24718 10268
rect 24776 10268 25736 10306
rect 24776 10251 24978 10268
rect 24516 10234 24532 10251
rect 23944 10218 24532 10234
rect 24962 10234 24978 10251
rect 25534 10251 25736 10268
rect 25794 10268 26754 10306
rect 25794 10251 25996 10268
rect 25534 10234 25550 10251
rect 24962 10218 25550 10234
rect 25980 10234 25996 10251
rect 26552 10251 26754 10268
rect 26812 10268 27772 10306
rect 26812 10251 27014 10268
rect 26552 10234 26568 10251
rect 25980 10218 26568 10234
rect 26998 10234 27014 10251
rect 27570 10251 27772 10268
rect 27830 10268 28790 10306
rect 27830 10251 28032 10268
rect 27570 10234 27586 10251
rect 26998 10218 27586 10234
rect 28016 10234 28032 10251
rect 28588 10251 28790 10268
rect 28848 10268 29808 10306
rect 28848 10251 29050 10268
rect 28588 10234 28604 10251
rect 28016 10218 28604 10234
rect 29034 10234 29050 10251
rect 29606 10251 29808 10268
rect 29866 10268 30826 10306
rect 29866 10251 30068 10268
rect 29606 10234 29622 10251
rect 29034 10218 29622 10234
rect 30052 10234 30068 10251
rect 30624 10251 30826 10268
rect 30884 10268 31844 10306
rect 30884 10251 31086 10268
rect 30624 10234 30640 10251
rect 30052 10218 30640 10234
rect 31070 10234 31086 10251
rect 31642 10251 31844 10268
rect 31902 10268 32862 10306
rect 31902 10251 32104 10268
rect 31642 10234 31658 10251
rect 31070 10218 31658 10234
rect 32088 10234 32104 10251
rect 32660 10251 32862 10268
rect 32920 10268 33880 10306
rect 32920 10251 33122 10268
rect 32660 10234 32676 10251
rect 32088 10218 32676 10234
rect 33106 10234 33122 10251
rect 33678 10251 33880 10268
rect 33678 10234 33694 10251
rect 33106 10218 33694 10234
rect 1812 9948 2772 9986
rect 1812 9931 2014 9948
rect 1998 9914 2014 9931
rect 2570 9931 2772 9948
rect 2830 9948 3790 9986
rect 2830 9931 3032 9948
rect 2570 9914 2586 9931
rect 1998 9898 2586 9914
rect 3016 9914 3032 9931
rect 3588 9931 3790 9948
rect 3848 9948 4808 9986
rect 3848 9931 4050 9948
rect 3588 9914 3604 9931
rect 3016 9898 3604 9914
rect 1998 9840 2586 9856
rect 1998 9823 2014 9840
rect 1812 9806 2014 9823
rect 2570 9823 2586 9840
rect 4034 9914 4050 9931
rect 4606 9931 4808 9948
rect 4866 9948 5826 9986
rect 4866 9931 5068 9948
rect 4606 9914 4622 9931
rect 4034 9898 4622 9914
rect 3016 9840 3604 9856
rect 3016 9823 3032 9840
rect 2570 9806 2772 9823
rect 1812 9768 2772 9806
rect 2830 9806 3032 9823
rect 3588 9823 3604 9840
rect 5052 9914 5068 9931
rect 5624 9931 5826 9948
rect 5884 9948 6844 9986
rect 5884 9931 6086 9948
rect 5624 9914 5640 9931
rect 5052 9898 5640 9914
rect 4034 9840 4622 9856
rect 4034 9823 4050 9840
rect 3588 9806 3790 9823
rect 2830 9768 3790 9806
rect 3848 9806 4050 9823
rect 4606 9823 4622 9840
rect 6070 9914 6086 9931
rect 6642 9931 6844 9948
rect 6902 9948 7862 9986
rect 6902 9931 7104 9948
rect 6642 9914 6658 9931
rect 6070 9898 6658 9914
rect 5052 9840 5640 9856
rect 5052 9823 5068 9840
rect 4606 9806 4808 9823
rect 3848 9768 4808 9806
rect 4866 9806 5068 9823
rect 5624 9823 5640 9840
rect 7088 9914 7104 9931
rect 7660 9931 7862 9948
rect 7920 9948 8880 9986
rect 7920 9931 8122 9948
rect 7660 9914 7676 9931
rect 7088 9898 7676 9914
rect 6070 9840 6658 9856
rect 6070 9823 6086 9840
rect 5624 9806 5826 9823
rect 4866 9768 5826 9806
rect 5884 9806 6086 9823
rect 6642 9823 6658 9840
rect 8106 9914 8122 9931
rect 8678 9931 8880 9948
rect 8938 9948 9898 9986
rect 8938 9931 9140 9948
rect 8678 9914 8694 9931
rect 8106 9898 8694 9914
rect 7088 9840 7676 9856
rect 7088 9823 7104 9840
rect 6642 9806 6844 9823
rect 5884 9768 6844 9806
rect 6902 9806 7104 9823
rect 7660 9823 7676 9840
rect 9124 9914 9140 9931
rect 9696 9931 9898 9948
rect 9956 9948 10916 9986
rect 9956 9931 10158 9948
rect 9696 9914 9712 9931
rect 9124 9898 9712 9914
rect 8106 9840 8694 9856
rect 8106 9823 8122 9840
rect 7660 9806 7862 9823
rect 6902 9768 7862 9806
rect 7920 9806 8122 9823
rect 8678 9823 8694 9840
rect 10142 9914 10158 9931
rect 10714 9931 10916 9948
rect 10714 9914 10730 9931
rect 10142 9898 10730 9914
rect 9124 9840 9712 9856
rect 9124 9823 9140 9840
rect 8678 9806 8880 9823
rect 7920 9768 8880 9806
rect 8938 9806 9140 9823
rect 9696 9823 9712 9840
rect 10142 9840 10730 9856
rect 10142 9823 10158 9840
rect 9696 9806 9898 9823
rect 8938 9768 9898 9806
rect 9956 9806 10158 9823
rect 10714 9823 10730 9840
rect 10714 9806 10916 9823
rect 9956 9768 10916 9806
rect 13762 9744 14350 9760
rect 13762 9727 13778 9744
rect 13576 9710 13778 9727
rect 14334 9727 14350 9744
rect 14780 9744 15368 9760
rect 14780 9727 14796 9744
rect 14334 9710 14536 9727
rect 13576 9672 14536 9710
rect 14594 9710 14796 9727
rect 15352 9727 15368 9744
rect 15798 9744 16386 9760
rect 15798 9727 15814 9744
rect 15352 9710 15554 9727
rect 14594 9672 15554 9710
rect 15612 9710 15814 9727
rect 16370 9727 16386 9744
rect 16816 9744 17404 9760
rect 16816 9727 16832 9744
rect 16370 9710 16572 9727
rect 15612 9672 16572 9710
rect 16630 9710 16832 9727
rect 17388 9727 17404 9744
rect 17834 9744 18422 9760
rect 17834 9727 17850 9744
rect 17388 9710 17590 9727
rect 16630 9672 17590 9710
rect 17648 9710 17850 9727
rect 18406 9727 18422 9744
rect 18852 9744 19440 9760
rect 18852 9727 18868 9744
rect 18406 9710 18608 9727
rect 17648 9672 18608 9710
rect 18666 9710 18868 9727
rect 19424 9727 19440 9744
rect 19870 9744 20458 9760
rect 19870 9727 19886 9744
rect 19424 9710 19626 9727
rect 18666 9672 19626 9710
rect 19684 9710 19886 9727
rect 20442 9727 20458 9744
rect 20888 9744 21476 9760
rect 20888 9727 20904 9744
rect 20442 9710 20644 9727
rect 19684 9672 20644 9710
rect 20702 9710 20904 9727
rect 21460 9727 21476 9744
rect 21906 9744 22494 9760
rect 21906 9727 21922 9744
rect 21460 9710 21662 9727
rect 20702 9672 21662 9710
rect 21720 9710 21922 9727
rect 22478 9727 22494 9744
rect 22924 9744 23512 9760
rect 22924 9727 22940 9744
rect 22478 9710 22680 9727
rect 21720 9672 22680 9710
rect 22738 9710 22940 9727
rect 23496 9727 23512 9744
rect 23942 9744 24530 9760
rect 23942 9727 23958 9744
rect 23496 9710 23698 9727
rect 22738 9672 23698 9710
rect 23756 9710 23958 9727
rect 24514 9727 24530 9744
rect 24960 9744 25548 9760
rect 24960 9727 24976 9744
rect 24514 9710 24716 9727
rect 23756 9672 24716 9710
rect 24774 9710 24976 9727
rect 25532 9727 25548 9744
rect 25978 9744 26566 9760
rect 25978 9727 25994 9744
rect 25532 9710 25734 9727
rect 24774 9672 25734 9710
rect 25792 9710 25994 9727
rect 26550 9727 26566 9744
rect 26996 9744 27584 9760
rect 26996 9727 27012 9744
rect 26550 9710 26752 9727
rect 25792 9672 26752 9710
rect 26810 9710 27012 9727
rect 27568 9727 27584 9744
rect 28014 9744 28602 9760
rect 28014 9727 28030 9744
rect 27568 9710 27770 9727
rect 26810 9672 27770 9710
rect 27828 9710 28030 9727
rect 28586 9727 28602 9744
rect 29032 9744 29620 9760
rect 29032 9727 29048 9744
rect 28586 9710 28788 9727
rect 27828 9672 28788 9710
rect 28846 9710 29048 9727
rect 29604 9727 29620 9744
rect 30050 9744 30638 9760
rect 30050 9727 30066 9744
rect 29604 9710 29806 9727
rect 28846 9672 29806 9710
rect 29864 9710 30066 9727
rect 30622 9727 30638 9744
rect 31068 9744 31656 9760
rect 31068 9727 31084 9744
rect 30622 9710 30824 9727
rect 29864 9672 30824 9710
rect 30882 9710 31084 9727
rect 31640 9727 31656 9744
rect 32086 9744 32674 9760
rect 32086 9727 32102 9744
rect 31640 9710 31842 9727
rect 30882 9672 31842 9710
rect 31900 9710 32102 9727
rect 32658 9727 32674 9744
rect 33104 9744 33692 9760
rect 33104 9727 33120 9744
rect 32658 9710 32860 9727
rect 31900 9672 32860 9710
rect 32918 9710 33120 9727
rect 33676 9727 33692 9744
rect 33676 9710 33878 9727
rect 32918 9672 33878 9710
rect 1812 9130 2772 9168
rect 1812 9113 2014 9130
rect 1998 9096 2014 9113
rect 2570 9113 2772 9130
rect 2830 9130 3790 9168
rect 2830 9113 3032 9130
rect 2570 9096 2586 9113
rect 1998 9080 2586 9096
rect 3016 9096 3032 9113
rect 3588 9113 3790 9130
rect 3848 9130 4808 9168
rect 3848 9113 4050 9130
rect 3588 9096 3604 9113
rect 3016 9080 3604 9096
rect 1998 9022 2586 9038
rect 1998 9005 2014 9022
rect 1812 8988 2014 9005
rect 2570 9005 2586 9022
rect 4034 9096 4050 9113
rect 4606 9113 4808 9130
rect 4866 9130 5826 9168
rect 4866 9113 5068 9130
rect 4606 9096 4622 9113
rect 4034 9080 4622 9096
rect 3016 9022 3604 9038
rect 3016 9005 3032 9022
rect 2570 8988 2772 9005
rect 1812 8950 2772 8988
rect 2830 8988 3032 9005
rect 3588 9005 3604 9022
rect 5052 9096 5068 9113
rect 5624 9113 5826 9130
rect 5884 9130 6844 9168
rect 5884 9113 6086 9130
rect 5624 9096 5640 9113
rect 5052 9080 5640 9096
rect 4034 9022 4622 9038
rect 4034 9005 4050 9022
rect 3588 8988 3790 9005
rect 2830 8950 3790 8988
rect 3848 8988 4050 9005
rect 4606 9005 4622 9022
rect 6070 9096 6086 9113
rect 6642 9113 6844 9130
rect 6902 9130 7862 9168
rect 6902 9113 7104 9130
rect 6642 9096 6658 9113
rect 6070 9080 6658 9096
rect 5052 9022 5640 9038
rect 5052 9005 5068 9022
rect 4606 8988 4808 9005
rect 3848 8950 4808 8988
rect 4866 8988 5068 9005
rect 5624 9005 5640 9022
rect 7088 9096 7104 9113
rect 7660 9113 7862 9130
rect 7920 9130 8880 9168
rect 7920 9113 8122 9130
rect 7660 9096 7676 9113
rect 7088 9080 7676 9096
rect 6070 9022 6658 9038
rect 6070 9005 6086 9022
rect 5624 8988 5826 9005
rect 4866 8950 5826 8988
rect 5884 8988 6086 9005
rect 6642 9005 6658 9022
rect 8106 9096 8122 9113
rect 8678 9113 8880 9130
rect 8938 9130 9898 9168
rect 8938 9113 9140 9130
rect 8678 9096 8694 9113
rect 8106 9080 8694 9096
rect 7088 9022 7676 9038
rect 7088 9005 7104 9022
rect 6642 8988 6844 9005
rect 5884 8950 6844 8988
rect 6902 8988 7104 9005
rect 7660 9005 7676 9022
rect 9124 9096 9140 9113
rect 9696 9113 9898 9130
rect 9956 9130 10916 9168
rect 9956 9113 10158 9130
rect 9696 9096 9712 9113
rect 9124 9080 9712 9096
rect 8106 9022 8694 9038
rect 8106 9005 8122 9022
rect 7660 8988 7862 9005
rect 6902 8950 7862 8988
rect 7920 8988 8122 9005
rect 8678 9005 8694 9022
rect 10142 9096 10158 9113
rect 10714 9113 10916 9130
rect 10714 9096 10730 9113
rect 10142 9080 10730 9096
rect 9124 9022 9712 9038
rect 9124 9005 9140 9022
rect 8678 8988 8880 9005
rect 7920 8950 8880 8988
rect 8938 8988 9140 9005
rect 9696 9005 9712 9022
rect 10142 9022 10730 9038
rect 10142 9005 10158 9022
rect 9696 8988 9898 9005
rect 8938 8950 9898 8988
rect 9956 8988 10158 9005
rect 10714 9005 10730 9022
rect 13576 9034 14536 9072
rect 13576 9017 13778 9034
rect 10714 8988 10916 9005
rect 9956 8950 10916 8988
rect 13762 9000 13778 9017
rect 14334 9017 14536 9034
rect 14594 9034 15554 9072
rect 14594 9017 14796 9034
rect 14334 9000 14350 9017
rect 13762 8984 14350 9000
rect 14780 9000 14796 9017
rect 15352 9017 15554 9034
rect 15612 9034 16572 9072
rect 15612 9017 15814 9034
rect 15352 9000 15368 9017
rect 14780 8984 15368 9000
rect 15798 9000 15814 9017
rect 16370 9017 16572 9034
rect 16630 9034 17590 9072
rect 16630 9017 16832 9034
rect 16370 9000 16386 9017
rect 15798 8984 16386 9000
rect 16816 9000 16832 9017
rect 17388 9017 17590 9034
rect 17648 9034 18608 9072
rect 17648 9017 17850 9034
rect 17388 9000 17404 9017
rect 16816 8984 17404 9000
rect 17834 9000 17850 9017
rect 18406 9017 18608 9034
rect 18666 9034 19626 9072
rect 18666 9017 18868 9034
rect 18406 9000 18422 9017
rect 17834 8984 18422 9000
rect 18852 9000 18868 9017
rect 19424 9017 19626 9034
rect 19684 9034 20644 9072
rect 19684 9017 19886 9034
rect 19424 9000 19440 9017
rect 18852 8984 19440 9000
rect 19870 9000 19886 9017
rect 20442 9017 20644 9034
rect 20702 9034 21662 9072
rect 20702 9017 20904 9034
rect 20442 9000 20458 9017
rect 19870 8984 20458 9000
rect 20888 9000 20904 9017
rect 21460 9017 21662 9034
rect 21720 9034 22680 9072
rect 21720 9017 21922 9034
rect 21460 9000 21476 9017
rect 20888 8984 21476 9000
rect 21906 9000 21922 9017
rect 22478 9017 22680 9034
rect 22738 9034 23698 9072
rect 22738 9017 22940 9034
rect 22478 9000 22494 9017
rect 21906 8984 22494 9000
rect 22924 9000 22940 9017
rect 23496 9017 23698 9034
rect 23756 9034 24716 9072
rect 23756 9017 23958 9034
rect 23496 9000 23512 9017
rect 22924 8984 23512 9000
rect 23942 9000 23958 9017
rect 24514 9017 24716 9034
rect 24774 9034 25734 9072
rect 24774 9017 24976 9034
rect 24514 9000 24530 9017
rect 23942 8984 24530 9000
rect 24960 9000 24976 9017
rect 25532 9017 25734 9034
rect 25792 9034 26752 9072
rect 25792 9017 25994 9034
rect 25532 9000 25548 9017
rect 24960 8984 25548 9000
rect 25978 9000 25994 9017
rect 26550 9017 26752 9034
rect 26810 9034 27770 9072
rect 26810 9017 27012 9034
rect 26550 9000 26566 9017
rect 25978 8984 26566 9000
rect 26996 9000 27012 9017
rect 27568 9017 27770 9034
rect 27828 9034 28788 9072
rect 27828 9017 28030 9034
rect 27568 9000 27584 9017
rect 26996 8984 27584 9000
rect 28014 9000 28030 9017
rect 28586 9017 28788 9034
rect 28846 9034 29806 9072
rect 28846 9017 29048 9034
rect 28586 9000 28602 9017
rect 28014 8984 28602 9000
rect 29032 9000 29048 9017
rect 29604 9017 29806 9034
rect 29864 9034 30824 9072
rect 29864 9017 30066 9034
rect 29604 9000 29620 9017
rect 29032 8984 29620 9000
rect 30050 9000 30066 9017
rect 30622 9017 30824 9034
rect 30882 9034 31842 9072
rect 30882 9017 31084 9034
rect 30622 9000 30638 9017
rect 30050 8984 30638 9000
rect 31068 9000 31084 9017
rect 31640 9017 31842 9034
rect 31900 9034 32860 9072
rect 31900 9017 32102 9034
rect 31640 9000 31656 9017
rect 31068 8984 31656 9000
rect 32086 9000 32102 9017
rect 32658 9017 32860 9034
rect 32918 9034 33878 9072
rect 32918 9017 33120 9034
rect 32658 9000 32674 9017
rect 32086 8984 32674 9000
rect 33104 9000 33120 9017
rect 33676 9017 33878 9034
rect 33676 9000 33692 9017
rect 33104 8984 33692 9000
rect 13762 8510 14350 8526
rect 13762 8493 13778 8510
rect 13576 8476 13778 8493
rect 14334 8493 14350 8510
rect 14780 8510 15368 8526
rect 14780 8493 14796 8510
rect 14334 8476 14536 8493
rect 13576 8438 14536 8476
rect 14594 8476 14796 8493
rect 15352 8493 15368 8510
rect 15798 8510 16386 8526
rect 15798 8493 15814 8510
rect 15352 8476 15554 8493
rect 14594 8438 15554 8476
rect 15612 8476 15814 8493
rect 16370 8493 16386 8510
rect 16816 8510 17404 8526
rect 16816 8493 16832 8510
rect 16370 8476 16572 8493
rect 15612 8438 16572 8476
rect 16630 8476 16832 8493
rect 17388 8493 17404 8510
rect 17834 8510 18422 8526
rect 17834 8493 17850 8510
rect 17388 8476 17590 8493
rect 16630 8438 17590 8476
rect 17648 8476 17850 8493
rect 18406 8493 18422 8510
rect 18852 8510 19440 8526
rect 18852 8493 18868 8510
rect 18406 8476 18608 8493
rect 17648 8438 18608 8476
rect 18666 8476 18868 8493
rect 19424 8493 19440 8510
rect 19870 8510 20458 8526
rect 19870 8493 19886 8510
rect 19424 8476 19626 8493
rect 18666 8438 19626 8476
rect 19684 8476 19886 8493
rect 20442 8493 20458 8510
rect 20888 8510 21476 8526
rect 20888 8493 20904 8510
rect 20442 8476 20644 8493
rect 19684 8438 20644 8476
rect 20702 8476 20904 8493
rect 21460 8493 21476 8510
rect 21906 8510 22494 8526
rect 21906 8493 21922 8510
rect 21460 8476 21662 8493
rect 20702 8438 21662 8476
rect 21720 8476 21922 8493
rect 22478 8493 22494 8510
rect 22924 8510 23512 8526
rect 22924 8493 22940 8510
rect 22478 8476 22680 8493
rect 21720 8438 22680 8476
rect 22738 8476 22940 8493
rect 23496 8493 23512 8510
rect 23942 8510 24530 8526
rect 23942 8493 23958 8510
rect 23496 8476 23698 8493
rect 22738 8438 23698 8476
rect 23756 8476 23958 8493
rect 24514 8493 24530 8510
rect 24960 8510 25548 8526
rect 24960 8493 24976 8510
rect 24514 8476 24716 8493
rect 23756 8438 24716 8476
rect 24774 8476 24976 8493
rect 25532 8493 25548 8510
rect 25978 8510 26566 8526
rect 25978 8493 25994 8510
rect 25532 8476 25734 8493
rect 24774 8438 25734 8476
rect 25792 8476 25994 8493
rect 26550 8493 26566 8510
rect 26996 8510 27584 8526
rect 26996 8493 27012 8510
rect 26550 8476 26752 8493
rect 25792 8438 26752 8476
rect 26810 8476 27012 8493
rect 27568 8493 27584 8510
rect 28014 8510 28602 8526
rect 28014 8493 28030 8510
rect 27568 8476 27770 8493
rect 26810 8438 27770 8476
rect 27828 8476 28030 8493
rect 28586 8493 28602 8510
rect 29032 8510 29620 8526
rect 29032 8493 29048 8510
rect 28586 8476 28788 8493
rect 27828 8438 28788 8476
rect 28846 8476 29048 8493
rect 29604 8493 29620 8510
rect 30050 8510 30638 8526
rect 30050 8493 30066 8510
rect 29604 8476 29806 8493
rect 28846 8438 29806 8476
rect 29864 8476 30066 8493
rect 30622 8493 30638 8510
rect 31068 8510 31656 8526
rect 31068 8493 31084 8510
rect 30622 8476 30824 8493
rect 29864 8438 30824 8476
rect 30882 8476 31084 8493
rect 31640 8493 31656 8510
rect 32086 8510 32674 8526
rect 32086 8493 32102 8510
rect 31640 8476 31842 8493
rect 30882 8438 31842 8476
rect 31900 8476 32102 8493
rect 32658 8493 32674 8510
rect 33104 8510 33692 8526
rect 33104 8493 33120 8510
rect 32658 8476 32860 8493
rect 31900 8438 32860 8476
rect 32918 8476 33120 8493
rect 33676 8493 33692 8510
rect 33676 8476 33878 8493
rect 32918 8438 33878 8476
rect 1812 8312 2772 8350
rect 1812 8295 2014 8312
rect 1998 8278 2014 8295
rect 2570 8295 2772 8312
rect 2830 8312 3790 8350
rect 2830 8295 3032 8312
rect 2570 8278 2586 8295
rect 1998 8262 2586 8278
rect 3016 8278 3032 8295
rect 3588 8295 3790 8312
rect 3848 8312 4808 8350
rect 3848 8295 4050 8312
rect 3588 8278 3604 8295
rect 3016 8262 3604 8278
rect 1998 8204 2586 8220
rect 1998 8187 2014 8204
rect 1812 8170 2014 8187
rect 2570 8187 2586 8204
rect 4034 8278 4050 8295
rect 4606 8295 4808 8312
rect 4866 8312 5826 8350
rect 4866 8295 5068 8312
rect 4606 8278 4622 8295
rect 4034 8262 4622 8278
rect 3016 8204 3604 8220
rect 3016 8187 3032 8204
rect 2570 8170 2772 8187
rect 1812 8132 2772 8170
rect 2830 8170 3032 8187
rect 3588 8187 3604 8204
rect 5052 8278 5068 8295
rect 5624 8295 5826 8312
rect 5884 8312 6844 8350
rect 5884 8295 6086 8312
rect 5624 8278 5640 8295
rect 5052 8262 5640 8278
rect 4034 8204 4622 8220
rect 4034 8187 4050 8204
rect 3588 8170 3790 8187
rect 2830 8132 3790 8170
rect 3848 8170 4050 8187
rect 4606 8187 4622 8204
rect 6070 8278 6086 8295
rect 6642 8295 6844 8312
rect 6902 8312 7862 8350
rect 6902 8295 7104 8312
rect 6642 8278 6658 8295
rect 6070 8262 6658 8278
rect 5052 8204 5640 8220
rect 5052 8187 5068 8204
rect 4606 8170 4808 8187
rect 3848 8132 4808 8170
rect 4866 8170 5068 8187
rect 5624 8187 5640 8204
rect 7088 8278 7104 8295
rect 7660 8295 7862 8312
rect 7920 8312 8880 8350
rect 7920 8295 8122 8312
rect 7660 8278 7676 8295
rect 7088 8262 7676 8278
rect 6070 8204 6658 8220
rect 6070 8187 6086 8204
rect 5624 8170 5826 8187
rect 4866 8132 5826 8170
rect 5884 8170 6086 8187
rect 6642 8187 6658 8204
rect 8106 8278 8122 8295
rect 8678 8295 8880 8312
rect 8938 8312 9898 8350
rect 8938 8295 9140 8312
rect 8678 8278 8694 8295
rect 8106 8262 8694 8278
rect 7088 8204 7676 8220
rect 7088 8187 7104 8204
rect 6642 8170 6844 8187
rect 5884 8132 6844 8170
rect 6902 8170 7104 8187
rect 7660 8187 7676 8204
rect 9124 8278 9140 8295
rect 9696 8295 9898 8312
rect 9956 8312 10916 8350
rect 9956 8295 10158 8312
rect 9696 8278 9712 8295
rect 9124 8262 9712 8278
rect 8106 8204 8694 8220
rect 8106 8187 8122 8204
rect 7660 8170 7862 8187
rect 6902 8132 7862 8170
rect 7920 8170 8122 8187
rect 8678 8187 8694 8204
rect 10142 8278 10158 8295
rect 10714 8295 10916 8312
rect 10714 8278 10730 8295
rect 10142 8262 10730 8278
rect 9124 8204 9712 8220
rect 9124 8187 9140 8204
rect 8678 8170 8880 8187
rect 7920 8132 8880 8170
rect 8938 8170 9140 8187
rect 9696 8187 9712 8204
rect 10142 8204 10730 8220
rect 10142 8187 10158 8204
rect 9696 8170 9898 8187
rect 8938 8132 9898 8170
rect 9956 8170 10158 8187
rect 10714 8187 10730 8204
rect 10714 8170 10916 8187
rect 9956 8132 10916 8170
rect 13576 7800 14536 7838
rect 13576 7783 13778 7800
rect 13762 7766 13778 7783
rect 14334 7783 14536 7800
rect 14594 7800 15554 7838
rect 14594 7783 14796 7800
rect 14334 7766 14350 7783
rect 13762 7750 14350 7766
rect 14780 7766 14796 7783
rect 15352 7783 15554 7800
rect 15612 7800 16572 7838
rect 15612 7783 15814 7800
rect 15352 7766 15368 7783
rect 14780 7750 15368 7766
rect 15798 7766 15814 7783
rect 16370 7783 16572 7800
rect 16630 7800 17590 7838
rect 16630 7783 16832 7800
rect 16370 7766 16386 7783
rect 15798 7750 16386 7766
rect 16816 7766 16832 7783
rect 17388 7783 17590 7800
rect 17648 7800 18608 7838
rect 17648 7783 17850 7800
rect 17388 7766 17404 7783
rect 16816 7750 17404 7766
rect 17834 7766 17850 7783
rect 18406 7783 18608 7800
rect 18666 7800 19626 7838
rect 18666 7783 18868 7800
rect 18406 7766 18422 7783
rect 17834 7750 18422 7766
rect 18852 7766 18868 7783
rect 19424 7783 19626 7800
rect 19684 7800 20644 7838
rect 19684 7783 19886 7800
rect 19424 7766 19440 7783
rect 18852 7750 19440 7766
rect 19870 7766 19886 7783
rect 20442 7783 20644 7800
rect 20702 7800 21662 7838
rect 20702 7783 20904 7800
rect 20442 7766 20458 7783
rect 19870 7750 20458 7766
rect 20888 7766 20904 7783
rect 21460 7783 21662 7800
rect 21720 7800 22680 7838
rect 21720 7783 21922 7800
rect 21460 7766 21476 7783
rect 20888 7750 21476 7766
rect 21906 7766 21922 7783
rect 22478 7783 22680 7800
rect 22738 7800 23698 7838
rect 22738 7783 22940 7800
rect 22478 7766 22494 7783
rect 21906 7750 22494 7766
rect 22924 7766 22940 7783
rect 23496 7783 23698 7800
rect 23756 7800 24716 7838
rect 23756 7783 23958 7800
rect 23496 7766 23512 7783
rect 22924 7750 23512 7766
rect 23942 7766 23958 7783
rect 24514 7783 24716 7800
rect 24774 7800 25734 7838
rect 24774 7783 24976 7800
rect 24514 7766 24530 7783
rect 23942 7750 24530 7766
rect 24960 7766 24976 7783
rect 25532 7783 25734 7800
rect 25792 7800 26752 7838
rect 25792 7783 25994 7800
rect 25532 7766 25548 7783
rect 24960 7750 25548 7766
rect 25978 7766 25994 7783
rect 26550 7783 26752 7800
rect 26810 7800 27770 7838
rect 26810 7783 27012 7800
rect 26550 7766 26566 7783
rect 25978 7750 26566 7766
rect 26996 7766 27012 7783
rect 27568 7783 27770 7800
rect 27828 7800 28788 7838
rect 27828 7783 28030 7800
rect 27568 7766 27584 7783
rect 26996 7750 27584 7766
rect 28014 7766 28030 7783
rect 28586 7783 28788 7800
rect 28846 7800 29806 7838
rect 28846 7783 29048 7800
rect 28586 7766 28602 7783
rect 28014 7750 28602 7766
rect 29032 7766 29048 7783
rect 29604 7783 29806 7800
rect 29864 7800 30824 7838
rect 29864 7783 30066 7800
rect 29604 7766 29620 7783
rect 29032 7750 29620 7766
rect 30050 7766 30066 7783
rect 30622 7783 30824 7800
rect 30882 7800 31842 7838
rect 30882 7783 31084 7800
rect 30622 7766 30638 7783
rect 30050 7750 30638 7766
rect 31068 7766 31084 7783
rect 31640 7783 31842 7800
rect 31900 7800 32860 7838
rect 31900 7783 32102 7800
rect 31640 7766 31656 7783
rect 31068 7750 31656 7766
rect 32086 7766 32102 7783
rect 32658 7783 32860 7800
rect 32918 7800 33878 7838
rect 32918 7783 33120 7800
rect 32658 7766 32674 7783
rect 32086 7750 32674 7766
rect 33104 7766 33120 7783
rect 33676 7783 33878 7800
rect 33676 7766 33692 7783
rect 33104 7750 33692 7766
rect 1812 7494 2772 7532
rect 1812 7477 2014 7494
rect 1998 7460 2014 7477
rect 2570 7477 2772 7494
rect 2830 7494 3790 7532
rect 2830 7477 3032 7494
rect 2570 7460 2586 7477
rect 1998 7444 2586 7460
rect 3016 7460 3032 7477
rect 3588 7477 3790 7494
rect 3848 7494 4808 7532
rect 3848 7477 4050 7494
rect 3588 7460 3604 7477
rect 3016 7444 3604 7460
rect 4034 7460 4050 7477
rect 4606 7477 4808 7494
rect 4866 7494 5826 7532
rect 4866 7477 5068 7494
rect 4606 7460 4622 7477
rect 4034 7444 4622 7460
rect 5052 7460 5068 7477
rect 5624 7477 5826 7494
rect 5884 7494 6844 7532
rect 5884 7477 6086 7494
rect 5624 7460 5640 7477
rect 5052 7444 5640 7460
rect 6070 7460 6086 7477
rect 6642 7477 6844 7494
rect 6902 7494 7862 7532
rect 6902 7477 7104 7494
rect 6642 7460 6658 7477
rect 6070 7444 6658 7460
rect 7088 7460 7104 7477
rect 7660 7477 7862 7494
rect 7920 7494 8880 7532
rect 7920 7477 8122 7494
rect 7660 7460 7676 7477
rect 7088 7444 7676 7460
rect 8106 7460 8122 7477
rect 8678 7477 8880 7494
rect 8938 7494 9898 7532
rect 8938 7477 9140 7494
rect 8678 7460 8694 7477
rect 8106 7444 8694 7460
rect 9124 7460 9140 7477
rect 9696 7477 9898 7494
rect 9956 7494 10916 7532
rect 9956 7477 10158 7494
rect 9696 7460 9712 7477
rect 9124 7444 9712 7460
rect 10142 7460 10158 7477
rect 10714 7477 10916 7494
rect 10714 7460 10730 7477
rect 10142 7444 10730 7460
rect 13762 7278 14350 7294
rect 13762 7261 13778 7278
rect 13576 7244 13778 7261
rect 14334 7261 14350 7278
rect 14780 7278 15368 7294
rect 14780 7261 14796 7278
rect 14334 7244 14536 7261
rect 13576 7206 14536 7244
rect 14594 7244 14796 7261
rect 15352 7261 15368 7278
rect 15798 7278 16386 7294
rect 15798 7261 15814 7278
rect 15352 7244 15554 7261
rect 14594 7206 15554 7244
rect 15612 7244 15814 7261
rect 16370 7261 16386 7278
rect 16816 7278 17404 7294
rect 16816 7261 16832 7278
rect 16370 7244 16572 7261
rect 15612 7206 16572 7244
rect 16630 7244 16832 7261
rect 17388 7261 17404 7278
rect 17834 7278 18422 7294
rect 17834 7261 17850 7278
rect 17388 7244 17590 7261
rect 16630 7206 17590 7244
rect 17648 7244 17850 7261
rect 18406 7261 18422 7278
rect 18852 7278 19440 7294
rect 18852 7261 18868 7278
rect 18406 7244 18608 7261
rect 17648 7206 18608 7244
rect 18666 7244 18868 7261
rect 19424 7261 19440 7278
rect 19870 7278 20458 7294
rect 19870 7261 19886 7278
rect 19424 7244 19626 7261
rect 18666 7206 19626 7244
rect 19684 7244 19886 7261
rect 20442 7261 20458 7278
rect 20888 7278 21476 7294
rect 20888 7261 20904 7278
rect 20442 7244 20644 7261
rect 19684 7206 20644 7244
rect 20702 7244 20904 7261
rect 21460 7261 21476 7278
rect 21906 7278 22494 7294
rect 21906 7261 21922 7278
rect 21460 7244 21662 7261
rect 20702 7206 21662 7244
rect 21720 7244 21922 7261
rect 22478 7261 22494 7278
rect 22924 7278 23512 7294
rect 22924 7261 22940 7278
rect 22478 7244 22680 7261
rect 21720 7206 22680 7244
rect 22738 7244 22940 7261
rect 23496 7261 23512 7278
rect 23942 7278 24530 7294
rect 23942 7261 23958 7278
rect 23496 7244 23698 7261
rect 22738 7206 23698 7244
rect 23756 7244 23958 7261
rect 24514 7261 24530 7278
rect 24960 7278 25548 7294
rect 24960 7261 24976 7278
rect 24514 7244 24716 7261
rect 23756 7206 24716 7244
rect 24774 7244 24976 7261
rect 25532 7261 25548 7278
rect 25978 7278 26566 7294
rect 25978 7261 25994 7278
rect 25532 7244 25734 7261
rect 24774 7206 25734 7244
rect 25792 7244 25994 7261
rect 26550 7261 26566 7278
rect 26996 7278 27584 7294
rect 26996 7261 27012 7278
rect 26550 7244 26752 7261
rect 25792 7206 26752 7244
rect 26810 7244 27012 7261
rect 27568 7261 27584 7278
rect 28014 7278 28602 7294
rect 28014 7261 28030 7278
rect 27568 7244 27770 7261
rect 26810 7206 27770 7244
rect 27828 7244 28030 7261
rect 28586 7261 28602 7278
rect 29032 7278 29620 7294
rect 29032 7261 29048 7278
rect 28586 7244 28788 7261
rect 27828 7206 28788 7244
rect 28846 7244 29048 7261
rect 29604 7261 29620 7278
rect 30050 7278 30638 7294
rect 30050 7261 30066 7278
rect 29604 7244 29806 7261
rect 28846 7206 29806 7244
rect 29864 7244 30066 7261
rect 30622 7261 30638 7278
rect 31068 7278 31656 7294
rect 31068 7261 31084 7278
rect 30622 7244 30824 7261
rect 29864 7206 30824 7244
rect 30882 7244 31084 7261
rect 31640 7261 31656 7278
rect 32086 7278 32674 7294
rect 32086 7261 32102 7278
rect 31640 7244 31842 7261
rect 30882 7206 31842 7244
rect 31900 7244 32102 7261
rect 32658 7261 32674 7278
rect 33104 7278 33692 7294
rect 33104 7261 33120 7278
rect 32658 7244 32860 7261
rect 31900 7206 32860 7244
rect 32918 7244 33120 7261
rect 33676 7261 33692 7278
rect 33676 7244 33878 7261
rect 32918 7206 33878 7244
rect 13576 6568 14536 6606
rect 13576 6551 13778 6568
rect 13762 6534 13778 6551
rect 14334 6551 14536 6568
rect 14594 6568 15554 6606
rect 14594 6551 14796 6568
rect 14334 6534 14350 6551
rect 13762 6518 14350 6534
rect 14780 6534 14796 6551
rect 15352 6551 15554 6568
rect 15612 6568 16572 6606
rect 15612 6551 15814 6568
rect 15352 6534 15368 6551
rect 14780 6518 15368 6534
rect 15798 6534 15814 6551
rect 16370 6551 16572 6568
rect 16630 6568 17590 6606
rect 16630 6551 16832 6568
rect 16370 6534 16386 6551
rect 15798 6518 16386 6534
rect 16816 6534 16832 6551
rect 17388 6551 17590 6568
rect 17648 6568 18608 6606
rect 17648 6551 17850 6568
rect 17388 6534 17404 6551
rect 16816 6518 17404 6534
rect 17834 6534 17850 6551
rect 18406 6551 18608 6568
rect 18666 6568 19626 6606
rect 18666 6551 18868 6568
rect 18406 6534 18422 6551
rect 17834 6518 18422 6534
rect 18852 6534 18868 6551
rect 19424 6551 19626 6568
rect 19684 6568 20644 6606
rect 19684 6551 19886 6568
rect 19424 6534 19440 6551
rect 18852 6518 19440 6534
rect 19870 6534 19886 6551
rect 20442 6551 20644 6568
rect 20702 6568 21662 6606
rect 20702 6551 20904 6568
rect 20442 6534 20458 6551
rect 19870 6518 20458 6534
rect 20888 6534 20904 6551
rect 21460 6551 21662 6568
rect 21720 6568 22680 6606
rect 21720 6551 21922 6568
rect 21460 6534 21476 6551
rect 20888 6518 21476 6534
rect 21906 6534 21922 6551
rect 22478 6551 22680 6568
rect 22738 6568 23698 6606
rect 22738 6551 22940 6568
rect 22478 6534 22494 6551
rect 21906 6518 22494 6534
rect 22924 6534 22940 6551
rect 23496 6551 23698 6568
rect 23756 6568 24716 6606
rect 23756 6551 23958 6568
rect 23496 6534 23512 6551
rect 22924 6518 23512 6534
rect 23942 6534 23958 6551
rect 24514 6551 24716 6568
rect 24774 6568 25734 6606
rect 24774 6551 24976 6568
rect 24514 6534 24530 6551
rect 23942 6518 24530 6534
rect 24960 6534 24976 6551
rect 25532 6551 25734 6568
rect 25792 6568 26752 6606
rect 25792 6551 25994 6568
rect 25532 6534 25548 6551
rect 24960 6518 25548 6534
rect 25978 6534 25994 6551
rect 26550 6551 26752 6568
rect 26810 6568 27770 6606
rect 26810 6551 27012 6568
rect 26550 6534 26566 6551
rect 25978 6518 26566 6534
rect 26996 6534 27012 6551
rect 27568 6551 27770 6568
rect 27828 6568 28788 6606
rect 27828 6551 28030 6568
rect 27568 6534 27584 6551
rect 26996 6518 27584 6534
rect 28014 6534 28030 6551
rect 28586 6551 28788 6568
rect 28846 6568 29806 6606
rect 28846 6551 29048 6568
rect 28586 6534 28602 6551
rect 28014 6518 28602 6534
rect 29032 6534 29048 6551
rect 29604 6551 29806 6568
rect 29864 6568 30824 6606
rect 29864 6551 30066 6568
rect 29604 6534 29620 6551
rect 29032 6518 29620 6534
rect 30050 6534 30066 6551
rect 30622 6551 30824 6568
rect 30882 6568 31842 6606
rect 30882 6551 31084 6568
rect 30622 6534 30638 6551
rect 30050 6518 30638 6534
rect 31068 6534 31084 6551
rect 31640 6551 31842 6568
rect 31900 6568 32860 6606
rect 31900 6551 32102 6568
rect 31640 6534 31656 6551
rect 31068 6518 31656 6534
rect 32086 6534 32102 6551
rect 32658 6551 32860 6568
rect 32918 6568 33878 6606
rect 32918 6551 33120 6568
rect 32658 6534 32674 6551
rect 32086 6518 32674 6534
rect 33104 6534 33120 6551
rect 33676 6551 33878 6568
rect 33676 6534 33692 6551
rect 33104 6518 33692 6534
rect 674 6180 1262 6196
rect 674 6163 690 6180
rect 488 6146 690 6163
rect 1246 6163 1262 6180
rect 1692 6180 2280 6196
rect 1692 6163 1708 6180
rect 1246 6146 1448 6163
rect 488 6108 1448 6146
rect 1506 6146 1708 6163
rect 2264 6163 2280 6180
rect 2710 6180 3298 6196
rect 2710 6163 2726 6180
rect 2264 6146 2466 6163
rect 1506 6108 2466 6146
rect 2524 6146 2726 6163
rect 3282 6163 3298 6180
rect 3728 6180 4316 6196
rect 3728 6163 3744 6180
rect 3282 6146 3484 6163
rect 2524 6108 3484 6146
rect 3542 6146 3744 6163
rect 4300 6163 4316 6180
rect 4746 6180 5334 6196
rect 4746 6163 4762 6180
rect 4300 6146 4502 6163
rect 3542 6108 4502 6146
rect 4560 6146 4762 6163
rect 5318 6163 5334 6180
rect 5764 6180 6352 6196
rect 5764 6163 5780 6180
rect 5318 6146 5520 6163
rect 4560 6108 5520 6146
rect 5578 6146 5780 6163
rect 6336 6163 6352 6180
rect 6782 6180 7370 6196
rect 6782 6163 6798 6180
rect 6336 6146 6538 6163
rect 5578 6108 6538 6146
rect 6596 6146 6798 6163
rect 7354 6163 7370 6180
rect 7800 6180 8388 6196
rect 7800 6163 7816 6180
rect 7354 6146 7556 6163
rect 6596 6108 7556 6146
rect 7614 6146 7816 6163
rect 8372 6163 8388 6180
rect 8818 6180 9406 6196
rect 8818 6163 8834 6180
rect 8372 6146 8574 6163
rect 7614 6108 8574 6146
rect 8632 6146 8834 6163
rect 9390 6163 9406 6180
rect 9836 6180 10424 6196
rect 9836 6163 9852 6180
rect 9390 6146 9592 6163
rect 8632 6108 9592 6146
rect 9650 6146 9852 6163
rect 10408 6163 10424 6180
rect 10854 6180 11442 6196
rect 10854 6163 10870 6180
rect 10408 6146 10610 6163
rect 9650 6108 10610 6146
rect 10668 6146 10870 6163
rect 11426 6163 11442 6180
rect 11426 6146 11628 6163
rect 10668 6108 11628 6146
rect 13762 6044 14350 6060
rect 13762 6027 13778 6044
rect 13576 6010 13778 6027
rect 14334 6027 14350 6044
rect 14780 6044 15368 6060
rect 14780 6027 14796 6044
rect 14334 6010 14536 6027
rect 13576 5972 14536 6010
rect 14594 6010 14796 6027
rect 15352 6027 15368 6044
rect 15798 6044 16386 6060
rect 15798 6027 15814 6044
rect 15352 6010 15554 6027
rect 14594 5972 15554 6010
rect 15612 6010 15814 6027
rect 16370 6027 16386 6044
rect 16816 6044 17404 6060
rect 16816 6027 16832 6044
rect 16370 6010 16572 6027
rect 15612 5972 16572 6010
rect 16630 6010 16832 6027
rect 17388 6027 17404 6044
rect 17834 6044 18422 6060
rect 17834 6027 17850 6044
rect 17388 6010 17590 6027
rect 16630 5972 17590 6010
rect 17648 6010 17850 6027
rect 18406 6027 18422 6044
rect 18852 6044 19440 6060
rect 18852 6027 18868 6044
rect 18406 6010 18608 6027
rect 17648 5972 18608 6010
rect 18666 6010 18868 6027
rect 19424 6027 19440 6044
rect 19870 6044 20458 6060
rect 19870 6027 19886 6044
rect 19424 6010 19626 6027
rect 18666 5972 19626 6010
rect 19684 6010 19886 6027
rect 20442 6027 20458 6044
rect 20888 6044 21476 6060
rect 20888 6027 20904 6044
rect 20442 6010 20644 6027
rect 19684 5972 20644 6010
rect 20702 6010 20904 6027
rect 21460 6027 21476 6044
rect 21906 6044 22494 6060
rect 21906 6027 21922 6044
rect 21460 6010 21662 6027
rect 20702 5972 21662 6010
rect 21720 6010 21922 6027
rect 22478 6027 22494 6044
rect 22924 6044 23512 6060
rect 22924 6027 22940 6044
rect 22478 6010 22680 6027
rect 21720 5972 22680 6010
rect 22738 6010 22940 6027
rect 23496 6027 23512 6044
rect 23942 6044 24530 6060
rect 23942 6027 23958 6044
rect 23496 6010 23698 6027
rect 22738 5972 23698 6010
rect 23756 6010 23958 6027
rect 24514 6027 24530 6044
rect 24960 6044 25548 6060
rect 24960 6027 24976 6044
rect 24514 6010 24716 6027
rect 23756 5972 24716 6010
rect 24774 6010 24976 6027
rect 25532 6027 25548 6044
rect 25978 6044 26566 6060
rect 25978 6027 25994 6044
rect 25532 6010 25734 6027
rect 24774 5972 25734 6010
rect 25792 6010 25994 6027
rect 26550 6027 26566 6044
rect 26996 6044 27584 6060
rect 26996 6027 27012 6044
rect 26550 6010 26752 6027
rect 25792 5972 26752 6010
rect 26810 6010 27012 6027
rect 27568 6027 27584 6044
rect 28014 6044 28602 6060
rect 28014 6027 28030 6044
rect 27568 6010 27770 6027
rect 26810 5972 27770 6010
rect 27828 6010 28030 6027
rect 28586 6027 28602 6044
rect 29032 6044 29620 6060
rect 29032 6027 29048 6044
rect 28586 6010 28788 6027
rect 27828 5972 28788 6010
rect 28846 6010 29048 6027
rect 29604 6027 29620 6044
rect 30050 6044 30638 6060
rect 30050 6027 30066 6044
rect 29604 6010 29806 6027
rect 28846 5972 29806 6010
rect 29864 6010 30066 6027
rect 30622 6027 30638 6044
rect 31068 6044 31656 6060
rect 31068 6027 31084 6044
rect 30622 6010 30824 6027
rect 29864 5972 30824 6010
rect 30882 6010 31084 6027
rect 31640 6027 31656 6044
rect 32086 6044 32674 6060
rect 32086 6027 32102 6044
rect 31640 6010 31842 6027
rect 30882 5972 31842 6010
rect 31900 6010 32102 6027
rect 32658 6027 32674 6044
rect 33104 6044 33692 6060
rect 33104 6027 33120 6044
rect 32658 6010 32860 6027
rect 31900 5972 32860 6010
rect 32918 6010 33120 6027
rect 33676 6027 33692 6044
rect 33676 6010 33878 6027
rect 32918 5972 33878 6010
rect 488 5470 1448 5508
rect 488 5453 690 5470
rect 674 5436 690 5453
rect 1246 5453 1448 5470
rect 1506 5470 2466 5508
rect 1506 5453 1708 5470
rect 1246 5436 1262 5453
rect 674 5420 1262 5436
rect 1692 5436 1708 5453
rect 2264 5453 2466 5470
rect 2524 5470 3484 5508
rect 2524 5453 2726 5470
rect 2264 5436 2280 5453
rect 1692 5420 2280 5436
rect 2710 5436 2726 5453
rect 3282 5453 3484 5470
rect 3542 5470 4502 5508
rect 3542 5453 3744 5470
rect 3282 5436 3298 5453
rect 2710 5420 3298 5436
rect 3728 5436 3744 5453
rect 4300 5453 4502 5470
rect 4560 5470 5520 5508
rect 4560 5453 4762 5470
rect 4300 5436 4316 5453
rect 3728 5420 4316 5436
rect 4746 5436 4762 5453
rect 5318 5453 5520 5470
rect 5578 5470 6538 5508
rect 5578 5453 5780 5470
rect 5318 5436 5334 5453
rect 4746 5420 5334 5436
rect 5764 5436 5780 5453
rect 6336 5453 6538 5470
rect 6596 5470 7556 5508
rect 6596 5453 6798 5470
rect 6336 5436 6352 5453
rect 5764 5420 6352 5436
rect 6782 5436 6798 5453
rect 7354 5453 7556 5470
rect 7614 5470 8574 5508
rect 7614 5453 7816 5470
rect 7354 5436 7370 5453
rect 6782 5420 7370 5436
rect 7800 5436 7816 5453
rect 8372 5453 8574 5470
rect 8632 5470 9592 5508
rect 8632 5453 8834 5470
rect 8372 5436 8388 5453
rect 7800 5420 8388 5436
rect 8818 5436 8834 5453
rect 9390 5453 9592 5470
rect 9650 5470 10610 5508
rect 9650 5453 9852 5470
rect 9390 5436 9406 5453
rect 8818 5420 9406 5436
rect 9836 5436 9852 5453
rect 10408 5453 10610 5470
rect 10668 5470 11628 5508
rect 10668 5453 10870 5470
rect 10408 5436 10424 5453
rect 9836 5420 10424 5436
rect 10854 5436 10870 5453
rect 11426 5453 11628 5470
rect 11426 5436 11442 5453
rect 10854 5420 11442 5436
rect 13576 5334 14536 5372
rect 13576 5317 13778 5334
rect 13762 5300 13778 5317
rect 14334 5317 14536 5334
rect 14594 5334 15554 5372
rect 14594 5317 14796 5334
rect 14334 5300 14350 5317
rect 13762 5284 14350 5300
rect 14780 5300 14796 5317
rect 15352 5317 15554 5334
rect 15612 5334 16572 5372
rect 15612 5317 15814 5334
rect 15352 5300 15368 5317
rect 14780 5284 15368 5300
rect 15798 5300 15814 5317
rect 16370 5317 16572 5334
rect 16630 5334 17590 5372
rect 16630 5317 16832 5334
rect 16370 5300 16386 5317
rect 15798 5284 16386 5300
rect 16816 5300 16832 5317
rect 17388 5317 17590 5334
rect 17648 5334 18608 5372
rect 17648 5317 17850 5334
rect 17388 5300 17404 5317
rect 16816 5284 17404 5300
rect 17834 5300 17850 5317
rect 18406 5317 18608 5334
rect 18666 5334 19626 5372
rect 18666 5317 18868 5334
rect 18406 5300 18422 5317
rect 17834 5284 18422 5300
rect 18852 5300 18868 5317
rect 19424 5317 19626 5334
rect 19684 5334 20644 5372
rect 19684 5317 19886 5334
rect 19424 5300 19440 5317
rect 18852 5284 19440 5300
rect 19870 5300 19886 5317
rect 20442 5317 20644 5334
rect 20702 5334 21662 5372
rect 20702 5317 20904 5334
rect 20442 5300 20458 5317
rect 19870 5284 20458 5300
rect 20888 5300 20904 5317
rect 21460 5317 21662 5334
rect 21720 5334 22680 5372
rect 21720 5317 21922 5334
rect 21460 5300 21476 5317
rect 20888 5284 21476 5300
rect 21906 5300 21922 5317
rect 22478 5317 22680 5334
rect 22738 5334 23698 5372
rect 22738 5317 22940 5334
rect 22478 5300 22494 5317
rect 21906 5284 22494 5300
rect 22924 5300 22940 5317
rect 23496 5317 23698 5334
rect 23756 5334 24716 5372
rect 23756 5317 23958 5334
rect 23496 5300 23512 5317
rect 22924 5284 23512 5300
rect 23942 5300 23958 5317
rect 24514 5317 24716 5334
rect 24774 5334 25734 5372
rect 24774 5317 24976 5334
rect 24514 5300 24530 5317
rect 23942 5284 24530 5300
rect 24960 5300 24976 5317
rect 25532 5317 25734 5334
rect 25792 5334 26752 5372
rect 25792 5317 25994 5334
rect 25532 5300 25548 5317
rect 24960 5284 25548 5300
rect 25978 5300 25994 5317
rect 26550 5317 26752 5334
rect 26810 5334 27770 5372
rect 26810 5317 27012 5334
rect 26550 5300 26566 5317
rect 25978 5284 26566 5300
rect 26996 5300 27012 5317
rect 27568 5317 27770 5334
rect 27828 5334 28788 5372
rect 27828 5317 28030 5334
rect 27568 5300 27584 5317
rect 26996 5284 27584 5300
rect 28014 5300 28030 5317
rect 28586 5317 28788 5334
rect 28846 5334 29806 5372
rect 28846 5317 29048 5334
rect 28586 5300 28602 5317
rect 28014 5284 28602 5300
rect 29032 5300 29048 5317
rect 29604 5317 29806 5334
rect 29864 5334 30824 5372
rect 29864 5317 30066 5334
rect 29604 5300 29620 5317
rect 29032 5284 29620 5300
rect 30050 5300 30066 5317
rect 30622 5317 30824 5334
rect 30882 5334 31842 5372
rect 30882 5317 31084 5334
rect 30622 5300 30638 5317
rect 30050 5284 30638 5300
rect 31068 5300 31084 5317
rect 31640 5317 31842 5334
rect 31900 5334 32860 5372
rect 31900 5317 32102 5334
rect 31640 5300 31656 5317
rect 31068 5284 31656 5300
rect 32086 5300 32102 5317
rect 32658 5317 32860 5334
rect 32918 5334 33878 5372
rect 32918 5317 33120 5334
rect 32658 5300 32674 5317
rect 32086 5284 32674 5300
rect 33104 5300 33120 5317
rect 33676 5317 33878 5334
rect 33676 5300 33692 5317
rect 33104 5284 33692 5300
rect 674 5068 1262 5084
rect 674 5051 690 5068
rect 488 5034 690 5051
rect 1246 5051 1262 5068
rect 1692 5068 2280 5084
rect 1692 5051 1708 5068
rect 1246 5034 1448 5051
rect 488 4996 1448 5034
rect 1506 5034 1708 5051
rect 2264 5051 2280 5068
rect 2710 5068 3298 5084
rect 2710 5051 2726 5068
rect 2264 5034 2466 5051
rect 1506 4996 2466 5034
rect 2524 5034 2726 5051
rect 3282 5051 3298 5068
rect 3728 5068 4316 5084
rect 3728 5051 3744 5068
rect 3282 5034 3484 5051
rect 2524 4996 3484 5034
rect 3542 5034 3744 5051
rect 4300 5051 4316 5068
rect 4746 5068 5334 5084
rect 4746 5051 4762 5068
rect 4300 5034 4502 5051
rect 3542 4996 4502 5034
rect 4560 5034 4762 5051
rect 5318 5051 5334 5068
rect 5764 5068 6352 5084
rect 5764 5051 5780 5068
rect 5318 5034 5520 5051
rect 4560 4996 5520 5034
rect 5578 5034 5780 5051
rect 6336 5051 6352 5068
rect 6782 5068 7370 5084
rect 6782 5051 6798 5068
rect 6336 5034 6538 5051
rect 5578 4996 6538 5034
rect 6596 5034 6798 5051
rect 7354 5051 7370 5068
rect 7800 5068 8388 5084
rect 7800 5051 7816 5068
rect 7354 5034 7556 5051
rect 6596 4996 7556 5034
rect 7614 5034 7816 5051
rect 8372 5051 8388 5068
rect 8818 5068 9406 5084
rect 8818 5051 8834 5068
rect 8372 5034 8574 5051
rect 7614 4996 8574 5034
rect 8632 5034 8834 5051
rect 9390 5051 9406 5068
rect 9836 5068 10424 5084
rect 9836 5051 9852 5068
rect 9390 5034 9592 5051
rect 8632 4996 9592 5034
rect 9650 5034 9852 5051
rect 10408 5051 10424 5068
rect 10854 5068 11442 5084
rect 10854 5051 10870 5068
rect 10408 5034 10610 5051
rect 9650 4996 10610 5034
rect 10668 5034 10870 5051
rect 11426 5051 11442 5068
rect 11426 5034 11628 5051
rect 10668 4996 11628 5034
rect 13762 4810 14350 4826
rect 13762 4793 13778 4810
rect 13576 4776 13778 4793
rect 14334 4793 14350 4810
rect 14780 4810 15368 4826
rect 14780 4793 14796 4810
rect 14334 4776 14536 4793
rect 13576 4738 14536 4776
rect 14594 4776 14796 4793
rect 15352 4793 15368 4810
rect 15798 4810 16386 4826
rect 15798 4793 15814 4810
rect 15352 4776 15554 4793
rect 14594 4738 15554 4776
rect 15612 4776 15814 4793
rect 16370 4793 16386 4810
rect 16816 4810 17404 4826
rect 16816 4793 16832 4810
rect 16370 4776 16572 4793
rect 15612 4738 16572 4776
rect 16630 4776 16832 4793
rect 17388 4793 17404 4810
rect 17834 4810 18422 4826
rect 17834 4793 17850 4810
rect 17388 4776 17590 4793
rect 16630 4738 17590 4776
rect 17648 4776 17850 4793
rect 18406 4793 18422 4810
rect 18852 4810 19440 4826
rect 18852 4793 18868 4810
rect 18406 4776 18608 4793
rect 17648 4738 18608 4776
rect 18666 4776 18868 4793
rect 19424 4793 19440 4810
rect 19870 4810 20458 4826
rect 19870 4793 19886 4810
rect 19424 4776 19626 4793
rect 18666 4738 19626 4776
rect 19684 4776 19886 4793
rect 20442 4793 20458 4810
rect 20888 4810 21476 4826
rect 20888 4793 20904 4810
rect 20442 4776 20644 4793
rect 19684 4738 20644 4776
rect 20702 4776 20904 4793
rect 21460 4793 21476 4810
rect 21906 4810 22494 4826
rect 21906 4793 21922 4810
rect 21460 4776 21662 4793
rect 20702 4738 21662 4776
rect 21720 4776 21922 4793
rect 22478 4793 22494 4810
rect 22924 4810 23512 4826
rect 22924 4793 22940 4810
rect 22478 4776 22680 4793
rect 21720 4738 22680 4776
rect 22738 4776 22940 4793
rect 23496 4793 23512 4810
rect 23942 4810 24530 4826
rect 23942 4793 23958 4810
rect 23496 4776 23698 4793
rect 22738 4738 23698 4776
rect 23756 4776 23958 4793
rect 24514 4793 24530 4810
rect 24960 4810 25548 4826
rect 24960 4793 24976 4810
rect 24514 4776 24716 4793
rect 23756 4738 24716 4776
rect 24774 4776 24976 4793
rect 25532 4793 25548 4810
rect 25978 4810 26566 4826
rect 25978 4793 25994 4810
rect 25532 4776 25734 4793
rect 24774 4738 25734 4776
rect 25792 4776 25994 4793
rect 26550 4793 26566 4810
rect 26996 4810 27584 4826
rect 26996 4793 27012 4810
rect 26550 4776 26752 4793
rect 25792 4738 26752 4776
rect 26810 4776 27012 4793
rect 27568 4793 27584 4810
rect 28014 4810 28602 4826
rect 28014 4793 28030 4810
rect 27568 4776 27770 4793
rect 26810 4738 27770 4776
rect 27828 4776 28030 4793
rect 28586 4793 28602 4810
rect 29032 4810 29620 4826
rect 29032 4793 29048 4810
rect 28586 4776 28788 4793
rect 27828 4738 28788 4776
rect 28846 4776 29048 4793
rect 29604 4793 29620 4810
rect 30050 4810 30638 4826
rect 30050 4793 30066 4810
rect 29604 4776 29806 4793
rect 28846 4738 29806 4776
rect 29864 4776 30066 4793
rect 30622 4793 30638 4810
rect 31068 4810 31656 4826
rect 31068 4793 31084 4810
rect 30622 4776 30824 4793
rect 29864 4738 30824 4776
rect 30882 4776 31084 4793
rect 31640 4793 31656 4810
rect 32086 4810 32674 4826
rect 32086 4793 32102 4810
rect 31640 4776 31842 4793
rect 30882 4738 31842 4776
rect 31900 4776 32102 4793
rect 32658 4793 32674 4810
rect 33104 4810 33692 4826
rect 33104 4793 33120 4810
rect 32658 4776 32860 4793
rect 31900 4738 32860 4776
rect 32918 4776 33120 4793
rect 33676 4793 33692 4810
rect 33676 4776 33878 4793
rect 32918 4738 33878 4776
rect 488 4358 1448 4396
rect 488 4341 690 4358
rect 674 4324 690 4341
rect 1246 4341 1448 4358
rect 1506 4358 2466 4396
rect 1506 4341 1708 4358
rect 1246 4324 1262 4341
rect 674 4308 1262 4324
rect 1692 4324 1708 4341
rect 2264 4341 2466 4358
rect 2524 4358 3484 4396
rect 2524 4341 2726 4358
rect 2264 4324 2280 4341
rect 1692 4308 2280 4324
rect 2710 4324 2726 4341
rect 3282 4341 3484 4358
rect 3542 4358 4502 4396
rect 3542 4341 3744 4358
rect 3282 4324 3298 4341
rect 2710 4308 3298 4324
rect 3728 4324 3744 4341
rect 4300 4341 4502 4358
rect 4560 4358 5520 4396
rect 4560 4341 4762 4358
rect 4300 4324 4316 4341
rect 3728 4308 4316 4324
rect 4746 4324 4762 4341
rect 5318 4341 5520 4358
rect 5578 4358 6538 4396
rect 5578 4341 5780 4358
rect 5318 4324 5334 4341
rect 4746 4308 5334 4324
rect 5764 4324 5780 4341
rect 6336 4341 6538 4358
rect 6596 4358 7556 4396
rect 6596 4341 6798 4358
rect 6336 4324 6352 4341
rect 5764 4308 6352 4324
rect 6782 4324 6798 4341
rect 7354 4341 7556 4358
rect 7614 4358 8574 4396
rect 7614 4341 7816 4358
rect 7354 4324 7370 4341
rect 6782 4308 7370 4324
rect 7800 4324 7816 4341
rect 8372 4341 8574 4358
rect 8632 4358 9592 4396
rect 8632 4341 8834 4358
rect 8372 4324 8388 4341
rect 7800 4308 8388 4324
rect 8818 4324 8834 4341
rect 9390 4341 9592 4358
rect 9650 4358 10610 4396
rect 9650 4341 9852 4358
rect 9390 4324 9406 4341
rect 8818 4308 9406 4324
rect 9836 4324 9852 4341
rect 10408 4341 10610 4358
rect 10668 4358 11628 4396
rect 10668 4341 10870 4358
rect 10408 4324 10424 4341
rect 9836 4308 10424 4324
rect 10854 4324 10870 4341
rect 11426 4341 11628 4358
rect 11426 4324 11442 4341
rect 10854 4308 11442 4324
rect 13576 4100 14536 4138
rect 13576 4083 13778 4100
rect 13762 4066 13778 4083
rect 14334 4083 14536 4100
rect 14594 4100 15554 4138
rect 14594 4083 14796 4100
rect 14334 4066 14350 4083
rect 13762 4050 14350 4066
rect 14780 4066 14796 4083
rect 15352 4083 15554 4100
rect 15612 4100 16572 4138
rect 15612 4083 15814 4100
rect 15352 4066 15368 4083
rect 14780 4050 15368 4066
rect 15798 4066 15814 4083
rect 16370 4083 16572 4100
rect 16630 4100 17590 4138
rect 16630 4083 16832 4100
rect 16370 4066 16386 4083
rect 15798 4050 16386 4066
rect 16816 4066 16832 4083
rect 17388 4083 17590 4100
rect 17648 4100 18608 4138
rect 17648 4083 17850 4100
rect 17388 4066 17404 4083
rect 16816 4050 17404 4066
rect 17834 4066 17850 4083
rect 18406 4083 18608 4100
rect 18666 4100 19626 4138
rect 18666 4083 18868 4100
rect 18406 4066 18422 4083
rect 17834 4050 18422 4066
rect 18852 4066 18868 4083
rect 19424 4083 19626 4100
rect 19684 4100 20644 4138
rect 19684 4083 19886 4100
rect 19424 4066 19440 4083
rect 18852 4050 19440 4066
rect 19870 4066 19886 4083
rect 20442 4083 20644 4100
rect 20702 4100 21662 4138
rect 20702 4083 20904 4100
rect 20442 4066 20458 4083
rect 19870 4050 20458 4066
rect 20888 4066 20904 4083
rect 21460 4083 21662 4100
rect 21720 4100 22680 4138
rect 21720 4083 21922 4100
rect 21460 4066 21476 4083
rect 20888 4050 21476 4066
rect 21906 4066 21922 4083
rect 22478 4083 22680 4100
rect 22738 4100 23698 4138
rect 22738 4083 22940 4100
rect 22478 4066 22494 4083
rect 21906 4050 22494 4066
rect 22924 4066 22940 4083
rect 23496 4083 23698 4100
rect 23756 4100 24716 4138
rect 23756 4083 23958 4100
rect 23496 4066 23512 4083
rect 22924 4050 23512 4066
rect 23942 4066 23958 4083
rect 24514 4083 24716 4100
rect 24774 4100 25734 4138
rect 24774 4083 24976 4100
rect 24514 4066 24530 4083
rect 23942 4050 24530 4066
rect 24960 4066 24976 4083
rect 25532 4083 25734 4100
rect 25792 4100 26752 4138
rect 25792 4083 25994 4100
rect 25532 4066 25548 4083
rect 24960 4050 25548 4066
rect 25978 4066 25994 4083
rect 26550 4083 26752 4100
rect 26810 4100 27770 4138
rect 26810 4083 27012 4100
rect 26550 4066 26566 4083
rect 25978 4050 26566 4066
rect 26996 4066 27012 4083
rect 27568 4083 27770 4100
rect 27828 4100 28788 4138
rect 27828 4083 28030 4100
rect 27568 4066 27584 4083
rect 26996 4050 27584 4066
rect 28014 4066 28030 4083
rect 28586 4083 28788 4100
rect 28846 4100 29806 4138
rect 28846 4083 29048 4100
rect 28586 4066 28602 4083
rect 28014 4050 28602 4066
rect 29032 4066 29048 4083
rect 29604 4083 29806 4100
rect 29864 4100 30824 4138
rect 29864 4083 30066 4100
rect 29604 4066 29620 4083
rect 29032 4050 29620 4066
rect 30050 4066 30066 4083
rect 30622 4083 30824 4100
rect 30882 4100 31842 4138
rect 30882 4083 31084 4100
rect 30622 4066 30638 4083
rect 30050 4050 30638 4066
rect 31068 4066 31084 4083
rect 31640 4083 31842 4100
rect 31900 4100 32860 4138
rect 31900 4083 32102 4100
rect 31640 4066 31656 4083
rect 31068 4050 31656 4066
rect 32086 4066 32102 4083
rect 32658 4083 32860 4100
rect 32918 4100 33878 4138
rect 32918 4083 33120 4100
rect 32658 4066 32674 4083
rect 32086 4050 32674 4066
rect 33104 4066 33120 4083
rect 33676 4083 33878 4100
rect 33676 4066 33692 4083
rect 33104 4050 33692 4066
rect 674 3956 1262 3972
rect 674 3939 690 3956
rect 488 3922 690 3939
rect 1246 3939 1262 3956
rect 1692 3956 2280 3972
rect 1692 3939 1708 3956
rect 1246 3922 1448 3939
rect 488 3884 1448 3922
rect 1506 3922 1708 3939
rect 2264 3939 2280 3956
rect 2710 3956 3298 3972
rect 2710 3939 2726 3956
rect 2264 3922 2466 3939
rect 1506 3884 2466 3922
rect 2524 3922 2726 3939
rect 3282 3939 3298 3956
rect 3728 3956 4316 3972
rect 3728 3939 3744 3956
rect 3282 3922 3484 3939
rect 2524 3884 3484 3922
rect 3542 3922 3744 3939
rect 4300 3939 4316 3956
rect 4746 3956 5334 3972
rect 4746 3939 4762 3956
rect 4300 3922 4502 3939
rect 3542 3884 4502 3922
rect 4560 3922 4762 3939
rect 5318 3939 5334 3956
rect 5764 3956 6352 3972
rect 5764 3939 5780 3956
rect 5318 3922 5520 3939
rect 4560 3884 5520 3922
rect 5578 3922 5780 3939
rect 6336 3939 6352 3956
rect 6782 3956 7370 3972
rect 6782 3939 6798 3956
rect 6336 3922 6538 3939
rect 5578 3884 6538 3922
rect 6596 3922 6798 3939
rect 7354 3939 7370 3956
rect 7800 3956 8388 3972
rect 7800 3939 7816 3956
rect 7354 3922 7556 3939
rect 6596 3884 7556 3922
rect 7614 3922 7816 3939
rect 8372 3939 8388 3956
rect 8818 3956 9406 3972
rect 8818 3939 8834 3956
rect 8372 3922 8574 3939
rect 7614 3884 8574 3922
rect 8632 3922 8834 3939
rect 9390 3939 9406 3956
rect 9836 3956 10424 3972
rect 9836 3939 9852 3956
rect 9390 3922 9592 3939
rect 8632 3884 9592 3922
rect 9650 3922 9852 3939
rect 10408 3939 10424 3956
rect 10854 3956 11442 3972
rect 10854 3939 10870 3956
rect 10408 3922 10610 3939
rect 9650 3884 10610 3922
rect 10668 3922 10870 3939
rect 11426 3939 11442 3956
rect 11426 3922 11628 3939
rect 10668 3884 11628 3922
rect 13762 3578 14350 3594
rect 13762 3561 13778 3578
rect 13576 3544 13778 3561
rect 14334 3561 14350 3578
rect 14780 3578 15368 3594
rect 14780 3561 14796 3578
rect 14334 3544 14536 3561
rect 13576 3506 14536 3544
rect 14594 3544 14796 3561
rect 15352 3561 15368 3578
rect 15798 3578 16386 3594
rect 15798 3561 15814 3578
rect 15352 3544 15554 3561
rect 14594 3506 15554 3544
rect 15612 3544 15814 3561
rect 16370 3561 16386 3578
rect 16816 3578 17404 3594
rect 16816 3561 16832 3578
rect 16370 3544 16572 3561
rect 15612 3506 16572 3544
rect 16630 3544 16832 3561
rect 17388 3561 17404 3578
rect 17834 3578 18422 3594
rect 17834 3561 17850 3578
rect 17388 3544 17590 3561
rect 16630 3506 17590 3544
rect 17648 3544 17850 3561
rect 18406 3561 18422 3578
rect 18852 3578 19440 3594
rect 18852 3561 18868 3578
rect 18406 3544 18608 3561
rect 17648 3506 18608 3544
rect 18666 3544 18868 3561
rect 19424 3561 19440 3578
rect 19870 3578 20458 3594
rect 19870 3561 19886 3578
rect 19424 3544 19626 3561
rect 18666 3506 19626 3544
rect 19684 3544 19886 3561
rect 20442 3561 20458 3578
rect 20888 3578 21476 3594
rect 20888 3561 20904 3578
rect 20442 3544 20644 3561
rect 19684 3506 20644 3544
rect 20702 3544 20904 3561
rect 21460 3561 21476 3578
rect 21906 3578 22494 3594
rect 21906 3561 21922 3578
rect 21460 3544 21662 3561
rect 20702 3506 21662 3544
rect 21720 3544 21922 3561
rect 22478 3561 22494 3578
rect 22924 3578 23512 3594
rect 22924 3561 22940 3578
rect 22478 3544 22680 3561
rect 21720 3506 22680 3544
rect 22738 3544 22940 3561
rect 23496 3561 23512 3578
rect 23942 3578 24530 3594
rect 23942 3561 23958 3578
rect 23496 3544 23698 3561
rect 22738 3506 23698 3544
rect 23756 3544 23958 3561
rect 24514 3561 24530 3578
rect 24960 3578 25548 3594
rect 24960 3561 24976 3578
rect 24514 3544 24716 3561
rect 23756 3506 24716 3544
rect 24774 3544 24976 3561
rect 25532 3561 25548 3578
rect 25978 3578 26566 3594
rect 25978 3561 25994 3578
rect 25532 3544 25734 3561
rect 24774 3506 25734 3544
rect 25792 3544 25994 3561
rect 26550 3561 26566 3578
rect 26996 3578 27584 3594
rect 26996 3561 27012 3578
rect 26550 3544 26752 3561
rect 25792 3506 26752 3544
rect 26810 3544 27012 3561
rect 27568 3561 27584 3578
rect 28014 3578 28602 3594
rect 28014 3561 28030 3578
rect 27568 3544 27770 3561
rect 26810 3506 27770 3544
rect 27828 3544 28030 3561
rect 28586 3561 28602 3578
rect 29032 3578 29620 3594
rect 29032 3561 29048 3578
rect 28586 3544 28788 3561
rect 27828 3506 28788 3544
rect 28846 3544 29048 3561
rect 29604 3561 29620 3578
rect 30050 3578 30638 3594
rect 30050 3561 30066 3578
rect 29604 3544 29806 3561
rect 28846 3506 29806 3544
rect 29864 3544 30066 3561
rect 30622 3561 30638 3578
rect 31068 3578 31656 3594
rect 31068 3561 31084 3578
rect 30622 3544 30824 3561
rect 29864 3506 30824 3544
rect 30882 3544 31084 3561
rect 31640 3561 31656 3578
rect 32086 3578 32674 3594
rect 32086 3561 32102 3578
rect 31640 3544 31842 3561
rect 30882 3506 31842 3544
rect 31900 3544 32102 3561
rect 32658 3561 32674 3578
rect 33104 3578 33692 3594
rect 33104 3561 33120 3578
rect 32658 3544 32860 3561
rect 31900 3506 32860 3544
rect 32918 3544 33120 3561
rect 33676 3561 33692 3578
rect 33676 3544 33878 3561
rect 32918 3506 33878 3544
rect 488 3246 1448 3284
rect 488 3229 690 3246
rect 674 3212 690 3229
rect 1246 3229 1448 3246
rect 1506 3246 2466 3284
rect 1506 3229 1708 3246
rect 1246 3212 1262 3229
rect 674 3196 1262 3212
rect 1692 3212 1708 3229
rect 2264 3229 2466 3246
rect 2524 3246 3484 3284
rect 2524 3229 2726 3246
rect 2264 3212 2280 3229
rect 1692 3196 2280 3212
rect 2710 3212 2726 3229
rect 3282 3229 3484 3246
rect 3542 3246 4502 3284
rect 3542 3229 3744 3246
rect 3282 3212 3298 3229
rect 2710 3196 3298 3212
rect 3728 3212 3744 3229
rect 4300 3229 4502 3246
rect 4560 3246 5520 3284
rect 4560 3229 4762 3246
rect 4300 3212 4316 3229
rect 3728 3196 4316 3212
rect 4746 3212 4762 3229
rect 5318 3229 5520 3246
rect 5578 3246 6538 3284
rect 5578 3229 5780 3246
rect 5318 3212 5334 3229
rect 4746 3196 5334 3212
rect 5764 3212 5780 3229
rect 6336 3229 6538 3246
rect 6596 3246 7556 3284
rect 6596 3229 6798 3246
rect 6336 3212 6352 3229
rect 5764 3196 6352 3212
rect 6782 3212 6798 3229
rect 7354 3229 7556 3246
rect 7614 3246 8574 3284
rect 7614 3229 7816 3246
rect 7354 3212 7370 3229
rect 6782 3196 7370 3212
rect 7800 3212 7816 3229
rect 8372 3229 8574 3246
rect 8632 3246 9592 3284
rect 8632 3229 8834 3246
rect 8372 3212 8388 3229
rect 7800 3196 8388 3212
rect 8818 3212 8834 3229
rect 9390 3229 9592 3246
rect 9650 3246 10610 3284
rect 9650 3229 9852 3246
rect 9390 3212 9406 3229
rect 8818 3196 9406 3212
rect 9836 3212 9852 3229
rect 10408 3229 10610 3246
rect 10668 3246 11628 3284
rect 10668 3229 10870 3246
rect 10408 3212 10424 3229
rect 9836 3196 10424 3212
rect 10854 3212 10870 3229
rect 11426 3229 11628 3246
rect 11426 3212 11442 3229
rect 10854 3196 11442 3212
rect 13576 2868 14536 2906
rect 674 2844 1262 2860
rect 674 2827 690 2844
rect 488 2810 690 2827
rect 1246 2827 1262 2844
rect 1692 2844 2280 2860
rect 1692 2827 1708 2844
rect 1246 2810 1448 2827
rect 488 2772 1448 2810
rect 1506 2810 1708 2827
rect 2264 2827 2280 2844
rect 2710 2844 3298 2860
rect 2710 2827 2726 2844
rect 2264 2810 2466 2827
rect 1506 2772 2466 2810
rect 2524 2810 2726 2827
rect 3282 2827 3298 2844
rect 3728 2844 4316 2860
rect 3728 2827 3744 2844
rect 3282 2810 3484 2827
rect 2524 2772 3484 2810
rect 3542 2810 3744 2827
rect 4300 2827 4316 2844
rect 4746 2844 5334 2860
rect 4746 2827 4762 2844
rect 4300 2810 4502 2827
rect 3542 2772 4502 2810
rect 4560 2810 4762 2827
rect 5318 2827 5334 2844
rect 5764 2844 6352 2860
rect 5764 2827 5780 2844
rect 5318 2810 5520 2827
rect 4560 2772 5520 2810
rect 5578 2810 5780 2827
rect 6336 2827 6352 2844
rect 6782 2844 7370 2860
rect 6782 2827 6798 2844
rect 6336 2810 6538 2827
rect 5578 2772 6538 2810
rect 6596 2810 6798 2827
rect 7354 2827 7370 2844
rect 7800 2844 8388 2860
rect 7800 2827 7816 2844
rect 7354 2810 7556 2827
rect 6596 2772 7556 2810
rect 7614 2810 7816 2827
rect 8372 2827 8388 2844
rect 8818 2844 9406 2860
rect 8818 2827 8834 2844
rect 8372 2810 8574 2827
rect 7614 2772 8574 2810
rect 8632 2810 8834 2827
rect 9390 2827 9406 2844
rect 9836 2844 10424 2860
rect 9836 2827 9852 2844
rect 9390 2810 9592 2827
rect 8632 2772 9592 2810
rect 9650 2810 9852 2827
rect 10408 2827 10424 2844
rect 10854 2844 11442 2860
rect 13576 2851 13778 2868
rect 10854 2827 10870 2844
rect 10408 2810 10610 2827
rect 9650 2772 10610 2810
rect 10668 2810 10870 2827
rect 11426 2827 11442 2844
rect 13762 2834 13778 2851
rect 14334 2851 14536 2868
rect 14594 2868 15554 2906
rect 14594 2851 14796 2868
rect 14334 2834 14350 2851
rect 11426 2810 11628 2827
rect 13762 2818 14350 2834
rect 14780 2834 14796 2851
rect 15352 2851 15554 2868
rect 15612 2868 16572 2906
rect 15612 2851 15814 2868
rect 15352 2834 15368 2851
rect 14780 2818 15368 2834
rect 15798 2834 15814 2851
rect 16370 2851 16572 2868
rect 16630 2868 17590 2906
rect 16630 2851 16832 2868
rect 16370 2834 16386 2851
rect 15798 2818 16386 2834
rect 16816 2834 16832 2851
rect 17388 2851 17590 2868
rect 17648 2868 18608 2906
rect 17648 2851 17850 2868
rect 17388 2834 17404 2851
rect 16816 2818 17404 2834
rect 17834 2834 17850 2851
rect 18406 2851 18608 2868
rect 18666 2868 19626 2906
rect 18666 2851 18868 2868
rect 18406 2834 18422 2851
rect 17834 2818 18422 2834
rect 18852 2834 18868 2851
rect 19424 2851 19626 2868
rect 19684 2868 20644 2906
rect 19684 2851 19886 2868
rect 19424 2834 19440 2851
rect 18852 2818 19440 2834
rect 19870 2834 19886 2851
rect 20442 2851 20644 2868
rect 20702 2868 21662 2906
rect 20702 2851 20904 2868
rect 20442 2834 20458 2851
rect 19870 2818 20458 2834
rect 20888 2834 20904 2851
rect 21460 2851 21662 2868
rect 21720 2868 22680 2906
rect 21720 2851 21922 2868
rect 21460 2834 21476 2851
rect 20888 2818 21476 2834
rect 21906 2834 21922 2851
rect 22478 2851 22680 2868
rect 22738 2868 23698 2906
rect 22738 2851 22940 2868
rect 22478 2834 22494 2851
rect 21906 2818 22494 2834
rect 22924 2834 22940 2851
rect 23496 2851 23698 2868
rect 23756 2868 24716 2906
rect 23756 2851 23958 2868
rect 23496 2834 23512 2851
rect 22924 2818 23512 2834
rect 23942 2834 23958 2851
rect 24514 2851 24716 2868
rect 24774 2868 25734 2906
rect 24774 2851 24976 2868
rect 24514 2834 24530 2851
rect 23942 2818 24530 2834
rect 24960 2834 24976 2851
rect 25532 2851 25734 2868
rect 25792 2868 26752 2906
rect 25792 2851 25994 2868
rect 25532 2834 25548 2851
rect 24960 2818 25548 2834
rect 25978 2834 25994 2851
rect 26550 2851 26752 2868
rect 26810 2868 27770 2906
rect 26810 2851 27012 2868
rect 26550 2834 26566 2851
rect 25978 2818 26566 2834
rect 26996 2834 27012 2851
rect 27568 2851 27770 2868
rect 27828 2868 28788 2906
rect 27828 2851 28030 2868
rect 27568 2834 27584 2851
rect 26996 2818 27584 2834
rect 28014 2834 28030 2851
rect 28586 2851 28788 2868
rect 28846 2868 29806 2906
rect 28846 2851 29048 2868
rect 28586 2834 28602 2851
rect 28014 2818 28602 2834
rect 29032 2834 29048 2851
rect 29604 2851 29806 2868
rect 29864 2868 30824 2906
rect 29864 2851 30066 2868
rect 29604 2834 29620 2851
rect 29032 2818 29620 2834
rect 30050 2834 30066 2851
rect 30622 2851 30824 2868
rect 30882 2868 31842 2906
rect 30882 2851 31084 2868
rect 30622 2834 30638 2851
rect 30050 2818 30638 2834
rect 31068 2834 31084 2851
rect 31640 2851 31842 2868
rect 31900 2868 32860 2906
rect 31900 2851 32102 2868
rect 31640 2834 31656 2851
rect 31068 2818 31656 2834
rect 32086 2834 32102 2851
rect 32658 2851 32860 2868
rect 32918 2868 33878 2906
rect 32918 2851 33120 2868
rect 32658 2834 32674 2851
rect 32086 2818 32674 2834
rect 33104 2834 33120 2851
rect 33676 2851 33878 2868
rect 33676 2834 33692 2851
rect 33104 2818 33692 2834
rect 10668 2772 11628 2810
rect 13762 2344 14350 2360
rect 13762 2327 13778 2344
rect 13576 2310 13778 2327
rect 14334 2327 14350 2344
rect 14780 2344 15368 2360
rect 14780 2327 14796 2344
rect 14334 2310 14536 2327
rect 13576 2272 14536 2310
rect 14594 2310 14796 2327
rect 15352 2327 15368 2344
rect 15798 2344 16386 2360
rect 15798 2327 15814 2344
rect 15352 2310 15554 2327
rect 14594 2272 15554 2310
rect 15612 2310 15814 2327
rect 16370 2327 16386 2344
rect 16816 2344 17404 2360
rect 16816 2327 16832 2344
rect 16370 2310 16572 2327
rect 15612 2272 16572 2310
rect 16630 2310 16832 2327
rect 17388 2327 17404 2344
rect 17834 2344 18422 2360
rect 17834 2327 17850 2344
rect 17388 2310 17590 2327
rect 16630 2272 17590 2310
rect 17648 2310 17850 2327
rect 18406 2327 18422 2344
rect 18852 2344 19440 2360
rect 18852 2327 18868 2344
rect 18406 2310 18608 2327
rect 17648 2272 18608 2310
rect 18666 2310 18868 2327
rect 19424 2327 19440 2344
rect 19870 2344 20458 2360
rect 19870 2327 19886 2344
rect 19424 2310 19626 2327
rect 18666 2272 19626 2310
rect 19684 2310 19886 2327
rect 20442 2327 20458 2344
rect 20888 2344 21476 2360
rect 20888 2327 20904 2344
rect 20442 2310 20644 2327
rect 19684 2272 20644 2310
rect 20702 2310 20904 2327
rect 21460 2327 21476 2344
rect 21906 2344 22494 2360
rect 21906 2327 21922 2344
rect 21460 2310 21662 2327
rect 20702 2272 21662 2310
rect 21720 2310 21922 2327
rect 22478 2327 22494 2344
rect 22924 2344 23512 2360
rect 22924 2327 22940 2344
rect 22478 2310 22680 2327
rect 21720 2272 22680 2310
rect 22738 2310 22940 2327
rect 23496 2327 23512 2344
rect 23942 2344 24530 2360
rect 23942 2327 23958 2344
rect 23496 2310 23698 2327
rect 22738 2272 23698 2310
rect 23756 2310 23958 2327
rect 24514 2327 24530 2344
rect 24960 2344 25548 2360
rect 24960 2327 24976 2344
rect 24514 2310 24716 2327
rect 23756 2272 24716 2310
rect 24774 2310 24976 2327
rect 25532 2327 25548 2344
rect 25978 2344 26566 2360
rect 25978 2327 25994 2344
rect 25532 2310 25734 2327
rect 24774 2272 25734 2310
rect 25792 2310 25994 2327
rect 26550 2327 26566 2344
rect 26996 2344 27584 2360
rect 26996 2327 27012 2344
rect 26550 2310 26752 2327
rect 25792 2272 26752 2310
rect 26810 2310 27012 2327
rect 27568 2327 27584 2344
rect 28014 2344 28602 2360
rect 28014 2327 28030 2344
rect 27568 2310 27770 2327
rect 26810 2272 27770 2310
rect 27828 2310 28030 2327
rect 28586 2327 28602 2344
rect 29032 2344 29620 2360
rect 29032 2327 29048 2344
rect 28586 2310 28788 2327
rect 27828 2272 28788 2310
rect 28846 2310 29048 2327
rect 29604 2327 29620 2344
rect 30050 2344 30638 2360
rect 30050 2327 30066 2344
rect 29604 2310 29806 2327
rect 28846 2272 29806 2310
rect 29864 2310 30066 2327
rect 30622 2327 30638 2344
rect 31068 2344 31656 2360
rect 31068 2327 31084 2344
rect 30622 2310 30824 2327
rect 29864 2272 30824 2310
rect 30882 2310 31084 2327
rect 31640 2327 31656 2344
rect 32086 2344 32674 2360
rect 32086 2327 32102 2344
rect 31640 2310 31842 2327
rect 30882 2272 31842 2310
rect 31900 2310 32102 2327
rect 32658 2327 32674 2344
rect 33104 2344 33692 2360
rect 33104 2327 33120 2344
rect 32658 2310 32860 2327
rect 31900 2272 32860 2310
rect 32918 2310 33120 2327
rect 33676 2327 33692 2344
rect 33676 2310 33878 2327
rect 32918 2272 33878 2310
rect 488 2134 1448 2172
rect 488 2117 690 2134
rect 674 2100 690 2117
rect 1246 2117 1448 2134
rect 1506 2134 2466 2172
rect 1506 2117 1708 2134
rect 1246 2100 1262 2117
rect 674 2084 1262 2100
rect 1692 2100 1708 2117
rect 2264 2117 2466 2134
rect 2524 2134 3484 2172
rect 2524 2117 2726 2134
rect 2264 2100 2280 2117
rect 1692 2084 2280 2100
rect 2710 2100 2726 2117
rect 3282 2117 3484 2134
rect 3542 2134 4502 2172
rect 3542 2117 3744 2134
rect 3282 2100 3298 2117
rect 2710 2084 3298 2100
rect 3728 2100 3744 2117
rect 4300 2117 4502 2134
rect 4560 2134 5520 2172
rect 4560 2117 4762 2134
rect 4300 2100 4316 2117
rect 3728 2084 4316 2100
rect 4746 2100 4762 2117
rect 5318 2117 5520 2134
rect 5578 2134 6538 2172
rect 5578 2117 5780 2134
rect 5318 2100 5334 2117
rect 4746 2084 5334 2100
rect 5764 2100 5780 2117
rect 6336 2117 6538 2134
rect 6596 2134 7556 2172
rect 6596 2117 6798 2134
rect 6336 2100 6352 2117
rect 5764 2084 6352 2100
rect 6782 2100 6798 2117
rect 7354 2117 7556 2134
rect 7614 2134 8574 2172
rect 7614 2117 7816 2134
rect 7354 2100 7370 2117
rect 6782 2084 7370 2100
rect 7800 2100 7816 2117
rect 8372 2117 8574 2134
rect 8632 2134 9592 2172
rect 8632 2117 8834 2134
rect 8372 2100 8388 2117
rect 7800 2084 8388 2100
rect 8818 2100 8834 2117
rect 9390 2117 9592 2134
rect 9650 2134 10610 2172
rect 9650 2117 9852 2134
rect 9390 2100 9406 2117
rect 8818 2084 9406 2100
rect 9836 2100 9852 2117
rect 10408 2117 10610 2134
rect 10668 2134 11628 2172
rect 10668 2117 10870 2134
rect 10408 2100 10424 2117
rect 9836 2084 10424 2100
rect 10854 2100 10870 2117
rect 11426 2117 11628 2134
rect 11426 2100 11442 2117
rect 10854 2084 11442 2100
rect 13576 1634 14536 1672
rect 13576 1617 13778 1634
rect 13762 1600 13778 1617
rect 14334 1617 14536 1634
rect 14594 1634 15554 1672
rect 14594 1617 14796 1634
rect 14334 1600 14350 1617
rect 13762 1584 14350 1600
rect 14780 1600 14796 1617
rect 15352 1617 15554 1634
rect 15612 1634 16572 1672
rect 15612 1617 15814 1634
rect 15352 1600 15368 1617
rect 14780 1584 15368 1600
rect 15798 1600 15814 1617
rect 16370 1617 16572 1634
rect 16630 1634 17590 1672
rect 16630 1617 16832 1634
rect 16370 1600 16386 1617
rect 15798 1584 16386 1600
rect 16816 1600 16832 1617
rect 17388 1617 17590 1634
rect 17648 1634 18608 1672
rect 17648 1617 17850 1634
rect 17388 1600 17404 1617
rect 16816 1584 17404 1600
rect 17834 1600 17850 1617
rect 18406 1617 18608 1634
rect 18666 1634 19626 1672
rect 18666 1617 18868 1634
rect 18406 1600 18422 1617
rect 17834 1584 18422 1600
rect 18852 1600 18868 1617
rect 19424 1617 19626 1634
rect 19684 1634 20644 1672
rect 19684 1617 19886 1634
rect 19424 1600 19440 1617
rect 18852 1584 19440 1600
rect 19870 1600 19886 1617
rect 20442 1617 20644 1634
rect 20702 1634 21662 1672
rect 20702 1617 20904 1634
rect 20442 1600 20458 1617
rect 19870 1584 20458 1600
rect 20888 1600 20904 1617
rect 21460 1617 21662 1634
rect 21720 1634 22680 1672
rect 21720 1617 21922 1634
rect 21460 1600 21476 1617
rect 20888 1584 21476 1600
rect 21906 1600 21922 1617
rect 22478 1617 22680 1634
rect 22738 1634 23698 1672
rect 22738 1617 22940 1634
rect 22478 1600 22494 1617
rect 21906 1584 22494 1600
rect 22924 1600 22940 1617
rect 23496 1617 23698 1634
rect 23756 1634 24716 1672
rect 23756 1617 23958 1634
rect 23496 1600 23512 1617
rect 22924 1584 23512 1600
rect 23942 1600 23958 1617
rect 24514 1617 24716 1634
rect 24774 1634 25734 1672
rect 24774 1617 24976 1634
rect 24514 1600 24530 1617
rect 23942 1584 24530 1600
rect 24960 1600 24976 1617
rect 25532 1617 25734 1634
rect 25792 1634 26752 1672
rect 25792 1617 25994 1634
rect 25532 1600 25548 1617
rect 24960 1584 25548 1600
rect 25978 1600 25994 1617
rect 26550 1617 26752 1634
rect 26810 1634 27770 1672
rect 26810 1617 27012 1634
rect 26550 1600 26566 1617
rect 25978 1584 26566 1600
rect 26996 1600 27012 1617
rect 27568 1617 27770 1634
rect 27828 1634 28788 1672
rect 27828 1617 28030 1634
rect 27568 1600 27584 1617
rect 26996 1584 27584 1600
rect 28014 1600 28030 1617
rect 28586 1617 28788 1634
rect 28846 1634 29806 1672
rect 28846 1617 29048 1634
rect 28586 1600 28602 1617
rect 28014 1584 28602 1600
rect 29032 1600 29048 1617
rect 29604 1617 29806 1634
rect 29864 1634 30824 1672
rect 29864 1617 30066 1634
rect 29604 1600 29620 1617
rect 29032 1584 29620 1600
rect 30050 1600 30066 1617
rect 30622 1617 30824 1634
rect 30882 1634 31842 1672
rect 30882 1617 31084 1634
rect 30622 1600 30638 1617
rect 30050 1584 30638 1600
rect 31068 1600 31084 1617
rect 31640 1617 31842 1634
rect 31900 1634 32860 1672
rect 31900 1617 32102 1634
rect 31640 1600 31656 1617
rect 31068 1584 31656 1600
rect 32086 1600 32102 1617
rect 32658 1617 32860 1634
rect 32918 1634 33878 1672
rect 32918 1617 33120 1634
rect 32658 1600 32674 1617
rect 32086 1584 32674 1600
rect 33104 1600 33120 1617
rect 33676 1617 33878 1634
rect 33676 1600 33692 1617
rect 33104 1584 33692 1600
rect 1132 1302 1720 1318
rect 1132 1285 1148 1302
rect 946 1268 1148 1285
rect 1704 1285 1720 1302
rect 2150 1302 2738 1318
rect 2150 1285 2166 1302
rect 1704 1268 1906 1285
rect 946 1230 1906 1268
rect 1964 1268 2166 1285
rect 2722 1285 2738 1302
rect 3168 1302 3756 1318
rect 3168 1285 3184 1302
rect 2722 1268 2924 1285
rect 1964 1230 2924 1268
rect 2982 1268 3184 1285
rect 3740 1285 3756 1302
rect 4186 1302 4774 1318
rect 4186 1285 4202 1302
rect 3740 1268 3942 1285
rect 2982 1230 3942 1268
rect 4000 1268 4202 1285
rect 4758 1285 4774 1302
rect 5204 1302 5792 1318
rect 5204 1285 5220 1302
rect 4758 1268 4960 1285
rect 4000 1230 4960 1268
rect 5018 1268 5220 1285
rect 5776 1285 5792 1302
rect 6222 1302 6810 1318
rect 6222 1285 6238 1302
rect 5776 1268 5978 1285
rect 5018 1230 5978 1268
rect 6036 1268 6238 1285
rect 6794 1285 6810 1302
rect 7240 1302 7828 1318
rect 7240 1285 7256 1302
rect 6794 1268 6996 1285
rect 6036 1230 6996 1268
rect 7054 1268 7256 1285
rect 7812 1285 7828 1302
rect 8258 1302 8846 1318
rect 8258 1285 8274 1302
rect 7812 1268 8014 1285
rect 7054 1230 8014 1268
rect 8072 1268 8274 1285
rect 8830 1285 8846 1302
rect 9276 1302 9864 1318
rect 9276 1285 9292 1302
rect 8830 1268 9032 1285
rect 8072 1230 9032 1268
rect 9090 1268 9292 1285
rect 9848 1285 9864 1302
rect 10294 1302 10882 1318
rect 10294 1285 10310 1302
rect 9848 1268 10050 1285
rect 9090 1230 10050 1268
rect 10108 1268 10310 1285
rect 10866 1285 10882 1302
rect 10866 1268 11068 1285
rect 10108 1230 11068 1268
rect 13762 1112 14350 1128
rect 13762 1095 13778 1112
rect 13576 1078 13778 1095
rect 14334 1095 14350 1112
rect 14780 1112 15368 1128
rect 14780 1095 14796 1112
rect 14334 1078 14536 1095
rect 13576 1040 14536 1078
rect 14594 1078 14796 1095
rect 15352 1095 15368 1112
rect 15798 1112 16386 1128
rect 15798 1095 15814 1112
rect 15352 1078 15554 1095
rect 14594 1040 15554 1078
rect 15612 1078 15814 1095
rect 16370 1095 16386 1112
rect 16816 1112 17404 1128
rect 16816 1095 16832 1112
rect 16370 1078 16572 1095
rect 15612 1040 16572 1078
rect 16630 1078 16832 1095
rect 17388 1095 17404 1112
rect 17834 1112 18422 1128
rect 17834 1095 17850 1112
rect 17388 1078 17590 1095
rect 16630 1040 17590 1078
rect 17648 1078 17850 1095
rect 18406 1095 18422 1112
rect 18852 1112 19440 1128
rect 18852 1095 18868 1112
rect 18406 1078 18608 1095
rect 17648 1040 18608 1078
rect 18666 1078 18868 1095
rect 19424 1095 19440 1112
rect 19870 1112 20458 1128
rect 19870 1095 19886 1112
rect 19424 1078 19626 1095
rect 18666 1040 19626 1078
rect 19684 1078 19886 1095
rect 20442 1095 20458 1112
rect 20888 1112 21476 1128
rect 20888 1095 20904 1112
rect 20442 1078 20644 1095
rect 19684 1040 20644 1078
rect 20702 1078 20904 1095
rect 21460 1095 21476 1112
rect 21906 1112 22494 1128
rect 21906 1095 21922 1112
rect 21460 1078 21662 1095
rect 20702 1040 21662 1078
rect 21720 1078 21922 1095
rect 22478 1095 22494 1112
rect 22924 1112 23512 1128
rect 22924 1095 22940 1112
rect 22478 1078 22680 1095
rect 21720 1040 22680 1078
rect 22738 1078 22940 1095
rect 23496 1095 23512 1112
rect 23942 1112 24530 1128
rect 23942 1095 23958 1112
rect 23496 1078 23698 1095
rect 22738 1040 23698 1078
rect 23756 1078 23958 1095
rect 24514 1095 24530 1112
rect 24960 1112 25548 1128
rect 24960 1095 24976 1112
rect 24514 1078 24716 1095
rect 23756 1040 24716 1078
rect 24774 1078 24976 1095
rect 25532 1095 25548 1112
rect 25978 1112 26566 1128
rect 25978 1095 25994 1112
rect 25532 1078 25734 1095
rect 24774 1040 25734 1078
rect 25792 1078 25994 1095
rect 26550 1095 26566 1112
rect 26996 1112 27584 1128
rect 26996 1095 27012 1112
rect 26550 1078 26752 1095
rect 25792 1040 26752 1078
rect 26810 1078 27012 1095
rect 27568 1095 27584 1112
rect 28014 1112 28602 1128
rect 28014 1095 28030 1112
rect 27568 1078 27770 1095
rect 26810 1040 27770 1078
rect 27828 1078 28030 1095
rect 28586 1095 28602 1112
rect 29032 1112 29620 1128
rect 29032 1095 29048 1112
rect 28586 1078 28788 1095
rect 27828 1040 28788 1078
rect 28846 1078 29048 1095
rect 29604 1095 29620 1112
rect 30050 1112 30638 1128
rect 30050 1095 30066 1112
rect 29604 1078 29806 1095
rect 28846 1040 29806 1078
rect 29864 1078 30066 1095
rect 30622 1095 30638 1112
rect 31068 1112 31656 1128
rect 31068 1095 31084 1112
rect 30622 1078 30824 1095
rect 29864 1040 30824 1078
rect 30882 1078 31084 1095
rect 31640 1095 31656 1112
rect 32086 1112 32674 1128
rect 32086 1095 32102 1112
rect 31640 1078 31842 1095
rect 30882 1040 31842 1078
rect 31900 1078 32102 1095
rect 32658 1095 32674 1112
rect 33104 1112 33692 1128
rect 33104 1095 33120 1112
rect 32658 1078 32860 1095
rect 31900 1040 32860 1078
rect 32918 1078 33120 1095
rect 33676 1095 33692 1112
rect 33676 1078 33878 1095
rect 32918 1040 33878 1078
rect 946 592 1906 630
rect 946 575 1148 592
rect 1132 558 1148 575
rect 1704 575 1906 592
rect 1964 592 2924 630
rect 1964 575 2166 592
rect 1704 558 1720 575
rect 1132 542 1720 558
rect 2150 558 2166 575
rect 2722 575 2924 592
rect 2982 592 3942 630
rect 2982 575 3184 592
rect 2722 558 2738 575
rect 2150 542 2738 558
rect 3168 558 3184 575
rect 3740 575 3942 592
rect 4000 592 4960 630
rect 4000 575 4202 592
rect 3740 558 3756 575
rect 3168 542 3756 558
rect 4186 558 4202 575
rect 4758 575 4960 592
rect 5018 592 5978 630
rect 5018 575 5220 592
rect 4758 558 4774 575
rect 4186 542 4774 558
rect 5204 558 5220 575
rect 5776 575 5978 592
rect 6036 592 6996 630
rect 6036 575 6238 592
rect 5776 558 5792 575
rect 5204 542 5792 558
rect 6222 558 6238 575
rect 6794 575 6996 592
rect 7054 592 8014 630
rect 7054 575 7256 592
rect 6794 558 6810 575
rect 6222 542 6810 558
rect 7240 558 7256 575
rect 7812 575 8014 592
rect 8072 592 9032 630
rect 8072 575 8274 592
rect 7812 558 7828 575
rect 7240 542 7828 558
rect 8258 558 8274 575
rect 8830 575 9032 592
rect 9090 592 10050 630
rect 9090 575 9292 592
rect 8830 558 8846 575
rect 8258 542 8846 558
rect 9276 558 9292 575
rect 9848 575 10050 592
rect 10108 592 11068 630
rect 10108 575 10310 592
rect 9848 558 9864 575
rect 9276 542 9864 558
rect 10294 558 10310 575
rect 10866 575 11068 592
rect 10866 558 10882 575
rect 10294 542 10882 558
rect 13576 402 14536 440
rect 13576 385 13778 402
rect -1046 274 -980 290
rect -1046 240 -1030 274
rect -996 240 -980 274
rect -1046 224 -980 240
rect -1028 202 -998 224
rect 13762 368 13778 385
rect 14334 385 14536 402
rect 14594 402 15554 440
rect 14594 385 14796 402
rect 14334 368 14350 385
rect 13762 352 14350 368
rect 14780 368 14796 385
rect 15352 385 15554 402
rect 15612 402 16572 440
rect 15612 385 15814 402
rect 15352 368 15368 385
rect 14780 352 15368 368
rect 15798 368 15814 385
rect 16370 385 16572 402
rect 16630 402 17590 440
rect 16630 385 16832 402
rect 16370 368 16386 385
rect 15798 352 16386 368
rect 16816 368 16832 385
rect 17388 385 17590 402
rect 17648 402 18608 440
rect 17648 385 17850 402
rect 17388 368 17404 385
rect 16816 352 17404 368
rect 17834 368 17850 385
rect 18406 385 18608 402
rect 18666 402 19626 440
rect 18666 385 18868 402
rect 18406 368 18422 385
rect 17834 352 18422 368
rect 18852 368 18868 385
rect 19424 385 19626 402
rect 19684 402 20644 440
rect 19684 385 19886 402
rect 19424 368 19440 385
rect 18852 352 19440 368
rect 19870 368 19886 385
rect 20442 385 20644 402
rect 20702 402 21662 440
rect 20702 385 20904 402
rect 20442 368 20458 385
rect 19870 352 20458 368
rect 20888 368 20904 385
rect 21460 385 21662 402
rect 21720 402 22680 440
rect 21720 385 21922 402
rect 21460 368 21476 385
rect 20888 352 21476 368
rect 21906 368 21922 385
rect 22478 385 22680 402
rect 22738 402 23698 440
rect 22738 385 22940 402
rect 22478 368 22494 385
rect 21906 352 22494 368
rect 22924 368 22940 385
rect 23496 385 23698 402
rect 23756 402 24716 440
rect 23756 385 23958 402
rect 23496 368 23512 385
rect 22924 352 23512 368
rect 23942 368 23958 385
rect 24514 385 24716 402
rect 24774 402 25734 440
rect 24774 385 24976 402
rect 24514 368 24530 385
rect 23942 352 24530 368
rect 24960 368 24976 385
rect 25532 385 25734 402
rect 25792 402 26752 440
rect 25792 385 25994 402
rect 25532 368 25548 385
rect 24960 352 25548 368
rect 25978 368 25994 385
rect 26550 385 26752 402
rect 26810 402 27770 440
rect 26810 385 27012 402
rect 26550 368 26566 385
rect 25978 352 26566 368
rect 26996 368 27012 385
rect 27568 385 27770 402
rect 27828 402 28788 440
rect 27828 385 28030 402
rect 27568 368 27584 385
rect 26996 352 27584 368
rect 28014 368 28030 385
rect 28586 385 28788 402
rect 28846 402 29806 440
rect 28846 385 29048 402
rect 28586 368 28602 385
rect 28014 352 28602 368
rect 29032 368 29048 385
rect 29604 385 29806 402
rect 29864 402 30824 440
rect 29864 385 30066 402
rect 29604 368 29620 385
rect 29032 352 29620 368
rect 30050 368 30066 385
rect 30622 385 30824 402
rect 30882 402 31842 440
rect 30882 385 31084 402
rect 30622 368 30638 385
rect 30050 352 30638 368
rect 31068 368 31084 385
rect 31640 385 31842 402
rect 31900 402 32860 440
rect 31900 385 32102 402
rect 31640 368 31656 385
rect 31068 352 31656 368
rect 32086 368 32102 385
rect 32658 385 32860 402
rect 32918 402 33878 440
rect 32918 385 33120 402
rect 32658 368 32674 385
rect 32086 352 32674 368
rect 33104 368 33120 385
rect 33676 385 33878 402
rect 33676 368 33692 385
rect 33104 352 33692 368
rect -1028 50 -998 72
rect -1046 34 -980 50
rect -1046 0 -1030 34
rect -996 0 -980 34
rect -1046 -16 -980 0
rect 36990 13079 37122 13095
rect 36990 13062 37006 13079
rect 36956 13045 37006 13062
rect 37106 13062 37122 13079
rect 37248 13079 37380 13095
rect 37248 13062 37264 13079
rect 37106 13045 37156 13062
rect 36956 12998 37156 13045
rect 37214 13045 37264 13062
rect 37364 13062 37380 13079
rect 37506 13079 37638 13095
rect 37506 13062 37522 13079
rect 37364 13045 37414 13062
rect 37214 12998 37414 13045
rect 37472 13045 37522 13062
rect 37622 13062 37638 13079
rect 37764 13079 37896 13095
rect 37764 13062 37780 13079
rect 37622 13045 37672 13062
rect 37472 12998 37672 13045
rect 37730 13045 37780 13062
rect 37880 13062 37896 13079
rect 38022 13079 38154 13095
rect 38022 13062 38038 13079
rect 37880 13045 37930 13062
rect 37730 12998 37930 13045
rect 37988 13045 38038 13062
rect 38138 13062 38154 13079
rect 38280 13079 38412 13095
rect 38280 13062 38296 13079
rect 38138 13045 38188 13062
rect 37988 12998 38188 13045
rect 38246 13045 38296 13062
rect 38396 13062 38412 13079
rect 38396 13045 38446 13062
rect 38246 12998 38446 13045
rect 36956 12751 37156 12798
rect 36956 12734 37006 12751
rect 36990 12717 37006 12734
rect 37106 12734 37156 12751
rect 37214 12751 37414 12798
rect 37214 12734 37264 12751
rect 37106 12717 37122 12734
rect 36990 12701 37122 12717
rect 37248 12717 37264 12734
rect 37364 12734 37414 12751
rect 37472 12751 37672 12798
rect 37472 12734 37522 12751
rect 37364 12717 37380 12734
rect 37248 12701 37380 12717
rect 37506 12717 37522 12734
rect 37622 12734 37672 12751
rect 37730 12751 37930 12798
rect 37730 12734 37780 12751
rect 37622 12717 37638 12734
rect 37506 12701 37638 12717
rect 37764 12717 37780 12734
rect 37880 12734 37930 12751
rect 37988 12751 38188 12798
rect 37988 12734 38038 12751
rect 37880 12717 37896 12734
rect 37764 12701 37896 12717
rect 38022 12717 38038 12734
rect 38138 12734 38188 12751
rect 38246 12751 38446 12798
rect 38246 12734 38296 12751
rect 38138 12717 38154 12734
rect 38022 12701 38154 12717
rect 38280 12717 38296 12734
rect 38396 12734 38446 12751
rect 38396 12717 38412 12734
rect 38280 12701 38412 12717
rect 54764 14406 55352 14422
rect 54764 14389 54780 14406
rect 54578 14372 54780 14389
rect 55336 14389 55352 14406
rect 55782 14406 56370 14422
rect 55782 14389 55798 14406
rect 55336 14372 55538 14389
rect 54578 14334 55538 14372
rect 55596 14372 55798 14389
rect 56354 14389 56370 14406
rect 56800 14406 57388 14422
rect 56800 14389 56816 14406
rect 56354 14372 56556 14389
rect 55596 14334 56556 14372
rect 56614 14372 56816 14389
rect 57372 14389 57388 14406
rect 57818 14406 58406 14422
rect 57818 14389 57834 14406
rect 57372 14372 57574 14389
rect 56614 14334 57574 14372
rect 57632 14372 57834 14389
rect 58390 14389 58406 14406
rect 58836 14406 59424 14422
rect 58836 14389 58852 14406
rect 58390 14372 58592 14389
rect 57632 14334 58592 14372
rect 58650 14372 58852 14389
rect 59408 14389 59424 14406
rect 59854 14406 60442 14422
rect 59854 14389 59870 14406
rect 59408 14372 59610 14389
rect 58650 14334 59610 14372
rect 59668 14372 59870 14389
rect 60426 14389 60442 14406
rect 60872 14406 61460 14422
rect 60872 14389 60888 14406
rect 60426 14372 60628 14389
rect 59668 14334 60628 14372
rect 60686 14372 60888 14389
rect 61444 14389 61460 14406
rect 61890 14406 62478 14422
rect 61890 14389 61906 14406
rect 61444 14372 61646 14389
rect 60686 14334 61646 14372
rect 61704 14372 61906 14389
rect 62462 14389 62478 14406
rect 62908 14406 63496 14422
rect 62908 14389 62924 14406
rect 62462 14372 62664 14389
rect 61704 14334 62664 14372
rect 62722 14372 62924 14389
rect 63480 14389 63496 14406
rect 63926 14406 64514 14422
rect 63926 14389 63942 14406
rect 63480 14372 63682 14389
rect 62722 14334 63682 14372
rect 63740 14372 63942 14389
rect 64498 14389 64514 14406
rect 64944 14406 65532 14422
rect 64944 14389 64960 14406
rect 64498 14372 64700 14389
rect 63740 14334 64700 14372
rect 64758 14372 64960 14389
rect 65516 14389 65532 14406
rect 65962 14406 66550 14422
rect 65962 14389 65978 14406
rect 65516 14372 65718 14389
rect 64758 14334 65718 14372
rect 65776 14372 65978 14389
rect 66534 14389 66550 14406
rect 66980 14406 67568 14422
rect 66980 14389 66996 14406
rect 66534 14372 66736 14389
rect 65776 14334 66736 14372
rect 66794 14372 66996 14389
rect 67552 14389 67568 14406
rect 67998 14406 68586 14422
rect 67998 14389 68014 14406
rect 67552 14372 67754 14389
rect 66794 14334 67754 14372
rect 67812 14372 68014 14389
rect 68570 14389 68586 14406
rect 69016 14406 69604 14422
rect 69016 14389 69032 14406
rect 68570 14372 68772 14389
rect 67812 14334 68772 14372
rect 68830 14372 69032 14389
rect 69588 14389 69604 14406
rect 70034 14406 70622 14422
rect 70034 14389 70050 14406
rect 69588 14372 69790 14389
rect 68830 14334 69790 14372
rect 69848 14372 70050 14389
rect 70606 14389 70622 14406
rect 71052 14406 71640 14422
rect 71052 14389 71068 14406
rect 70606 14372 70808 14389
rect 69848 14334 70808 14372
rect 70866 14372 71068 14389
rect 71624 14389 71640 14406
rect 72070 14406 72658 14422
rect 72070 14389 72086 14406
rect 71624 14372 71826 14389
rect 70866 14334 71826 14372
rect 71884 14372 72086 14389
rect 72642 14389 72658 14406
rect 73088 14406 73676 14422
rect 73088 14389 73104 14406
rect 72642 14372 72844 14389
rect 71884 14334 72844 14372
rect 72902 14372 73104 14389
rect 73660 14389 73676 14406
rect 74106 14406 74694 14422
rect 74106 14389 74122 14406
rect 73660 14372 73862 14389
rect 72902 14334 73862 14372
rect 73920 14372 74122 14389
rect 74678 14389 74694 14406
rect 74678 14372 74880 14389
rect 73920 14334 74880 14372
rect 42998 13930 43586 13946
rect 42998 13913 43014 13930
rect 42812 13896 43014 13913
rect 43570 13913 43586 13930
rect 44016 13930 44604 13946
rect 44016 13913 44032 13930
rect 43570 13896 43772 13913
rect 42812 13858 43772 13896
rect 43830 13896 44032 13913
rect 44588 13913 44604 13930
rect 45034 13930 45622 13946
rect 45034 13913 45050 13930
rect 44588 13896 44790 13913
rect 43830 13858 44790 13896
rect 44848 13896 45050 13913
rect 45606 13913 45622 13930
rect 46052 13930 46640 13946
rect 46052 13913 46068 13930
rect 45606 13896 45808 13913
rect 44848 13858 45808 13896
rect 45866 13896 46068 13913
rect 46624 13913 46640 13930
rect 47070 13930 47658 13946
rect 47070 13913 47086 13930
rect 46624 13896 46826 13913
rect 45866 13858 46826 13896
rect 46884 13896 47086 13913
rect 47642 13913 47658 13930
rect 48088 13930 48676 13946
rect 48088 13913 48104 13930
rect 47642 13896 47844 13913
rect 46884 13858 47844 13896
rect 47902 13896 48104 13913
rect 48660 13913 48676 13930
rect 49106 13930 49694 13946
rect 49106 13913 49122 13930
rect 48660 13896 48862 13913
rect 47902 13858 48862 13896
rect 48920 13896 49122 13913
rect 49678 13913 49694 13930
rect 50124 13930 50712 13946
rect 50124 13913 50140 13930
rect 49678 13896 49880 13913
rect 48920 13858 49880 13896
rect 49938 13896 50140 13913
rect 50696 13913 50712 13930
rect 51142 13930 51730 13946
rect 51142 13913 51158 13930
rect 50696 13896 50898 13913
rect 49938 13858 50898 13896
rect 50956 13896 51158 13913
rect 51714 13913 51730 13930
rect 51714 13896 51916 13913
rect 50956 13858 51916 13896
rect 54578 13696 55538 13734
rect 54578 13679 54780 13696
rect 54764 13662 54780 13679
rect 55336 13679 55538 13696
rect 55596 13696 56556 13734
rect 55596 13679 55798 13696
rect 55336 13662 55352 13679
rect 54764 13646 55352 13662
rect 55782 13662 55798 13679
rect 56354 13679 56556 13696
rect 56614 13696 57574 13734
rect 56614 13679 56816 13696
rect 56354 13662 56370 13679
rect 55782 13646 56370 13662
rect 56800 13662 56816 13679
rect 57372 13679 57574 13696
rect 57632 13696 58592 13734
rect 57632 13679 57834 13696
rect 57372 13662 57388 13679
rect 56800 13646 57388 13662
rect 57818 13662 57834 13679
rect 58390 13679 58592 13696
rect 58650 13696 59610 13734
rect 58650 13679 58852 13696
rect 58390 13662 58406 13679
rect 57818 13646 58406 13662
rect 58836 13662 58852 13679
rect 59408 13679 59610 13696
rect 59668 13696 60628 13734
rect 59668 13679 59870 13696
rect 59408 13662 59424 13679
rect 58836 13646 59424 13662
rect 59854 13662 59870 13679
rect 60426 13679 60628 13696
rect 60686 13696 61646 13734
rect 60686 13679 60888 13696
rect 60426 13662 60442 13679
rect 59854 13646 60442 13662
rect 60872 13662 60888 13679
rect 61444 13679 61646 13696
rect 61704 13696 62664 13734
rect 61704 13679 61906 13696
rect 61444 13662 61460 13679
rect 60872 13646 61460 13662
rect 61890 13662 61906 13679
rect 62462 13679 62664 13696
rect 62722 13696 63682 13734
rect 62722 13679 62924 13696
rect 62462 13662 62478 13679
rect 61890 13646 62478 13662
rect 62908 13662 62924 13679
rect 63480 13679 63682 13696
rect 63740 13696 64700 13734
rect 63740 13679 63942 13696
rect 63480 13662 63496 13679
rect 62908 13646 63496 13662
rect 63926 13662 63942 13679
rect 64498 13679 64700 13696
rect 64758 13696 65718 13734
rect 64758 13679 64960 13696
rect 64498 13662 64514 13679
rect 63926 13646 64514 13662
rect 64944 13662 64960 13679
rect 65516 13679 65718 13696
rect 65776 13696 66736 13734
rect 65776 13679 65978 13696
rect 65516 13662 65532 13679
rect 64944 13646 65532 13662
rect 65962 13662 65978 13679
rect 66534 13679 66736 13696
rect 66794 13696 67754 13734
rect 66794 13679 66996 13696
rect 66534 13662 66550 13679
rect 65962 13646 66550 13662
rect 66980 13662 66996 13679
rect 67552 13679 67754 13696
rect 67812 13696 68772 13734
rect 67812 13679 68014 13696
rect 67552 13662 67568 13679
rect 66980 13646 67568 13662
rect 67998 13662 68014 13679
rect 68570 13679 68772 13696
rect 68830 13696 69790 13734
rect 68830 13679 69032 13696
rect 68570 13662 68586 13679
rect 67998 13646 68586 13662
rect 69016 13662 69032 13679
rect 69588 13679 69790 13696
rect 69848 13696 70808 13734
rect 69848 13679 70050 13696
rect 69588 13662 69604 13679
rect 69016 13646 69604 13662
rect 70034 13662 70050 13679
rect 70606 13679 70808 13696
rect 70866 13696 71826 13734
rect 70866 13679 71068 13696
rect 70606 13662 70622 13679
rect 70034 13646 70622 13662
rect 71052 13662 71068 13679
rect 71624 13679 71826 13696
rect 71884 13696 72844 13734
rect 71884 13679 72086 13696
rect 71624 13662 71640 13679
rect 71052 13646 71640 13662
rect 72070 13662 72086 13679
rect 72642 13679 72844 13696
rect 72902 13696 73862 13734
rect 72902 13679 73104 13696
rect 72642 13662 72658 13679
rect 72070 13646 72658 13662
rect 73088 13662 73104 13679
rect 73660 13679 73862 13696
rect 73920 13696 74880 13734
rect 73920 13679 74122 13696
rect 73660 13662 73676 13679
rect 73088 13646 73676 13662
rect 74106 13662 74122 13679
rect 74678 13679 74880 13696
rect 74678 13662 74694 13679
rect 74106 13646 74694 13662
rect 54764 13588 55352 13604
rect 54764 13571 54780 13588
rect 54578 13554 54780 13571
rect 55336 13571 55352 13588
rect 55782 13588 56370 13604
rect 55782 13571 55798 13588
rect 55336 13554 55538 13571
rect 54578 13516 55538 13554
rect 55596 13554 55798 13571
rect 56354 13571 56370 13588
rect 56800 13588 57388 13604
rect 56800 13571 56816 13588
rect 56354 13554 56556 13571
rect 55596 13516 56556 13554
rect 56614 13554 56816 13571
rect 57372 13571 57388 13588
rect 57818 13588 58406 13604
rect 57818 13571 57834 13588
rect 57372 13554 57574 13571
rect 56614 13516 57574 13554
rect 57632 13554 57834 13571
rect 58390 13571 58406 13588
rect 58836 13588 59424 13604
rect 58836 13571 58852 13588
rect 58390 13554 58592 13571
rect 57632 13516 58592 13554
rect 58650 13554 58852 13571
rect 59408 13571 59424 13588
rect 59854 13588 60442 13604
rect 59854 13571 59870 13588
rect 59408 13554 59610 13571
rect 58650 13516 59610 13554
rect 59668 13554 59870 13571
rect 60426 13571 60442 13588
rect 60872 13588 61460 13604
rect 60872 13571 60888 13588
rect 60426 13554 60628 13571
rect 59668 13516 60628 13554
rect 60686 13554 60888 13571
rect 61444 13571 61460 13588
rect 61890 13588 62478 13604
rect 61890 13571 61906 13588
rect 61444 13554 61646 13571
rect 60686 13516 61646 13554
rect 61704 13554 61906 13571
rect 62462 13571 62478 13588
rect 62908 13588 63496 13604
rect 62908 13571 62924 13588
rect 62462 13554 62664 13571
rect 61704 13516 62664 13554
rect 62722 13554 62924 13571
rect 63480 13571 63496 13588
rect 63926 13588 64514 13604
rect 63926 13571 63942 13588
rect 63480 13554 63682 13571
rect 62722 13516 63682 13554
rect 63740 13554 63942 13571
rect 64498 13571 64514 13588
rect 64944 13588 65532 13604
rect 64944 13571 64960 13588
rect 64498 13554 64700 13571
rect 63740 13516 64700 13554
rect 64758 13554 64960 13571
rect 65516 13571 65532 13588
rect 65962 13588 66550 13604
rect 65962 13571 65978 13588
rect 65516 13554 65718 13571
rect 64758 13516 65718 13554
rect 65776 13554 65978 13571
rect 66534 13571 66550 13588
rect 66980 13588 67568 13604
rect 66980 13571 66996 13588
rect 66534 13554 66736 13571
rect 65776 13516 66736 13554
rect 66794 13554 66996 13571
rect 67552 13571 67568 13588
rect 67998 13588 68586 13604
rect 67998 13571 68014 13588
rect 67552 13554 67754 13571
rect 66794 13516 67754 13554
rect 67812 13554 68014 13571
rect 68570 13571 68586 13588
rect 69016 13588 69604 13604
rect 69016 13571 69032 13588
rect 68570 13554 68772 13571
rect 67812 13516 68772 13554
rect 68830 13554 69032 13571
rect 69588 13571 69604 13588
rect 70034 13588 70622 13604
rect 70034 13571 70050 13588
rect 69588 13554 69790 13571
rect 68830 13516 69790 13554
rect 69848 13554 70050 13571
rect 70606 13571 70622 13588
rect 71052 13588 71640 13604
rect 71052 13571 71068 13588
rect 70606 13554 70808 13571
rect 69848 13516 70808 13554
rect 70866 13554 71068 13571
rect 71624 13571 71640 13588
rect 72070 13588 72658 13604
rect 72070 13571 72086 13588
rect 71624 13554 71826 13571
rect 70866 13516 71826 13554
rect 71884 13554 72086 13571
rect 72642 13571 72658 13588
rect 73088 13588 73676 13604
rect 73088 13571 73104 13588
rect 72642 13554 72844 13571
rect 71884 13516 72844 13554
rect 72902 13554 73104 13571
rect 73660 13571 73676 13588
rect 74106 13588 74694 13604
rect 74106 13571 74122 13588
rect 73660 13554 73862 13571
rect 72902 13516 73862 13554
rect 73920 13554 74122 13571
rect 74678 13571 74694 13588
rect 74678 13554 74880 13571
rect 73920 13516 74880 13554
rect 42812 13220 43772 13258
rect 42812 13203 43014 13220
rect 42998 13186 43014 13203
rect 43570 13203 43772 13220
rect 43830 13220 44790 13258
rect 43830 13203 44032 13220
rect 43570 13186 43586 13203
rect 42998 13170 43586 13186
rect 44016 13186 44032 13203
rect 44588 13203 44790 13220
rect 44848 13220 45808 13258
rect 44848 13203 45050 13220
rect 44588 13186 44604 13203
rect 44016 13170 44604 13186
rect 42998 13112 43586 13128
rect 42998 13095 43014 13112
rect 42812 13078 43014 13095
rect 43570 13095 43586 13112
rect 45034 13186 45050 13203
rect 45606 13203 45808 13220
rect 45866 13220 46826 13258
rect 45866 13203 46068 13220
rect 45606 13186 45622 13203
rect 45034 13170 45622 13186
rect 44016 13112 44604 13128
rect 44016 13095 44032 13112
rect 43570 13078 43772 13095
rect 42812 13040 43772 13078
rect 43830 13078 44032 13095
rect 44588 13095 44604 13112
rect 46052 13186 46068 13203
rect 46624 13203 46826 13220
rect 46884 13220 47844 13258
rect 46884 13203 47086 13220
rect 46624 13186 46640 13203
rect 46052 13170 46640 13186
rect 45034 13112 45622 13128
rect 45034 13095 45050 13112
rect 44588 13078 44790 13095
rect 43830 13040 44790 13078
rect 44848 13078 45050 13095
rect 45606 13095 45622 13112
rect 47070 13186 47086 13203
rect 47642 13203 47844 13220
rect 47902 13220 48862 13258
rect 47902 13203 48104 13220
rect 47642 13186 47658 13203
rect 47070 13170 47658 13186
rect 46052 13112 46640 13128
rect 46052 13095 46068 13112
rect 45606 13078 45808 13095
rect 44848 13040 45808 13078
rect 45866 13078 46068 13095
rect 46624 13095 46640 13112
rect 48088 13186 48104 13203
rect 48660 13203 48862 13220
rect 48920 13220 49880 13258
rect 48920 13203 49122 13220
rect 48660 13186 48676 13203
rect 48088 13170 48676 13186
rect 47070 13112 47658 13128
rect 47070 13095 47086 13112
rect 46624 13078 46826 13095
rect 45866 13040 46826 13078
rect 46884 13078 47086 13095
rect 47642 13095 47658 13112
rect 49106 13186 49122 13203
rect 49678 13203 49880 13220
rect 49938 13220 50898 13258
rect 49938 13203 50140 13220
rect 49678 13186 49694 13203
rect 49106 13170 49694 13186
rect 48088 13112 48676 13128
rect 48088 13095 48104 13112
rect 47642 13078 47844 13095
rect 46884 13040 47844 13078
rect 47902 13078 48104 13095
rect 48660 13095 48676 13112
rect 50124 13186 50140 13203
rect 50696 13203 50898 13220
rect 50956 13220 51916 13258
rect 50956 13203 51158 13220
rect 50696 13186 50712 13203
rect 50124 13170 50712 13186
rect 49106 13112 49694 13128
rect 49106 13095 49122 13112
rect 48660 13078 48862 13095
rect 47902 13040 48862 13078
rect 48920 13078 49122 13095
rect 49678 13095 49694 13112
rect 51142 13186 51158 13203
rect 51714 13203 51916 13220
rect 51714 13186 51730 13203
rect 51142 13170 51730 13186
rect 50124 13112 50712 13128
rect 50124 13095 50140 13112
rect 49678 13078 49880 13095
rect 48920 13040 49880 13078
rect 49938 13078 50140 13095
rect 50696 13095 50712 13112
rect 51142 13112 51730 13128
rect 51142 13095 51158 13112
rect 50696 13078 50898 13095
rect 49938 13040 50898 13078
rect 50956 13078 51158 13095
rect 51714 13095 51730 13112
rect 51714 13078 51916 13095
rect 50956 13040 51916 13078
rect 54578 12878 55538 12916
rect 54578 12861 54780 12878
rect 54764 12844 54780 12861
rect 55336 12861 55538 12878
rect 55596 12878 56556 12916
rect 55596 12861 55798 12878
rect 55336 12844 55352 12861
rect 54764 12828 55352 12844
rect 55782 12844 55798 12861
rect 56354 12861 56556 12878
rect 56614 12878 57574 12916
rect 56614 12861 56816 12878
rect 56354 12844 56370 12861
rect 55782 12828 56370 12844
rect 56800 12844 56816 12861
rect 57372 12861 57574 12878
rect 57632 12878 58592 12916
rect 57632 12861 57834 12878
rect 57372 12844 57388 12861
rect 56800 12828 57388 12844
rect 57818 12844 57834 12861
rect 58390 12861 58592 12878
rect 58650 12878 59610 12916
rect 58650 12861 58852 12878
rect 58390 12844 58406 12861
rect 57818 12828 58406 12844
rect 58836 12844 58852 12861
rect 59408 12861 59610 12878
rect 59668 12878 60628 12916
rect 59668 12861 59870 12878
rect 59408 12844 59424 12861
rect 58836 12828 59424 12844
rect 59854 12844 59870 12861
rect 60426 12861 60628 12878
rect 60686 12878 61646 12916
rect 60686 12861 60888 12878
rect 60426 12844 60442 12861
rect 59854 12828 60442 12844
rect 60872 12844 60888 12861
rect 61444 12861 61646 12878
rect 61704 12878 62664 12916
rect 61704 12861 61906 12878
rect 61444 12844 61460 12861
rect 60872 12828 61460 12844
rect 61890 12844 61906 12861
rect 62462 12861 62664 12878
rect 62722 12878 63682 12916
rect 62722 12861 62924 12878
rect 62462 12844 62478 12861
rect 61890 12828 62478 12844
rect 62908 12844 62924 12861
rect 63480 12861 63682 12878
rect 63740 12878 64700 12916
rect 63740 12861 63942 12878
rect 63480 12844 63496 12861
rect 62908 12828 63496 12844
rect 63926 12844 63942 12861
rect 64498 12861 64700 12878
rect 64758 12878 65718 12916
rect 64758 12861 64960 12878
rect 64498 12844 64514 12861
rect 63926 12828 64514 12844
rect 64944 12844 64960 12861
rect 65516 12861 65718 12878
rect 65776 12878 66736 12916
rect 65776 12861 65978 12878
rect 65516 12844 65532 12861
rect 64944 12828 65532 12844
rect 65962 12844 65978 12861
rect 66534 12861 66736 12878
rect 66794 12878 67754 12916
rect 66794 12861 66996 12878
rect 66534 12844 66550 12861
rect 65962 12828 66550 12844
rect 66980 12844 66996 12861
rect 67552 12861 67754 12878
rect 67812 12878 68772 12916
rect 67812 12861 68014 12878
rect 67552 12844 67568 12861
rect 66980 12828 67568 12844
rect 67998 12844 68014 12861
rect 68570 12861 68772 12878
rect 68830 12878 69790 12916
rect 68830 12861 69032 12878
rect 68570 12844 68586 12861
rect 67998 12828 68586 12844
rect 69016 12844 69032 12861
rect 69588 12861 69790 12878
rect 69848 12878 70808 12916
rect 69848 12861 70050 12878
rect 69588 12844 69604 12861
rect 69016 12828 69604 12844
rect 70034 12844 70050 12861
rect 70606 12861 70808 12878
rect 70866 12878 71826 12916
rect 70866 12861 71068 12878
rect 70606 12844 70622 12861
rect 70034 12828 70622 12844
rect 71052 12844 71068 12861
rect 71624 12861 71826 12878
rect 71884 12878 72844 12916
rect 71884 12861 72086 12878
rect 71624 12844 71640 12861
rect 71052 12828 71640 12844
rect 72070 12844 72086 12861
rect 72642 12861 72844 12878
rect 72902 12878 73862 12916
rect 72902 12861 73104 12878
rect 72642 12844 72658 12861
rect 72070 12828 72658 12844
rect 73088 12844 73104 12861
rect 73660 12861 73862 12878
rect 73920 12878 74880 12916
rect 73920 12861 74122 12878
rect 73660 12844 73676 12861
rect 73088 12828 73676 12844
rect 74106 12844 74122 12861
rect 74678 12861 74880 12878
rect 74678 12844 74694 12861
rect 74106 12828 74694 12844
rect 42812 12402 43772 12440
rect 42812 12385 43014 12402
rect 42998 12368 43014 12385
rect 43570 12385 43772 12402
rect 43830 12402 44790 12440
rect 43830 12385 44032 12402
rect 43570 12368 43586 12385
rect 42998 12352 43586 12368
rect 44016 12368 44032 12385
rect 44588 12385 44790 12402
rect 44848 12402 45808 12440
rect 44848 12385 45050 12402
rect 44588 12368 44604 12385
rect 44016 12352 44604 12368
rect 42998 12294 43586 12310
rect 42998 12277 43014 12294
rect 42812 12260 43014 12277
rect 43570 12277 43586 12294
rect 45034 12368 45050 12385
rect 45606 12385 45808 12402
rect 45866 12402 46826 12440
rect 45866 12385 46068 12402
rect 45606 12368 45622 12385
rect 45034 12352 45622 12368
rect 44016 12294 44604 12310
rect 44016 12277 44032 12294
rect 43570 12260 43772 12277
rect 42812 12222 43772 12260
rect 43830 12260 44032 12277
rect 44588 12277 44604 12294
rect 46052 12368 46068 12385
rect 46624 12385 46826 12402
rect 46884 12402 47844 12440
rect 46884 12385 47086 12402
rect 46624 12368 46640 12385
rect 46052 12352 46640 12368
rect 45034 12294 45622 12310
rect 45034 12277 45050 12294
rect 44588 12260 44790 12277
rect 43830 12222 44790 12260
rect 44848 12260 45050 12277
rect 45606 12277 45622 12294
rect 47070 12368 47086 12385
rect 47642 12385 47844 12402
rect 47902 12402 48862 12440
rect 47902 12385 48104 12402
rect 47642 12368 47658 12385
rect 47070 12352 47658 12368
rect 46052 12294 46640 12310
rect 46052 12277 46068 12294
rect 45606 12260 45808 12277
rect 44848 12222 45808 12260
rect 45866 12260 46068 12277
rect 46624 12277 46640 12294
rect 48088 12368 48104 12385
rect 48660 12385 48862 12402
rect 48920 12402 49880 12440
rect 48920 12385 49122 12402
rect 48660 12368 48676 12385
rect 48088 12352 48676 12368
rect 47070 12294 47658 12310
rect 47070 12277 47086 12294
rect 46624 12260 46826 12277
rect 45866 12222 46826 12260
rect 46884 12260 47086 12277
rect 47642 12277 47658 12294
rect 49106 12368 49122 12385
rect 49678 12385 49880 12402
rect 49938 12402 50898 12440
rect 49938 12385 50140 12402
rect 49678 12368 49694 12385
rect 49106 12352 49694 12368
rect 48088 12294 48676 12310
rect 48088 12277 48104 12294
rect 47642 12260 47844 12277
rect 46884 12222 47844 12260
rect 47902 12260 48104 12277
rect 48660 12277 48676 12294
rect 50124 12368 50140 12385
rect 50696 12385 50898 12402
rect 50956 12402 51916 12440
rect 50956 12385 51158 12402
rect 50696 12368 50712 12385
rect 50124 12352 50712 12368
rect 49106 12294 49694 12310
rect 49106 12277 49122 12294
rect 48660 12260 48862 12277
rect 47902 12222 48862 12260
rect 48920 12260 49122 12277
rect 49678 12277 49694 12294
rect 51142 12368 51158 12385
rect 51714 12385 51916 12402
rect 51714 12368 51730 12385
rect 51142 12352 51730 12368
rect 50124 12294 50712 12310
rect 50124 12277 50140 12294
rect 49678 12260 49880 12277
rect 48920 12222 49880 12260
rect 49938 12260 50140 12277
rect 50696 12277 50712 12294
rect 51142 12294 51730 12310
rect 51142 12277 51158 12294
rect 50696 12260 50898 12277
rect 49938 12222 50898 12260
rect 50956 12260 51158 12277
rect 51714 12277 51730 12294
rect 51714 12260 51916 12277
rect 50956 12222 51916 12260
rect 54764 12210 55352 12226
rect 54764 12193 54780 12210
rect 54578 12176 54780 12193
rect 55336 12193 55352 12210
rect 55782 12210 56370 12226
rect 55782 12193 55798 12210
rect 55336 12176 55538 12193
rect 54578 12138 55538 12176
rect 55596 12176 55798 12193
rect 56354 12193 56370 12210
rect 56800 12210 57388 12226
rect 56800 12193 56816 12210
rect 56354 12176 56556 12193
rect 55596 12138 56556 12176
rect 56614 12176 56816 12193
rect 57372 12193 57388 12210
rect 57818 12210 58406 12226
rect 57818 12193 57834 12210
rect 57372 12176 57574 12193
rect 56614 12138 57574 12176
rect 57632 12176 57834 12193
rect 58390 12193 58406 12210
rect 58836 12210 59424 12226
rect 58836 12193 58852 12210
rect 58390 12176 58592 12193
rect 57632 12138 58592 12176
rect 58650 12176 58852 12193
rect 59408 12193 59424 12210
rect 59854 12210 60442 12226
rect 59854 12193 59870 12210
rect 59408 12176 59610 12193
rect 58650 12138 59610 12176
rect 59668 12176 59870 12193
rect 60426 12193 60442 12210
rect 60872 12210 61460 12226
rect 60872 12193 60888 12210
rect 60426 12176 60628 12193
rect 59668 12138 60628 12176
rect 60686 12176 60888 12193
rect 61444 12193 61460 12210
rect 61890 12210 62478 12226
rect 61890 12193 61906 12210
rect 61444 12176 61646 12193
rect 60686 12138 61646 12176
rect 61704 12176 61906 12193
rect 62462 12193 62478 12210
rect 62908 12210 63496 12226
rect 62908 12193 62924 12210
rect 62462 12176 62664 12193
rect 61704 12138 62664 12176
rect 62722 12176 62924 12193
rect 63480 12193 63496 12210
rect 63926 12210 64514 12226
rect 63926 12193 63942 12210
rect 63480 12176 63682 12193
rect 62722 12138 63682 12176
rect 63740 12176 63942 12193
rect 64498 12193 64514 12210
rect 64944 12210 65532 12226
rect 64944 12193 64960 12210
rect 64498 12176 64700 12193
rect 63740 12138 64700 12176
rect 64758 12176 64960 12193
rect 65516 12193 65532 12210
rect 65962 12210 66550 12226
rect 65962 12193 65978 12210
rect 65516 12176 65718 12193
rect 64758 12138 65718 12176
rect 65776 12176 65978 12193
rect 66534 12193 66550 12210
rect 66980 12210 67568 12226
rect 66980 12193 66996 12210
rect 66534 12176 66736 12193
rect 65776 12138 66736 12176
rect 66794 12176 66996 12193
rect 67552 12193 67568 12210
rect 67998 12210 68586 12226
rect 67998 12193 68014 12210
rect 67552 12176 67754 12193
rect 66794 12138 67754 12176
rect 67812 12176 68014 12193
rect 68570 12193 68586 12210
rect 69016 12210 69604 12226
rect 69016 12193 69032 12210
rect 68570 12176 68772 12193
rect 67812 12138 68772 12176
rect 68830 12176 69032 12193
rect 69588 12193 69604 12210
rect 70034 12210 70622 12226
rect 70034 12193 70050 12210
rect 69588 12176 69790 12193
rect 68830 12138 69790 12176
rect 69848 12176 70050 12193
rect 70606 12193 70622 12210
rect 71052 12210 71640 12226
rect 71052 12193 71068 12210
rect 70606 12176 70808 12193
rect 69848 12138 70808 12176
rect 70866 12176 71068 12193
rect 71624 12193 71640 12210
rect 72070 12210 72658 12226
rect 72070 12193 72086 12210
rect 71624 12176 71826 12193
rect 70866 12138 71826 12176
rect 71884 12176 72086 12193
rect 72642 12193 72658 12210
rect 73088 12210 73676 12226
rect 73088 12193 73104 12210
rect 72642 12176 72844 12193
rect 71884 12138 72844 12176
rect 72902 12176 73104 12193
rect 73660 12193 73676 12210
rect 74106 12210 74694 12226
rect 74106 12193 74122 12210
rect 73660 12176 73862 12193
rect 72902 12138 73862 12176
rect 73920 12176 74122 12193
rect 74678 12193 74694 12210
rect 74678 12176 74880 12193
rect 73920 12138 74880 12176
rect 42812 11584 43772 11622
rect 42812 11567 43014 11584
rect 42998 11550 43014 11567
rect 43570 11567 43772 11584
rect 43830 11584 44790 11622
rect 43830 11567 44032 11584
rect 43570 11550 43586 11567
rect 42998 11534 43586 11550
rect 44016 11550 44032 11567
rect 44588 11567 44790 11584
rect 44848 11584 45808 11622
rect 44848 11567 45050 11584
rect 44588 11550 44604 11567
rect 44016 11534 44604 11550
rect 42998 11476 43586 11492
rect 42998 11459 43014 11476
rect 42812 11442 43014 11459
rect 43570 11459 43586 11476
rect 45034 11550 45050 11567
rect 45606 11567 45808 11584
rect 45866 11584 46826 11622
rect 45866 11567 46068 11584
rect 45606 11550 45622 11567
rect 45034 11534 45622 11550
rect 44016 11476 44604 11492
rect 44016 11459 44032 11476
rect 43570 11442 43772 11459
rect 42812 11404 43772 11442
rect 43830 11442 44032 11459
rect 44588 11459 44604 11476
rect 46052 11550 46068 11567
rect 46624 11567 46826 11584
rect 46884 11584 47844 11622
rect 46884 11567 47086 11584
rect 46624 11550 46640 11567
rect 46052 11534 46640 11550
rect 45034 11476 45622 11492
rect 45034 11459 45050 11476
rect 44588 11442 44790 11459
rect 43830 11404 44790 11442
rect 44848 11442 45050 11459
rect 45606 11459 45622 11476
rect 47070 11550 47086 11567
rect 47642 11567 47844 11584
rect 47902 11584 48862 11622
rect 47902 11567 48104 11584
rect 47642 11550 47658 11567
rect 47070 11534 47658 11550
rect 46052 11476 46640 11492
rect 46052 11459 46068 11476
rect 45606 11442 45808 11459
rect 44848 11404 45808 11442
rect 45866 11442 46068 11459
rect 46624 11459 46640 11476
rect 48088 11550 48104 11567
rect 48660 11567 48862 11584
rect 48920 11584 49880 11622
rect 48920 11567 49122 11584
rect 48660 11550 48676 11567
rect 48088 11534 48676 11550
rect 47070 11476 47658 11492
rect 47070 11459 47086 11476
rect 46624 11442 46826 11459
rect 45866 11404 46826 11442
rect 46884 11442 47086 11459
rect 47642 11459 47658 11476
rect 49106 11550 49122 11567
rect 49678 11567 49880 11584
rect 49938 11584 50898 11622
rect 49938 11567 50140 11584
rect 49678 11550 49694 11567
rect 49106 11534 49694 11550
rect 48088 11476 48676 11492
rect 48088 11459 48104 11476
rect 47642 11442 47844 11459
rect 46884 11404 47844 11442
rect 47902 11442 48104 11459
rect 48660 11459 48676 11476
rect 50124 11550 50140 11567
rect 50696 11567 50898 11584
rect 50956 11584 51916 11622
rect 50956 11567 51158 11584
rect 50696 11550 50712 11567
rect 50124 11534 50712 11550
rect 49106 11476 49694 11492
rect 49106 11459 49122 11476
rect 48660 11442 48862 11459
rect 47902 11404 48862 11442
rect 48920 11442 49122 11459
rect 49678 11459 49694 11476
rect 51142 11550 51158 11567
rect 51714 11567 51916 11584
rect 51714 11550 51730 11567
rect 51142 11534 51730 11550
rect 50124 11476 50712 11492
rect 50124 11459 50140 11476
rect 49678 11442 49880 11459
rect 48920 11404 49880 11442
rect 49938 11442 50140 11459
rect 50696 11459 50712 11476
rect 51142 11476 51730 11492
rect 51142 11459 51158 11476
rect 50696 11442 50898 11459
rect 49938 11404 50898 11442
rect 50956 11442 51158 11459
rect 51714 11459 51730 11476
rect 54578 11500 55538 11538
rect 54578 11483 54780 11500
rect 54764 11466 54780 11483
rect 55336 11483 55538 11500
rect 55596 11500 56556 11538
rect 55596 11483 55798 11500
rect 55336 11466 55352 11483
rect 51714 11442 51916 11459
rect 54764 11450 55352 11466
rect 55782 11466 55798 11483
rect 56354 11483 56556 11500
rect 56614 11500 57574 11538
rect 56614 11483 56816 11500
rect 56354 11466 56370 11483
rect 55782 11450 56370 11466
rect 56800 11466 56816 11483
rect 57372 11483 57574 11500
rect 57632 11500 58592 11538
rect 57632 11483 57834 11500
rect 57372 11466 57388 11483
rect 56800 11450 57388 11466
rect 57818 11466 57834 11483
rect 58390 11483 58592 11500
rect 58650 11500 59610 11538
rect 58650 11483 58852 11500
rect 58390 11466 58406 11483
rect 57818 11450 58406 11466
rect 58836 11466 58852 11483
rect 59408 11483 59610 11500
rect 59668 11500 60628 11538
rect 59668 11483 59870 11500
rect 59408 11466 59424 11483
rect 58836 11450 59424 11466
rect 59854 11466 59870 11483
rect 60426 11483 60628 11500
rect 60686 11500 61646 11538
rect 60686 11483 60888 11500
rect 60426 11466 60442 11483
rect 59854 11450 60442 11466
rect 60872 11466 60888 11483
rect 61444 11483 61646 11500
rect 61704 11500 62664 11538
rect 61704 11483 61906 11500
rect 61444 11466 61460 11483
rect 60872 11450 61460 11466
rect 61890 11466 61906 11483
rect 62462 11483 62664 11500
rect 62722 11500 63682 11538
rect 62722 11483 62924 11500
rect 62462 11466 62478 11483
rect 61890 11450 62478 11466
rect 62908 11466 62924 11483
rect 63480 11483 63682 11500
rect 63740 11500 64700 11538
rect 63740 11483 63942 11500
rect 63480 11466 63496 11483
rect 62908 11450 63496 11466
rect 63926 11466 63942 11483
rect 64498 11483 64700 11500
rect 64758 11500 65718 11538
rect 64758 11483 64960 11500
rect 64498 11466 64514 11483
rect 63926 11450 64514 11466
rect 64944 11466 64960 11483
rect 65516 11483 65718 11500
rect 65776 11500 66736 11538
rect 65776 11483 65978 11500
rect 65516 11466 65532 11483
rect 64944 11450 65532 11466
rect 65962 11466 65978 11483
rect 66534 11483 66736 11500
rect 66794 11500 67754 11538
rect 66794 11483 66996 11500
rect 66534 11466 66550 11483
rect 65962 11450 66550 11466
rect 66980 11466 66996 11483
rect 67552 11483 67754 11500
rect 67812 11500 68772 11538
rect 67812 11483 68014 11500
rect 67552 11466 67568 11483
rect 66980 11450 67568 11466
rect 67998 11466 68014 11483
rect 68570 11483 68772 11500
rect 68830 11500 69790 11538
rect 68830 11483 69032 11500
rect 68570 11466 68586 11483
rect 67998 11450 68586 11466
rect 69016 11466 69032 11483
rect 69588 11483 69790 11500
rect 69848 11500 70808 11538
rect 69848 11483 70050 11500
rect 69588 11466 69604 11483
rect 69016 11450 69604 11466
rect 70034 11466 70050 11483
rect 70606 11483 70808 11500
rect 70866 11500 71826 11538
rect 70866 11483 71068 11500
rect 70606 11466 70622 11483
rect 70034 11450 70622 11466
rect 71052 11466 71068 11483
rect 71624 11483 71826 11500
rect 71884 11500 72844 11538
rect 71884 11483 72086 11500
rect 71624 11466 71640 11483
rect 71052 11450 71640 11466
rect 72070 11466 72086 11483
rect 72642 11483 72844 11500
rect 72902 11500 73862 11538
rect 72902 11483 73104 11500
rect 72642 11466 72658 11483
rect 72070 11450 72658 11466
rect 73088 11466 73104 11483
rect 73660 11483 73862 11500
rect 73920 11500 74880 11538
rect 73920 11483 74122 11500
rect 73660 11466 73676 11483
rect 73088 11450 73676 11466
rect 74106 11466 74122 11483
rect 74678 11483 74880 11500
rect 74678 11466 74694 11483
rect 74106 11450 74694 11466
rect 50956 11404 51916 11442
rect 54764 10978 55352 10994
rect 54764 10961 54780 10978
rect 54578 10944 54780 10961
rect 55336 10961 55352 10978
rect 55782 10978 56370 10994
rect 55782 10961 55798 10978
rect 55336 10944 55538 10961
rect 54578 10906 55538 10944
rect 55596 10944 55798 10961
rect 56354 10961 56370 10978
rect 56800 10978 57388 10994
rect 56800 10961 56816 10978
rect 56354 10944 56556 10961
rect 55596 10906 56556 10944
rect 56614 10944 56816 10961
rect 57372 10961 57388 10978
rect 57818 10978 58406 10994
rect 57818 10961 57834 10978
rect 57372 10944 57574 10961
rect 56614 10906 57574 10944
rect 57632 10944 57834 10961
rect 58390 10961 58406 10978
rect 58836 10978 59424 10994
rect 58836 10961 58852 10978
rect 58390 10944 58592 10961
rect 57632 10906 58592 10944
rect 58650 10944 58852 10961
rect 59408 10961 59424 10978
rect 59854 10978 60442 10994
rect 59854 10961 59870 10978
rect 59408 10944 59610 10961
rect 58650 10906 59610 10944
rect 59668 10944 59870 10961
rect 60426 10961 60442 10978
rect 60872 10978 61460 10994
rect 60872 10961 60888 10978
rect 60426 10944 60628 10961
rect 59668 10906 60628 10944
rect 60686 10944 60888 10961
rect 61444 10961 61460 10978
rect 61890 10978 62478 10994
rect 61890 10961 61906 10978
rect 61444 10944 61646 10961
rect 60686 10906 61646 10944
rect 61704 10944 61906 10961
rect 62462 10961 62478 10978
rect 62908 10978 63496 10994
rect 62908 10961 62924 10978
rect 62462 10944 62664 10961
rect 61704 10906 62664 10944
rect 62722 10944 62924 10961
rect 63480 10961 63496 10978
rect 63926 10978 64514 10994
rect 63926 10961 63942 10978
rect 63480 10944 63682 10961
rect 62722 10906 63682 10944
rect 63740 10944 63942 10961
rect 64498 10961 64514 10978
rect 64944 10978 65532 10994
rect 64944 10961 64960 10978
rect 64498 10944 64700 10961
rect 63740 10906 64700 10944
rect 64758 10944 64960 10961
rect 65516 10961 65532 10978
rect 65962 10978 66550 10994
rect 65962 10961 65978 10978
rect 65516 10944 65718 10961
rect 64758 10906 65718 10944
rect 65776 10944 65978 10961
rect 66534 10961 66550 10978
rect 66980 10978 67568 10994
rect 66980 10961 66996 10978
rect 66534 10944 66736 10961
rect 65776 10906 66736 10944
rect 66794 10944 66996 10961
rect 67552 10961 67568 10978
rect 67998 10978 68586 10994
rect 67998 10961 68014 10978
rect 67552 10944 67754 10961
rect 66794 10906 67754 10944
rect 67812 10944 68014 10961
rect 68570 10961 68586 10978
rect 69016 10978 69604 10994
rect 69016 10961 69032 10978
rect 68570 10944 68772 10961
rect 67812 10906 68772 10944
rect 68830 10944 69032 10961
rect 69588 10961 69604 10978
rect 70034 10978 70622 10994
rect 70034 10961 70050 10978
rect 69588 10944 69790 10961
rect 68830 10906 69790 10944
rect 69848 10944 70050 10961
rect 70606 10961 70622 10978
rect 71052 10978 71640 10994
rect 71052 10961 71068 10978
rect 70606 10944 70808 10961
rect 69848 10906 70808 10944
rect 70866 10944 71068 10961
rect 71624 10961 71640 10978
rect 72070 10978 72658 10994
rect 72070 10961 72086 10978
rect 71624 10944 71826 10961
rect 70866 10906 71826 10944
rect 71884 10944 72086 10961
rect 72642 10961 72658 10978
rect 73088 10978 73676 10994
rect 73088 10961 73104 10978
rect 72642 10944 72844 10961
rect 71884 10906 72844 10944
rect 72902 10944 73104 10961
rect 73660 10961 73676 10978
rect 74106 10978 74694 10994
rect 74106 10961 74122 10978
rect 73660 10944 73862 10961
rect 72902 10906 73862 10944
rect 73920 10944 74122 10961
rect 74678 10961 74694 10978
rect 74678 10944 74880 10961
rect 73920 10906 74880 10944
rect 42812 10766 43772 10804
rect 42812 10749 43014 10766
rect 42998 10732 43014 10749
rect 43570 10749 43772 10766
rect 43830 10766 44790 10804
rect 43830 10749 44032 10766
rect 43570 10732 43586 10749
rect 42998 10716 43586 10732
rect 44016 10732 44032 10749
rect 44588 10749 44790 10766
rect 44848 10766 45808 10804
rect 44848 10749 45050 10766
rect 44588 10732 44604 10749
rect 44016 10716 44604 10732
rect 42998 10658 43586 10674
rect 42998 10641 43014 10658
rect 42812 10624 43014 10641
rect 43570 10641 43586 10658
rect 45034 10732 45050 10749
rect 45606 10749 45808 10766
rect 45866 10766 46826 10804
rect 45866 10749 46068 10766
rect 45606 10732 45622 10749
rect 45034 10716 45622 10732
rect 44016 10658 44604 10674
rect 44016 10641 44032 10658
rect 43570 10624 43772 10641
rect 42812 10586 43772 10624
rect 43830 10624 44032 10641
rect 44588 10641 44604 10658
rect 46052 10732 46068 10749
rect 46624 10749 46826 10766
rect 46884 10766 47844 10804
rect 46884 10749 47086 10766
rect 46624 10732 46640 10749
rect 46052 10716 46640 10732
rect 45034 10658 45622 10674
rect 45034 10641 45050 10658
rect 44588 10624 44790 10641
rect 43830 10586 44790 10624
rect 44848 10624 45050 10641
rect 45606 10641 45622 10658
rect 47070 10732 47086 10749
rect 47642 10749 47844 10766
rect 47902 10766 48862 10804
rect 47902 10749 48104 10766
rect 47642 10732 47658 10749
rect 47070 10716 47658 10732
rect 46052 10658 46640 10674
rect 46052 10641 46068 10658
rect 45606 10624 45808 10641
rect 44848 10586 45808 10624
rect 45866 10624 46068 10641
rect 46624 10641 46640 10658
rect 48088 10732 48104 10749
rect 48660 10749 48862 10766
rect 48920 10766 49880 10804
rect 48920 10749 49122 10766
rect 48660 10732 48676 10749
rect 48088 10716 48676 10732
rect 47070 10658 47658 10674
rect 47070 10641 47086 10658
rect 46624 10624 46826 10641
rect 45866 10586 46826 10624
rect 46884 10624 47086 10641
rect 47642 10641 47658 10658
rect 49106 10732 49122 10749
rect 49678 10749 49880 10766
rect 49938 10766 50898 10804
rect 49938 10749 50140 10766
rect 49678 10732 49694 10749
rect 49106 10716 49694 10732
rect 48088 10658 48676 10674
rect 48088 10641 48104 10658
rect 47642 10624 47844 10641
rect 46884 10586 47844 10624
rect 47902 10624 48104 10641
rect 48660 10641 48676 10658
rect 50124 10732 50140 10749
rect 50696 10749 50898 10766
rect 50956 10766 51916 10804
rect 50956 10749 51158 10766
rect 50696 10732 50712 10749
rect 50124 10716 50712 10732
rect 49106 10658 49694 10674
rect 49106 10641 49122 10658
rect 48660 10624 48862 10641
rect 47902 10586 48862 10624
rect 48920 10624 49122 10641
rect 49678 10641 49694 10658
rect 51142 10732 51158 10749
rect 51714 10749 51916 10766
rect 51714 10732 51730 10749
rect 51142 10716 51730 10732
rect 50124 10658 50712 10674
rect 50124 10641 50140 10658
rect 49678 10624 49880 10641
rect 48920 10586 49880 10624
rect 49938 10624 50140 10641
rect 50696 10641 50712 10658
rect 51142 10658 51730 10674
rect 51142 10641 51158 10658
rect 50696 10624 50898 10641
rect 49938 10586 50898 10624
rect 50956 10624 51158 10641
rect 51714 10641 51730 10658
rect 51714 10624 51916 10641
rect 50956 10586 51916 10624
rect 54578 10268 55538 10306
rect 54578 10251 54780 10268
rect 54764 10234 54780 10251
rect 55336 10251 55538 10268
rect 55596 10268 56556 10306
rect 55596 10251 55798 10268
rect 55336 10234 55352 10251
rect 54764 10218 55352 10234
rect 55782 10234 55798 10251
rect 56354 10251 56556 10268
rect 56614 10268 57574 10306
rect 56614 10251 56816 10268
rect 56354 10234 56370 10251
rect 55782 10218 56370 10234
rect 56800 10234 56816 10251
rect 57372 10251 57574 10268
rect 57632 10268 58592 10306
rect 57632 10251 57834 10268
rect 57372 10234 57388 10251
rect 56800 10218 57388 10234
rect 57818 10234 57834 10251
rect 58390 10251 58592 10268
rect 58650 10268 59610 10306
rect 58650 10251 58852 10268
rect 58390 10234 58406 10251
rect 57818 10218 58406 10234
rect 58836 10234 58852 10251
rect 59408 10251 59610 10268
rect 59668 10268 60628 10306
rect 59668 10251 59870 10268
rect 59408 10234 59424 10251
rect 58836 10218 59424 10234
rect 59854 10234 59870 10251
rect 60426 10251 60628 10268
rect 60686 10268 61646 10306
rect 60686 10251 60888 10268
rect 60426 10234 60442 10251
rect 59854 10218 60442 10234
rect 60872 10234 60888 10251
rect 61444 10251 61646 10268
rect 61704 10268 62664 10306
rect 61704 10251 61906 10268
rect 61444 10234 61460 10251
rect 60872 10218 61460 10234
rect 61890 10234 61906 10251
rect 62462 10251 62664 10268
rect 62722 10268 63682 10306
rect 62722 10251 62924 10268
rect 62462 10234 62478 10251
rect 61890 10218 62478 10234
rect 62908 10234 62924 10251
rect 63480 10251 63682 10268
rect 63740 10268 64700 10306
rect 63740 10251 63942 10268
rect 63480 10234 63496 10251
rect 62908 10218 63496 10234
rect 63926 10234 63942 10251
rect 64498 10251 64700 10268
rect 64758 10268 65718 10306
rect 64758 10251 64960 10268
rect 64498 10234 64514 10251
rect 63926 10218 64514 10234
rect 64944 10234 64960 10251
rect 65516 10251 65718 10268
rect 65776 10268 66736 10306
rect 65776 10251 65978 10268
rect 65516 10234 65532 10251
rect 64944 10218 65532 10234
rect 65962 10234 65978 10251
rect 66534 10251 66736 10268
rect 66794 10268 67754 10306
rect 66794 10251 66996 10268
rect 66534 10234 66550 10251
rect 65962 10218 66550 10234
rect 66980 10234 66996 10251
rect 67552 10251 67754 10268
rect 67812 10268 68772 10306
rect 67812 10251 68014 10268
rect 67552 10234 67568 10251
rect 66980 10218 67568 10234
rect 67998 10234 68014 10251
rect 68570 10251 68772 10268
rect 68830 10268 69790 10306
rect 68830 10251 69032 10268
rect 68570 10234 68586 10251
rect 67998 10218 68586 10234
rect 69016 10234 69032 10251
rect 69588 10251 69790 10268
rect 69848 10268 70808 10306
rect 69848 10251 70050 10268
rect 69588 10234 69604 10251
rect 69016 10218 69604 10234
rect 70034 10234 70050 10251
rect 70606 10251 70808 10268
rect 70866 10268 71826 10306
rect 70866 10251 71068 10268
rect 70606 10234 70622 10251
rect 70034 10218 70622 10234
rect 71052 10234 71068 10251
rect 71624 10251 71826 10268
rect 71884 10268 72844 10306
rect 71884 10251 72086 10268
rect 71624 10234 71640 10251
rect 71052 10218 71640 10234
rect 72070 10234 72086 10251
rect 72642 10251 72844 10268
rect 72902 10268 73862 10306
rect 72902 10251 73104 10268
rect 72642 10234 72658 10251
rect 72070 10218 72658 10234
rect 73088 10234 73104 10251
rect 73660 10251 73862 10268
rect 73920 10268 74880 10306
rect 73920 10251 74122 10268
rect 73660 10234 73676 10251
rect 73088 10218 73676 10234
rect 74106 10234 74122 10251
rect 74678 10251 74880 10268
rect 74678 10234 74694 10251
rect 74106 10218 74694 10234
rect 42812 9948 43772 9986
rect 42812 9931 43014 9948
rect 42998 9914 43014 9931
rect 43570 9931 43772 9948
rect 43830 9948 44790 9986
rect 43830 9931 44032 9948
rect 43570 9914 43586 9931
rect 42998 9898 43586 9914
rect 44016 9914 44032 9931
rect 44588 9931 44790 9948
rect 44848 9948 45808 9986
rect 44848 9931 45050 9948
rect 44588 9914 44604 9931
rect 44016 9898 44604 9914
rect 42998 9840 43586 9856
rect 42998 9823 43014 9840
rect 42812 9806 43014 9823
rect 43570 9823 43586 9840
rect 45034 9914 45050 9931
rect 45606 9931 45808 9948
rect 45866 9948 46826 9986
rect 45866 9931 46068 9948
rect 45606 9914 45622 9931
rect 45034 9898 45622 9914
rect 44016 9840 44604 9856
rect 44016 9823 44032 9840
rect 43570 9806 43772 9823
rect 42812 9768 43772 9806
rect 43830 9806 44032 9823
rect 44588 9823 44604 9840
rect 46052 9914 46068 9931
rect 46624 9931 46826 9948
rect 46884 9948 47844 9986
rect 46884 9931 47086 9948
rect 46624 9914 46640 9931
rect 46052 9898 46640 9914
rect 45034 9840 45622 9856
rect 45034 9823 45050 9840
rect 44588 9806 44790 9823
rect 43830 9768 44790 9806
rect 44848 9806 45050 9823
rect 45606 9823 45622 9840
rect 47070 9914 47086 9931
rect 47642 9931 47844 9948
rect 47902 9948 48862 9986
rect 47902 9931 48104 9948
rect 47642 9914 47658 9931
rect 47070 9898 47658 9914
rect 46052 9840 46640 9856
rect 46052 9823 46068 9840
rect 45606 9806 45808 9823
rect 44848 9768 45808 9806
rect 45866 9806 46068 9823
rect 46624 9823 46640 9840
rect 48088 9914 48104 9931
rect 48660 9931 48862 9948
rect 48920 9948 49880 9986
rect 48920 9931 49122 9948
rect 48660 9914 48676 9931
rect 48088 9898 48676 9914
rect 47070 9840 47658 9856
rect 47070 9823 47086 9840
rect 46624 9806 46826 9823
rect 45866 9768 46826 9806
rect 46884 9806 47086 9823
rect 47642 9823 47658 9840
rect 49106 9914 49122 9931
rect 49678 9931 49880 9948
rect 49938 9948 50898 9986
rect 49938 9931 50140 9948
rect 49678 9914 49694 9931
rect 49106 9898 49694 9914
rect 48088 9840 48676 9856
rect 48088 9823 48104 9840
rect 47642 9806 47844 9823
rect 46884 9768 47844 9806
rect 47902 9806 48104 9823
rect 48660 9823 48676 9840
rect 50124 9914 50140 9931
rect 50696 9931 50898 9948
rect 50956 9948 51916 9986
rect 50956 9931 51158 9948
rect 50696 9914 50712 9931
rect 50124 9898 50712 9914
rect 49106 9840 49694 9856
rect 49106 9823 49122 9840
rect 48660 9806 48862 9823
rect 47902 9768 48862 9806
rect 48920 9806 49122 9823
rect 49678 9823 49694 9840
rect 51142 9914 51158 9931
rect 51714 9931 51916 9948
rect 51714 9914 51730 9931
rect 51142 9898 51730 9914
rect 50124 9840 50712 9856
rect 50124 9823 50140 9840
rect 49678 9806 49880 9823
rect 48920 9768 49880 9806
rect 49938 9806 50140 9823
rect 50696 9823 50712 9840
rect 51142 9840 51730 9856
rect 51142 9823 51158 9840
rect 50696 9806 50898 9823
rect 49938 9768 50898 9806
rect 50956 9806 51158 9823
rect 51714 9823 51730 9840
rect 51714 9806 51916 9823
rect 50956 9768 51916 9806
rect 54762 9744 55350 9760
rect 54762 9727 54778 9744
rect 54576 9710 54778 9727
rect 55334 9727 55350 9744
rect 55780 9744 56368 9760
rect 55780 9727 55796 9744
rect 55334 9710 55536 9727
rect 54576 9672 55536 9710
rect 55594 9710 55796 9727
rect 56352 9727 56368 9744
rect 56798 9744 57386 9760
rect 56798 9727 56814 9744
rect 56352 9710 56554 9727
rect 55594 9672 56554 9710
rect 56612 9710 56814 9727
rect 57370 9727 57386 9744
rect 57816 9744 58404 9760
rect 57816 9727 57832 9744
rect 57370 9710 57572 9727
rect 56612 9672 57572 9710
rect 57630 9710 57832 9727
rect 58388 9727 58404 9744
rect 58834 9744 59422 9760
rect 58834 9727 58850 9744
rect 58388 9710 58590 9727
rect 57630 9672 58590 9710
rect 58648 9710 58850 9727
rect 59406 9727 59422 9744
rect 59852 9744 60440 9760
rect 59852 9727 59868 9744
rect 59406 9710 59608 9727
rect 58648 9672 59608 9710
rect 59666 9710 59868 9727
rect 60424 9727 60440 9744
rect 60870 9744 61458 9760
rect 60870 9727 60886 9744
rect 60424 9710 60626 9727
rect 59666 9672 60626 9710
rect 60684 9710 60886 9727
rect 61442 9727 61458 9744
rect 61888 9744 62476 9760
rect 61888 9727 61904 9744
rect 61442 9710 61644 9727
rect 60684 9672 61644 9710
rect 61702 9710 61904 9727
rect 62460 9727 62476 9744
rect 62906 9744 63494 9760
rect 62906 9727 62922 9744
rect 62460 9710 62662 9727
rect 61702 9672 62662 9710
rect 62720 9710 62922 9727
rect 63478 9727 63494 9744
rect 63924 9744 64512 9760
rect 63924 9727 63940 9744
rect 63478 9710 63680 9727
rect 62720 9672 63680 9710
rect 63738 9710 63940 9727
rect 64496 9727 64512 9744
rect 64942 9744 65530 9760
rect 64942 9727 64958 9744
rect 64496 9710 64698 9727
rect 63738 9672 64698 9710
rect 64756 9710 64958 9727
rect 65514 9727 65530 9744
rect 65960 9744 66548 9760
rect 65960 9727 65976 9744
rect 65514 9710 65716 9727
rect 64756 9672 65716 9710
rect 65774 9710 65976 9727
rect 66532 9727 66548 9744
rect 66978 9744 67566 9760
rect 66978 9727 66994 9744
rect 66532 9710 66734 9727
rect 65774 9672 66734 9710
rect 66792 9710 66994 9727
rect 67550 9727 67566 9744
rect 67996 9744 68584 9760
rect 67996 9727 68012 9744
rect 67550 9710 67752 9727
rect 66792 9672 67752 9710
rect 67810 9710 68012 9727
rect 68568 9727 68584 9744
rect 69014 9744 69602 9760
rect 69014 9727 69030 9744
rect 68568 9710 68770 9727
rect 67810 9672 68770 9710
rect 68828 9710 69030 9727
rect 69586 9727 69602 9744
rect 70032 9744 70620 9760
rect 70032 9727 70048 9744
rect 69586 9710 69788 9727
rect 68828 9672 69788 9710
rect 69846 9710 70048 9727
rect 70604 9727 70620 9744
rect 71050 9744 71638 9760
rect 71050 9727 71066 9744
rect 70604 9710 70806 9727
rect 69846 9672 70806 9710
rect 70864 9710 71066 9727
rect 71622 9727 71638 9744
rect 72068 9744 72656 9760
rect 72068 9727 72084 9744
rect 71622 9710 71824 9727
rect 70864 9672 71824 9710
rect 71882 9710 72084 9727
rect 72640 9727 72656 9744
rect 73086 9744 73674 9760
rect 73086 9727 73102 9744
rect 72640 9710 72842 9727
rect 71882 9672 72842 9710
rect 72900 9710 73102 9727
rect 73658 9727 73674 9744
rect 74104 9744 74692 9760
rect 74104 9727 74120 9744
rect 73658 9710 73860 9727
rect 72900 9672 73860 9710
rect 73918 9710 74120 9727
rect 74676 9727 74692 9744
rect 74676 9710 74878 9727
rect 73918 9672 74878 9710
rect 42812 9130 43772 9168
rect 42812 9113 43014 9130
rect 42998 9096 43014 9113
rect 43570 9113 43772 9130
rect 43830 9130 44790 9168
rect 43830 9113 44032 9130
rect 43570 9096 43586 9113
rect 42998 9080 43586 9096
rect 44016 9096 44032 9113
rect 44588 9113 44790 9130
rect 44848 9130 45808 9168
rect 44848 9113 45050 9130
rect 44588 9096 44604 9113
rect 44016 9080 44604 9096
rect 42998 9022 43586 9038
rect 42998 9005 43014 9022
rect 42812 8988 43014 9005
rect 43570 9005 43586 9022
rect 45034 9096 45050 9113
rect 45606 9113 45808 9130
rect 45866 9130 46826 9168
rect 45866 9113 46068 9130
rect 45606 9096 45622 9113
rect 45034 9080 45622 9096
rect 44016 9022 44604 9038
rect 44016 9005 44032 9022
rect 43570 8988 43772 9005
rect 42812 8950 43772 8988
rect 43830 8988 44032 9005
rect 44588 9005 44604 9022
rect 46052 9096 46068 9113
rect 46624 9113 46826 9130
rect 46884 9130 47844 9168
rect 46884 9113 47086 9130
rect 46624 9096 46640 9113
rect 46052 9080 46640 9096
rect 45034 9022 45622 9038
rect 45034 9005 45050 9022
rect 44588 8988 44790 9005
rect 43830 8950 44790 8988
rect 44848 8988 45050 9005
rect 45606 9005 45622 9022
rect 47070 9096 47086 9113
rect 47642 9113 47844 9130
rect 47902 9130 48862 9168
rect 47902 9113 48104 9130
rect 47642 9096 47658 9113
rect 47070 9080 47658 9096
rect 46052 9022 46640 9038
rect 46052 9005 46068 9022
rect 45606 8988 45808 9005
rect 44848 8950 45808 8988
rect 45866 8988 46068 9005
rect 46624 9005 46640 9022
rect 48088 9096 48104 9113
rect 48660 9113 48862 9130
rect 48920 9130 49880 9168
rect 48920 9113 49122 9130
rect 48660 9096 48676 9113
rect 48088 9080 48676 9096
rect 47070 9022 47658 9038
rect 47070 9005 47086 9022
rect 46624 8988 46826 9005
rect 45866 8950 46826 8988
rect 46884 8988 47086 9005
rect 47642 9005 47658 9022
rect 49106 9096 49122 9113
rect 49678 9113 49880 9130
rect 49938 9130 50898 9168
rect 49938 9113 50140 9130
rect 49678 9096 49694 9113
rect 49106 9080 49694 9096
rect 48088 9022 48676 9038
rect 48088 9005 48104 9022
rect 47642 8988 47844 9005
rect 46884 8950 47844 8988
rect 47902 8988 48104 9005
rect 48660 9005 48676 9022
rect 50124 9096 50140 9113
rect 50696 9113 50898 9130
rect 50956 9130 51916 9168
rect 50956 9113 51158 9130
rect 50696 9096 50712 9113
rect 50124 9080 50712 9096
rect 49106 9022 49694 9038
rect 49106 9005 49122 9022
rect 48660 8988 48862 9005
rect 47902 8950 48862 8988
rect 48920 8988 49122 9005
rect 49678 9005 49694 9022
rect 51142 9096 51158 9113
rect 51714 9113 51916 9130
rect 51714 9096 51730 9113
rect 51142 9080 51730 9096
rect 50124 9022 50712 9038
rect 50124 9005 50140 9022
rect 49678 8988 49880 9005
rect 48920 8950 49880 8988
rect 49938 8988 50140 9005
rect 50696 9005 50712 9022
rect 51142 9022 51730 9038
rect 51142 9005 51158 9022
rect 50696 8988 50898 9005
rect 49938 8950 50898 8988
rect 50956 8988 51158 9005
rect 51714 9005 51730 9022
rect 54576 9034 55536 9072
rect 54576 9017 54778 9034
rect 51714 8988 51916 9005
rect 50956 8950 51916 8988
rect 54762 9000 54778 9017
rect 55334 9017 55536 9034
rect 55594 9034 56554 9072
rect 55594 9017 55796 9034
rect 55334 9000 55350 9017
rect 54762 8984 55350 9000
rect 55780 9000 55796 9017
rect 56352 9017 56554 9034
rect 56612 9034 57572 9072
rect 56612 9017 56814 9034
rect 56352 9000 56368 9017
rect 55780 8984 56368 9000
rect 56798 9000 56814 9017
rect 57370 9017 57572 9034
rect 57630 9034 58590 9072
rect 57630 9017 57832 9034
rect 57370 9000 57386 9017
rect 56798 8984 57386 9000
rect 57816 9000 57832 9017
rect 58388 9017 58590 9034
rect 58648 9034 59608 9072
rect 58648 9017 58850 9034
rect 58388 9000 58404 9017
rect 57816 8984 58404 9000
rect 58834 9000 58850 9017
rect 59406 9017 59608 9034
rect 59666 9034 60626 9072
rect 59666 9017 59868 9034
rect 59406 9000 59422 9017
rect 58834 8984 59422 9000
rect 59852 9000 59868 9017
rect 60424 9017 60626 9034
rect 60684 9034 61644 9072
rect 60684 9017 60886 9034
rect 60424 9000 60440 9017
rect 59852 8984 60440 9000
rect 60870 9000 60886 9017
rect 61442 9017 61644 9034
rect 61702 9034 62662 9072
rect 61702 9017 61904 9034
rect 61442 9000 61458 9017
rect 60870 8984 61458 9000
rect 61888 9000 61904 9017
rect 62460 9017 62662 9034
rect 62720 9034 63680 9072
rect 62720 9017 62922 9034
rect 62460 9000 62476 9017
rect 61888 8984 62476 9000
rect 62906 9000 62922 9017
rect 63478 9017 63680 9034
rect 63738 9034 64698 9072
rect 63738 9017 63940 9034
rect 63478 9000 63494 9017
rect 62906 8984 63494 9000
rect 63924 9000 63940 9017
rect 64496 9017 64698 9034
rect 64756 9034 65716 9072
rect 64756 9017 64958 9034
rect 64496 9000 64512 9017
rect 63924 8984 64512 9000
rect 64942 9000 64958 9017
rect 65514 9017 65716 9034
rect 65774 9034 66734 9072
rect 65774 9017 65976 9034
rect 65514 9000 65530 9017
rect 64942 8984 65530 9000
rect 65960 9000 65976 9017
rect 66532 9017 66734 9034
rect 66792 9034 67752 9072
rect 66792 9017 66994 9034
rect 66532 9000 66548 9017
rect 65960 8984 66548 9000
rect 66978 9000 66994 9017
rect 67550 9017 67752 9034
rect 67810 9034 68770 9072
rect 67810 9017 68012 9034
rect 67550 9000 67566 9017
rect 66978 8984 67566 9000
rect 67996 9000 68012 9017
rect 68568 9017 68770 9034
rect 68828 9034 69788 9072
rect 68828 9017 69030 9034
rect 68568 9000 68584 9017
rect 67996 8984 68584 9000
rect 69014 9000 69030 9017
rect 69586 9017 69788 9034
rect 69846 9034 70806 9072
rect 69846 9017 70048 9034
rect 69586 9000 69602 9017
rect 69014 8984 69602 9000
rect 70032 9000 70048 9017
rect 70604 9017 70806 9034
rect 70864 9034 71824 9072
rect 70864 9017 71066 9034
rect 70604 9000 70620 9017
rect 70032 8984 70620 9000
rect 71050 9000 71066 9017
rect 71622 9017 71824 9034
rect 71882 9034 72842 9072
rect 71882 9017 72084 9034
rect 71622 9000 71638 9017
rect 71050 8984 71638 9000
rect 72068 9000 72084 9017
rect 72640 9017 72842 9034
rect 72900 9034 73860 9072
rect 72900 9017 73102 9034
rect 72640 9000 72656 9017
rect 72068 8984 72656 9000
rect 73086 9000 73102 9017
rect 73658 9017 73860 9034
rect 73918 9034 74878 9072
rect 73918 9017 74120 9034
rect 73658 9000 73674 9017
rect 73086 8984 73674 9000
rect 74104 9000 74120 9017
rect 74676 9017 74878 9034
rect 74676 9000 74692 9017
rect 74104 8984 74692 9000
rect 54762 8510 55350 8526
rect 54762 8493 54778 8510
rect 54576 8476 54778 8493
rect 55334 8493 55350 8510
rect 55780 8510 56368 8526
rect 55780 8493 55796 8510
rect 55334 8476 55536 8493
rect 54576 8438 55536 8476
rect 55594 8476 55796 8493
rect 56352 8493 56368 8510
rect 56798 8510 57386 8526
rect 56798 8493 56814 8510
rect 56352 8476 56554 8493
rect 55594 8438 56554 8476
rect 56612 8476 56814 8493
rect 57370 8493 57386 8510
rect 57816 8510 58404 8526
rect 57816 8493 57832 8510
rect 57370 8476 57572 8493
rect 56612 8438 57572 8476
rect 57630 8476 57832 8493
rect 58388 8493 58404 8510
rect 58834 8510 59422 8526
rect 58834 8493 58850 8510
rect 58388 8476 58590 8493
rect 57630 8438 58590 8476
rect 58648 8476 58850 8493
rect 59406 8493 59422 8510
rect 59852 8510 60440 8526
rect 59852 8493 59868 8510
rect 59406 8476 59608 8493
rect 58648 8438 59608 8476
rect 59666 8476 59868 8493
rect 60424 8493 60440 8510
rect 60870 8510 61458 8526
rect 60870 8493 60886 8510
rect 60424 8476 60626 8493
rect 59666 8438 60626 8476
rect 60684 8476 60886 8493
rect 61442 8493 61458 8510
rect 61888 8510 62476 8526
rect 61888 8493 61904 8510
rect 61442 8476 61644 8493
rect 60684 8438 61644 8476
rect 61702 8476 61904 8493
rect 62460 8493 62476 8510
rect 62906 8510 63494 8526
rect 62906 8493 62922 8510
rect 62460 8476 62662 8493
rect 61702 8438 62662 8476
rect 62720 8476 62922 8493
rect 63478 8493 63494 8510
rect 63924 8510 64512 8526
rect 63924 8493 63940 8510
rect 63478 8476 63680 8493
rect 62720 8438 63680 8476
rect 63738 8476 63940 8493
rect 64496 8493 64512 8510
rect 64942 8510 65530 8526
rect 64942 8493 64958 8510
rect 64496 8476 64698 8493
rect 63738 8438 64698 8476
rect 64756 8476 64958 8493
rect 65514 8493 65530 8510
rect 65960 8510 66548 8526
rect 65960 8493 65976 8510
rect 65514 8476 65716 8493
rect 64756 8438 65716 8476
rect 65774 8476 65976 8493
rect 66532 8493 66548 8510
rect 66978 8510 67566 8526
rect 66978 8493 66994 8510
rect 66532 8476 66734 8493
rect 65774 8438 66734 8476
rect 66792 8476 66994 8493
rect 67550 8493 67566 8510
rect 67996 8510 68584 8526
rect 67996 8493 68012 8510
rect 67550 8476 67752 8493
rect 66792 8438 67752 8476
rect 67810 8476 68012 8493
rect 68568 8493 68584 8510
rect 69014 8510 69602 8526
rect 69014 8493 69030 8510
rect 68568 8476 68770 8493
rect 67810 8438 68770 8476
rect 68828 8476 69030 8493
rect 69586 8493 69602 8510
rect 70032 8510 70620 8526
rect 70032 8493 70048 8510
rect 69586 8476 69788 8493
rect 68828 8438 69788 8476
rect 69846 8476 70048 8493
rect 70604 8493 70620 8510
rect 71050 8510 71638 8526
rect 71050 8493 71066 8510
rect 70604 8476 70806 8493
rect 69846 8438 70806 8476
rect 70864 8476 71066 8493
rect 71622 8493 71638 8510
rect 72068 8510 72656 8526
rect 72068 8493 72084 8510
rect 71622 8476 71824 8493
rect 70864 8438 71824 8476
rect 71882 8476 72084 8493
rect 72640 8493 72656 8510
rect 73086 8510 73674 8526
rect 73086 8493 73102 8510
rect 72640 8476 72842 8493
rect 71882 8438 72842 8476
rect 72900 8476 73102 8493
rect 73658 8493 73674 8510
rect 74104 8510 74692 8526
rect 74104 8493 74120 8510
rect 73658 8476 73860 8493
rect 72900 8438 73860 8476
rect 73918 8476 74120 8493
rect 74676 8493 74692 8510
rect 74676 8476 74878 8493
rect 73918 8438 74878 8476
rect 42812 8312 43772 8350
rect 42812 8295 43014 8312
rect 42998 8278 43014 8295
rect 43570 8295 43772 8312
rect 43830 8312 44790 8350
rect 43830 8295 44032 8312
rect 43570 8278 43586 8295
rect 42998 8262 43586 8278
rect 44016 8278 44032 8295
rect 44588 8295 44790 8312
rect 44848 8312 45808 8350
rect 44848 8295 45050 8312
rect 44588 8278 44604 8295
rect 44016 8262 44604 8278
rect 42998 8204 43586 8220
rect 42998 8187 43014 8204
rect 42812 8170 43014 8187
rect 43570 8187 43586 8204
rect 45034 8278 45050 8295
rect 45606 8295 45808 8312
rect 45866 8312 46826 8350
rect 45866 8295 46068 8312
rect 45606 8278 45622 8295
rect 45034 8262 45622 8278
rect 44016 8204 44604 8220
rect 44016 8187 44032 8204
rect 43570 8170 43772 8187
rect 42812 8132 43772 8170
rect 43830 8170 44032 8187
rect 44588 8187 44604 8204
rect 46052 8278 46068 8295
rect 46624 8295 46826 8312
rect 46884 8312 47844 8350
rect 46884 8295 47086 8312
rect 46624 8278 46640 8295
rect 46052 8262 46640 8278
rect 45034 8204 45622 8220
rect 45034 8187 45050 8204
rect 44588 8170 44790 8187
rect 43830 8132 44790 8170
rect 44848 8170 45050 8187
rect 45606 8187 45622 8204
rect 47070 8278 47086 8295
rect 47642 8295 47844 8312
rect 47902 8312 48862 8350
rect 47902 8295 48104 8312
rect 47642 8278 47658 8295
rect 47070 8262 47658 8278
rect 46052 8204 46640 8220
rect 46052 8187 46068 8204
rect 45606 8170 45808 8187
rect 44848 8132 45808 8170
rect 45866 8170 46068 8187
rect 46624 8187 46640 8204
rect 48088 8278 48104 8295
rect 48660 8295 48862 8312
rect 48920 8312 49880 8350
rect 48920 8295 49122 8312
rect 48660 8278 48676 8295
rect 48088 8262 48676 8278
rect 47070 8204 47658 8220
rect 47070 8187 47086 8204
rect 46624 8170 46826 8187
rect 45866 8132 46826 8170
rect 46884 8170 47086 8187
rect 47642 8187 47658 8204
rect 49106 8278 49122 8295
rect 49678 8295 49880 8312
rect 49938 8312 50898 8350
rect 49938 8295 50140 8312
rect 49678 8278 49694 8295
rect 49106 8262 49694 8278
rect 48088 8204 48676 8220
rect 48088 8187 48104 8204
rect 47642 8170 47844 8187
rect 46884 8132 47844 8170
rect 47902 8170 48104 8187
rect 48660 8187 48676 8204
rect 50124 8278 50140 8295
rect 50696 8295 50898 8312
rect 50956 8312 51916 8350
rect 50956 8295 51158 8312
rect 50696 8278 50712 8295
rect 50124 8262 50712 8278
rect 49106 8204 49694 8220
rect 49106 8187 49122 8204
rect 48660 8170 48862 8187
rect 47902 8132 48862 8170
rect 48920 8170 49122 8187
rect 49678 8187 49694 8204
rect 51142 8278 51158 8295
rect 51714 8295 51916 8312
rect 51714 8278 51730 8295
rect 51142 8262 51730 8278
rect 50124 8204 50712 8220
rect 50124 8187 50140 8204
rect 49678 8170 49880 8187
rect 48920 8132 49880 8170
rect 49938 8170 50140 8187
rect 50696 8187 50712 8204
rect 51142 8204 51730 8220
rect 51142 8187 51158 8204
rect 50696 8170 50898 8187
rect 49938 8132 50898 8170
rect 50956 8170 51158 8187
rect 51714 8187 51730 8204
rect 51714 8170 51916 8187
rect 50956 8132 51916 8170
rect 54576 7800 55536 7838
rect 54576 7783 54778 7800
rect 54762 7766 54778 7783
rect 55334 7783 55536 7800
rect 55594 7800 56554 7838
rect 55594 7783 55796 7800
rect 55334 7766 55350 7783
rect 54762 7750 55350 7766
rect 55780 7766 55796 7783
rect 56352 7783 56554 7800
rect 56612 7800 57572 7838
rect 56612 7783 56814 7800
rect 56352 7766 56368 7783
rect 55780 7750 56368 7766
rect 56798 7766 56814 7783
rect 57370 7783 57572 7800
rect 57630 7800 58590 7838
rect 57630 7783 57832 7800
rect 57370 7766 57386 7783
rect 56798 7750 57386 7766
rect 57816 7766 57832 7783
rect 58388 7783 58590 7800
rect 58648 7800 59608 7838
rect 58648 7783 58850 7800
rect 58388 7766 58404 7783
rect 57816 7750 58404 7766
rect 58834 7766 58850 7783
rect 59406 7783 59608 7800
rect 59666 7800 60626 7838
rect 59666 7783 59868 7800
rect 59406 7766 59422 7783
rect 58834 7750 59422 7766
rect 59852 7766 59868 7783
rect 60424 7783 60626 7800
rect 60684 7800 61644 7838
rect 60684 7783 60886 7800
rect 60424 7766 60440 7783
rect 59852 7750 60440 7766
rect 60870 7766 60886 7783
rect 61442 7783 61644 7800
rect 61702 7800 62662 7838
rect 61702 7783 61904 7800
rect 61442 7766 61458 7783
rect 60870 7750 61458 7766
rect 61888 7766 61904 7783
rect 62460 7783 62662 7800
rect 62720 7800 63680 7838
rect 62720 7783 62922 7800
rect 62460 7766 62476 7783
rect 61888 7750 62476 7766
rect 62906 7766 62922 7783
rect 63478 7783 63680 7800
rect 63738 7800 64698 7838
rect 63738 7783 63940 7800
rect 63478 7766 63494 7783
rect 62906 7750 63494 7766
rect 63924 7766 63940 7783
rect 64496 7783 64698 7800
rect 64756 7800 65716 7838
rect 64756 7783 64958 7800
rect 64496 7766 64512 7783
rect 63924 7750 64512 7766
rect 64942 7766 64958 7783
rect 65514 7783 65716 7800
rect 65774 7800 66734 7838
rect 65774 7783 65976 7800
rect 65514 7766 65530 7783
rect 64942 7750 65530 7766
rect 65960 7766 65976 7783
rect 66532 7783 66734 7800
rect 66792 7800 67752 7838
rect 66792 7783 66994 7800
rect 66532 7766 66548 7783
rect 65960 7750 66548 7766
rect 66978 7766 66994 7783
rect 67550 7783 67752 7800
rect 67810 7800 68770 7838
rect 67810 7783 68012 7800
rect 67550 7766 67566 7783
rect 66978 7750 67566 7766
rect 67996 7766 68012 7783
rect 68568 7783 68770 7800
rect 68828 7800 69788 7838
rect 68828 7783 69030 7800
rect 68568 7766 68584 7783
rect 67996 7750 68584 7766
rect 69014 7766 69030 7783
rect 69586 7783 69788 7800
rect 69846 7800 70806 7838
rect 69846 7783 70048 7800
rect 69586 7766 69602 7783
rect 69014 7750 69602 7766
rect 70032 7766 70048 7783
rect 70604 7783 70806 7800
rect 70864 7800 71824 7838
rect 70864 7783 71066 7800
rect 70604 7766 70620 7783
rect 70032 7750 70620 7766
rect 71050 7766 71066 7783
rect 71622 7783 71824 7800
rect 71882 7800 72842 7838
rect 71882 7783 72084 7800
rect 71622 7766 71638 7783
rect 71050 7750 71638 7766
rect 72068 7766 72084 7783
rect 72640 7783 72842 7800
rect 72900 7800 73860 7838
rect 72900 7783 73102 7800
rect 72640 7766 72656 7783
rect 72068 7750 72656 7766
rect 73086 7766 73102 7783
rect 73658 7783 73860 7800
rect 73918 7800 74878 7838
rect 73918 7783 74120 7800
rect 73658 7766 73674 7783
rect 73086 7750 73674 7766
rect 74104 7766 74120 7783
rect 74676 7783 74878 7800
rect 74676 7766 74692 7783
rect 74104 7750 74692 7766
rect 42812 7494 43772 7532
rect 42812 7477 43014 7494
rect 42998 7460 43014 7477
rect 43570 7477 43772 7494
rect 43830 7494 44790 7532
rect 43830 7477 44032 7494
rect 43570 7460 43586 7477
rect 42998 7444 43586 7460
rect 44016 7460 44032 7477
rect 44588 7477 44790 7494
rect 44848 7494 45808 7532
rect 44848 7477 45050 7494
rect 44588 7460 44604 7477
rect 44016 7444 44604 7460
rect 45034 7460 45050 7477
rect 45606 7477 45808 7494
rect 45866 7494 46826 7532
rect 45866 7477 46068 7494
rect 45606 7460 45622 7477
rect 45034 7444 45622 7460
rect 46052 7460 46068 7477
rect 46624 7477 46826 7494
rect 46884 7494 47844 7532
rect 46884 7477 47086 7494
rect 46624 7460 46640 7477
rect 46052 7444 46640 7460
rect 47070 7460 47086 7477
rect 47642 7477 47844 7494
rect 47902 7494 48862 7532
rect 47902 7477 48104 7494
rect 47642 7460 47658 7477
rect 47070 7444 47658 7460
rect 48088 7460 48104 7477
rect 48660 7477 48862 7494
rect 48920 7494 49880 7532
rect 48920 7477 49122 7494
rect 48660 7460 48676 7477
rect 48088 7444 48676 7460
rect 49106 7460 49122 7477
rect 49678 7477 49880 7494
rect 49938 7494 50898 7532
rect 49938 7477 50140 7494
rect 49678 7460 49694 7477
rect 49106 7444 49694 7460
rect 50124 7460 50140 7477
rect 50696 7477 50898 7494
rect 50956 7494 51916 7532
rect 50956 7477 51158 7494
rect 50696 7460 50712 7477
rect 50124 7444 50712 7460
rect 51142 7460 51158 7477
rect 51714 7477 51916 7494
rect 51714 7460 51730 7477
rect 51142 7444 51730 7460
rect 54762 7278 55350 7294
rect 54762 7261 54778 7278
rect 54576 7244 54778 7261
rect 55334 7261 55350 7278
rect 55780 7278 56368 7294
rect 55780 7261 55796 7278
rect 55334 7244 55536 7261
rect 54576 7206 55536 7244
rect 55594 7244 55796 7261
rect 56352 7261 56368 7278
rect 56798 7278 57386 7294
rect 56798 7261 56814 7278
rect 56352 7244 56554 7261
rect 55594 7206 56554 7244
rect 56612 7244 56814 7261
rect 57370 7261 57386 7278
rect 57816 7278 58404 7294
rect 57816 7261 57832 7278
rect 57370 7244 57572 7261
rect 56612 7206 57572 7244
rect 57630 7244 57832 7261
rect 58388 7261 58404 7278
rect 58834 7278 59422 7294
rect 58834 7261 58850 7278
rect 58388 7244 58590 7261
rect 57630 7206 58590 7244
rect 58648 7244 58850 7261
rect 59406 7261 59422 7278
rect 59852 7278 60440 7294
rect 59852 7261 59868 7278
rect 59406 7244 59608 7261
rect 58648 7206 59608 7244
rect 59666 7244 59868 7261
rect 60424 7261 60440 7278
rect 60870 7278 61458 7294
rect 60870 7261 60886 7278
rect 60424 7244 60626 7261
rect 59666 7206 60626 7244
rect 60684 7244 60886 7261
rect 61442 7261 61458 7278
rect 61888 7278 62476 7294
rect 61888 7261 61904 7278
rect 61442 7244 61644 7261
rect 60684 7206 61644 7244
rect 61702 7244 61904 7261
rect 62460 7261 62476 7278
rect 62906 7278 63494 7294
rect 62906 7261 62922 7278
rect 62460 7244 62662 7261
rect 61702 7206 62662 7244
rect 62720 7244 62922 7261
rect 63478 7261 63494 7278
rect 63924 7278 64512 7294
rect 63924 7261 63940 7278
rect 63478 7244 63680 7261
rect 62720 7206 63680 7244
rect 63738 7244 63940 7261
rect 64496 7261 64512 7278
rect 64942 7278 65530 7294
rect 64942 7261 64958 7278
rect 64496 7244 64698 7261
rect 63738 7206 64698 7244
rect 64756 7244 64958 7261
rect 65514 7261 65530 7278
rect 65960 7278 66548 7294
rect 65960 7261 65976 7278
rect 65514 7244 65716 7261
rect 64756 7206 65716 7244
rect 65774 7244 65976 7261
rect 66532 7261 66548 7278
rect 66978 7278 67566 7294
rect 66978 7261 66994 7278
rect 66532 7244 66734 7261
rect 65774 7206 66734 7244
rect 66792 7244 66994 7261
rect 67550 7261 67566 7278
rect 67996 7278 68584 7294
rect 67996 7261 68012 7278
rect 67550 7244 67752 7261
rect 66792 7206 67752 7244
rect 67810 7244 68012 7261
rect 68568 7261 68584 7278
rect 69014 7278 69602 7294
rect 69014 7261 69030 7278
rect 68568 7244 68770 7261
rect 67810 7206 68770 7244
rect 68828 7244 69030 7261
rect 69586 7261 69602 7278
rect 70032 7278 70620 7294
rect 70032 7261 70048 7278
rect 69586 7244 69788 7261
rect 68828 7206 69788 7244
rect 69846 7244 70048 7261
rect 70604 7261 70620 7278
rect 71050 7278 71638 7294
rect 71050 7261 71066 7278
rect 70604 7244 70806 7261
rect 69846 7206 70806 7244
rect 70864 7244 71066 7261
rect 71622 7261 71638 7278
rect 72068 7278 72656 7294
rect 72068 7261 72084 7278
rect 71622 7244 71824 7261
rect 70864 7206 71824 7244
rect 71882 7244 72084 7261
rect 72640 7261 72656 7278
rect 73086 7278 73674 7294
rect 73086 7261 73102 7278
rect 72640 7244 72842 7261
rect 71882 7206 72842 7244
rect 72900 7244 73102 7261
rect 73658 7261 73674 7278
rect 74104 7278 74692 7294
rect 74104 7261 74120 7278
rect 73658 7244 73860 7261
rect 72900 7206 73860 7244
rect 73918 7244 74120 7261
rect 74676 7261 74692 7278
rect 74676 7244 74878 7261
rect 73918 7206 74878 7244
rect 54576 6568 55536 6606
rect 54576 6551 54778 6568
rect 54762 6534 54778 6551
rect 55334 6551 55536 6568
rect 55594 6568 56554 6606
rect 55594 6551 55796 6568
rect 55334 6534 55350 6551
rect 54762 6518 55350 6534
rect 55780 6534 55796 6551
rect 56352 6551 56554 6568
rect 56612 6568 57572 6606
rect 56612 6551 56814 6568
rect 56352 6534 56368 6551
rect 55780 6518 56368 6534
rect 56798 6534 56814 6551
rect 57370 6551 57572 6568
rect 57630 6568 58590 6606
rect 57630 6551 57832 6568
rect 57370 6534 57386 6551
rect 56798 6518 57386 6534
rect 57816 6534 57832 6551
rect 58388 6551 58590 6568
rect 58648 6568 59608 6606
rect 58648 6551 58850 6568
rect 58388 6534 58404 6551
rect 57816 6518 58404 6534
rect 58834 6534 58850 6551
rect 59406 6551 59608 6568
rect 59666 6568 60626 6606
rect 59666 6551 59868 6568
rect 59406 6534 59422 6551
rect 58834 6518 59422 6534
rect 59852 6534 59868 6551
rect 60424 6551 60626 6568
rect 60684 6568 61644 6606
rect 60684 6551 60886 6568
rect 60424 6534 60440 6551
rect 59852 6518 60440 6534
rect 60870 6534 60886 6551
rect 61442 6551 61644 6568
rect 61702 6568 62662 6606
rect 61702 6551 61904 6568
rect 61442 6534 61458 6551
rect 60870 6518 61458 6534
rect 61888 6534 61904 6551
rect 62460 6551 62662 6568
rect 62720 6568 63680 6606
rect 62720 6551 62922 6568
rect 62460 6534 62476 6551
rect 61888 6518 62476 6534
rect 62906 6534 62922 6551
rect 63478 6551 63680 6568
rect 63738 6568 64698 6606
rect 63738 6551 63940 6568
rect 63478 6534 63494 6551
rect 62906 6518 63494 6534
rect 63924 6534 63940 6551
rect 64496 6551 64698 6568
rect 64756 6568 65716 6606
rect 64756 6551 64958 6568
rect 64496 6534 64512 6551
rect 63924 6518 64512 6534
rect 64942 6534 64958 6551
rect 65514 6551 65716 6568
rect 65774 6568 66734 6606
rect 65774 6551 65976 6568
rect 65514 6534 65530 6551
rect 64942 6518 65530 6534
rect 65960 6534 65976 6551
rect 66532 6551 66734 6568
rect 66792 6568 67752 6606
rect 66792 6551 66994 6568
rect 66532 6534 66548 6551
rect 65960 6518 66548 6534
rect 66978 6534 66994 6551
rect 67550 6551 67752 6568
rect 67810 6568 68770 6606
rect 67810 6551 68012 6568
rect 67550 6534 67566 6551
rect 66978 6518 67566 6534
rect 67996 6534 68012 6551
rect 68568 6551 68770 6568
rect 68828 6568 69788 6606
rect 68828 6551 69030 6568
rect 68568 6534 68584 6551
rect 67996 6518 68584 6534
rect 69014 6534 69030 6551
rect 69586 6551 69788 6568
rect 69846 6568 70806 6606
rect 69846 6551 70048 6568
rect 69586 6534 69602 6551
rect 69014 6518 69602 6534
rect 70032 6534 70048 6551
rect 70604 6551 70806 6568
rect 70864 6568 71824 6606
rect 70864 6551 71066 6568
rect 70604 6534 70620 6551
rect 70032 6518 70620 6534
rect 71050 6534 71066 6551
rect 71622 6551 71824 6568
rect 71882 6568 72842 6606
rect 71882 6551 72084 6568
rect 71622 6534 71638 6551
rect 71050 6518 71638 6534
rect 72068 6534 72084 6551
rect 72640 6551 72842 6568
rect 72900 6568 73860 6606
rect 72900 6551 73102 6568
rect 72640 6534 72656 6551
rect 72068 6518 72656 6534
rect 73086 6534 73102 6551
rect 73658 6551 73860 6568
rect 73918 6568 74878 6606
rect 73918 6551 74120 6568
rect 73658 6534 73674 6551
rect 73086 6518 73674 6534
rect 74104 6534 74120 6551
rect 74676 6551 74878 6568
rect 74676 6534 74692 6551
rect 74104 6518 74692 6534
rect 41674 6180 42262 6196
rect 41674 6163 41690 6180
rect 41488 6146 41690 6163
rect 42246 6163 42262 6180
rect 42692 6180 43280 6196
rect 42692 6163 42708 6180
rect 42246 6146 42448 6163
rect 41488 6108 42448 6146
rect 42506 6146 42708 6163
rect 43264 6163 43280 6180
rect 43710 6180 44298 6196
rect 43710 6163 43726 6180
rect 43264 6146 43466 6163
rect 42506 6108 43466 6146
rect 43524 6146 43726 6163
rect 44282 6163 44298 6180
rect 44728 6180 45316 6196
rect 44728 6163 44744 6180
rect 44282 6146 44484 6163
rect 43524 6108 44484 6146
rect 44542 6146 44744 6163
rect 45300 6163 45316 6180
rect 45746 6180 46334 6196
rect 45746 6163 45762 6180
rect 45300 6146 45502 6163
rect 44542 6108 45502 6146
rect 45560 6146 45762 6163
rect 46318 6163 46334 6180
rect 46764 6180 47352 6196
rect 46764 6163 46780 6180
rect 46318 6146 46520 6163
rect 45560 6108 46520 6146
rect 46578 6146 46780 6163
rect 47336 6163 47352 6180
rect 47782 6180 48370 6196
rect 47782 6163 47798 6180
rect 47336 6146 47538 6163
rect 46578 6108 47538 6146
rect 47596 6146 47798 6163
rect 48354 6163 48370 6180
rect 48800 6180 49388 6196
rect 48800 6163 48816 6180
rect 48354 6146 48556 6163
rect 47596 6108 48556 6146
rect 48614 6146 48816 6163
rect 49372 6163 49388 6180
rect 49818 6180 50406 6196
rect 49818 6163 49834 6180
rect 49372 6146 49574 6163
rect 48614 6108 49574 6146
rect 49632 6146 49834 6163
rect 50390 6163 50406 6180
rect 50836 6180 51424 6196
rect 50836 6163 50852 6180
rect 50390 6146 50592 6163
rect 49632 6108 50592 6146
rect 50650 6146 50852 6163
rect 51408 6163 51424 6180
rect 51854 6180 52442 6196
rect 51854 6163 51870 6180
rect 51408 6146 51610 6163
rect 50650 6108 51610 6146
rect 51668 6146 51870 6163
rect 52426 6163 52442 6180
rect 52426 6146 52628 6163
rect 51668 6108 52628 6146
rect 54762 6044 55350 6060
rect 54762 6027 54778 6044
rect 54576 6010 54778 6027
rect 55334 6027 55350 6044
rect 55780 6044 56368 6060
rect 55780 6027 55796 6044
rect 55334 6010 55536 6027
rect 54576 5972 55536 6010
rect 55594 6010 55796 6027
rect 56352 6027 56368 6044
rect 56798 6044 57386 6060
rect 56798 6027 56814 6044
rect 56352 6010 56554 6027
rect 55594 5972 56554 6010
rect 56612 6010 56814 6027
rect 57370 6027 57386 6044
rect 57816 6044 58404 6060
rect 57816 6027 57832 6044
rect 57370 6010 57572 6027
rect 56612 5972 57572 6010
rect 57630 6010 57832 6027
rect 58388 6027 58404 6044
rect 58834 6044 59422 6060
rect 58834 6027 58850 6044
rect 58388 6010 58590 6027
rect 57630 5972 58590 6010
rect 58648 6010 58850 6027
rect 59406 6027 59422 6044
rect 59852 6044 60440 6060
rect 59852 6027 59868 6044
rect 59406 6010 59608 6027
rect 58648 5972 59608 6010
rect 59666 6010 59868 6027
rect 60424 6027 60440 6044
rect 60870 6044 61458 6060
rect 60870 6027 60886 6044
rect 60424 6010 60626 6027
rect 59666 5972 60626 6010
rect 60684 6010 60886 6027
rect 61442 6027 61458 6044
rect 61888 6044 62476 6060
rect 61888 6027 61904 6044
rect 61442 6010 61644 6027
rect 60684 5972 61644 6010
rect 61702 6010 61904 6027
rect 62460 6027 62476 6044
rect 62906 6044 63494 6060
rect 62906 6027 62922 6044
rect 62460 6010 62662 6027
rect 61702 5972 62662 6010
rect 62720 6010 62922 6027
rect 63478 6027 63494 6044
rect 63924 6044 64512 6060
rect 63924 6027 63940 6044
rect 63478 6010 63680 6027
rect 62720 5972 63680 6010
rect 63738 6010 63940 6027
rect 64496 6027 64512 6044
rect 64942 6044 65530 6060
rect 64942 6027 64958 6044
rect 64496 6010 64698 6027
rect 63738 5972 64698 6010
rect 64756 6010 64958 6027
rect 65514 6027 65530 6044
rect 65960 6044 66548 6060
rect 65960 6027 65976 6044
rect 65514 6010 65716 6027
rect 64756 5972 65716 6010
rect 65774 6010 65976 6027
rect 66532 6027 66548 6044
rect 66978 6044 67566 6060
rect 66978 6027 66994 6044
rect 66532 6010 66734 6027
rect 65774 5972 66734 6010
rect 66792 6010 66994 6027
rect 67550 6027 67566 6044
rect 67996 6044 68584 6060
rect 67996 6027 68012 6044
rect 67550 6010 67752 6027
rect 66792 5972 67752 6010
rect 67810 6010 68012 6027
rect 68568 6027 68584 6044
rect 69014 6044 69602 6060
rect 69014 6027 69030 6044
rect 68568 6010 68770 6027
rect 67810 5972 68770 6010
rect 68828 6010 69030 6027
rect 69586 6027 69602 6044
rect 70032 6044 70620 6060
rect 70032 6027 70048 6044
rect 69586 6010 69788 6027
rect 68828 5972 69788 6010
rect 69846 6010 70048 6027
rect 70604 6027 70620 6044
rect 71050 6044 71638 6060
rect 71050 6027 71066 6044
rect 70604 6010 70806 6027
rect 69846 5972 70806 6010
rect 70864 6010 71066 6027
rect 71622 6027 71638 6044
rect 72068 6044 72656 6060
rect 72068 6027 72084 6044
rect 71622 6010 71824 6027
rect 70864 5972 71824 6010
rect 71882 6010 72084 6027
rect 72640 6027 72656 6044
rect 73086 6044 73674 6060
rect 73086 6027 73102 6044
rect 72640 6010 72842 6027
rect 71882 5972 72842 6010
rect 72900 6010 73102 6027
rect 73658 6027 73674 6044
rect 74104 6044 74692 6060
rect 74104 6027 74120 6044
rect 73658 6010 73860 6027
rect 72900 5972 73860 6010
rect 73918 6010 74120 6027
rect 74676 6027 74692 6044
rect 74676 6010 74878 6027
rect 73918 5972 74878 6010
rect 41488 5470 42448 5508
rect 41488 5453 41690 5470
rect 41674 5436 41690 5453
rect 42246 5453 42448 5470
rect 42506 5470 43466 5508
rect 42506 5453 42708 5470
rect 42246 5436 42262 5453
rect 41674 5420 42262 5436
rect 42692 5436 42708 5453
rect 43264 5453 43466 5470
rect 43524 5470 44484 5508
rect 43524 5453 43726 5470
rect 43264 5436 43280 5453
rect 42692 5420 43280 5436
rect 43710 5436 43726 5453
rect 44282 5453 44484 5470
rect 44542 5470 45502 5508
rect 44542 5453 44744 5470
rect 44282 5436 44298 5453
rect 43710 5420 44298 5436
rect 44728 5436 44744 5453
rect 45300 5453 45502 5470
rect 45560 5470 46520 5508
rect 45560 5453 45762 5470
rect 45300 5436 45316 5453
rect 44728 5420 45316 5436
rect 45746 5436 45762 5453
rect 46318 5453 46520 5470
rect 46578 5470 47538 5508
rect 46578 5453 46780 5470
rect 46318 5436 46334 5453
rect 45746 5420 46334 5436
rect 46764 5436 46780 5453
rect 47336 5453 47538 5470
rect 47596 5470 48556 5508
rect 47596 5453 47798 5470
rect 47336 5436 47352 5453
rect 46764 5420 47352 5436
rect 47782 5436 47798 5453
rect 48354 5453 48556 5470
rect 48614 5470 49574 5508
rect 48614 5453 48816 5470
rect 48354 5436 48370 5453
rect 47782 5420 48370 5436
rect 48800 5436 48816 5453
rect 49372 5453 49574 5470
rect 49632 5470 50592 5508
rect 49632 5453 49834 5470
rect 49372 5436 49388 5453
rect 48800 5420 49388 5436
rect 49818 5436 49834 5453
rect 50390 5453 50592 5470
rect 50650 5470 51610 5508
rect 50650 5453 50852 5470
rect 50390 5436 50406 5453
rect 49818 5420 50406 5436
rect 50836 5436 50852 5453
rect 51408 5453 51610 5470
rect 51668 5470 52628 5508
rect 51668 5453 51870 5470
rect 51408 5436 51424 5453
rect 50836 5420 51424 5436
rect 51854 5436 51870 5453
rect 52426 5453 52628 5470
rect 52426 5436 52442 5453
rect 51854 5420 52442 5436
rect 54576 5334 55536 5372
rect 54576 5317 54778 5334
rect 54762 5300 54778 5317
rect 55334 5317 55536 5334
rect 55594 5334 56554 5372
rect 55594 5317 55796 5334
rect 55334 5300 55350 5317
rect 54762 5284 55350 5300
rect 55780 5300 55796 5317
rect 56352 5317 56554 5334
rect 56612 5334 57572 5372
rect 56612 5317 56814 5334
rect 56352 5300 56368 5317
rect 55780 5284 56368 5300
rect 56798 5300 56814 5317
rect 57370 5317 57572 5334
rect 57630 5334 58590 5372
rect 57630 5317 57832 5334
rect 57370 5300 57386 5317
rect 56798 5284 57386 5300
rect 57816 5300 57832 5317
rect 58388 5317 58590 5334
rect 58648 5334 59608 5372
rect 58648 5317 58850 5334
rect 58388 5300 58404 5317
rect 57816 5284 58404 5300
rect 58834 5300 58850 5317
rect 59406 5317 59608 5334
rect 59666 5334 60626 5372
rect 59666 5317 59868 5334
rect 59406 5300 59422 5317
rect 58834 5284 59422 5300
rect 59852 5300 59868 5317
rect 60424 5317 60626 5334
rect 60684 5334 61644 5372
rect 60684 5317 60886 5334
rect 60424 5300 60440 5317
rect 59852 5284 60440 5300
rect 60870 5300 60886 5317
rect 61442 5317 61644 5334
rect 61702 5334 62662 5372
rect 61702 5317 61904 5334
rect 61442 5300 61458 5317
rect 60870 5284 61458 5300
rect 61888 5300 61904 5317
rect 62460 5317 62662 5334
rect 62720 5334 63680 5372
rect 62720 5317 62922 5334
rect 62460 5300 62476 5317
rect 61888 5284 62476 5300
rect 62906 5300 62922 5317
rect 63478 5317 63680 5334
rect 63738 5334 64698 5372
rect 63738 5317 63940 5334
rect 63478 5300 63494 5317
rect 62906 5284 63494 5300
rect 63924 5300 63940 5317
rect 64496 5317 64698 5334
rect 64756 5334 65716 5372
rect 64756 5317 64958 5334
rect 64496 5300 64512 5317
rect 63924 5284 64512 5300
rect 64942 5300 64958 5317
rect 65514 5317 65716 5334
rect 65774 5334 66734 5372
rect 65774 5317 65976 5334
rect 65514 5300 65530 5317
rect 64942 5284 65530 5300
rect 65960 5300 65976 5317
rect 66532 5317 66734 5334
rect 66792 5334 67752 5372
rect 66792 5317 66994 5334
rect 66532 5300 66548 5317
rect 65960 5284 66548 5300
rect 66978 5300 66994 5317
rect 67550 5317 67752 5334
rect 67810 5334 68770 5372
rect 67810 5317 68012 5334
rect 67550 5300 67566 5317
rect 66978 5284 67566 5300
rect 67996 5300 68012 5317
rect 68568 5317 68770 5334
rect 68828 5334 69788 5372
rect 68828 5317 69030 5334
rect 68568 5300 68584 5317
rect 67996 5284 68584 5300
rect 69014 5300 69030 5317
rect 69586 5317 69788 5334
rect 69846 5334 70806 5372
rect 69846 5317 70048 5334
rect 69586 5300 69602 5317
rect 69014 5284 69602 5300
rect 70032 5300 70048 5317
rect 70604 5317 70806 5334
rect 70864 5334 71824 5372
rect 70864 5317 71066 5334
rect 70604 5300 70620 5317
rect 70032 5284 70620 5300
rect 71050 5300 71066 5317
rect 71622 5317 71824 5334
rect 71882 5334 72842 5372
rect 71882 5317 72084 5334
rect 71622 5300 71638 5317
rect 71050 5284 71638 5300
rect 72068 5300 72084 5317
rect 72640 5317 72842 5334
rect 72900 5334 73860 5372
rect 72900 5317 73102 5334
rect 72640 5300 72656 5317
rect 72068 5284 72656 5300
rect 73086 5300 73102 5317
rect 73658 5317 73860 5334
rect 73918 5334 74878 5372
rect 73918 5317 74120 5334
rect 73658 5300 73674 5317
rect 73086 5284 73674 5300
rect 74104 5300 74120 5317
rect 74676 5317 74878 5334
rect 74676 5300 74692 5317
rect 74104 5284 74692 5300
rect 41674 5068 42262 5084
rect 41674 5051 41690 5068
rect 41488 5034 41690 5051
rect 42246 5051 42262 5068
rect 42692 5068 43280 5084
rect 42692 5051 42708 5068
rect 42246 5034 42448 5051
rect 41488 4996 42448 5034
rect 42506 5034 42708 5051
rect 43264 5051 43280 5068
rect 43710 5068 44298 5084
rect 43710 5051 43726 5068
rect 43264 5034 43466 5051
rect 42506 4996 43466 5034
rect 43524 5034 43726 5051
rect 44282 5051 44298 5068
rect 44728 5068 45316 5084
rect 44728 5051 44744 5068
rect 44282 5034 44484 5051
rect 43524 4996 44484 5034
rect 44542 5034 44744 5051
rect 45300 5051 45316 5068
rect 45746 5068 46334 5084
rect 45746 5051 45762 5068
rect 45300 5034 45502 5051
rect 44542 4996 45502 5034
rect 45560 5034 45762 5051
rect 46318 5051 46334 5068
rect 46764 5068 47352 5084
rect 46764 5051 46780 5068
rect 46318 5034 46520 5051
rect 45560 4996 46520 5034
rect 46578 5034 46780 5051
rect 47336 5051 47352 5068
rect 47782 5068 48370 5084
rect 47782 5051 47798 5068
rect 47336 5034 47538 5051
rect 46578 4996 47538 5034
rect 47596 5034 47798 5051
rect 48354 5051 48370 5068
rect 48800 5068 49388 5084
rect 48800 5051 48816 5068
rect 48354 5034 48556 5051
rect 47596 4996 48556 5034
rect 48614 5034 48816 5051
rect 49372 5051 49388 5068
rect 49818 5068 50406 5084
rect 49818 5051 49834 5068
rect 49372 5034 49574 5051
rect 48614 4996 49574 5034
rect 49632 5034 49834 5051
rect 50390 5051 50406 5068
rect 50836 5068 51424 5084
rect 50836 5051 50852 5068
rect 50390 5034 50592 5051
rect 49632 4996 50592 5034
rect 50650 5034 50852 5051
rect 51408 5051 51424 5068
rect 51854 5068 52442 5084
rect 51854 5051 51870 5068
rect 51408 5034 51610 5051
rect 50650 4996 51610 5034
rect 51668 5034 51870 5051
rect 52426 5051 52442 5068
rect 52426 5034 52628 5051
rect 51668 4996 52628 5034
rect 54762 4810 55350 4826
rect 54762 4793 54778 4810
rect 54576 4776 54778 4793
rect 55334 4793 55350 4810
rect 55780 4810 56368 4826
rect 55780 4793 55796 4810
rect 55334 4776 55536 4793
rect 54576 4738 55536 4776
rect 55594 4776 55796 4793
rect 56352 4793 56368 4810
rect 56798 4810 57386 4826
rect 56798 4793 56814 4810
rect 56352 4776 56554 4793
rect 55594 4738 56554 4776
rect 56612 4776 56814 4793
rect 57370 4793 57386 4810
rect 57816 4810 58404 4826
rect 57816 4793 57832 4810
rect 57370 4776 57572 4793
rect 56612 4738 57572 4776
rect 57630 4776 57832 4793
rect 58388 4793 58404 4810
rect 58834 4810 59422 4826
rect 58834 4793 58850 4810
rect 58388 4776 58590 4793
rect 57630 4738 58590 4776
rect 58648 4776 58850 4793
rect 59406 4793 59422 4810
rect 59852 4810 60440 4826
rect 59852 4793 59868 4810
rect 59406 4776 59608 4793
rect 58648 4738 59608 4776
rect 59666 4776 59868 4793
rect 60424 4793 60440 4810
rect 60870 4810 61458 4826
rect 60870 4793 60886 4810
rect 60424 4776 60626 4793
rect 59666 4738 60626 4776
rect 60684 4776 60886 4793
rect 61442 4793 61458 4810
rect 61888 4810 62476 4826
rect 61888 4793 61904 4810
rect 61442 4776 61644 4793
rect 60684 4738 61644 4776
rect 61702 4776 61904 4793
rect 62460 4793 62476 4810
rect 62906 4810 63494 4826
rect 62906 4793 62922 4810
rect 62460 4776 62662 4793
rect 61702 4738 62662 4776
rect 62720 4776 62922 4793
rect 63478 4793 63494 4810
rect 63924 4810 64512 4826
rect 63924 4793 63940 4810
rect 63478 4776 63680 4793
rect 62720 4738 63680 4776
rect 63738 4776 63940 4793
rect 64496 4793 64512 4810
rect 64942 4810 65530 4826
rect 64942 4793 64958 4810
rect 64496 4776 64698 4793
rect 63738 4738 64698 4776
rect 64756 4776 64958 4793
rect 65514 4793 65530 4810
rect 65960 4810 66548 4826
rect 65960 4793 65976 4810
rect 65514 4776 65716 4793
rect 64756 4738 65716 4776
rect 65774 4776 65976 4793
rect 66532 4793 66548 4810
rect 66978 4810 67566 4826
rect 66978 4793 66994 4810
rect 66532 4776 66734 4793
rect 65774 4738 66734 4776
rect 66792 4776 66994 4793
rect 67550 4793 67566 4810
rect 67996 4810 68584 4826
rect 67996 4793 68012 4810
rect 67550 4776 67752 4793
rect 66792 4738 67752 4776
rect 67810 4776 68012 4793
rect 68568 4793 68584 4810
rect 69014 4810 69602 4826
rect 69014 4793 69030 4810
rect 68568 4776 68770 4793
rect 67810 4738 68770 4776
rect 68828 4776 69030 4793
rect 69586 4793 69602 4810
rect 70032 4810 70620 4826
rect 70032 4793 70048 4810
rect 69586 4776 69788 4793
rect 68828 4738 69788 4776
rect 69846 4776 70048 4793
rect 70604 4793 70620 4810
rect 71050 4810 71638 4826
rect 71050 4793 71066 4810
rect 70604 4776 70806 4793
rect 69846 4738 70806 4776
rect 70864 4776 71066 4793
rect 71622 4793 71638 4810
rect 72068 4810 72656 4826
rect 72068 4793 72084 4810
rect 71622 4776 71824 4793
rect 70864 4738 71824 4776
rect 71882 4776 72084 4793
rect 72640 4793 72656 4810
rect 73086 4810 73674 4826
rect 73086 4793 73102 4810
rect 72640 4776 72842 4793
rect 71882 4738 72842 4776
rect 72900 4776 73102 4793
rect 73658 4793 73674 4810
rect 74104 4810 74692 4826
rect 74104 4793 74120 4810
rect 73658 4776 73860 4793
rect 72900 4738 73860 4776
rect 73918 4776 74120 4793
rect 74676 4793 74692 4810
rect 74676 4776 74878 4793
rect 73918 4738 74878 4776
rect 41488 4358 42448 4396
rect 41488 4341 41690 4358
rect 41674 4324 41690 4341
rect 42246 4341 42448 4358
rect 42506 4358 43466 4396
rect 42506 4341 42708 4358
rect 42246 4324 42262 4341
rect 41674 4308 42262 4324
rect 42692 4324 42708 4341
rect 43264 4341 43466 4358
rect 43524 4358 44484 4396
rect 43524 4341 43726 4358
rect 43264 4324 43280 4341
rect 42692 4308 43280 4324
rect 43710 4324 43726 4341
rect 44282 4341 44484 4358
rect 44542 4358 45502 4396
rect 44542 4341 44744 4358
rect 44282 4324 44298 4341
rect 43710 4308 44298 4324
rect 44728 4324 44744 4341
rect 45300 4341 45502 4358
rect 45560 4358 46520 4396
rect 45560 4341 45762 4358
rect 45300 4324 45316 4341
rect 44728 4308 45316 4324
rect 45746 4324 45762 4341
rect 46318 4341 46520 4358
rect 46578 4358 47538 4396
rect 46578 4341 46780 4358
rect 46318 4324 46334 4341
rect 45746 4308 46334 4324
rect 46764 4324 46780 4341
rect 47336 4341 47538 4358
rect 47596 4358 48556 4396
rect 47596 4341 47798 4358
rect 47336 4324 47352 4341
rect 46764 4308 47352 4324
rect 47782 4324 47798 4341
rect 48354 4341 48556 4358
rect 48614 4358 49574 4396
rect 48614 4341 48816 4358
rect 48354 4324 48370 4341
rect 47782 4308 48370 4324
rect 48800 4324 48816 4341
rect 49372 4341 49574 4358
rect 49632 4358 50592 4396
rect 49632 4341 49834 4358
rect 49372 4324 49388 4341
rect 48800 4308 49388 4324
rect 49818 4324 49834 4341
rect 50390 4341 50592 4358
rect 50650 4358 51610 4396
rect 50650 4341 50852 4358
rect 50390 4324 50406 4341
rect 49818 4308 50406 4324
rect 50836 4324 50852 4341
rect 51408 4341 51610 4358
rect 51668 4358 52628 4396
rect 51668 4341 51870 4358
rect 51408 4324 51424 4341
rect 50836 4308 51424 4324
rect 51854 4324 51870 4341
rect 52426 4341 52628 4358
rect 52426 4324 52442 4341
rect 51854 4308 52442 4324
rect 54576 4100 55536 4138
rect 54576 4083 54778 4100
rect 54762 4066 54778 4083
rect 55334 4083 55536 4100
rect 55594 4100 56554 4138
rect 55594 4083 55796 4100
rect 55334 4066 55350 4083
rect 54762 4050 55350 4066
rect 55780 4066 55796 4083
rect 56352 4083 56554 4100
rect 56612 4100 57572 4138
rect 56612 4083 56814 4100
rect 56352 4066 56368 4083
rect 55780 4050 56368 4066
rect 56798 4066 56814 4083
rect 57370 4083 57572 4100
rect 57630 4100 58590 4138
rect 57630 4083 57832 4100
rect 57370 4066 57386 4083
rect 56798 4050 57386 4066
rect 57816 4066 57832 4083
rect 58388 4083 58590 4100
rect 58648 4100 59608 4138
rect 58648 4083 58850 4100
rect 58388 4066 58404 4083
rect 57816 4050 58404 4066
rect 58834 4066 58850 4083
rect 59406 4083 59608 4100
rect 59666 4100 60626 4138
rect 59666 4083 59868 4100
rect 59406 4066 59422 4083
rect 58834 4050 59422 4066
rect 59852 4066 59868 4083
rect 60424 4083 60626 4100
rect 60684 4100 61644 4138
rect 60684 4083 60886 4100
rect 60424 4066 60440 4083
rect 59852 4050 60440 4066
rect 60870 4066 60886 4083
rect 61442 4083 61644 4100
rect 61702 4100 62662 4138
rect 61702 4083 61904 4100
rect 61442 4066 61458 4083
rect 60870 4050 61458 4066
rect 61888 4066 61904 4083
rect 62460 4083 62662 4100
rect 62720 4100 63680 4138
rect 62720 4083 62922 4100
rect 62460 4066 62476 4083
rect 61888 4050 62476 4066
rect 62906 4066 62922 4083
rect 63478 4083 63680 4100
rect 63738 4100 64698 4138
rect 63738 4083 63940 4100
rect 63478 4066 63494 4083
rect 62906 4050 63494 4066
rect 63924 4066 63940 4083
rect 64496 4083 64698 4100
rect 64756 4100 65716 4138
rect 64756 4083 64958 4100
rect 64496 4066 64512 4083
rect 63924 4050 64512 4066
rect 64942 4066 64958 4083
rect 65514 4083 65716 4100
rect 65774 4100 66734 4138
rect 65774 4083 65976 4100
rect 65514 4066 65530 4083
rect 64942 4050 65530 4066
rect 65960 4066 65976 4083
rect 66532 4083 66734 4100
rect 66792 4100 67752 4138
rect 66792 4083 66994 4100
rect 66532 4066 66548 4083
rect 65960 4050 66548 4066
rect 66978 4066 66994 4083
rect 67550 4083 67752 4100
rect 67810 4100 68770 4138
rect 67810 4083 68012 4100
rect 67550 4066 67566 4083
rect 66978 4050 67566 4066
rect 67996 4066 68012 4083
rect 68568 4083 68770 4100
rect 68828 4100 69788 4138
rect 68828 4083 69030 4100
rect 68568 4066 68584 4083
rect 67996 4050 68584 4066
rect 69014 4066 69030 4083
rect 69586 4083 69788 4100
rect 69846 4100 70806 4138
rect 69846 4083 70048 4100
rect 69586 4066 69602 4083
rect 69014 4050 69602 4066
rect 70032 4066 70048 4083
rect 70604 4083 70806 4100
rect 70864 4100 71824 4138
rect 70864 4083 71066 4100
rect 70604 4066 70620 4083
rect 70032 4050 70620 4066
rect 71050 4066 71066 4083
rect 71622 4083 71824 4100
rect 71882 4100 72842 4138
rect 71882 4083 72084 4100
rect 71622 4066 71638 4083
rect 71050 4050 71638 4066
rect 72068 4066 72084 4083
rect 72640 4083 72842 4100
rect 72900 4100 73860 4138
rect 72900 4083 73102 4100
rect 72640 4066 72656 4083
rect 72068 4050 72656 4066
rect 73086 4066 73102 4083
rect 73658 4083 73860 4100
rect 73918 4100 74878 4138
rect 73918 4083 74120 4100
rect 73658 4066 73674 4083
rect 73086 4050 73674 4066
rect 74104 4066 74120 4083
rect 74676 4083 74878 4100
rect 74676 4066 74692 4083
rect 74104 4050 74692 4066
rect 41674 3956 42262 3972
rect 41674 3939 41690 3956
rect 41488 3922 41690 3939
rect 42246 3939 42262 3956
rect 42692 3956 43280 3972
rect 42692 3939 42708 3956
rect 42246 3922 42448 3939
rect 41488 3884 42448 3922
rect 42506 3922 42708 3939
rect 43264 3939 43280 3956
rect 43710 3956 44298 3972
rect 43710 3939 43726 3956
rect 43264 3922 43466 3939
rect 42506 3884 43466 3922
rect 43524 3922 43726 3939
rect 44282 3939 44298 3956
rect 44728 3956 45316 3972
rect 44728 3939 44744 3956
rect 44282 3922 44484 3939
rect 43524 3884 44484 3922
rect 44542 3922 44744 3939
rect 45300 3939 45316 3956
rect 45746 3956 46334 3972
rect 45746 3939 45762 3956
rect 45300 3922 45502 3939
rect 44542 3884 45502 3922
rect 45560 3922 45762 3939
rect 46318 3939 46334 3956
rect 46764 3956 47352 3972
rect 46764 3939 46780 3956
rect 46318 3922 46520 3939
rect 45560 3884 46520 3922
rect 46578 3922 46780 3939
rect 47336 3939 47352 3956
rect 47782 3956 48370 3972
rect 47782 3939 47798 3956
rect 47336 3922 47538 3939
rect 46578 3884 47538 3922
rect 47596 3922 47798 3939
rect 48354 3939 48370 3956
rect 48800 3956 49388 3972
rect 48800 3939 48816 3956
rect 48354 3922 48556 3939
rect 47596 3884 48556 3922
rect 48614 3922 48816 3939
rect 49372 3939 49388 3956
rect 49818 3956 50406 3972
rect 49818 3939 49834 3956
rect 49372 3922 49574 3939
rect 48614 3884 49574 3922
rect 49632 3922 49834 3939
rect 50390 3939 50406 3956
rect 50836 3956 51424 3972
rect 50836 3939 50852 3956
rect 50390 3922 50592 3939
rect 49632 3884 50592 3922
rect 50650 3922 50852 3939
rect 51408 3939 51424 3956
rect 51854 3956 52442 3972
rect 51854 3939 51870 3956
rect 51408 3922 51610 3939
rect 50650 3884 51610 3922
rect 51668 3922 51870 3939
rect 52426 3939 52442 3956
rect 52426 3922 52628 3939
rect 51668 3884 52628 3922
rect 54762 3578 55350 3594
rect 54762 3561 54778 3578
rect 54576 3544 54778 3561
rect 55334 3561 55350 3578
rect 55780 3578 56368 3594
rect 55780 3561 55796 3578
rect 55334 3544 55536 3561
rect 54576 3506 55536 3544
rect 55594 3544 55796 3561
rect 56352 3561 56368 3578
rect 56798 3578 57386 3594
rect 56798 3561 56814 3578
rect 56352 3544 56554 3561
rect 55594 3506 56554 3544
rect 56612 3544 56814 3561
rect 57370 3561 57386 3578
rect 57816 3578 58404 3594
rect 57816 3561 57832 3578
rect 57370 3544 57572 3561
rect 56612 3506 57572 3544
rect 57630 3544 57832 3561
rect 58388 3561 58404 3578
rect 58834 3578 59422 3594
rect 58834 3561 58850 3578
rect 58388 3544 58590 3561
rect 57630 3506 58590 3544
rect 58648 3544 58850 3561
rect 59406 3561 59422 3578
rect 59852 3578 60440 3594
rect 59852 3561 59868 3578
rect 59406 3544 59608 3561
rect 58648 3506 59608 3544
rect 59666 3544 59868 3561
rect 60424 3561 60440 3578
rect 60870 3578 61458 3594
rect 60870 3561 60886 3578
rect 60424 3544 60626 3561
rect 59666 3506 60626 3544
rect 60684 3544 60886 3561
rect 61442 3561 61458 3578
rect 61888 3578 62476 3594
rect 61888 3561 61904 3578
rect 61442 3544 61644 3561
rect 60684 3506 61644 3544
rect 61702 3544 61904 3561
rect 62460 3561 62476 3578
rect 62906 3578 63494 3594
rect 62906 3561 62922 3578
rect 62460 3544 62662 3561
rect 61702 3506 62662 3544
rect 62720 3544 62922 3561
rect 63478 3561 63494 3578
rect 63924 3578 64512 3594
rect 63924 3561 63940 3578
rect 63478 3544 63680 3561
rect 62720 3506 63680 3544
rect 63738 3544 63940 3561
rect 64496 3561 64512 3578
rect 64942 3578 65530 3594
rect 64942 3561 64958 3578
rect 64496 3544 64698 3561
rect 63738 3506 64698 3544
rect 64756 3544 64958 3561
rect 65514 3561 65530 3578
rect 65960 3578 66548 3594
rect 65960 3561 65976 3578
rect 65514 3544 65716 3561
rect 64756 3506 65716 3544
rect 65774 3544 65976 3561
rect 66532 3561 66548 3578
rect 66978 3578 67566 3594
rect 66978 3561 66994 3578
rect 66532 3544 66734 3561
rect 65774 3506 66734 3544
rect 66792 3544 66994 3561
rect 67550 3561 67566 3578
rect 67996 3578 68584 3594
rect 67996 3561 68012 3578
rect 67550 3544 67752 3561
rect 66792 3506 67752 3544
rect 67810 3544 68012 3561
rect 68568 3561 68584 3578
rect 69014 3578 69602 3594
rect 69014 3561 69030 3578
rect 68568 3544 68770 3561
rect 67810 3506 68770 3544
rect 68828 3544 69030 3561
rect 69586 3561 69602 3578
rect 70032 3578 70620 3594
rect 70032 3561 70048 3578
rect 69586 3544 69788 3561
rect 68828 3506 69788 3544
rect 69846 3544 70048 3561
rect 70604 3561 70620 3578
rect 71050 3578 71638 3594
rect 71050 3561 71066 3578
rect 70604 3544 70806 3561
rect 69846 3506 70806 3544
rect 70864 3544 71066 3561
rect 71622 3561 71638 3578
rect 72068 3578 72656 3594
rect 72068 3561 72084 3578
rect 71622 3544 71824 3561
rect 70864 3506 71824 3544
rect 71882 3544 72084 3561
rect 72640 3561 72656 3578
rect 73086 3578 73674 3594
rect 73086 3561 73102 3578
rect 72640 3544 72842 3561
rect 71882 3506 72842 3544
rect 72900 3544 73102 3561
rect 73658 3561 73674 3578
rect 74104 3578 74692 3594
rect 74104 3561 74120 3578
rect 73658 3544 73860 3561
rect 72900 3506 73860 3544
rect 73918 3544 74120 3561
rect 74676 3561 74692 3578
rect 74676 3544 74878 3561
rect 73918 3506 74878 3544
rect 41488 3246 42448 3284
rect 41488 3229 41690 3246
rect 41674 3212 41690 3229
rect 42246 3229 42448 3246
rect 42506 3246 43466 3284
rect 42506 3229 42708 3246
rect 42246 3212 42262 3229
rect 41674 3196 42262 3212
rect 42692 3212 42708 3229
rect 43264 3229 43466 3246
rect 43524 3246 44484 3284
rect 43524 3229 43726 3246
rect 43264 3212 43280 3229
rect 42692 3196 43280 3212
rect 43710 3212 43726 3229
rect 44282 3229 44484 3246
rect 44542 3246 45502 3284
rect 44542 3229 44744 3246
rect 44282 3212 44298 3229
rect 43710 3196 44298 3212
rect 44728 3212 44744 3229
rect 45300 3229 45502 3246
rect 45560 3246 46520 3284
rect 45560 3229 45762 3246
rect 45300 3212 45316 3229
rect 44728 3196 45316 3212
rect 45746 3212 45762 3229
rect 46318 3229 46520 3246
rect 46578 3246 47538 3284
rect 46578 3229 46780 3246
rect 46318 3212 46334 3229
rect 45746 3196 46334 3212
rect 46764 3212 46780 3229
rect 47336 3229 47538 3246
rect 47596 3246 48556 3284
rect 47596 3229 47798 3246
rect 47336 3212 47352 3229
rect 46764 3196 47352 3212
rect 47782 3212 47798 3229
rect 48354 3229 48556 3246
rect 48614 3246 49574 3284
rect 48614 3229 48816 3246
rect 48354 3212 48370 3229
rect 47782 3196 48370 3212
rect 48800 3212 48816 3229
rect 49372 3229 49574 3246
rect 49632 3246 50592 3284
rect 49632 3229 49834 3246
rect 49372 3212 49388 3229
rect 48800 3196 49388 3212
rect 49818 3212 49834 3229
rect 50390 3229 50592 3246
rect 50650 3246 51610 3284
rect 50650 3229 50852 3246
rect 50390 3212 50406 3229
rect 49818 3196 50406 3212
rect 50836 3212 50852 3229
rect 51408 3229 51610 3246
rect 51668 3246 52628 3284
rect 51668 3229 51870 3246
rect 51408 3212 51424 3229
rect 50836 3196 51424 3212
rect 51854 3212 51870 3229
rect 52426 3229 52628 3246
rect 52426 3212 52442 3229
rect 51854 3196 52442 3212
rect 54576 2868 55536 2906
rect 41674 2844 42262 2860
rect 41674 2827 41690 2844
rect 41488 2810 41690 2827
rect 42246 2827 42262 2844
rect 42692 2844 43280 2860
rect 42692 2827 42708 2844
rect 42246 2810 42448 2827
rect 41488 2772 42448 2810
rect 42506 2810 42708 2827
rect 43264 2827 43280 2844
rect 43710 2844 44298 2860
rect 43710 2827 43726 2844
rect 43264 2810 43466 2827
rect 42506 2772 43466 2810
rect 43524 2810 43726 2827
rect 44282 2827 44298 2844
rect 44728 2844 45316 2860
rect 44728 2827 44744 2844
rect 44282 2810 44484 2827
rect 43524 2772 44484 2810
rect 44542 2810 44744 2827
rect 45300 2827 45316 2844
rect 45746 2844 46334 2860
rect 45746 2827 45762 2844
rect 45300 2810 45502 2827
rect 44542 2772 45502 2810
rect 45560 2810 45762 2827
rect 46318 2827 46334 2844
rect 46764 2844 47352 2860
rect 46764 2827 46780 2844
rect 46318 2810 46520 2827
rect 45560 2772 46520 2810
rect 46578 2810 46780 2827
rect 47336 2827 47352 2844
rect 47782 2844 48370 2860
rect 47782 2827 47798 2844
rect 47336 2810 47538 2827
rect 46578 2772 47538 2810
rect 47596 2810 47798 2827
rect 48354 2827 48370 2844
rect 48800 2844 49388 2860
rect 48800 2827 48816 2844
rect 48354 2810 48556 2827
rect 47596 2772 48556 2810
rect 48614 2810 48816 2827
rect 49372 2827 49388 2844
rect 49818 2844 50406 2860
rect 49818 2827 49834 2844
rect 49372 2810 49574 2827
rect 48614 2772 49574 2810
rect 49632 2810 49834 2827
rect 50390 2827 50406 2844
rect 50836 2844 51424 2860
rect 50836 2827 50852 2844
rect 50390 2810 50592 2827
rect 49632 2772 50592 2810
rect 50650 2810 50852 2827
rect 51408 2827 51424 2844
rect 51854 2844 52442 2860
rect 54576 2851 54778 2868
rect 51854 2827 51870 2844
rect 51408 2810 51610 2827
rect 50650 2772 51610 2810
rect 51668 2810 51870 2827
rect 52426 2827 52442 2844
rect 54762 2834 54778 2851
rect 55334 2851 55536 2868
rect 55594 2868 56554 2906
rect 55594 2851 55796 2868
rect 55334 2834 55350 2851
rect 52426 2810 52628 2827
rect 54762 2818 55350 2834
rect 55780 2834 55796 2851
rect 56352 2851 56554 2868
rect 56612 2868 57572 2906
rect 56612 2851 56814 2868
rect 56352 2834 56368 2851
rect 55780 2818 56368 2834
rect 56798 2834 56814 2851
rect 57370 2851 57572 2868
rect 57630 2868 58590 2906
rect 57630 2851 57832 2868
rect 57370 2834 57386 2851
rect 56798 2818 57386 2834
rect 57816 2834 57832 2851
rect 58388 2851 58590 2868
rect 58648 2868 59608 2906
rect 58648 2851 58850 2868
rect 58388 2834 58404 2851
rect 57816 2818 58404 2834
rect 58834 2834 58850 2851
rect 59406 2851 59608 2868
rect 59666 2868 60626 2906
rect 59666 2851 59868 2868
rect 59406 2834 59422 2851
rect 58834 2818 59422 2834
rect 59852 2834 59868 2851
rect 60424 2851 60626 2868
rect 60684 2868 61644 2906
rect 60684 2851 60886 2868
rect 60424 2834 60440 2851
rect 59852 2818 60440 2834
rect 60870 2834 60886 2851
rect 61442 2851 61644 2868
rect 61702 2868 62662 2906
rect 61702 2851 61904 2868
rect 61442 2834 61458 2851
rect 60870 2818 61458 2834
rect 61888 2834 61904 2851
rect 62460 2851 62662 2868
rect 62720 2868 63680 2906
rect 62720 2851 62922 2868
rect 62460 2834 62476 2851
rect 61888 2818 62476 2834
rect 62906 2834 62922 2851
rect 63478 2851 63680 2868
rect 63738 2868 64698 2906
rect 63738 2851 63940 2868
rect 63478 2834 63494 2851
rect 62906 2818 63494 2834
rect 63924 2834 63940 2851
rect 64496 2851 64698 2868
rect 64756 2868 65716 2906
rect 64756 2851 64958 2868
rect 64496 2834 64512 2851
rect 63924 2818 64512 2834
rect 64942 2834 64958 2851
rect 65514 2851 65716 2868
rect 65774 2868 66734 2906
rect 65774 2851 65976 2868
rect 65514 2834 65530 2851
rect 64942 2818 65530 2834
rect 65960 2834 65976 2851
rect 66532 2851 66734 2868
rect 66792 2868 67752 2906
rect 66792 2851 66994 2868
rect 66532 2834 66548 2851
rect 65960 2818 66548 2834
rect 66978 2834 66994 2851
rect 67550 2851 67752 2868
rect 67810 2868 68770 2906
rect 67810 2851 68012 2868
rect 67550 2834 67566 2851
rect 66978 2818 67566 2834
rect 67996 2834 68012 2851
rect 68568 2851 68770 2868
rect 68828 2868 69788 2906
rect 68828 2851 69030 2868
rect 68568 2834 68584 2851
rect 67996 2818 68584 2834
rect 69014 2834 69030 2851
rect 69586 2851 69788 2868
rect 69846 2868 70806 2906
rect 69846 2851 70048 2868
rect 69586 2834 69602 2851
rect 69014 2818 69602 2834
rect 70032 2834 70048 2851
rect 70604 2851 70806 2868
rect 70864 2868 71824 2906
rect 70864 2851 71066 2868
rect 70604 2834 70620 2851
rect 70032 2818 70620 2834
rect 71050 2834 71066 2851
rect 71622 2851 71824 2868
rect 71882 2868 72842 2906
rect 71882 2851 72084 2868
rect 71622 2834 71638 2851
rect 71050 2818 71638 2834
rect 72068 2834 72084 2851
rect 72640 2851 72842 2868
rect 72900 2868 73860 2906
rect 72900 2851 73102 2868
rect 72640 2834 72656 2851
rect 72068 2818 72656 2834
rect 73086 2834 73102 2851
rect 73658 2851 73860 2868
rect 73918 2868 74878 2906
rect 73918 2851 74120 2868
rect 73658 2834 73674 2851
rect 73086 2818 73674 2834
rect 74104 2834 74120 2851
rect 74676 2851 74878 2868
rect 74676 2834 74692 2851
rect 74104 2818 74692 2834
rect 51668 2772 52628 2810
rect 54762 2344 55350 2360
rect 54762 2327 54778 2344
rect 54576 2310 54778 2327
rect 55334 2327 55350 2344
rect 55780 2344 56368 2360
rect 55780 2327 55796 2344
rect 55334 2310 55536 2327
rect 54576 2272 55536 2310
rect 55594 2310 55796 2327
rect 56352 2327 56368 2344
rect 56798 2344 57386 2360
rect 56798 2327 56814 2344
rect 56352 2310 56554 2327
rect 55594 2272 56554 2310
rect 56612 2310 56814 2327
rect 57370 2327 57386 2344
rect 57816 2344 58404 2360
rect 57816 2327 57832 2344
rect 57370 2310 57572 2327
rect 56612 2272 57572 2310
rect 57630 2310 57832 2327
rect 58388 2327 58404 2344
rect 58834 2344 59422 2360
rect 58834 2327 58850 2344
rect 58388 2310 58590 2327
rect 57630 2272 58590 2310
rect 58648 2310 58850 2327
rect 59406 2327 59422 2344
rect 59852 2344 60440 2360
rect 59852 2327 59868 2344
rect 59406 2310 59608 2327
rect 58648 2272 59608 2310
rect 59666 2310 59868 2327
rect 60424 2327 60440 2344
rect 60870 2344 61458 2360
rect 60870 2327 60886 2344
rect 60424 2310 60626 2327
rect 59666 2272 60626 2310
rect 60684 2310 60886 2327
rect 61442 2327 61458 2344
rect 61888 2344 62476 2360
rect 61888 2327 61904 2344
rect 61442 2310 61644 2327
rect 60684 2272 61644 2310
rect 61702 2310 61904 2327
rect 62460 2327 62476 2344
rect 62906 2344 63494 2360
rect 62906 2327 62922 2344
rect 62460 2310 62662 2327
rect 61702 2272 62662 2310
rect 62720 2310 62922 2327
rect 63478 2327 63494 2344
rect 63924 2344 64512 2360
rect 63924 2327 63940 2344
rect 63478 2310 63680 2327
rect 62720 2272 63680 2310
rect 63738 2310 63940 2327
rect 64496 2327 64512 2344
rect 64942 2344 65530 2360
rect 64942 2327 64958 2344
rect 64496 2310 64698 2327
rect 63738 2272 64698 2310
rect 64756 2310 64958 2327
rect 65514 2327 65530 2344
rect 65960 2344 66548 2360
rect 65960 2327 65976 2344
rect 65514 2310 65716 2327
rect 64756 2272 65716 2310
rect 65774 2310 65976 2327
rect 66532 2327 66548 2344
rect 66978 2344 67566 2360
rect 66978 2327 66994 2344
rect 66532 2310 66734 2327
rect 65774 2272 66734 2310
rect 66792 2310 66994 2327
rect 67550 2327 67566 2344
rect 67996 2344 68584 2360
rect 67996 2327 68012 2344
rect 67550 2310 67752 2327
rect 66792 2272 67752 2310
rect 67810 2310 68012 2327
rect 68568 2327 68584 2344
rect 69014 2344 69602 2360
rect 69014 2327 69030 2344
rect 68568 2310 68770 2327
rect 67810 2272 68770 2310
rect 68828 2310 69030 2327
rect 69586 2327 69602 2344
rect 70032 2344 70620 2360
rect 70032 2327 70048 2344
rect 69586 2310 69788 2327
rect 68828 2272 69788 2310
rect 69846 2310 70048 2327
rect 70604 2327 70620 2344
rect 71050 2344 71638 2360
rect 71050 2327 71066 2344
rect 70604 2310 70806 2327
rect 69846 2272 70806 2310
rect 70864 2310 71066 2327
rect 71622 2327 71638 2344
rect 72068 2344 72656 2360
rect 72068 2327 72084 2344
rect 71622 2310 71824 2327
rect 70864 2272 71824 2310
rect 71882 2310 72084 2327
rect 72640 2327 72656 2344
rect 73086 2344 73674 2360
rect 73086 2327 73102 2344
rect 72640 2310 72842 2327
rect 71882 2272 72842 2310
rect 72900 2310 73102 2327
rect 73658 2327 73674 2344
rect 74104 2344 74692 2360
rect 74104 2327 74120 2344
rect 73658 2310 73860 2327
rect 72900 2272 73860 2310
rect 73918 2310 74120 2327
rect 74676 2327 74692 2344
rect 74676 2310 74878 2327
rect 73918 2272 74878 2310
rect 41488 2134 42448 2172
rect 41488 2117 41690 2134
rect 41674 2100 41690 2117
rect 42246 2117 42448 2134
rect 42506 2134 43466 2172
rect 42506 2117 42708 2134
rect 42246 2100 42262 2117
rect 41674 2084 42262 2100
rect 42692 2100 42708 2117
rect 43264 2117 43466 2134
rect 43524 2134 44484 2172
rect 43524 2117 43726 2134
rect 43264 2100 43280 2117
rect 42692 2084 43280 2100
rect 43710 2100 43726 2117
rect 44282 2117 44484 2134
rect 44542 2134 45502 2172
rect 44542 2117 44744 2134
rect 44282 2100 44298 2117
rect 43710 2084 44298 2100
rect 44728 2100 44744 2117
rect 45300 2117 45502 2134
rect 45560 2134 46520 2172
rect 45560 2117 45762 2134
rect 45300 2100 45316 2117
rect 44728 2084 45316 2100
rect 45746 2100 45762 2117
rect 46318 2117 46520 2134
rect 46578 2134 47538 2172
rect 46578 2117 46780 2134
rect 46318 2100 46334 2117
rect 45746 2084 46334 2100
rect 46764 2100 46780 2117
rect 47336 2117 47538 2134
rect 47596 2134 48556 2172
rect 47596 2117 47798 2134
rect 47336 2100 47352 2117
rect 46764 2084 47352 2100
rect 47782 2100 47798 2117
rect 48354 2117 48556 2134
rect 48614 2134 49574 2172
rect 48614 2117 48816 2134
rect 48354 2100 48370 2117
rect 47782 2084 48370 2100
rect 48800 2100 48816 2117
rect 49372 2117 49574 2134
rect 49632 2134 50592 2172
rect 49632 2117 49834 2134
rect 49372 2100 49388 2117
rect 48800 2084 49388 2100
rect 49818 2100 49834 2117
rect 50390 2117 50592 2134
rect 50650 2134 51610 2172
rect 50650 2117 50852 2134
rect 50390 2100 50406 2117
rect 49818 2084 50406 2100
rect 50836 2100 50852 2117
rect 51408 2117 51610 2134
rect 51668 2134 52628 2172
rect 51668 2117 51870 2134
rect 51408 2100 51424 2117
rect 50836 2084 51424 2100
rect 51854 2100 51870 2117
rect 52426 2117 52628 2134
rect 52426 2100 52442 2117
rect 51854 2084 52442 2100
rect 54576 1634 55536 1672
rect 54576 1617 54778 1634
rect 54762 1600 54778 1617
rect 55334 1617 55536 1634
rect 55594 1634 56554 1672
rect 55594 1617 55796 1634
rect 55334 1600 55350 1617
rect 54762 1584 55350 1600
rect 55780 1600 55796 1617
rect 56352 1617 56554 1634
rect 56612 1634 57572 1672
rect 56612 1617 56814 1634
rect 56352 1600 56368 1617
rect 55780 1584 56368 1600
rect 56798 1600 56814 1617
rect 57370 1617 57572 1634
rect 57630 1634 58590 1672
rect 57630 1617 57832 1634
rect 57370 1600 57386 1617
rect 56798 1584 57386 1600
rect 57816 1600 57832 1617
rect 58388 1617 58590 1634
rect 58648 1634 59608 1672
rect 58648 1617 58850 1634
rect 58388 1600 58404 1617
rect 57816 1584 58404 1600
rect 58834 1600 58850 1617
rect 59406 1617 59608 1634
rect 59666 1634 60626 1672
rect 59666 1617 59868 1634
rect 59406 1600 59422 1617
rect 58834 1584 59422 1600
rect 59852 1600 59868 1617
rect 60424 1617 60626 1634
rect 60684 1634 61644 1672
rect 60684 1617 60886 1634
rect 60424 1600 60440 1617
rect 59852 1584 60440 1600
rect 60870 1600 60886 1617
rect 61442 1617 61644 1634
rect 61702 1634 62662 1672
rect 61702 1617 61904 1634
rect 61442 1600 61458 1617
rect 60870 1584 61458 1600
rect 61888 1600 61904 1617
rect 62460 1617 62662 1634
rect 62720 1634 63680 1672
rect 62720 1617 62922 1634
rect 62460 1600 62476 1617
rect 61888 1584 62476 1600
rect 62906 1600 62922 1617
rect 63478 1617 63680 1634
rect 63738 1634 64698 1672
rect 63738 1617 63940 1634
rect 63478 1600 63494 1617
rect 62906 1584 63494 1600
rect 63924 1600 63940 1617
rect 64496 1617 64698 1634
rect 64756 1634 65716 1672
rect 64756 1617 64958 1634
rect 64496 1600 64512 1617
rect 63924 1584 64512 1600
rect 64942 1600 64958 1617
rect 65514 1617 65716 1634
rect 65774 1634 66734 1672
rect 65774 1617 65976 1634
rect 65514 1600 65530 1617
rect 64942 1584 65530 1600
rect 65960 1600 65976 1617
rect 66532 1617 66734 1634
rect 66792 1634 67752 1672
rect 66792 1617 66994 1634
rect 66532 1600 66548 1617
rect 65960 1584 66548 1600
rect 66978 1600 66994 1617
rect 67550 1617 67752 1634
rect 67810 1634 68770 1672
rect 67810 1617 68012 1634
rect 67550 1600 67566 1617
rect 66978 1584 67566 1600
rect 67996 1600 68012 1617
rect 68568 1617 68770 1634
rect 68828 1634 69788 1672
rect 68828 1617 69030 1634
rect 68568 1600 68584 1617
rect 67996 1584 68584 1600
rect 69014 1600 69030 1617
rect 69586 1617 69788 1634
rect 69846 1634 70806 1672
rect 69846 1617 70048 1634
rect 69586 1600 69602 1617
rect 69014 1584 69602 1600
rect 70032 1600 70048 1617
rect 70604 1617 70806 1634
rect 70864 1634 71824 1672
rect 70864 1617 71066 1634
rect 70604 1600 70620 1617
rect 70032 1584 70620 1600
rect 71050 1600 71066 1617
rect 71622 1617 71824 1634
rect 71882 1634 72842 1672
rect 71882 1617 72084 1634
rect 71622 1600 71638 1617
rect 71050 1584 71638 1600
rect 72068 1600 72084 1617
rect 72640 1617 72842 1634
rect 72900 1634 73860 1672
rect 72900 1617 73102 1634
rect 72640 1600 72656 1617
rect 72068 1584 72656 1600
rect 73086 1600 73102 1617
rect 73658 1617 73860 1634
rect 73918 1634 74878 1672
rect 73918 1617 74120 1634
rect 73658 1600 73674 1617
rect 73086 1584 73674 1600
rect 74104 1600 74120 1617
rect 74676 1617 74878 1634
rect 74676 1600 74692 1617
rect 74104 1584 74692 1600
rect 42132 1302 42720 1318
rect 42132 1285 42148 1302
rect 41946 1268 42148 1285
rect 42704 1285 42720 1302
rect 43150 1302 43738 1318
rect 43150 1285 43166 1302
rect 42704 1268 42906 1285
rect 41946 1230 42906 1268
rect 42964 1268 43166 1285
rect 43722 1285 43738 1302
rect 44168 1302 44756 1318
rect 44168 1285 44184 1302
rect 43722 1268 43924 1285
rect 42964 1230 43924 1268
rect 43982 1268 44184 1285
rect 44740 1285 44756 1302
rect 45186 1302 45774 1318
rect 45186 1285 45202 1302
rect 44740 1268 44942 1285
rect 43982 1230 44942 1268
rect 45000 1268 45202 1285
rect 45758 1285 45774 1302
rect 46204 1302 46792 1318
rect 46204 1285 46220 1302
rect 45758 1268 45960 1285
rect 45000 1230 45960 1268
rect 46018 1268 46220 1285
rect 46776 1285 46792 1302
rect 47222 1302 47810 1318
rect 47222 1285 47238 1302
rect 46776 1268 46978 1285
rect 46018 1230 46978 1268
rect 47036 1268 47238 1285
rect 47794 1285 47810 1302
rect 48240 1302 48828 1318
rect 48240 1285 48256 1302
rect 47794 1268 47996 1285
rect 47036 1230 47996 1268
rect 48054 1268 48256 1285
rect 48812 1285 48828 1302
rect 49258 1302 49846 1318
rect 49258 1285 49274 1302
rect 48812 1268 49014 1285
rect 48054 1230 49014 1268
rect 49072 1268 49274 1285
rect 49830 1285 49846 1302
rect 50276 1302 50864 1318
rect 50276 1285 50292 1302
rect 49830 1268 50032 1285
rect 49072 1230 50032 1268
rect 50090 1268 50292 1285
rect 50848 1285 50864 1302
rect 51294 1302 51882 1318
rect 51294 1285 51310 1302
rect 50848 1268 51050 1285
rect 50090 1230 51050 1268
rect 51108 1268 51310 1285
rect 51866 1285 51882 1302
rect 51866 1268 52068 1285
rect 51108 1230 52068 1268
rect 54762 1112 55350 1128
rect 54762 1095 54778 1112
rect 54576 1078 54778 1095
rect 55334 1095 55350 1112
rect 55780 1112 56368 1128
rect 55780 1095 55796 1112
rect 55334 1078 55536 1095
rect 54576 1040 55536 1078
rect 55594 1078 55796 1095
rect 56352 1095 56368 1112
rect 56798 1112 57386 1128
rect 56798 1095 56814 1112
rect 56352 1078 56554 1095
rect 55594 1040 56554 1078
rect 56612 1078 56814 1095
rect 57370 1095 57386 1112
rect 57816 1112 58404 1128
rect 57816 1095 57832 1112
rect 57370 1078 57572 1095
rect 56612 1040 57572 1078
rect 57630 1078 57832 1095
rect 58388 1095 58404 1112
rect 58834 1112 59422 1128
rect 58834 1095 58850 1112
rect 58388 1078 58590 1095
rect 57630 1040 58590 1078
rect 58648 1078 58850 1095
rect 59406 1095 59422 1112
rect 59852 1112 60440 1128
rect 59852 1095 59868 1112
rect 59406 1078 59608 1095
rect 58648 1040 59608 1078
rect 59666 1078 59868 1095
rect 60424 1095 60440 1112
rect 60870 1112 61458 1128
rect 60870 1095 60886 1112
rect 60424 1078 60626 1095
rect 59666 1040 60626 1078
rect 60684 1078 60886 1095
rect 61442 1095 61458 1112
rect 61888 1112 62476 1128
rect 61888 1095 61904 1112
rect 61442 1078 61644 1095
rect 60684 1040 61644 1078
rect 61702 1078 61904 1095
rect 62460 1095 62476 1112
rect 62906 1112 63494 1128
rect 62906 1095 62922 1112
rect 62460 1078 62662 1095
rect 61702 1040 62662 1078
rect 62720 1078 62922 1095
rect 63478 1095 63494 1112
rect 63924 1112 64512 1128
rect 63924 1095 63940 1112
rect 63478 1078 63680 1095
rect 62720 1040 63680 1078
rect 63738 1078 63940 1095
rect 64496 1095 64512 1112
rect 64942 1112 65530 1128
rect 64942 1095 64958 1112
rect 64496 1078 64698 1095
rect 63738 1040 64698 1078
rect 64756 1078 64958 1095
rect 65514 1095 65530 1112
rect 65960 1112 66548 1128
rect 65960 1095 65976 1112
rect 65514 1078 65716 1095
rect 64756 1040 65716 1078
rect 65774 1078 65976 1095
rect 66532 1095 66548 1112
rect 66978 1112 67566 1128
rect 66978 1095 66994 1112
rect 66532 1078 66734 1095
rect 65774 1040 66734 1078
rect 66792 1078 66994 1095
rect 67550 1095 67566 1112
rect 67996 1112 68584 1128
rect 67996 1095 68012 1112
rect 67550 1078 67752 1095
rect 66792 1040 67752 1078
rect 67810 1078 68012 1095
rect 68568 1095 68584 1112
rect 69014 1112 69602 1128
rect 69014 1095 69030 1112
rect 68568 1078 68770 1095
rect 67810 1040 68770 1078
rect 68828 1078 69030 1095
rect 69586 1095 69602 1112
rect 70032 1112 70620 1128
rect 70032 1095 70048 1112
rect 69586 1078 69788 1095
rect 68828 1040 69788 1078
rect 69846 1078 70048 1095
rect 70604 1095 70620 1112
rect 71050 1112 71638 1128
rect 71050 1095 71066 1112
rect 70604 1078 70806 1095
rect 69846 1040 70806 1078
rect 70864 1078 71066 1095
rect 71622 1095 71638 1112
rect 72068 1112 72656 1128
rect 72068 1095 72084 1112
rect 71622 1078 71824 1095
rect 70864 1040 71824 1078
rect 71882 1078 72084 1095
rect 72640 1095 72656 1112
rect 73086 1112 73674 1128
rect 73086 1095 73102 1112
rect 72640 1078 72842 1095
rect 71882 1040 72842 1078
rect 72900 1078 73102 1095
rect 73658 1095 73674 1112
rect 74104 1112 74692 1128
rect 74104 1095 74120 1112
rect 73658 1078 73860 1095
rect 72900 1040 73860 1078
rect 73918 1078 74120 1095
rect 74676 1095 74692 1112
rect 74676 1078 74878 1095
rect 73918 1040 74878 1078
rect 41946 592 42906 630
rect 41946 575 42148 592
rect 42132 558 42148 575
rect 42704 575 42906 592
rect 42964 592 43924 630
rect 42964 575 43166 592
rect 42704 558 42720 575
rect 42132 542 42720 558
rect 43150 558 43166 575
rect 43722 575 43924 592
rect 43982 592 44942 630
rect 43982 575 44184 592
rect 43722 558 43738 575
rect 43150 542 43738 558
rect 44168 558 44184 575
rect 44740 575 44942 592
rect 45000 592 45960 630
rect 45000 575 45202 592
rect 44740 558 44756 575
rect 44168 542 44756 558
rect 45186 558 45202 575
rect 45758 575 45960 592
rect 46018 592 46978 630
rect 46018 575 46220 592
rect 45758 558 45774 575
rect 45186 542 45774 558
rect 46204 558 46220 575
rect 46776 575 46978 592
rect 47036 592 47996 630
rect 47036 575 47238 592
rect 46776 558 46792 575
rect 46204 542 46792 558
rect 47222 558 47238 575
rect 47794 575 47996 592
rect 48054 592 49014 630
rect 48054 575 48256 592
rect 47794 558 47810 575
rect 47222 542 47810 558
rect 48240 558 48256 575
rect 48812 575 49014 592
rect 49072 592 50032 630
rect 49072 575 49274 592
rect 48812 558 48828 575
rect 48240 542 48828 558
rect 49258 558 49274 575
rect 49830 575 50032 592
rect 50090 592 51050 630
rect 50090 575 50292 592
rect 49830 558 49846 575
rect 49258 542 49846 558
rect 50276 558 50292 575
rect 50848 575 51050 592
rect 51108 592 52068 630
rect 51108 575 51310 592
rect 50848 558 50864 575
rect 50276 542 50864 558
rect 51294 558 51310 575
rect 51866 575 52068 592
rect 51866 558 51882 575
rect 51294 542 51882 558
rect 54576 402 55536 440
rect 54576 385 54778 402
rect 54762 368 54778 385
rect 55334 385 55536 402
rect 55594 402 56554 440
rect 55594 385 55796 402
rect 55334 368 55350 385
rect 54762 352 55350 368
rect 55780 368 55796 385
rect 56352 385 56554 402
rect 56612 402 57572 440
rect 56612 385 56814 402
rect 56352 368 56368 385
rect 55780 352 56368 368
rect 56798 368 56814 385
rect 57370 385 57572 402
rect 57630 402 58590 440
rect 57630 385 57832 402
rect 57370 368 57386 385
rect 56798 352 57386 368
rect 57816 368 57832 385
rect 58388 385 58590 402
rect 58648 402 59608 440
rect 58648 385 58850 402
rect 58388 368 58404 385
rect 57816 352 58404 368
rect 58834 368 58850 385
rect 59406 385 59608 402
rect 59666 402 60626 440
rect 59666 385 59868 402
rect 59406 368 59422 385
rect 58834 352 59422 368
rect 59852 368 59868 385
rect 60424 385 60626 402
rect 60684 402 61644 440
rect 60684 385 60886 402
rect 60424 368 60440 385
rect 59852 352 60440 368
rect 60870 368 60886 385
rect 61442 385 61644 402
rect 61702 402 62662 440
rect 61702 385 61904 402
rect 61442 368 61458 385
rect 60870 352 61458 368
rect 61888 368 61904 385
rect 62460 385 62662 402
rect 62720 402 63680 440
rect 62720 385 62922 402
rect 62460 368 62476 385
rect 61888 352 62476 368
rect 62906 368 62922 385
rect 63478 385 63680 402
rect 63738 402 64698 440
rect 63738 385 63940 402
rect 63478 368 63494 385
rect 62906 352 63494 368
rect 63924 368 63940 385
rect 64496 385 64698 402
rect 64756 402 65716 440
rect 64756 385 64958 402
rect 64496 368 64512 385
rect 63924 352 64512 368
rect 64942 368 64958 385
rect 65514 385 65716 402
rect 65774 402 66734 440
rect 65774 385 65976 402
rect 65514 368 65530 385
rect 64942 352 65530 368
rect 65960 368 65976 385
rect 66532 385 66734 402
rect 66792 402 67752 440
rect 66792 385 66994 402
rect 66532 368 66548 385
rect 65960 352 66548 368
rect 66978 368 66994 385
rect 67550 385 67752 402
rect 67810 402 68770 440
rect 67810 385 68012 402
rect 67550 368 67566 385
rect 66978 352 67566 368
rect 67996 368 68012 385
rect 68568 385 68770 402
rect 68828 402 69788 440
rect 68828 385 69030 402
rect 68568 368 68584 385
rect 67996 352 68584 368
rect 69014 368 69030 385
rect 69586 385 69788 402
rect 69846 402 70806 440
rect 69846 385 70048 402
rect 69586 368 69602 385
rect 69014 352 69602 368
rect 70032 368 70048 385
rect 70604 385 70806 402
rect 70864 402 71824 440
rect 70864 385 71066 402
rect 70604 368 70620 385
rect 70032 352 70620 368
rect 71050 368 71066 385
rect 71622 385 71824 402
rect 71882 402 72842 440
rect 71882 385 72084 402
rect 71622 368 71638 385
rect 71050 352 71638 368
rect 72068 368 72084 385
rect 72640 385 72842 402
rect 72900 402 73860 440
rect 72900 385 73102 402
rect 72640 368 72656 385
rect 72068 352 72656 368
rect 73086 368 73102 385
rect 73658 385 73860 402
rect 73918 402 74878 440
rect 73918 385 74120 402
rect 73658 368 73674 385
rect 73086 352 73674 368
rect 74104 368 74120 385
rect 74676 385 74878 402
rect 74676 368 74692 385
rect 74104 352 74692 368
<< polycont >>
rect 17686 27891 18242 27925
rect 18704 27891 19260 27925
rect 19722 27891 20278 27925
rect 20740 27891 21296 27925
rect 21758 27891 22314 27925
rect 22776 27891 23332 27925
rect 23794 27891 24350 27925
rect 24812 27891 25368 27925
rect 25830 27891 26386 27925
rect 26848 27891 27404 27925
rect 27866 27891 28422 27925
rect 28884 27891 29440 27925
rect 29902 27891 30458 27925
rect 30920 27891 31476 27925
rect 31938 27891 32494 27925
rect 32956 27891 33512 27925
rect 17686 27163 18242 27197
rect 18704 27163 19260 27197
rect 19722 27163 20278 27197
rect 20740 27163 21296 27197
rect 21758 27163 22314 27197
rect 22776 27163 23332 27197
rect 23794 27163 24350 27197
rect 24812 27163 25368 27197
rect 25830 27163 26386 27197
rect 26848 27163 27404 27197
rect 27866 27163 28422 27197
rect 28884 27163 29440 27197
rect 29902 27163 30458 27197
rect 30920 27163 31476 27197
rect 31938 27163 32494 27197
rect 32956 27163 33512 27197
rect 17686 26755 18242 26789
rect 18704 26755 19260 26789
rect 19722 26755 20278 26789
rect 20740 26755 21296 26789
rect 21758 26755 22314 26789
rect 22776 26755 23332 26789
rect 23794 26755 24350 26789
rect 24812 26755 25368 26789
rect 25830 26755 26386 26789
rect 26848 26755 27404 26789
rect 27866 26755 28422 26789
rect 28884 26755 29440 26789
rect 29902 26755 30458 26789
rect 30920 26755 31476 26789
rect 31938 26755 32494 26789
rect 32956 26755 33512 26789
rect 17686 26027 18242 26061
rect 18704 26027 19260 26061
rect 19722 26027 20278 26061
rect 20740 26027 21296 26061
rect 21758 26027 22314 26061
rect 22776 26027 23332 26061
rect 23794 26027 24350 26061
rect 24812 26027 25368 26061
rect 25830 26027 26386 26061
rect 26848 26027 27404 26061
rect 27866 26027 28422 26061
rect 28884 26027 29440 26061
rect 29902 26027 30458 26061
rect 30920 26027 31476 26061
rect 31938 26027 32494 26061
rect 32956 26027 33512 26061
rect 17686 25619 18242 25653
rect 18704 25619 19260 25653
rect 19722 25619 20278 25653
rect 20740 25619 21296 25653
rect 21758 25619 22314 25653
rect 22776 25619 23332 25653
rect 23794 25619 24350 25653
rect 24812 25619 25368 25653
rect 25830 25619 26386 25653
rect 26848 25619 27404 25653
rect 27866 25619 28422 25653
rect 28884 25619 29440 25653
rect 29902 25619 30458 25653
rect 30920 25619 31476 25653
rect 31938 25619 32494 25653
rect 32956 25619 33512 25653
rect 17686 24891 18242 24925
rect 18704 24891 19260 24925
rect 19722 24891 20278 24925
rect 20740 24891 21296 24925
rect 21758 24891 22314 24925
rect 22776 24891 23332 24925
rect 23794 24891 24350 24925
rect 24812 24891 25368 24925
rect 25830 24891 26386 24925
rect 26848 24891 27404 24925
rect 27866 24891 28422 24925
rect 28884 24891 29440 24925
rect 29902 24891 30458 24925
rect 30920 24891 31476 24925
rect 31938 24891 32494 24925
rect 32956 24891 33512 24925
rect 18880 23981 19436 24015
rect 19898 23981 20454 24015
rect 20916 23981 21472 24015
rect 21934 23981 22490 24015
rect 22952 23981 23508 24015
rect 23970 23981 24526 24015
rect 24988 23981 25544 24015
rect 26006 23981 26562 24015
rect 27024 23981 27580 24015
rect 28042 23981 28598 24015
rect 29060 23981 29616 24015
rect 30078 23981 30634 24015
rect 31096 23981 31652 24015
rect 32114 23981 32670 24015
rect 18880 23253 19436 23287
rect 19898 23253 20454 23287
rect 20916 23253 21472 23287
rect 21934 23253 22490 23287
rect 22952 23253 23508 23287
rect 23970 23253 24526 23287
rect 24988 23253 25544 23287
rect 26006 23253 26562 23287
rect 27024 23253 27580 23287
rect 28042 23253 28598 23287
rect 29060 23253 29616 23287
rect 30078 23253 30634 23287
rect 31096 23253 31652 23287
rect 32114 23253 32670 23287
rect 18880 22949 19436 22983
rect 19898 22949 20454 22983
rect 20916 22949 21472 22983
rect 21934 22949 22490 22983
rect 22952 22949 23508 22983
rect 23970 22949 24526 22983
rect 24988 22949 25544 22983
rect 26006 22949 26562 22983
rect 27024 22949 27580 22983
rect 28042 22949 28598 22983
rect 29060 22949 29616 22983
rect 30078 22949 30634 22983
rect 31096 22949 31652 22983
rect 32114 22949 32670 22983
rect 18880 22221 19436 22255
rect 19898 22221 20454 22255
rect 20916 22221 21472 22255
rect 21934 22221 22490 22255
rect 22952 22221 23508 22255
rect 23970 22221 24526 22255
rect 24988 22221 25544 22255
rect 26006 22221 26562 22255
rect 27024 22221 27580 22255
rect 28042 22221 28598 22255
rect 29060 22221 29616 22255
rect 30078 22221 30634 22255
rect 31096 22221 31652 22255
rect 32114 22221 32670 22255
rect 18672 21345 19228 21379
rect 19690 21345 20246 21379
rect 20708 21345 21264 21379
rect 21726 21345 22282 21379
rect 22744 21345 23300 21379
rect 23762 21345 24318 21379
rect 24780 21345 25336 21379
rect 25798 21345 26354 21379
rect 26816 21345 27372 21379
rect 27834 21345 28390 21379
rect 28852 21345 29408 21379
rect 29870 21345 30426 21379
rect 30888 21345 31444 21379
rect 31906 21345 32462 21379
rect 32924 21345 33480 21379
rect 13368 21241 13924 21275
rect 14386 21241 14942 21275
rect 15404 21241 15960 21275
rect 16422 21241 16978 21275
rect 18672 20617 19228 20651
rect 19690 20617 20246 20651
rect 20708 20617 21264 20651
rect 21726 20617 22282 20651
rect 22744 20617 23300 20651
rect 23762 20617 24318 20651
rect 24780 20617 25336 20651
rect 25798 20617 26354 20651
rect 26816 20617 27372 20651
rect 27834 20617 28390 20651
rect 28852 20617 29408 20651
rect 29870 20617 30426 20651
rect 30888 20617 31444 20651
rect 31906 20617 32462 20651
rect 32924 20617 33480 20651
rect 13368 20513 13924 20547
rect 14386 20513 14942 20547
rect 15404 20513 15960 20547
rect 16422 20513 16978 20547
rect 13368 20209 13924 20243
rect 14386 20209 14942 20243
rect 15404 20209 15960 20243
rect 16422 20209 16978 20243
rect 18672 20089 19228 20123
rect 19690 20089 20246 20123
rect 20708 20089 21264 20123
rect 21726 20089 22282 20123
rect 22744 20089 23300 20123
rect 23762 20089 24318 20123
rect 24780 20089 25336 20123
rect 25798 20089 26354 20123
rect 26816 20089 27372 20123
rect 27834 20089 28390 20123
rect 28852 20089 29408 20123
rect 29870 20089 30426 20123
rect 30888 20089 31444 20123
rect 31906 20089 32462 20123
rect 32924 20089 33480 20123
rect 13368 19481 13924 19515
rect 14386 19481 14942 19515
rect 15404 19481 15960 19515
rect 16422 19481 16978 19515
rect 18672 19361 19228 19395
rect 19690 19361 20246 19395
rect 20708 19361 21264 19395
rect 21726 19361 22282 19395
rect 22744 19361 23300 19395
rect 23762 19361 24318 19395
rect 24780 19361 25336 19395
rect 25798 19361 26354 19395
rect 26816 19361 27372 19395
rect 27834 19361 28390 19395
rect 28852 19361 29408 19395
rect 29870 19361 30426 19395
rect 30888 19361 31444 19395
rect 31906 19361 32462 19395
rect 32924 19361 33480 19395
rect 13368 19177 13924 19211
rect 14386 19177 14942 19211
rect 15404 19177 15960 19211
rect 16422 19177 16978 19211
rect 18672 18833 19228 18867
rect 19690 18833 20246 18867
rect 20708 18833 21264 18867
rect 21726 18833 22282 18867
rect 22744 18833 23300 18867
rect 23762 18833 24318 18867
rect 24780 18833 25336 18867
rect 25798 18833 26354 18867
rect 26816 18833 27372 18867
rect 27834 18833 28390 18867
rect 28852 18833 29408 18867
rect 29870 18833 30426 18867
rect 30888 18833 31444 18867
rect 31906 18833 32462 18867
rect 32924 18833 33480 18867
rect 13368 18449 13924 18483
rect 14386 18449 14942 18483
rect 15404 18449 15960 18483
rect 16422 18449 16978 18483
rect 13368 18145 13924 18179
rect 14386 18145 14942 18179
rect 15404 18145 15960 18179
rect 16422 18145 16978 18179
rect 18672 18105 19228 18139
rect 19690 18105 20246 18139
rect 20708 18105 21264 18139
rect 21726 18105 22282 18139
rect 22744 18105 23300 18139
rect 23762 18105 24318 18139
rect 24780 18105 25336 18139
rect 25798 18105 26354 18139
rect 26816 18105 27372 18139
rect 27834 18105 28390 18139
rect 28852 18105 29408 18139
rect 29870 18105 30426 18139
rect 30888 18105 31444 18139
rect 31906 18105 32462 18139
rect 32924 18105 33480 18139
rect 18672 17577 19228 17611
rect 19690 17577 20246 17611
rect 20708 17577 21264 17611
rect 21726 17577 22282 17611
rect 22744 17577 23300 17611
rect 23762 17577 24318 17611
rect 24780 17577 25336 17611
rect 25798 17577 26354 17611
rect 26816 17577 27372 17611
rect 27834 17577 28390 17611
rect 28852 17577 29408 17611
rect 29870 17577 30426 17611
rect 30888 17577 31444 17611
rect 31906 17577 32462 17611
rect 32924 17577 33480 17611
rect 13368 17417 13924 17451
rect 14386 17417 14942 17451
rect 15404 17417 15960 17451
rect 16422 17417 16978 17451
rect 18672 16849 19228 16883
rect 19690 16849 20246 16883
rect 20708 16849 21264 16883
rect 21726 16849 22282 16883
rect 22744 16849 23300 16883
rect 23762 16849 24318 16883
rect 24780 16849 25336 16883
rect 25798 16849 26354 16883
rect 26816 16849 27372 16883
rect 27834 16849 28390 16883
rect 28852 16849 29408 16883
rect 29870 16849 30426 16883
rect 30888 16849 31444 16883
rect 31906 16849 32462 16883
rect 32924 16849 33480 16883
rect 58686 27891 59242 27925
rect 59704 27891 60260 27925
rect 60722 27891 61278 27925
rect 61740 27891 62296 27925
rect 62758 27891 63314 27925
rect 63776 27891 64332 27925
rect 64794 27891 65350 27925
rect 65812 27891 66368 27925
rect 66830 27891 67386 27925
rect 67848 27891 68404 27925
rect 68866 27891 69422 27925
rect 69884 27891 70440 27925
rect 70902 27891 71458 27925
rect 71920 27891 72476 27925
rect 72938 27891 73494 27925
rect 73956 27891 74512 27925
rect 58686 27163 59242 27197
rect 59704 27163 60260 27197
rect 60722 27163 61278 27197
rect 61740 27163 62296 27197
rect 62758 27163 63314 27197
rect 63776 27163 64332 27197
rect 64794 27163 65350 27197
rect 65812 27163 66368 27197
rect 66830 27163 67386 27197
rect 67848 27163 68404 27197
rect 68866 27163 69422 27197
rect 69884 27163 70440 27197
rect 70902 27163 71458 27197
rect 71920 27163 72476 27197
rect 72938 27163 73494 27197
rect 73956 27163 74512 27197
rect 58686 26755 59242 26789
rect 59704 26755 60260 26789
rect 60722 26755 61278 26789
rect 61740 26755 62296 26789
rect 62758 26755 63314 26789
rect 63776 26755 64332 26789
rect 64794 26755 65350 26789
rect 65812 26755 66368 26789
rect 66830 26755 67386 26789
rect 67848 26755 68404 26789
rect 68866 26755 69422 26789
rect 69884 26755 70440 26789
rect 70902 26755 71458 26789
rect 71920 26755 72476 26789
rect 72938 26755 73494 26789
rect 73956 26755 74512 26789
rect 58686 26027 59242 26061
rect 59704 26027 60260 26061
rect 60722 26027 61278 26061
rect 61740 26027 62296 26061
rect 62758 26027 63314 26061
rect 63776 26027 64332 26061
rect 64794 26027 65350 26061
rect 65812 26027 66368 26061
rect 66830 26027 67386 26061
rect 67848 26027 68404 26061
rect 68866 26027 69422 26061
rect 69884 26027 70440 26061
rect 70902 26027 71458 26061
rect 71920 26027 72476 26061
rect 72938 26027 73494 26061
rect 73956 26027 74512 26061
rect 58686 25619 59242 25653
rect 59704 25619 60260 25653
rect 60722 25619 61278 25653
rect 61740 25619 62296 25653
rect 62758 25619 63314 25653
rect 63776 25619 64332 25653
rect 64794 25619 65350 25653
rect 65812 25619 66368 25653
rect 66830 25619 67386 25653
rect 67848 25619 68404 25653
rect 68866 25619 69422 25653
rect 69884 25619 70440 25653
rect 70902 25619 71458 25653
rect 71920 25619 72476 25653
rect 72938 25619 73494 25653
rect 73956 25619 74512 25653
rect 58686 24891 59242 24925
rect 59704 24891 60260 24925
rect 60722 24891 61278 24925
rect 61740 24891 62296 24925
rect 62758 24891 63314 24925
rect 63776 24891 64332 24925
rect 64794 24891 65350 24925
rect 65812 24891 66368 24925
rect 66830 24891 67386 24925
rect 67848 24891 68404 24925
rect 68866 24891 69422 24925
rect 69884 24891 70440 24925
rect 70902 24891 71458 24925
rect 71920 24891 72476 24925
rect 72938 24891 73494 24925
rect 73956 24891 74512 24925
rect 59880 23981 60436 24015
rect 60898 23981 61454 24015
rect 61916 23981 62472 24015
rect 62934 23981 63490 24015
rect 63952 23981 64508 24015
rect 64970 23981 65526 24015
rect 65988 23981 66544 24015
rect 67006 23981 67562 24015
rect 68024 23981 68580 24015
rect 69042 23981 69598 24015
rect 70060 23981 70616 24015
rect 71078 23981 71634 24015
rect 72096 23981 72652 24015
rect 73114 23981 73670 24015
rect 59880 23253 60436 23287
rect 60898 23253 61454 23287
rect 61916 23253 62472 23287
rect 62934 23253 63490 23287
rect 63952 23253 64508 23287
rect 64970 23253 65526 23287
rect 65988 23253 66544 23287
rect 67006 23253 67562 23287
rect 68024 23253 68580 23287
rect 69042 23253 69598 23287
rect 70060 23253 70616 23287
rect 71078 23253 71634 23287
rect 72096 23253 72652 23287
rect 73114 23253 73670 23287
rect 59880 22949 60436 22983
rect 60898 22949 61454 22983
rect 61916 22949 62472 22983
rect 62934 22949 63490 22983
rect 63952 22949 64508 22983
rect 64970 22949 65526 22983
rect 65988 22949 66544 22983
rect 67006 22949 67562 22983
rect 68024 22949 68580 22983
rect 69042 22949 69598 22983
rect 70060 22949 70616 22983
rect 71078 22949 71634 22983
rect 72096 22949 72652 22983
rect 73114 22949 73670 22983
rect 59880 22221 60436 22255
rect 60898 22221 61454 22255
rect 61916 22221 62472 22255
rect 62934 22221 63490 22255
rect 63952 22221 64508 22255
rect 64970 22221 65526 22255
rect 65988 22221 66544 22255
rect 67006 22221 67562 22255
rect 68024 22221 68580 22255
rect 69042 22221 69598 22255
rect 70060 22221 70616 22255
rect 71078 22221 71634 22255
rect 72096 22221 72652 22255
rect 73114 22221 73670 22255
rect 59672 21345 60228 21379
rect 60690 21345 61246 21379
rect 61708 21345 62264 21379
rect 62726 21345 63282 21379
rect 63744 21345 64300 21379
rect 64762 21345 65318 21379
rect 65780 21345 66336 21379
rect 66798 21345 67354 21379
rect 67816 21345 68372 21379
rect 68834 21345 69390 21379
rect 69852 21345 70408 21379
rect 70870 21345 71426 21379
rect 71888 21345 72444 21379
rect 72906 21345 73462 21379
rect 73924 21345 74480 21379
rect 54368 21241 54924 21275
rect 55386 21241 55942 21275
rect 56404 21241 56960 21275
rect 57422 21241 57978 21275
rect 59672 20617 60228 20651
rect 60690 20617 61246 20651
rect 61708 20617 62264 20651
rect 62726 20617 63282 20651
rect 63744 20617 64300 20651
rect 64762 20617 65318 20651
rect 65780 20617 66336 20651
rect 66798 20617 67354 20651
rect 67816 20617 68372 20651
rect 68834 20617 69390 20651
rect 69852 20617 70408 20651
rect 70870 20617 71426 20651
rect 71888 20617 72444 20651
rect 72906 20617 73462 20651
rect 73924 20617 74480 20651
rect 54368 20513 54924 20547
rect 55386 20513 55942 20547
rect 56404 20513 56960 20547
rect 57422 20513 57978 20547
rect 54368 20209 54924 20243
rect 55386 20209 55942 20243
rect 56404 20209 56960 20243
rect 57422 20209 57978 20243
rect 59672 20089 60228 20123
rect 60690 20089 61246 20123
rect 61708 20089 62264 20123
rect 62726 20089 63282 20123
rect 63744 20089 64300 20123
rect 64762 20089 65318 20123
rect 65780 20089 66336 20123
rect 66798 20089 67354 20123
rect 67816 20089 68372 20123
rect 68834 20089 69390 20123
rect 69852 20089 70408 20123
rect 70870 20089 71426 20123
rect 71888 20089 72444 20123
rect 72906 20089 73462 20123
rect 73924 20089 74480 20123
rect 54368 19481 54924 19515
rect 55386 19481 55942 19515
rect 56404 19481 56960 19515
rect 57422 19481 57978 19515
rect 59672 19361 60228 19395
rect 60690 19361 61246 19395
rect 61708 19361 62264 19395
rect 62726 19361 63282 19395
rect 63744 19361 64300 19395
rect 64762 19361 65318 19395
rect 65780 19361 66336 19395
rect 66798 19361 67354 19395
rect 67816 19361 68372 19395
rect 68834 19361 69390 19395
rect 69852 19361 70408 19395
rect 70870 19361 71426 19395
rect 71888 19361 72444 19395
rect 72906 19361 73462 19395
rect 73924 19361 74480 19395
rect 54368 19177 54924 19211
rect 55386 19177 55942 19211
rect 56404 19177 56960 19211
rect 57422 19177 57978 19211
rect 59672 18833 60228 18867
rect 60690 18833 61246 18867
rect 61708 18833 62264 18867
rect 62726 18833 63282 18867
rect 63744 18833 64300 18867
rect 64762 18833 65318 18867
rect 65780 18833 66336 18867
rect 66798 18833 67354 18867
rect 67816 18833 68372 18867
rect 68834 18833 69390 18867
rect 69852 18833 70408 18867
rect 70870 18833 71426 18867
rect 71888 18833 72444 18867
rect 72906 18833 73462 18867
rect 73924 18833 74480 18867
rect 54368 18449 54924 18483
rect 55386 18449 55942 18483
rect 56404 18449 56960 18483
rect 57422 18449 57978 18483
rect 54368 18145 54924 18179
rect 55386 18145 55942 18179
rect 56404 18145 56960 18179
rect 57422 18145 57978 18179
rect 59672 18105 60228 18139
rect 60690 18105 61246 18139
rect 61708 18105 62264 18139
rect 62726 18105 63282 18139
rect 63744 18105 64300 18139
rect 64762 18105 65318 18139
rect 65780 18105 66336 18139
rect 66798 18105 67354 18139
rect 67816 18105 68372 18139
rect 68834 18105 69390 18139
rect 69852 18105 70408 18139
rect 70870 18105 71426 18139
rect 71888 18105 72444 18139
rect 72906 18105 73462 18139
rect 73924 18105 74480 18139
rect 59672 17577 60228 17611
rect 60690 17577 61246 17611
rect 61708 17577 62264 17611
rect 62726 17577 63282 17611
rect 63744 17577 64300 17611
rect 64762 17577 65318 17611
rect 65780 17577 66336 17611
rect 66798 17577 67354 17611
rect 67816 17577 68372 17611
rect 68834 17577 69390 17611
rect 69852 17577 70408 17611
rect 70870 17577 71426 17611
rect 71888 17577 72444 17611
rect 72906 17577 73462 17611
rect 73924 17577 74480 17611
rect 54368 17417 54924 17451
rect 55386 17417 55942 17451
rect 56404 17417 56960 17451
rect 57422 17417 57978 17451
rect 59672 16849 60228 16883
rect 60690 16849 61246 16883
rect 61708 16849 62264 16883
rect 62726 16849 63282 16883
rect 63744 16849 64300 16883
rect 64762 16849 65318 16883
rect 65780 16849 66336 16883
rect 66798 16849 67354 16883
rect 67816 16849 68372 16883
rect 68834 16849 69390 16883
rect 69852 16849 70408 16883
rect 70870 16849 71426 16883
rect 71888 16849 72444 16883
rect 72906 16849 73462 16883
rect 73924 16849 74480 16883
rect 13780 14372 14336 14406
rect 14798 14372 15354 14406
rect 15816 14372 16372 14406
rect 16834 14372 17390 14406
rect 17852 14372 18408 14406
rect 18870 14372 19426 14406
rect 19888 14372 20444 14406
rect 20906 14372 21462 14406
rect 21924 14372 22480 14406
rect 22942 14372 23498 14406
rect 23960 14372 24516 14406
rect 24978 14372 25534 14406
rect 25996 14372 26552 14406
rect 27014 14372 27570 14406
rect 28032 14372 28588 14406
rect 29050 14372 29606 14406
rect 30068 14372 30624 14406
rect 31086 14372 31642 14406
rect 32104 14372 32660 14406
rect 33122 14372 33678 14406
rect 2014 13896 2570 13930
rect 3032 13896 3588 13930
rect 4050 13896 4606 13930
rect 5068 13896 5624 13930
rect 6086 13896 6642 13930
rect 7104 13896 7660 13930
rect 8122 13896 8678 13930
rect 9140 13896 9696 13930
rect 10158 13896 10714 13930
rect 13780 13662 14336 13696
rect 14798 13662 15354 13696
rect 15816 13662 16372 13696
rect 16834 13662 17390 13696
rect 17852 13662 18408 13696
rect 18870 13662 19426 13696
rect 19888 13662 20444 13696
rect 20906 13662 21462 13696
rect 21924 13662 22480 13696
rect 22942 13662 23498 13696
rect 23960 13662 24516 13696
rect 24978 13662 25534 13696
rect 25996 13662 26552 13696
rect 27014 13662 27570 13696
rect 28032 13662 28588 13696
rect 29050 13662 29606 13696
rect 30068 13662 30624 13696
rect 31086 13662 31642 13696
rect 32104 13662 32660 13696
rect 33122 13662 33678 13696
rect 13780 13554 14336 13588
rect 14798 13554 15354 13588
rect 15816 13554 16372 13588
rect 16834 13554 17390 13588
rect 17852 13554 18408 13588
rect 18870 13554 19426 13588
rect 19888 13554 20444 13588
rect 20906 13554 21462 13588
rect 21924 13554 22480 13588
rect 22942 13554 23498 13588
rect 23960 13554 24516 13588
rect 24978 13554 25534 13588
rect 25996 13554 26552 13588
rect 27014 13554 27570 13588
rect 28032 13554 28588 13588
rect 29050 13554 29606 13588
rect 30068 13554 30624 13588
rect 31086 13554 31642 13588
rect 32104 13554 32660 13588
rect 33122 13554 33678 13588
rect 2014 13186 2570 13220
rect 3032 13186 3588 13220
rect 2014 13078 2570 13112
rect 4050 13186 4606 13220
rect 3032 13078 3588 13112
rect 5068 13186 5624 13220
rect 4050 13078 4606 13112
rect 6086 13186 6642 13220
rect 5068 13078 5624 13112
rect 7104 13186 7660 13220
rect 6086 13078 6642 13112
rect 8122 13186 8678 13220
rect 7104 13078 7660 13112
rect 9140 13186 9696 13220
rect 8122 13078 8678 13112
rect 10158 13186 10714 13220
rect 9140 13078 9696 13112
rect 10158 13078 10714 13112
rect 13780 12844 14336 12878
rect 14798 12844 15354 12878
rect 15816 12844 16372 12878
rect 16834 12844 17390 12878
rect 17852 12844 18408 12878
rect 18870 12844 19426 12878
rect 19888 12844 20444 12878
rect 20906 12844 21462 12878
rect 21924 12844 22480 12878
rect 22942 12844 23498 12878
rect 23960 12844 24516 12878
rect 24978 12844 25534 12878
rect 25996 12844 26552 12878
rect 27014 12844 27570 12878
rect 28032 12844 28588 12878
rect 29050 12844 29606 12878
rect 30068 12844 30624 12878
rect 31086 12844 31642 12878
rect 32104 12844 32660 12878
rect 33122 12844 33678 12878
rect 2014 12368 2570 12402
rect 3032 12368 3588 12402
rect 2014 12260 2570 12294
rect 4050 12368 4606 12402
rect 3032 12260 3588 12294
rect 5068 12368 5624 12402
rect 4050 12260 4606 12294
rect 6086 12368 6642 12402
rect 5068 12260 5624 12294
rect 7104 12368 7660 12402
rect 6086 12260 6642 12294
rect 8122 12368 8678 12402
rect 7104 12260 7660 12294
rect 9140 12368 9696 12402
rect 8122 12260 8678 12294
rect 10158 12368 10714 12402
rect 9140 12260 9696 12294
rect 10158 12260 10714 12294
rect 13780 12176 14336 12210
rect 14798 12176 15354 12210
rect 15816 12176 16372 12210
rect 16834 12176 17390 12210
rect 17852 12176 18408 12210
rect 18870 12176 19426 12210
rect 19888 12176 20444 12210
rect 20906 12176 21462 12210
rect 21924 12176 22480 12210
rect 22942 12176 23498 12210
rect 23960 12176 24516 12210
rect 24978 12176 25534 12210
rect 25996 12176 26552 12210
rect 27014 12176 27570 12210
rect 28032 12176 28588 12210
rect 29050 12176 29606 12210
rect 30068 12176 30624 12210
rect 31086 12176 31642 12210
rect 32104 12176 32660 12210
rect 33122 12176 33678 12210
rect 2014 11550 2570 11584
rect 3032 11550 3588 11584
rect 2014 11442 2570 11476
rect 4050 11550 4606 11584
rect 3032 11442 3588 11476
rect 5068 11550 5624 11584
rect 4050 11442 4606 11476
rect 6086 11550 6642 11584
rect 5068 11442 5624 11476
rect 7104 11550 7660 11584
rect 6086 11442 6642 11476
rect 8122 11550 8678 11584
rect 7104 11442 7660 11476
rect 9140 11550 9696 11584
rect 8122 11442 8678 11476
rect 10158 11550 10714 11584
rect 9140 11442 9696 11476
rect 10158 11442 10714 11476
rect 13780 11466 14336 11500
rect 14798 11466 15354 11500
rect 15816 11466 16372 11500
rect 16834 11466 17390 11500
rect 17852 11466 18408 11500
rect 18870 11466 19426 11500
rect 19888 11466 20444 11500
rect 20906 11466 21462 11500
rect 21924 11466 22480 11500
rect 22942 11466 23498 11500
rect 23960 11466 24516 11500
rect 24978 11466 25534 11500
rect 25996 11466 26552 11500
rect 27014 11466 27570 11500
rect 28032 11466 28588 11500
rect 29050 11466 29606 11500
rect 30068 11466 30624 11500
rect 31086 11466 31642 11500
rect 32104 11466 32660 11500
rect 33122 11466 33678 11500
rect 13780 10944 14336 10978
rect 14798 10944 15354 10978
rect 15816 10944 16372 10978
rect 16834 10944 17390 10978
rect 17852 10944 18408 10978
rect 18870 10944 19426 10978
rect 19888 10944 20444 10978
rect 20906 10944 21462 10978
rect 21924 10944 22480 10978
rect 22942 10944 23498 10978
rect 23960 10944 24516 10978
rect 24978 10944 25534 10978
rect 25996 10944 26552 10978
rect 27014 10944 27570 10978
rect 28032 10944 28588 10978
rect 29050 10944 29606 10978
rect 30068 10944 30624 10978
rect 31086 10944 31642 10978
rect 32104 10944 32660 10978
rect 33122 10944 33678 10978
rect 2014 10732 2570 10766
rect 3032 10732 3588 10766
rect 2014 10624 2570 10658
rect 4050 10732 4606 10766
rect 3032 10624 3588 10658
rect 5068 10732 5624 10766
rect 4050 10624 4606 10658
rect 6086 10732 6642 10766
rect 5068 10624 5624 10658
rect 7104 10732 7660 10766
rect 6086 10624 6642 10658
rect 8122 10732 8678 10766
rect 7104 10624 7660 10658
rect 9140 10732 9696 10766
rect 8122 10624 8678 10658
rect 10158 10732 10714 10766
rect 9140 10624 9696 10658
rect 10158 10624 10714 10658
rect 13780 10234 14336 10268
rect 14798 10234 15354 10268
rect 15816 10234 16372 10268
rect 16834 10234 17390 10268
rect 17852 10234 18408 10268
rect 18870 10234 19426 10268
rect 19888 10234 20444 10268
rect 20906 10234 21462 10268
rect 21924 10234 22480 10268
rect 22942 10234 23498 10268
rect 23960 10234 24516 10268
rect 24978 10234 25534 10268
rect 25996 10234 26552 10268
rect 27014 10234 27570 10268
rect 28032 10234 28588 10268
rect 29050 10234 29606 10268
rect 30068 10234 30624 10268
rect 31086 10234 31642 10268
rect 32104 10234 32660 10268
rect 33122 10234 33678 10268
rect 2014 9914 2570 9948
rect 3032 9914 3588 9948
rect 2014 9806 2570 9840
rect 4050 9914 4606 9948
rect 3032 9806 3588 9840
rect 5068 9914 5624 9948
rect 4050 9806 4606 9840
rect 6086 9914 6642 9948
rect 5068 9806 5624 9840
rect 7104 9914 7660 9948
rect 6086 9806 6642 9840
rect 8122 9914 8678 9948
rect 7104 9806 7660 9840
rect 9140 9914 9696 9948
rect 8122 9806 8678 9840
rect 10158 9914 10714 9948
rect 9140 9806 9696 9840
rect 10158 9806 10714 9840
rect 13778 9710 14334 9744
rect 14796 9710 15352 9744
rect 15814 9710 16370 9744
rect 16832 9710 17388 9744
rect 17850 9710 18406 9744
rect 18868 9710 19424 9744
rect 19886 9710 20442 9744
rect 20904 9710 21460 9744
rect 21922 9710 22478 9744
rect 22940 9710 23496 9744
rect 23958 9710 24514 9744
rect 24976 9710 25532 9744
rect 25994 9710 26550 9744
rect 27012 9710 27568 9744
rect 28030 9710 28586 9744
rect 29048 9710 29604 9744
rect 30066 9710 30622 9744
rect 31084 9710 31640 9744
rect 32102 9710 32658 9744
rect 33120 9710 33676 9744
rect 2014 9096 2570 9130
rect 3032 9096 3588 9130
rect 2014 8988 2570 9022
rect 4050 9096 4606 9130
rect 3032 8988 3588 9022
rect 5068 9096 5624 9130
rect 4050 8988 4606 9022
rect 6086 9096 6642 9130
rect 5068 8988 5624 9022
rect 7104 9096 7660 9130
rect 6086 8988 6642 9022
rect 8122 9096 8678 9130
rect 7104 8988 7660 9022
rect 9140 9096 9696 9130
rect 8122 8988 8678 9022
rect 10158 9096 10714 9130
rect 9140 8988 9696 9022
rect 10158 8988 10714 9022
rect 13778 9000 14334 9034
rect 14796 9000 15352 9034
rect 15814 9000 16370 9034
rect 16832 9000 17388 9034
rect 17850 9000 18406 9034
rect 18868 9000 19424 9034
rect 19886 9000 20442 9034
rect 20904 9000 21460 9034
rect 21922 9000 22478 9034
rect 22940 9000 23496 9034
rect 23958 9000 24514 9034
rect 24976 9000 25532 9034
rect 25994 9000 26550 9034
rect 27012 9000 27568 9034
rect 28030 9000 28586 9034
rect 29048 9000 29604 9034
rect 30066 9000 30622 9034
rect 31084 9000 31640 9034
rect 32102 9000 32658 9034
rect 33120 9000 33676 9034
rect 13778 8476 14334 8510
rect 14796 8476 15352 8510
rect 15814 8476 16370 8510
rect 16832 8476 17388 8510
rect 17850 8476 18406 8510
rect 18868 8476 19424 8510
rect 19886 8476 20442 8510
rect 20904 8476 21460 8510
rect 21922 8476 22478 8510
rect 22940 8476 23496 8510
rect 23958 8476 24514 8510
rect 24976 8476 25532 8510
rect 25994 8476 26550 8510
rect 27012 8476 27568 8510
rect 28030 8476 28586 8510
rect 29048 8476 29604 8510
rect 30066 8476 30622 8510
rect 31084 8476 31640 8510
rect 32102 8476 32658 8510
rect 33120 8476 33676 8510
rect 2014 8278 2570 8312
rect 3032 8278 3588 8312
rect 2014 8170 2570 8204
rect 4050 8278 4606 8312
rect 3032 8170 3588 8204
rect 5068 8278 5624 8312
rect 4050 8170 4606 8204
rect 6086 8278 6642 8312
rect 5068 8170 5624 8204
rect 7104 8278 7660 8312
rect 6086 8170 6642 8204
rect 8122 8278 8678 8312
rect 7104 8170 7660 8204
rect 9140 8278 9696 8312
rect 8122 8170 8678 8204
rect 10158 8278 10714 8312
rect 9140 8170 9696 8204
rect 10158 8170 10714 8204
rect 13778 7766 14334 7800
rect 14796 7766 15352 7800
rect 15814 7766 16370 7800
rect 16832 7766 17388 7800
rect 17850 7766 18406 7800
rect 18868 7766 19424 7800
rect 19886 7766 20442 7800
rect 20904 7766 21460 7800
rect 21922 7766 22478 7800
rect 22940 7766 23496 7800
rect 23958 7766 24514 7800
rect 24976 7766 25532 7800
rect 25994 7766 26550 7800
rect 27012 7766 27568 7800
rect 28030 7766 28586 7800
rect 29048 7766 29604 7800
rect 30066 7766 30622 7800
rect 31084 7766 31640 7800
rect 32102 7766 32658 7800
rect 33120 7766 33676 7800
rect 2014 7460 2570 7494
rect 3032 7460 3588 7494
rect 4050 7460 4606 7494
rect 5068 7460 5624 7494
rect 6086 7460 6642 7494
rect 7104 7460 7660 7494
rect 8122 7460 8678 7494
rect 9140 7460 9696 7494
rect 10158 7460 10714 7494
rect 13778 7244 14334 7278
rect 14796 7244 15352 7278
rect 15814 7244 16370 7278
rect 16832 7244 17388 7278
rect 17850 7244 18406 7278
rect 18868 7244 19424 7278
rect 19886 7244 20442 7278
rect 20904 7244 21460 7278
rect 21922 7244 22478 7278
rect 22940 7244 23496 7278
rect 23958 7244 24514 7278
rect 24976 7244 25532 7278
rect 25994 7244 26550 7278
rect 27012 7244 27568 7278
rect 28030 7244 28586 7278
rect 29048 7244 29604 7278
rect 30066 7244 30622 7278
rect 31084 7244 31640 7278
rect 32102 7244 32658 7278
rect 33120 7244 33676 7278
rect 13778 6534 14334 6568
rect 14796 6534 15352 6568
rect 15814 6534 16370 6568
rect 16832 6534 17388 6568
rect 17850 6534 18406 6568
rect 18868 6534 19424 6568
rect 19886 6534 20442 6568
rect 20904 6534 21460 6568
rect 21922 6534 22478 6568
rect 22940 6534 23496 6568
rect 23958 6534 24514 6568
rect 24976 6534 25532 6568
rect 25994 6534 26550 6568
rect 27012 6534 27568 6568
rect 28030 6534 28586 6568
rect 29048 6534 29604 6568
rect 30066 6534 30622 6568
rect 31084 6534 31640 6568
rect 32102 6534 32658 6568
rect 33120 6534 33676 6568
rect 690 6146 1246 6180
rect 1708 6146 2264 6180
rect 2726 6146 3282 6180
rect 3744 6146 4300 6180
rect 4762 6146 5318 6180
rect 5780 6146 6336 6180
rect 6798 6146 7354 6180
rect 7816 6146 8372 6180
rect 8834 6146 9390 6180
rect 9852 6146 10408 6180
rect 10870 6146 11426 6180
rect 13778 6010 14334 6044
rect 14796 6010 15352 6044
rect 15814 6010 16370 6044
rect 16832 6010 17388 6044
rect 17850 6010 18406 6044
rect 18868 6010 19424 6044
rect 19886 6010 20442 6044
rect 20904 6010 21460 6044
rect 21922 6010 22478 6044
rect 22940 6010 23496 6044
rect 23958 6010 24514 6044
rect 24976 6010 25532 6044
rect 25994 6010 26550 6044
rect 27012 6010 27568 6044
rect 28030 6010 28586 6044
rect 29048 6010 29604 6044
rect 30066 6010 30622 6044
rect 31084 6010 31640 6044
rect 32102 6010 32658 6044
rect 33120 6010 33676 6044
rect 690 5436 1246 5470
rect 1708 5436 2264 5470
rect 2726 5436 3282 5470
rect 3744 5436 4300 5470
rect 4762 5436 5318 5470
rect 5780 5436 6336 5470
rect 6798 5436 7354 5470
rect 7816 5436 8372 5470
rect 8834 5436 9390 5470
rect 9852 5436 10408 5470
rect 10870 5436 11426 5470
rect 13778 5300 14334 5334
rect 14796 5300 15352 5334
rect 15814 5300 16370 5334
rect 16832 5300 17388 5334
rect 17850 5300 18406 5334
rect 18868 5300 19424 5334
rect 19886 5300 20442 5334
rect 20904 5300 21460 5334
rect 21922 5300 22478 5334
rect 22940 5300 23496 5334
rect 23958 5300 24514 5334
rect 24976 5300 25532 5334
rect 25994 5300 26550 5334
rect 27012 5300 27568 5334
rect 28030 5300 28586 5334
rect 29048 5300 29604 5334
rect 30066 5300 30622 5334
rect 31084 5300 31640 5334
rect 32102 5300 32658 5334
rect 33120 5300 33676 5334
rect 690 5034 1246 5068
rect 1708 5034 2264 5068
rect 2726 5034 3282 5068
rect 3744 5034 4300 5068
rect 4762 5034 5318 5068
rect 5780 5034 6336 5068
rect 6798 5034 7354 5068
rect 7816 5034 8372 5068
rect 8834 5034 9390 5068
rect 9852 5034 10408 5068
rect 10870 5034 11426 5068
rect 13778 4776 14334 4810
rect 14796 4776 15352 4810
rect 15814 4776 16370 4810
rect 16832 4776 17388 4810
rect 17850 4776 18406 4810
rect 18868 4776 19424 4810
rect 19886 4776 20442 4810
rect 20904 4776 21460 4810
rect 21922 4776 22478 4810
rect 22940 4776 23496 4810
rect 23958 4776 24514 4810
rect 24976 4776 25532 4810
rect 25994 4776 26550 4810
rect 27012 4776 27568 4810
rect 28030 4776 28586 4810
rect 29048 4776 29604 4810
rect 30066 4776 30622 4810
rect 31084 4776 31640 4810
rect 32102 4776 32658 4810
rect 33120 4776 33676 4810
rect 690 4324 1246 4358
rect 1708 4324 2264 4358
rect 2726 4324 3282 4358
rect 3744 4324 4300 4358
rect 4762 4324 5318 4358
rect 5780 4324 6336 4358
rect 6798 4324 7354 4358
rect 7816 4324 8372 4358
rect 8834 4324 9390 4358
rect 9852 4324 10408 4358
rect 10870 4324 11426 4358
rect 13778 4066 14334 4100
rect 14796 4066 15352 4100
rect 15814 4066 16370 4100
rect 16832 4066 17388 4100
rect 17850 4066 18406 4100
rect 18868 4066 19424 4100
rect 19886 4066 20442 4100
rect 20904 4066 21460 4100
rect 21922 4066 22478 4100
rect 22940 4066 23496 4100
rect 23958 4066 24514 4100
rect 24976 4066 25532 4100
rect 25994 4066 26550 4100
rect 27012 4066 27568 4100
rect 28030 4066 28586 4100
rect 29048 4066 29604 4100
rect 30066 4066 30622 4100
rect 31084 4066 31640 4100
rect 32102 4066 32658 4100
rect 33120 4066 33676 4100
rect 690 3922 1246 3956
rect 1708 3922 2264 3956
rect 2726 3922 3282 3956
rect 3744 3922 4300 3956
rect 4762 3922 5318 3956
rect 5780 3922 6336 3956
rect 6798 3922 7354 3956
rect 7816 3922 8372 3956
rect 8834 3922 9390 3956
rect 9852 3922 10408 3956
rect 10870 3922 11426 3956
rect 13778 3544 14334 3578
rect 14796 3544 15352 3578
rect 15814 3544 16370 3578
rect 16832 3544 17388 3578
rect 17850 3544 18406 3578
rect 18868 3544 19424 3578
rect 19886 3544 20442 3578
rect 20904 3544 21460 3578
rect 21922 3544 22478 3578
rect 22940 3544 23496 3578
rect 23958 3544 24514 3578
rect 24976 3544 25532 3578
rect 25994 3544 26550 3578
rect 27012 3544 27568 3578
rect 28030 3544 28586 3578
rect 29048 3544 29604 3578
rect 30066 3544 30622 3578
rect 31084 3544 31640 3578
rect 32102 3544 32658 3578
rect 33120 3544 33676 3578
rect 690 3212 1246 3246
rect 1708 3212 2264 3246
rect 2726 3212 3282 3246
rect 3744 3212 4300 3246
rect 4762 3212 5318 3246
rect 5780 3212 6336 3246
rect 6798 3212 7354 3246
rect 7816 3212 8372 3246
rect 8834 3212 9390 3246
rect 9852 3212 10408 3246
rect 10870 3212 11426 3246
rect 690 2810 1246 2844
rect 1708 2810 2264 2844
rect 2726 2810 3282 2844
rect 3744 2810 4300 2844
rect 4762 2810 5318 2844
rect 5780 2810 6336 2844
rect 6798 2810 7354 2844
rect 7816 2810 8372 2844
rect 8834 2810 9390 2844
rect 9852 2810 10408 2844
rect 10870 2810 11426 2844
rect 13778 2834 14334 2868
rect 14796 2834 15352 2868
rect 15814 2834 16370 2868
rect 16832 2834 17388 2868
rect 17850 2834 18406 2868
rect 18868 2834 19424 2868
rect 19886 2834 20442 2868
rect 20904 2834 21460 2868
rect 21922 2834 22478 2868
rect 22940 2834 23496 2868
rect 23958 2834 24514 2868
rect 24976 2834 25532 2868
rect 25994 2834 26550 2868
rect 27012 2834 27568 2868
rect 28030 2834 28586 2868
rect 29048 2834 29604 2868
rect 30066 2834 30622 2868
rect 31084 2834 31640 2868
rect 32102 2834 32658 2868
rect 33120 2834 33676 2868
rect 13778 2310 14334 2344
rect 14796 2310 15352 2344
rect 15814 2310 16370 2344
rect 16832 2310 17388 2344
rect 17850 2310 18406 2344
rect 18868 2310 19424 2344
rect 19886 2310 20442 2344
rect 20904 2310 21460 2344
rect 21922 2310 22478 2344
rect 22940 2310 23496 2344
rect 23958 2310 24514 2344
rect 24976 2310 25532 2344
rect 25994 2310 26550 2344
rect 27012 2310 27568 2344
rect 28030 2310 28586 2344
rect 29048 2310 29604 2344
rect 30066 2310 30622 2344
rect 31084 2310 31640 2344
rect 32102 2310 32658 2344
rect 33120 2310 33676 2344
rect 690 2100 1246 2134
rect 1708 2100 2264 2134
rect 2726 2100 3282 2134
rect 3744 2100 4300 2134
rect 4762 2100 5318 2134
rect 5780 2100 6336 2134
rect 6798 2100 7354 2134
rect 7816 2100 8372 2134
rect 8834 2100 9390 2134
rect 9852 2100 10408 2134
rect 10870 2100 11426 2134
rect 13778 1600 14334 1634
rect 14796 1600 15352 1634
rect 15814 1600 16370 1634
rect 16832 1600 17388 1634
rect 17850 1600 18406 1634
rect 18868 1600 19424 1634
rect 19886 1600 20442 1634
rect 20904 1600 21460 1634
rect 21922 1600 22478 1634
rect 22940 1600 23496 1634
rect 23958 1600 24514 1634
rect 24976 1600 25532 1634
rect 25994 1600 26550 1634
rect 27012 1600 27568 1634
rect 28030 1600 28586 1634
rect 29048 1600 29604 1634
rect 30066 1600 30622 1634
rect 31084 1600 31640 1634
rect 32102 1600 32658 1634
rect 33120 1600 33676 1634
rect 1148 1268 1704 1302
rect 2166 1268 2722 1302
rect 3184 1268 3740 1302
rect 4202 1268 4758 1302
rect 5220 1268 5776 1302
rect 6238 1268 6794 1302
rect 7256 1268 7812 1302
rect 8274 1268 8830 1302
rect 9292 1268 9848 1302
rect 10310 1268 10866 1302
rect 13778 1078 14334 1112
rect 14796 1078 15352 1112
rect 15814 1078 16370 1112
rect 16832 1078 17388 1112
rect 17850 1078 18406 1112
rect 18868 1078 19424 1112
rect 19886 1078 20442 1112
rect 20904 1078 21460 1112
rect 21922 1078 22478 1112
rect 22940 1078 23496 1112
rect 23958 1078 24514 1112
rect 24976 1078 25532 1112
rect 25994 1078 26550 1112
rect 27012 1078 27568 1112
rect 28030 1078 28586 1112
rect 29048 1078 29604 1112
rect 30066 1078 30622 1112
rect 31084 1078 31640 1112
rect 32102 1078 32658 1112
rect 33120 1078 33676 1112
rect 1148 558 1704 592
rect 2166 558 2722 592
rect 3184 558 3740 592
rect 4202 558 4758 592
rect 5220 558 5776 592
rect 6238 558 6794 592
rect 7256 558 7812 592
rect 8274 558 8830 592
rect 9292 558 9848 592
rect 10310 558 10866 592
rect -1030 240 -996 274
rect 13778 368 14334 402
rect 14796 368 15352 402
rect 15814 368 16370 402
rect 16832 368 17388 402
rect 17850 368 18406 402
rect 18868 368 19424 402
rect 19886 368 20442 402
rect 20904 368 21460 402
rect 21922 368 22478 402
rect 22940 368 23496 402
rect 23958 368 24514 402
rect 24976 368 25532 402
rect 25994 368 26550 402
rect 27012 368 27568 402
rect 28030 368 28586 402
rect 29048 368 29604 402
rect 30066 368 30622 402
rect 31084 368 31640 402
rect 32102 368 32658 402
rect 33120 368 33676 402
rect -1030 0 -996 34
rect 37006 13045 37106 13079
rect 37264 13045 37364 13079
rect 37522 13045 37622 13079
rect 37780 13045 37880 13079
rect 38038 13045 38138 13079
rect 38296 13045 38396 13079
rect 37006 12717 37106 12751
rect 37264 12717 37364 12751
rect 37522 12717 37622 12751
rect 37780 12717 37880 12751
rect 38038 12717 38138 12751
rect 38296 12717 38396 12751
rect 54780 14372 55336 14406
rect 55798 14372 56354 14406
rect 56816 14372 57372 14406
rect 57834 14372 58390 14406
rect 58852 14372 59408 14406
rect 59870 14372 60426 14406
rect 60888 14372 61444 14406
rect 61906 14372 62462 14406
rect 62924 14372 63480 14406
rect 63942 14372 64498 14406
rect 64960 14372 65516 14406
rect 65978 14372 66534 14406
rect 66996 14372 67552 14406
rect 68014 14372 68570 14406
rect 69032 14372 69588 14406
rect 70050 14372 70606 14406
rect 71068 14372 71624 14406
rect 72086 14372 72642 14406
rect 73104 14372 73660 14406
rect 74122 14372 74678 14406
rect 43014 13896 43570 13930
rect 44032 13896 44588 13930
rect 45050 13896 45606 13930
rect 46068 13896 46624 13930
rect 47086 13896 47642 13930
rect 48104 13896 48660 13930
rect 49122 13896 49678 13930
rect 50140 13896 50696 13930
rect 51158 13896 51714 13930
rect 54780 13662 55336 13696
rect 55798 13662 56354 13696
rect 56816 13662 57372 13696
rect 57834 13662 58390 13696
rect 58852 13662 59408 13696
rect 59870 13662 60426 13696
rect 60888 13662 61444 13696
rect 61906 13662 62462 13696
rect 62924 13662 63480 13696
rect 63942 13662 64498 13696
rect 64960 13662 65516 13696
rect 65978 13662 66534 13696
rect 66996 13662 67552 13696
rect 68014 13662 68570 13696
rect 69032 13662 69588 13696
rect 70050 13662 70606 13696
rect 71068 13662 71624 13696
rect 72086 13662 72642 13696
rect 73104 13662 73660 13696
rect 74122 13662 74678 13696
rect 54780 13554 55336 13588
rect 55798 13554 56354 13588
rect 56816 13554 57372 13588
rect 57834 13554 58390 13588
rect 58852 13554 59408 13588
rect 59870 13554 60426 13588
rect 60888 13554 61444 13588
rect 61906 13554 62462 13588
rect 62924 13554 63480 13588
rect 63942 13554 64498 13588
rect 64960 13554 65516 13588
rect 65978 13554 66534 13588
rect 66996 13554 67552 13588
rect 68014 13554 68570 13588
rect 69032 13554 69588 13588
rect 70050 13554 70606 13588
rect 71068 13554 71624 13588
rect 72086 13554 72642 13588
rect 73104 13554 73660 13588
rect 74122 13554 74678 13588
rect 43014 13186 43570 13220
rect 44032 13186 44588 13220
rect 43014 13078 43570 13112
rect 45050 13186 45606 13220
rect 44032 13078 44588 13112
rect 46068 13186 46624 13220
rect 45050 13078 45606 13112
rect 47086 13186 47642 13220
rect 46068 13078 46624 13112
rect 48104 13186 48660 13220
rect 47086 13078 47642 13112
rect 49122 13186 49678 13220
rect 48104 13078 48660 13112
rect 50140 13186 50696 13220
rect 49122 13078 49678 13112
rect 51158 13186 51714 13220
rect 50140 13078 50696 13112
rect 51158 13078 51714 13112
rect 54780 12844 55336 12878
rect 55798 12844 56354 12878
rect 56816 12844 57372 12878
rect 57834 12844 58390 12878
rect 58852 12844 59408 12878
rect 59870 12844 60426 12878
rect 60888 12844 61444 12878
rect 61906 12844 62462 12878
rect 62924 12844 63480 12878
rect 63942 12844 64498 12878
rect 64960 12844 65516 12878
rect 65978 12844 66534 12878
rect 66996 12844 67552 12878
rect 68014 12844 68570 12878
rect 69032 12844 69588 12878
rect 70050 12844 70606 12878
rect 71068 12844 71624 12878
rect 72086 12844 72642 12878
rect 73104 12844 73660 12878
rect 74122 12844 74678 12878
rect 43014 12368 43570 12402
rect 44032 12368 44588 12402
rect 43014 12260 43570 12294
rect 45050 12368 45606 12402
rect 44032 12260 44588 12294
rect 46068 12368 46624 12402
rect 45050 12260 45606 12294
rect 47086 12368 47642 12402
rect 46068 12260 46624 12294
rect 48104 12368 48660 12402
rect 47086 12260 47642 12294
rect 49122 12368 49678 12402
rect 48104 12260 48660 12294
rect 50140 12368 50696 12402
rect 49122 12260 49678 12294
rect 51158 12368 51714 12402
rect 50140 12260 50696 12294
rect 51158 12260 51714 12294
rect 54780 12176 55336 12210
rect 55798 12176 56354 12210
rect 56816 12176 57372 12210
rect 57834 12176 58390 12210
rect 58852 12176 59408 12210
rect 59870 12176 60426 12210
rect 60888 12176 61444 12210
rect 61906 12176 62462 12210
rect 62924 12176 63480 12210
rect 63942 12176 64498 12210
rect 64960 12176 65516 12210
rect 65978 12176 66534 12210
rect 66996 12176 67552 12210
rect 68014 12176 68570 12210
rect 69032 12176 69588 12210
rect 70050 12176 70606 12210
rect 71068 12176 71624 12210
rect 72086 12176 72642 12210
rect 73104 12176 73660 12210
rect 74122 12176 74678 12210
rect 43014 11550 43570 11584
rect 44032 11550 44588 11584
rect 43014 11442 43570 11476
rect 45050 11550 45606 11584
rect 44032 11442 44588 11476
rect 46068 11550 46624 11584
rect 45050 11442 45606 11476
rect 47086 11550 47642 11584
rect 46068 11442 46624 11476
rect 48104 11550 48660 11584
rect 47086 11442 47642 11476
rect 49122 11550 49678 11584
rect 48104 11442 48660 11476
rect 50140 11550 50696 11584
rect 49122 11442 49678 11476
rect 51158 11550 51714 11584
rect 50140 11442 50696 11476
rect 51158 11442 51714 11476
rect 54780 11466 55336 11500
rect 55798 11466 56354 11500
rect 56816 11466 57372 11500
rect 57834 11466 58390 11500
rect 58852 11466 59408 11500
rect 59870 11466 60426 11500
rect 60888 11466 61444 11500
rect 61906 11466 62462 11500
rect 62924 11466 63480 11500
rect 63942 11466 64498 11500
rect 64960 11466 65516 11500
rect 65978 11466 66534 11500
rect 66996 11466 67552 11500
rect 68014 11466 68570 11500
rect 69032 11466 69588 11500
rect 70050 11466 70606 11500
rect 71068 11466 71624 11500
rect 72086 11466 72642 11500
rect 73104 11466 73660 11500
rect 74122 11466 74678 11500
rect 54780 10944 55336 10978
rect 55798 10944 56354 10978
rect 56816 10944 57372 10978
rect 57834 10944 58390 10978
rect 58852 10944 59408 10978
rect 59870 10944 60426 10978
rect 60888 10944 61444 10978
rect 61906 10944 62462 10978
rect 62924 10944 63480 10978
rect 63942 10944 64498 10978
rect 64960 10944 65516 10978
rect 65978 10944 66534 10978
rect 66996 10944 67552 10978
rect 68014 10944 68570 10978
rect 69032 10944 69588 10978
rect 70050 10944 70606 10978
rect 71068 10944 71624 10978
rect 72086 10944 72642 10978
rect 73104 10944 73660 10978
rect 74122 10944 74678 10978
rect 43014 10732 43570 10766
rect 44032 10732 44588 10766
rect 43014 10624 43570 10658
rect 45050 10732 45606 10766
rect 44032 10624 44588 10658
rect 46068 10732 46624 10766
rect 45050 10624 45606 10658
rect 47086 10732 47642 10766
rect 46068 10624 46624 10658
rect 48104 10732 48660 10766
rect 47086 10624 47642 10658
rect 49122 10732 49678 10766
rect 48104 10624 48660 10658
rect 50140 10732 50696 10766
rect 49122 10624 49678 10658
rect 51158 10732 51714 10766
rect 50140 10624 50696 10658
rect 51158 10624 51714 10658
rect 54780 10234 55336 10268
rect 55798 10234 56354 10268
rect 56816 10234 57372 10268
rect 57834 10234 58390 10268
rect 58852 10234 59408 10268
rect 59870 10234 60426 10268
rect 60888 10234 61444 10268
rect 61906 10234 62462 10268
rect 62924 10234 63480 10268
rect 63942 10234 64498 10268
rect 64960 10234 65516 10268
rect 65978 10234 66534 10268
rect 66996 10234 67552 10268
rect 68014 10234 68570 10268
rect 69032 10234 69588 10268
rect 70050 10234 70606 10268
rect 71068 10234 71624 10268
rect 72086 10234 72642 10268
rect 73104 10234 73660 10268
rect 74122 10234 74678 10268
rect 43014 9914 43570 9948
rect 44032 9914 44588 9948
rect 43014 9806 43570 9840
rect 45050 9914 45606 9948
rect 44032 9806 44588 9840
rect 46068 9914 46624 9948
rect 45050 9806 45606 9840
rect 47086 9914 47642 9948
rect 46068 9806 46624 9840
rect 48104 9914 48660 9948
rect 47086 9806 47642 9840
rect 49122 9914 49678 9948
rect 48104 9806 48660 9840
rect 50140 9914 50696 9948
rect 49122 9806 49678 9840
rect 51158 9914 51714 9948
rect 50140 9806 50696 9840
rect 51158 9806 51714 9840
rect 54778 9710 55334 9744
rect 55796 9710 56352 9744
rect 56814 9710 57370 9744
rect 57832 9710 58388 9744
rect 58850 9710 59406 9744
rect 59868 9710 60424 9744
rect 60886 9710 61442 9744
rect 61904 9710 62460 9744
rect 62922 9710 63478 9744
rect 63940 9710 64496 9744
rect 64958 9710 65514 9744
rect 65976 9710 66532 9744
rect 66994 9710 67550 9744
rect 68012 9710 68568 9744
rect 69030 9710 69586 9744
rect 70048 9710 70604 9744
rect 71066 9710 71622 9744
rect 72084 9710 72640 9744
rect 73102 9710 73658 9744
rect 74120 9710 74676 9744
rect 43014 9096 43570 9130
rect 44032 9096 44588 9130
rect 43014 8988 43570 9022
rect 45050 9096 45606 9130
rect 44032 8988 44588 9022
rect 46068 9096 46624 9130
rect 45050 8988 45606 9022
rect 47086 9096 47642 9130
rect 46068 8988 46624 9022
rect 48104 9096 48660 9130
rect 47086 8988 47642 9022
rect 49122 9096 49678 9130
rect 48104 8988 48660 9022
rect 50140 9096 50696 9130
rect 49122 8988 49678 9022
rect 51158 9096 51714 9130
rect 50140 8988 50696 9022
rect 51158 8988 51714 9022
rect 54778 9000 55334 9034
rect 55796 9000 56352 9034
rect 56814 9000 57370 9034
rect 57832 9000 58388 9034
rect 58850 9000 59406 9034
rect 59868 9000 60424 9034
rect 60886 9000 61442 9034
rect 61904 9000 62460 9034
rect 62922 9000 63478 9034
rect 63940 9000 64496 9034
rect 64958 9000 65514 9034
rect 65976 9000 66532 9034
rect 66994 9000 67550 9034
rect 68012 9000 68568 9034
rect 69030 9000 69586 9034
rect 70048 9000 70604 9034
rect 71066 9000 71622 9034
rect 72084 9000 72640 9034
rect 73102 9000 73658 9034
rect 74120 9000 74676 9034
rect 54778 8476 55334 8510
rect 55796 8476 56352 8510
rect 56814 8476 57370 8510
rect 57832 8476 58388 8510
rect 58850 8476 59406 8510
rect 59868 8476 60424 8510
rect 60886 8476 61442 8510
rect 61904 8476 62460 8510
rect 62922 8476 63478 8510
rect 63940 8476 64496 8510
rect 64958 8476 65514 8510
rect 65976 8476 66532 8510
rect 66994 8476 67550 8510
rect 68012 8476 68568 8510
rect 69030 8476 69586 8510
rect 70048 8476 70604 8510
rect 71066 8476 71622 8510
rect 72084 8476 72640 8510
rect 73102 8476 73658 8510
rect 74120 8476 74676 8510
rect 43014 8278 43570 8312
rect 44032 8278 44588 8312
rect 43014 8170 43570 8204
rect 45050 8278 45606 8312
rect 44032 8170 44588 8204
rect 46068 8278 46624 8312
rect 45050 8170 45606 8204
rect 47086 8278 47642 8312
rect 46068 8170 46624 8204
rect 48104 8278 48660 8312
rect 47086 8170 47642 8204
rect 49122 8278 49678 8312
rect 48104 8170 48660 8204
rect 50140 8278 50696 8312
rect 49122 8170 49678 8204
rect 51158 8278 51714 8312
rect 50140 8170 50696 8204
rect 51158 8170 51714 8204
rect 54778 7766 55334 7800
rect 55796 7766 56352 7800
rect 56814 7766 57370 7800
rect 57832 7766 58388 7800
rect 58850 7766 59406 7800
rect 59868 7766 60424 7800
rect 60886 7766 61442 7800
rect 61904 7766 62460 7800
rect 62922 7766 63478 7800
rect 63940 7766 64496 7800
rect 64958 7766 65514 7800
rect 65976 7766 66532 7800
rect 66994 7766 67550 7800
rect 68012 7766 68568 7800
rect 69030 7766 69586 7800
rect 70048 7766 70604 7800
rect 71066 7766 71622 7800
rect 72084 7766 72640 7800
rect 73102 7766 73658 7800
rect 74120 7766 74676 7800
rect 43014 7460 43570 7494
rect 44032 7460 44588 7494
rect 45050 7460 45606 7494
rect 46068 7460 46624 7494
rect 47086 7460 47642 7494
rect 48104 7460 48660 7494
rect 49122 7460 49678 7494
rect 50140 7460 50696 7494
rect 51158 7460 51714 7494
rect 54778 7244 55334 7278
rect 55796 7244 56352 7278
rect 56814 7244 57370 7278
rect 57832 7244 58388 7278
rect 58850 7244 59406 7278
rect 59868 7244 60424 7278
rect 60886 7244 61442 7278
rect 61904 7244 62460 7278
rect 62922 7244 63478 7278
rect 63940 7244 64496 7278
rect 64958 7244 65514 7278
rect 65976 7244 66532 7278
rect 66994 7244 67550 7278
rect 68012 7244 68568 7278
rect 69030 7244 69586 7278
rect 70048 7244 70604 7278
rect 71066 7244 71622 7278
rect 72084 7244 72640 7278
rect 73102 7244 73658 7278
rect 74120 7244 74676 7278
rect 54778 6534 55334 6568
rect 55796 6534 56352 6568
rect 56814 6534 57370 6568
rect 57832 6534 58388 6568
rect 58850 6534 59406 6568
rect 59868 6534 60424 6568
rect 60886 6534 61442 6568
rect 61904 6534 62460 6568
rect 62922 6534 63478 6568
rect 63940 6534 64496 6568
rect 64958 6534 65514 6568
rect 65976 6534 66532 6568
rect 66994 6534 67550 6568
rect 68012 6534 68568 6568
rect 69030 6534 69586 6568
rect 70048 6534 70604 6568
rect 71066 6534 71622 6568
rect 72084 6534 72640 6568
rect 73102 6534 73658 6568
rect 74120 6534 74676 6568
rect 41690 6146 42246 6180
rect 42708 6146 43264 6180
rect 43726 6146 44282 6180
rect 44744 6146 45300 6180
rect 45762 6146 46318 6180
rect 46780 6146 47336 6180
rect 47798 6146 48354 6180
rect 48816 6146 49372 6180
rect 49834 6146 50390 6180
rect 50852 6146 51408 6180
rect 51870 6146 52426 6180
rect 54778 6010 55334 6044
rect 55796 6010 56352 6044
rect 56814 6010 57370 6044
rect 57832 6010 58388 6044
rect 58850 6010 59406 6044
rect 59868 6010 60424 6044
rect 60886 6010 61442 6044
rect 61904 6010 62460 6044
rect 62922 6010 63478 6044
rect 63940 6010 64496 6044
rect 64958 6010 65514 6044
rect 65976 6010 66532 6044
rect 66994 6010 67550 6044
rect 68012 6010 68568 6044
rect 69030 6010 69586 6044
rect 70048 6010 70604 6044
rect 71066 6010 71622 6044
rect 72084 6010 72640 6044
rect 73102 6010 73658 6044
rect 74120 6010 74676 6044
rect 41690 5436 42246 5470
rect 42708 5436 43264 5470
rect 43726 5436 44282 5470
rect 44744 5436 45300 5470
rect 45762 5436 46318 5470
rect 46780 5436 47336 5470
rect 47798 5436 48354 5470
rect 48816 5436 49372 5470
rect 49834 5436 50390 5470
rect 50852 5436 51408 5470
rect 51870 5436 52426 5470
rect 54778 5300 55334 5334
rect 55796 5300 56352 5334
rect 56814 5300 57370 5334
rect 57832 5300 58388 5334
rect 58850 5300 59406 5334
rect 59868 5300 60424 5334
rect 60886 5300 61442 5334
rect 61904 5300 62460 5334
rect 62922 5300 63478 5334
rect 63940 5300 64496 5334
rect 64958 5300 65514 5334
rect 65976 5300 66532 5334
rect 66994 5300 67550 5334
rect 68012 5300 68568 5334
rect 69030 5300 69586 5334
rect 70048 5300 70604 5334
rect 71066 5300 71622 5334
rect 72084 5300 72640 5334
rect 73102 5300 73658 5334
rect 74120 5300 74676 5334
rect 41690 5034 42246 5068
rect 42708 5034 43264 5068
rect 43726 5034 44282 5068
rect 44744 5034 45300 5068
rect 45762 5034 46318 5068
rect 46780 5034 47336 5068
rect 47798 5034 48354 5068
rect 48816 5034 49372 5068
rect 49834 5034 50390 5068
rect 50852 5034 51408 5068
rect 51870 5034 52426 5068
rect 54778 4776 55334 4810
rect 55796 4776 56352 4810
rect 56814 4776 57370 4810
rect 57832 4776 58388 4810
rect 58850 4776 59406 4810
rect 59868 4776 60424 4810
rect 60886 4776 61442 4810
rect 61904 4776 62460 4810
rect 62922 4776 63478 4810
rect 63940 4776 64496 4810
rect 64958 4776 65514 4810
rect 65976 4776 66532 4810
rect 66994 4776 67550 4810
rect 68012 4776 68568 4810
rect 69030 4776 69586 4810
rect 70048 4776 70604 4810
rect 71066 4776 71622 4810
rect 72084 4776 72640 4810
rect 73102 4776 73658 4810
rect 74120 4776 74676 4810
rect 41690 4324 42246 4358
rect 42708 4324 43264 4358
rect 43726 4324 44282 4358
rect 44744 4324 45300 4358
rect 45762 4324 46318 4358
rect 46780 4324 47336 4358
rect 47798 4324 48354 4358
rect 48816 4324 49372 4358
rect 49834 4324 50390 4358
rect 50852 4324 51408 4358
rect 51870 4324 52426 4358
rect 54778 4066 55334 4100
rect 55796 4066 56352 4100
rect 56814 4066 57370 4100
rect 57832 4066 58388 4100
rect 58850 4066 59406 4100
rect 59868 4066 60424 4100
rect 60886 4066 61442 4100
rect 61904 4066 62460 4100
rect 62922 4066 63478 4100
rect 63940 4066 64496 4100
rect 64958 4066 65514 4100
rect 65976 4066 66532 4100
rect 66994 4066 67550 4100
rect 68012 4066 68568 4100
rect 69030 4066 69586 4100
rect 70048 4066 70604 4100
rect 71066 4066 71622 4100
rect 72084 4066 72640 4100
rect 73102 4066 73658 4100
rect 74120 4066 74676 4100
rect 41690 3922 42246 3956
rect 42708 3922 43264 3956
rect 43726 3922 44282 3956
rect 44744 3922 45300 3956
rect 45762 3922 46318 3956
rect 46780 3922 47336 3956
rect 47798 3922 48354 3956
rect 48816 3922 49372 3956
rect 49834 3922 50390 3956
rect 50852 3922 51408 3956
rect 51870 3922 52426 3956
rect 54778 3544 55334 3578
rect 55796 3544 56352 3578
rect 56814 3544 57370 3578
rect 57832 3544 58388 3578
rect 58850 3544 59406 3578
rect 59868 3544 60424 3578
rect 60886 3544 61442 3578
rect 61904 3544 62460 3578
rect 62922 3544 63478 3578
rect 63940 3544 64496 3578
rect 64958 3544 65514 3578
rect 65976 3544 66532 3578
rect 66994 3544 67550 3578
rect 68012 3544 68568 3578
rect 69030 3544 69586 3578
rect 70048 3544 70604 3578
rect 71066 3544 71622 3578
rect 72084 3544 72640 3578
rect 73102 3544 73658 3578
rect 74120 3544 74676 3578
rect 41690 3212 42246 3246
rect 42708 3212 43264 3246
rect 43726 3212 44282 3246
rect 44744 3212 45300 3246
rect 45762 3212 46318 3246
rect 46780 3212 47336 3246
rect 47798 3212 48354 3246
rect 48816 3212 49372 3246
rect 49834 3212 50390 3246
rect 50852 3212 51408 3246
rect 51870 3212 52426 3246
rect 41690 2810 42246 2844
rect 42708 2810 43264 2844
rect 43726 2810 44282 2844
rect 44744 2810 45300 2844
rect 45762 2810 46318 2844
rect 46780 2810 47336 2844
rect 47798 2810 48354 2844
rect 48816 2810 49372 2844
rect 49834 2810 50390 2844
rect 50852 2810 51408 2844
rect 51870 2810 52426 2844
rect 54778 2834 55334 2868
rect 55796 2834 56352 2868
rect 56814 2834 57370 2868
rect 57832 2834 58388 2868
rect 58850 2834 59406 2868
rect 59868 2834 60424 2868
rect 60886 2834 61442 2868
rect 61904 2834 62460 2868
rect 62922 2834 63478 2868
rect 63940 2834 64496 2868
rect 64958 2834 65514 2868
rect 65976 2834 66532 2868
rect 66994 2834 67550 2868
rect 68012 2834 68568 2868
rect 69030 2834 69586 2868
rect 70048 2834 70604 2868
rect 71066 2834 71622 2868
rect 72084 2834 72640 2868
rect 73102 2834 73658 2868
rect 74120 2834 74676 2868
rect 54778 2310 55334 2344
rect 55796 2310 56352 2344
rect 56814 2310 57370 2344
rect 57832 2310 58388 2344
rect 58850 2310 59406 2344
rect 59868 2310 60424 2344
rect 60886 2310 61442 2344
rect 61904 2310 62460 2344
rect 62922 2310 63478 2344
rect 63940 2310 64496 2344
rect 64958 2310 65514 2344
rect 65976 2310 66532 2344
rect 66994 2310 67550 2344
rect 68012 2310 68568 2344
rect 69030 2310 69586 2344
rect 70048 2310 70604 2344
rect 71066 2310 71622 2344
rect 72084 2310 72640 2344
rect 73102 2310 73658 2344
rect 74120 2310 74676 2344
rect 41690 2100 42246 2134
rect 42708 2100 43264 2134
rect 43726 2100 44282 2134
rect 44744 2100 45300 2134
rect 45762 2100 46318 2134
rect 46780 2100 47336 2134
rect 47798 2100 48354 2134
rect 48816 2100 49372 2134
rect 49834 2100 50390 2134
rect 50852 2100 51408 2134
rect 51870 2100 52426 2134
rect 54778 1600 55334 1634
rect 55796 1600 56352 1634
rect 56814 1600 57370 1634
rect 57832 1600 58388 1634
rect 58850 1600 59406 1634
rect 59868 1600 60424 1634
rect 60886 1600 61442 1634
rect 61904 1600 62460 1634
rect 62922 1600 63478 1634
rect 63940 1600 64496 1634
rect 64958 1600 65514 1634
rect 65976 1600 66532 1634
rect 66994 1600 67550 1634
rect 68012 1600 68568 1634
rect 69030 1600 69586 1634
rect 70048 1600 70604 1634
rect 71066 1600 71622 1634
rect 72084 1600 72640 1634
rect 73102 1600 73658 1634
rect 74120 1600 74676 1634
rect 42148 1268 42704 1302
rect 43166 1268 43722 1302
rect 44184 1268 44740 1302
rect 45202 1268 45758 1302
rect 46220 1268 46776 1302
rect 47238 1268 47794 1302
rect 48256 1268 48812 1302
rect 49274 1268 49830 1302
rect 50292 1268 50848 1302
rect 51310 1268 51866 1302
rect 54778 1078 55334 1112
rect 55796 1078 56352 1112
rect 56814 1078 57370 1112
rect 57832 1078 58388 1112
rect 58850 1078 59406 1112
rect 59868 1078 60424 1112
rect 60886 1078 61442 1112
rect 61904 1078 62460 1112
rect 62922 1078 63478 1112
rect 63940 1078 64496 1112
rect 64958 1078 65514 1112
rect 65976 1078 66532 1112
rect 66994 1078 67550 1112
rect 68012 1078 68568 1112
rect 69030 1078 69586 1112
rect 70048 1078 70604 1112
rect 71066 1078 71622 1112
rect 72084 1078 72640 1112
rect 73102 1078 73658 1112
rect 74120 1078 74676 1112
rect 42148 558 42704 592
rect 43166 558 43722 592
rect 44184 558 44740 592
rect 45202 558 45758 592
rect 46220 558 46776 592
rect 47238 558 47794 592
rect 48256 558 48812 592
rect 49274 558 49830 592
rect 50292 558 50848 592
rect 51310 558 51866 592
rect 54778 368 55334 402
rect 55796 368 56352 402
rect 56814 368 57370 402
rect 57832 368 58388 402
rect 58850 368 59406 402
rect 59868 368 60424 402
rect 60886 368 61442 402
rect 61904 368 62460 402
rect 62922 368 63478 402
rect 63940 368 64496 402
rect 64958 368 65514 402
rect 65976 368 66532 402
rect 66994 368 67550 402
rect 68012 368 68568 402
rect 69030 368 69586 402
rect 70048 368 70604 402
rect 71066 368 71622 402
rect 72084 368 72640 402
rect 73102 368 73658 402
rect 74120 368 74676 402
<< locali >>
rect 11328 30530 11428 30692
rect 35672 30530 35772 30692
rect 17918 28148 18008 28178
rect 17918 28114 17946 28148
rect 17980 28114 18008 28148
rect 17918 28086 18008 28114
rect 18936 28148 19026 28178
rect 18936 28114 18964 28148
rect 18998 28114 19026 28148
rect 18936 28086 19026 28114
rect 19954 28148 20044 28178
rect 19954 28114 19982 28148
rect 20016 28114 20044 28148
rect 19954 28086 20044 28114
rect 20972 28148 21062 28178
rect 20972 28114 21000 28148
rect 21034 28114 21062 28148
rect 20972 28086 21062 28114
rect 21990 28148 22080 28178
rect 21990 28114 22018 28148
rect 22052 28114 22080 28148
rect 21990 28086 22080 28114
rect 23008 28148 23098 28178
rect 23008 28114 23036 28148
rect 23070 28114 23098 28148
rect 23008 28086 23098 28114
rect 24026 28148 24116 28178
rect 24026 28114 24054 28148
rect 24088 28114 24116 28148
rect 24026 28086 24116 28114
rect 25044 28148 25134 28178
rect 25044 28114 25072 28148
rect 25106 28114 25134 28148
rect 25044 28086 25134 28114
rect 26062 28148 26152 28178
rect 26062 28114 26090 28148
rect 26124 28114 26152 28148
rect 26062 28086 26152 28114
rect 27080 28148 27170 28178
rect 27080 28114 27108 28148
rect 27142 28114 27170 28148
rect 27080 28086 27170 28114
rect 28098 28148 28188 28178
rect 28098 28114 28126 28148
rect 28160 28114 28188 28148
rect 28098 28086 28188 28114
rect 29116 28148 29206 28178
rect 29116 28114 29144 28148
rect 29178 28114 29206 28148
rect 29116 28086 29206 28114
rect 30134 28148 30224 28178
rect 30134 28114 30162 28148
rect 30196 28114 30224 28148
rect 30134 28086 30224 28114
rect 31152 28148 31242 28178
rect 31152 28114 31180 28148
rect 31214 28114 31242 28148
rect 31152 28086 31242 28114
rect 32170 28148 32260 28178
rect 32170 28114 32198 28148
rect 32232 28114 32260 28148
rect 32170 28086 32260 28114
rect 33188 28148 33278 28178
rect 33188 28114 33216 28148
rect 33250 28114 33278 28148
rect 33188 28086 33278 28114
rect 17670 27891 17686 27925
rect 18242 27891 18258 27925
rect 18688 27891 18704 27925
rect 19260 27891 19276 27925
rect 19706 27891 19722 27925
rect 20278 27891 20294 27925
rect 20724 27891 20740 27925
rect 21296 27891 21312 27925
rect 21742 27891 21758 27925
rect 22314 27891 22330 27925
rect 22760 27891 22776 27925
rect 23332 27891 23348 27925
rect 23778 27891 23794 27925
rect 24350 27891 24366 27925
rect 24796 27891 24812 27925
rect 25368 27891 25384 27925
rect 25814 27891 25830 27925
rect 26386 27891 26402 27925
rect 26832 27891 26848 27925
rect 27404 27891 27420 27925
rect 27850 27891 27866 27925
rect 28422 27891 28438 27925
rect 28868 27891 28884 27925
rect 29440 27891 29456 27925
rect 29886 27891 29902 27925
rect 30458 27891 30474 27925
rect 30904 27891 30920 27925
rect 31476 27891 31492 27925
rect 31922 27891 31938 27925
rect 32494 27891 32510 27925
rect 32940 27891 32956 27925
rect 33512 27891 33528 27925
rect 17438 27832 17472 27848
rect 17438 27240 17472 27256
rect 18456 27832 18490 27848
rect 18456 27240 18490 27256
rect 19474 27832 19508 27848
rect 19474 27240 19508 27256
rect 20492 27832 20526 27848
rect 20492 27240 20526 27256
rect 21510 27832 21544 27848
rect 21510 27240 21544 27256
rect 22528 27832 22562 27848
rect 22528 27240 22562 27256
rect 23546 27832 23580 27848
rect 23546 27240 23580 27256
rect 24564 27832 24598 27848
rect 24564 27240 24598 27256
rect 25582 27832 25616 27848
rect 25582 27240 25616 27256
rect 26600 27832 26634 27848
rect 26600 27240 26634 27256
rect 27618 27832 27652 27848
rect 27618 27240 27652 27256
rect 28636 27832 28670 27848
rect 28636 27240 28670 27256
rect 29654 27832 29688 27848
rect 29654 27240 29688 27256
rect 30672 27832 30706 27848
rect 30672 27240 30706 27256
rect 31690 27832 31724 27848
rect 31690 27240 31724 27256
rect 32708 27832 32742 27848
rect 32708 27240 32742 27256
rect 33726 27832 33760 27848
rect 33726 27240 33760 27256
rect 17670 27163 17686 27197
rect 18242 27163 18258 27197
rect 18688 27163 18704 27197
rect 19260 27163 19276 27197
rect 19706 27163 19722 27197
rect 20278 27163 20294 27197
rect 20724 27163 20740 27197
rect 21296 27163 21312 27197
rect 21742 27163 21758 27197
rect 22314 27163 22330 27197
rect 22760 27163 22776 27197
rect 23332 27163 23348 27197
rect 23778 27163 23794 27197
rect 24350 27163 24366 27197
rect 24796 27163 24812 27197
rect 25368 27163 25384 27197
rect 25814 27163 25830 27197
rect 26386 27163 26402 27197
rect 26832 27163 26848 27197
rect 27404 27163 27420 27197
rect 27850 27163 27866 27197
rect 28422 27163 28438 27197
rect 28868 27163 28884 27197
rect 29440 27163 29456 27197
rect 29886 27163 29902 27197
rect 30458 27163 30474 27197
rect 30904 27163 30920 27197
rect 31476 27163 31492 27197
rect 31922 27163 31938 27197
rect 32494 27163 32510 27197
rect 32940 27163 32956 27197
rect 33512 27163 33528 27197
rect 17940 26994 18030 27024
rect 17940 26960 17968 26994
rect 18002 26960 18030 26994
rect 17940 26932 18030 26960
rect 18958 26994 19048 27024
rect 18958 26960 18986 26994
rect 19020 26960 19048 26994
rect 18958 26932 19048 26960
rect 19976 26994 20066 27024
rect 19976 26960 20004 26994
rect 20038 26960 20066 26994
rect 19976 26932 20066 26960
rect 20994 26994 21084 27024
rect 20994 26960 21022 26994
rect 21056 26960 21084 26994
rect 20994 26932 21084 26960
rect 22012 26994 22102 27024
rect 22012 26960 22040 26994
rect 22074 26960 22102 26994
rect 22012 26932 22102 26960
rect 23030 26994 23120 27024
rect 23030 26960 23058 26994
rect 23092 26960 23120 26994
rect 23030 26932 23120 26960
rect 24048 26994 24138 27024
rect 24048 26960 24076 26994
rect 24110 26960 24138 26994
rect 24048 26932 24138 26960
rect 25066 26994 25156 27024
rect 25066 26960 25094 26994
rect 25128 26960 25156 26994
rect 25066 26932 25156 26960
rect 26084 26994 26174 27024
rect 26084 26960 26112 26994
rect 26146 26960 26174 26994
rect 26084 26932 26174 26960
rect 27102 26994 27192 27024
rect 27102 26960 27130 26994
rect 27164 26960 27192 26994
rect 27102 26932 27192 26960
rect 28120 26994 28210 27024
rect 28120 26960 28148 26994
rect 28182 26960 28210 26994
rect 28120 26932 28210 26960
rect 29138 26994 29228 27024
rect 29138 26960 29166 26994
rect 29200 26960 29228 26994
rect 29138 26932 29228 26960
rect 30156 26994 30246 27024
rect 30156 26960 30184 26994
rect 30218 26960 30246 26994
rect 30156 26932 30246 26960
rect 31174 26994 31264 27024
rect 31174 26960 31202 26994
rect 31236 26960 31264 26994
rect 31174 26932 31264 26960
rect 32192 26994 32282 27024
rect 32192 26960 32220 26994
rect 32254 26960 32282 26994
rect 32192 26932 32282 26960
rect 33210 26994 33300 27024
rect 33210 26960 33238 26994
rect 33272 26960 33300 26994
rect 33210 26932 33300 26960
rect 17670 26755 17686 26789
rect 18242 26755 18258 26789
rect 18688 26755 18704 26789
rect 19260 26755 19276 26789
rect 19706 26755 19722 26789
rect 20278 26755 20294 26789
rect 20724 26755 20740 26789
rect 21296 26755 21312 26789
rect 21742 26755 21758 26789
rect 22314 26755 22330 26789
rect 22760 26755 22776 26789
rect 23332 26755 23348 26789
rect 23778 26755 23794 26789
rect 24350 26755 24366 26789
rect 24796 26755 24812 26789
rect 25368 26755 25384 26789
rect 25814 26755 25830 26789
rect 26386 26755 26402 26789
rect 26832 26755 26848 26789
rect 27404 26755 27420 26789
rect 27850 26755 27866 26789
rect 28422 26755 28438 26789
rect 28868 26755 28884 26789
rect 29440 26755 29456 26789
rect 29886 26755 29902 26789
rect 30458 26755 30474 26789
rect 30904 26755 30920 26789
rect 31476 26755 31492 26789
rect 31922 26755 31938 26789
rect 32494 26755 32510 26789
rect 32940 26755 32956 26789
rect 33512 26755 33528 26789
rect 17438 26696 17472 26712
rect 17438 26104 17472 26120
rect 18456 26696 18490 26712
rect 18456 26104 18490 26120
rect 19474 26696 19508 26712
rect 19474 26104 19508 26120
rect 20492 26696 20526 26712
rect 20492 26104 20526 26120
rect 21510 26696 21544 26712
rect 21510 26104 21544 26120
rect 22528 26696 22562 26712
rect 22528 26104 22562 26120
rect 23546 26696 23580 26712
rect 23546 26104 23580 26120
rect 24564 26696 24598 26712
rect 24564 26104 24598 26120
rect 25582 26696 25616 26712
rect 25582 26104 25616 26120
rect 26600 26696 26634 26712
rect 26600 26104 26634 26120
rect 27618 26696 27652 26712
rect 27618 26104 27652 26120
rect 28636 26696 28670 26712
rect 28636 26104 28670 26120
rect 29654 26696 29688 26712
rect 29654 26104 29688 26120
rect 30672 26696 30706 26712
rect 30672 26104 30706 26120
rect 31690 26696 31724 26712
rect 31690 26104 31724 26120
rect 32708 26696 32742 26712
rect 32708 26104 32742 26120
rect 33726 26696 33760 26712
rect 33726 26104 33760 26120
rect 17670 26027 17686 26061
rect 18242 26027 18258 26061
rect 18688 26027 18704 26061
rect 19260 26027 19276 26061
rect 19706 26027 19722 26061
rect 20278 26027 20294 26061
rect 20724 26027 20740 26061
rect 21296 26027 21312 26061
rect 21742 26027 21758 26061
rect 22314 26027 22330 26061
rect 22760 26027 22776 26061
rect 23332 26027 23348 26061
rect 23778 26027 23794 26061
rect 24350 26027 24366 26061
rect 24796 26027 24812 26061
rect 25368 26027 25384 26061
rect 25814 26027 25830 26061
rect 26386 26027 26402 26061
rect 26832 26027 26848 26061
rect 27404 26027 27420 26061
rect 27850 26027 27866 26061
rect 28422 26027 28438 26061
rect 28868 26027 28884 26061
rect 29440 26027 29456 26061
rect 29886 26027 29902 26061
rect 30458 26027 30474 26061
rect 30904 26027 30920 26061
rect 31476 26027 31492 26061
rect 31922 26027 31938 26061
rect 32494 26027 32510 26061
rect 32940 26027 32956 26061
rect 33512 26027 33528 26061
rect 17918 25862 18008 25892
rect 17918 25828 17946 25862
rect 17980 25828 18008 25862
rect 17918 25800 18008 25828
rect 18936 25862 19026 25892
rect 18936 25828 18964 25862
rect 18998 25828 19026 25862
rect 18936 25800 19026 25828
rect 19954 25862 20044 25892
rect 19954 25828 19982 25862
rect 20016 25828 20044 25862
rect 19954 25800 20044 25828
rect 20972 25862 21062 25892
rect 20972 25828 21000 25862
rect 21034 25828 21062 25862
rect 20972 25800 21062 25828
rect 21990 25862 22080 25892
rect 21990 25828 22018 25862
rect 22052 25828 22080 25862
rect 21990 25800 22080 25828
rect 23008 25862 23098 25892
rect 23008 25828 23036 25862
rect 23070 25828 23098 25862
rect 23008 25800 23098 25828
rect 24026 25862 24116 25892
rect 24026 25828 24054 25862
rect 24088 25828 24116 25862
rect 24026 25800 24116 25828
rect 25044 25862 25134 25892
rect 25044 25828 25072 25862
rect 25106 25828 25134 25862
rect 25044 25800 25134 25828
rect 26062 25862 26152 25892
rect 26062 25828 26090 25862
rect 26124 25828 26152 25862
rect 26062 25800 26152 25828
rect 27080 25862 27170 25892
rect 27080 25828 27108 25862
rect 27142 25828 27170 25862
rect 27080 25800 27170 25828
rect 28098 25862 28188 25892
rect 28098 25828 28126 25862
rect 28160 25828 28188 25862
rect 28098 25800 28188 25828
rect 29116 25862 29206 25892
rect 29116 25828 29144 25862
rect 29178 25828 29206 25862
rect 29116 25800 29206 25828
rect 30134 25862 30224 25892
rect 30134 25828 30162 25862
rect 30196 25828 30224 25862
rect 30134 25800 30224 25828
rect 31152 25862 31242 25892
rect 31152 25828 31180 25862
rect 31214 25828 31242 25862
rect 31152 25800 31242 25828
rect 32170 25862 32260 25892
rect 32170 25828 32198 25862
rect 32232 25828 32260 25862
rect 32170 25800 32260 25828
rect 33188 25862 33278 25892
rect 33188 25828 33216 25862
rect 33250 25828 33278 25862
rect 33188 25800 33278 25828
rect 17670 25619 17686 25653
rect 18242 25619 18258 25653
rect 18688 25619 18704 25653
rect 19260 25619 19276 25653
rect 19706 25619 19722 25653
rect 20278 25619 20294 25653
rect 20724 25619 20740 25653
rect 21296 25619 21312 25653
rect 21742 25619 21758 25653
rect 22314 25619 22330 25653
rect 22760 25619 22776 25653
rect 23332 25619 23348 25653
rect 23778 25619 23794 25653
rect 24350 25619 24366 25653
rect 24796 25619 24812 25653
rect 25368 25619 25384 25653
rect 25814 25619 25830 25653
rect 26386 25619 26402 25653
rect 26832 25619 26848 25653
rect 27404 25619 27420 25653
rect 27850 25619 27866 25653
rect 28422 25619 28438 25653
rect 28868 25619 28884 25653
rect 29440 25619 29456 25653
rect 29886 25619 29902 25653
rect 30458 25619 30474 25653
rect 30904 25619 30920 25653
rect 31476 25619 31492 25653
rect 31922 25619 31938 25653
rect 32494 25619 32510 25653
rect 32940 25619 32956 25653
rect 33512 25619 33528 25653
rect 17438 25560 17472 25576
rect 17438 24968 17472 24984
rect 18456 25560 18490 25576
rect 18456 24968 18490 24984
rect 19474 25560 19508 25576
rect 19474 24968 19508 24984
rect 20492 25560 20526 25576
rect 20492 24968 20526 24984
rect 21510 25560 21544 25576
rect 21510 24968 21544 24984
rect 22528 25560 22562 25576
rect 22528 24968 22562 24984
rect 23546 25560 23580 25576
rect 23546 24968 23580 24984
rect 24564 25560 24598 25576
rect 24564 24968 24598 24984
rect 25582 25560 25616 25576
rect 25582 24968 25616 24984
rect 26600 25560 26634 25576
rect 26600 24968 26634 24984
rect 27618 25560 27652 25576
rect 27618 24968 27652 24984
rect 28636 25560 28670 25576
rect 28636 24968 28670 24984
rect 29654 25560 29688 25576
rect 29654 24968 29688 24984
rect 30672 25560 30706 25576
rect 30672 24968 30706 24984
rect 31690 25560 31724 25576
rect 31690 24968 31724 24984
rect 32708 25560 32742 25576
rect 32708 24968 32742 24984
rect 33726 25560 33760 25576
rect 33726 24968 33760 24984
rect 17670 24891 17686 24925
rect 18242 24891 18258 24925
rect 18688 24891 18704 24925
rect 19260 24891 19276 24925
rect 19706 24891 19722 24925
rect 20278 24891 20294 24925
rect 20724 24891 20740 24925
rect 21296 24891 21312 24925
rect 21742 24891 21758 24925
rect 22314 24891 22330 24925
rect 22760 24891 22776 24925
rect 23332 24891 23348 24925
rect 23778 24891 23794 24925
rect 24350 24891 24366 24925
rect 24796 24891 24812 24925
rect 25368 24891 25384 24925
rect 25814 24891 25830 24925
rect 26386 24891 26402 24925
rect 26832 24891 26848 24925
rect 27404 24891 27420 24925
rect 27850 24891 27866 24925
rect 28422 24891 28438 24925
rect 28868 24891 28884 24925
rect 29440 24891 29456 24925
rect 29886 24891 29902 24925
rect 30458 24891 30474 24925
rect 30904 24891 30920 24925
rect 31476 24891 31492 24925
rect 31922 24891 31938 24925
rect 32494 24891 32510 24925
rect 32940 24891 32956 24925
rect 33512 24891 33528 24925
rect 17918 24480 18008 24510
rect 17918 24446 17946 24480
rect 17980 24446 18008 24480
rect 17918 24418 18008 24446
rect 18936 24480 19026 24510
rect 18936 24446 18964 24480
rect 18998 24446 19026 24480
rect 18936 24418 19026 24446
rect 19954 24480 20044 24510
rect 19954 24446 19982 24480
rect 20016 24446 20044 24480
rect 19954 24418 20044 24446
rect 20972 24480 21062 24510
rect 20972 24446 21000 24480
rect 21034 24446 21062 24480
rect 20972 24418 21062 24446
rect 21990 24480 22080 24510
rect 21990 24446 22018 24480
rect 22052 24446 22080 24480
rect 21990 24418 22080 24446
rect 23008 24480 23098 24510
rect 23008 24446 23036 24480
rect 23070 24446 23098 24480
rect 23008 24418 23098 24446
rect 24026 24480 24116 24510
rect 24026 24446 24054 24480
rect 24088 24446 24116 24480
rect 24026 24418 24116 24446
rect 25044 24480 25134 24510
rect 25044 24446 25072 24480
rect 25106 24446 25134 24480
rect 25044 24418 25134 24446
rect 26062 24480 26152 24510
rect 26062 24446 26090 24480
rect 26124 24446 26152 24480
rect 26062 24418 26152 24446
rect 27080 24480 27170 24510
rect 27080 24446 27108 24480
rect 27142 24446 27170 24480
rect 27080 24418 27170 24446
rect 28098 24480 28188 24510
rect 28098 24446 28126 24480
rect 28160 24446 28188 24480
rect 28098 24418 28188 24446
rect 29116 24480 29206 24510
rect 29116 24446 29144 24480
rect 29178 24446 29206 24480
rect 29116 24418 29206 24446
rect 30134 24480 30224 24510
rect 30134 24446 30162 24480
rect 30196 24446 30224 24480
rect 30134 24418 30224 24446
rect 31152 24480 31242 24510
rect 31152 24446 31180 24480
rect 31214 24446 31242 24480
rect 31152 24418 31242 24446
rect 32170 24480 32260 24510
rect 32170 24446 32198 24480
rect 32232 24446 32260 24480
rect 32170 24418 32260 24446
rect 33188 24480 33278 24510
rect 33188 24446 33216 24480
rect 33250 24446 33278 24480
rect 33188 24418 33278 24446
rect 18864 23981 18880 24015
rect 19436 23981 19452 24015
rect 19882 23981 19898 24015
rect 20454 23981 20470 24015
rect 20900 23981 20916 24015
rect 21472 23981 21488 24015
rect 21918 23981 21934 24015
rect 22490 23981 22506 24015
rect 22936 23981 22952 24015
rect 23508 23981 23524 24015
rect 23954 23981 23970 24015
rect 24526 23981 24542 24015
rect 24972 23981 24988 24015
rect 25544 23981 25560 24015
rect 25990 23981 26006 24015
rect 26562 23981 26578 24015
rect 27008 23981 27024 24015
rect 27580 23981 27596 24015
rect 28026 23981 28042 24015
rect 28598 23981 28614 24015
rect 29044 23981 29060 24015
rect 29616 23981 29632 24015
rect 30062 23981 30078 24015
rect 30634 23981 30650 24015
rect 31080 23981 31096 24015
rect 31652 23981 31668 24015
rect 32098 23981 32114 24015
rect 32670 23981 32686 24015
rect 18632 23922 18666 23938
rect 18632 23330 18666 23346
rect 19650 23922 19684 23938
rect 19650 23330 19684 23346
rect 20668 23922 20702 23938
rect 20668 23330 20702 23346
rect 21686 23922 21720 23938
rect 21686 23330 21720 23346
rect 22704 23922 22738 23938
rect 22704 23330 22738 23346
rect 23722 23922 23756 23938
rect 23722 23330 23756 23346
rect 24740 23922 24774 23938
rect 24740 23330 24774 23346
rect 25758 23922 25792 23938
rect 25758 23330 25792 23346
rect 26776 23922 26810 23938
rect 26776 23330 26810 23346
rect 27794 23922 27828 23938
rect 27794 23330 27828 23346
rect 28812 23922 28846 23938
rect 28812 23330 28846 23346
rect 29830 23922 29864 23938
rect 29830 23330 29864 23346
rect 30848 23922 30882 23938
rect 30848 23330 30882 23346
rect 31866 23922 31900 23938
rect 31866 23330 31900 23346
rect 32884 23922 32918 23938
rect 32884 23330 32918 23346
rect 18864 23253 18880 23287
rect 19436 23253 19452 23287
rect 19882 23253 19898 23287
rect 20454 23253 20470 23287
rect 20900 23253 20916 23287
rect 21472 23253 21488 23287
rect 21918 23253 21934 23287
rect 22490 23253 22506 23287
rect 22936 23253 22952 23287
rect 23508 23253 23524 23287
rect 23954 23253 23970 23287
rect 24526 23253 24542 23287
rect 24972 23253 24988 23287
rect 25544 23253 25560 23287
rect 25990 23253 26006 23287
rect 26562 23253 26578 23287
rect 27008 23253 27024 23287
rect 27580 23253 27596 23287
rect 28026 23253 28042 23287
rect 28598 23253 28614 23287
rect 29044 23253 29060 23287
rect 29616 23253 29632 23287
rect 30062 23253 30078 23287
rect 30634 23253 30650 23287
rect 31080 23253 31096 23287
rect 31652 23253 31668 23287
rect 32098 23253 32114 23287
rect 32670 23253 32686 23287
rect 18606 23132 18696 23162
rect 18606 23098 18634 23132
rect 18668 23098 18696 23132
rect 18606 23070 18696 23098
rect 19624 23132 19714 23162
rect 19624 23098 19652 23132
rect 19686 23098 19714 23132
rect 19624 23070 19714 23098
rect 20642 23132 20732 23162
rect 20642 23098 20670 23132
rect 20704 23098 20732 23132
rect 20642 23070 20732 23098
rect 21660 23132 21750 23162
rect 21660 23098 21688 23132
rect 21722 23098 21750 23132
rect 21660 23070 21750 23098
rect 22678 23132 22768 23162
rect 22678 23098 22706 23132
rect 22740 23098 22768 23132
rect 22678 23070 22768 23098
rect 23696 23132 23786 23162
rect 23696 23098 23724 23132
rect 23758 23098 23786 23132
rect 23696 23070 23786 23098
rect 24714 23132 24804 23162
rect 24714 23098 24742 23132
rect 24776 23098 24804 23132
rect 24714 23070 24804 23098
rect 25732 23132 25822 23162
rect 25732 23098 25760 23132
rect 25794 23098 25822 23132
rect 25732 23070 25822 23098
rect 26750 23132 26840 23162
rect 26750 23098 26778 23132
rect 26812 23098 26840 23132
rect 26750 23070 26840 23098
rect 27768 23132 27858 23162
rect 27768 23098 27796 23132
rect 27830 23098 27858 23132
rect 27768 23070 27858 23098
rect 28786 23132 28876 23162
rect 28786 23098 28814 23132
rect 28848 23098 28876 23132
rect 28786 23070 28876 23098
rect 29804 23132 29894 23162
rect 29804 23098 29832 23132
rect 29866 23098 29894 23132
rect 29804 23070 29894 23098
rect 30822 23132 30912 23162
rect 30822 23098 30850 23132
rect 30884 23098 30912 23132
rect 30822 23070 30912 23098
rect 31840 23132 31930 23162
rect 31840 23098 31868 23132
rect 31902 23098 31930 23132
rect 31840 23070 31930 23098
rect 32858 23132 32948 23162
rect 32858 23098 32886 23132
rect 32920 23098 32948 23132
rect 32858 23070 32948 23098
rect 18864 22949 18880 22983
rect 19436 22949 19452 22983
rect 19882 22949 19898 22983
rect 20454 22949 20470 22983
rect 20900 22949 20916 22983
rect 21472 22949 21488 22983
rect 21918 22949 21934 22983
rect 22490 22949 22506 22983
rect 22936 22949 22952 22983
rect 23508 22949 23524 22983
rect 23954 22949 23970 22983
rect 24526 22949 24542 22983
rect 24972 22949 24988 22983
rect 25544 22949 25560 22983
rect 25990 22949 26006 22983
rect 26562 22949 26578 22983
rect 27008 22949 27024 22983
rect 27580 22949 27596 22983
rect 28026 22949 28042 22983
rect 28598 22949 28614 22983
rect 29044 22949 29060 22983
rect 29616 22949 29632 22983
rect 30062 22949 30078 22983
rect 30634 22949 30650 22983
rect 31080 22949 31096 22983
rect 31652 22949 31668 22983
rect 32098 22949 32114 22983
rect 32670 22949 32686 22983
rect 18632 22890 18666 22906
rect 18632 22298 18666 22314
rect 19650 22890 19684 22906
rect 19650 22298 19684 22314
rect 20668 22890 20702 22906
rect 20668 22298 20702 22314
rect 21686 22890 21720 22906
rect 21686 22298 21720 22314
rect 22704 22890 22738 22906
rect 22704 22298 22738 22314
rect 23722 22890 23756 22906
rect 23722 22298 23756 22314
rect 24740 22890 24774 22906
rect 24740 22298 24774 22314
rect 25758 22890 25792 22906
rect 25758 22298 25792 22314
rect 26776 22890 26810 22906
rect 26776 22298 26810 22314
rect 27794 22890 27828 22906
rect 27794 22298 27828 22314
rect 28812 22890 28846 22906
rect 28812 22298 28846 22314
rect 29830 22890 29864 22906
rect 29830 22298 29864 22314
rect 30848 22890 30882 22906
rect 30848 22298 30882 22314
rect 31866 22890 31900 22906
rect 31866 22298 31900 22314
rect 32884 22890 32918 22906
rect 32884 22298 32918 22314
rect 18864 22221 18880 22255
rect 19436 22221 19452 22255
rect 19882 22221 19898 22255
rect 20454 22221 20470 22255
rect 20900 22221 20916 22255
rect 21472 22221 21488 22255
rect 21918 22221 21934 22255
rect 22490 22221 22506 22255
rect 22936 22221 22952 22255
rect 23508 22221 23524 22255
rect 23954 22221 23970 22255
rect 24526 22221 24542 22255
rect 24972 22221 24988 22255
rect 25544 22221 25560 22255
rect 25990 22221 26006 22255
rect 26562 22221 26578 22255
rect 27008 22221 27024 22255
rect 27580 22221 27596 22255
rect 28026 22221 28042 22255
rect 28598 22221 28614 22255
rect 29044 22221 29060 22255
rect 29616 22221 29632 22255
rect 30062 22221 30078 22255
rect 30634 22221 30650 22255
rect 31080 22221 31096 22255
rect 31652 22221 31668 22255
rect 32098 22221 32114 22255
rect 32670 22221 32686 22255
rect 18212 21854 18302 21884
rect 18212 21820 18240 21854
rect 18274 21820 18302 21854
rect 18212 21792 18302 21820
rect 19230 21854 19320 21884
rect 19230 21820 19258 21854
rect 19292 21820 19320 21854
rect 19230 21792 19320 21820
rect 20248 21854 20338 21884
rect 20248 21820 20276 21854
rect 20310 21820 20338 21854
rect 20248 21792 20338 21820
rect 21266 21854 21356 21884
rect 21266 21820 21294 21854
rect 21328 21820 21356 21854
rect 21266 21792 21356 21820
rect 22284 21854 22374 21884
rect 22284 21820 22312 21854
rect 22346 21820 22374 21854
rect 22284 21792 22374 21820
rect 23302 21854 23392 21884
rect 23302 21820 23330 21854
rect 23364 21820 23392 21854
rect 23302 21792 23392 21820
rect 24320 21854 24410 21884
rect 24320 21820 24348 21854
rect 24382 21820 24410 21854
rect 24320 21792 24410 21820
rect 25338 21854 25428 21884
rect 25338 21820 25366 21854
rect 25400 21820 25428 21854
rect 25338 21792 25428 21820
rect 26356 21854 26446 21884
rect 26356 21820 26384 21854
rect 26418 21820 26446 21854
rect 26356 21792 26446 21820
rect 27374 21854 27464 21884
rect 27374 21820 27402 21854
rect 27436 21820 27464 21854
rect 27374 21792 27464 21820
rect 28392 21854 28482 21884
rect 28392 21820 28420 21854
rect 28454 21820 28482 21854
rect 28392 21792 28482 21820
rect 29410 21854 29500 21884
rect 29410 21820 29438 21854
rect 29472 21820 29500 21854
rect 29410 21792 29500 21820
rect 30428 21854 30518 21884
rect 30428 21820 30456 21854
rect 30490 21820 30518 21854
rect 30428 21792 30518 21820
rect 31446 21854 31536 21884
rect 31446 21820 31474 21854
rect 31508 21820 31536 21854
rect 31446 21792 31536 21820
rect 32464 21854 32554 21884
rect 32464 21820 32492 21854
rect 32526 21820 32554 21854
rect 32464 21792 32554 21820
rect 33482 21854 33572 21884
rect 33482 21820 33510 21854
rect 33544 21820 33572 21854
rect 33482 21792 33572 21820
rect 13614 21544 13704 21574
rect 13614 21510 13642 21544
rect 13676 21510 13704 21544
rect 13614 21482 13704 21510
rect 14632 21544 14722 21574
rect 14632 21510 14660 21544
rect 14694 21510 14722 21544
rect 14632 21482 14722 21510
rect 15650 21544 15740 21574
rect 15650 21510 15678 21544
rect 15712 21510 15740 21544
rect 15650 21482 15740 21510
rect 16668 21544 16758 21574
rect 16668 21510 16696 21544
rect 16730 21510 16758 21544
rect 16668 21482 16758 21510
rect 18656 21345 18672 21379
rect 19228 21345 19244 21379
rect 19674 21345 19690 21379
rect 20246 21345 20262 21379
rect 20692 21345 20708 21379
rect 21264 21345 21280 21379
rect 21710 21345 21726 21379
rect 22282 21345 22298 21379
rect 22728 21345 22744 21379
rect 23300 21345 23316 21379
rect 23746 21345 23762 21379
rect 24318 21345 24334 21379
rect 24764 21345 24780 21379
rect 25336 21345 25352 21379
rect 25782 21345 25798 21379
rect 26354 21345 26370 21379
rect 26800 21345 26816 21379
rect 27372 21345 27388 21379
rect 27818 21345 27834 21379
rect 28390 21345 28406 21379
rect 28836 21345 28852 21379
rect 29408 21345 29424 21379
rect 29854 21345 29870 21379
rect 30426 21345 30442 21379
rect 30872 21345 30888 21379
rect 31444 21345 31460 21379
rect 31890 21345 31906 21379
rect 32462 21345 32478 21379
rect 32908 21345 32924 21379
rect 33480 21345 33496 21379
rect 18424 21286 18458 21302
rect 13352 21241 13368 21275
rect 13924 21241 13940 21275
rect 14370 21241 14386 21275
rect 14942 21241 14958 21275
rect 15388 21241 15404 21275
rect 15960 21241 15976 21275
rect 16406 21241 16422 21275
rect 16978 21241 16994 21275
rect 13120 21182 13154 21198
rect 13120 20590 13154 20606
rect 14138 21182 14172 21198
rect 14138 20590 14172 20606
rect 15156 21182 15190 21198
rect 15156 20590 15190 20606
rect 16174 21182 16208 21198
rect 16174 20590 16208 20606
rect 17192 21182 17226 21198
rect 18424 20694 18458 20710
rect 19442 21286 19476 21302
rect 19442 20694 19476 20710
rect 20460 21286 20494 21302
rect 20460 20694 20494 20710
rect 21478 21286 21512 21302
rect 21478 20694 21512 20710
rect 22496 21286 22530 21302
rect 22496 20694 22530 20710
rect 23514 21286 23548 21302
rect 23514 20694 23548 20710
rect 24532 21286 24566 21302
rect 24532 20694 24566 20710
rect 25550 21286 25584 21302
rect 25550 20694 25584 20710
rect 26568 21286 26602 21302
rect 26568 20694 26602 20710
rect 27586 21286 27620 21302
rect 27586 20694 27620 20710
rect 28604 21286 28638 21302
rect 28604 20694 28638 20710
rect 29622 21286 29656 21302
rect 29622 20694 29656 20710
rect 30640 21286 30674 21302
rect 30640 20694 30674 20710
rect 31658 21286 31692 21302
rect 31658 20694 31692 20710
rect 32676 21286 32710 21302
rect 32676 20694 32710 20710
rect 33694 21286 33728 21302
rect 33694 20694 33728 20710
rect 18656 20617 18672 20651
rect 19228 20617 19244 20651
rect 19674 20617 19690 20651
rect 20246 20617 20262 20651
rect 20692 20617 20708 20651
rect 21264 20617 21280 20651
rect 21710 20617 21726 20651
rect 22282 20617 22298 20651
rect 22728 20617 22744 20651
rect 23300 20617 23316 20651
rect 23746 20617 23762 20651
rect 24318 20617 24334 20651
rect 24764 20617 24780 20651
rect 25336 20617 25352 20651
rect 25782 20617 25798 20651
rect 26354 20617 26370 20651
rect 26800 20617 26816 20651
rect 27372 20617 27388 20651
rect 27818 20617 27834 20651
rect 28390 20617 28406 20651
rect 28836 20617 28852 20651
rect 29408 20617 29424 20651
rect 29854 20617 29870 20651
rect 30426 20617 30442 20651
rect 30872 20617 30888 20651
rect 31444 20617 31460 20651
rect 31890 20617 31906 20651
rect 32462 20617 32478 20651
rect 32908 20617 32924 20651
rect 33480 20617 33496 20651
rect 17192 20590 17226 20606
rect 13352 20513 13368 20547
rect 13924 20513 13940 20547
rect 14370 20513 14386 20547
rect 14942 20513 14958 20547
rect 15388 20513 15404 20547
rect 15960 20513 15976 20547
rect 16406 20513 16422 20547
rect 16978 20513 16994 20547
rect 13090 20390 13180 20420
rect 13090 20356 13118 20390
rect 13152 20356 13180 20390
rect 13090 20328 13180 20356
rect 14108 20390 14198 20420
rect 14108 20356 14136 20390
rect 14170 20356 14198 20390
rect 14108 20328 14198 20356
rect 15126 20390 15216 20420
rect 15126 20356 15154 20390
rect 15188 20356 15216 20390
rect 15126 20328 15216 20356
rect 16144 20390 16234 20420
rect 16144 20356 16172 20390
rect 16206 20356 16234 20390
rect 16144 20328 16234 20356
rect 18302 20406 18392 20436
rect 18302 20372 18330 20406
rect 18364 20372 18392 20406
rect 18302 20344 18392 20372
rect 19320 20406 19410 20436
rect 19320 20372 19348 20406
rect 19382 20372 19410 20406
rect 19320 20344 19410 20372
rect 20338 20406 20428 20436
rect 20338 20372 20366 20406
rect 20400 20372 20428 20406
rect 20338 20344 20428 20372
rect 21356 20406 21446 20436
rect 21356 20372 21384 20406
rect 21418 20372 21446 20406
rect 21356 20344 21446 20372
rect 22374 20406 22464 20436
rect 22374 20372 22402 20406
rect 22436 20372 22464 20406
rect 22374 20344 22464 20372
rect 23392 20406 23482 20436
rect 23392 20372 23420 20406
rect 23454 20372 23482 20406
rect 23392 20344 23482 20372
rect 24410 20406 24500 20436
rect 24410 20372 24438 20406
rect 24472 20372 24500 20406
rect 24410 20344 24500 20372
rect 25428 20406 25518 20436
rect 25428 20372 25456 20406
rect 25490 20372 25518 20406
rect 25428 20344 25518 20372
rect 26446 20406 26536 20436
rect 26446 20372 26474 20406
rect 26508 20372 26536 20406
rect 26446 20344 26536 20372
rect 27464 20406 27554 20436
rect 27464 20372 27492 20406
rect 27526 20372 27554 20406
rect 27464 20344 27554 20372
rect 28482 20406 28572 20436
rect 28482 20372 28510 20406
rect 28544 20372 28572 20406
rect 28482 20344 28572 20372
rect 29500 20406 29590 20436
rect 29500 20372 29528 20406
rect 29562 20372 29590 20406
rect 29500 20344 29590 20372
rect 30518 20406 30608 20436
rect 30518 20372 30546 20406
rect 30580 20372 30608 20406
rect 30518 20344 30608 20372
rect 31536 20406 31626 20436
rect 31536 20372 31564 20406
rect 31598 20372 31626 20406
rect 31536 20344 31626 20372
rect 32554 20406 32644 20436
rect 32554 20372 32582 20406
rect 32616 20372 32644 20406
rect 32554 20344 32644 20372
rect 33572 20406 33662 20436
rect 33572 20372 33600 20406
rect 33634 20372 33662 20406
rect 33572 20344 33662 20372
rect 13352 20209 13368 20243
rect 13924 20209 13940 20243
rect 14370 20209 14386 20243
rect 14942 20209 14958 20243
rect 15388 20209 15404 20243
rect 15960 20209 15976 20243
rect 16406 20209 16422 20243
rect 16978 20209 16994 20243
rect 13120 20150 13154 20166
rect 13120 19558 13154 19574
rect 14138 20150 14172 20166
rect 14138 19558 14172 19574
rect 15156 20150 15190 20166
rect 15156 19558 15190 19574
rect 16174 20150 16208 20166
rect 16174 19558 16208 19574
rect 17192 20150 17226 20166
rect 18656 20089 18672 20123
rect 19228 20089 19244 20123
rect 19674 20089 19690 20123
rect 20246 20089 20262 20123
rect 20692 20089 20708 20123
rect 21264 20089 21280 20123
rect 21710 20089 21726 20123
rect 22282 20089 22298 20123
rect 22728 20089 22744 20123
rect 23300 20089 23316 20123
rect 23746 20089 23762 20123
rect 24318 20089 24334 20123
rect 24764 20089 24780 20123
rect 25336 20089 25352 20123
rect 25782 20089 25798 20123
rect 26354 20089 26370 20123
rect 26800 20089 26816 20123
rect 27372 20089 27388 20123
rect 27818 20089 27834 20123
rect 28390 20089 28406 20123
rect 28836 20089 28852 20123
rect 29408 20089 29424 20123
rect 29854 20089 29870 20123
rect 30426 20089 30442 20123
rect 30872 20089 30888 20123
rect 31444 20089 31460 20123
rect 31890 20089 31906 20123
rect 32462 20089 32478 20123
rect 32908 20089 32924 20123
rect 33480 20089 33496 20123
rect 17192 19558 17226 19574
rect 18424 20030 18458 20046
rect 13352 19481 13368 19515
rect 13924 19481 13940 19515
rect 14370 19481 14386 19515
rect 14942 19481 14958 19515
rect 15388 19481 15404 19515
rect 15960 19481 15976 19515
rect 16406 19481 16422 19515
rect 16978 19481 16994 19515
rect 18424 19438 18458 19454
rect 19442 20030 19476 20046
rect 19442 19438 19476 19454
rect 20460 20030 20494 20046
rect 20460 19438 20494 19454
rect 21478 20030 21512 20046
rect 21478 19438 21512 19454
rect 22496 20030 22530 20046
rect 22496 19438 22530 19454
rect 23514 20030 23548 20046
rect 23514 19438 23548 19454
rect 24532 20030 24566 20046
rect 24532 19438 24566 19454
rect 25550 20030 25584 20046
rect 25550 19438 25584 19454
rect 26568 20030 26602 20046
rect 26568 19438 26602 19454
rect 27586 20030 27620 20046
rect 27586 19438 27620 19454
rect 28604 20030 28638 20046
rect 28604 19438 28638 19454
rect 29622 20030 29656 20046
rect 29622 19438 29656 19454
rect 30640 20030 30674 20046
rect 30640 19438 30674 19454
rect 31658 20030 31692 20046
rect 31658 19438 31692 19454
rect 32676 20030 32710 20046
rect 32676 19438 32710 19454
rect 33694 20030 33728 20046
rect 33694 19438 33728 19454
rect 13100 19362 13190 19392
rect 13100 19328 13128 19362
rect 13162 19328 13190 19362
rect 13100 19300 13190 19328
rect 14118 19362 14208 19392
rect 14118 19328 14146 19362
rect 14180 19328 14208 19362
rect 14118 19300 14208 19328
rect 15136 19362 15226 19392
rect 15136 19328 15164 19362
rect 15198 19328 15226 19362
rect 15136 19300 15226 19328
rect 16154 19362 16244 19392
rect 16154 19328 16182 19362
rect 16216 19328 16244 19362
rect 18656 19361 18672 19395
rect 19228 19361 19244 19395
rect 19674 19361 19690 19395
rect 20246 19361 20262 19395
rect 20692 19361 20708 19395
rect 21264 19361 21280 19395
rect 21710 19361 21726 19395
rect 22282 19361 22298 19395
rect 22728 19361 22744 19395
rect 23300 19361 23316 19395
rect 23746 19361 23762 19395
rect 24318 19361 24334 19395
rect 24764 19361 24780 19395
rect 25336 19361 25352 19395
rect 25782 19361 25798 19395
rect 26354 19361 26370 19395
rect 26800 19361 26816 19395
rect 27372 19361 27388 19395
rect 27818 19361 27834 19395
rect 28390 19361 28406 19395
rect 28836 19361 28852 19395
rect 29408 19361 29424 19395
rect 29854 19361 29870 19395
rect 30426 19361 30442 19395
rect 30872 19361 30888 19395
rect 31444 19361 31460 19395
rect 31890 19361 31906 19395
rect 32462 19361 32478 19395
rect 32908 19361 32924 19395
rect 33480 19361 33496 19395
rect 16154 19300 16244 19328
rect 13352 19177 13368 19211
rect 13924 19177 13940 19211
rect 14370 19177 14386 19211
rect 14942 19177 14958 19211
rect 15388 19177 15404 19211
rect 15960 19177 15976 19211
rect 16406 19177 16422 19211
rect 16978 19177 16994 19211
rect 18326 19138 18416 19168
rect 13120 19118 13154 19134
rect 13120 18526 13154 18542
rect 14138 19118 14172 19134
rect 14138 18526 14172 18542
rect 15156 19118 15190 19134
rect 15156 18526 15190 18542
rect 16174 19118 16208 19134
rect 16174 18526 16208 18542
rect 17192 19118 17226 19134
rect 18326 19104 18354 19138
rect 18388 19104 18416 19138
rect 18326 19076 18416 19104
rect 19344 19138 19434 19168
rect 19344 19104 19372 19138
rect 19406 19104 19434 19138
rect 19344 19076 19434 19104
rect 20362 19138 20452 19168
rect 20362 19104 20390 19138
rect 20424 19104 20452 19138
rect 20362 19076 20452 19104
rect 21380 19138 21470 19168
rect 21380 19104 21408 19138
rect 21442 19104 21470 19138
rect 21380 19076 21470 19104
rect 22398 19138 22488 19168
rect 22398 19104 22426 19138
rect 22460 19104 22488 19138
rect 22398 19076 22488 19104
rect 23416 19138 23506 19168
rect 23416 19104 23444 19138
rect 23478 19104 23506 19138
rect 23416 19076 23506 19104
rect 24434 19138 24524 19168
rect 24434 19104 24462 19138
rect 24496 19104 24524 19138
rect 24434 19076 24524 19104
rect 25452 19138 25542 19168
rect 25452 19104 25480 19138
rect 25514 19104 25542 19138
rect 25452 19076 25542 19104
rect 26470 19138 26560 19168
rect 26470 19104 26498 19138
rect 26532 19104 26560 19138
rect 26470 19076 26560 19104
rect 27488 19138 27578 19168
rect 27488 19104 27516 19138
rect 27550 19104 27578 19138
rect 27488 19076 27578 19104
rect 28506 19138 28596 19168
rect 28506 19104 28534 19138
rect 28568 19104 28596 19138
rect 28506 19076 28596 19104
rect 29524 19138 29614 19168
rect 29524 19104 29552 19138
rect 29586 19104 29614 19138
rect 29524 19076 29614 19104
rect 30542 19138 30632 19168
rect 30542 19104 30570 19138
rect 30604 19104 30632 19138
rect 30542 19076 30632 19104
rect 31560 19138 31650 19168
rect 31560 19104 31588 19138
rect 31622 19104 31650 19138
rect 31560 19076 31650 19104
rect 32578 19138 32668 19168
rect 32578 19104 32606 19138
rect 32640 19104 32668 19138
rect 32578 19076 32668 19104
rect 33596 19138 33686 19168
rect 33596 19104 33624 19138
rect 33658 19104 33686 19138
rect 33596 19076 33686 19104
rect 18656 18833 18672 18867
rect 19228 18833 19244 18867
rect 19674 18833 19690 18867
rect 20246 18833 20262 18867
rect 20692 18833 20708 18867
rect 21264 18833 21280 18867
rect 21710 18833 21726 18867
rect 22282 18833 22298 18867
rect 22728 18833 22744 18867
rect 23300 18833 23316 18867
rect 23746 18833 23762 18867
rect 24318 18833 24334 18867
rect 24764 18833 24780 18867
rect 25336 18833 25352 18867
rect 25782 18833 25798 18867
rect 26354 18833 26370 18867
rect 26800 18833 26816 18867
rect 27372 18833 27388 18867
rect 27818 18833 27834 18867
rect 28390 18833 28406 18867
rect 28836 18833 28852 18867
rect 29408 18833 29424 18867
rect 29854 18833 29870 18867
rect 30426 18833 30442 18867
rect 30872 18833 30888 18867
rect 31444 18833 31460 18867
rect 31890 18833 31906 18867
rect 32462 18833 32478 18867
rect 32908 18833 32924 18867
rect 33480 18833 33496 18867
rect 17192 18526 17226 18542
rect 18424 18774 18458 18790
rect 13352 18449 13368 18483
rect 13924 18449 13940 18483
rect 14370 18449 14386 18483
rect 14942 18449 14958 18483
rect 15388 18449 15404 18483
rect 15960 18449 15976 18483
rect 16406 18449 16422 18483
rect 16978 18449 16994 18483
rect 13090 18334 13180 18364
rect 13090 18300 13118 18334
rect 13152 18300 13180 18334
rect 13090 18272 13180 18300
rect 14108 18334 14198 18364
rect 14108 18300 14136 18334
rect 14170 18300 14198 18334
rect 14108 18272 14198 18300
rect 15126 18334 15216 18364
rect 15126 18300 15154 18334
rect 15188 18300 15216 18334
rect 15126 18272 15216 18300
rect 16144 18334 16234 18364
rect 16144 18300 16172 18334
rect 16206 18300 16234 18334
rect 16144 18272 16234 18300
rect 18424 18182 18458 18198
rect 19442 18774 19476 18790
rect 19442 18182 19476 18198
rect 20460 18774 20494 18790
rect 20460 18182 20494 18198
rect 21478 18774 21512 18790
rect 21478 18182 21512 18198
rect 22496 18774 22530 18790
rect 22496 18182 22530 18198
rect 23514 18774 23548 18790
rect 23514 18182 23548 18198
rect 24532 18774 24566 18790
rect 24532 18182 24566 18198
rect 25550 18774 25584 18790
rect 25550 18182 25584 18198
rect 26568 18774 26602 18790
rect 26568 18182 26602 18198
rect 27586 18774 27620 18790
rect 27586 18182 27620 18198
rect 28604 18774 28638 18790
rect 28604 18182 28638 18198
rect 29622 18774 29656 18790
rect 29622 18182 29656 18198
rect 30640 18774 30674 18790
rect 30640 18182 30674 18198
rect 31658 18774 31692 18790
rect 31658 18182 31692 18198
rect 32676 18774 32710 18790
rect 32676 18182 32710 18198
rect 33694 18774 33728 18790
rect 33694 18182 33728 18198
rect 13352 18145 13368 18179
rect 13924 18145 13940 18179
rect 14370 18145 14386 18179
rect 14942 18145 14958 18179
rect 15388 18145 15404 18179
rect 15960 18145 15976 18179
rect 16406 18145 16422 18179
rect 16978 18145 16994 18179
rect 18656 18105 18672 18139
rect 19228 18105 19244 18139
rect 19674 18105 19690 18139
rect 20246 18105 20262 18139
rect 20692 18105 20708 18139
rect 21264 18105 21280 18139
rect 21710 18105 21726 18139
rect 22282 18105 22298 18139
rect 22728 18105 22744 18139
rect 23300 18105 23316 18139
rect 23746 18105 23762 18139
rect 24318 18105 24334 18139
rect 24764 18105 24780 18139
rect 25336 18105 25352 18139
rect 25782 18105 25798 18139
rect 26354 18105 26370 18139
rect 26800 18105 26816 18139
rect 27372 18105 27388 18139
rect 27818 18105 27834 18139
rect 28390 18105 28406 18139
rect 28836 18105 28852 18139
rect 29408 18105 29424 18139
rect 29854 18105 29870 18139
rect 30426 18105 30442 18139
rect 30872 18105 30888 18139
rect 31444 18105 31460 18139
rect 31890 18105 31906 18139
rect 32462 18105 32478 18139
rect 32908 18105 32924 18139
rect 33480 18105 33496 18139
rect 13120 18086 13154 18102
rect 13120 17494 13154 17510
rect 14138 18086 14172 18102
rect 14138 17494 14172 17510
rect 15156 18086 15190 18102
rect 15156 17494 15190 17510
rect 16174 18086 16208 18102
rect 16174 17494 16208 17510
rect 17192 18086 17226 18102
rect 18190 17894 18280 17924
rect 18190 17860 18218 17894
rect 18252 17860 18280 17894
rect 18190 17832 18280 17860
rect 19208 17894 19298 17924
rect 19208 17860 19236 17894
rect 19270 17860 19298 17894
rect 19208 17832 19298 17860
rect 20226 17894 20316 17924
rect 20226 17860 20254 17894
rect 20288 17860 20316 17894
rect 20226 17832 20316 17860
rect 21244 17894 21334 17924
rect 21244 17860 21272 17894
rect 21306 17860 21334 17894
rect 21244 17832 21334 17860
rect 22262 17894 22352 17924
rect 22262 17860 22290 17894
rect 22324 17860 22352 17894
rect 22262 17832 22352 17860
rect 23280 17894 23370 17924
rect 23280 17860 23308 17894
rect 23342 17860 23370 17894
rect 23280 17832 23370 17860
rect 24298 17894 24388 17924
rect 24298 17860 24326 17894
rect 24360 17860 24388 17894
rect 24298 17832 24388 17860
rect 25316 17894 25406 17924
rect 25316 17860 25344 17894
rect 25378 17860 25406 17894
rect 25316 17832 25406 17860
rect 26334 17894 26424 17924
rect 26334 17860 26362 17894
rect 26396 17860 26424 17894
rect 26334 17832 26424 17860
rect 27352 17894 27442 17924
rect 27352 17860 27380 17894
rect 27414 17860 27442 17894
rect 27352 17832 27442 17860
rect 28370 17894 28460 17924
rect 28370 17860 28398 17894
rect 28432 17860 28460 17894
rect 28370 17832 28460 17860
rect 29388 17894 29478 17924
rect 29388 17860 29416 17894
rect 29450 17860 29478 17894
rect 29388 17832 29478 17860
rect 30406 17894 30496 17924
rect 30406 17860 30434 17894
rect 30468 17860 30496 17894
rect 30406 17832 30496 17860
rect 31424 17894 31514 17924
rect 31424 17860 31452 17894
rect 31486 17860 31514 17894
rect 31424 17832 31514 17860
rect 32442 17894 32532 17924
rect 32442 17860 32470 17894
rect 32504 17860 32532 17894
rect 32442 17832 32532 17860
rect 33460 17894 33550 17924
rect 33460 17860 33488 17894
rect 33522 17860 33550 17894
rect 33460 17832 33550 17860
rect 18656 17577 18672 17611
rect 19228 17577 19244 17611
rect 19674 17577 19690 17611
rect 20246 17577 20262 17611
rect 20692 17577 20708 17611
rect 21264 17577 21280 17611
rect 21710 17577 21726 17611
rect 22282 17577 22298 17611
rect 22728 17577 22744 17611
rect 23300 17577 23316 17611
rect 23746 17577 23762 17611
rect 24318 17577 24334 17611
rect 24764 17577 24780 17611
rect 25336 17577 25352 17611
rect 25782 17577 25798 17611
rect 26354 17577 26370 17611
rect 26800 17577 26816 17611
rect 27372 17577 27388 17611
rect 27818 17577 27834 17611
rect 28390 17577 28406 17611
rect 28836 17577 28852 17611
rect 29408 17577 29424 17611
rect 29854 17577 29870 17611
rect 30426 17577 30442 17611
rect 30872 17577 30888 17611
rect 31444 17577 31460 17611
rect 31890 17577 31906 17611
rect 32462 17577 32478 17611
rect 32908 17577 32924 17611
rect 33480 17577 33496 17611
rect 17192 17494 17226 17510
rect 18424 17518 18458 17534
rect 13352 17417 13368 17451
rect 13924 17417 13940 17451
rect 14370 17417 14386 17451
rect 14942 17417 14958 17451
rect 15388 17417 15404 17451
rect 15960 17417 15976 17451
rect 16406 17417 16422 17451
rect 16978 17417 16994 17451
rect 13614 17182 13704 17212
rect 13614 17148 13642 17182
rect 13676 17148 13704 17182
rect 13614 17120 13704 17148
rect 14632 17182 14722 17212
rect 14632 17148 14660 17182
rect 14694 17148 14722 17182
rect 14632 17120 14722 17148
rect 15650 17182 15740 17212
rect 15650 17148 15678 17182
rect 15712 17148 15740 17182
rect 15650 17120 15740 17148
rect 16668 17182 16758 17212
rect 16668 17148 16696 17182
rect 16730 17148 16758 17182
rect 16668 17120 16758 17148
rect 18424 16926 18458 16942
rect 19442 17518 19476 17534
rect 19442 16926 19476 16942
rect 20460 17518 20494 17534
rect 20460 16926 20494 16942
rect 21478 17518 21512 17534
rect 21478 16926 21512 16942
rect 22496 17518 22530 17534
rect 22496 16926 22530 16942
rect 23514 17518 23548 17534
rect 23514 16926 23548 16942
rect 24532 17518 24566 17534
rect 24532 16926 24566 16942
rect 25550 17518 25584 17534
rect 25550 16926 25584 16942
rect 26568 17518 26602 17534
rect 26568 16926 26602 16942
rect 27586 17518 27620 17534
rect 27586 16926 27620 16942
rect 28604 17518 28638 17534
rect 28604 16926 28638 16942
rect 29622 17518 29656 17534
rect 29622 16926 29656 16942
rect 30640 17518 30674 17534
rect 30640 16926 30674 16942
rect 31658 17518 31692 17534
rect 31658 16926 31692 16942
rect 32676 17518 32710 17534
rect 32676 16926 32710 16942
rect 33694 17518 33728 17534
rect 33694 16926 33728 16942
rect 18656 16849 18672 16883
rect 19228 16849 19244 16883
rect 19674 16849 19690 16883
rect 20246 16849 20262 16883
rect 20692 16849 20708 16883
rect 21264 16849 21280 16883
rect 21710 16849 21726 16883
rect 22282 16849 22298 16883
rect 22728 16849 22744 16883
rect 23300 16849 23316 16883
rect 23746 16849 23762 16883
rect 24318 16849 24334 16883
rect 24764 16849 24780 16883
rect 25336 16849 25352 16883
rect 25782 16849 25798 16883
rect 26354 16849 26370 16883
rect 26800 16849 26816 16883
rect 27372 16849 27388 16883
rect 27818 16849 27834 16883
rect 28390 16849 28406 16883
rect 28836 16849 28852 16883
rect 29408 16849 29424 16883
rect 29854 16849 29870 16883
rect 30426 16849 30442 16883
rect 30872 16849 30888 16883
rect 31444 16849 31460 16883
rect 31890 16849 31906 16883
rect 32462 16849 32478 16883
rect 32908 16849 32924 16883
rect 33480 16849 33496 16883
rect 11328 16022 11428 16184
rect 35672 16022 35772 16184
rect 52328 30530 52428 30692
rect 76672 30530 76772 30692
rect 58918 28148 59008 28178
rect 58918 28114 58946 28148
rect 58980 28114 59008 28148
rect 58918 28086 59008 28114
rect 59936 28148 60026 28178
rect 59936 28114 59964 28148
rect 59998 28114 60026 28148
rect 59936 28086 60026 28114
rect 60954 28148 61044 28178
rect 60954 28114 60982 28148
rect 61016 28114 61044 28148
rect 60954 28086 61044 28114
rect 61972 28148 62062 28178
rect 61972 28114 62000 28148
rect 62034 28114 62062 28148
rect 61972 28086 62062 28114
rect 62990 28148 63080 28178
rect 62990 28114 63018 28148
rect 63052 28114 63080 28148
rect 62990 28086 63080 28114
rect 64008 28148 64098 28178
rect 64008 28114 64036 28148
rect 64070 28114 64098 28148
rect 64008 28086 64098 28114
rect 65026 28148 65116 28178
rect 65026 28114 65054 28148
rect 65088 28114 65116 28148
rect 65026 28086 65116 28114
rect 66044 28148 66134 28178
rect 66044 28114 66072 28148
rect 66106 28114 66134 28148
rect 66044 28086 66134 28114
rect 67062 28148 67152 28178
rect 67062 28114 67090 28148
rect 67124 28114 67152 28148
rect 67062 28086 67152 28114
rect 68080 28148 68170 28178
rect 68080 28114 68108 28148
rect 68142 28114 68170 28148
rect 68080 28086 68170 28114
rect 69098 28148 69188 28178
rect 69098 28114 69126 28148
rect 69160 28114 69188 28148
rect 69098 28086 69188 28114
rect 70116 28148 70206 28178
rect 70116 28114 70144 28148
rect 70178 28114 70206 28148
rect 70116 28086 70206 28114
rect 71134 28148 71224 28178
rect 71134 28114 71162 28148
rect 71196 28114 71224 28148
rect 71134 28086 71224 28114
rect 72152 28148 72242 28178
rect 72152 28114 72180 28148
rect 72214 28114 72242 28148
rect 72152 28086 72242 28114
rect 73170 28148 73260 28178
rect 73170 28114 73198 28148
rect 73232 28114 73260 28148
rect 73170 28086 73260 28114
rect 74188 28148 74278 28178
rect 74188 28114 74216 28148
rect 74250 28114 74278 28148
rect 74188 28086 74278 28114
rect 58670 27891 58686 27925
rect 59242 27891 59258 27925
rect 59688 27891 59704 27925
rect 60260 27891 60276 27925
rect 60706 27891 60722 27925
rect 61278 27891 61294 27925
rect 61724 27891 61740 27925
rect 62296 27891 62312 27925
rect 62742 27891 62758 27925
rect 63314 27891 63330 27925
rect 63760 27891 63776 27925
rect 64332 27891 64348 27925
rect 64778 27891 64794 27925
rect 65350 27891 65366 27925
rect 65796 27891 65812 27925
rect 66368 27891 66384 27925
rect 66814 27891 66830 27925
rect 67386 27891 67402 27925
rect 67832 27891 67848 27925
rect 68404 27891 68420 27925
rect 68850 27891 68866 27925
rect 69422 27891 69438 27925
rect 69868 27891 69884 27925
rect 70440 27891 70456 27925
rect 70886 27891 70902 27925
rect 71458 27891 71474 27925
rect 71904 27891 71920 27925
rect 72476 27891 72492 27925
rect 72922 27891 72938 27925
rect 73494 27891 73510 27925
rect 73940 27891 73956 27925
rect 74512 27891 74528 27925
rect 58438 27832 58472 27848
rect 58438 27240 58472 27256
rect 59456 27832 59490 27848
rect 59456 27240 59490 27256
rect 60474 27832 60508 27848
rect 60474 27240 60508 27256
rect 61492 27832 61526 27848
rect 61492 27240 61526 27256
rect 62510 27832 62544 27848
rect 62510 27240 62544 27256
rect 63528 27832 63562 27848
rect 63528 27240 63562 27256
rect 64546 27832 64580 27848
rect 64546 27240 64580 27256
rect 65564 27832 65598 27848
rect 65564 27240 65598 27256
rect 66582 27832 66616 27848
rect 66582 27240 66616 27256
rect 67600 27832 67634 27848
rect 67600 27240 67634 27256
rect 68618 27832 68652 27848
rect 68618 27240 68652 27256
rect 69636 27832 69670 27848
rect 69636 27240 69670 27256
rect 70654 27832 70688 27848
rect 70654 27240 70688 27256
rect 71672 27832 71706 27848
rect 71672 27240 71706 27256
rect 72690 27832 72724 27848
rect 72690 27240 72724 27256
rect 73708 27832 73742 27848
rect 73708 27240 73742 27256
rect 74726 27832 74760 27848
rect 74726 27240 74760 27256
rect 58670 27163 58686 27197
rect 59242 27163 59258 27197
rect 59688 27163 59704 27197
rect 60260 27163 60276 27197
rect 60706 27163 60722 27197
rect 61278 27163 61294 27197
rect 61724 27163 61740 27197
rect 62296 27163 62312 27197
rect 62742 27163 62758 27197
rect 63314 27163 63330 27197
rect 63760 27163 63776 27197
rect 64332 27163 64348 27197
rect 64778 27163 64794 27197
rect 65350 27163 65366 27197
rect 65796 27163 65812 27197
rect 66368 27163 66384 27197
rect 66814 27163 66830 27197
rect 67386 27163 67402 27197
rect 67832 27163 67848 27197
rect 68404 27163 68420 27197
rect 68850 27163 68866 27197
rect 69422 27163 69438 27197
rect 69868 27163 69884 27197
rect 70440 27163 70456 27197
rect 70886 27163 70902 27197
rect 71458 27163 71474 27197
rect 71904 27163 71920 27197
rect 72476 27163 72492 27197
rect 72922 27163 72938 27197
rect 73494 27163 73510 27197
rect 73940 27163 73956 27197
rect 74512 27163 74528 27197
rect 58940 26994 59030 27024
rect 58940 26960 58968 26994
rect 59002 26960 59030 26994
rect 58940 26932 59030 26960
rect 59958 26994 60048 27024
rect 59958 26960 59986 26994
rect 60020 26960 60048 26994
rect 59958 26932 60048 26960
rect 60976 26994 61066 27024
rect 60976 26960 61004 26994
rect 61038 26960 61066 26994
rect 60976 26932 61066 26960
rect 61994 26994 62084 27024
rect 61994 26960 62022 26994
rect 62056 26960 62084 26994
rect 61994 26932 62084 26960
rect 63012 26994 63102 27024
rect 63012 26960 63040 26994
rect 63074 26960 63102 26994
rect 63012 26932 63102 26960
rect 64030 26994 64120 27024
rect 64030 26960 64058 26994
rect 64092 26960 64120 26994
rect 64030 26932 64120 26960
rect 65048 26994 65138 27024
rect 65048 26960 65076 26994
rect 65110 26960 65138 26994
rect 65048 26932 65138 26960
rect 66066 26994 66156 27024
rect 66066 26960 66094 26994
rect 66128 26960 66156 26994
rect 66066 26932 66156 26960
rect 67084 26994 67174 27024
rect 67084 26960 67112 26994
rect 67146 26960 67174 26994
rect 67084 26932 67174 26960
rect 68102 26994 68192 27024
rect 68102 26960 68130 26994
rect 68164 26960 68192 26994
rect 68102 26932 68192 26960
rect 69120 26994 69210 27024
rect 69120 26960 69148 26994
rect 69182 26960 69210 26994
rect 69120 26932 69210 26960
rect 70138 26994 70228 27024
rect 70138 26960 70166 26994
rect 70200 26960 70228 26994
rect 70138 26932 70228 26960
rect 71156 26994 71246 27024
rect 71156 26960 71184 26994
rect 71218 26960 71246 26994
rect 71156 26932 71246 26960
rect 72174 26994 72264 27024
rect 72174 26960 72202 26994
rect 72236 26960 72264 26994
rect 72174 26932 72264 26960
rect 73192 26994 73282 27024
rect 73192 26960 73220 26994
rect 73254 26960 73282 26994
rect 73192 26932 73282 26960
rect 74210 26994 74300 27024
rect 74210 26960 74238 26994
rect 74272 26960 74300 26994
rect 74210 26932 74300 26960
rect 58670 26755 58686 26789
rect 59242 26755 59258 26789
rect 59688 26755 59704 26789
rect 60260 26755 60276 26789
rect 60706 26755 60722 26789
rect 61278 26755 61294 26789
rect 61724 26755 61740 26789
rect 62296 26755 62312 26789
rect 62742 26755 62758 26789
rect 63314 26755 63330 26789
rect 63760 26755 63776 26789
rect 64332 26755 64348 26789
rect 64778 26755 64794 26789
rect 65350 26755 65366 26789
rect 65796 26755 65812 26789
rect 66368 26755 66384 26789
rect 66814 26755 66830 26789
rect 67386 26755 67402 26789
rect 67832 26755 67848 26789
rect 68404 26755 68420 26789
rect 68850 26755 68866 26789
rect 69422 26755 69438 26789
rect 69868 26755 69884 26789
rect 70440 26755 70456 26789
rect 70886 26755 70902 26789
rect 71458 26755 71474 26789
rect 71904 26755 71920 26789
rect 72476 26755 72492 26789
rect 72922 26755 72938 26789
rect 73494 26755 73510 26789
rect 73940 26755 73956 26789
rect 74512 26755 74528 26789
rect 58438 26696 58472 26712
rect 58438 26104 58472 26120
rect 59456 26696 59490 26712
rect 59456 26104 59490 26120
rect 60474 26696 60508 26712
rect 60474 26104 60508 26120
rect 61492 26696 61526 26712
rect 61492 26104 61526 26120
rect 62510 26696 62544 26712
rect 62510 26104 62544 26120
rect 63528 26696 63562 26712
rect 63528 26104 63562 26120
rect 64546 26696 64580 26712
rect 64546 26104 64580 26120
rect 65564 26696 65598 26712
rect 65564 26104 65598 26120
rect 66582 26696 66616 26712
rect 66582 26104 66616 26120
rect 67600 26696 67634 26712
rect 67600 26104 67634 26120
rect 68618 26696 68652 26712
rect 68618 26104 68652 26120
rect 69636 26696 69670 26712
rect 69636 26104 69670 26120
rect 70654 26696 70688 26712
rect 70654 26104 70688 26120
rect 71672 26696 71706 26712
rect 71672 26104 71706 26120
rect 72690 26696 72724 26712
rect 72690 26104 72724 26120
rect 73708 26696 73742 26712
rect 73708 26104 73742 26120
rect 74726 26696 74760 26712
rect 74726 26104 74760 26120
rect 58670 26027 58686 26061
rect 59242 26027 59258 26061
rect 59688 26027 59704 26061
rect 60260 26027 60276 26061
rect 60706 26027 60722 26061
rect 61278 26027 61294 26061
rect 61724 26027 61740 26061
rect 62296 26027 62312 26061
rect 62742 26027 62758 26061
rect 63314 26027 63330 26061
rect 63760 26027 63776 26061
rect 64332 26027 64348 26061
rect 64778 26027 64794 26061
rect 65350 26027 65366 26061
rect 65796 26027 65812 26061
rect 66368 26027 66384 26061
rect 66814 26027 66830 26061
rect 67386 26027 67402 26061
rect 67832 26027 67848 26061
rect 68404 26027 68420 26061
rect 68850 26027 68866 26061
rect 69422 26027 69438 26061
rect 69868 26027 69884 26061
rect 70440 26027 70456 26061
rect 70886 26027 70902 26061
rect 71458 26027 71474 26061
rect 71904 26027 71920 26061
rect 72476 26027 72492 26061
rect 72922 26027 72938 26061
rect 73494 26027 73510 26061
rect 73940 26027 73956 26061
rect 74512 26027 74528 26061
rect 58918 25862 59008 25892
rect 58918 25828 58946 25862
rect 58980 25828 59008 25862
rect 58918 25800 59008 25828
rect 59936 25862 60026 25892
rect 59936 25828 59964 25862
rect 59998 25828 60026 25862
rect 59936 25800 60026 25828
rect 60954 25862 61044 25892
rect 60954 25828 60982 25862
rect 61016 25828 61044 25862
rect 60954 25800 61044 25828
rect 61972 25862 62062 25892
rect 61972 25828 62000 25862
rect 62034 25828 62062 25862
rect 61972 25800 62062 25828
rect 62990 25862 63080 25892
rect 62990 25828 63018 25862
rect 63052 25828 63080 25862
rect 62990 25800 63080 25828
rect 64008 25862 64098 25892
rect 64008 25828 64036 25862
rect 64070 25828 64098 25862
rect 64008 25800 64098 25828
rect 65026 25862 65116 25892
rect 65026 25828 65054 25862
rect 65088 25828 65116 25862
rect 65026 25800 65116 25828
rect 66044 25862 66134 25892
rect 66044 25828 66072 25862
rect 66106 25828 66134 25862
rect 66044 25800 66134 25828
rect 67062 25862 67152 25892
rect 67062 25828 67090 25862
rect 67124 25828 67152 25862
rect 67062 25800 67152 25828
rect 68080 25862 68170 25892
rect 68080 25828 68108 25862
rect 68142 25828 68170 25862
rect 68080 25800 68170 25828
rect 69098 25862 69188 25892
rect 69098 25828 69126 25862
rect 69160 25828 69188 25862
rect 69098 25800 69188 25828
rect 70116 25862 70206 25892
rect 70116 25828 70144 25862
rect 70178 25828 70206 25862
rect 70116 25800 70206 25828
rect 71134 25862 71224 25892
rect 71134 25828 71162 25862
rect 71196 25828 71224 25862
rect 71134 25800 71224 25828
rect 72152 25862 72242 25892
rect 72152 25828 72180 25862
rect 72214 25828 72242 25862
rect 72152 25800 72242 25828
rect 73170 25862 73260 25892
rect 73170 25828 73198 25862
rect 73232 25828 73260 25862
rect 73170 25800 73260 25828
rect 74188 25862 74278 25892
rect 74188 25828 74216 25862
rect 74250 25828 74278 25862
rect 74188 25800 74278 25828
rect 58670 25619 58686 25653
rect 59242 25619 59258 25653
rect 59688 25619 59704 25653
rect 60260 25619 60276 25653
rect 60706 25619 60722 25653
rect 61278 25619 61294 25653
rect 61724 25619 61740 25653
rect 62296 25619 62312 25653
rect 62742 25619 62758 25653
rect 63314 25619 63330 25653
rect 63760 25619 63776 25653
rect 64332 25619 64348 25653
rect 64778 25619 64794 25653
rect 65350 25619 65366 25653
rect 65796 25619 65812 25653
rect 66368 25619 66384 25653
rect 66814 25619 66830 25653
rect 67386 25619 67402 25653
rect 67832 25619 67848 25653
rect 68404 25619 68420 25653
rect 68850 25619 68866 25653
rect 69422 25619 69438 25653
rect 69868 25619 69884 25653
rect 70440 25619 70456 25653
rect 70886 25619 70902 25653
rect 71458 25619 71474 25653
rect 71904 25619 71920 25653
rect 72476 25619 72492 25653
rect 72922 25619 72938 25653
rect 73494 25619 73510 25653
rect 73940 25619 73956 25653
rect 74512 25619 74528 25653
rect 58438 25560 58472 25576
rect 58438 24968 58472 24984
rect 59456 25560 59490 25576
rect 59456 24968 59490 24984
rect 60474 25560 60508 25576
rect 60474 24968 60508 24984
rect 61492 25560 61526 25576
rect 61492 24968 61526 24984
rect 62510 25560 62544 25576
rect 62510 24968 62544 24984
rect 63528 25560 63562 25576
rect 63528 24968 63562 24984
rect 64546 25560 64580 25576
rect 64546 24968 64580 24984
rect 65564 25560 65598 25576
rect 65564 24968 65598 24984
rect 66582 25560 66616 25576
rect 66582 24968 66616 24984
rect 67600 25560 67634 25576
rect 67600 24968 67634 24984
rect 68618 25560 68652 25576
rect 68618 24968 68652 24984
rect 69636 25560 69670 25576
rect 69636 24968 69670 24984
rect 70654 25560 70688 25576
rect 70654 24968 70688 24984
rect 71672 25560 71706 25576
rect 71672 24968 71706 24984
rect 72690 25560 72724 25576
rect 72690 24968 72724 24984
rect 73708 25560 73742 25576
rect 73708 24968 73742 24984
rect 74726 25560 74760 25576
rect 74726 24968 74760 24984
rect 58670 24891 58686 24925
rect 59242 24891 59258 24925
rect 59688 24891 59704 24925
rect 60260 24891 60276 24925
rect 60706 24891 60722 24925
rect 61278 24891 61294 24925
rect 61724 24891 61740 24925
rect 62296 24891 62312 24925
rect 62742 24891 62758 24925
rect 63314 24891 63330 24925
rect 63760 24891 63776 24925
rect 64332 24891 64348 24925
rect 64778 24891 64794 24925
rect 65350 24891 65366 24925
rect 65796 24891 65812 24925
rect 66368 24891 66384 24925
rect 66814 24891 66830 24925
rect 67386 24891 67402 24925
rect 67832 24891 67848 24925
rect 68404 24891 68420 24925
rect 68850 24891 68866 24925
rect 69422 24891 69438 24925
rect 69868 24891 69884 24925
rect 70440 24891 70456 24925
rect 70886 24891 70902 24925
rect 71458 24891 71474 24925
rect 71904 24891 71920 24925
rect 72476 24891 72492 24925
rect 72922 24891 72938 24925
rect 73494 24891 73510 24925
rect 73940 24891 73956 24925
rect 74512 24891 74528 24925
rect 58918 24480 59008 24510
rect 58918 24446 58946 24480
rect 58980 24446 59008 24480
rect 58918 24418 59008 24446
rect 59936 24480 60026 24510
rect 59936 24446 59964 24480
rect 59998 24446 60026 24480
rect 59936 24418 60026 24446
rect 60954 24480 61044 24510
rect 60954 24446 60982 24480
rect 61016 24446 61044 24480
rect 60954 24418 61044 24446
rect 61972 24480 62062 24510
rect 61972 24446 62000 24480
rect 62034 24446 62062 24480
rect 61972 24418 62062 24446
rect 62990 24480 63080 24510
rect 62990 24446 63018 24480
rect 63052 24446 63080 24480
rect 62990 24418 63080 24446
rect 64008 24480 64098 24510
rect 64008 24446 64036 24480
rect 64070 24446 64098 24480
rect 64008 24418 64098 24446
rect 65026 24480 65116 24510
rect 65026 24446 65054 24480
rect 65088 24446 65116 24480
rect 65026 24418 65116 24446
rect 66044 24480 66134 24510
rect 66044 24446 66072 24480
rect 66106 24446 66134 24480
rect 66044 24418 66134 24446
rect 67062 24480 67152 24510
rect 67062 24446 67090 24480
rect 67124 24446 67152 24480
rect 67062 24418 67152 24446
rect 68080 24480 68170 24510
rect 68080 24446 68108 24480
rect 68142 24446 68170 24480
rect 68080 24418 68170 24446
rect 69098 24480 69188 24510
rect 69098 24446 69126 24480
rect 69160 24446 69188 24480
rect 69098 24418 69188 24446
rect 70116 24480 70206 24510
rect 70116 24446 70144 24480
rect 70178 24446 70206 24480
rect 70116 24418 70206 24446
rect 71134 24480 71224 24510
rect 71134 24446 71162 24480
rect 71196 24446 71224 24480
rect 71134 24418 71224 24446
rect 72152 24480 72242 24510
rect 72152 24446 72180 24480
rect 72214 24446 72242 24480
rect 72152 24418 72242 24446
rect 73170 24480 73260 24510
rect 73170 24446 73198 24480
rect 73232 24446 73260 24480
rect 73170 24418 73260 24446
rect 74188 24480 74278 24510
rect 74188 24446 74216 24480
rect 74250 24446 74278 24480
rect 74188 24418 74278 24446
rect 59864 23981 59880 24015
rect 60436 23981 60452 24015
rect 60882 23981 60898 24015
rect 61454 23981 61470 24015
rect 61900 23981 61916 24015
rect 62472 23981 62488 24015
rect 62918 23981 62934 24015
rect 63490 23981 63506 24015
rect 63936 23981 63952 24015
rect 64508 23981 64524 24015
rect 64954 23981 64970 24015
rect 65526 23981 65542 24015
rect 65972 23981 65988 24015
rect 66544 23981 66560 24015
rect 66990 23981 67006 24015
rect 67562 23981 67578 24015
rect 68008 23981 68024 24015
rect 68580 23981 68596 24015
rect 69026 23981 69042 24015
rect 69598 23981 69614 24015
rect 70044 23981 70060 24015
rect 70616 23981 70632 24015
rect 71062 23981 71078 24015
rect 71634 23981 71650 24015
rect 72080 23981 72096 24015
rect 72652 23981 72668 24015
rect 73098 23981 73114 24015
rect 73670 23981 73686 24015
rect 59632 23922 59666 23938
rect 59632 23330 59666 23346
rect 60650 23922 60684 23938
rect 60650 23330 60684 23346
rect 61668 23922 61702 23938
rect 61668 23330 61702 23346
rect 62686 23922 62720 23938
rect 62686 23330 62720 23346
rect 63704 23922 63738 23938
rect 63704 23330 63738 23346
rect 64722 23922 64756 23938
rect 64722 23330 64756 23346
rect 65740 23922 65774 23938
rect 65740 23330 65774 23346
rect 66758 23922 66792 23938
rect 66758 23330 66792 23346
rect 67776 23922 67810 23938
rect 67776 23330 67810 23346
rect 68794 23922 68828 23938
rect 68794 23330 68828 23346
rect 69812 23922 69846 23938
rect 69812 23330 69846 23346
rect 70830 23922 70864 23938
rect 70830 23330 70864 23346
rect 71848 23922 71882 23938
rect 71848 23330 71882 23346
rect 72866 23922 72900 23938
rect 72866 23330 72900 23346
rect 73884 23922 73918 23938
rect 73884 23330 73918 23346
rect 59864 23253 59880 23287
rect 60436 23253 60452 23287
rect 60882 23253 60898 23287
rect 61454 23253 61470 23287
rect 61900 23253 61916 23287
rect 62472 23253 62488 23287
rect 62918 23253 62934 23287
rect 63490 23253 63506 23287
rect 63936 23253 63952 23287
rect 64508 23253 64524 23287
rect 64954 23253 64970 23287
rect 65526 23253 65542 23287
rect 65972 23253 65988 23287
rect 66544 23253 66560 23287
rect 66990 23253 67006 23287
rect 67562 23253 67578 23287
rect 68008 23253 68024 23287
rect 68580 23253 68596 23287
rect 69026 23253 69042 23287
rect 69598 23253 69614 23287
rect 70044 23253 70060 23287
rect 70616 23253 70632 23287
rect 71062 23253 71078 23287
rect 71634 23253 71650 23287
rect 72080 23253 72096 23287
rect 72652 23253 72668 23287
rect 73098 23253 73114 23287
rect 73670 23253 73686 23287
rect 59606 23132 59696 23162
rect 59606 23098 59634 23132
rect 59668 23098 59696 23132
rect 59606 23070 59696 23098
rect 60624 23132 60714 23162
rect 60624 23098 60652 23132
rect 60686 23098 60714 23132
rect 60624 23070 60714 23098
rect 61642 23132 61732 23162
rect 61642 23098 61670 23132
rect 61704 23098 61732 23132
rect 61642 23070 61732 23098
rect 62660 23132 62750 23162
rect 62660 23098 62688 23132
rect 62722 23098 62750 23132
rect 62660 23070 62750 23098
rect 63678 23132 63768 23162
rect 63678 23098 63706 23132
rect 63740 23098 63768 23132
rect 63678 23070 63768 23098
rect 64696 23132 64786 23162
rect 64696 23098 64724 23132
rect 64758 23098 64786 23132
rect 64696 23070 64786 23098
rect 65714 23132 65804 23162
rect 65714 23098 65742 23132
rect 65776 23098 65804 23132
rect 65714 23070 65804 23098
rect 66732 23132 66822 23162
rect 66732 23098 66760 23132
rect 66794 23098 66822 23132
rect 66732 23070 66822 23098
rect 67750 23132 67840 23162
rect 67750 23098 67778 23132
rect 67812 23098 67840 23132
rect 67750 23070 67840 23098
rect 68768 23132 68858 23162
rect 68768 23098 68796 23132
rect 68830 23098 68858 23132
rect 68768 23070 68858 23098
rect 69786 23132 69876 23162
rect 69786 23098 69814 23132
rect 69848 23098 69876 23132
rect 69786 23070 69876 23098
rect 70804 23132 70894 23162
rect 70804 23098 70832 23132
rect 70866 23098 70894 23132
rect 70804 23070 70894 23098
rect 71822 23132 71912 23162
rect 71822 23098 71850 23132
rect 71884 23098 71912 23132
rect 71822 23070 71912 23098
rect 72840 23132 72930 23162
rect 72840 23098 72868 23132
rect 72902 23098 72930 23132
rect 72840 23070 72930 23098
rect 73858 23132 73948 23162
rect 73858 23098 73886 23132
rect 73920 23098 73948 23132
rect 73858 23070 73948 23098
rect 59864 22949 59880 22983
rect 60436 22949 60452 22983
rect 60882 22949 60898 22983
rect 61454 22949 61470 22983
rect 61900 22949 61916 22983
rect 62472 22949 62488 22983
rect 62918 22949 62934 22983
rect 63490 22949 63506 22983
rect 63936 22949 63952 22983
rect 64508 22949 64524 22983
rect 64954 22949 64970 22983
rect 65526 22949 65542 22983
rect 65972 22949 65988 22983
rect 66544 22949 66560 22983
rect 66990 22949 67006 22983
rect 67562 22949 67578 22983
rect 68008 22949 68024 22983
rect 68580 22949 68596 22983
rect 69026 22949 69042 22983
rect 69598 22949 69614 22983
rect 70044 22949 70060 22983
rect 70616 22949 70632 22983
rect 71062 22949 71078 22983
rect 71634 22949 71650 22983
rect 72080 22949 72096 22983
rect 72652 22949 72668 22983
rect 73098 22949 73114 22983
rect 73670 22949 73686 22983
rect 59632 22890 59666 22906
rect 59632 22298 59666 22314
rect 60650 22890 60684 22906
rect 60650 22298 60684 22314
rect 61668 22890 61702 22906
rect 61668 22298 61702 22314
rect 62686 22890 62720 22906
rect 62686 22298 62720 22314
rect 63704 22890 63738 22906
rect 63704 22298 63738 22314
rect 64722 22890 64756 22906
rect 64722 22298 64756 22314
rect 65740 22890 65774 22906
rect 65740 22298 65774 22314
rect 66758 22890 66792 22906
rect 66758 22298 66792 22314
rect 67776 22890 67810 22906
rect 67776 22298 67810 22314
rect 68794 22890 68828 22906
rect 68794 22298 68828 22314
rect 69812 22890 69846 22906
rect 69812 22298 69846 22314
rect 70830 22890 70864 22906
rect 70830 22298 70864 22314
rect 71848 22890 71882 22906
rect 71848 22298 71882 22314
rect 72866 22890 72900 22906
rect 72866 22298 72900 22314
rect 73884 22890 73918 22906
rect 73884 22298 73918 22314
rect 59864 22221 59880 22255
rect 60436 22221 60452 22255
rect 60882 22221 60898 22255
rect 61454 22221 61470 22255
rect 61900 22221 61916 22255
rect 62472 22221 62488 22255
rect 62918 22221 62934 22255
rect 63490 22221 63506 22255
rect 63936 22221 63952 22255
rect 64508 22221 64524 22255
rect 64954 22221 64970 22255
rect 65526 22221 65542 22255
rect 65972 22221 65988 22255
rect 66544 22221 66560 22255
rect 66990 22221 67006 22255
rect 67562 22221 67578 22255
rect 68008 22221 68024 22255
rect 68580 22221 68596 22255
rect 69026 22221 69042 22255
rect 69598 22221 69614 22255
rect 70044 22221 70060 22255
rect 70616 22221 70632 22255
rect 71062 22221 71078 22255
rect 71634 22221 71650 22255
rect 72080 22221 72096 22255
rect 72652 22221 72668 22255
rect 73098 22221 73114 22255
rect 73670 22221 73686 22255
rect 59212 21854 59302 21884
rect 59212 21820 59240 21854
rect 59274 21820 59302 21854
rect 59212 21792 59302 21820
rect 60230 21854 60320 21884
rect 60230 21820 60258 21854
rect 60292 21820 60320 21854
rect 60230 21792 60320 21820
rect 61248 21854 61338 21884
rect 61248 21820 61276 21854
rect 61310 21820 61338 21854
rect 61248 21792 61338 21820
rect 62266 21854 62356 21884
rect 62266 21820 62294 21854
rect 62328 21820 62356 21854
rect 62266 21792 62356 21820
rect 63284 21854 63374 21884
rect 63284 21820 63312 21854
rect 63346 21820 63374 21854
rect 63284 21792 63374 21820
rect 64302 21854 64392 21884
rect 64302 21820 64330 21854
rect 64364 21820 64392 21854
rect 64302 21792 64392 21820
rect 65320 21854 65410 21884
rect 65320 21820 65348 21854
rect 65382 21820 65410 21854
rect 65320 21792 65410 21820
rect 66338 21854 66428 21884
rect 66338 21820 66366 21854
rect 66400 21820 66428 21854
rect 66338 21792 66428 21820
rect 67356 21854 67446 21884
rect 67356 21820 67384 21854
rect 67418 21820 67446 21854
rect 67356 21792 67446 21820
rect 68374 21854 68464 21884
rect 68374 21820 68402 21854
rect 68436 21820 68464 21854
rect 68374 21792 68464 21820
rect 69392 21854 69482 21884
rect 69392 21820 69420 21854
rect 69454 21820 69482 21854
rect 69392 21792 69482 21820
rect 70410 21854 70500 21884
rect 70410 21820 70438 21854
rect 70472 21820 70500 21854
rect 70410 21792 70500 21820
rect 71428 21854 71518 21884
rect 71428 21820 71456 21854
rect 71490 21820 71518 21854
rect 71428 21792 71518 21820
rect 72446 21854 72536 21884
rect 72446 21820 72474 21854
rect 72508 21820 72536 21854
rect 72446 21792 72536 21820
rect 73464 21854 73554 21884
rect 73464 21820 73492 21854
rect 73526 21820 73554 21854
rect 73464 21792 73554 21820
rect 74482 21854 74572 21884
rect 74482 21820 74510 21854
rect 74544 21820 74572 21854
rect 74482 21792 74572 21820
rect 54614 21544 54704 21574
rect 54614 21510 54642 21544
rect 54676 21510 54704 21544
rect 54614 21482 54704 21510
rect 55632 21544 55722 21574
rect 55632 21510 55660 21544
rect 55694 21510 55722 21544
rect 55632 21482 55722 21510
rect 56650 21544 56740 21574
rect 56650 21510 56678 21544
rect 56712 21510 56740 21544
rect 56650 21482 56740 21510
rect 57668 21544 57758 21574
rect 57668 21510 57696 21544
rect 57730 21510 57758 21544
rect 57668 21482 57758 21510
rect 59656 21345 59672 21379
rect 60228 21345 60244 21379
rect 60674 21345 60690 21379
rect 61246 21345 61262 21379
rect 61692 21345 61708 21379
rect 62264 21345 62280 21379
rect 62710 21345 62726 21379
rect 63282 21345 63298 21379
rect 63728 21345 63744 21379
rect 64300 21345 64316 21379
rect 64746 21345 64762 21379
rect 65318 21345 65334 21379
rect 65764 21345 65780 21379
rect 66336 21345 66352 21379
rect 66782 21345 66798 21379
rect 67354 21345 67370 21379
rect 67800 21345 67816 21379
rect 68372 21345 68388 21379
rect 68818 21345 68834 21379
rect 69390 21345 69406 21379
rect 69836 21345 69852 21379
rect 70408 21345 70424 21379
rect 70854 21345 70870 21379
rect 71426 21345 71442 21379
rect 71872 21345 71888 21379
rect 72444 21345 72460 21379
rect 72890 21345 72906 21379
rect 73462 21345 73478 21379
rect 73908 21345 73924 21379
rect 74480 21345 74496 21379
rect 59424 21286 59458 21302
rect 54352 21241 54368 21275
rect 54924 21241 54940 21275
rect 55370 21241 55386 21275
rect 55942 21241 55958 21275
rect 56388 21241 56404 21275
rect 56960 21241 56976 21275
rect 57406 21241 57422 21275
rect 57978 21241 57994 21275
rect 54120 21182 54154 21198
rect 54120 20590 54154 20606
rect 55138 21182 55172 21198
rect 55138 20590 55172 20606
rect 56156 21182 56190 21198
rect 56156 20590 56190 20606
rect 57174 21182 57208 21198
rect 57174 20590 57208 20606
rect 58192 21182 58226 21198
rect 59424 20694 59458 20710
rect 60442 21286 60476 21302
rect 60442 20694 60476 20710
rect 61460 21286 61494 21302
rect 61460 20694 61494 20710
rect 62478 21286 62512 21302
rect 62478 20694 62512 20710
rect 63496 21286 63530 21302
rect 63496 20694 63530 20710
rect 64514 21286 64548 21302
rect 64514 20694 64548 20710
rect 65532 21286 65566 21302
rect 65532 20694 65566 20710
rect 66550 21286 66584 21302
rect 66550 20694 66584 20710
rect 67568 21286 67602 21302
rect 67568 20694 67602 20710
rect 68586 21286 68620 21302
rect 68586 20694 68620 20710
rect 69604 21286 69638 21302
rect 69604 20694 69638 20710
rect 70622 21286 70656 21302
rect 70622 20694 70656 20710
rect 71640 21286 71674 21302
rect 71640 20694 71674 20710
rect 72658 21286 72692 21302
rect 72658 20694 72692 20710
rect 73676 21286 73710 21302
rect 73676 20694 73710 20710
rect 74694 21286 74728 21302
rect 74694 20694 74728 20710
rect 59656 20617 59672 20651
rect 60228 20617 60244 20651
rect 60674 20617 60690 20651
rect 61246 20617 61262 20651
rect 61692 20617 61708 20651
rect 62264 20617 62280 20651
rect 62710 20617 62726 20651
rect 63282 20617 63298 20651
rect 63728 20617 63744 20651
rect 64300 20617 64316 20651
rect 64746 20617 64762 20651
rect 65318 20617 65334 20651
rect 65764 20617 65780 20651
rect 66336 20617 66352 20651
rect 66782 20617 66798 20651
rect 67354 20617 67370 20651
rect 67800 20617 67816 20651
rect 68372 20617 68388 20651
rect 68818 20617 68834 20651
rect 69390 20617 69406 20651
rect 69836 20617 69852 20651
rect 70408 20617 70424 20651
rect 70854 20617 70870 20651
rect 71426 20617 71442 20651
rect 71872 20617 71888 20651
rect 72444 20617 72460 20651
rect 72890 20617 72906 20651
rect 73462 20617 73478 20651
rect 73908 20617 73924 20651
rect 74480 20617 74496 20651
rect 58192 20590 58226 20606
rect 54352 20513 54368 20547
rect 54924 20513 54940 20547
rect 55370 20513 55386 20547
rect 55942 20513 55958 20547
rect 56388 20513 56404 20547
rect 56960 20513 56976 20547
rect 57406 20513 57422 20547
rect 57978 20513 57994 20547
rect 54090 20390 54180 20420
rect 54090 20356 54118 20390
rect 54152 20356 54180 20390
rect 54090 20328 54180 20356
rect 55108 20390 55198 20420
rect 55108 20356 55136 20390
rect 55170 20356 55198 20390
rect 55108 20328 55198 20356
rect 56126 20390 56216 20420
rect 56126 20356 56154 20390
rect 56188 20356 56216 20390
rect 56126 20328 56216 20356
rect 57144 20390 57234 20420
rect 57144 20356 57172 20390
rect 57206 20356 57234 20390
rect 57144 20328 57234 20356
rect 59302 20406 59392 20436
rect 59302 20372 59330 20406
rect 59364 20372 59392 20406
rect 59302 20344 59392 20372
rect 60320 20406 60410 20436
rect 60320 20372 60348 20406
rect 60382 20372 60410 20406
rect 60320 20344 60410 20372
rect 61338 20406 61428 20436
rect 61338 20372 61366 20406
rect 61400 20372 61428 20406
rect 61338 20344 61428 20372
rect 62356 20406 62446 20436
rect 62356 20372 62384 20406
rect 62418 20372 62446 20406
rect 62356 20344 62446 20372
rect 63374 20406 63464 20436
rect 63374 20372 63402 20406
rect 63436 20372 63464 20406
rect 63374 20344 63464 20372
rect 64392 20406 64482 20436
rect 64392 20372 64420 20406
rect 64454 20372 64482 20406
rect 64392 20344 64482 20372
rect 65410 20406 65500 20436
rect 65410 20372 65438 20406
rect 65472 20372 65500 20406
rect 65410 20344 65500 20372
rect 66428 20406 66518 20436
rect 66428 20372 66456 20406
rect 66490 20372 66518 20406
rect 66428 20344 66518 20372
rect 67446 20406 67536 20436
rect 67446 20372 67474 20406
rect 67508 20372 67536 20406
rect 67446 20344 67536 20372
rect 68464 20406 68554 20436
rect 68464 20372 68492 20406
rect 68526 20372 68554 20406
rect 68464 20344 68554 20372
rect 69482 20406 69572 20436
rect 69482 20372 69510 20406
rect 69544 20372 69572 20406
rect 69482 20344 69572 20372
rect 70500 20406 70590 20436
rect 70500 20372 70528 20406
rect 70562 20372 70590 20406
rect 70500 20344 70590 20372
rect 71518 20406 71608 20436
rect 71518 20372 71546 20406
rect 71580 20372 71608 20406
rect 71518 20344 71608 20372
rect 72536 20406 72626 20436
rect 72536 20372 72564 20406
rect 72598 20372 72626 20406
rect 72536 20344 72626 20372
rect 73554 20406 73644 20436
rect 73554 20372 73582 20406
rect 73616 20372 73644 20406
rect 73554 20344 73644 20372
rect 74572 20406 74662 20436
rect 74572 20372 74600 20406
rect 74634 20372 74662 20406
rect 74572 20344 74662 20372
rect 54352 20209 54368 20243
rect 54924 20209 54940 20243
rect 55370 20209 55386 20243
rect 55942 20209 55958 20243
rect 56388 20209 56404 20243
rect 56960 20209 56976 20243
rect 57406 20209 57422 20243
rect 57978 20209 57994 20243
rect 54120 20150 54154 20166
rect 54120 19558 54154 19574
rect 55138 20150 55172 20166
rect 55138 19558 55172 19574
rect 56156 20150 56190 20166
rect 56156 19558 56190 19574
rect 57174 20150 57208 20166
rect 57174 19558 57208 19574
rect 58192 20150 58226 20166
rect 59656 20089 59672 20123
rect 60228 20089 60244 20123
rect 60674 20089 60690 20123
rect 61246 20089 61262 20123
rect 61692 20089 61708 20123
rect 62264 20089 62280 20123
rect 62710 20089 62726 20123
rect 63282 20089 63298 20123
rect 63728 20089 63744 20123
rect 64300 20089 64316 20123
rect 64746 20089 64762 20123
rect 65318 20089 65334 20123
rect 65764 20089 65780 20123
rect 66336 20089 66352 20123
rect 66782 20089 66798 20123
rect 67354 20089 67370 20123
rect 67800 20089 67816 20123
rect 68372 20089 68388 20123
rect 68818 20089 68834 20123
rect 69390 20089 69406 20123
rect 69836 20089 69852 20123
rect 70408 20089 70424 20123
rect 70854 20089 70870 20123
rect 71426 20089 71442 20123
rect 71872 20089 71888 20123
rect 72444 20089 72460 20123
rect 72890 20089 72906 20123
rect 73462 20089 73478 20123
rect 73908 20089 73924 20123
rect 74480 20089 74496 20123
rect 58192 19558 58226 19574
rect 59424 20030 59458 20046
rect 54352 19481 54368 19515
rect 54924 19481 54940 19515
rect 55370 19481 55386 19515
rect 55942 19481 55958 19515
rect 56388 19481 56404 19515
rect 56960 19481 56976 19515
rect 57406 19481 57422 19515
rect 57978 19481 57994 19515
rect 59424 19438 59458 19454
rect 60442 20030 60476 20046
rect 60442 19438 60476 19454
rect 61460 20030 61494 20046
rect 61460 19438 61494 19454
rect 62478 20030 62512 20046
rect 62478 19438 62512 19454
rect 63496 20030 63530 20046
rect 63496 19438 63530 19454
rect 64514 20030 64548 20046
rect 64514 19438 64548 19454
rect 65532 20030 65566 20046
rect 65532 19438 65566 19454
rect 66550 20030 66584 20046
rect 66550 19438 66584 19454
rect 67568 20030 67602 20046
rect 67568 19438 67602 19454
rect 68586 20030 68620 20046
rect 68586 19438 68620 19454
rect 69604 20030 69638 20046
rect 69604 19438 69638 19454
rect 70622 20030 70656 20046
rect 70622 19438 70656 19454
rect 71640 20030 71674 20046
rect 71640 19438 71674 19454
rect 72658 20030 72692 20046
rect 72658 19438 72692 19454
rect 73676 20030 73710 20046
rect 73676 19438 73710 19454
rect 74694 20030 74728 20046
rect 74694 19438 74728 19454
rect 54100 19362 54190 19392
rect 54100 19328 54128 19362
rect 54162 19328 54190 19362
rect 54100 19300 54190 19328
rect 55118 19362 55208 19392
rect 55118 19328 55146 19362
rect 55180 19328 55208 19362
rect 55118 19300 55208 19328
rect 56136 19362 56226 19392
rect 56136 19328 56164 19362
rect 56198 19328 56226 19362
rect 56136 19300 56226 19328
rect 57154 19362 57244 19392
rect 57154 19328 57182 19362
rect 57216 19328 57244 19362
rect 59656 19361 59672 19395
rect 60228 19361 60244 19395
rect 60674 19361 60690 19395
rect 61246 19361 61262 19395
rect 61692 19361 61708 19395
rect 62264 19361 62280 19395
rect 62710 19361 62726 19395
rect 63282 19361 63298 19395
rect 63728 19361 63744 19395
rect 64300 19361 64316 19395
rect 64746 19361 64762 19395
rect 65318 19361 65334 19395
rect 65764 19361 65780 19395
rect 66336 19361 66352 19395
rect 66782 19361 66798 19395
rect 67354 19361 67370 19395
rect 67800 19361 67816 19395
rect 68372 19361 68388 19395
rect 68818 19361 68834 19395
rect 69390 19361 69406 19395
rect 69836 19361 69852 19395
rect 70408 19361 70424 19395
rect 70854 19361 70870 19395
rect 71426 19361 71442 19395
rect 71872 19361 71888 19395
rect 72444 19361 72460 19395
rect 72890 19361 72906 19395
rect 73462 19361 73478 19395
rect 73908 19361 73924 19395
rect 74480 19361 74496 19395
rect 57154 19300 57244 19328
rect 54352 19177 54368 19211
rect 54924 19177 54940 19211
rect 55370 19177 55386 19211
rect 55942 19177 55958 19211
rect 56388 19177 56404 19211
rect 56960 19177 56976 19211
rect 57406 19177 57422 19211
rect 57978 19177 57994 19211
rect 59326 19138 59416 19168
rect 54120 19118 54154 19134
rect 54120 18526 54154 18542
rect 55138 19118 55172 19134
rect 55138 18526 55172 18542
rect 56156 19118 56190 19134
rect 56156 18526 56190 18542
rect 57174 19118 57208 19134
rect 57174 18526 57208 18542
rect 58192 19118 58226 19134
rect 59326 19104 59354 19138
rect 59388 19104 59416 19138
rect 59326 19076 59416 19104
rect 60344 19138 60434 19168
rect 60344 19104 60372 19138
rect 60406 19104 60434 19138
rect 60344 19076 60434 19104
rect 61362 19138 61452 19168
rect 61362 19104 61390 19138
rect 61424 19104 61452 19138
rect 61362 19076 61452 19104
rect 62380 19138 62470 19168
rect 62380 19104 62408 19138
rect 62442 19104 62470 19138
rect 62380 19076 62470 19104
rect 63398 19138 63488 19168
rect 63398 19104 63426 19138
rect 63460 19104 63488 19138
rect 63398 19076 63488 19104
rect 64416 19138 64506 19168
rect 64416 19104 64444 19138
rect 64478 19104 64506 19138
rect 64416 19076 64506 19104
rect 65434 19138 65524 19168
rect 65434 19104 65462 19138
rect 65496 19104 65524 19138
rect 65434 19076 65524 19104
rect 66452 19138 66542 19168
rect 66452 19104 66480 19138
rect 66514 19104 66542 19138
rect 66452 19076 66542 19104
rect 67470 19138 67560 19168
rect 67470 19104 67498 19138
rect 67532 19104 67560 19138
rect 67470 19076 67560 19104
rect 68488 19138 68578 19168
rect 68488 19104 68516 19138
rect 68550 19104 68578 19138
rect 68488 19076 68578 19104
rect 69506 19138 69596 19168
rect 69506 19104 69534 19138
rect 69568 19104 69596 19138
rect 69506 19076 69596 19104
rect 70524 19138 70614 19168
rect 70524 19104 70552 19138
rect 70586 19104 70614 19138
rect 70524 19076 70614 19104
rect 71542 19138 71632 19168
rect 71542 19104 71570 19138
rect 71604 19104 71632 19138
rect 71542 19076 71632 19104
rect 72560 19138 72650 19168
rect 72560 19104 72588 19138
rect 72622 19104 72650 19138
rect 72560 19076 72650 19104
rect 73578 19138 73668 19168
rect 73578 19104 73606 19138
rect 73640 19104 73668 19138
rect 73578 19076 73668 19104
rect 74596 19138 74686 19168
rect 74596 19104 74624 19138
rect 74658 19104 74686 19138
rect 74596 19076 74686 19104
rect 59656 18833 59672 18867
rect 60228 18833 60244 18867
rect 60674 18833 60690 18867
rect 61246 18833 61262 18867
rect 61692 18833 61708 18867
rect 62264 18833 62280 18867
rect 62710 18833 62726 18867
rect 63282 18833 63298 18867
rect 63728 18833 63744 18867
rect 64300 18833 64316 18867
rect 64746 18833 64762 18867
rect 65318 18833 65334 18867
rect 65764 18833 65780 18867
rect 66336 18833 66352 18867
rect 66782 18833 66798 18867
rect 67354 18833 67370 18867
rect 67800 18833 67816 18867
rect 68372 18833 68388 18867
rect 68818 18833 68834 18867
rect 69390 18833 69406 18867
rect 69836 18833 69852 18867
rect 70408 18833 70424 18867
rect 70854 18833 70870 18867
rect 71426 18833 71442 18867
rect 71872 18833 71888 18867
rect 72444 18833 72460 18867
rect 72890 18833 72906 18867
rect 73462 18833 73478 18867
rect 73908 18833 73924 18867
rect 74480 18833 74496 18867
rect 58192 18526 58226 18542
rect 59424 18774 59458 18790
rect 54352 18449 54368 18483
rect 54924 18449 54940 18483
rect 55370 18449 55386 18483
rect 55942 18449 55958 18483
rect 56388 18449 56404 18483
rect 56960 18449 56976 18483
rect 57406 18449 57422 18483
rect 57978 18449 57994 18483
rect 54090 18334 54180 18364
rect 54090 18300 54118 18334
rect 54152 18300 54180 18334
rect 54090 18272 54180 18300
rect 55108 18334 55198 18364
rect 55108 18300 55136 18334
rect 55170 18300 55198 18334
rect 55108 18272 55198 18300
rect 56126 18334 56216 18364
rect 56126 18300 56154 18334
rect 56188 18300 56216 18334
rect 56126 18272 56216 18300
rect 57144 18334 57234 18364
rect 57144 18300 57172 18334
rect 57206 18300 57234 18334
rect 57144 18272 57234 18300
rect 59424 18182 59458 18198
rect 60442 18774 60476 18790
rect 60442 18182 60476 18198
rect 61460 18774 61494 18790
rect 61460 18182 61494 18198
rect 62478 18774 62512 18790
rect 62478 18182 62512 18198
rect 63496 18774 63530 18790
rect 63496 18182 63530 18198
rect 64514 18774 64548 18790
rect 64514 18182 64548 18198
rect 65532 18774 65566 18790
rect 65532 18182 65566 18198
rect 66550 18774 66584 18790
rect 66550 18182 66584 18198
rect 67568 18774 67602 18790
rect 67568 18182 67602 18198
rect 68586 18774 68620 18790
rect 68586 18182 68620 18198
rect 69604 18774 69638 18790
rect 69604 18182 69638 18198
rect 70622 18774 70656 18790
rect 70622 18182 70656 18198
rect 71640 18774 71674 18790
rect 71640 18182 71674 18198
rect 72658 18774 72692 18790
rect 72658 18182 72692 18198
rect 73676 18774 73710 18790
rect 73676 18182 73710 18198
rect 74694 18774 74728 18790
rect 74694 18182 74728 18198
rect 54352 18145 54368 18179
rect 54924 18145 54940 18179
rect 55370 18145 55386 18179
rect 55942 18145 55958 18179
rect 56388 18145 56404 18179
rect 56960 18145 56976 18179
rect 57406 18145 57422 18179
rect 57978 18145 57994 18179
rect 59656 18105 59672 18139
rect 60228 18105 60244 18139
rect 60674 18105 60690 18139
rect 61246 18105 61262 18139
rect 61692 18105 61708 18139
rect 62264 18105 62280 18139
rect 62710 18105 62726 18139
rect 63282 18105 63298 18139
rect 63728 18105 63744 18139
rect 64300 18105 64316 18139
rect 64746 18105 64762 18139
rect 65318 18105 65334 18139
rect 65764 18105 65780 18139
rect 66336 18105 66352 18139
rect 66782 18105 66798 18139
rect 67354 18105 67370 18139
rect 67800 18105 67816 18139
rect 68372 18105 68388 18139
rect 68818 18105 68834 18139
rect 69390 18105 69406 18139
rect 69836 18105 69852 18139
rect 70408 18105 70424 18139
rect 70854 18105 70870 18139
rect 71426 18105 71442 18139
rect 71872 18105 71888 18139
rect 72444 18105 72460 18139
rect 72890 18105 72906 18139
rect 73462 18105 73478 18139
rect 73908 18105 73924 18139
rect 74480 18105 74496 18139
rect 54120 18086 54154 18102
rect 54120 17494 54154 17510
rect 55138 18086 55172 18102
rect 55138 17494 55172 17510
rect 56156 18086 56190 18102
rect 56156 17494 56190 17510
rect 57174 18086 57208 18102
rect 57174 17494 57208 17510
rect 58192 18086 58226 18102
rect 59190 17894 59280 17924
rect 59190 17860 59218 17894
rect 59252 17860 59280 17894
rect 59190 17832 59280 17860
rect 60208 17894 60298 17924
rect 60208 17860 60236 17894
rect 60270 17860 60298 17894
rect 60208 17832 60298 17860
rect 61226 17894 61316 17924
rect 61226 17860 61254 17894
rect 61288 17860 61316 17894
rect 61226 17832 61316 17860
rect 62244 17894 62334 17924
rect 62244 17860 62272 17894
rect 62306 17860 62334 17894
rect 62244 17832 62334 17860
rect 63262 17894 63352 17924
rect 63262 17860 63290 17894
rect 63324 17860 63352 17894
rect 63262 17832 63352 17860
rect 64280 17894 64370 17924
rect 64280 17860 64308 17894
rect 64342 17860 64370 17894
rect 64280 17832 64370 17860
rect 65298 17894 65388 17924
rect 65298 17860 65326 17894
rect 65360 17860 65388 17894
rect 65298 17832 65388 17860
rect 66316 17894 66406 17924
rect 66316 17860 66344 17894
rect 66378 17860 66406 17894
rect 66316 17832 66406 17860
rect 67334 17894 67424 17924
rect 67334 17860 67362 17894
rect 67396 17860 67424 17894
rect 67334 17832 67424 17860
rect 68352 17894 68442 17924
rect 68352 17860 68380 17894
rect 68414 17860 68442 17894
rect 68352 17832 68442 17860
rect 69370 17894 69460 17924
rect 69370 17860 69398 17894
rect 69432 17860 69460 17894
rect 69370 17832 69460 17860
rect 70388 17894 70478 17924
rect 70388 17860 70416 17894
rect 70450 17860 70478 17894
rect 70388 17832 70478 17860
rect 71406 17894 71496 17924
rect 71406 17860 71434 17894
rect 71468 17860 71496 17894
rect 71406 17832 71496 17860
rect 72424 17894 72514 17924
rect 72424 17860 72452 17894
rect 72486 17860 72514 17894
rect 72424 17832 72514 17860
rect 73442 17894 73532 17924
rect 73442 17860 73470 17894
rect 73504 17860 73532 17894
rect 73442 17832 73532 17860
rect 74460 17894 74550 17924
rect 74460 17860 74488 17894
rect 74522 17860 74550 17894
rect 74460 17832 74550 17860
rect 59656 17577 59672 17611
rect 60228 17577 60244 17611
rect 60674 17577 60690 17611
rect 61246 17577 61262 17611
rect 61692 17577 61708 17611
rect 62264 17577 62280 17611
rect 62710 17577 62726 17611
rect 63282 17577 63298 17611
rect 63728 17577 63744 17611
rect 64300 17577 64316 17611
rect 64746 17577 64762 17611
rect 65318 17577 65334 17611
rect 65764 17577 65780 17611
rect 66336 17577 66352 17611
rect 66782 17577 66798 17611
rect 67354 17577 67370 17611
rect 67800 17577 67816 17611
rect 68372 17577 68388 17611
rect 68818 17577 68834 17611
rect 69390 17577 69406 17611
rect 69836 17577 69852 17611
rect 70408 17577 70424 17611
rect 70854 17577 70870 17611
rect 71426 17577 71442 17611
rect 71872 17577 71888 17611
rect 72444 17577 72460 17611
rect 72890 17577 72906 17611
rect 73462 17577 73478 17611
rect 73908 17577 73924 17611
rect 74480 17577 74496 17611
rect 58192 17494 58226 17510
rect 59424 17518 59458 17534
rect 54352 17417 54368 17451
rect 54924 17417 54940 17451
rect 55370 17417 55386 17451
rect 55942 17417 55958 17451
rect 56388 17417 56404 17451
rect 56960 17417 56976 17451
rect 57406 17417 57422 17451
rect 57978 17417 57994 17451
rect 54614 17182 54704 17212
rect 54614 17148 54642 17182
rect 54676 17148 54704 17182
rect 54614 17120 54704 17148
rect 55632 17182 55722 17212
rect 55632 17148 55660 17182
rect 55694 17148 55722 17182
rect 55632 17120 55722 17148
rect 56650 17182 56740 17212
rect 56650 17148 56678 17182
rect 56712 17148 56740 17182
rect 56650 17120 56740 17148
rect 57668 17182 57758 17212
rect 57668 17148 57696 17182
rect 57730 17148 57758 17182
rect 57668 17120 57758 17148
rect 59424 16926 59458 16942
rect 60442 17518 60476 17534
rect 60442 16926 60476 16942
rect 61460 17518 61494 17534
rect 61460 16926 61494 16942
rect 62478 17518 62512 17534
rect 62478 16926 62512 16942
rect 63496 17518 63530 17534
rect 63496 16926 63530 16942
rect 64514 17518 64548 17534
rect 64514 16926 64548 16942
rect 65532 17518 65566 17534
rect 65532 16926 65566 16942
rect 66550 17518 66584 17534
rect 66550 16926 66584 16942
rect 67568 17518 67602 17534
rect 67568 16926 67602 16942
rect 68586 17518 68620 17534
rect 68586 16926 68620 16942
rect 69604 17518 69638 17534
rect 69604 16926 69638 16942
rect 70622 17518 70656 17534
rect 70622 16926 70656 16942
rect 71640 17518 71674 17534
rect 71640 16926 71674 16942
rect 72658 17518 72692 17534
rect 72658 16926 72692 16942
rect 73676 17518 73710 17534
rect 73676 16926 73710 16942
rect 74694 17518 74728 17534
rect 74694 16926 74728 16942
rect 59656 16849 59672 16883
rect 60228 16849 60244 16883
rect 60674 16849 60690 16883
rect 61246 16849 61262 16883
rect 61692 16849 61708 16883
rect 62264 16849 62280 16883
rect 62710 16849 62726 16883
rect 63282 16849 63298 16883
rect 63728 16849 63744 16883
rect 64300 16849 64316 16883
rect 64746 16849 64762 16883
rect 65318 16849 65334 16883
rect 65764 16849 65780 16883
rect 66336 16849 66352 16883
rect 66782 16849 66798 16883
rect 67354 16849 67370 16883
rect 67800 16849 67816 16883
rect 68372 16849 68388 16883
rect 68818 16849 68834 16883
rect 69390 16849 69406 16883
rect 69836 16849 69852 16883
rect 70408 16849 70424 16883
rect 70854 16849 70870 16883
rect 71426 16849 71442 16883
rect 71872 16849 71888 16883
rect 72444 16849 72460 16883
rect 72890 16849 72906 16883
rect 73462 16849 73478 16883
rect 73908 16849 73924 16883
rect 74480 16849 74496 16883
rect 52328 16022 52428 16184
rect 76672 16022 76772 16184
rect -1372 15030 -1272 15192
rect 35772 15030 35872 15192
rect 14036 14586 14118 14610
rect 14036 14552 14060 14586
rect 14094 14552 14118 14586
rect 14036 14528 14118 14552
rect 15054 14586 15136 14610
rect 15054 14552 15078 14586
rect 15112 14552 15136 14586
rect 15054 14528 15136 14552
rect 16072 14586 16154 14610
rect 16072 14552 16096 14586
rect 16130 14552 16154 14586
rect 16072 14528 16154 14552
rect 17090 14586 17172 14610
rect 17090 14552 17114 14586
rect 17148 14552 17172 14586
rect 17090 14528 17172 14552
rect 18108 14586 18190 14610
rect 18108 14552 18132 14586
rect 18166 14552 18190 14586
rect 18108 14528 18190 14552
rect 19126 14586 19208 14610
rect 19126 14552 19150 14586
rect 19184 14552 19208 14586
rect 19126 14528 19208 14552
rect 20144 14586 20226 14610
rect 20144 14552 20168 14586
rect 20202 14552 20226 14586
rect 20144 14528 20226 14552
rect 21162 14586 21244 14610
rect 21162 14552 21186 14586
rect 21220 14552 21244 14586
rect 21162 14528 21244 14552
rect 22180 14586 22262 14610
rect 22180 14552 22204 14586
rect 22238 14552 22262 14586
rect 22180 14528 22262 14552
rect 23198 14586 23280 14610
rect 23198 14552 23222 14586
rect 23256 14552 23280 14586
rect 23198 14528 23280 14552
rect 24216 14586 24298 14610
rect 24216 14552 24240 14586
rect 24274 14552 24298 14586
rect 24216 14528 24298 14552
rect 25234 14586 25316 14610
rect 25234 14552 25258 14586
rect 25292 14552 25316 14586
rect 25234 14528 25316 14552
rect 26252 14586 26334 14610
rect 26252 14552 26276 14586
rect 26310 14552 26334 14586
rect 26252 14528 26334 14552
rect 27270 14586 27352 14610
rect 27270 14552 27294 14586
rect 27328 14552 27352 14586
rect 27270 14528 27352 14552
rect 28288 14586 28370 14610
rect 28288 14552 28312 14586
rect 28346 14552 28370 14586
rect 28288 14528 28370 14552
rect 29306 14586 29388 14610
rect 29306 14552 29330 14586
rect 29364 14552 29388 14586
rect 29306 14528 29388 14552
rect 30324 14586 30406 14610
rect 30324 14552 30348 14586
rect 30382 14552 30406 14586
rect 30324 14528 30406 14552
rect 31342 14586 31424 14610
rect 31342 14552 31366 14586
rect 31400 14552 31424 14586
rect 31342 14528 31424 14552
rect 32360 14586 32442 14610
rect 32360 14552 32384 14586
rect 32418 14552 32442 14586
rect 32360 14528 32442 14552
rect 33378 14586 33460 14610
rect 33378 14552 33402 14586
rect 33436 14552 33460 14586
rect 33378 14528 33460 14552
rect 13764 14372 13780 14406
rect 14336 14372 14352 14406
rect 14782 14372 14798 14406
rect 15354 14372 15370 14406
rect 15800 14372 15816 14406
rect 16372 14372 16388 14406
rect 16818 14372 16834 14406
rect 17390 14372 17406 14406
rect 17836 14372 17852 14406
rect 18408 14372 18424 14406
rect 18854 14372 18870 14406
rect 19426 14372 19442 14406
rect 19872 14372 19888 14406
rect 20444 14372 20460 14406
rect 20890 14372 20906 14406
rect 21462 14372 21478 14406
rect 21908 14372 21924 14406
rect 22480 14372 22496 14406
rect 22926 14372 22942 14406
rect 23498 14372 23514 14406
rect 23944 14372 23960 14406
rect 24516 14372 24532 14406
rect 24962 14372 24978 14406
rect 25534 14372 25550 14406
rect 25980 14372 25996 14406
rect 26552 14372 26568 14406
rect 26998 14372 27014 14406
rect 27570 14372 27586 14406
rect 28016 14372 28032 14406
rect 28588 14372 28604 14406
rect 29034 14372 29050 14406
rect 29606 14372 29622 14406
rect 30052 14372 30068 14406
rect 30624 14372 30640 14406
rect 31070 14372 31086 14406
rect 31642 14372 31658 14406
rect 32088 14372 32104 14406
rect 32660 14372 32676 14406
rect 33106 14372 33122 14406
rect 33678 14372 33694 14406
rect 13532 14322 13566 14338
rect 1742 13984 1824 14008
rect 1742 13950 1766 13984
rect 1800 13950 1824 13984
rect 1742 13926 1824 13950
rect 2760 13984 2842 14008
rect 2760 13950 2784 13984
rect 2818 13950 2842 13984
rect 1998 13896 2014 13930
rect 2570 13896 2586 13930
rect 2760 13926 2842 13950
rect 3778 13984 3860 14008
rect 3778 13950 3802 13984
rect 3836 13950 3860 13984
rect 3016 13896 3032 13930
rect 3588 13896 3604 13930
rect 3778 13926 3860 13950
rect 4796 13984 4878 14008
rect 4796 13950 4820 13984
rect 4854 13950 4878 13984
rect 4034 13896 4050 13930
rect 4606 13896 4622 13930
rect 4796 13926 4878 13950
rect 5814 13984 5896 14008
rect 5814 13950 5838 13984
rect 5872 13950 5896 13984
rect 5052 13896 5068 13930
rect 5624 13896 5640 13930
rect 5814 13926 5896 13950
rect 6832 13984 6914 14008
rect 6832 13950 6856 13984
rect 6890 13950 6914 13984
rect 6070 13896 6086 13930
rect 6642 13896 6658 13930
rect 6832 13926 6914 13950
rect 7850 13984 7932 14008
rect 7850 13950 7874 13984
rect 7908 13950 7932 13984
rect 7088 13896 7104 13930
rect 7660 13896 7676 13930
rect 7850 13926 7932 13950
rect 8868 13984 8950 14008
rect 8868 13950 8892 13984
rect 8926 13950 8950 13984
rect 8106 13896 8122 13930
rect 8678 13896 8694 13930
rect 8868 13926 8950 13950
rect 9886 13984 9968 14008
rect 9886 13950 9910 13984
rect 9944 13950 9968 13984
rect 9124 13896 9140 13930
rect 9696 13896 9712 13930
rect 9886 13926 9968 13950
rect 10914 13984 10996 14008
rect 10914 13950 10938 13984
rect 10972 13950 10996 13984
rect 10142 13896 10158 13930
rect 10714 13896 10730 13930
rect 10914 13926 10996 13950
rect 1766 13846 1800 13862
rect 1766 13254 1800 13270
rect 2784 13846 2818 13862
rect 2784 13254 2818 13270
rect 3802 13846 3836 13862
rect 3802 13254 3836 13270
rect 4820 13846 4854 13862
rect 4820 13254 4854 13270
rect 5838 13846 5872 13862
rect 5838 13254 5872 13270
rect 6856 13846 6890 13862
rect 6856 13254 6890 13270
rect 7874 13846 7908 13862
rect 7874 13254 7908 13270
rect 8892 13846 8926 13862
rect 8892 13254 8926 13270
rect 9910 13846 9944 13862
rect 9910 13254 9944 13270
rect 10928 13846 10962 13862
rect 13532 13730 13566 13746
rect 14550 14322 14584 14338
rect 14550 13730 14584 13746
rect 15568 14322 15602 14338
rect 15568 13730 15602 13746
rect 16586 14322 16620 14338
rect 16586 13730 16620 13746
rect 17604 14322 17638 14338
rect 17604 13730 17638 13746
rect 18622 14322 18656 14338
rect 18622 13730 18656 13746
rect 19640 14322 19674 14338
rect 19640 13730 19674 13746
rect 20658 14322 20692 14338
rect 20658 13730 20692 13746
rect 21676 14322 21710 14338
rect 21676 13730 21710 13746
rect 22694 14322 22728 14338
rect 22694 13730 22728 13746
rect 23712 14322 23746 14338
rect 23712 13730 23746 13746
rect 24730 14322 24764 14338
rect 24730 13730 24764 13746
rect 25748 14322 25782 14338
rect 25748 13730 25782 13746
rect 26766 14322 26800 14338
rect 26766 13730 26800 13746
rect 27784 14322 27818 14338
rect 27784 13730 27818 13746
rect 28802 14322 28836 14338
rect 28802 13730 28836 13746
rect 29820 14322 29854 14338
rect 29820 13730 29854 13746
rect 30838 14322 30872 14338
rect 30838 13730 30872 13746
rect 31856 14322 31890 14338
rect 31856 13730 31890 13746
rect 32874 14322 32908 14338
rect 32874 13730 32908 13746
rect 33892 14322 33926 14338
rect 33892 13730 33926 13746
rect 13764 13662 13780 13696
rect 14336 13662 14352 13696
rect 14782 13662 14798 13696
rect 15354 13662 15370 13696
rect 15800 13662 15816 13696
rect 16372 13662 16388 13696
rect 16818 13662 16834 13696
rect 17390 13662 17406 13696
rect 17836 13662 17852 13696
rect 18408 13662 18424 13696
rect 18854 13662 18870 13696
rect 19426 13662 19442 13696
rect 19872 13662 19888 13696
rect 20444 13662 20460 13696
rect 20890 13662 20906 13696
rect 21462 13662 21478 13696
rect 21908 13662 21924 13696
rect 22480 13662 22496 13696
rect 22926 13662 22942 13696
rect 23498 13662 23514 13696
rect 23944 13662 23960 13696
rect 24516 13662 24532 13696
rect 24962 13662 24978 13696
rect 25534 13662 25550 13696
rect 25980 13662 25996 13696
rect 26552 13662 26568 13696
rect 26998 13662 27014 13696
rect 27570 13662 27586 13696
rect 28016 13662 28032 13696
rect 28588 13662 28604 13696
rect 29034 13662 29050 13696
rect 29606 13662 29622 13696
rect 30052 13662 30068 13696
rect 30624 13662 30640 13696
rect 31070 13662 31086 13696
rect 31642 13662 31658 13696
rect 32088 13662 32104 13696
rect 32660 13662 32676 13696
rect 33106 13662 33122 13696
rect 33678 13662 33694 13696
rect 13764 13554 13780 13588
rect 14336 13554 14352 13588
rect 14782 13554 14798 13588
rect 15354 13554 15370 13588
rect 15800 13554 15816 13588
rect 16372 13554 16388 13588
rect 16818 13554 16834 13588
rect 17390 13554 17406 13588
rect 17836 13554 17852 13588
rect 18408 13554 18424 13588
rect 18854 13554 18870 13588
rect 19426 13554 19442 13588
rect 19872 13554 19888 13588
rect 20444 13554 20460 13588
rect 20890 13554 20906 13588
rect 21462 13554 21478 13588
rect 21908 13554 21924 13588
rect 22480 13554 22496 13588
rect 22926 13554 22942 13588
rect 23498 13554 23514 13588
rect 23944 13554 23960 13588
rect 24516 13554 24532 13588
rect 24962 13554 24978 13588
rect 25534 13554 25550 13588
rect 25980 13554 25996 13588
rect 26552 13554 26568 13588
rect 26998 13554 27014 13588
rect 27570 13554 27586 13588
rect 28016 13554 28032 13588
rect 28588 13554 28604 13588
rect 29034 13554 29050 13588
rect 29606 13554 29622 13588
rect 30052 13554 30068 13588
rect 30624 13554 30640 13588
rect 31070 13554 31086 13588
rect 31642 13554 31658 13588
rect 32088 13554 32104 13588
rect 32660 13554 32676 13588
rect 33106 13554 33122 13588
rect 33678 13554 33694 13588
rect 10928 13254 10962 13270
rect 13532 13504 13566 13520
rect 1742 13166 1824 13190
rect 1998 13186 2014 13220
rect 2570 13186 2586 13220
rect 1742 13132 1766 13166
rect 1800 13132 1824 13166
rect 1742 13108 1824 13132
rect 2760 13166 2842 13190
rect 3016 13186 3032 13220
rect 3588 13186 3604 13220
rect 2760 13132 2784 13166
rect 2818 13132 2842 13166
rect 1998 13078 2014 13112
rect 2570 13078 2586 13112
rect 2760 13108 2842 13132
rect 3778 13166 3860 13190
rect 4034 13186 4050 13220
rect 4606 13186 4622 13220
rect 3778 13132 3802 13166
rect 3836 13132 3860 13166
rect 3016 13078 3032 13112
rect 3588 13078 3604 13112
rect 3778 13108 3860 13132
rect 4796 13166 4878 13190
rect 5052 13186 5068 13220
rect 5624 13186 5640 13220
rect 4796 13132 4820 13166
rect 4854 13132 4878 13166
rect 4034 13078 4050 13112
rect 4606 13078 4622 13112
rect 4796 13108 4878 13132
rect 5814 13166 5896 13190
rect 6070 13186 6086 13220
rect 6642 13186 6658 13220
rect 5814 13132 5838 13166
rect 5872 13132 5896 13166
rect 5052 13078 5068 13112
rect 5624 13078 5640 13112
rect 5814 13108 5896 13132
rect 6832 13166 6914 13190
rect 7088 13186 7104 13220
rect 7660 13186 7676 13220
rect 6832 13132 6856 13166
rect 6890 13132 6914 13166
rect 6070 13078 6086 13112
rect 6642 13078 6658 13112
rect 6832 13108 6914 13132
rect 7850 13166 7932 13190
rect 8106 13186 8122 13220
rect 8678 13186 8694 13220
rect 7850 13132 7874 13166
rect 7908 13132 7932 13166
rect 7088 13078 7104 13112
rect 7660 13078 7676 13112
rect 7850 13108 7932 13132
rect 8868 13166 8950 13190
rect 9124 13186 9140 13220
rect 9696 13186 9712 13220
rect 8868 13132 8892 13166
rect 8926 13132 8950 13166
rect 8106 13078 8122 13112
rect 8678 13078 8694 13112
rect 8868 13108 8950 13132
rect 9886 13166 9968 13190
rect 10142 13186 10158 13220
rect 10714 13186 10730 13220
rect 9886 13132 9910 13166
rect 9944 13132 9968 13166
rect 9124 13078 9140 13112
rect 9696 13078 9712 13112
rect 9886 13108 9968 13132
rect 10914 13166 10996 13190
rect 10914 13132 10938 13166
rect 10972 13132 10996 13166
rect 10142 13078 10158 13112
rect 10714 13078 10730 13112
rect 10914 13108 10996 13132
rect 7358 13076 7418 13078
rect 1766 13028 1800 13044
rect 1766 12436 1800 12452
rect 2784 13028 2818 13044
rect 2784 12436 2818 12452
rect 3802 13028 3836 13044
rect 3802 12436 3836 12452
rect 4820 13028 4854 13044
rect 4820 12436 4854 12452
rect 5838 13028 5872 13044
rect 5838 12436 5872 12452
rect 6856 13028 6890 13044
rect 6856 12436 6890 12452
rect 7874 13028 7908 13044
rect 7874 12436 7908 12452
rect 8892 13028 8926 13044
rect 8892 12436 8926 12452
rect 9910 13028 9944 13044
rect 9910 12436 9944 12452
rect 10928 13028 10962 13044
rect 13532 12912 13566 12928
rect 14550 13504 14584 13520
rect 14550 12912 14584 12928
rect 15568 13504 15602 13520
rect 15568 12912 15602 12928
rect 16586 13504 16620 13520
rect 16586 12912 16620 12928
rect 17604 13504 17638 13520
rect 17604 12912 17638 12928
rect 18622 13504 18656 13520
rect 18622 12912 18656 12928
rect 19640 13504 19674 13520
rect 19640 12912 19674 12928
rect 20658 13504 20692 13520
rect 20658 12912 20692 12928
rect 21676 13504 21710 13520
rect 21676 12912 21710 12928
rect 22694 13504 22728 13520
rect 22694 12912 22728 12928
rect 23712 13504 23746 13520
rect 23712 12912 23746 12928
rect 24730 13504 24764 13520
rect 24730 12912 24764 12928
rect 25748 13504 25782 13520
rect 25748 12912 25782 12928
rect 26766 13504 26800 13520
rect 26766 12912 26800 12928
rect 27784 13504 27818 13520
rect 27784 12912 27818 12928
rect 28802 13504 28836 13520
rect 28802 12912 28836 12928
rect 29820 13504 29854 13520
rect 29820 12912 29854 12928
rect 30838 13504 30872 13520
rect 30838 12912 30872 12928
rect 31856 13504 31890 13520
rect 31856 12912 31890 12928
rect 32874 13504 32908 13520
rect 32874 12912 32908 12928
rect 33892 13504 33926 13520
rect 33892 12912 33926 12928
rect 13764 12844 13780 12878
rect 14336 12844 14352 12878
rect 14782 12844 14798 12878
rect 15354 12844 15370 12878
rect 15800 12844 15816 12878
rect 16372 12844 16388 12878
rect 16818 12844 16834 12878
rect 17390 12844 17406 12878
rect 17836 12844 17852 12878
rect 18408 12844 18424 12878
rect 18854 12844 18870 12878
rect 19426 12844 19442 12878
rect 19872 12844 19888 12878
rect 20444 12844 20460 12878
rect 20890 12844 20906 12878
rect 21462 12844 21478 12878
rect 21908 12844 21924 12878
rect 22480 12844 22496 12878
rect 22926 12844 22942 12878
rect 23498 12844 23514 12878
rect 23944 12844 23960 12878
rect 24516 12844 24532 12878
rect 24962 12844 24978 12878
rect 25534 12844 25550 12878
rect 25980 12844 25996 12878
rect 26552 12844 26568 12878
rect 26998 12844 27014 12878
rect 27570 12844 27586 12878
rect 28016 12844 28032 12878
rect 28588 12844 28604 12878
rect 29034 12844 29050 12878
rect 29606 12844 29622 12878
rect 30052 12844 30068 12878
rect 30624 12844 30640 12878
rect 31070 12844 31086 12878
rect 31642 12844 31658 12878
rect 32088 12844 32104 12878
rect 32660 12844 32676 12878
rect 33106 12844 33122 12878
rect 33678 12844 33694 12878
rect 14048 12560 14130 12584
rect 14048 12526 14072 12560
rect 14106 12526 14130 12560
rect 14048 12502 14130 12526
rect 15066 12560 15148 12584
rect 15066 12526 15090 12560
rect 15124 12526 15148 12560
rect 15066 12502 15148 12526
rect 16084 12560 16166 12584
rect 16084 12526 16108 12560
rect 16142 12526 16166 12560
rect 16084 12502 16166 12526
rect 17102 12560 17184 12584
rect 17102 12526 17126 12560
rect 17160 12526 17184 12560
rect 17102 12502 17184 12526
rect 18120 12560 18202 12584
rect 18120 12526 18144 12560
rect 18178 12526 18202 12560
rect 18120 12502 18202 12526
rect 19138 12560 19220 12584
rect 19138 12526 19162 12560
rect 19196 12526 19220 12560
rect 19138 12502 19220 12526
rect 20156 12560 20238 12584
rect 20156 12526 20180 12560
rect 20214 12526 20238 12560
rect 20156 12502 20238 12526
rect 21174 12560 21256 12584
rect 21174 12526 21198 12560
rect 21232 12526 21256 12560
rect 21174 12502 21256 12526
rect 22192 12560 22274 12584
rect 22192 12526 22216 12560
rect 22250 12526 22274 12560
rect 22192 12502 22274 12526
rect 23210 12560 23292 12584
rect 23210 12526 23234 12560
rect 23268 12526 23292 12560
rect 23210 12502 23292 12526
rect 24228 12560 24310 12584
rect 24228 12526 24252 12560
rect 24286 12526 24310 12560
rect 24228 12502 24310 12526
rect 25246 12560 25328 12584
rect 25246 12526 25270 12560
rect 25304 12526 25328 12560
rect 25246 12502 25328 12526
rect 26264 12560 26346 12584
rect 26264 12526 26288 12560
rect 26322 12526 26346 12560
rect 26264 12502 26346 12526
rect 27282 12560 27364 12584
rect 27282 12526 27306 12560
rect 27340 12526 27364 12560
rect 27282 12502 27364 12526
rect 28300 12560 28382 12584
rect 28300 12526 28324 12560
rect 28358 12526 28382 12560
rect 28300 12502 28382 12526
rect 29318 12560 29400 12584
rect 29318 12526 29342 12560
rect 29376 12526 29400 12560
rect 29318 12502 29400 12526
rect 30336 12560 30418 12584
rect 30336 12526 30360 12560
rect 30394 12526 30418 12560
rect 30336 12502 30418 12526
rect 31354 12560 31436 12584
rect 31354 12526 31378 12560
rect 31412 12526 31436 12560
rect 31354 12502 31436 12526
rect 32372 12560 32454 12584
rect 32372 12526 32396 12560
rect 32430 12526 32454 12560
rect 32372 12502 32454 12526
rect 33390 12560 33472 12584
rect 33390 12526 33414 12560
rect 33448 12526 33472 12560
rect 33390 12502 33472 12526
rect 10928 12436 10962 12452
rect 3290 12402 3350 12404
rect 4304 12402 4364 12404
rect 8378 12402 8438 12404
rect 9394 12402 9454 12404
rect 1742 12348 1824 12372
rect 1998 12368 2014 12402
rect 2570 12368 2586 12402
rect 1742 12314 1766 12348
rect 1800 12314 1824 12348
rect 1742 12290 1824 12314
rect 2760 12348 2842 12372
rect 3016 12368 3032 12402
rect 3588 12368 3604 12402
rect 2760 12314 2784 12348
rect 2818 12314 2842 12348
rect 1998 12260 2014 12294
rect 2570 12260 2586 12294
rect 2760 12290 2842 12314
rect 3778 12348 3860 12372
rect 4034 12368 4050 12402
rect 4606 12368 4622 12402
rect 3778 12314 3802 12348
rect 3836 12314 3860 12348
rect 3016 12260 3032 12294
rect 3588 12260 3604 12294
rect 3778 12290 3860 12314
rect 4796 12348 4878 12372
rect 5052 12368 5068 12402
rect 5624 12368 5640 12402
rect 4796 12314 4820 12348
rect 4854 12314 4878 12348
rect 4034 12260 4050 12294
rect 4606 12260 4622 12294
rect 4796 12290 4878 12314
rect 5814 12348 5896 12372
rect 6070 12368 6086 12402
rect 6642 12368 6658 12402
rect 5814 12314 5838 12348
rect 5872 12314 5896 12348
rect 5052 12260 5068 12294
rect 5624 12260 5640 12294
rect 5814 12290 5896 12314
rect 6832 12348 6914 12372
rect 7088 12368 7104 12402
rect 7660 12368 7676 12402
rect 6832 12314 6856 12348
rect 6890 12314 6914 12348
rect 6070 12260 6086 12294
rect 6642 12260 6658 12294
rect 6832 12290 6914 12314
rect 7850 12348 7932 12372
rect 8106 12368 8122 12402
rect 8678 12368 8694 12402
rect 7850 12314 7874 12348
rect 7908 12314 7932 12348
rect 7088 12260 7104 12294
rect 7660 12260 7676 12294
rect 7850 12290 7932 12314
rect 8868 12348 8950 12372
rect 9124 12368 9140 12402
rect 9696 12368 9712 12402
rect 8868 12314 8892 12348
rect 8926 12314 8950 12348
rect 8106 12260 8122 12294
rect 8678 12260 8694 12294
rect 8868 12290 8950 12314
rect 9886 12348 9968 12372
rect 10142 12368 10158 12402
rect 10714 12368 10730 12402
rect 9886 12314 9910 12348
rect 9944 12314 9968 12348
rect 9124 12260 9140 12294
rect 9696 12260 9712 12294
rect 9886 12290 9968 12314
rect 10914 12348 10996 12372
rect 10914 12314 10938 12348
rect 10972 12314 10996 12348
rect 10142 12260 10158 12294
rect 10714 12260 10730 12294
rect 10914 12290 10996 12314
rect 1766 12210 1800 12226
rect 1766 11618 1800 11634
rect 2784 12210 2818 12226
rect 2784 11618 2818 11634
rect 3802 12210 3836 12226
rect 3802 11618 3836 11634
rect 4820 12210 4854 12226
rect 4820 11618 4854 11634
rect 5838 12210 5872 12226
rect 5838 11618 5872 11634
rect 6856 12210 6890 12226
rect 6856 11618 6890 11634
rect 7874 12210 7908 12226
rect 7874 11618 7908 11634
rect 8892 12210 8926 12226
rect 8892 11618 8926 11634
rect 9910 12210 9944 12226
rect 9910 11618 9944 11634
rect 10928 12210 10962 12226
rect 13764 12176 13780 12210
rect 14336 12176 14352 12210
rect 14782 12176 14798 12210
rect 15354 12176 15370 12210
rect 15800 12176 15816 12210
rect 16372 12176 16388 12210
rect 16818 12176 16834 12210
rect 17390 12176 17406 12210
rect 17836 12176 17852 12210
rect 18408 12176 18424 12210
rect 18854 12176 18870 12210
rect 19426 12176 19442 12210
rect 19872 12176 19888 12210
rect 20444 12176 20460 12210
rect 20890 12176 20906 12210
rect 21462 12176 21478 12210
rect 21908 12176 21924 12210
rect 22480 12176 22496 12210
rect 22926 12176 22942 12210
rect 23498 12176 23514 12210
rect 23944 12176 23960 12210
rect 24516 12176 24532 12210
rect 24962 12176 24978 12210
rect 25534 12176 25550 12210
rect 25980 12176 25996 12210
rect 26552 12176 26568 12210
rect 26998 12176 27014 12210
rect 27570 12176 27586 12210
rect 28016 12176 28032 12210
rect 28588 12176 28604 12210
rect 29034 12176 29050 12210
rect 29606 12176 29622 12210
rect 30052 12176 30068 12210
rect 30624 12176 30640 12210
rect 31070 12176 31086 12210
rect 31642 12176 31658 12210
rect 32088 12176 32104 12210
rect 32660 12176 32676 12210
rect 33106 12176 33122 12210
rect 33678 12176 33694 12210
rect 23188 12170 23248 12176
rect 10928 11618 10962 11634
rect 13532 12126 13566 12142
rect 3294 11584 3354 11586
rect 4308 11584 4368 11586
rect 8382 11584 8442 11586
rect 9398 11584 9458 11586
rect 1742 11530 1824 11554
rect 1998 11550 2014 11584
rect 2570 11550 2586 11584
rect 1742 11496 1766 11530
rect 1800 11496 1824 11530
rect 1742 11472 1824 11496
rect 2760 11530 2842 11554
rect 3016 11550 3032 11584
rect 3588 11550 3604 11584
rect 2760 11496 2784 11530
rect 2818 11496 2842 11530
rect 1998 11442 2014 11476
rect 2570 11442 2586 11476
rect 2760 11472 2842 11496
rect 3778 11530 3860 11554
rect 4034 11550 4050 11584
rect 4606 11550 4622 11584
rect 3778 11496 3802 11530
rect 3836 11496 3860 11530
rect 3016 11442 3032 11476
rect 3588 11442 3604 11476
rect 3778 11472 3860 11496
rect 4796 11530 4878 11554
rect 5052 11550 5068 11584
rect 5624 11550 5640 11584
rect 4796 11496 4820 11530
rect 4854 11496 4878 11530
rect 4034 11442 4050 11476
rect 4606 11442 4622 11476
rect 4796 11472 4878 11496
rect 5814 11530 5896 11554
rect 6070 11550 6086 11584
rect 6642 11550 6658 11584
rect 5814 11496 5838 11530
rect 5872 11496 5896 11530
rect 5052 11442 5068 11476
rect 5624 11442 5640 11476
rect 5814 11472 5896 11496
rect 6832 11530 6914 11554
rect 7088 11550 7104 11584
rect 7660 11550 7676 11584
rect 6832 11496 6856 11530
rect 6890 11496 6914 11530
rect 6070 11442 6086 11476
rect 6642 11442 6658 11476
rect 6832 11472 6914 11496
rect 7850 11530 7932 11554
rect 8106 11550 8122 11584
rect 8678 11550 8694 11584
rect 7850 11496 7874 11530
rect 7908 11496 7932 11530
rect 7088 11442 7104 11476
rect 7660 11442 7676 11476
rect 7850 11472 7932 11496
rect 8868 11530 8950 11554
rect 9124 11550 9140 11584
rect 9696 11550 9712 11584
rect 8868 11496 8892 11530
rect 8926 11496 8950 11530
rect 8106 11442 8122 11476
rect 8678 11442 8694 11476
rect 8868 11472 8950 11496
rect 9886 11530 9968 11554
rect 10142 11550 10158 11584
rect 10714 11550 10730 11584
rect 9886 11496 9910 11530
rect 9944 11496 9968 11530
rect 9124 11442 9140 11476
rect 9696 11442 9712 11476
rect 9886 11472 9968 11496
rect 10914 11530 10996 11554
rect 13532 11534 13566 11550
rect 14550 12126 14584 12142
rect 14550 11534 14584 11550
rect 15568 12126 15602 12142
rect 15568 11534 15602 11550
rect 16586 12126 16620 12142
rect 16586 11534 16620 11550
rect 17604 12126 17638 12142
rect 17604 11534 17638 11550
rect 18622 12126 18656 12142
rect 18622 11534 18656 11550
rect 19640 12126 19674 12142
rect 19640 11534 19674 11550
rect 20658 12126 20692 12142
rect 20658 11534 20692 11550
rect 21676 12126 21710 12142
rect 21676 11534 21710 11550
rect 22694 12126 22728 12142
rect 22694 11534 22728 11550
rect 23712 12126 23746 12142
rect 23712 11534 23746 11550
rect 24730 12126 24764 12142
rect 24730 11534 24764 11550
rect 25748 12126 25782 12142
rect 25748 11534 25782 11550
rect 26766 12126 26800 12142
rect 26766 11534 26800 11550
rect 27784 12126 27818 12142
rect 27784 11534 27818 11550
rect 28802 12126 28836 12142
rect 28802 11534 28836 11550
rect 29820 12126 29854 12142
rect 29820 11534 29854 11550
rect 30838 12126 30872 12142
rect 30838 11534 30872 11550
rect 31856 12126 31890 12142
rect 31856 11534 31890 11550
rect 32874 12126 32908 12142
rect 32874 11534 32908 11550
rect 33892 12126 33926 12142
rect 33892 11534 33926 11550
rect 10914 11496 10938 11530
rect 10972 11496 10996 11530
rect 19116 11500 19176 11506
rect 21152 11500 21212 11506
rect 22172 11500 22232 11506
rect 27244 11500 27304 11506
rect 10142 11442 10158 11476
rect 10714 11442 10730 11476
rect 10914 11472 10996 11496
rect 13764 11466 13780 11500
rect 14336 11466 14352 11500
rect 14782 11466 14798 11500
rect 15354 11466 15370 11500
rect 15800 11466 15816 11500
rect 16372 11466 16388 11500
rect 16818 11466 16834 11500
rect 17390 11466 17406 11500
rect 17836 11466 17852 11500
rect 18408 11466 18424 11500
rect 18854 11466 18870 11500
rect 19426 11466 19442 11500
rect 19872 11466 19888 11500
rect 20444 11466 20460 11500
rect 20890 11466 20906 11500
rect 21462 11466 21478 11500
rect 21908 11466 21924 11500
rect 22480 11466 22496 11500
rect 22926 11466 22942 11500
rect 23498 11466 23514 11500
rect 23944 11466 23960 11500
rect 24516 11466 24532 11500
rect 24962 11466 24978 11500
rect 25534 11466 25550 11500
rect 25980 11466 25996 11500
rect 26552 11466 26568 11500
rect 26998 11466 27014 11500
rect 27570 11466 27586 11500
rect 28016 11466 28032 11500
rect 28588 11466 28604 11500
rect 29034 11466 29050 11500
rect 29606 11466 29622 11500
rect 30052 11466 30068 11500
rect 30624 11466 30640 11500
rect 31070 11466 31086 11500
rect 31642 11466 31658 11500
rect 32088 11466 32104 11500
rect 32660 11466 32676 11500
rect 33106 11466 33122 11500
rect 33678 11466 33694 11500
rect 1766 11392 1800 11408
rect 1766 10800 1800 10816
rect 2784 11392 2818 11408
rect 2784 10800 2818 10816
rect 3802 11392 3836 11408
rect 3802 10800 3836 10816
rect 4820 11392 4854 11408
rect 4820 10800 4854 10816
rect 5838 11392 5872 11408
rect 5838 10800 5872 10816
rect 6856 11392 6890 11408
rect 6856 10800 6890 10816
rect 7874 11392 7908 11408
rect 7874 10800 7908 10816
rect 8892 11392 8926 11408
rect 8892 10800 8926 10816
rect 9910 11392 9944 11408
rect 9910 10800 9944 10816
rect 10928 11392 10962 11408
rect 14036 11254 14118 11278
rect 14036 11220 14060 11254
rect 14094 11220 14118 11254
rect 14036 11196 14118 11220
rect 15054 11254 15136 11278
rect 15054 11220 15078 11254
rect 15112 11220 15136 11254
rect 15054 11196 15136 11220
rect 16072 11254 16154 11278
rect 16072 11220 16096 11254
rect 16130 11220 16154 11254
rect 16072 11196 16154 11220
rect 17090 11254 17172 11278
rect 17090 11220 17114 11254
rect 17148 11220 17172 11254
rect 17090 11196 17172 11220
rect 18108 11254 18190 11278
rect 18108 11220 18132 11254
rect 18166 11220 18190 11254
rect 18108 11196 18190 11220
rect 19126 11254 19208 11278
rect 19126 11220 19150 11254
rect 19184 11220 19208 11254
rect 19126 11196 19208 11220
rect 20144 11254 20226 11278
rect 20144 11220 20168 11254
rect 20202 11220 20226 11254
rect 20144 11196 20226 11220
rect 21162 11254 21244 11278
rect 21162 11220 21186 11254
rect 21220 11220 21244 11254
rect 21162 11196 21244 11220
rect 22180 11254 22262 11278
rect 22180 11220 22204 11254
rect 22238 11220 22262 11254
rect 22180 11196 22262 11220
rect 23198 11254 23280 11278
rect 23198 11220 23222 11254
rect 23256 11220 23280 11254
rect 23198 11196 23280 11220
rect 24216 11254 24298 11278
rect 24216 11220 24240 11254
rect 24274 11220 24298 11254
rect 24216 11196 24298 11220
rect 25234 11254 25316 11278
rect 25234 11220 25258 11254
rect 25292 11220 25316 11254
rect 25234 11196 25316 11220
rect 26252 11254 26334 11278
rect 26252 11220 26276 11254
rect 26310 11220 26334 11254
rect 26252 11196 26334 11220
rect 27270 11254 27352 11278
rect 27270 11220 27294 11254
rect 27328 11220 27352 11254
rect 27270 11196 27352 11220
rect 28288 11254 28370 11278
rect 28288 11220 28312 11254
rect 28346 11220 28370 11254
rect 28288 11196 28370 11220
rect 29306 11254 29388 11278
rect 29306 11220 29330 11254
rect 29364 11220 29388 11254
rect 29306 11196 29388 11220
rect 30324 11254 30406 11278
rect 30324 11220 30348 11254
rect 30382 11220 30406 11254
rect 30324 11196 30406 11220
rect 31342 11254 31424 11278
rect 31342 11220 31366 11254
rect 31400 11220 31424 11254
rect 31342 11196 31424 11220
rect 32360 11254 32442 11278
rect 32360 11220 32384 11254
rect 32418 11220 32442 11254
rect 32360 11196 32442 11220
rect 33378 11254 33460 11278
rect 33378 11220 33402 11254
rect 33436 11220 33460 11254
rect 33378 11196 33460 11220
rect 13764 10944 13780 10978
rect 14336 10944 14352 10978
rect 14782 10944 14798 10978
rect 15354 10944 15370 10978
rect 15800 10944 15816 10978
rect 16372 10944 16388 10978
rect 16818 10944 16834 10978
rect 17390 10944 17406 10978
rect 17836 10944 17852 10978
rect 18408 10944 18424 10978
rect 18854 10944 18870 10978
rect 19426 10944 19442 10978
rect 19872 10944 19888 10978
rect 20444 10944 20460 10978
rect 20890 10944 20906 10978
rect 21462 10944 21478 10978
rect 21908 10944 21924 10978
rect 22480 10944 22496 10978
rect 22926 10944 22942 10978
rect 23498 10944 23514 10978
rect 23944 10944 23960 10978
rect 24516 10944 24532 10978
rect 24962 10944 24978 10978
rect 25534 10944 25550 10978
rect 25980 10944 25996 10978
rect 26552 10944 26568 10978
rect 26998 10944 27014 10978
rect 27570 10944 27586 10978
rect 28016 10944 28032 10978
rect 28588 10944 28604 10978
rect 29034 10944 29050 10978
rect 29606 10944 29622 10978
rect 30052 10944 30068 10978
rect 30624 10944 30640 10978
rect 31070 10944 31086 10978
rect 31642 10944 31658 10978
rect 32088 10944 32104 10978
rect 32660 10944 32676 10978
rect 33106 10944 33122 10978
rect 33678 10944 33694 10978
rect 15050 10940 15110 10944
rect 16066 10940 16126 10944
rect 20142 10936 20202 10944
rect 24208 10940 24268 10944
rect 26242 10940 26302 10944
rect 32354 10940 32414 10944
rect 10928 10800 10962 10816
rect 13532 10894 13566 10910
rect 1742 10712 1824 10736
rect 1998 10732 2014 10766
rect 2570 10732 2586 10766
rect 1742 10678 1766 10712
rect 1800 10678 1824 10712
rect 1742 10654 1824 10678
rect 2760 10712 2842 10736
rect 3016 10732 3032 10766
rect 3588 10732 3604 10766
rect 2760 10678 2784 10712
rect 2818 10678 2842 10712
rect 1998 10624 2014 10658
rect 2570 10624 2586 10658
rect 2760 10654 2842 10678
rect 3778 10712 3860 10736
rect 4034 10732 4050 10766
rect 4606 10732 4622 10766
rect 3778 10678 3802 10712
rect 3836 10678 3860 10712
rect 3016 10624 3032 10658
rect 3588 10624 3604 10658
rect 3778 10654 3860 10678
rect 4796 10712 4878 10736
rect 5052 10732 5068 10766
rect 5624 10732 5640 10766
rect 4796 10678 4820 10712
rect 4854 10678 4878 10712
rect 4034 10624 4050 10658
rect 4606 10624 4622 10658
rect 4796 10654 4878 10678
rect 5814 10712 5896 10736
rect 6070 10732 6086 10766
rect 6642 10732 6658 10766
rect 5814 10678 5838 10712
rect 5872 10678 5896 10712
rect 5052 10624 5068 10658
rect 5624 10624 5640 10658
rect 5814 10654 5896 10678
rect 6832 10712 6914 10736
rect 7088 10732 7104 10766
rect 7660 10732 7676 10766
rect 6832 10678 6856 10712
rect 6890 10678 6914 10712
rect 6070 10624 6086 10658
rect 6642 10624 6658 10658
rect 6832 10654 6914 10678
rect 7850 10712 7932 10736
rect 8106 10732 8122 10766
rect 8678 10732 8694 10766
rect 7850 10678 7874 10712
rect 7908 10678 7932 10712
rect 7088 10624 7104 10658
rect 7660 10624 7676 10658
rect 7850 10654 7932 10678
rect 8868 10712 8950 10736
rect 9124 10732 9140 10766
rect 9696 10732 9712 10766
rect 8868 10678 8892 10712
rect 8926 10678 8950 10712
rect 8106 10624 8122 10658
rect 8678 10624 8694 10658
rect 8868 10654 8950 10678
rect 9886 10712 9968 10736
rect 10142 10732 10158 10766
rect 10714 10732 10730 10766
rect 9886 10678 9910 10712
rect 9944 10678 9968 10712
rect 9124 10624 9140 10658
rect 9696 10624 9712 10658
rect 9886 10654 9968 10678
rect 10914 10712 10996 10736
rect 10914 10678 10938 10712
rect 10972 10678 10996 10712
rect 10142 10624 10158 10658
rect 10714 10624 10730 10658
rect 10914 10654 10996 10678
rect 7354 10622 7414 10624
rect 1766 10574 1800 10590
rect 1766 9982 1800 9998
rect 2784 10574 2818 10590
rect 2784 9982 2818 9998
rect 3802 10574 3836 10590
rect 3802 9982 3836 9998
rect 4820 10574 4854 10590
rect 4820 9982 4854 9998
rect 5838 10574 5872 10590
rect 5838 9982 5872 9998
rect 6856 10574 6890 10590
rect 6856 9982 6890 9998
rect 7874 10574 7908 10590
rect 7874 9982 7908 9998
rect 8892 10574 8926 10590
rect 8892 9982 8926 9998
rect 9910 10574 9944 10590
rect 9910 9982 9944 9998
rect 10928 10574 10962 10590
rect 13532 10302 13566 10318
rect 14550 10894 14584 10910
rect 14550 10302 14584 10318
rect 15568 10894 15602 10910
rect 15568 10302 15602 10318
rect 16586 10894 16620 10910
rect 16586 10302 16620 10318
rect 17604 10894 17638 10910
rect 17604 10302 17638 10318
rect 18622 10894 18656 10910
rect 18622 10302 18656 10318
rect 19640 10894 19674 10910
rect 19640 10302 19674 10318
rect 20658 10894 20692 10910
rect 20658 10302 20692 10318
rect 21676 10894 21710 10910
rect 21676 10302 21710 10318
rect 22694 10894 22728 10910
rect 22694 10302 22728 10318
rect 23712 10894 23746 10910
rect 23712 10302 23746 10318
rect 24730 10894 24764 10910
rect 24730 10302 24764 10318
rect 25748 10894 25782 10910
rect 25748 10302 25782 10318
rect 26766 10894 26800 10910
rect 26766 10302 26800 10318
rect 27784 10894 27818 10910
rect 27784 10302 27818 10318
rect 28802 10894 28836 10910
rect 28802 10302 28836 10318
rect 29820 10894 29854 10910
rect 29820 10302 29854 10318
rect 30838 10894 30872 10910
rect 30838 10302 30872 10318
rect 31856 10894 31890 10910
rect 31856 10302 31890 10318
rect 32874 10894 32908 10910
rect 32874 10302 32908 10318
rect 33892 10894 33926 10910
rect 33926 10318 33932 10366
rect 33892 10302 33926 10318
rect 17076 10268 17136 10270
rect 13764 10234 13780 10268
rect 14336 10234 14352 10268
rect 14782 10234 14798 10268
rect 15354 10234 15370 10268
rect 15800 10234 15816 10268
rect 16372 10234 16388 10268
rect 16818 10234 16834 10268
rect 17390 10234 17406 10268
rect 17836 10234 17852 10268
rect 18408 10234 18424 10268
rect 18854 10234 18870 10268
rect 19426 10234 19442 10268
rect 19872 10234 19888 10268
rect 20444 10234 20460 10268
rect 20890 10234 20906 10268
rect 21462 10234 21478 10268
rect 21908 10234 21924 10268
rect 22480 10234 22496 10268
rect 22926 10234 22942 10268
rect 23498 10234 23514 10268
rect 23944 10234 23960 10268
rect 24516 10234 24532 10268
rect 24962 10234 24978 10268
rect 25534 10234 25550 10268
rect 25980 10234 25996 10268
rect 26552 10234 26568 10268
rect 26998 10234 27014 10268
rect 27570 10234 27586 10268
rect 28016 10234 28032 10268
rect 28588 10234 28604 10268
rect 29034 10234 29050 10268
rect 29606 10234 29622 10268
rect 30052 10234 30068 10268
rect 30624 10234 30640 10268
rect 31070 10234 31086 10268
rect 31642 10234 31658 10268
rect 32088 10234 32104 10268
rect 32660 10234 32676 10268
rect 33106 10234 33122 10268
rect 33678 10234 33694 10268
rect 19110 10230 19170 10234
rect 28268 10220 28328 10234
rect 29302 10220 29362 10234
rect 10928 9982 10962 9998
rect 14024 10018 14106 10042
rect 14024 9984 14048 10018
rect 14082 9984 14106 10018
rect 14024 9960 14106 9984
rect 15042 10018 15124 10042
rect 15042 9984 15066 10018
rect 15100 9984 15124 10018
rect 15042 9960 15124 9984
rect 16060 10018 16142 10042
rect 16060 9984 16084 10018
rect 16118 9984 16142 10018
rect 16060 9960 16142 9984
rect 17078 10018 17160 10042
rect 17078 9984 17102 10018
rect 17136 9984 17160 10018
rect 17078 9960 17160 9984
rect 18096 10018 18178 10042
rect 18096 9984 18120 10018
rect 18154 9984 18178 10018
rect 18096 9960 18178 9984
rect 19114 10018 19196 10042
rect 19114 9984 19138 10018
rect 19172 9984 19196 10018
rect 19114 9960 19196 9984
rect 20132 10018 20214 10042
rect 20132 9984 20156 10018
rect 20190 9984 20214 10018
rect 20132 9960 20214 9984
rect 21150 10018 21232 10042
rect 21150 9984 21174 10018
rect 21208 9984 21232 10018
rect 21150 9960 21232 9984
rect 22168 10018 22250 10042
rect 22168 9984 22192 10018
rect 22226 9984 22250 10018
rect 22168 9960 22250 9984
rect 23186 10018 23268 10042
rect 23186 9984 23210 10018
rect 23244 9984 23268 10018
rect 23186 9960 23268 9984
rect 24204 10018 24286 10042
rect 24204 9984 24228 10018
rect 24262 9984 24286 10018
rect 24204 9960 24286 9984
rect 25222 10018 25304 10042
rect 25222 9984 25246 10018
rect 25280 9984 25304 10018
rect 25222 9960 25304 9984
rect 26240 10018 26322 10042
rect 26240 9984 26264 10018
rect 26298 9984 26322 10018
rect 26240 9960 26322 9984
rect 27258 10018 27340 10042
rect 27258 9984 27282 10018
rect 27316 9984 27340 10018
rect 27258 9960 27340 9984
rect 28276 10018 28358 10042
rect 28276 9984 28300 10018
rect 28334 9984 28358 10018
rect 28276 9960 28358 9984
rect 29294 10018 29376 10042
rect 29294 9984 29318 10018
rect 29352 9984 29376 10018
rect 29294 9960 29376 9984
rect 30312 10018 30394 10042
rect 30312 9984 30336 10018
rect 30370 9984 30394 10018
rect 30312 9960 30394 9984
rect 31330 10018 31412 10042
rect 31330 9984 31354 10018
rect 31388 9984 31412 10018
rect 31330 9960 31412 9984
rect 32348 10018 32430 10042
rect 32348 9984 32372 10018
rect 32406 9984 32430 10018
rect 32348 9960 32430 9984
rect 33366 10018 33448 10042
rect 33366 9984 33390 10018
rect 33424 9984 33448 10018
rect 33366 9960 33448 9984
rect 3280 9948 3340 9950
rect 4294 9948 4354 9950
rect 8368 9948 8428 9950
rect 9384 9948 9444 9950
rect 1742 9894 1824 9918
rect 1998 9914 2014 9948
rect 2570 9914 2586 9948
rect 1742 9860 1766 9894
rect 1800 9860 1824 9894
rect 1742 9836 1824 9860
rect 2760 9894 2842 9918
rect 3016 9914 3032 9948
rect 3588 9914 3604 9948
rect 2760 9860 2784 9894
rect 2818 9860 2842 9894
rect 1998 9806 2014 9840
rect 2570 9806 2586 9840
rect 2760 9836 2842 9860
rect 3778 9894 3860 9918
rect 4034 9914 4050 9948
rect 4606 9914 4622 9948
rect 3778 9860 3802 9894
rect 3836 9860 3860 9894
rect 3016 9806 3032 9840
rect 3588 9806 3604 9840
rect 3778 9836 3860 9860
rect 4796 9894 4878 9918
rect 5052 9914 5068 9948
rect 5624 9914 5640 9948
rect 4796 9860 4820 9894
rect 4854 9860 4878 9894
rect 4034 9806 4050 9840
rect 4606 9806 4622 9840
rect 4796 9836 4878 9860
rect 5814 9894 5896 9918
rect 6070 9914 6086 9948
rect 6642 9914 6658 9948
rect 5814 9860 5838 9894
rect 5872 9860 5896 9894
rect 5052 9806 5068 9840
rect 5624 9806 5640 9840
rect 5814 9836 5896 9860
rect 6832 9894 6914 9918
rect 7088 9914 7104 9948
rect 7660 9914 7676 9948
rect 6832 9860 6856 9894
rect 6890 9860 6914 9894
rect 6070 9806 6086 9840
rect 6642 9806 6658 9840
rect 6832 9836 6914 9860
rect 7850 9894 7932 9918
rect 8106 9914 8122 9948
rect 8678 9914 8694 9948
rect 7850 9860 7874 9894
rect 7908 9860 7932 9894
rect 7088 9806 7104 9840
rect 7660 9806 7676 9840
rect 7850 9836 7932 9860
rect 8868 9894 8950 9918
rect 9124 9914 9140 9948
rect 9696 9914 9712 9948
rect 8868 9860 8892 9894
rect 8926 9860 8950 9894
rect 8106 9806 8122 9840
rect 8678 9806 8694 9840
rect 8868 9836 8950 9860
rect 9886 9894 9968 9918
rect 10142 9914 10158 9948
rect 10714 9914 10730 9948
rect 9886 9860 9910 9894
rect 9944 9860 9968 9894
rect 9124 9806 9140 9840
rect 9696 9806 9712 9840
rect 9886 9836 9968 9860
rect 10914 9894 10996 9918
rect 10914 9860 10938 9894
rect 10972 9860 10996 9894
rect 10142 9806 10158 9840
rect 10714 9806 10730 9840
rect 10914 9836 10996 9860
rect 1766 9756 1800 9772
rect 1766 9164 1800 9180
rect 2784 9756 2818 9772
rect 2784 9164 2818 9180
rect 3802 9756 3836 9772
rect 3802 9164 3836 9180
rect 4820 9756 4854 9772
rect 4820 9164 4854 9180
rect 5838 9756 5872 9772
rect 5838 9164 5872 9180
rect 6856 9756 6890 9772
rect 6856 9164 6890 9180
rect 7874 9756 7908 9772
rect 7874 9164 7908 9180
rect 8892 9756 8926 9772
rect 8892 9164 8926 9180
rect 9910 9756 9944 9772
rect 9910 9164 9944 9180
rect 10928 9756 10962 9772
rect 13762 9710 13778 9744
rect 14334 9710 14350 9744
rect 14780 9710 14796 9744
rect 15352 9710 15368 9744
rect 15798 9710 15814 9744
rect 16370 9710 16386 9744
rect 16816 9710 16832 9744
rect 17388 9710 17404 9744
rect 17834 9710 17850 9744
rect 18406 9710 18422 9744
rect 18852 9710 18868 9744
rect 19424 9710 19440 9744
rect 19870 9710 19886 9744
rect 20442 9710 20458 9744
rect 20888 9710 20904 9744
rect 21460 9710 21476 9744
rect 21906 9710 21922 9744
rect 22478 9710 22494 9744
rect 22924 9710 22940 9744
rect 23496 9710 23512 9744
rect 23942 9710 23958 9744
rect 24514 9710 24530 9744
rect 24960 9710 24976 9744
rect 25532 9710 25548 9744
rect 25978 9710 25994 9744
rect 26550 9710 26566 9744
rect 26996 9710 27012 9744
rect 27568 9710 27584 9744
rect 28014 9710 28030 9744
rect 28586 9710 28602 9744
rect 29032 9710 29048 9744
rect 29604 9710 29620 9744
rect 30050 9710 30066 9744
rect 30622 9710 30638 9744
rect 31068 9710 31084 9744
rect 31640 9710 31656 9744
rect 32086 9710 32102 9744
rect 32658 9710 32674 9744
rect 33104 9710 33120 9744
rect 33676 9710 33692 9744
rect 16072 9706 16132 9710
rect 10928 9164 10962 9180
rect 13530 9660 13564 9676
rect 3284 9130 3344 9132
rect 4298 9130 4358 9132
rect 8372 9130 8432 9132
rect 9388 9130 9448 9132
rect 1742 9076 1824 9100
rect 1998 9096 2014 9130
rect 2570 9096 2586 9130
rect 1742 9042 1766 9076
rect 1800 9042 1824 9076
rect 1742 9018 1824 9042
rect 2760 9076 2842 9100
rect 3016 9096 3032 9130
rect 3588 9096 3604 9130
rect 2760 9042 2784 9076
rect 2818 9042 2842 9076
rect 1998 8988 2014 9022
rect 2570 8988 2586 9022
rect 2760 9018 2842 9042
rect 3778 9076 3860 9100
rect 4034 9096 4050 9130
rect 4606 9096 4622 9130
rect 3778 9042 3802 9076
rect 3836 9042 3860 9076
rect 3016 8988 3032 9022
rect 3588 8988 3604 9022
rect 3778 9018 3860 9042
rect 4796 9076 4878 9100
rect 5052 9096 5068 9130
rect 5624 9096 5640 9130
rect 4796 9042 4820 9076
rect 4854 9042 4878 9076
rect 4034 8988 4050 9022
rect 4606 8988 4622 9022
rect 4796 9018 4878 9042
rect 5814 9076 5896 9100
rect 6070 9096 6086 9130
rect 6642 9096 6658 9130
rect 5814 9042 5838 9076
rect 5872 9042 5896 9076
rect 5052 8988 5068 9022
rect 5624 8988 5640 9022
rect 5814 9018 5896 9042
rect 6832 9076 6914 9100
rect 7088 9096 7104 9130
rect 7660 9096 7676 9130
rect 6832 9042 6856 9076
rect 6890 9042 6914 9076
rect 6070 8988 6086 9022
rect 6642 8988 6658 9022
rect 6832 9018 6914 9042
rect 7850 9076 7932 9100
rect 8106 9096 8122 9130
rect 8678 9096 8694 9130
rect 7850 9042 7874 9076
rect 7908 9042 7932 9076
rect 7088 8988 7104 9022
rect 7660 8988 7676 9022
rect 7850 9018 7932 9042
rect 8868 9076 8950 9100
rect 9124 9096 9140 9130
rect 9696 9096 9712 9130
rect 8868 9042 8892 9076
rect 8926 9042 8950 9076
rect 8106 8988 8122 9022
rect 8678 8988 8694 9022
rect 8868 9018 8950 9042
rect 9886 9076 9968 9100
rect 10142 9096 10158 9130
rect 10714 9096 10730 9130
rect 9886 9042 9910 9076
rect 9944 9042 9968 9076
rect 9124 8988 9140 9022
rect 9696 8988 9712 9022
rect 9886 9018 9968 9042
rect 10914 9076 10996 9100
rect 10914 9042 10938 9076
rect 10972 9042 10996 9076
rect 13530 9068 13564 9084
rect 14548 9660 14582 9676
rect 14548 9068 14582 9084
rect 15566 9660 15600 9676
rect 15566 9068 15600 9084
rect 16584 9660 16618 9676
rect 16584 9068 16618 9084
rect 17602 9660 17636 9676
rect 17602 9068 17636 9084
rect 18620 9660 18654 9676
rect 18620 9068 18654 9084
rect 19638 9660 19672 9676
rect 19638 9068 19672 9084
rect 20656 9660 20690 9676
rect 20656 9068 20690 9084
rect 21674 9660 21708 9676
rect 21674 9068 21708 9084
rect 22692 9660 22726 9676
rect 22692 9068 22726 9084
rect 23710 9660 23744 9676
rect 23710 9068 23744 9084
rect 24728 9660 24762 9676
rect 24728 9068 24762 9084
rect 25746 9660 25780 9676
rect 25746 9068 25780 9084
rect 26764 9660 26798 9676
rect 26764 9068 26798 9084
rect 27782 9660 27816 9676
rect 27782 9068 27816 9084
rect 28800 9660 28834 9676
rect 28800 9068 28834 9084
rect 29818 9660 29852 9676
rect 29818 9068 29852 9084
rect 30836 9660 30870 9676
rect 30836 9068 30870 9084
rect 31854 9660 31888 9676
rect 31854 9068 31888 9084
rect 32872 9660 32906 9676
rect 32872 9068 32906 9084
rect 33890 9660 33924 9676
rect 33890 9068 33924 9084
rect 10142 8988 10158 9022
rect 10714 8988 10730 9022
rect 10914 9018 10996 9042
rect 21140 9034 21200 9038
rect 22168 9034 22228 9036
rect 24212 9034 24272 9038
rect 13762 9000 13778 9034
rect 14334 9000 14350 9034
rect 14780 9000 14796 9034
rect 15352 9000 15368 9034
rect 15798 9000 15814 9034
rect 16370 9000 16386 9034
rect 16816 9000 16832 9034
rect 17388 9000 17404 9034
rect 17834 9000 17850 9034
rect 18406 9000 18422 9034
rect 18852 9000 18868 9034
rect 19424 9000 19440 9034
rect 19870 9000 19886 9034
rect 20442 9000 20458 9034
rect 20888 9000 20904 9034
rect 21460 9000 21476 9034
rect 21906 9000 21922 9034
rect 22478 9000 22494 9034
rect 22924 9000 22940 9034
rect 23496 9000 23512 9034
rect 23942 9000 23958 9034
rect 24514 9000 24530 9034
rect 24960 9000 24976 9034
rect 25532 9000 25548 9034
rect 25978 9000 25994 9034
rect 26550 9000 26566 9034
rect 26996 9000 27012 9034
rect 27568 9000 27584 9034
rect 28014 9000 28030 9034
rect 28586 9000 28602 9034
rect 29032 9000 29048 9034
rect 29604 9000 29620 9034
rect 30050 9000 30066 9034
rect 30622 9000 30638 9034
rect 31068 9000 31084 9034
rect 31640 9000 31656 9034
rect 32086 9000 32102 9034
rect 32658 9000 32674 9034
rect 33104 9000 33120 9034
rect 33676 9000 33692 9034
rect 1766 8938 1800 8954
rect 1766 8346 1800 8362
rect 2784 8938 2818 8954
rect 2784 8346 2818 8362
rect 3802 8938 3836 8954
rect 3802 8346 3836 8362
rect 4820 8938 4854 8954
rect 4820 8346 4854 8362
rect 5838 8938 5872 8954
rect 5838 8346 5872 8362
rect 6856 8938 6890 8954
rect 6856 8346 6890 8362
rect 7874 8938 7908 8954
rect 7874 8346 7908 8362
rect 8892 8938 8926 8954
rect 8892 8346 8926 8362
rect 9910 8938 9944 8954
rect 9910 8346 9944 8362
rect 10928 8938 10962 8954
rect 14024 8794 14106 8818
rect 14024 8760 14048 8794
rect 14082 8760 14106 8794
rect 14024 8736 14106 8760
rect 15042 8794 15124 8818
rect 15042 8760 15066 8794
rect 15100 8760 15124 8794
rect 15042 8736 15124 8760
rect 16060 8794 16142 8818
rect 16060 8760 16084 8794
rect 16118 8760 16142 8794
rect 16060 8736 16142 8760
rect 17078 8794 17160 8818
rect 17078 8760 17102 8794
rect 17136 8760 17160 8794
rect 17078 8736 17160 8760
rect 18096 8794 18178 8818
rect 18096 8760 18120 8794
rect 18154 8760 18178 8794
rect 18096 8736 18178 8760
rect 19114 8794 19196 8818
rect 19114 8760 19138 8794
rect 19172 8760 19196 8794
rect 19114 8736 19196 8760
rect 20132 8794 20214 8818
rect 20132 8760 20156 8794
rect 20190 8760 20214 8794
rect 20132 8736 20214 8760
rect 21150 8794 21232 8818
rect 21150 8760 21174 8794
rect 21208 8760 21232 8794
rect 21150 8736 21232 8760
rect 22168 8794 22250 8818
rect 22168 8760 22192 8794
rect 22226 8760 22250 8794
rect 22168 8736 22250 8760
rect 23186 8794 23268 8818
rect 23186 8760 23210 8794
rect 23244 8760 23268 8794
rect 23186 8736 23268 8760
rect 24204 8794 24286 8818
rect 24204 8760 24228 8794
rect 24262 8760 24286 8794
rect 24204 8736 24286 8760
rect 25222 8794 25304 8818
rect 25222 8760 25246 8794
rect 25280 8760 25304 8794
rect 25222 8736 25304 8760
rect 26240 8794 26322 8818
rect 26240 8760 26264 8794
rect 26298 8760 26322 8794
rect 26240 8736 26322 8760
rect 27258 8794 27340 8818
rect 27258 8760 27282 8794
rect 27316 8760 27340 8794
rect 27258 8736 27340 8760
rect 28276 8794 28358 8818
rect 28276 8760 28300 8794
rect 28334 8760 28358 8794
rect 28276 8736 28358 8760
rect 29294 8794 29376 8818
rect 29294 8760 29318 8794
rect 29352 8760 29376 8794
rect 29294 8736 29376 8760
rect 30312 8794 30394 8818
rect 30312 8760 30336 8794
rect 30370 8760 30394 8794
rect 30312 8736 30394 8760
rect 31330 8794 31412 8818
rect 31330 8760 31354 8794
rect 31388 8760 31412 8794
rect 31330 8736 31412 8760
rect 32348 8794 32430 8818
rect 32348 8760 32372 8794
rect 32406 8760 32430 8794
rect 32348 8736 32430 8760
rect 33366 8794 33448 8818
rect 33366 8760 33390 8794
rect 33424 8760 33448 8794
rect 33366 8736 33448 8760
rect 13762 8476 13778 8510
rect 14334 8476 14350 8510
rect 14780 8476 14796 8510
rect 15352 8476 15368 8510
rect 15798 8476 15814 8510
rect 16370 8476 16386 8510
rect 16816 8476 16832 8510
rect 17388 8476 17404 8510
rect 17834 8476 17850 8510
rect 18406 8476 18422 8510
rect 18852 8476 18868 8510
rect 19424 8476 19440 8510
rect 19870 8476 19886 8510
rect 20442 8476 20458 8510
rect 20888 8476 20904 8510
rect 21460 8476 21476 8510
rect 21906 8476 21922 8510
rect 22478 8476 22494 8510
rect 22924 8476 22940 8510
rect 23496 8476 23512 8510
rect 23942 8476 23958 8510
rect 24514 8476 24530 8510
rect 24960 8476 24976 8510
rect 25532 8476 25548 8510
rect 25978 8476 25994 8510
rect 26550 8476 26566 8510
rect 26996 8476 27012 8510
rect 27568 8476 27584 8510
rect 28014 8476 28030 8510
rect 28586 8476 28602 8510
rect 29032 8476 29048 8510
rect 29604 8476 29620 8510
rect 30050 8476 30066 8510
rect 30622 8476 30638 8510
rect 31068 8476 31084 8510
rect 31640 8476 31656 8510
rect 32086 8476 32102 8510
rect 32658 8476 32674 8510
rect 33104 8476 33120 8510
rect 33676 8476 33692 8510
rect 10928 8346 10962 8362
rect 13530 8426 13564 8442
rect 2258 8312 2318 8314
rect 3284 8312 3344 8316
rect 4298 8312 4358 8316
rect 5318 8312 5378 8314
rect 6340 8312 6400 8314
rect 8372 8312 8432 8316
rect 9388 8312 9448 8316
rect 10408 8312 10468 8314
rect 1742 8258 1824 8282
rect 1998 8278 2014 8312
rect 2570 8278 2586 8312
rect 1742 8224 1766 8258
rect 1800 8224 1824 8258
rect 1742 8200 1824 8224
rect 2760 8258 2842 8282
rect 3016 8278 3032 8312
rect 3588 8278 3604 8312
rect 2760 8224 2784 8258
rect 2818 8224 2842 8258
rect 1998 8170 2014 8204
rect 2570 8170 2586 8204
rect 2760 8200 2842 8224
rect 3778 8258 3860 8282
rect 4034 8278 4050 8312
rect 4606 8278 4622 8312
rect 3778 8224 3802 8258
rect 3836 8224 3860 8258
rect 3016 8170 3032 8204
rect 3588 8170 3604 8204
rect 3778 8200 3860 8224
rect 4796 8258 4878 8282
rect 5052 8278 5068 8312
rect 5624 8278 5640 8312
rect 4796 8224 4820 8258
rect 4854 8224 4878 8258
rect 4034 8170 4050 8204
rect 4606 8170 4622 8204
rect 4796 8200 4878 8224
rect 5814 8258 5896 8282
rect 6070 8278 6086 8312
rect 6642 8278 6658 8312
rect 5814 8224 5838 8258
rect 5872 8224 5896 8258
rect 5052 8170 5068 8204
rect 5624 8170 5640 8204
rect 5814 8200 5896 8224
rect 6832 8258 6914 8282
rect 7088 8278 7104 8312
rect 7660 8278 7676 8312
rect 6832 8224 6856 8258
rect 6890 8224 6914 8258
rect 6070 8170 6086 8204
rect 6642 8170 6658 8204
rect 6832 8200 6914 8224
rect 7850 8258 7932 8282
rect 8106 8278 8122 8312
rect 8678 8278 8694 8312
rect 7850 8224 7874 8258
rect 7908 8224 7932 8258
rect 7088 8170 7104 8204
rect 7660 8170 7676 8204
rect 7850 8200 7932 8224
rect 8868 8258 8950 8282
rect 9124 8278 9140 8312
rect 9696 8278 9712 8312
rect 8868 8224 8892 8258
rect 8926 8224 8950 8258
rect 8106 8170 8122 8204
rect 8678 8170 8694 8204
rect 8868 8200 8950 8224
rect 9886 8258 9968 8282
rect 10142 8278 10158 8312
rect 10714 8278 10730 8312
rect 9886 8224 9910 8258
rect 9944 8224 9968 8258
rect 9124 8170 9140 8204
rect 9696 8170 9712 8204
rect 9886 8200 9968 8224
rect 10914 8258 10996 8282
rect 10914 8224 10938 8258
rect 10972 8224 10996 8258
rect 10142 8170 10158 8204
rect 10714 8170 10730 8204
rect 10914 8200 10996 8224
rect 1766 8120 1800 8136
rect 1766 7528 1800 7544
rect 2784 8120 2818 8136
rect 2784 7528 2818 7544
rect 3802 8120 3836 8136
rect 3802 7528 3836 7544
rect 4820 8120 4854 8136
rect 4820 7528 4854 7544
rect 5838 8120 5872 8136
rect 5838 7528 5872 7544
rect 6856 8120 6890 8136
rect 6856 7528 6890 7544
rect 7874 8120 7908 8136
rect 7874 7528 7908 7544
rect 8892 8120 8926 8136
rect 8892 7528 8926 7544
rect 9910 8120 9944 8136
rect 9910 7528 9944 7544
rect 10928 8120 10962 8136
rect 13530 7834 13564 7850
rect 14548 8426 14582 8442
rect 14548 7834 14582 7850
rect 15566 8426 15600 8442
rect 15566 7834 15600 7850
rect 16584 8426 16618 8442
rect 16584 7834 16618 7850
rect 17602 8426 17636 8442
rect 17602 7834 17636 7850
rect 18620 8426 18654 8442
rect 18620 7834 18654 7850
rect 19638 8426 19672 8442
rect 19638 7834 19672 7850
rect 20656 8426 20690 8442
rect 20656 7834 20690 7850
rect 21674 8426 21708 8442
rect 21674 7834 21708 7850
rect 22692 8426 22726 8442
rect 22692 7834 22726 7850
rect 23710 8426 23744 8442
rect 23710 7834 23744 7850
rect 24728 8426 24762 8442
rect 24728 7834 24762 7850
rect 25746 8426 25780 8442
rect 25746 7834 25780 7850
rect 26764 8426 26798 8442
rect 26764 7834 26798 7850
rect 27782 8426 27816 8442
rect 27782 7834 27816 7850
rect 28800 8426 28834 8442
rect 28800 7834 28834 7850
rect 29818 8426 29852 8442
rect 29818 7834 29852 7850
rect 30836 8426 30870 8442
rect 30836 7834 30870 7850
rect 31854 8426 31888 8442
rect 31854 7834 31888 7850
rect 32872 8426 32906 8442
rect 32872 7834 32906 7850
rect 33890 8426 33924 8442
rect 33890 7834 33924 7850
rect 13762 7766 13778 7800
rect 14334 7766 14350 7800
rect 14780 7766 14796 7800
rect 15352 7766 15368 7800
rect 15798 7766 15814 7800
rect 16370 7766 16386 7800
rect 16816 7766 16832 7800
rect 17388 7766 17404 7800
rect 17834 7766 17850 7800
rect 18406 7766 18422 7800
rect 18852 7766 18868 7800
rect 19424 7766 19440 7800
rect 19870 7766 19886 7800
rect 20442 7766 20458 7800
rect 20888 7766 20904 7800
rect 21460 7766 21476 7800
rect 21906 7766 21922 7800
rect 22478 7766 22494 7800
rect 22924 7766 22940 7800
rect 23496 7766 23512 7800
rect 23942 7766 23958 7800
rect 24514 7766 24530 7800
rect 24960 7766 24976 7800
rect 25532 7766 25548 7800
rect 25978 7766 25994 7800
rect 26550 7766 26566 7800
rect 26996 7766 27012 7800
rect 27568 7766 27584 7800
rect 28014 7766 28030 7800
rect 28586 7766 28602 7800
rect 29032 7766 29048 7800
rect 29604 7766 29620 7800
rect 30050 7766 30066 7800
rect 30622 7766 30638 7800
rect 31068 7766 31084 7800
rect 31640 7766 31656 7800
rect 32086 7766 32102 7800
rect 32658 7766 32674 7800
rect 33104 7766 33120 7800
rect 33676 7766 33692 7800
rect 10928 7528 10962 7544
rect 14036 7558 14118 7582
rect 14036 7524 14060 7558
rect 14094 7524 14118 7558
rect 14036 7500 14118 7524
rect 15054 7558 15136 7582
rect 15054 7524 15078 7558
rect 15112 7524 15136 7558
rect 15054 7500 15136 7524
rect 16072 7558 16154 7582
rect 16072 7524 16096 7558
rect 16130 7524 16154 7558
rect 16072 7500 16154 7524
rect 17090 7558 17172 7582
rect 17090 7524 17114 7558
rect 17148 7524 17172 7558
rect 17090 7500 17172 7524
rect 18108 7558 18190 7582
rect 18108 7524 18132 7558
rect 18166 7524 18190 7558
rect 18108 7500 18190 7524
rect 19126 7558 19208 7582
rect 19126 7524 19150 7558
rect 19184 7524 19208 7558
rect 19126 7500 19208 7524
rect 20144 7558 20226 7582
rect 20144 7524 20168 7558
rect 20202 7524 20226 7558
rect 20144 7500 20226 7524
rect 21162 7558 21244 7582
rect 21162 7524 21186 7558
rect 21220 7524 21244 7558
rect 21162 7500 21244 7524
rect 22180 7558 22262 7582
rect 22180 7524 22204 7558
rect 22238 7524 22262 7558
rect 22180 7500 22262 7524
rect 23198 7558 23280 7582
rect 23198 7524 23222 7558
rect 23256 7524 23280 7558
rect 23198 7500 23280 7524
rect 24216 7558 24298 7582
rect 24216 7524 24240 7558
rect 24274 7524 24298 7558
rect 24216 7500 24298 7524
rect 25234 7558 25316 7582
rect 25234 7524 25258 7558
rect 25292 7524 25316 7558
rect 25234 7500 25316 7524
rect 26252 7558 26334 7582
rect 26252 7524 26276 7558
rect 26310 7524 26334 7558
rect 26252 7500 26334 7524
rect 27270 7558 27352 7582
rect 27270 7524 27294 7558
rect 27328 7524 27352 7558
rect 27270 7500 27352 7524
rect 28288 7558 28370 7582
rect 28288 7524 28312 7558
rect 28346 7524 28370 7558
rect 28288 7500 28370 7524
rect 29306 7558 29388 7582
rect 29306 7524 29330 7558
rect 29364 7524 29388 7558
rect 29306 7500 29388 7524
rect 30324 7558 30406 7582
rect 30324 7524 30348 7558
rect 30382 7524 30406 7558
rect 30324 7500 30406 7524
rect 31342 7558 31424 7582
rect 31342 7524 31366 7558
rect 31400 7524 31424 7558
rect 31342 7500 31424 7524
rect 32360 7558 32442 7582
rect 32360 7524 32384 7558
rect 32418 7524 32442 7558
rect 32360 7500 32442 7524
rect 33378 7558 33460 7582
rect 33378 7524 33402 7558
rect 33436 7524 33460 7558
rect 33378 7500 33460 7524
rect 1998 7460 2014 7494
rect 2570 7460 2586 7494
rect 3016 7460 3032 7494
rect 3588 7460 3604 7494
rect 4034 7460 4050 7494
rect 4606 7460 4622 7494
rect 5052 7460 5068 7494
rect 5624 7460 5640 7494
rect 6070 7460 6086 7494
rect 6642 7460 6658 7494
rect 7088 7460 7104 7494
rect 7660 7460 7676 7494
rect 8106 7460 8122 7494
rect 8678 7460 8694 7494
rect 9124 7460 9140 7494
rect 9696 7460 9712 7494
rect 10142 7460 10158 7494
rect 10714 7460 10730 7494
rect 1730 7364 1812 7388
rect 1730 7330 1754 7364
rect 1788 7330 1812 7364
rect 1730 7306 1812 7330
rect 2748 7364 2830 7388
rect 2748 7330 2772 7364
rect 2806 7330 2830 7364
rect 2748 7306 2830 7330
rect 3766 7364 3848 7388
rect 3766 7330 3790 7364
rect 3824 7330 3848 7364
rect 3766 7306 3848 7330
rect 4784 7364 4866 7388
rect 4784 7330 4808 7364
rect 4842 7330 4866 7364
rect 4784 7306 4866 7330
rect 5802 7364 5884 7388
rect 5802 7330 5826 7364
rect 5860 7330 5884 7364
rect 5802 7306 5884 7330
rect 6820 7364 6902 7388
rect 6820 7330 6844 7364
rect 6878 7330 6902 7364
rect 6820 7306 6902 7330
rect 7838 7364 7920 7388
rect 7838 7330 7862 7364
rect 7896 7330 7920 7364
rect 7838 7306 7920 7330
rect 8856 7364 8938 7388
rect 8856 7330 8880 7364
rect 8914 7330 8938 7364
rect 8856 7306 8938 7330
rect 9874 7364 9956 7388
rect 9874 7330 9898 7364
rect 9932 7330 9956 7364
rect 9874 7306 9956 7330
rect 10902 7364 10984 7388
rect 10902 7330 10926 7364
rect 10960 7330 10984 7364
rect 10902 7306 10984 7330
rect 13762 7244 13778 7278
rect 14334 7244 14350 7278
rect 14780 7244 14796 7278
rect 15352 7244 15368 7278
rect 15798 7244 15814 7278
rect 16370 7244 16386 7278
rect 16816 7244 16832 7278
rect 17388 7244 17404 7278
rect 17834 7244 17850 7278
rect 18406 7244 18422 7278
rect 18852 7244 18868 7278
rect 19424 7244 19440 7278
rect 19870 7244 19886 7278
rect 20442 7244 20458 7278
rect 20888 7244 20904 7278
rect 21460 7244 21476 7278
rect 21906 7244 21922 7278
rect 22478 7244 22494 7278
rect 22924 7244 22940 7278
rect 23496 7244 23512 7278
rect 23942 7244 23958 7278
rect 24514 7244 24530 7278
rect 24960 7244 24976 7278
rect 25532 7244 25548 7278
rect 25978 7244 25994 7278
rect 26550 7244 26566 7278
rect 26996 7244 27012 7278
rect 27568 7244 27584 7278
rect 28014 7244 28030 7278
rect 28586 7244 28602 7278
rect 29032 7244 29048 7278
rect 29604 7244 29620 7278
rect 30050 7244 30066 7278
rect 30622 7244 30638 7278
rect 31068 7244 31084 7278
rect 31640 7244 31656 7278
rect 32086 7244 32102 7278
rect 32658 7244 32674 7278
rect 33104 7244 33120 7278
rect 33676 7244 33692 7278
rect 13530 7194 13564 7210
rect 13530 6602 13564 6618
rect 14548 7194 14582 7210
rect 14548 6602 14582 6618
rect 15566 7194 15600 7210
rect 15566 6602 15600 6618
rect 16584 7194 16618 7210
rect 16584 6602 16618 6618
rect 17602 7194 17636 7210
rect 17602 6602 17636 6618
rect 18620 7194 18654 7210
rect 18620 6602 18654 6618
rect 19638 7194 19672 7210
rect 19638 6602 19672 6618
rect 20656 7194 20690 7210
rect 20656 6602 20690 6618
rect 21674 7194 21708 7210
rect 21674 6602 21708 6618
rect 22692 7194 22726 7210
rect 22692 6602 22726 6618
rect 23710 7194 23744 7210
rect 23710 6602 23744 6618
rect 24728 7194 24762 7210
rect 24728 6602 24762 6618
rect 25746 7194 25780 7210
rect 25746 6602 25780 6618
rect 26764 7194 26798 7210
rect 26764 6602 26798 6618
rect 27782 7194 27816 7210
rect 27782 6602 27816 6618
rect 28800 7194 28834 7210
rect 28800 6602 28834 6618
rect 29818 7194 29852 7210
rect 29818 6602 29852 6618
rect 30836 7194 30870 7210
rect 30836 6602 30870 6618
rect 31854 7194 31888 7210
rect 31854 6602 31888 6618
rect 32872 7194 32906 7210
rect 32872 6602 32906 6618
rect 33890 7194 33924 7210
rect 33890 6602 33924 6618
rect 22180 6568 22240 6570
rect 24224 6568 24284 6572
rect 32358 6568 32418 6570
rect 13762 6534 13778 6568
rect 14334 6534 14350 6568
rect 14780 6534 14796 6568
rect 15352 6534 15368 6568
rect 15798 6534 15814 6568
rect 16370 6534 16386 6568
rect 16816 6534 16832 6568
rect 17388 6534 17404 6568
rect 17834 6534 17850 6568
rect 18406 6534 18422 6568
rect 18852 6534 18868 6568
rect 19424 6534 19440 6568
rect 19870 6534 19886 6568
rect 20442 6534 20458 6568
rect 20888 6534 20904 6568
rect 21460 6534 21476 6568
rect 21906 6534 21922 6568
rect 22478 6534 22494 6568
rect 22924 6534 22940 6568
rect 23496 6534 23512 6568
rect 23942 6534 23958 6568
rect 24514 6534 24530 6568
rect 24960 6534 24976 6568
rect 25532 6534 25548 6568
rect 25978 6534 25994 6568
rect 26550 6534 26566 6568
rect 26996 6534 27012 6568
rect 27568 6534 27584 6568
rect 28014 6534 28030 6568
rect 28586 6534 28602 6568
rect 29032 6534 29048 6568
rect 29604 6534 29620 6568
rect 30050 6534 30066 6568
rect 30622 6534 30638 6568
rect 31068 6534 31084 6568
rect 31640 6534 31656 6568
rect 32086 6534 32102 6568
rect 32658 6534 32674 6568
rect 33104 6534 33120 6568
rect 33676 6534 33692 6568
rect 934 6416 1016 6440
rect 934 6382 958 6416
rect 992 6382 1016 6416
rect 934 6358 1016 6382
rect 1952 6416 2034 6440
rect 1952 6382 1976 6416
rect 2010 6382 2034 6416
rect 1952 6358 2034 6382
rect 2970 6416 3052 6440
rect 2970 6382 2994 6416
rect 3028 6382 3052 6416
rect 2970 6358 3052 6382
rect 3988 6416 4070 6440
rect 3988 6382 4012 6416
rect 4046 6382 4070 6416
rect 3988 6358 4070 6382
rect 5006 6416 5088 6440
rect 5006 6382 5030 6416
rect 5064 6382 5088 6416
rect 5006 6358 5088 6382
rect 6024 6416 6106 6440
rect 6024 6382 6048 6416
rect 6082 6382 6106 6416
rect 6024 6358 6106 6382
rect 7042 6416 7124 6440
rect 7042 6382 7066 6416
rect 7100 6382 7124 6416
rect 7042 6358 7124 6382
rect 8060 6416 8142 6440
rect 8060 6382 8084 6416
rect 8118 6382 8142 6416
rect 8060 6358 8142 6382
rect 9078 6416 9160 6440
rect 9078 6382 9102 6416
rect 9136 6382 9160 6416
rect 9078 6358 9160 6382
rect 10096 6416 10178 6440
rect 10096 6382 10120 6416
rect 10154 6382 10178 6416
rect 10096 6358 10178 6382
rect 11114 6416 11196 6440
rect 11114 6382 11138 6416
rect 11172 6382 11196 6416
rect 11114 6358 11196 6382
rect 14036 6310 14118 6334
rect 14036 6276 14060 6310
rect 14094 6276 14118 6310
rect 14036 6252 14118 6276
rect 15054 6310 15136 6334
rect 15054 6276 15078 6310
rect 15112 6276 15136 6310
rect 15054 6252 15136 6276
rect 16072 6310 16154 6334
rect 16072 6276 16096 6310
rect 16130 6276 16154 6310
rect 16072 6252 16154 6276
rect 17090 6310 17172 6334
rect 17090 6276 17114 6310
rect 17148 6276 17172 6310
rect 17090 6252 17172 6276
rect 18108 6310 18190 6334
rect 18108 6276 18132 6310
rect 18166 6276 18190 6310
rect 18108 6252 18190 6276
rect 19126 6310 19208 6334
rect 19126 6276 19150 6310
rect 19184 6276 19208 6310
rect 19126 6252 19208 6276
rect 20144 6310 20226 6334
rect 20144 6276 20168 6310
rect 20202 6276 20226 6310
rect 20144 6252 20226 6276
rect 21162 6310 21244 6334
rect 21162 6276 21186 6310
rect 21220 6276 21244 6310
rect 21162 6252 21244 6276
rect 22180 6310 22262 6334
rect 22180 6276 22204 6310
rect 22238 6276 22262 6310
rect 22180 6252 22262 6276
rect 23198 6310 23280 6334
rect 23198 6276 23222 6310
rect 23256 6276 23280 6310
rect 23198 6252 23280 6276
rect 24216 6310 24298 6334
rect 24216 6276 24240 6310
rect 24274 6276 24298 6310
rect 24216 6252 24298 6276
rect 25234 6310 25316 6334
rect 25234 6276 25258 6310
rect 25292 6276 25316 6310
rect 25234 6252 25316 6276
rect 26252 6310 26334 6334
rect 26252 6276 26276 6310
rect 26310 6276 26334 6310
rect 26252 6252 26334 6276
rect 27270 6310 27352 6334
rect 27270 6276 27294 6310
rect 27328 6276 27352 6310
rect 27270 6252 27352 6276
rect 28288 6310 28370 6334
rect 28288 6276 28312 6310
rect 28346 6276 28370 6310
rect 28288 6252 28370 6276
rect 29306 6310 29388 6334
rect 29306 6276 29330 6310
rect 29364 6276 29388 6310
rect 29306 6252 29388 6276
rect 30324 6310 30406 6334
rect 30324 6276 30348 6310
rect 30382 6276 30406 6310
rect 30324 6252 30406 6276
rect 31342 6310 31424 6334
rect 31342 6276 31366 6310
rect 31400 6276 31424 6310
rect 31342 6252 31424 6276
rect 32360 6310 32442 6334
rect 32360 6276 32384 6310
rect 32418 6276 32442 6310
rect 32360 6252 32442 6276
rect 33378 6310 33460 6334
rect 33378 6276 33402 6310
rect 33436 6276 33460 6310
rect 33378 6252 33460 6276
rect 674 6146 690 6180
rect 1246 6146 1262 6180
rect 1692 6146 1708 6180
rect 2264 6146 2280 6180
rect 2710 6146 2726 6180
rect 3282 6146 3298 6180
rect 3728 6146 3744 6180
rect 4300 6146 4316 6180
rect 4746 6146 4762 6180
rect 5318 6146 5334 6180
rect 5764 6146 5780 6180
rect 6336 6146 6352 6180
rect 6782 6146 6798 6180
rect 7354 6146 7370 6180
rect 7800 6146 7816 6180
rect 8372 6146 8388 6180
rect 8818 6146 8834 6180
rect 9390 6146 9406 6180
rect 9836 6146 9852 6180
rect 10408 6146 10424 6180
rect 10854 6146 10870 6180
rect 11426 6146 11442 6180
rect 442 6096 476 6112
rect 442 5504 476 5520
rect 1460 6096 1494 6112
rect 1460 5504 1494 5520
rect 2478 6096 2512 6112
rect 2478 5504 2512 5520
rect 3496 6096 3530 6112
rect 3496 5504 3530 5520
rect 4514 6096 4548 6112
rect 4514 5504 4548 5520
rect 5532 6096 5566 6112
rect 5532 5504 5566 5520
rect 6550 6096 6584 6112
rect 6550 5504 6584 5520
rect 7568 6096 7602 6112
rect 7568 5504 7602 5520
rect 8586 6096 8620 6112
rect 8586 5504 8620 5520
rect 9604 6096 9638 6112
rect 9604 5504 9638 5520
rect 10622 6096 10656 6112
rect 10622 5504 10656 5520
rect 11640 6096 11674 6112
rect 13762 6010 13778 6044
rect 14334 6010 14350 6044
rect 14780 6010 14796 6044
rect 15352 6010 15368 6044
rect 15798 6010 15814 6044
rect 16370 6010 16386 6044
rect 16816 6010 16832 6044
rect 17388 6010 17404 6044
rect 17834 6010 17850 6044
rect 18406 6010 18422 6044
rect 18852 6010 18868 6044
rect 19424 6010 19440 6044
rect 19870 6010 19886 6044
rect 20442 6010 20458 6044
rect 20888 6010 20904 6044
rect 21460 6010 21476 6044
rect 21906 6010 21922 6044
rect 22478 6010 22494 6044
rect 22924 6010 22940 6044
rect 23496 6010 23512 6044
rect 23942 6010 23958 6044
rect 24514 6010 24530 6044
rect 24960 6010 24976 6044
rect 25532 6010 25548 6044
rect 25978 6010 25994 6044
rect 26550 6010 26566 6044
rect 26996 6010 27012 6044
rect 27568 6010 27584 6044
rect 28014 6010 28030 6044
rect 28586 6010 28602 6044
rect 29032 6010 29048 6044
rect 29604 6010 29620 6044
rect 30050 6010 30066 6044
rect 30622 6010 30638 6044
rect 31068 6010 31084 6044
rect 31640 6010 31656 6044
rect 32086 6010 32102 6044
rect 32658 6010 32674 6044
rect 33104 6010 33120 6044
rect 33676 6010 33692 6044
rect 11640 5504 11674 5520
rect 13530 5960 13564 5976
rect 674 5436 690 5470
rect 1246 5436 1262 5470
rect 1692 5436 1708 5470
rect 2264 5436 2280 5470
rect 2710 5436 2726 5470
rect 3282 5436 3298 5470
rect 3728 5436 3744 5470
rect 4300 5436 4316 5470
rect 4746 5436 4762 5470
rect 5318 5436 5334 5470
rect 5764 5436 5780 5470
rect 6336 5436 6352 5470
rect 6782 5436 6798 5470
rect 7354 5436 7370 5470
rect 7800 5436 7816 5470
rect 8372 5436 8388 5470
rect 8818 5436 8834 5470
rect 9390 5436 9406 5470
rect 9836 5436 9852 5470
rect 10408 5436 10424 5470
rect 10854 5436 10870 5470
rect 11426 5436 11442 5470
rect 13530 5368 13564 5384
rect 14548 5960 14582 5976
rect 14548 5368 14582 5384
rect 15566 5960 15600 5976
rect 15566 5368 15600 5384
rect 16584 5960 16618 5976
rect 16584 5368 16618 5384
rect 17602 5960 17636 5976
rect 17602 5368 17636 5384
rect 18620 5960 18654 5976
rect 18620 5368 18654 5384
rect 19638 5960 19672 5976
rect 19638 5368 19672 5384
rect 20656 5960 20690 5976
rect 20656 5368 20690 5384
rect 21674 5960 21708 5976
rect 21674 5368 21708 5384
rect 22692 5960 22726 5976
rect 22692 5368 22726 5384
rect 23710 5960 23744 5976
rect 23710 5368 23744 5384
rect 24728 5960 24762 5976
rect 24728 5368 24762 5384
rect 25746 5960 25780 5976
rect 25746 5368 25780 5384
rect 26764 5960 26798 5976
rect 26764 5368 26798 5384
rect 27782 5960 27816 5976
rect 27782 5368 27816 5384
rect 28800 5960 28834 5976
rect 28800 5368 28834 5384
rect 29818 5960 29852 5976
rect 29818 5368 29852 5384
rect 30836 5960 30870 5976
rect 30836 5368 30870 5384
rect 31854 5960 31888 5976
rect 31854 5368 31888 5384
rect 32872 5960 32906 5976
rect 32872 5368 32906 5384
rect 33890 5960 33924 5976
rect 33890 5368 33924 5384
rect 16056 5334 16116 5338
rect 13762 5300 13778 5334
rect 14334 5300 14350 5334
rect 14780 5300 14796 5334
rect 15352 5300 15368 5334
rect 15798 5300 15814 5334
rect 16370 5300 16386 5334
rect 16816 5300 16832 5334
rect 17388 5300 17404 5334
rect 17834 5300 17850 5334
rect 18406 5300 18422 5334
rect 18852 5300 18868 5334
rect 19424 5300 19440 5334
rect 19870 5300 19886 5334
rect 20442 5300 20458 5334
rect 20888 5300 20904 5334
rect 21460 5300 21476 5334
rect 21906 5300 21922 5334
rect 22478 5300 22494 5334
rect 22924 5300 22940 5334
rect 23496 5300 23512 5334
rect 23942 5300 23958 5334
rect 24514 5300 24530 5334
rect 24960 5300 24976 5334
rect 25532 5300 25548 5334
rect 25978 5300 25994 5334
rect 26550 5300 26566 5334
rect 26996 5300 27012 5334
rect 27568 5300 27584 5334
rect 28014 5300 28030 5334
rect 28586 5300 28602 5334
rect 29032 5300 29048 5334
rect 29604 5300 29620 5334
rect 30050 5300 30066 5334
rect 30622 5300 30638 5334
rect 31068 5300 31084 5334
rect 31640 5300 31656 5334
rect 32086 5300 32102 5334
rect 32658 5300 32674 5334
rect 33104 5300 33120 5334
rect 33676 5300 33692 5334
rect 946 5274 1028 5298
rect 946 5240 970 5274
rect 1004 5240 1028 5274
rect 946 5216 1028 5240
rect 1964 5274 2046 5298
rect 1964 5240 1988 5274
rect 2022 5240 2046 5274
rect 1964 5216 2046 5240
rect 2982 5274 3064 5298
rect 2982 5240 3006 5274
rect 3040 5240 3064 5274
rect 2982 5216 3064 5240
rect 4000 5274 4082 5298
rect 4000 5240 4024 5274
rect 4058 5240 4082 5274
rect 4000 5216 4082 5240
rect 5018 5274 5100 5298
rect 5018 5240 5042 5274
rect 5076 5240 5100 5274
rect 5018 5216 5100 5240
rect 6036 5274 6118 5298
rect 6036 5240 6060 5274
rect 6094 5240 6118 5274
rect 6036 5216 6118 5240
rect 7054 5274 7136 5298
rect 7054 5240 7078 5274
rect 7112 5240 7136 5274
rect 7054 5216 7136 5240
rect 8072 5274 8154 5298
rect 8072 5240 8096 5274
rect 8130 5240 8154 5274
rect 8072 5216 8154 5240
rect 9090 5274 9172 5298
rect 9090 5240 9114 5274
rect 9148 5240 9172 5274
rect 9090 5216 9172 5240
rect 10108 5274 10190 5298
rect 10108 5240 10132 5274
rect 10166 5240 10190 5274
rect 10108 5216 10190 5240
rect 11126 5274 11208 5298
rect 11126 5240 11150 5274
rect 11184 5240 11208 5274
rect 11126 5216 11208 5240
rect 14012 5074 14094 5098
rect 674 5034 690 5068
rect 1246 5034 1262 5068
rect 1692 5034 1708 5068
rect 2264 5034 2280 5068
rect 2710 5034 2726 5068
rect 3282 5034 3298 5068
rect 3728 5034 3744 5068
rect 4300 5034 4316 5068
rect 4746 5034 4762 5068
rect 5318 5034 5334 5068
rect 5764 5034 5780 5068
rect 6336 5034 6352 5068
rect 6782 5034 6798 5068
rect 7354 5034 7370 5068
rect 7800 5034 7816 5068
rect 8372 5034 8388 5068
rect 8818 5034 8834 5068
rect 9390 5034 9406 5068
rect 9836 5034 9852 5068
rect 10408 5034 10424 5068
rect 10854 5034 10870 5068
rect 11426 5034 11442 5068
rect 14012 5040 14036 5074
rect 14070 5040 14094 5074
rect 14012 5016 14094 5040
rect 15030 5074 15112 5098
rect 15030 5040 15054 5074
rect 15088 5040 15112 5074
rect 15030 5016 15112 5040
rect 16048 5074 16130 5098
rect 16048 5040 16072 5074
rect 16106 5040 16130 5074
rect 16048 5016 16130 5040
rect 17066 5074 17148 5098
rect 17066 5040 17090 5074
rect 17124 5040 17148 5074
rect 17066 5016 17148 5040
rect 18084 5074 18166 5098
rect 18084 5040 18108 5074
rect 18142 5040 18166 5074
rect 18084 5016 18166 5040
rect 19102 5074 19184 5098
rect 19102 5040 19126 5074
rect 19160 5040 19184 5074
rect 19102 5016 19184 5040
rect 20120 5074 20202 5098
rect 20120 5040 20144 5074
rect 20178 5040 20202 5074
rect 20120 5016 20202 5040
rect 21138 5074 21220 5098
rect 21138 5040 21162 5074
rect 21196 5040 21220 5074
rect 21138 5016 21220 5040
rect 22156 5074 22238 5098
rect 22156 5040 22180 5074
rect 22214 5040 22238 5074
rect 22156 5016 22238 5040
rect 23174 5074 23256 5098
rect 23174 5040 23198 5074
rect 23232 5040 23256 5074
rect 23174 5016 23256 5040
rect 24192 5074 24274 5098
rect 24192 5040 24216 5074
rect 24250 5040 24274 5074
rect 24192 5016 24274 5040
rect 25210 5074 25292 5098
rect 25210 5040 25234 5074
rect 25268 5040 25292 5074
rect 25210 5016 25292 5040
rect 26228 5074 26310 5098
rect 26228 5040 26252 5074
rect 26286 5040 26310 5074
rect 26228 5016 26310 5040
rect 27246 5074 27328 5098
rect 27246 5040 27270 5074
rect 27304 5040 27328 5074
rect 27246 5016 27328 5040
rect 28264 5074 28346 5098
rect 28264 5040 28288 5074
rect 28322 5040 28346 5074
rect 28264 5016 28346 5040
rect 29282 5074 29364 5098
rect 29282 5040 29306 5074
rect 29340 5040 29364 5074
rect 29282 5016 29364 5040
rect 30300 5074 30382 5098
rect 30300 5040 30324 5074
rect 30358 5040 30382 5074
rect 30300 5016 30382 5040
rect 31318 5074 31400 5098
rect 31318 5040 31342 5074
rect 31376 5040 31400 5074
rect 31318 5016 31400 5040
rect 32336 5074 32418 5098
rect 32336 5040 32360 5074
rect 32394 5040 32418 5074
rect 32336 5016 32418 5040
rect 33354 5074 33436 5098
rect 33354 5040 33378 5074
rect 33412 5040 33436 5074
rect 33354 5016 33436 5040
rect 442 4984 476 5000
rect 442 4392 476 4408
rect 1460 4984 1494 5000
rect 1460 4392 1494 4408
rect 2478 4984 2512 5000
rect 2478 4392 2512 4408
rect 3496 4984 3530 5000
rect 3496 4392 3530 4408
rect 4514 4984 4548 5000
rect 4514 4392 4548 4408
rect 5532 4984 5566 5000
rect 5532 4392 5566 4408
rect 6550 4984 6584 5000
rect 6550 4392 6584 4408
rect 7568 4984 7602 5000
rect 7568 4392 7602 4408
rect 8586 4984 8620 5000
rect 8586 4392 8620 4408
rect 9604 4984 9638 5000
rect 9604 4392 9638 4408
rect 10622 4984 10656 5000
rect 10622 4392 10656 4408
rect 11640 4984 11674 5000
rect 13762 4776 13778 4810
rect 14334 4776 14350 4810
rect 14780 4776 14796 4810
rect 15352 4776 15368 4810
rect 15798 4776 15814 4810
rect 16370 4776 16386 4810
rect 16816 4776 16832 4810
rect 17388 4776 17404 4810
rect 17834 4776 17850 4810
rect 18406 4776 18422 4810
rect 18852 4776 18868 4810
rect 19424 4776 19440 4810
rect 19870 4776 19886 4810
rect 20442 4776 20458 4810
rect 20888 4776 20904 4810
rect 21460 4776 21476 4810
rect 21906 4776 21922 4810
rect 22478 4776 22494 4810
rect 22924 4776 22940 4810
rect 23496 4776 23512 4810
rect 23942 4776 23958 4810
rect 24514 4776 24530 4810
rect 24960 4776 24976 4810
rect 25532 4776 25548 4810
rect 25978 4776 25994 4810
rect 26550 4776 26566 4810
rect 26996 4776 27012 4810
rect 27568 4776 27584 4810
rect 28014 4776 28030 4810
rect 28586 4776 28602 4810
rect 29032 4776 29048 4810
rect 29604 4776 29620 4810
rect 30050 4776 30066 4810
rect 30622 4776 30638 4810
rect 31068 4776 31084 4810
rect 31640 4776 31656 4810
rect 32086 4776 32102 4810
rect 32658 4776 32674 4810
rect 33104 4776 33120 4810
rect 33676 4776 33692 4810
rect 11640 4392 11674 4408
rect 13530 4726 13564 4742
rect 674 4324 690 4358
rect 1246 4324 1262 4358
rect 1692 4324 1708 4358
rect 2264 4324 2280 4358
rect 2710 4324 2726 4358
rect 3282 4324 3298 4358
rect 3728 4324 3744 4358
rect 4300 4324 4316 4358
rect 4746 4324 4762 4358
rect 5318 4324 5334 4358
rect 5764 4324 5780 4358
rect 6336 4324 6352 4358
rect 6782 4324 6798 4358
rect 7354 4324 7370 4358
rect 7800 4324 7816 4358
rect 8372 4324 8388 4358
rect 8818 4324 8834 4358
rect 9390 4324 9406 4358
rect 9836 4324 9852 4358
rect 10408 4324 10424 4358
rect 10854 4324 10870 4358
rect 11426 4324 11442 4358
rect 924 4166 1006 4190
rect 924 4132 948 4166
rect 982 4132 1006 4166
rect 924 4108 1006 4132
rect 1942 4166 2024 4190
rect 1942 4132 1966 4166
rect 2000 4132 2024 4166
rect 1942 4108 2024 4132
rect 2960 4166 3042 4190
rect 2960 4132 2984 4166
rect 3018 4132 3042 4166
rect 2960 4108 3042 4132
rect 3978 4166 4060 4190
rect 3978 4132 4002 4166
rect 4036 4132 4060 4166
rect 3978 4108 4060 4132
rect 4996 4166 5078 4190
rect 4996 4132 5020 4166
rect 5054 4132 5078 4166
rect 4996 4108 5078 4132
rect 6014 4166 6096 4190
rect 6014 4132 6038 4166
rect 6072 4132 6096 4166
rect 6014 4108 6096 4132
rect 7032 4166 7114 4190
rect 7032 4132 7056 4166
rect 7090 4132 7114 4166
rect 7032 4108 7114 4132
rect 8050 4166 8132 4190
rect 8050 4132 8074 4166
rect 8108 4132 8132 4166
rect 8050 4108 8132 4132
rect 9068 4166 9150 4190
rect 9068 4132 9092 4166
rect 9126 4132 9150 4166
rect 9068 4108 9150 4132
rect 10086 4166 10168 4190
rect 10086 4132 10110 4166
rect 10144 4132 10168 4166
rect 10086 4108 10168 4132
rect 11104 4166 11186 4190
rect 11104 4132 11128 4166
rect 11162 4132 11186 4166
rect 13530 4134 13564 4150
rect 14548 4726 14582 4742
rect 14548 4134 14582 4150
rect 15566 4726 15600 4742
rect 15566 4134 15600 4150
rect 16584 4726 16618 4742
rect 16584 4134 16618 4150
rect 17602 4726 17636 4742
rect 17602 4134 17636 4150
rect 18620 4726 18654 4742
rect 18620 4134 18654 4150
rect 19638 4726 19672 4742
rect 19638 4134 19672 4150
rect 20656 4726 20690 4742
rect 20656 4134 20690 4150
rect 21674 4726 21708 4742
rect 21674 4134 21708 4150
rect 22692 4726 22726 4742
rect 22692 4134 22726 4150
rect 23710 4726 23744 4742
rect 23710 4134 23744 4150
rect 24728 4726 24762 4742
rect 24728 4134 24762 4150
rect 25746 4726 25780 4742
rect 25746 4134 25780 4150
rect 26764 4726 26798 4742
rect 26764 4134 26798 4150
rect 27782 4726 27816 4742
rect 27782 4134 27816 4150
rect 28800 4726 28834 4742
rect 28800 4134 28834 4150
rect 29818 4726 29852 4742
rect 29818 4134 29852 4150
rect 30836 4726 30870 4742
rect 30836 4134 30870 4150
rect 31854 4726 31888 4742
rect 31854 4134 31888 4150
rect 32872 4726 32906 4742
rect 32872 4134 32906 4150
rect 33890 4726 33924 4742
rect 33890 4134 33924 4150
rect 11104 4108 11186 4132
rect 22180 4100 22240 4102
rect 24224 4100 24284 4104
rect 27262 4100 27322 4104
rect 13762 4066 13778 4100
rect 14334 4066 14350 4100
rect 14780 4066 14796 4100
rect 15352 4066 15368 4100
rect 15798 4066 15814 4100
rect 16370 4066 16386 4100
rect 16816 4066 16832 4100
rect 17388 4066 17404 4100
rect 17834 4066 17850 4100
rect 18406 4066 18422 4100
rect 18852 4066 18868 4100
rect 19424 4066 19440 4100
rect 19870 4066 19886 4100
rect 20442 4066 20458 4100
rect 20888 4066 20904 4100
rect 21460 4066 21476 4100
rect 21906 4066 21922 4100
rect 22478 4066 22494 4100
rect 22924 4066 22940 4100
rect 23496 4066 23512 4100
rect 23942 4066 23958 4100
rect 24514 4066 24530 4100
rect 24960 4066 24976 4100
rect 25532 4066 25548 4100
rect 25978 4066 25994 4100
rect 26550 4066 26566 4100
rect 26996 4066 27012 4100
rect 27568 4066 27584 4100
rect 28014 4066 28030 4100
rect 28586 4066 28602 4100
rect 29032 4066 29048 4100
rect 29604 4066 29620 4100
rect 30050 4066 30066 4100
rect 30622 4066 30638 4100
rect 31068 4066 31084 4100
rect 31640 4066 31656 4100
rect 32086 4066 32102 4100
rect 32658 4066 32674 4100
rect 33104 4066 33120 4100
rect 33676 4066 33692 4100
rect 674 3922 690 3956
rect 1246 3922 1262 3956
rect 1692 3922 1708 3956
rect 2264 3922 2280 3956
rect 2710 3922 2726 3956
rect 3282 3922 3298 3956
rect 3728 3922 3744 3956
rect 4300 3922 4316 3956
rect 4746 3922 4762 3956
rect 5318 3922 5334 3956
rect 5764 3922 5780 3956
rect 6336 3922 6352 3956
rect 6782 3922 6798 3956
rect 7354 3922 7370 3956
rect 7800 3922 7816 3956
rect 8372 3922 8388 3956
rect 8818 3922 8834 3956
rect 9390 3922 9406 3956
rect 9836 3922 9852 3956
rect 10408 3922 10424 3956
rect 10854 3922 10870 3956
rect 11426 3922 11442 3956
rect 442 3872 476 3888
rect 442 3280 476 3296
rect 1460 3872 1494 3888
rect 1460 3280 1494 3296
rect 2478 3872 2512 3888
rect 2478 3280 2512 3296
rect 3496 3872 3530 3888
rect 3496 3280 3530 3296
rect 4514 3872 4548 3888
rect 4514 3280 4548 3296
rect 5532 3872 5566 3888
rect 5532 3280 5566 3296
rect 6550 3872 6584 3888
rect 6550 3280 6584 3296
rect 7568 3872 7602 3888
rect 7568 3280 7602 3296
rect 8586 3872 8620 3888
rect 8586 3280 8620 3296
rect 9604 3872 9638 3888
rect 9604 3280 9638 3296
rect 10622 3872 10656 3888
rect 10622 3280 10656 3296
rect 11640 3872 11674 3888
rect 14024 3850 14106 3874
rect 14024 3816 14048 3850
rect 14082 3816 14106 3850
rect 14024 3792 14106 3816
rect 15042 3850 15124 3874
rect 15042 3816 15066 3850
rect 15100 3816 15124 3850
rect 15042 3792 15124 3816
rect 16060 3850 16142 3874
rect 16060 3816 16084 3850
rect 16118 3816 16142 3850
rect 16060 3792 16142 3816
rect 17078 3850 17160 3874
rect 17078 3816 17102 3850
rect 17136 3816 17160 3850
rect 17078 3792 17160 3816
rect 18096 3850 18178 3874
rect 18096 3816 18120 3850
rect 18154 3816 18178 3850
rect 18096 3792 18178 3816
rect 19114 3850 19196 3874
rect 19114 3816 19138 3850
rect 19172 3816 19196 3850
rect 19114 3792 19196 3816
rect 20132 3850 20214 3874
rect 20132 3816 20156 3850
rect 20190 3816 20214 3850
rect 20132 3792 20214 3816
rect 21150 3850 21232 3874
rect 21150 3816 21174 3850
rect 21208 3816 21232 3850
rect 21150 3792 21232 3816
rect 22168 3850 22250 3874
rect 22168 3816 22192 3850
rect 22226 3816 22250 3850
rect 22168 3792 22250 3816
rect 23186 3850 23268 3874
rect 23186 3816 23210 3850
rect 23244 3816 23268 3850
rect 23186 3792 23268 3816
rect 24204 3850 24286 3874
rect 24204 3816 24228 3850
rect 24262 3816 24286 3850
rect 24204 3792 24286 3816
rect 25222 3850 25304 3874
rect 25222 3816 25246 3850
rect 25280 3816 25304 3850
rect 25222 3792 25304 3816
rect 26240 3850 26322 3874
rect 26240 3816 26264 3850
rect 26298 3816 26322 3850
rect 26240 3792 26322 3816
rect 27258 3850 27340 3874
rect 27258 3816 27282 3850
rect 27316 3816 27340 3850
rect 27258 3792 27340 3816
rect 28276 3850 28358 3874
rect 28276 3816 28300 3850
rect 28334 3816 28358 3850
rect 28276 3792 28358 3816
rect 29294 3850 29376 3874
rect 29294 3816 29318 3850
rect 29352 3816 29376 3850
rect 29294 3792 29376 3816
rect 30312 3850 30394 3874
rect 30312 3816 30336 3850
rect 30370 3816 30394 3850
rect 30312 3792 30394 3816
rect 31330 3850 31412 3874
rect 31330 3816 31354 3850
rect 31388 3816 31412 3850
rect 31330 3792 31412 3816
rect 32348 3850 32430 3874
rect 32348 3816 32372 3850
rect 32406 3816 32430 3850
rect 32348 3792 32430 3816
rect 33366 3850 33448 3874
rect 33366 3816 33390 3850
rect 33424 3816 33448 3850
rect 33366 3792 33448 3816
rect 13762 3544 13778 3578
rect 14334 3544 14350 3578
rect 14780 3544 14796 3578
rect 15352 3544 15368 3578
rect 15798 3544 15814 3578
rect 16370 3544 16386 3578
rect 16816 3544 16832 3578
rect 17388 3544 17404 3578
rect 17834 3544 17850 3578
rect 18406 3544 18422 3578
rect 18852 3544 18868 3578
rect 19424 3544 19440 3578
rect 19870 3544 19886 3578
rect 20442 3544 20458 3578
rect 20888 3544 20904 3578
rect 21460 3544 21476 3578
rect 21906 3544 21922 3578
rect 22478 3544 22494 3578
rect 22924 3544 22940 3578
rect 23496 3544 23512 3578
rect 23942 3544 23958 3578
rect 24514 3544 24530 3578
rect 24960 3544 24976 3578
rect 25532 3544 25548 3578
rect 25978 3544 25994 3578
rect 26550 3544 26566 3578
rect 26996 3544 27012 3578
rect 27568 3544 27584 3578
rect 28014 3544 28030 3578
rect 28586 3544 28602 3578
rect 29032 3544 29048 3578
rect 29604 3544 29620 3578
rect 30050 3544 30066 3578
rect 30622 3544 30638 3578
rect 31068 3544 31084 3578
rect 31640 3544 31656 3578
rect 32086 3544 32102 3578
rect 32658 3544 32674 3578
rect 33104 3544 33120 3578
rect 33676 3544 33692 3578
rect 17084 3542 17144 3544
rect 11640 3280 11674 3296
rect 13530 3494 13564 3510
rect 674 3212 690 3246
rect 1246 3212 1262 3246
rect 1692 3212 1708 3246
rect 2264 3212 2280 3246
rect 2710 3212 2726 3246
rect 3282 3212 3298 3246
rect 3728 3212 3744 3246
rect 4300 3212 4316 3246
rect 4746 3212 4762 3246
rect 5318 3212 5334 3246
rect 5764 3212 5780 3246
rect 6336 3212 6352 3246
rect 6782 3212 6798 3246
rect 7354 3212 7370 3246
rect 7800 3212 7816 3246
rect 8372 3212 8388 3246
rect 8818 3212 8834 3246
rect 9390 3212 9406 3246
rect 9836 3212 9852 3246
rect 10408 3212 10424 3246
rect 10854 3212 10870 3246
rect 11426 3212 11442 3246
rect 924 3060 1006 3084
rect 924 3026 948 3060
rect 982 3026 1006 3060
rect 924 3002 1006 3026
rect 1942 3060 2024 3084
rect 1942 3026 1966 3060
rect 2000 3026 2024 3060
rect 1942 3002 2024 3026
rect 2960 3060 3042 3084
rect 2960 3026 2984 3060
rect 3018 3026 3042 3060
rect 2960 3002 3042 3026
rect 3978 3060 4060 3084
rect 3978 3026 4002 3060
rect 4036 3026 4060 3060
rect 3978 3002 4060 3026
rect 4996 3060 5078 3084
rect 4996 3026 5020 3060
rect 5054 3026 5078 3060
rect 4996 3002 5078 3026
rect 6014 3060 6096 3084
rect 6014 3026 6038 3060
rect 6072 3026 6096 3060
rect 6014 3002 6096 3026
rect 7032 3060 7114 3084
rect 7032 3026 7056 3060
rect 7090 3026 7114 3060
rect 7032 3002 7114 3026
rect 8050 3060 8132 3084
rect 8050 3026 8074 3060
rect 8108 3026 8132 3060
rect 8050 3002 8132 3026
rect 9068 3060 9150 3084
rect 9068 3026 9092 3060
rect 9126 3026 9150 3060
rect 9068 3002 9150 3026
rect 10086 3060 10168 3084
rect 10086 3026 10110 3060
rect 10144 3026 10168 3060
rect 10086 3002 10168 3026
rect 11104 3060 11186 3084
rect 11104 3026 11128 3060
rect 11162 3026 11186 3060
rect 11104 3002 11186 3026
rect 13530 2902 13564 2918
rect 14548 3494 14582 3510
rect 14548 2902 14582 2918
rect 15566 3494 15600 3510
rect 15566 2902 15600 2918
rect 16584 3494 16618 3510
rect 16584 2902 16618 2918
rect 17602 3494 17636 3510
rect 17602 2902 17636 2918
rect 18620 3494 18654 3510
rect 18620 2902 18654 2918
rect 19638 3494 19672 3510
rect 19638 2902 19672 2918
rect 20656 3494 20690 3510
rect 20656 2902 20690 2918
rect 21674 3494 21708 3510
rect 21674 2902 21708 2918
rect 22692 3494 22726 3510
rect 22692 2902 22726 2918
rect 23710 3494 23744 3510
rect 23710 2902 23744 2918
rect 24728 3494 24762 3510
rect 24728 2902 24762 2918
rect 25746 3494 25780 3510
rect 25746 2902 25780 2918
rect 26764 3494 26798 3510
rect 26764 2902 26798 2918
rect 27782 3494 27816 3510
rect 27782 2902 27816 2918
rect 28800 3494 28834 3510
rect 28800 2902 28834 2918
rect 29818 3494 29852 3510
rect 29818 2902 29852 2918
rect 30836 3494 30870 3510
rect 30836 2902 30870 2918
rect 31854 3494 31888 3510
rect 31854 2902 31888 2918
rect 32872 3494 32906 3510
rect 32872 2902 32906 2918
rect 33890 3494 33924 3510
rect 33890 2902 33924 2918
rect 21156 2868 21216 2878
rect 674 2810 690 2844
rect 1246 2810 1262 2844
rect 1692 2810 1708 2844
rect 2264 2810 2280 2844
rect 2710 2810 2726 2844
rect 3282 2810 3298 2844
rect 3728 2810 3744 2844
rect 4300 2810 4316 2844
rect 4746 2810 4762 2844
rect 5318 2810 5334 2844
rect 5764 2810 5780 2844
rect 6336 2810 6352 2844
rect 6782 2810 6798 2844
rect 7354 2810 7370 2844
rect 7800 2810 7816 2844
rect 8372 2810 8388 2844
rect 8818 2810 8834 2844
rect 9390 2810 9406 2844
rect 9836 2810 9852 2844
rect 10408 2810 10424 2844
rect 10854 2810 10870 2844
rect 11426 2810 11442 2844
rect 13762 2834 13778 2868
rect 14334 2834 14350 2868
rect 14780 2834 14796 2868
rect 15352 2834 15368 2868
rect 15798 2834 15814 2868
rect 16370 2834 16386 2868
rect 16816 2834 16832 2868
rect 17388 2834 17404 2868
rect 17834 2834 17850 2868
rect 18406 2834 18422 2868
rect 18852 2834 18868 2868
rect 19424 2834 19440 2868
rect 19870 2834 19886 2868
rect 20442 2834 20458 2868
rect 20888 2834 20904 2868
rect 21460 2834 21476 2868
rect 21906 2834 21922 2868
rect 22478 2834 22494 2868
rect 22924 2834 22940 2868
rect 23496 2834 23512 2868
rect 23942 2834 23958 2868
rect 24514 2834 24530 2868
rect 24960 2834 24976 2868
rect 25532 2834 25548 2868
rect 25978 2834 25994 2868
rect 26550 2834 26566 2868
rect 26996 2834 27012 2868
rect 27568 2834 27584 2868
rect 28014 2834 28030 2868
rect 28586 2834 28602 2868
rect 29032 2834 29048 2868
rect 29604 2834 29620 2868
rect 30050 2834 30066 2868
rect 30622 2834 30638 2868
rect 31068 2834 31084 2868
rect 31640 2834 31656 2868
rect 32086 2834 32102 2868
rect 32658 2834 32674 2868
rect 33104 2834 33120 2868
rect 33676 2834 33692 2868
rect 442 2760 476 2776
rect 442 2168 476 2184
rect 1460 2760 1494 2776
rect 1460 2168 1494 2184
rect 2478 2760 2512 2776
rect 2478 2168 2512 2184
rect 3496 2760 3530 2776
rect 3496 2168 3530 2184
rect 4514 2760 4548 2776
rect 4514 2168 4548 2184
rect 5532 2760 5566 2776
rect 5532 2168 5566 2184
rect 6550 2760 6584 2776
rect 6550 2168 6584 2184
rect 7568 2760 7602 2776
rect 7568 2168 7602 2184
rect 8586 2760 8620 2776
rect 8586 2168 8620 2184
rect 9604 2760 9638 2776
rect 9604 2168 9638 2184
rect 10622 2760 10656 2776
rect 10622 2168 10656 2184
rect 11640 2760 11674 2776
rect 14024 2614 14106 2638
rect 14024 2580 14048 2614
rect 14082 2580 14106 2614
rect 14024 2556 14106 2580
rect 15042 2614 15124 2638
rect 15042 2580 15066 2614
rect 15100 2580 15124 2614
rect 15042 2556 15124 2580
rect 16060 2614 16142 2638
rect 16060 2580 16084 2614
rect 16118 2580 16142 2614
rect 16060 2556 16142 2580
rect 17078 2614 17160 2638
rect 17078 2580 17102 2614
rect 17136 2580 17160 2614
rect 17078 2556 17160 2580
rect 18096 2614 18178 2638
rect 18096 2580 18120 2614
rect 18154 2580 18178 2614
rect 18096 2556 18178 2580
rect 19114 2614 19196 2638
rect 19114 2580 19138 2614
rect 19172 2580 19196 2614
rect 19114 2556 19196 2580
rect 20132 2614 20214 2638
rect 20132 2580 20156 2614
rect 20190 2580 20214 2614
rect 20132 2556 20214 2580
rect 21150 2614 21232 2638
rect 21150 2580 21174 2614
rect 21208 2580 21232 2614
rect 21150 2556 21232 2580
rect 22168 2614 22250 2638
rect 22168 2580 22192 2614
rect 22226 2580 22250 2614
rect 22168 2556 22250 2580
rect 23186 2614 23268 2638
rect 23186 2580 23210 2614
rect 23244 2580 23268 2614
rect 23186 2556 23268 2580
rect 24204 2614 24286 2638
rect 24204 2580 24228 2614
rect 24262 2580 24286 2614
rect 24204 2556 24286 2580
rect 25222 2614 25304 2638
rect 25222 2580 25246 2614
rect 25280 2580 25304 2614
rect 25222 2556 25304 2580
rect 26240 2614 26322 2638
rect 26240 2580 26264 2614
rect 26298 2580 26322 2614
rect 26240 2556 26322 2580
rect 27258 2614 27340 2638
rect 27258 2580 27282 2614
rect 27316 2580 27340 2614
rect 27258 2556 27340 2580
rect 28276 2614 28358 2638
rect 28276 2580 28300 2614
rect 28334 2580 28358 2614
rect 28276 2556 28358 2580
rect 29294 2614 29376 2638
rect 29294 2580 29318 2614
rect 29352 2580 29376 2614
rect 29294 2556 29376 2580
rect 30312 2614 30394 2638
rect 30312 2580 30336 2614
rect 30370 2580 30394 2614
rect 30312 2556 30394 2580
rect 31330 2614 31412 2638
rect 31330 2580 31354 2614
rect 31388 2580 31412 2614
rect 31330 2556 31412 2580
rect 32348 2614 32430 2638
rect 32348 2580 32372 2614
rect 32406 2580 32430 2614
rect 32348 2556 32430 2580
rect 33366 2614 33448 2638
rect 33366 2580 33390 2614
rect 33424 2580 33448 2614
rect 33366 2556 33448 2580
rect 13762 2310 13778 2344
rect 14334 2310 14350 2344
rect 14780 2310 14796 2344
rect 15352 2310 15368 2344
rect 15798 2310 15814 2344
rect 16370 2310 16386 2344
rect 16816 2310 16832 2344
rect 17388 2310 17404 2344
rect 17834 2310 17850 2344
rect 18406 2310 18422 2344
rect 18852 2310 18868 2344
rect 19424 2310 19440 2344
rect 19870 2310 19886 2344
rect 20442 2310 20458 2344
rect 20888 2310 20904 2344
rect 21460 2310 21476 2344
rect 21906 2310 21922 2344
rect 22478 2310 22494 2344
rect 22924 2310 22940 2344
rect 23496 2310 23512 2344
rect 23942 2310 23958 2344
rect 24514 2310 24530 2344
rect 24960 2310 24976 2344
rect 25532 2310 25548 2344
rect 25978 2310 25994 2344
rect 26550 2310 26566 2344
rect 26996 2310 27012 2344
rect 27568 2310 27584 2344
rect 28014 2310 28030 2344
rect 28586 2310 28602 2344
rect 29032 2310 29048 2344
rect 29604 2310 29620 2344
rect 30050 2310 30066 2344
rect 30622 2310 30638 2344
rect 31068 2310 31084 2344
rect 31640 2310 31656 2344
rect 32086 2310 32102 2344
rect 32658 2310 32674 2344
rect 33104 2310 33120 2344
rect 33676 2310 33692 2344
rect 17070 2308 17130 2310
rect 11640 2168 11674 2184
rect 13530 2260 13564 2276
rect 674 2100 690 2134
rect 1246 2100 1262 2134
rect 1692 2100 1708 2134
rect 2264 2100 2280 2134
rect 2710 2100 2726 2134
rect 3282 2100 3298 2134
rect 3728 2100 3744 2134
rect 4300 2100 4316 2134
rect 4746 2100 4762 2134
rect 5318 2100 5334 2134
rect 5764 2100 5780 2134
rect 6336 2100 6352 2134
rect 6782 2100 6798 2134
rect 7354 2100 7370 2134
rect 7800 2100 7816 2134
rect 8372 2100 8388 2134
rect 8818 2100 8834 2134
rect 9390 2100 9406 2134
rect 9836 2100 9852 2134
rect 10408 2100 10424 2134
rect 10854 2100 10870 2134
rect 11426 2100 11442 2134
rect 924 1718 1006 1742
rect 924 1684 948 1718
rect 982 1684 1006 1718
rect 924 1660 1006 1684
rect 1942 1718 2024 1742
rect 1942 1684 1966 1718
rect 2000 1684 2024 1718
rect 1942 1660 2024 1684
rect 2960 1718 3042 1742
rect 2960 1684 2984 1718
rect 3018 1684 3042 1718
rect 2960 1660 3042 1684
rect 3978 1718 4060 1742
rect 3978 1684 4002 1718
rect 4036 1684 4060 1718
rect 3978 1660 4060 1684
rect 4996 1718 5078 1742
rect 4996 1684 5020 1718
rect 5054 1684 5078 1718
rect 4996 1660 5078 1684
rect 6014 1718 6096 1742
rect 6014 1684 6038 1718
rect 6072 1684 6096 1718
rect 6014 1660 6096 1684
rect 7032 1718 7114 1742
rect 7032 1684 7056 1718
rect 7090 1684 7114 1718
rect 7032 1660 7114 1684
rect 8050 1718 8132 1742
rect 8050 1684 8074 1718
rect 8108 1684 8132 1718
rect 8050 1660 8132 1684
rect 9068 1718 9150 1742
rect 9068 1684 9092 1718
rect 9126 1684 9150 1718
rect 9068 1660 9150 1684
rect 10086 1718 10168 1742
rect 10086 1684 10110 1718
rect 10144 1684 10168 1718
rect 10086 1660 10168 1684
rect 11104 1718 11186 1742
rect 11104 1684 11128 1718
rect 11162 1684 11186 1718
rect 11104 1660 11186 1684
rect 13530 1668 13564 1684
rect 14548 2260 14582 2276
rect 14548 1668 14582 1684
rect 15566 2260 15600 2276
rect 15566 1668 15600 1684
rect 16584 2260 16618 2276
rect 16584 1668 16618 1684
rect 17602 2260 17636 2276
rect 17602 1668 17636 1684
rect 18620 2260 18654 2276
rect 18620 1668 18654 1684
rect 19638 2260 19672 2276
rect 19638 1668 19672 1684
rect 20656 2260 20690 2276
rect 20656 1668 20690 1684
rect 21674 2260 21708 2276
rect 21674 1668 21708 1684
rect 22692 2260 22726 2276
rect 22692 1668 22726 1684
rect 23710 2260 23744 2276
rect 23710 1668 23744 1684
rect 24728 2260 24762 2276
rect 24728 1668 24762 1684
rect 25746 2260 25780 2276
rect 25746 1668 25780 1684
rect 26764 2260 26798 2276
rect 26764 1668 26798 1684
rect 27782 2260 27816 2276
rect 27782 1668 27816 1684
rect 28800 2260 28834 2276
rect 28800 1668 28834 1684
rect 29818 2260 29852 2276
rect 29818 1668 29852 1684
rect 30836 2260 30870 2276
rect 30836 1668 30870 1684
rect 31854 2260 31888 2276
rect 31854 1668 31888 1684
rect 32872 2260 32906 2276
rect 32872 1668 32906 1684
rect 33890 2260 33924 2276
rect 33890 1668 33924 1684
rect 15038 1634 15098 1636
rect 21150 1634 21210 1636
rect 23184 1634 23244 1636
rect 27250 1634 27310 1640
rect 31326 1634 31386 1636
rect 32342 1634 32402 1636
rect 13762 1600 13778 1634
rect 14334 1600 14350 1634
rect 14780 1600 14796 1634
rect 15352 1600 15368 1634
rect 15798 1600 15814 1634
rect 16370 1600 16386 1634
rect 16816 1600 16832 1634
rect 17388 1600 17404 1634
rect 17834 1600 17850 1634
rect 18406 1600 18422 1634
rect 18852 1600 18868 1634
rect 19424 1600 19440 1634
rect 19870 1600 19886 1634
rect 20442 1600 20458 1634
rect 20888 1600 20904 1634
rect 21460 1600 21476 1634
rect 21906 1600 21922 1634
rect 22478 1600 22494 1634
rect 22924 1600 22940 1634
rect 23496 1600 23512 1634
rect 23942 1600 23958 1634
rect 24514 1600 24530 1634
rect 24960 1600 24976 1634
rect 25532 1600 25548 1634
rect 25978 1600 25994 1634
rect 26550 1600 26566 1634
rect 26996 1600 27012 1634
rect 27568 1600 27584 1634
rect 28014 1600 28030 1634
rect 28586 1600 28602 1634
rect 29032 1600 29048 1634
rect 29604 1600 29620 1634
rect 30050 1600 30066 1634
rect 30622 1600 30638 1634
rect 31068 1600 31084 1634
rect 31640 1600 31656 1634
rect 32086 1600 32102 1634
rect 32658 1600 32674 1634
rect 33104 1600 33120 1634
rect 33676 1600 33692 1634
rect 14036 1368 14118 1392
rect 14036 1334 14060 1368
rect 14094 1334 14118 1368
rect 14036 1310 14118 1334
rect 15054 1368 15136 1392
rect 15054 1334 15078 1368
rect 15112 1334 15136 1368
rect 15054 1310 15136 1334
rect 16072 1368 16154 1392
rect 16072 1334 16096 1368
rect 16130 1334 16154 1368
rect 16072 1310 16154 1334
rect 17090 1368 17172 1392
rect 17090 1334 17114 1368
rect 17148 1334 17172 1368
rect 17090 1310 17172 1334
rect 18108 1368 18190 1392
rect 18108 1334 18132 1368
rect 18166 1334 18190 1368
rect 18108 1310 18190 1334
rect 19126 1368 19208 1392
rect 19126 1334 19150 1368
rect 19184 1334 19208 1368
rect 19126 1310 19208 1334
rect 20144 1368 20226 1392
rect 20144 1334 20168 1368
rect 20202 1334 20226 1368
rect 20144 1310 20226 1334
rect 21162 1368 21244 1392
rect 21162 1334 21186 1368
rect 21220 1334 21244 1368
rect 21162 1310 21244 1334
rect 22180 1368 22262 1392
rect 22180 1334 22204 1368
rect 22238 1334 22262 1368
rect 22180 1310 22262 1334
rect 23198 1368 23280 1392
rect 23198 1334 23222 1368
rect 23256 1334 23280 1368
rect 23198 1310 23280 1334
rect 24216 1368 24298 1392
rect 24216 1334 24240 1368
rect 24274 1334 24298 1368
rect 24216 1310 24298 1334
rect 25234 1368 25316 1392
rect 25234 1334 25258 1368
rect 25292 1334 25316 1368
rect 25234 1310 25316 1334
rect 26252 1368 26334 1392
rect 26252 1334 26276 1368
rect 26310 1334 26334 1368
rect 26252 1310 26334 1334
rect 27270 1368 27352 1392
rect 27270 1334 27294 1368
rect 27328 1334 27352 1368
rect 27270 1310 27352 1334
rect 28288 1368 28370 1392
rect 28288 1334 28312 1368
rect 28346 1334 28370 1368
rect 28288 1310 28370 1334
rect 29306 1368 29388 1392
rect 29306 1334 29330 1368
rect 29364 1334 29388 1368
rect 29306 1310 29388 1334
rect 30324 1368 30406 1392
rect 30324 1334 30348 1368
rect 30382 1334 30406 1368
rect 30324 1310 30406 1334
rect 31342 1368 31424 1392
rect 31342 1334 31366 1368
rect 31400 1334 31424 1368
rect 31342 1310 31424 1334
rect 32360 1368 32442 1392
rect 32360 1334 32384 1368
rect 32418 1334 32442 1368
rect 32360 1310 32442 1334
rect 33378 1368 33460 1392
rect 33378 1334 33402 1368
rect 33436 1334 33460 1368
rect 33378 1310 33460 1334
rect 1132 1268 1148 1302
rect 1704 1268 1720 1302
rect 2150 1268 2166 1302
rect 2722 1268 2738 1302
rect 3168 1268 3184 1302
rect 3740 1268 3756 1302
rect 4186 1268 4202 1302
rect 4758 1268 4774 1302
rect 5204 1268 5220 1302
rect 5776 1268 5792 1302
rect 6222 1268 6238 1302
rect 6794 1268 6810 1302
rect 7240 1268 7256 1302
rect 7812 1268 7828 1302
rect 8258 1268 8274 1302
rect 8830 1268 8846 1302
rect 9276 1268 9292 1302
rect 9848 1268 9864 1302
rect 10294 1268 10310 1302
rect 10866 1268 10882 1302
rect 900 1218 934 1234
rect 900 626 934 642
rect 1918 1218 1952 1234
rect 1918 626 1952 642
rect 2936 1218 2970 1234
rect 2936 626 2970 642
rect 3954 1218 3988 1234
rect 3954 626 3988 642
rect 4972 1218 5006 1234
rect 4972 626 5006 642
rect 5990 1218 6024 1234
rect 5990 626 6024 642
rect 7008 1218 7042 1234
rect 7008 626 7042 642
rect 8026 1218 8060 1234
rect 8026 626 8060 642
rect 9044 1218 9078 1234
rect 9044 626 9078 642
rect 10062 1218 10096 1234
rect 10062 626 10096 642
rect 11080 1218 11114 1234
rect 13762 1078 13778 1112
rect 14334 1078 14350 1112
rect 14780 1078 14796 1112
rect 15352 1078 15368 1112
rect 15798 1078 15814 1112
rect 16370 1078 16386 1112
rect 16816 1078 16832 1112
rect 17388 1078 17404 1112
rect 17834 1078 17850 1112
rect 18406 1078 18422 1112
rect 18852 1078 18868 1112
rect 19424 1078 19440 1112
rect 19870 1078 19886 1112
rect 20442 1078 20458 1112
rect 20888 1078 20904 1112
rect 21460 1078 21476 1112
rect 21906 1078 21922 1112
rect 22478 1078 22494 1112
rect 22924 1078 22940 1112
rect 23496 1078 23512 1112
rect 23942 1078 23958 1112
rect 24514 1078 24530 1112
rect 24960 1078 24976 1112
rect 25532 1078 25548 1112
rect 25978 1078 25994 1112
rect 26550 1078 26566 1112
rect 26996 1078 27012 1112
rect 27568 1078 27584 1112
rect 28014 1078 28030 1112
rect 28586 1078 28602 1112
rect 29032 1078 29048 1112
rect 29604 1078 29620 1112
rect 30050 1078 30066 1112
rect 30622 1078 30638 1112
rect 31068 1078 31084 1112
rect 31640 1078 31656 1112
rect 32086 1078 32102 1112
rect 32658 1078 32674 1112
rect 33104 1078 33120 1112
rect 33676 1078 33692 1112
rect 11080 626 11114 642
rect 13530 1028 13564 1044
rect 1132 558 1148 592
rect 1704 558 1720 592
rect 2150 558 2166 592
rect 2722 558 2738 592
rect 3168 558 3184 592
rect 3740 558 3756 592
rect 4186 558 4202 592
rect 4758 558 4774 592
rect 5204 558 5220 592
rect 5776 558 5792 592
rect 6222 558 6238 592
rect 6794 558 6810 592
rect 7240 558 7256 592
rect 7812 558 7828 592
rect 8258 558 8274 592
rect 8830 558 8846 592
rect 9276 558 9292 592
rect 9848 558 9864 592
rect 10294 558 10310 592
rect 10866 558 10882 592
rect 13530 436 13564 452
rect 14548 1028 14582 1044
rect 14548 436 14582 452
rect 15566 1028 15600 1044
rect 15566 436 15600 452
rect 16584 1028 16618 1044
rect 16584 436 16618 452
rect 17602 1028 17636 1044
rect 17602 436 17636 452
rect 18620 1028 18654 1044
rect 18620 436 18654 452
rect 19638 1028 19672 1044
rect 19638 436 19672 452
rect 20656 1028 20690 1044
rect 20656 436 20690 452
rect 21674 1028 21708 1044
rect 21674 436 21708 452
rect 22692 1028 22726 1044
rect 22692 436 22726 452
rect 23710 1028 23744 1044
rect 23710 436 23744 452
rect 24728 1028 24762 1044
rect 24728 436 24762 452
rect 25746 1028 25780 1044
rect 25746 436 25780 452
rect 26764 1028 26798 1044
rect 26764 436 26798 452
rect 27782 1028 27816 1044
rect 27782 436 27816 452
rect 28800 1028 28834 1044
rect 28800 436 28834 452
rect 29818 1028 29852 1044
rect 29818 436 29852 452
rect 30836 1028 30870 1044
rect 30836 436 30870 452
rect 31854 1028 31888 1044
rect 31854 436 31888 452
rect 32872 1028 32906 1044
rect 32872 436 32906 452
rect 33890 1028 33924 1044
rect 33890 436 33924 452
rect -1188 362 -1114 396
rect -914 362 -838 396
rect 13762 368 13778 402
rect 14334 368 14350 402
rect 14780 368 14796 402
rect 15352 368 15368 402
rect 15798 368 15814 402
rect 16370 368 16386 402
rect 16816 368 16832 402
rect 17388 368 17404 402
rect 17834 368 17850 402
rect 18406 368 18422 402
rect 18852 368 18868 402
rect 19424 368 19440 402
rect 19870 368 19886 402
rect 20442 368 20458 402
rect 20888 368 20904 402
rect 21460 368 21476 402
rect 21906 368 21922 402
rect 22478 368 22494 402
rect 22924 368 22940 402
rect 23496 368 23512 402
rect 23942 368 23958 402
rect 24514 368 24530 402
rect 24960 368 24976 402
rect 25532 368 25548 402
rect 25978 368 25994 402
rect 26550 368 26566 402
rect 26996 368 27012 402
rect 27568 368 27584 402
rect 28014 368 28030 402
rect 28586 368 28602 402
rect 29032 368 29048 402
rect 29604 368 29620 402
rect 30050 368 30066 402
rect 30622 368 30638 402
rect 31068 368 31084 402
rect 31640 368 31656 402
rect 32086 368 32102 402
rect 32658 368 32674 402
rect 33104 368 33120 402
rect 33676 368 33692 402
rect -1188 360 -1154 362
rect -872 358 -838 362
rect -1046 240 -1030 274
rect -996 240 -980 274
rect -1074 190 -1040 206
rect -1074 68 -1040 84
rect -986 190 -952 206
rect -986 68 -952 84
rect 734 272 816 296
rect 734 238 758 272
rect 792 238 816 272
rect 734 214 816 238
rect 1752 272 1834 296
rect 1752 238 1776 272
rect 1810 238 1834 272
rect 1752 214 1834 238
rect 2770 272 2852 296
rect 2770 238 2794 272
rect 2828 238 2852 272
rect 2770 214 2852 238
rect 3788 272 3870 296
rect 3788 238 3812 272
rect 3846 238 3870 272
rect 3788 214 3870 238
rect 4806 272 4888 296
rect 4806 238 4830 272
rect 4864 238 4888 272
rect 4806 214 4888 238
rect 5824 272 5906 296
rect 5824 238 5848 272
rect 5882 238 5906 272
rect 5824 214 5906 238
rect 6842 272 6924 296
rect 6842 238 6866 272
rect 6900 238 6924 272
rect 6842 214 6924 238
rect 7860 272 7942 296
rect 7860 238 7884 272
rect 7918 238 7942 272
rect 7860 214 7942 238
rect 8878 272 8960 296
rect 8878 238 8902 272
rect 8936 238 8960 272
rect 8878 214 8960 238
rect 9896 272 9978 296
rect 9896 238 9920 272
rect 9954 238 9978 272
rect 9896 214 9978 238
rect 10914 272 10996 296
rect 10914 238 10938 272
rect 10972 238 10996 272
rect 10914 214 10996 238
rect 14024 190 14106 214
rect 14024 156 14048 190
rect 14082 156 14106 190
rect 14024 132 14106 156
rect 15042 190 15124 214
rect 15042 156 15066 190
rect 15100 156 15124 190
rect 15042 132 15124 156
rect 16060 190 16142 214
rect 16060 156 16084 190
rect 16118 156 16142 190
rect 16060 132 16142 156
rect 17078 190 17160 214
rect 17078 156 17102 190
rect 17136 156 17160 190
rect 17078 132 17160 156
rect 18096 190 18178 214
rect 18096 156 18120 190
rect 18154 156 18178 190
rect 18096 132 18178 156
rect 19114 190 19196 214
rect 19114 156 19138 190
rect 19172 156 19196 190
rect 19114 132 19196 156
rect 20132 190 20214 214
rect 20132 156 20156 190
rect 20190 156 20214 190
rect 20132 132 20214 156
rect 21150 190 21232 214
rect 21150 156 21174 190
rect 21208 156 21232 190
rect 21150 132 21232 156
rect 22168 190 22250 214
rect 22168 156 22192 190
rect 22226 156 22250 190
rect 22168 132 22250 156
rect 23186 190 23268 214
rect 23186 156 23210 190
rect 23244 156 23268 190
rect 23186 132 23268 156
rect 24204 190 24286 214
rect 24204 156 24228 190
rect 24262 156 24286 190
rect 24204 132 24286 156
rect 25222 190 25304 214
rect 25222 156 25246 190
rect 25280 156 25304 190
rect 25222 132 25304 156
rect 26240 190 26322 214
rect 26240 156 26264 190
rect 26298 156 26322 190
rect 26240 132 26322 156
rect 27258 190 27340 214
rect 27258 156 27282 190
rect 27316 156 27340 190
rect 27258 132 27340 156
rect 28276 190 28358 214
rect 28276 156 28300 190
rect 28334 156 28358 190
rect 28276 132 28358 156
rect 29294 190 29376 214
rect 29294 156 29318 190
rect 29352 156 29376 190
rect 29294 132 29376 156
rect 30312 190 30394 214
rect 30312 156 30336 190
rect 30370 156 30394 190
rect 30312 132 30394 156
rect 31330 190 31412 214
rect 31330 156 31354 190
rect 31388 156 31412 190
rect 31330 132 31412 156
rect 32348 190 32430 214
rect 32348 156 32372 190
rect 32406 156 32430 190
rect 32348 132 32430 156
rect 33366 190 33448 214
rect 33366 156 33390 190
rect 33424 156 33448 190
rect 33366 132 33448 156
rect -1046 0 -1030 34
rect -996 0 -980 34
rect -1188 -102 -1154 -100
rect 39628 15030 39728 15192
rect 76772 15030 76872 15192
rect 55036 14586 55118 14610
rect 55036 14552 55060 14586
rect 55094 14552 55118 14586
rect 55036 14528 55118 14552
rect 56054 14586 56136 14610
rect 56054 14552 56078 14586
rect 56112 14552 56136 14586
rect 56054 14528 56136 14552
rect 57072 14586 57154 14610
rect 57072 14552 57096 14586
rect 57130 14552 57154 14586
rect 57072 14528 57154 14552
rect 58090 14586 58172 14610
rect 58090 14552 58114 14586
rect 58148 14552 58172 14586
rect 58090 14528 58172 14552
rect 59108 14586 59190 14610
rect 59108 14552 59132 14586
rect 59166 14552 59190 14586
rect 59108 14528 59190 14552
rect 60126 14586 60208 14610
rect 60126 14552 60150 14586
rect 60184 14552 60208 14586
rect 60126 14528 60208 14552
rect 61144 14586 61226 14610
rect 61144 14552 61168 14586
rect 61202 14552 61226 14586
rect 61144 14528 61226 14552
rect 62162 14586 62244 14610
rect 62162 14552 62186 14586
rect 62220 14552 62244 14586
rect 62162 14528 62244 14552
rect 63180 14586 63262 14610
rect 63180 14552 63204 14586
rect 63238 14552 63262 14586
rect 63180 14528 63262 14552
rect 64198 14586 64280 14610
rect 64198 14552 64222 14586
rect 64256 14552 64280 14586
rect 64198 14528 64280 14552
rect 65216 14586 65298 14610
rect 65216 14552 65240 14586
rect 65274 14552 65298 14586
rect 65216 14528 65298 14552
rect 66234 14586 66316 14610
rect 66234 14552 66258 14586
rect 66292 14552 66316 14586
rect 66234 14528 66316 14552
rect 67252 14586 67334 14610
rect 67252 14552 67276 14586
rect 67310 14552 67334 14586
rect 67252 14528 67334 14552
rect 68270 14586 68352 14610
rect 68270 14552 68294 14586
rect 68328 14552 68352 14586
rect 68270 14528 68352 14552
rect 69288 14586 69370 14610
rect 69288 14552 69312 14586
rect 69346 14552 69370 14586
rect 69288 14528 69370 14552
rect 70306 14586 70388 14610
rect 70306 14552 70330 14586
rect 70364 14552 70388 14586
rect 70306 14528 70388 14552
rect 71324 14586 71406 14610
rect 71324 14552 71348 14586
rect 71382 14552 71406 14586
rect 71324 14528 71406 14552
rect 72342 14586 72424 14610
rect 72342 14552 72366 14586
rect 72400 14552 72424 14586
rect 72342 14528 72424 14552
rect 73360 14586 73442 14610
rect 73360 14552 73384 14586
rect 73418 14552 73442 14586
rect 73360 14528 73442 14552
rect 74378 14586 74460 14610
rect 74378 14552 74402 14586
rect 74436 14552 74460 14586
rect 74378 14528 74460 14552
rect 54764 14372 54780 14406
rect 55336 14372 55352 14406
rect 55782 14372 55798 14406
rect 56354 14372 56370 14406
rect 56800 14372 56816 14406
rect 57372 14372 57388 14406
rect 57818 14372 57834 14406
rect 58390 14372 58406 14406
rect 58836 14372 58852 14406
rect 59408 14372 59424 14406
rect 59854 14372 59870 14406
rect 60426 14372 60442 14406
rect 60872 14372 60888 14406
rect 61444 14372 61460 14406
rect 61890 14372 61906 14406
rect 62462 14372 62478 14406
rect 62908 14372 62924 14406
rect 63480 14372 63496 14406
rect 63926 14372 63942 14406
rect 64498 14372 64514 14406
rect 64944 14372 64960 14406
rect 65516 14372 65532 14406
rect 65962 14372 65978 14406
rect 66534 14372 66550 14406
rect 66980 14372 66996 14406
rect 67552 14372 67568 14406
rect 67998 14372 68014 14406
rect 68570 14372 68586 14406
rect 69016 14372 69032 14406
rect 69588 14372 69604 14406
rect 70034 14372 70050 14406
rect 70606 14372 70622 14406
rect 71052 14372 71068 14406
rect 71624 14372 71640 14406
rect 72070 14372 72086 14406
rect 72642 14372 72658 14406
rect 73088 14372 73104 14406
rect 73660 14372 73676 14406
rect 74106 14372 74122 14406
rect 74678 14372 74694 14406
rect 36718 13808 36818 13970
rect 38582 13808 38682 13970
rect 36990 13045 37006 13079
rect 37106 13045 37122 13079
rect 37248 13045 37264 13079
rect 37364 13045 37380 13079
rect 37506 13045 37522 13079
rect 37622 13045 37638 13079
rect 37764 13045 37780 13079
rect 37880 13045 37896 13079
rect 38022 13045 38038 13079
rect 38138 13045 38154 13079
rect 38280 13045 38296 13079
rect 38396 13045 38412 13079
rect 36910 12986 36944 13002
rect 36910 12794 36944 12810
rect 37168 12986 37202 13002
rect 37168 12794 37202 12810
rect 37426 12986 37460 13002
rect 37426 12794 37460 12810
rect 37684 12986 37718 13002
rect 37684 12794 37718 12810
rect 37942 12986 37976 13002
rect 37942 12794 37976 12810
rect 38200 12986 38234 13002
rect 38200 12794 38234 12810
rect 38458 12986 38492 13002
rect 38458 12794 38492 12810
rect 36990 12717 37006 12751
rect 37106 12717 37122 12751
rect 37248 12717 37264 12751
rect 37364 12717 37380 12751
rect 37506 12717 37522 12751
rect 37622 12717 37638 12751
rect 37764 12717 37780 12751
rect 37880 12717 37896 12751
rect 38022 12717 38038 12751
rect 38138 12717 38154 12751
rect 38280 12717 38296 12751
rect 38396 12717 38412 12751
rect 36718 12426 36818 12588
rect 38582 12426 38682 12588
rect -872 -102 -838 -96
rect -1188 -136 -1116 -102
rect -916 -136 -838 -102
rect -1372 -852 -1272 -690
rect 35772 -852 35872 -690
rect 54532 14322 54566 14338
rect 42742 13984 42824 14008
rect 42742 13950 42766 13984
rect 42800 13950 42824 13984
rect 42742 13926 42824 13950
rect 43760 13984 43842 14008
rect 43760 13950 43784 13984
rect 43818 13950 43842 13984
rect 42998 13896 43014 13930
rect 43570 13896 43586 13930
rect 43760 13926 43842 13950
rect 44778 13984 44860 14008
rect 44778 13950 44802 13984
rect 44836 13950 44860 13984
rect 44016 13896 44032 13930
rect 44588 13896 44604 13930
rect 44778 13926 44860 13950
rect 45796 13984 45878 14008
rect 45796 13950 45820 13984
rect 45854 13950 45878 13984
rect 45034 13896 45050 13930
rect 45606 13896 45622 13930
rect 45796 13926 45878 13950
rect 46814 13984 46896 14008
rect 46814 13950 46838 13984
rect 46872 13950 46896 13984
rect 46052 13896 46068 13930
rect 46624 13896 46640 13930
rect 46814 13926 46896 13950
rect 47832 13984 47914 14008
rect 47832 13950 47856 13984
rect 47890 13950 47914 13984
rect 47070 13896 47086 13930
rect 47642 13896 47658 13930
rect 47832 13926 47914 13950
rect 48850 13984 48932 14008
rect 48850 13950 48874 13984
rect 48908 13950 48932 13984
rect 48088 13896 48104 13930
rect 48660 13896 48676 13930
rect 48850 13926 48932 13950
rect 49868 13984 49950 14008
rect 49868 13950 49892 13984
rect 49926 13950 49950 13984
rect 49106 13896 49122 13930
rect 49678 13896 49694 13930
rect 49868 13926 49950 13950
rect 50886 13984 50968 14008
rect 50886 13950 50910 13984
rect 50944 13950 50968 13984
rect 50124 13896 50140 13930
rect 50696 13896 50712 13930
rect 50886 13926 50968 13950
rect 51914 13984 51996 14008
rect 51914 13950 51938 13984
rect 51972 13950 51996 13984
rect 51142 13896 51158 13930
rect 51714 13896 51730 13930
rect 51914 13926 51996 13950
rect 42766 13846 42800 13862
rect 42766 13254 42800 13270
rect 43784 13846 43818 13862
rect 43784 13254 43818 13270
rect 44802 13846 44836 13862
rect 44802 13254 44836 13270
rect 45820 13846 45854 13862
rect 45820 13254 45854 13270
rect 46838 13846 46872 13862
rect 46838 13254 46872 13270
rect 47856 13846 47890 13862
rect 47856 13254 47890 13270
rect 48874 13846 48908 13862
rect 48874 13254 48908 13270
rect 49892 13846 49926 13862
rect 49892 13254 49926 13270
rect 50910 13846 50944 13862
rect 50910 13254 50944 13270
rect 51928 13846 51962 13862
rect 54532 13730 54566 13746
rect 55550 14322 55584 14338
rect 55550 13730 55584 13746
rect 56568 14322 56602 14338
rect 56568 13730 56602 13746
rect 57586 14322 57620 14338
rect 57586 13730 57620 13746
rect 58604 14322 58638 14338
rect 58604 13730 58638 13746
rect 59622 14322 59656 14338
rect 59622 13730 59656 13746
rect 60640 14322 60674 14338
rect 60640 13730 60674 13746
rect 61658 14322 61692 14338
rect 61658 13730 61692 13746
rect 62676 14322 62710 14338
rect 62676 13730 62710 13746
rect 63694 14322 63728 14338
rect 63694 13730 63728 13746
rect 64712 14322 64746 14338
rect 64712 13730 64746 13746
rect 65730 14322 65764 14338
rect 65730 13730 65764 13746
rect 66748 14322 66782 14338
rect 66748 13730 66782 13746
rect 67766 14322 67800 14338
rect 67766 13730 67800 13746
rect 68784 14322 68818 14338
rect 68784 13730 68818 13746
rect 69802 14322 69836 14338
rect 69802 13730 69836 13746
rect 70820 14322 70854 14338
rect 70820 13730 70854 13746
rect 71838 14322 71872 14338
rect 71838 13730 71872 13746
rect 72856 14322 72890 14338
rect 72856 13730 72890 13746
rect 73874 14322 73908 14338
rect 73874 13730 73908 13746
rect 74892 14322 74926 14338
rect 74892 13730 74926 13746
rect 54764 13662 54780 13696
rect 55336 13662 55352 13696
rect 55782 13662 55798 13696
rect 56354 13662 56370 13696
rect 56800 13662 56816 13696
rect 57372 13662 57388 13696
rect 57818 13662 57834 13696
rect 58390 13662 58406 13696
rect 58836 13662 58852 13696
rect 59408 13662 59424 13696
rect 59854 13662 59870 13696
rect 60426 13662 60442 13696
rect 60872 13662 60888 13696
rect 61444 13662 61460 13696
rect 61890 13662 61906 13696
rect 62462 13662 62478 13696
rect 62908 13662 62924 13696
rect 63480 13662 63496 13696
rect 63926 13662 63942 13696
rect 64498 13662 64514 13696
rect 64944 13662 64960 13696
rect 65516 13662 65532 13696
rect 65962 13662 65978 13696
rect 66534 13662 66550 13696
rect 66980 13662 66996 13696
rect 67552 13662 67568 13696
rect 67998 13662 68014 13696
rect 68570 13662 68586 13696
rect 69016 13662 69032 13696
rect 69588 13662 69604 13696
rect 70034 13662 70050 13696
rect 70606 13662 70622 13696
rect 71052 13662 71068 13696
rect 71624 13662 71640 13696
rect 72070 13662 72086 13696
rect 72642 13662 72658 13696
rect 73088 13662 73104 13696
rect 73660 13662 73676 13696
rect 74106 13662 74122 13696
rect 74678 13662 74694 13696
rect 54764 13554 54780 13588
rect 55336 13554 55352 13588
rect 55782 13554 55798 13588
rect 56354 13554 56370 13588
rect 56800 13554 56816 13588
rect 57372 13554 57388 13588
rect 57818 13554 57834 13588
rect 58390 13554 58406 13588
rect 58836 13554 58852 13588
rect 59408 13554 59424 13588
rect 59854 13554 59870 13588
rect 60426 13554 60442 13588
rect 60872 13554 60888 13588
rect 61444 13554 61460 13588
rect 61890 13554 61906 13588
rect 62462 13554 62478 13588
rect 62908 13554 62924 13588
rect 63480 13554 63496 13588
rect 63926 13554 63942 13588
rect 64498 13554 64514 13588
rect 64944 13554 64960 13588
rect 65516 13554 65532 13588
rect 65962 13554 65978 13588
rect 66534 13554 66550 13588
rect 66980 13554 66996 13588
rect 67552 13554 67568 13588
rect 67998 13554 68014 13588
rect 68570 13554 68586 13588
rect 69016 13554 69032 13588
rect 69588 13554 69604 13588
rect 70034 13554 70050 13588
rect 70606 13554 70622 13588
rect 71052 13554 71068 13588
rect 71624 13554 71640 13588
rect 72070 13554 72086 13588
rect 72642 13554 72658 13588
rect 73088 13554 73104 13588
rect 73660 13554 73676 13588
rect 74106 13554 74122 13588
rect 74678 13554 74694 13588
rect 51928 13254 51962 13270
rect 54532 13504 54566 13520
rect 42742 13166 42824 13190
rect 42998 13186 43014 13220
rect 43570 13186 43586 13220
rect 42742 13132 42766 13166
rect 42800 13132 42824 13166
rect 42742 13108 42824 13132
rect 43760 13166 43842 13190
rect 44016 13186 44032 13220
rect 44588 13186 44604 13220
rect 43760 13132 43784 13166
rect 43818 13132 43842 13166
rect 42998 13078 43014 13112
rect 43570 13078 43586 13112
rect 43760 13108 43842 13132
rect 44778 13166 44860 13190
rect 45034 13186 45050 13220
rect 45606 13186 45622 13220
rect 44778 13132 44802 13166
rect 44836 13132 44860 13166
rect 44016 13078 44032 13112
rect 44588 13078 44604 13112
rect 44778 13108 44860 13132
rect 45796 13166 45878 13190
rect 46052 13186 46068 13220
rect 46624 13186 46640 13220
rect 45796 13132 45820 13166
rect 45854 13132 45878 13166
rect 45034 13078 45050 13112
rect 45606 13078 45622 13112
rect 45796 13108 45878 13132
rect 46814 13166 46896 13190
rect 47070 13186 47086 13220
rect 47642 13186 47658 13220
rect 46814 13132 46838 13166
rect 46872 13132 46896 13166
rect 46052 13078 46068 13112
rect 46624 13078 46640 13112
rect 46814 13108 46896 13132
rect 47832 13166 47914 13190
rect 48088 13186 48104 13220
rect 48660 13186 48676 13220
rect 47832 13132 47856 13166
rect 47890 13132 47914 13166
rect 47070 13078 47086 13112
rect 47642 13078 47658 13112
rect 47832 13108 47914 13132
rect 48850 13166 48932 13190
rect 49106 13186 49122 13220
rect 49678 13186 49694 13220
rect 48850 13132 48874 13166
rect 48908 13132 48932 13166
rect 48088 13078 48104 13112
rect 48660 13078 48676 13112
rect 48850 13108 48932 13132
rect 49868 13166 49950 13190
rect 50124 13186 50140 13220
rect 50696 13186 50712 13220
rect 49868 13132 49892 13166
rect 49926 13132 49950 13166
rect 49106 13078 49122 13112
rect 49678 13078 49694 13112
rect 49868 13108 49950 13132
rect 50886 13166 50968 13190
rect 51142 13186 51158 13220
rect 51714 13186 51730 13220
rect 50886 13132 50910 13166
rect 50944 13132 50968 13166
rect 50124 13078 50140 13112
rect 50696 13078 50712 13112
rect 50886 13108 50968 13132
rect 51914 13166 51996 13190
rect 51914 13132 51938 13166
rect 51972 13132 51996 13166
rect 51142 13078 51158 13112
rect 51714 13078 51730 13112
rect 51914 13108 51996 13132
rect 48358 13076 48418 13078
rect 42766 13028 42800 13044
rect 42766 12436 42800 12452
rect 43784 13028 43818 13044
rect 43784 12436 43818 12452
rect 44802 13028 44836 13044
rect 44802 12436 44836 12452
rect 45820 13028 45854 13044
rect 45820 12436 45854 12452
rect 46838 13028 46872 13044
rect 46838 12436 46872 12452
rect 47856 13028 47890 13044
rect 47856 12436 47890 12452
rect 48874 13028 48908 13044
rect 48874 12436 48908 12452
rect 49892 13028 49926 13044
rect 49892 12436 49926 12452
rect 50910 13028 50944 13044
rect 50910 12436 50944 12452
rect 51928 13028 51962 13044
rect 54532 12912 54566 12928
rect 55550 13504 55584 13520
rect 55550 12912 55584 12928
rect 56568 13504 56602 13520
rect 56568 12912 56602 12928
rect 57586 13504 57620 13520
rect 57586 12912 57620 12928
rect 58604 13504 58638 13520
rect 58604 12912 58638 12928
rect 59622 13504 59656 13520
rect 59622 12912 59656 12928
rect 60640 13504 60674 13520
rect 60640 12912 60674 12928
rect 61658 13504 61692 13520
rect 61658 12912 61692 12928
rect 62676 13504 62710 13520
rect 62676 12912 62710 12928
rect 63694 13504 63728 13520
rect 63694 12912 63728 12928
rect 64712 13504 64746 13520
rect 64712 12912 64746 12928
rect 65730 13504 65764 13520
rect 65730 12912 65764 12928
rect 66748 13504 66782 13520
rect 66748 12912 66782 12928
rect 67766 13504 67800 13520
rect 67766 12912 67800 12928
rect 68784 13504 68818 13520
rect 68784 12912 68818 12928
rect 69802 13504 69836 13520
rect 69802 12912 69836 12928
rect 70820 13504 70854 13520
rect 70820 12912 70854 12928
rect 71838 13504 71872 13520
rect 71838 12912 71872 12928
rect 72856 13504 72890 13520
rect 72856 12912 72890 12928
rect 73874 13504 73908 13520
rect 73874 12912 73908 12928
rect 74892 13504 74926 13520
rect 74892 12912 74926 12928
rect 54764 12844 54780 12878
rect 55336 12844 55352 12878
rect 55782 12844 55798 12878
rect 56354 12844 56370 12878
rect 56800 12844 56816 12878
rect 57372 12844 57388 12878
rect 57818 12844 57834 12878
rect 58390 12844 58406 12878
rect 58836 12844 58852 12878
rect 59408 12844 59424 12878
rect 59854 12844 59870 12878
rect 60426 12844 60442 12878
rect 60872 12844 60888 12878
rect 61444 12844 61460 12878
rect 61890 12844 61906 12878
rect 62462 12844 62478 12878
rect 62908 12844 62924 12878
rect 63480 12844 63496 12878
rect 63926 12844 63942 12878
rect 64498 12844 64514 12878
rect 64944 12844 64960 12878
rect 65516 12844 65532 12878
rect 65962 12844 65978 12878
rect 66534 12844 66550 12878
rect 66980 12844 66996 12878
rect 67552 12844 67568 12878
rect 67998 12844 68014 12878
rect 68570 12844 68586 12878
rect 69016 12844 69032 12878
rect 69588 12844 69604 12878
rect 70034 12844 70050 12878
rect 70606 12844 70622 12878
rect 71052 12844 71068 12878
rect 71624 12844 71640 12878
rect 72070 12844 72086 12878
rect 72642 12844 72658 12878
rect 73088 12844 73104 12878
rect 73660 12844 73676 12878
rect 74106 12844 74122 12878
rect 74678 12844 74694 12878
rect 55048 12560 55130 12584
rect 55048 12526 55072 12560
rect 55106 12526 55130 12560
rect 55048 12502 55130 12526
rect 56066 12560 56148 12584
rect 56066 12526 56090 12560
rect 56124 12526 56148 12560
rect 56066 12502 56148 12526
rect 57084 12560 57166 12584
rect 57084 12526 57108 12560
rect 57142 12526 57166 12560
rect 57084 12502 57166 12526
rect 58102 12560 58184 12584
rect 58102 12526 58126 12560
rect 58160 12526 58184 12560
rect 58102 12502 58184 12526
rect 59120 12560 59202 12584
rect 59120 12526 59144 12560
rect 59178 12526 59202 12560
rect 59120 12502 59202 12526
rect 60138 12560 60220 12584
rect 60138 12526 60162 12560
rect 60196 12526 60220 12560
rect 60138 12502 60220 12526
rect 61156 12560 61238 12584
rect 61156 12526 61180 12560
rect 61214 12526 61238 12560
rect 61156 12502 61238 12526
rect 62174 12560 62256 12584
rect 62174 12526 62198 12560
rect 62232 12526 62256 12560
rect 62174 12502 62256 12526
rect 63192 12560 63274 12584
rect 63192 12526 63216 12560
rect 63250 12526 63274 12560
rect 63192 12502 63274 12526
rect 64210 12560 64292 12584
rect 64210 12526 64234 12560
rect 64268 12526 64292 12560
rect 64210 12502 64292 12526
rect 65228 12560 65310 12584
rect 65228 12526 65252 12560
rect 65286 12526 65310 12560
rect 65228 12502 65310 12526
rect 66246 12560 66328 12584
rect 66246 12526 66270 12560
rect 66304 12526 66328 12560
rect 66246 12502 66328 12526
rect 67264 12560 67346 12584
rect 67264 12526 67288 12560
rect 67322 12526 67346 12560
rect 67264 12502 67346 12526
rect 68282 12560 68364 12584
rect 68282 12526 68306 12560
rect 68340 12526 68364 12560
rect 68282 12502 68364 12526
rect 69300 12560 69382 12584
rect 69300 12526 69324 12560
rect 69358 12526 69382 12560
rect 69300 12502 69382 12526
rect 70318 12560 70400 12584
rect 70318 12526 70342 12560
rect 70376 12526 70400 12560
rect 70318 12502 70400 12526
rect 71336 12560 71418 12584
rect 71336 12526 71360 12560
rect 71394 12526 71418 12560
rect 71336 12502 71418 12526
rect 72354 12560 72436 12584
rect 72354 12526 72378 12560
rect 72412 12526 72436 12560
rect 72354 12502 72436 12526
rect 73372 12560 73454 12584
rect 73372 12526 73396 12560
rect 73430 12526 73454 12560
rect 73372 12502 73454 12526
rect 74390 12560 74472 12584
rect 74390 12526 74414 12560
rect 74448 12526 74472 12560
rect 74390 12502 74472 12526
rect 51928 12436 51962 12452
rect 44290 12402 44350 12404
rect 45304 12402 45364 12404
rect 49378 12402 49438 12404
rect 50394 12402 50454 12404
rect 42742 12348 42824 12372
rect 42998 12368 43014 12402
rect 43570 12368 43586 12402
rect 42742 12314 42766 12348
rect 42800 12314 42824 12348
rect 42742 12290 42824 12314
rect 43760 12348 43842 12372
rect 44016 12368 44032 12402
rect 44588 12368 44604 12402
rect 43760 12314 43784 12348
rect 43818 12314 43842 12348
rect 42998 12260 43014 12294
rect 43570 12260 43586 12294
rect 43760 12290 43842 12314
rect 44778 12348 44860 12372
rect 45034 12368 45050 12402
rect 45606 12368 45622 12402
rect 44778 12314 44802 12348
rect 44836 12314 44860 12348
rect 44016 12260 44032 12294
rect 44588 12260 44604 12294
rect 44778 12290 44860 12314
rect 45796 12348 45878 12372
rect 46052 12368 46068 12402
rect 46624 12368 46640 12402
rect 45796 12314 45820 12348
rect 45854 12314 45878 12348
rect 45034 12260 45050 12294
rect 45606 12260 45622 12294
rect 45796 12290 45878 12314
rect 46814 12348 46896 12372
rect 47070 12368 47086 12402
rect 47642 12368 47658 12402
rect 46814 12314 46838 12348
rect 46872 12314 46896 12348
rect 46052 12260 46068 12294
rect 46624 12260 46640 12294
rect 46814 12290 46896 12314
rect 47832 12348 47914 12372
rect 48088 12368 48104 12402
rect 48660 12368 48676 12402
rect 47832 12314 47856 12348
rect 47890 12314 47914 12348
rect 47070 12260 47086 12294
rect 47642 12260 47658 12294
rect 47832 12290 47914 12314
rect 48850 12348 48932 12372
rect 49106 12368 49122 12402
rect 49678 12368 49694 12402
rect 48850 12314 48874 12348
rect 48908 12314 48932 12348
rect 48088 12260 48104 12294
rect 48660 12260 48676 12294
rect 48850 12290 48932 12314
rect 49868 12348 49950 12372
rect 50124 12368 50140 12402
rect 50696 12368 50712 12402
rect 49868 12314 49892 12348
rect 49926 12314 49950 12348
rect 49106 12260 49122 12294
rect 49678 12260 49694 12294
rect 49868 12290 49950 12314
rect 50886 12348 50968 12372
rect 51142 12368 51158 12402
rect 51714 12368 51730 12402
rect 50886 12314 50910 12348
rect 50944 12314 50968 12348
rect 50124 12260 50140 12294
rect 50696 12260 50712 12294
rect 50886 12290 50968 12314
rect 51914 12348 51996 12372
rect 51914 12314 51938 12348
rect 51972 12314 51996 12348
rect 51142 12260 51158 12294
rect 51714 12260 51730 12294
rect 51914 12290 51996 12314
rect 42766 12210 42800 12226
rect 42766 11618 42800 11634
rect 43784 12210 43818 12226
rect 43784 11618 43818 11634
rect 44802 12210 44836 12226
rect 44802 11618 44836 11634
rect 45820 12210 45854 12226
rect 45820 11618 45854 11634
rect 46838 12210 46872 12226
rect 46838 11618 46872 11634
rect 47856 12210 47890 12226
rect 47856 11618 47890 11634
rect 48874 12210 48908 12226
rect 48874 11618 48908 11634
rect 49892 12210 49926 12226
rect 49892 11618 49926 11634
rect 50910 12210 50944 12226
rect 50910 11618 50944 11634
rect 51928 12210 51962 12226
rect 54764 12176 54780 12210
rect 55336 12176 55352 12210
rect 55782 12176 55798 12210
rect 56354 12176 56370 12210
rect 56800 12176 56816 12210
rect 57372 12176 57388 12210
rect 57818 12176 57834 12210
rect 58390 12176 58406 12210
rect 58836 12176 58852 12210
rect 59408 12176 59424 12210
rect 59854 12176 59870 12210
rect 60426 12176 60442 12210
rect 60872 12176 60888 12210
rect 61444 12176 61460 12210
rect 61890 12176 61906 12210
rect 62462 12176 62478 12210
rect 62908 12176 62924 12210
rect 63480 12176 63496 12210
rect 63926 12176 63942 12210
rect 64498 12176 64514 12210
rect 64944 12176 64960 12210
rect 65516 12176 65532 12210
rect 65962 12176 65978 12210
rect 66534 12176 66550 12210
rect 66980 12176 66996 12210
rect 67552 12176 67568 12210
rect 67998 12176 68014 12210
rect 68570 12176 68586 12210
rect 69016 12176 69032 12210
rect 69588 12176 69604 12210
rect 70034 12176 70050 12210
rect 70606 12176 70622 12210
rect 71052 12176 71068 12210
rect 71624 12176 71640 12210
rect 72070 12176 72086 12210
rect 72642 12176 72658 12210
rect 73088 12176 73104 12210
rect 73660 12176 73676 12210
rect 74106 12176 74122 12210
rect 74678 12176 74694 12210
rect 64188 12170 64248 12176
rect 51928 11618 51962 11634
rect 54532 12126 54566 12142
rect 44294 11584 44354 11586
rect 45308 11584 45368 11586
rect 49382 11584 49442 11586
rect 50398 11584 50458 11586
rect 42742 11530 42824 11554
rect 42998 11550 43014 11584
rect 43570 11550 43586 11584
rect 42742 11496 42766 11530
rect 42800 11496 42824 11530
rect 42742 11472 42824 11496
rect 43760 11530 43842 11554
rect 44016 11550 44032 11584
rect 44588 11550 44604 11584
rect 43760 11496 43784 11530
rect 43818 11496 43842 11530
rect 42998 11442 43014 11476
rect 43570 11442 43586 11476
rect 43760 11472 43842 11496
rect 44778 11530 44860 11554
rect 45034 11550 45050 11584
rect 45606 11550 45622 11584
rect 44778 11496 44802 11530
rect 44836 11496 44860 11530
rect 44016 11442 44032 11476
rect 44588 11442 44604 11476
rect 44778 11472 44860 11496
rect 45796 11530 45878 11554
rect 46052 11550 46068 11584
rect 46624 11550 46640 11584
rect 45796 11496 45820 11530
rect 45854 11496 45878 11530
rect 45034 11442 45050 11476
rect 45606 11442 45622 11476
rect 45796 11472 45878 11496
rect 46814 11530 46896 11554
rect 47070 11550 47086 11584
rect 47642 11550 47658 11584
rect 46814 11496 46838 11530
rect 46872 11496 46896 11530
rect 46052 11442 46068 11476
rect 46624 11442 46640 11476
rect 46814 11472 46896 11496
rect 47832 11530 47914 11554
rect 48088 11550 48104 11584
rect 48660 11550 48676 11584
rect 47832 11496 47856 11530
rect 47890 11496 47914 11530
rect 47070 11442 47086 11476
rect 47642 11442 47658 11476
rect 47832 11472 47914 11496
rect 48850 11530 48932 11554
rect 49106 11550 49122 11584
rect 49678 11550 49694 11584
rect 48850 11496 48874 11530
rect 48908 11496 48932 11530
rect 48088 11442 48104 11476
rect 48660 11442 48676 11476
rect 48850 11472 48932 11496
rect 49868 11530 49950 11554
rect 50124 11550 50140 11584
rect 50696 11550 50712 11584
rect 49868 11496 49892 11530
rect 49926 11496 49950 11530
rect 49106 11442 49122 11476
rect 49678 11442 49694 11476
rect 49868 11472 49950 11496
rect 50886 11530 50968 11554
rect 51142 11550 51158 11584
rect 51714 11550 51730 11584
rect 50886 11496 50910 11530
rect 50944 11496 50968 11530
rect 50124 11442 50140 11476
rect 50696 11442 50712 11476
rect 50886 11472 50968 11496
rect 51914 11530 51996 11554
rect 54532 11534 54566 11550
rect 55550 12126 55584 12142
rect 55550 11534 55584 11550
rect 56568 12126 56602 12142
rect 56568 11534 56602 11550
rect 57586 12126 57620 12142
rect 57586 11534 57620 11550
rect 58604 12126 58638 12142
rect 58604 11534 58638 11550
rect 59622 12126 59656 12142
rect 59622 11534 59656 11550
rect 60640 12126 60674 12142
rect 60640 11534 60674 11550
rect 61658 12126 61692 12142
rect 61658 11534 61692 11550
rect 62676 12126 62710 12142
rect 62676 11534 62710 11550
rect 63694 12126 63728 12142
rect 63694 11534 63728 11550
rect 64712 12126 64746 12142
rect 64712 11534 64746 11550
rect 65730 12126 65764 12142
rect 65730 11534 65764 11550
rect 66748 12126 66782 12142
rect 66748 11534 66782 11550
rect 67766 12126 67800 12142
rect 67766 11534 67800 11550
rect 68784 12126 68818 12142
rect 68784 11534 68818 11550
rect 69802 12126 69836 12142
rect 69802 11534 69836 11550
rect 70820 12126 70854 12142
rect 70820 11534 70854 11550
rect 71838 12126 71872 12142
rect 71838 11534 71872 11550
rect 72856 12126 72890 12142
rect 72856 11534 72890 11550
rect 73874 12126 73908 12142
rect 73874 11534 73908 11550
rect 74892 12126 74926 12142
rect 74892 11534 74926 11550
rect 51914 11496 51938 11530
rect 51972 11496 51996 11530
rect 60116 11500 60176 11506
rect 62152 11500 62212 11506
rect 63172 11500 63232 11506
rect 68244 11500 68304 11506
rect 51142 11442 51158 11476
rect 51714 11442 51730 11476
rect 51914 11472 51996 11496
rect 54764 11466 54780 11500
rect 55336 11466 55352 11500
rect 55782 11466 55798 11500
rect 56354 11466 56370 11500
rect 56800 11466 56816 11500
rect 57372 11466 57388 11500
rect 57818 11466 57834 11500
rect 58390 11466 58406 11500
rect 58836 11466 58852 11500
rect 59408 11466 59424 11500
rect 59854 11466 59870 11500
rect 60426 11466 60442 11500
rect 60872 11466 60888 11500
rect 61444 11466 61460 11500
rect 61890 11466 61906 11500
rect 62462 11466 62478 11500
rect 62908 11466 62924 11500
rect 63480 11466 63496 11500
rect 63926 11466 63942 11500
rect 64498 11466 64514 11500
rect 64944 11466 64960 11500
rect 65516 11466 65532 11500
rect 65962 11466 65978 11500
rect 66534 11466 66550 11500
rect 66980 11466 66996 11500
rect 67552 11466 67568 11500
rect 67998 11466 68014 11500
rect 68570 11466 68586 11500
rect 69016 11466 69032 11500
rect 69588 11466 69604 11500
rect 70034 11466 70050 11500
rect 70606 11466 70622 11500
rect 71052 11466 71068 11500
rect 71624 11466 71640 11500
rect 72070 11466 72086 11500
rect 72642 11466 72658 11500
rect 73088 11466 73104 11500
rect 73660 11466 73676 11500
rect 74106 11466 74122 11500
rect 74678 11466 74694 11500
rect 42766 11392 42800 11408
rect 42766 10800 42800 10816
rect 43784 11392 43818 11408
rect 43784 10800 43818 10816
rect 44802 11392 44836 11408
rect 44802 10800 44836 10816
rect 45820 11392 45854 11408
rect 45820 10800 45854 10816
rect 46838 11392 46872 11408
rect 46838 10800 46872 10816
rect 47856 11392 47890 11408
rect 47856 10800 47890 10816
rect 48874 11392 48908 11408
rect 48874 10800 48908 10816
rect 49892 11392 49926 11408
rect 49892 10800 49926 10816
rect 50910 11392 50944 11408
rect 50910 10800 50944 10816
rect 51928 11392 51962 11408
rect 55036 11254 55118 11278
rect 55036 11220 55060 11254
rect 55094 11220 55118 11254
rect 55036 11196 55118 11220
rect 56054 11254 56136 11278
rect 56054 11220 56078 11254
rect 56112 11220 56136 11254
rect 56054 11196 56136 11220
rect 57072 11254 57154 11278
rect 57072 11220 57096 11254
rect 57130 11220 57154 11254
rect 57072 11196 57154 11220
rect 58090 11254 58172 11278
rect 58090 11220 58114 11254
rect 58148 11220 58172 11254
rect 58090 11196 58172 11220
rect 59108 11254 59190 11278
rect 59108 11220 59132 11254
rect 59166 11220 59190 11254
rect 59108 11196 59190 11220
rect 60126 11254 60208 11278
rect 60126 11220 60150 11254
rect 60184 11220 60208 11254
rect 60126 11196 60208 11220
rect 61144 11254 61226 11278
rect 61144 11220 61168 11254
rect 61202 11220 61226 11254
rect 61144 11196 61226 11220
rect 62162 11254 62244 11278
rect 62162 11220 62186 11254
rect 62220 11220 62244 11254
rect 62162 11196 62244 11220
rect 63180 11254 63262 11278
rect 63180 11220 63204 11254
rect 63238 11220 63262 11254
rect 63180 11196 63262 11220
rect 64198 11254 64280 11278
rect 64198 11220 64222 11254
rect 64256 11220 64280 11254
rect 64198 11196 64280 11220
rect 65216 11254 65298 11278
rect 65216 11220 65240 11254
rect 65274 11220 65298 11254
rect 65216 11196 65298 11220
rect 66234 11254 66316 11278
rect 66234 11220 66258 11254
rect 66292 11220 66316 11254
rect 66234 11196 66316 11220
rect 67252 11254 67334 11278
rect 67252 11220 67276 11254
rect 67310 11220 67334 11254
rect 67252 11196 67334 11220
rect 68270 11254 68352 11278
rect 68270 11220 68294 11254
rect 68328 11220 68352 11254
rect 68270 11196 68352 11220
rect 69288 11254 69370 11278
rect 69288 11220 69312 11254
rect 69346 11220 69370 11254
rect 69288 11196 69370 11220
rect 70306 11254 70388 11278
rect 70306 11220 70330 11254
rect 70364 11220 70388 11254
rect 70306 11196 70388 11220
rect 71324 11254 71406 11278
rect 71324 11220 71348 11254
rect 71382 11220 71406 11254
rect 71324 11196 71406 11220
rect 72342 11254 72424 11278
rect 72342 11220 72366 11254
rect 72400 11220 72424 11254
rect 72342 11196 72424 11220
rect 73360 11254 73442 11278
rect 73360 11220 73384 11254
rect 73418 11220 73442 11254
rect 73360 11196 73442 11220
rect 74378 11254 74460 11278
rect 74378 11220 74402 11254
rect 74436 11220 74460 11254
rect 74378 11196 74460 11220
rect 54764 10944 54780 10978
rect 55336 10944 55352 10978
rect 55782 10944 55798 10978
rect 56354 10944 56370 10978
rect 56800 10944 56816 10978
rect 57372 10944 57388 10978
rect 57818 10944 57834 10978
rect 58390 10944 58406 10978
rect 58836 10944 58852 10978
rect 59408 10944 59424 10978
rect 59854 10944 59870 10978
rect 60426 10944 60442 10978
rect 60872 10944 60888 10978
rect 61444 10944 61460 10978
rect 61890 10944 61906 10978
rect 62462 10944 62478 10978
rect 62908 10944 62924 10978
rect 63480 10944 63496 10978
rect 63926 10944 63942 10978
rect 64498 10944 64514 10978
rect 64944 10944 64960 10978
rect 65516 10944 65532 10978
rect 65962 10944 65978 10978
rect 66534 10944 66550 10978
rect 66980 10944 66996 10978
rect 67552 10944 67568 10978
rect 67998 10944 68014 10978
rect 68570 10944 68586 10978
rect 69016 10944 69032 10978
rect 69588 10944 69604 10978
rect 70034 10944 70050 10978
rect 70606 10944 70622 10978
rect 71052 10944 71068 10978
rect 71624 10944 71640 10978
rect 72070 10944 72086 10978
rect 72642 10944 72658 10978
rect 73088 10944 73104 10978
rect 73660 10944 73676 10978
rect 74106 10944 74122 10978
rect 74678 10944 74694 10978
rect 56050 10940 56110 10944
rect 57066 10940 57126 10944
rect 61142 10936 61202 10944
rect 65208 10940 65268 10944
rect 67242 10940 67302 10944
rect 73354 10940 73414 10944
rect 51928 10800 51962 10816
rect 54532 10894 54566 10910
rect 42742 10712 42824 10736
rect 42998 10732 43014 10766
rect 43570 10732 43586 10766
rect 42742 10678 42766 10712
rect 42800 10678 42824 10712
rect 42742 10654 42824 10678
rect 43760 10712 43842 10736
rect 44016 10732 44032 10766
rect 44588 10732 44604 10766
rect 43760 10678 43784 10712
rect 43818 10678 43842 10712
rect 42998 10624 43014 10658
rect 43570 10624 43586 10658
rect 43760 10654 43842 10678
rect 44778 10712 44860 10736
rect 45034 10732 45050 10766
rect 45606 10732 45622 10766
rect 44778 10678 44802 10712
rect 44836 10678 44860 10712
rect 44016 10624 44032 10658
rect 44588 10624 44604 10658
rect 44778 10654 44860 10678
rect 45796 10712 45878 10736
rect 46052 10732 46068 10766
rect 46624 10732 46640 10766
rect 45796 10678 45820 10712
rect 45854 10678 45878 10712
rect 45034 10624 45050 10658
rect 45606 10624 45622 10658
rect 45796 10654 45878 10678
rect 46814 10712 46896 10736
rect 47070 10732 47086 10766
rect 47642 10732 47658 10766
rect 46814 10678 46838 10712
rect 46872 10678 46896 10712
rect 46052 10624 46068 10658
rect 46624 10624 46640 10658
rect 46814 10654 46896 10678
rect 47832 10712 47914 10736
rect 48088 10732 48104 10766
rect 48660 10732 48676 10766
rect 47832 10678 47856 10712
rect 47890 10678 47914 10712
rect 47070 10624 47086 10658
rect 47642 10624 47658 10658
rect 47832 10654 47914 10678
rect 48850 10712 48932 10736
rect 49106 10732 49122 10766
rect 49678 10732 49694 10766
rect 48850 10678 48874 10712
rect 48908 10678 48932 10712
rect 48088 10624 48104 10658
rect 48660 10624 48676 10658
rect 48850 10654 48932 10678
rect 49868 10712 49950 10736
rect 50124 10732 50140 10766
rect 50696 10732 50712 10766
rect 49868 10678 49892 10712
rect 49926 10678 49950 10712
rect 49106 10624 49122 10658
rect 49678 10624 49694 10658
rect 49868 10654 49950 10678
rect 50886 10712 50968 10736
rect 51142 10732 51158 10766
rect 51714 10732 51730 10766
rect 50886 10678 50910 10712
rect 50944 10678 50968 10712
rect 50124 10624 50140 10658
rect 50696 10624 50712 10658
rect 50886 10654 50968 10678
rect 51914 10712 51996 10736
rect 51914 10678 51938 10712
rect 51972 10678 51996 10712
rect 51142 10624 51158 10658
rect 51714 10624 51730 10658
rect 51914 10654 51996 10678
rect 48354 10622 48414 10624
rect 42766 10574 42800 10590
rect 42766 9982 42800 9998
rect 43784 10574 43818 10590
rect 43784 9982 43818 9998
rect 44802 10574 44836 10590
rect 44802 9982 44836 9998
rect 45820 10574 45854 10590
rect 45820 9982 45854 9998
rect 46838 10574 46872 10590
rect 46838 9982 46872 9998
rect 47856 10574 47890 10590
rect 47856 9982 47890 9998
rect 48874 10574 48908 10590
rect 48874 9982 48908 9998
rect 49892 10574 49926 10590
rect 49892 9982 49926 9998
rect 50910 10574 50944 10590
rect 50910 9982 50944 9998
rect 51928 10574 51962 10590
rect 54532 10302 54566 10318
rect 55550 10894 55584 10910
rect 55550 10302 55584 10318
rect 56568 10894 56602 10910
rect 56568 10302 56602 10318
rect 57586 10894 57620 10910
rect 57586 10302 57620 10318
rect 58604 10894 58638 10910
rect 58604 10302 58638 10318
rect 59622 10894 59656 10910
rect 59622 10302 59656 10318
rect 60640 10894 60674 10910
rect 60640 10302 60674 10318
rect 61658 10894 61692 10910
rect 61658 10302 61692 10318
rect 62676 10894 62710 10910
rect 62676 10302 62710 10318
rect 63694 10894 63728 10910
rect 63694 10302 63728 10318
rect 64712 10894 64746 10910
rect 64712 10302 64746 10318
rect 65730 10894 65764 10910
rect 65730 10302 65764 10318
rect 66748 10894 66782 10910
rect 66748 10302 66782 10318
rect 67766 10894 67800 10910
rect 67766 10302 67800 10318
rect 68784 10894 68818 10910
rect 68784 10302 68818 10318
rect 69802 10894 69836 10910
rect 69802 10302 69836 10318
rect 70820 10894 70854 10910
rect 70820 10302 70854 10318
rect 71838 10894 71872 10910
rect 71838 10302 71872 10318
rect 72856 10894 72890 10910
rect 72856 10302 72890 10318
rect 73874 10894 73908 10910
rect 73874 10302 73908 10318
rect 74892 10894 74926 10910
rect 74926 10318 74932 10366
rect 74892 10302 74926 10318
rect 58076 10268 58136 10270
rect 54764 10234 54780 10268
rect 55336 10234 55352 10268
rect 55782 10234 55798 10268
rect 56354 10234 56370 10268
rect 56800 10234 56816 10268
rect 57372 10234 57388 10268
rect 57818 10234 57834 10268
rect 58390 10234 58406 10268
rect 58836 10234 58852 10268
rect 59408 10234 59424 10268
rect 59854 10234 59870 10268
rect 60426 10234 60442 10268
rect 60872 10234 60888 10268
rect 61444 10234 61460 10268
rect 61890 10234 61906 10268
rect 62462 10234 62478 10268
rect 62908 10234 62924 10268
rect 63480 10234 63496 10268
rect 63926 10234 63942 10268
rect 64498 10234 64514 10268
rect 64944 10234 64960 10268
rect 65516 10234 65532 10268
rect 65962 10234 65978 10268
rect 66534 10234 66550 10268
rect 66980 10234 66996 10268
rect 67552 10234 67568 10268
rect 67998 10234 68014 10268
rect 68570 10234 68586 10268
rect 69016 10234 69032 10268
rect 69588 10234 69604 10268
rect 70034 10234 70050 10268
rect 70606 10234 70622 10268
rect 71052 10234 71068 10268
rect 71624 10234 71640 10268
rect 72070 10234 72086 10268
rect 72642 10234 72658 10268
rect 73088 10234 73104 10268
rect 73660 10234 73676 10268
rect 74106 10234 74122 10268
rect 74678 10234 74694 10268
rect 60110 10230 60170 10234
rect 69268 10220 69328 10234
rect 70302 10220 70362 10234
rect 51928 9982 51962 9998
rect 55024 10018 55106 10042
rect 55024 9984 55048 10018
rect 55082 9984 55106 10018
rect 55024 9960 55106 9984
rect 56042 10018 56124 10042
rect 56042 9984 56066 10018
rect 56100 9984 56124 10018
rect 56042 9960 56124 9984
rect 57060 10018 57142 10042
rect 57060 9984 57084 10018
rect 57118 9984 57142 10018
rect 57060 9960 57142 9984
rect 58078 10018 58160 10042
rect 58078 9984 58102 10018
rect 58136 9984 58160 10018
rect 58078 9960 58160 9984
rect 59096 10018 59178 10042
rect 59096 9984 59120 10018
rect 59154 9984 59178 10018
rect 59096 9960 59178 9984
rect 60114 10018 60196 10042
rect 60114 9984 60138 10018
rect 60172 9984 60196 10018
rect 60114 9960 60196 9984
rect 61132 10018 61214 10042
rect 61132 9984 61156 10018
rect 61190 9984 61214 10018
rect 61132 9960 61214 9984
rect 62150 10018 62232 10042
rect 62150 9984 62174 10018
rect 62208 9984 62232 10018
rect 62150 9960 62232 9984
rect 63168 10018 63250 10042
rect 63168 9984 63192 10018
rect 63226 9984 63250 10018
rect 63168 9960 63250 9984
rect 64186 10018 64268 10042
rect 64186 9984 64210 10018
rect 64244 9984 64268 10018
rect 64186 9960 64268 9984
rect 65204 10018 65286 10042
rect 65204 9984 65228 10018
rect 65262 9984 65286 10018
rect 65204 9960 65286 9984
rect 66222 10018 66304 10042
rect 66222 9984 66246 10018
rect 66280 9984 66304 10018
rect 66222 9960 66304 9984
rect 67240 10018 67322 10042
rect 67240 9984 67264 10018
rect 67298 9984 67322 10018
rect 67240 9960 67322 9984
rect 68258 10018 68340 10042
rect 68258 9984 68282 10018
rect 68316 9984 68340 10018
rect 68258 9960 68340 9984
rect 69276 10018 69358 10042
rect 69276 9984 69300 10018
rect 69334 9984 69358 10018
rect 69276 9960 69358 9984
rect 70294 10018 70376 10042
rect 70294 9984 70318 10018
rect 70352 9984 70376 10018
rect 70294 9960 70376 9984
rect 71312 10018 71394 10042
rect 71312 9984 71336 10018
rect 71370 9984 71394 10018
rect 71312 9960 71394 9984
rect 72330 10018 72412 10042
rect 72330 9984 72354 10018
rect 72388 9984 72412 10018
rect 72330 9960 72412 9984
rect 73348 10018 73430 10042
rect 73348 9984 73372 10018
rect 73406 9984 73430 10018
rect 73348 9960 73430 9984
rect 74366 10018 74448 10042
rect 74366 9984 74390 10018
rect 74424 9984 74448 10018
rect 74366 9960 74448 9984
rect 44280 9948 44340 9950
rect 45294 9948 45354 9950
rect 49368 9948 49428 9950
rect 50384 9948 50444 9950
rect 42742 9894 42824 9918
rect 42998 9914 43014 9948
rect 43570 9914 43586 9948
rect 42742 9860 42766 9894
rect 42800 9860 42824 9894
rect 42742 9836 42824 9860
rect 43760 9894 43842 9918
rect 44016 9914 44032 9948
rect 44588 9914 44604 9948
rect 43760 9860 43784 9894
rect 43818 9860 43842 9894
rect 42998 9806 43014 9840
rect 43570 9806 43586 9840
rect 43760 9836 43842 9860
rect 44778 9894 44860 9918
rect 45034 9914 45050 9948
rect 45606 9914 45622 9948
rect 44778 9860 44802 9894
rect 44836 9860 44860 9894
rect 44016 9806 44032 9840
rect 44588 9806 44604 9840
rect 44778 9836 44860 9860
rect 45796 9894 45878 9918
rect 46052 9914 46068 9948
rect 46624 9914 46640 9948
rect 45796 9860 45820 9894
rect 45854 9860 45878 9894
rect 45034 9806 45050 9840
rect 45606 9806 45622 9840
rect 45796 9836 45878 9860
rect 46814 9894 46896 9918
rect 47070 9914 47086 9948
rect 47642 9914 47658 9948
rect 46814 9860 46838 9894
rect 46872 9860 46896 9894
rect 46052 9806 46068 9840
rect 46624 9806 46640 9840
rect 46814 9836 46896 9860
rect 47832 9894 47914 9918
rect 48088 9914 48104 9948
rect 48660 9914 48676 9948
rect 47832 9860 47856 9894
rect 47890 9860 47914 9894
rect 47070 9806 47086 9840
rect 47642 9806 47658 9840
rect 47832 9836 47914 9860
rect 48850 9894 48932 9918
rect 49106 9914 49122 9948
rect 49678 9914 49694 9948
rect 48850 9860 48874 9894
rect 48908 9860 48932 9894
rect 48088 9806 48104 9840
rect 48660 9806 48676 9840
rect 48850 9836 48932 9860
rect 49868 9894 49950 9918
rect 50124 9914 50140 9948
rect 50696 9914 50712 9948
rect 49868 9860 49892 9894
rect 49926 9860 49950 9894
rect 49106 9806 49122 9840
rect 49678 9806 49694 9840
rect 49868 9836 49950 9860
rect 50886 9894 50968 9918
rect 51142 9914 51158 9948
rect 51714 9914 51730 9948
rect 50886 9860 50910 9894
rect 50944 9860 50968 9894
rect 50124 9806 50140 9840
rect 50696 9806 50712 9840
rect 50886 9836 50968 9860
rect 51914 9894 51996 9918
rect 51914 9860 51938 9894
rect 51972 9860 51996 9894
rect 51142 9806 51158 9840
rect 51714 9806 51730 9840
rect 51914 9836 51996 9860
rect 42766 9756 42800 9772
rect 42766 9164 42800 9180
rect 43784 9756 43818 9772
rect 43784 9164 43818 9180
rect 44802 9756 44836 9772
rect 44802 9164 44836 9180
rect 45820 9756 45854 9772
rect 45820 9164 45854 9180
rect 46838 9756 46872 9772
rect 46838 9164 46872 9180
rect 47856 9756 47890 9772
rect 47856 9164 47890 9180
rect 48874 9756 48908 9772
rect 48874 9164 48908 9180
rect 49892 9756 49926 9772
rect 49892 9164 49926 9180
rect 50910 9756 50944 9772
rect 50910 9164 50944 9180
rect 51928 9756 51962 9772
rect 54762 9710 54778 9744
rect 55334 9710 55350 9744
rect 55780 9710 55796 9744
rect 56352 9710 56368 9744
rect 56798 9710 56814 9744
rect 57370 9710 57386 9744
rect 57816 9710 57832 9744
rect 58388 9710 58404 9744
rect 58834 9710 58850 9744
rect 59406 9710 59422 9744
rect 59852 9710 59868 9744
rect 60424 9710 60440 9744
rect 60870 9710 60886 9744
rect 61442 9710 61458 9744
rect 61888 9710 61904 9744
rect 62460 9710 62476 9744
rect 62906 9710 62922 9744
rect 63478 9710 63494 9744
rect 63924 9710 63940 9744
rect 64496 9710 64512 9744
rect 64942 9710 64958 9744
rect 65514 9710 65530 9744
rect 65960 9710 65976 9744
rect 66532 9710 66548 9744
rect 66978 9710 66994 9744
rect 67550 9710 67566 9744
rect 67996 9710 68012 9744
rect 68568 9710 68584 9744
rect 69014 9710 69030 9744
rect 69586 9710 69602 9744
rect 70032 9710 70048 9744
rect 70604 9710 70620 9744
rect 71050 9710 71066 9744
rect 71622 9710 71638 9744
rect 72068 9710 72084 9744
rect 72640 9710 72656 9744
rect 73086 9710 73102 9744
rect 73658 9710 73674 9744
rect 74104 9710 74120 9744
rect 74676 9710 74692 9744
rect 57072 9706 57132 9710
rect 51928 9164 51962 9180
rect 54530 9660 54564 9676
rect 44284 9130 44344 9132
rect 45298 9130 45358 9132
rect 49372 9130 49432 9132
rect 50388 9130 50448 9132
rect 42742 9076 42824 9100
rect 42998 9096 43014 9130
rect 43570 9096 43586 9130
rect 42742 9042 42766 9076
rect 42800 9042 42824 9076
rect 42742 9018 42824 9042
rect 43760 9076 43842 9100
rect 44016 9096 44032 9130
rect 44588 9096 44604 9130
rect 43760 9042 43784 9076
rect 43818 9042 43842 9076
rect 42998 8988 43014 9022
rect 43570 8988 43586 9022
rect 43760 9018 43842 9042
rect 44778 9076 44860 9100
rect 45034 9096 45050 9130
rect 45606 9096 45622 9130
rect 44778 9042 44802 9076
rect 44836 9042 44860 9076
rect 44016 8988 44032 9022
rect 44588 8988 44604 9022
rect 44778 9018 44860 9042
rect 45796 9076 45878 9100
rect 46052 9096 46068 9130
rect 46624 9096 46640 9130
rect 45796 9042 45820 9076
rect 45854 9042 45878 9076
rect 45034 8988 45050 9022
rect 45606 8988 45622 9022
rect 45796 9018 45878 9042
rect 46814 9076 46896 9100
rect 47070 9096 47086 9130
rect 47642 9096 47658 9130
rect 46814 9042 46838 9076
rect 46872 9042 46896 9076
rect 46052 8988 46068 9022
rect 46624 8988 46640 9022
rect 46814 9018 46896 9042
rect 47832 9076 47914 9100
rect 48088 9096 48104 9130
rect 48660 9096 48676 9130
rect 47832 9042 47856 9076
rect 47890 9042 47914 9076
rect 47070 8988 47086 9022
rect 47642 8988 47658 9022
rect 47832 9018 47914 9042
rect 48850 9076 48932 9100
rect 49106 9096 49122 9130
rect 49678 9096 49694 9130
rect 48850 9042 48874 9076
rect 48908 9042 48932 9076
rect 48088 8988 48104 9022
rect 48660 8988 48676 9022
rect 48850 9018 48932 9042
rect 49868 9076 49950 9100
rect 50124 9096 50140 9130
rect 50696 9096 50712 9130
rect 49868 9042 49892 9076
rect 49926 9042 49950 9076
rect 49106 8988 49122 9022
rect 49678 8988 49694 9022
rect 49868 9018 49950 9042
rect 50886 9076 50968 9100
rect 51142 9096 51158 9130
rect 51714 9096 51730 9130
rect 50886 9042 50910 9076
rect 50944 9042 50968 9076
rect 50124 8988 50140 9022
rect 50696 8988 50712 9022
rect 50886 9018 50968 9042
rect 51914 9076 51996 9100
rect 51914 9042 51938 9076
rect 51972 9042 51996 9076
rect 54530 9068 54564 9084
rect 55548 9660 55582 9676
rect 55548 9068 55582 9084
rect 56566 9660 56600 9676
rect 56566 9068 56600 9084
rect 57584 9660 57618 9676
rect 57584 9068 57618 9084
rect 58602 9660 58636 9676
rect 58602 9068 58636 9084
rect 59620 9660 59654 9676
rect 59620 9068 59654 9084
rect 60638 9660 60672 9676
rect 60638 9068 60672 9084
rect 61656 9660 61690 9676
rect 61656 9068 61690 9084
rect 62674 9660 62708 9676
rect 62674 9068 62708 9084
rect 63692 9660 63726 9676
rect 63692 9068 63726 9084
rect 64710 9660 64744 9676
rect 64710 9068 64744 9084
rect 65728 9660 65762 9676
rect 65728 9068 65762 9084
rect 66746 9660 66780 9676
rect 66746 9068 66780 9084
rect 67764 9660 67798 9676
rect 67764 9068 67798 9084
rect 68782 9660 68816 9676
rect 68782 9068 68816 9084
rect 69800 9660 69834 9676
rect 69800 9068 69834 9084
rect 70818 9660 70852 9676
rect 70818 9068 70852 9084
rect 71836 9660 71870 9676
rect 71836 9068 71870 9084
rect 72854 9660 72888 9676
rect 72854 9068 72888 9084
rect 73872 9660 73906 9676
rect 73872 9068 73906 9084
rect 74890 9660 74924 9676
rect 74890 9068 74924 9084
rect 51142 8988 51158 9022
rect 51714 8988 51730 9022
rect 51914 9018 51996 9042
rect 62140 9034 62200 9038
rect 63168 9034 63228 9036
rect 65212 9034 65272 9038
rect 54762 9000 54778 9034
rect 55334 9000 55350 9034
rect 55780 9000 55796 9034
rect 56352 9000 56368 9034
rect 56798 9000 56814 9034
rect 57370 9000 57386 9034
rect 57816 9000 57832 9034
rect 58388 9000 58404 9034
rect 58834 9000 58850 9034
rect 59406 9000 59422 9034
rect 59852 9000 59868 9034
rect 60424 9000 60440 9034
rect 60870 9000 60886 9034
rect 61442 9000 61458 9034
rect 61888 9000 61904 9034
rect 62460 9000 62476 9034
rect 62906 9000 62922 9034
rect 63478 9000 63494 9034
rect 63924 9000 63940 9034
rect 64496 9000 64512 9034
rect 64942 9000 64958 9034
rect 65514 9000 65530 9034
rect 65960 9000 65976 9034
rect 66532 9000 66548 9034
rect 66978 9000 66994 9034
rect 67550 9000 67566 9034
rect 67996 9000 68012 9034
rect 68568 9000 68584 9034
rect 69014 9000 69030 9034
rect 69586 9000 69602 9034
rect 70032 9000 70048 9034
rect 70604 9000 70620 9034
rect 71050 9000 71066 9034
rect 71622 9000 71638 9034
rect 72068 9000 72084 9034
rect 72640 9000 72656 9034
rect 73086 9000 73102 9034
rect 73658 9000 73674 9034
rect 74104 9000 74120 9034
rect 74676 9000 74692 9034
rect 42766 8938 42800 8954
rect 42766 8346 42800 8362
rect 43784 8938 43818 8954
rect 43784 8346 43818 8362
rect 44802 8938 44836 8954
rect 44802 8346 44836 8362
rect 45820 8938 45854 8954
rect 45820 8346 45854 8362
rect 46838 8938 46872 8954
rect 46838 8346 46872 8362
rect 47856 8938 47890 8954
rect 47856 8346 47890 8362
rect 48874 8938 48908 8954
rect 48874 8346 48908 8362
rect 49892 8938 49926 8954
rect 49892 8346 49926 8362
rect 50910 8938 50944 8954
rect 50910 8346 50944 8362
rect 51928 8938 51962 8954
rect 55024 8794 55106 8818
rect 55024 8760 55048 8794
rect 55082 8760 55106 8794
rect 55024 8736 55106 8760
rect 56042 8794 56124 8818
rect 56042 8760 56066 8794
rect 56100 8760 56124 8794
rect 56042 8736 56124 8760
rect 57060 8794 57142 8818
rect 57060 8760 57084 8794
rect 57118 8760 57142 8794
rect 57060 8736 57142 8760
rect 58078 8794 58160 8818
rect 58078 8760 58102 8794
rect 58136 8760 58160 8794
rect 58078 8736 58160 8760
rect 59096 8794 59178 8818
rect 59096 8760 59120 8794
rect 59154 8760 59178 8794
rect 59096 8736 59178 8760
rect 60114 8794 60196 8818
rect 60114 8760 60138 8794
rect 60172 8760 60196 8794
rect 60114 8736 60196 8760
rect 61132 8794 61214 8818
rect 61132 8760 61156 8794
rect 61190 8760 61214 8794
rect 61132 8736 61214 8760
rect 62150 8794 62232 8818
rect 62150 8760 62174 8794
rect 62208 8760 62232 8794
rect 62150 8736 62232 8760
rect 63168 8794 63250 8818
rect 63168 8760 63192 8794
rect 63226 8760 63250 8794
rect 63168 8736 63250 8760
rect 64186 8794 64268 8818
rect 64186 8760 64210 8794
rect 64244 8760 64268 8794
rect 64186 8736 64268 8760
rect 65204 8794 65286 8818
rect 65204 8760 65228 8794
rect 65262 8760 65286 8794
rect 65204 8736 65286 8760
rect 66222 8794 66304 8818
rect 66222 8760 66246 8794
rect 66280 8760 66304 8794
rect 66222 8736 66304 8760
rect 67240 8794 67322 8818
rect 67240 8760 67264 8794
rect 67298 8760 67322 8794
rect 67240 8736 67322 8760
rect 68258 8794 68340 8818
rect 68258 8760 68282 8794
rect 68316 8760 68340 8794
rect 68258 8736 68340 8760
rect 69276 8794 69358 8818
rect 69276 8760 69300 8794
rect 69334 8760 69358 8794
rect 69276 8736 69358 8760
rect 70294 8794 70376 8818
rect 70294 8760 70318 8794
rect 70352 8760 70376 8794
rect 70294 8736 70376 8760
rect 71312 8794 71394 8818
rect 71312 8760 71336 8794
rect 71370 8760 71394 8794
rect 71312 8736 71394 8760
rect 72330 8794 72412 8818
rect 72330 8760 72354 8794
rect 72388 8760 72412 8794
rect 72330 8736 72412 8760
rect 73348 8794 73430 8818
rect 73348 8760 73372 8794
rect 73406 8760 73430 8794
rect 73348 8736 73430 8760
rect 74366 8794 74448 8818
rect 74366 8760 74390 8794
rect 74424 8760 74448 8794
rect 74366 8736 74448 8760
rect 54762 8476 54778 8510
rect 55334 8476 55350 8510
rect 55780 8476 55796 8510
rect 56352 8476 56368 8510
rect 56798 8476 56814 8510
rect 57370 8476 57386 8510
rect 57816 8476 57832 8510
rect 58388 8476 58404 8510
rect 58834 8476 58850 8510
rect 59406 8476 59422 8510
rect 59852 8476 59868 8510
rect 60424 8476 60440 8510
rect 60870 8476 60886 8510
rect 61442 8476 61458 8510
rect 61888 8476 61904 8510
rect 62460 8476 62476 8510
rect 62906 8476 62922 8510
rect 63478 8476 63494 8510
rect 63924 8476 63940 8510
rect 64496 8476 64512 8510
rect 64942 8476 64958 8510
rect 65514 8476 65530 8510
rect 65960 8476 65976 8510
rect 66532 8476 66548 8510
rect 66978 8476 66994 8510
rect 67550 8476 67566 8510
rect 67996 8476 68012 8510
rect 68568 8476 68584 8510
rect 69014 8476 69030 8510
rect 69586 8476 69602 8510
rect 70032 8476 70048 8510
rect 70604 8476 70620 8510
rect 71050 8476 71066 8510
rect 71622 8476 71638 8510
rect 72068 8476 72084 8510
rect 72640 8476 72656 8510
rect 73086 8476 73102 8510
rect 73658 8476 73674 8510
rect 74104 8476 74120 8510
rect 74676 8476 74692 8510
rect 51928 8346 51962 8362
rect 54530 8426 54564 8442
rect 43258 8312 43318 8314
rect 44284 8312 44344 8316
rect 45298 8312 45358 8316
rect 46318 8312 46378 8314
rect 47340 8312 47400 8314
rect 49372 8312 49432 8316
rect 50388 8312 50448 8316
rect 51408 8312 51468 8314
rect 42742 8258 42824 8282
rect 42998 8278 43014 8312
rect 43570 8278 43586 8312
rect 42742 8224 42766 8258
rect 42800 8224 42824 8258
rect 42742 8200 42824 8224
rect 43760 8258 43842 8282
rect 44016 8278 44032 8312
rect 44588 8278 44604 8312
rect 43760 8224 43784 8258
rect 43818 8224 43842 8258
rect 42998 8170 43014 8204
rect 43570 8170 43586 8204
rect 43760 8200 43842 8224
rect 44778 8258 44860 8282
rect 45034 8278 45050 8312
rect 45606 8278 45622 8312
rect 44778 8224 44802 8258
rect 44836 8224 44860 8258
rect 44016 8170 44032 8204
rect 44588 8170 44604 8204
rect 44778 8200 44860 8224
rect 45796 8258 45878 8282
rect 46052 8278 46068 8312
rect 46624 8278 46640 8312
rect 45796 8224 45820 8258
rect 45854 8224 45878 8258
rect 45034 8170 45050 8204
rect 45606 8170 45622 8204
rect 45796 8200 45878 8224
rect 46814 8258 46896 8282
rect 47070 8278 47086 8312
rect 47642 8278 47658 8312
rect 46814 8224 46838 8258
rect 46872 8224 46896 8258
rect 46052 8170 46068 8204
rect 46624 8170 46640 8204
rect 46814 8200 46896 8224
rect 47832 8258 47914 8282
rect 48088 8278 48104 8312
rect 48660 8278 48676 8312
rect 47832 8224 47856 8258
rect 47890 8224 47914 8258
rect 47070 8170 47086 8204
rect 47642 8170 47658 8204
rect 47832 8200 47914 8224
rect 48850 8258 48932 8282
rect 49106 8278 49122 8312
rect 49678 8278 49694 8312
rect 48850 8224 48874 8258
rect 48908 8224 48932 8258
rect 48088 8170 48104 8204
rect 48660 8170 48676 8204
rect 48850 8200 48932 8224
rect 49868 8258 49950 8282
rect 50124 8278 50140 8312
rect 50696 8278 50712 8312
rect 49868 8224 49892 8258
rect 49926 8224 49950 8258
rect 49106 8170 49122 8204
rect 49678 8170 49694 8204
rect 49868 8200 49950 8224
rect 50886 8258 50968 8282
rect 51142 8278 51158 8312
rect 51714 8278 51730 8312
rect 50886 8224 50910 8258
rect 50944 8224 50968 8258
rect 50124 8170 50140 8204
rect 50696 8170 50712 8204
rect 50886 8200 50968 8224
rect 51914 8258 51996 8282
rect 51914 8224 51938 8258
rect 51972 8224 51996 8258
rect 51142 8170 51158 8204
rect 51714 8170 51730 8204
rect 51914 8200 51996 8224
rect 42766 8120 42800 8136
rect 42766 7528 42800 7544
rect 43784 8120 43818 8136
rect 43784 7528 43818 7544
rect 44802 8120 44836 8136
rect 44802 7528 44836 7544
rect 45820 8120 45854 8136
rect 45820 7528 45854 7544
rect 46838 8120 46872 8136
rect 46838 7528 46872 7544
rect 47856 8120 47890 8136
rect 47856 7528 47890 7544
rect 48874 8120 48908 8136
rect 48874 7528 48908 7544
rect 49892 8120 49926 8136
rect 49892 7528 49926 7544
rect 50910 8120 50944 8136
rect 50910 7528 50944 7544
rect 51928 8120 51962 8136
rect 54530 7834 54564 7850
rect 55548 8426 55582 8442
rect 55548 7834 55582 7850
rect 56566 8426 56600 8442
rect 56566 7834 56600 7850
rect 57584 8426 57618 8442
rect 57584 7834 57618 7850
rect 58602 8426 58636 8442
rect 58602 7834 58636 7850
rect 59620 8426 59654 8442
rect 59620 7834 59654 7850
rect 60638 8426 60672 8442
rect 60638 7834 60672 7850
rect 61656 8426 61690 8442
rect 61656 7834 61690 7850
rect 62674 8426 62708 8442
rect 62674 7834 62708 7850
rect 63692 8426 63726 8442
rect 63692 7834 63726 7850
rect 64710 8426 64744 8442
rect 64710 7834 64744 7850
rect 65728 8426 65762 8442
rect 65728 7834 65762 7850
rect 66746 8426 66780 8442
rect 66746 7834 66780 7850
rect 67764 8426 67798 8442
rect 67764 7834 67798 7850
rect 68782 8426 68816 8442
rect 68782 7834 68816 7850
rect 69800 8426 69834 8442
rect 69800 7834 69834 7850
rect 70818 8426 70852 8442
rect 70818 7834 70852 7850
rect 71836 8426 71870 8442
rect 71836 7834 71870 7850
rect 72854 8426 72888 8442
rect 72854 7834 72888 7850
rect 73872 8426 73906 8442
rect 73872 7834 73906 7850
rect 74890 8426 74924 8442
rect 74890 7834 74924 7850
rect 54762 7766 54778 7800
rect 55334 7766 55350 7800
rect 55780 7766 55796 7800
rect 56352 7766 56368 7800
rect 56798 7766 56814 7800
rect 57370 7766 57386 7800
rect 57816 7766 57832 7800
rect 58388 7766 58404 7800
rect 58834 7766 58850 7800
rect 59406 7766 59422 7800
rect 59852 7766 59868 7800
rect 60424 7766 60440 7800
rect 60870 7766 60886 7800
rect 61442 7766 61458 7800
rect 61888 7766 61904 7800
rect 62460 7766 62476 7800
rect 62906 7766 62922 7800
rect 63478 7766 63494 7800
rect 63924 7766 63940 7800
rect 64496 7766 64512 7800
rect 64942 7766 64958 7800
rect 65514 7766 65530 7800
rect 65960 7766 65976 7800
rect 66532 7766 66548 7800
rect 66978 7766 66994 7800
rect 67550 7766 67566 7800
rect 67996 7766 68012 7800
rect 68568 7766 68584 7800
rect 69014 7766 69030 7800
rect 69586 7766 69602 7800
rect 70032 7766 70048 7800
rect 70604 7766 70620 7800
rect 71050 7766 71066 7800
rect 71622 7766 71638 7800
rect 72068 7766 72084 7800
rect 72640 7766 72656 7800
rect 73086 7766 73102 7800
rect 73658 7766 73674 7800
rect 74104 7766 74120 7800
rect 74676 7766 74692 7800
rect 51928 7528 51962 7544
rect 55036 7558 55118 7582
rect 55036 7524 55060 7558
rect 55094 7524 55118 7558
rect 55036 7500 55118 7524
rect 56054 7558 56136 7582
rect 56054 7524 56078 7558
rect 56112 7524 56136 7558
rect 56054 7500 56136 7524
rect 57072 7558 57154 7582
rect 57072 7524 57096 7558
rect 57130 7524 57154 7558
rect 57072 7500 57154 7524
rect 58090 7558 58172 7582
rect 58090 7524 58114 7558
rect 58148 7524 58172 7558
rect 58090 7500 58172 7524
rect 59108 7558 59190 7582
rect 59108 7524 59132 7558
rect 59166 7524 59190 7558
rect 59108 7500 59190 7524
rect 60126 7558 60208 7582
rect 60126 7524 60150 7558
rect 60184 7524 60208 7558
rect 60126 7500 60208 7524
rect 61144 7558 61226 7582
rect 61144 7524 61168 7558
rect 61202 7524 61226 7558
rect 61144 7500 61226 7524
rect 62162 7558 62244 7582
rect 62162 7524 62186 7558
rect 62220 7524 62244 7558
rect 62162 7500 62244 7524
rect 63180 7558 63262 7582
rect 63180 7524 63204 7558
rect 63238 7524 63262 7558
rect 63180 7500 63262 7524
rect 64198 7558 64280 7582
rect 64198 7524 64222 7558
rect 64256 7524 64280 7558
rect 64198 7500 64280 7524
rect 65216 7558 65298 7582
rect 65216 7524 65240 7558
rect 65274 7524 65298 7558
rect 65216 7500 65298 7524
rect 66234 7558 66316 7582
rect 66234 7524 66258 7558
rect 66292 7524 66316 7558
rect 66234 7500 66316 7524
rect 67252 7558 67334 7582
rect 67252 7524 67276 7558
rect 67310 7524 67334 7558
rect 67252 7500 67334 7524
rect 68270 7558 68352 7582
rect 68270 7524 68294 7558
rect 68328 7524 68352 7558
rect 68270 7500 68352 7524
rect 69288 7558 69370 7582
rect 69288 7524 69312 7558
rect 69346 7524 69370 7558
rect 69288 7500 69370 7524
rect 70306 7558 70388 7582
rect 70306 7524 70330 7558
rect 70364 7524 70388 7558
rect 70306 7500 70388 7524
rect 71324 7558 71406 7582
rect 71324 7524 71348 7558
rect 71382 7524 71406 7558
rect 71324 7500 71406 7524
rect 72342 7558 72424 7582
rect 72342 7524 72366 7558
rect 72400 7524 72424 7558
rect 72342 7500 72424 7524
rect 73360 7558 73442 7582
rect 73360 7524 73384 7558
rect 73418 7524 73442 7558
rect 73360 7500 73442 7524
rect 74378 7558 74460 7582
rect 74378 7524 74402 7558
rect 74436 7524 74460 7558
rect 74378 7500 74460 7524
rect 42998 7460 43014 7494
rect 43570 7460 43586 7494
rect 44016 7460 44032 7494
rect 44588 7460 44604 7494
rect 45034 7460 45050 7494
rect 45606 7460 45622 7494
rect 46052 7460 46068 7494
rect 46624 7460 46640 7494
rect 47070 7460 47086 7494
rect 47642 7460 47658 7494
rect 48088 7460 48104 7494
rect 48660 7460 48676 7494
rect 49106 7460 49122 7494
rect 49678 7460 49694 7494
rect 50124 7460 50140 7494
rect 50696 7460 50712 7494
rect 51142 7460 51158 7494
rect 51714 7460 51730 7494
rect 42730 7364 42812 7388
rect 42730 7330 42754 7364
rect 42788 7330 42812 7364
rect 42730 7306 42812 7330
rect 43748 7364 43830 7388
rect 43748 7330 43772 7364
rect 43806 7330 43830 7364
rect 43748 7306 43830 7330
rect 44766 7364 44848 7388
rect 44766 7330 44790 7364
rect 44824 7330 44848 7364
rect 44766 7306 44848 7330
rect 45784 7364 45866 7388
rect 45784 7330 45808 7364
rect 45842 7330 45866 7364
rect 45784 7306 45866 7330
rect 46802 7364 46884 7388
rect 46802 7330 46826 7364
rect 46860 7330 46884 7364
rect 46802 7306 46884 7330
rect 47820 7364 47902 7388
rect 47820 7330 47844 7364
rect 47878 7330 47902 7364
rect 47820 7306 47902 7330
rect 48838 7364 48920 7388
rect 48838 7330 48862 7364
rect 48896 7330 48920 7364
rect 48838 7306 48920 7330
rect 49856 7364 49938 7388
rect 49856 7330 49880 7364
rect 49914 7330 49938 7364
rect 49856 7306 49938 7330
rect 50874 7364 50956 7388
rect 50874 7330 50898 7364
rect 50932 7330 50956 7364
rect 50874 7306 50956 7330
rect 51902 7364 51984 7388
rect 51902 7330 51926 7364
rect 51960 7330 51984 7364
rect 51902 7306 51984 7330
rect 54762 7244 54778 7278
rect 55334 7244 55350 7278
rect 55780 7244 55796 7278
rect 56352 7244 56368 7278
rect 56798 7244 56814 7278
rect 57370 7244 57386 7278
rect 57816 7244 57832 7278
rect 58388 7244 58404 7278
rect 58834 7244 58850 7278
rect 59406 7244 59422 7278
rect 59852 7244 59868 7278
rect 60424 7244 60440 7278
rect 60870 7244 60886 7278
rect 61442 7244 61458 7278
rect 61888 7244 61904 7278
rect 62460 7244 62476 7278
rect 62906 7244 62922 7278
rect 63478 7244 63494 7278
rect 63924 7244 63940 7278
rect 64496 7244 64512 7278
rect 64942 7244 64958 7278
rect 65514 7244 65530 7278
rect 65960 7244 65976 7278
rect 66532 7244 66548 7278
rect 66978 7244 66994 7278
rect 67550 7244 67566 7278
rect 67996 7244 68012 7278
rect 68568 7244 68584 7278
rect 69014 7244 69030 7278
rect 69586 7244 69602 7278
rect 70032 7244 70048 7278
rect 70604 7244 70620 7278
rect 71050 7244 71066 7278
rect 71622 7244 71638 7278
rect 72068 7244 72084 7278
rect 72640 7244 72656 7278
rect 73086 7244 73102 7278
rect 73658 7244 73674 7278
rect 74104 7244 74120 7278
rect 74676 7244 74692 7278
rect 54530 7194 54564 7210
rect 54530 6602 54564 6618
rect 55548 7194 55582 7210
rect 55548 6602 55582 6618
rect 56566 7194 56600 7210
rect 56566 6602 56600 6618
rect 57584 7194 57618 7210
rect 57584 6602 57618 6618
rect 58602 7194 58636 7210
rect 58602 6602 58636 6618
rect 59620 7194 59654 7210
rect 59620 6602 59654 6618
rect 60638 7194 60672 7210
rect 60638 6602 60672 6618
rect 61656 7194 61690 7210
rect 61656 6602 61690 6618
rect 62674 7194 62708 7210
rect 62674 6602 62708 6618
rect 63692 7194 63726 7210
rect 63692 6602 63726 6618
rect 64710 7194 64744 7210
rect 64710 6602 64744 6618
rect 65728 7194 65762 7210
rect 65728 6602 65762 6618
rect 66746 7194 66780 7210
rect 66746 6602 66780 6618
rect 67764 7194 67798 7210
rect 67764 6602 67798 6618
rect 68782 7194 68816 7210
rect 68782 6602 68816 6618
rect 69800 7194 69834 7210
rect 69800 6602 69834 6618
rect 70818 7194 70852 7210
rect 70818 6602 70852 6618
rect 71836 7194 71870 7210
rect 71836 6602 71870 6618
rect 72854 7194 72888 7210
rect 72854 6602 72888 6618
rect 73872 7194 73906 7210
rect 73872 6602 73906 6618
rect 74890 7194 74924 7210
rect 74890 6602 74924 6618
rect 63180 6568 63240 6570
rect 65224 6568 65284 6572
rect 73358 6568 73418 6570
rect 54762 6534 54778 6568
rect 55334 6534 55350 6568
rect 55780 6534 55796 6568
rect 56352 6534 56368 6568
rect 56798 6534 56814 6568
rect 57370 6534 57386 6568
rect 57816 6534 57832 6568
rect 58388 6534 58404 6568
rect 58834 6534 58850 6568
rect 59406 6534 59422 6568
rect 59852 6534 59868 6568
rect 60424 6534 60440 6568
rect 60870 6534 60886 6568
rect 61442 6534 61458 6568
rect 61888 6534 61904 6568
rect 62460 6534 62476 6568
rect 62906 6534 62922 6568
rect 63478 6534 63494 6568
rect 63924 6534 63940 6568
rect 64496 6534 64512 6568
rect 64942 6534 64958 6568
rect 65514 6534 65530 6568
rect 65960 6534 65976 6568
rect 66532 6534 66548 6568
rect 66978 6534 66994 6568
rect 67550 6534 67566 6568
rect 67996 6534 68012 6568
rect 68568 6534 68584 6568
rect 69014 6534 69030 6568
rect 69586 6534 69602 6568
rect 70032 6534 70048 6568
rect 70604 6534 70620 6568
rect 71050 6534 71066 6568
rect 71622 6534 71638 6568
rect 72068 6534 72084 6568
rect 72640 6534 72656 6568
rect 73086 6534 73102 6568
rect 73658 6534 73674 6568
rect 74104 6534 74120 6568
rect 74676 6534 74692 6568
rect 41934 6416 42016 6440
rect 41934 6382 41958 6416
rect 41992 6382 42016 6416
rect 41934 6358 42016 6382
rect 42952 6416 43034 6440
rect 42952 6382 42976 6416
rect 43010 6382 43034 6416
rect 42952 6358 43034 6382
rect 43970 6416 44052 6440
rect 43970 6382 43994 6416
rect 44028 6382 44052 6416
rect 43970 6358 44052 6382
rect 44988 6416 45070 6440
rect 44988 6382 45012 6416
rect 45046 6382 45070 6416
rect 44988 6358 45070 6382
rect 46006 6416 46088 6440
rect 46006 6382 46030 6416
rect 46064 6382 46088 6416
rect 46006 6358 46088 6382
rect 47024 6416 47106 6440
rect 47024 6382 47048 6416
rect 47082 6382 47106 6416
rect 47024 6358 47106 6382
rect 48042 6416 48124 6440
rect 48042 6382 48066 6416
rect 48100 6382 48124 6416
rect 48042 6358 48124 6382
rect 49060 6416 49142 6440
rect 49060 6382 49084 6416
rect 49118 6382 49142 6416
rect 49060 6358 49142 6382
rect 50078 6416 50160 6440
rect 50078 6382 50102 6416
rect 50136 6382 50160 6416
rect 50078 6358 50160 6382
rect 51096 6416 51178 6440
rect 51096 6382 51120 6416
rect 51154 6382 51178 6416
rect 51096 6358 51178 6382
rect 52114 6416 52196 6440
rect 52114 6382 52138 6416
rect 52172 6382 52196 6416
rect 52114 6358 52196 6382
rect 55036 6310 55118 6334
rect 55036 6276 55060 6310
rect 55094 6276 55118 6310
rect 55036 6252 55118 6276
rect 56054 6310 56136 6334
rect 56054 6276 56078 6310
rect 56112 6276 56136 6310
rect 56054 6252 56136 6276
rect 57072 6310 57154 6334
rect 57072 6276 57096 6310
rect 57130 6276 57154 6310
rect 57072 6252 57154 6276
rect 58090 6310 58172 6334
rect 58090 6276 58114 6310
rect 58148 6276 58172 6310
rect 58090 6252 58172 6276
rect 59108 6310 59190 6334
rect 59108 6276 59132 6310
rect 59166 6276 59190 6310
rect 59108 6252 59190 6276
rect 60126 6310 60208 6334
rect 60126 6276 60150 6310
rect 60184 6276 60208 6310
rect 60126 6252 60208 6276
rect 61144 6310 61226 6334
rect 61144 6276 61168 6310
rect 61202 6276 61226 6310
rect 61144 6252 61226 6276
rect 62162 6310 62244 6334
rect 62162 6276 62186 6310
rect 62220 6276 62244 6310
rect 62162 6252 62244 6276
rect 63180 6310 63262 6334
rect 63180 6276 63204 6310
rect 63238 6276 63262 6310
rect 63180 6252 63262 6276
rect 64198 6310 64280 6334
rect 64198 6276 64222 6310
rect 64256 6276 64280 6310
rect 64198 6252 64280 6276
rect 65216 6310 65298 6334
rect 65216 6276 65240 6310
rect 65274 6276 65298 6310
rect 65216 6252 65298 6276
rect 66234 6310 66316 6334
rect 66234 6276 66258 6310
rect 66292 6276 66316 6310
rect 66234 6252 66316 6276
rect 67252 6310 67334 6334
rect 67252 6276 67276 6310
rect 67310 6276 67334 6310
rect 67252 6252 67334 6276
rect 68270 6310 68352 6334
rect 68270 6276 68294 6310
rect 68328 6276 68352 6310
rect 68270 6252 68352 6276
rect 69288 6310 69370 6334
rect 69288 6276 69312 6310
rect 69346 6276 69370 6310
rect 69288 6252 69370 6276
rect 70306 6310 70388 6334
rect 70306 6276 70330 6310
rect 70364 6276 70388 6310
rect 70306 6252 70388 6276
rect 71324 6310 71406 6334
rect 71324 6276 71348 6310
rect 71382 6276 71406 6310
rect 71324 6252 71406 6276
rect 72342 6310 72424 6334
rect 72342 6276 72366 6310
rect 72400 6276 72424 6310
rect 72342 6252 72424 6276
rect 73360 6310 73442 6334
rect 73360 6276 73384 6310
rect 73418 6276 73442 6310
rect 73360 6252 73442 6276
rect 74378 6310 74460 6334
rect 74378 6276 74402 6310
rect 74436 6276 74460 6310
rect 74378 6252 74460 6276
rect 41674 6146 41690 6180
rect 42246 6146 42262 6180
rect 42692 6146 42708 6180
rect 43264 6146 43280 6180
rect 43710 6146 43726 6180
rect 44282 6146 44298 6180
rect 44728 6146 44744 6180
rect 45300 6146 45316 6180
rect 45746 6146 45762 6180
rect 46318 6146 46334 6180
rect 46764 6146 46780 6180
rect 47336 6146 47352 6180
rect 47782 6146 47798 6180
rect 48354 6146 48370 6180
rect 48800 6146 48816 6180
rect 49372 6146 49388 6180
rect 49818 6146 49834 6180
rect 50390 6146 50406 6180
rect 50836 6146 50852 6180
rect 51408 6146 51424 6180
rect 51854 6146 51870 6180
rect 52426 6146 52442 6180
rect 41442 6096 41476 6112
rect 41442 5504 41476 5520
rect 42460 6096 42494 6112
rect 42460 5504 42494 5520
rect 43478 6096 43512 6112
rect 43478 5504 43512 5520
rect 44496 6096 44530 6112
rect 44496 5504 44530 5520
rect 45514 6096 45548 6112
rect 45514 5504 45548 5520
rect 46532 6096 46566 6112
rect 46532 5504 46566 5520
rect 47550 6096 47584 6112
rect 47550 5504 47584 5520
rect 48568 6096 48602 6112
rect 48568 5504 48602 5520
rect 49586 6096 49620 6112
rect 49586 5504 49620 5520
rect 50604 6096 50638 6112
rect 50604 5504 50638 5520
rect 51622 6096 51656 6112
rect 51622 5504 51656 5520
rect 52640 6096 52674 6112
rect 54762 6010 54778 6044
rect 55334 6010 55350 6044
rect 55780 6010 55796 6044
rect 56352 6010 56368 6044
rect 56798 6010 56814 6044
rect 57370 6010 57386 6044
rect 57816 6010 57832 6044
rect 58388 6010 58404 6044
rect 58834 6010 58850 6044
rect 59406 6010 59422 6044
rect 59852 6010 59868 6044
rect 60424 6010 60440 6044
rect 60870 6010 60886 6044
rect 61442 6010 61458 6044
rect 61888 6010 61904 6044
rect 62460 6010 62476 6044
rect 62906 6010 62922 6044
rect 63478 6010 63494 6044
rect 63924 6010 63940 6044
rect 64496 6010 64512 6044
rect 64942 6010 64958 6044
rect 65514 6010 65530 6044
rect 65960 6010 65976 6044
rect 66532 6010 66548 6044
rect 66978 6010 66994 6044
rect 67550 6010 67566 6044
rect 67996 6010 68012 6044
rect 68568 6010 68584 6044
rect 69014 6010 69030 6044
rect 69586 6010 69602 6044
rect 70032 6010 70048 6044
rect 70604 6010 70620 6044
rect 71050 6010 71066 6044
rect 71622 6010 71638 6044
rect 72068 6010 72084 6044
rect 72640 6010 72656 6044
rect 73086 6010 73102 6044
rect 73658 6010 73674 6044
rect 74104 6010 74120 6044
rect 74676 6010 74692 6044
rect 52640 5504 52674 5520
rect 54530 5960 54564 5976
rect 41674 5436 41690 5470
rect 42246 5436 42262 5470
rect 42692 5436 42708 5470
rect 43264 5436 43280 5470
rect 43710 5436 43726 5470
rect 44282 5436 44298 5470
rect 44728 5436 44744 5470
rect 45300 5436 45316 5470
rect 45746 5436 45762 5470
rect 46318 5436 46334 5470
rect 46764 5436 46780 5470
rect 47336 5436 47352 5470
rect 47782 5436 47798 5470
rect 48354 5436 48370 5470
rect 48800 5436 48816 5470
rect 49372 5436 49388 5470
rect 49818 5436 49834 5470
rect 50390 5436 50406 5470
rect 50836 5436 50852 5470
rect 51408 5436 51424 5470
rect 51854 5436 51870 5470
rect 52426 5436 52442 5470
rect 54530 5368 54564 5384
rect 55548 5960 55582 5976
rect 55548 5368 55582 5384
rect 56566 5960 56600 5976
rect 56566 5368 56600 5384
rect 57584 5960 57618 5976
rect 57584 5368 57618 5384
rect 58602 5960 58636 5976
rect 58602 5368 58636 5384
rect 59620 5960 59654 5976
rect 59620 5368 59654 5384
rect 60638 5960 60672 5976
rect 60638 5368 60672 5384
rect 61656 5960 61690 5976
rect 61656 5368 61690 5384
rect 62674 5960 62708 5976
rect 62674 5368 62708 5384
rect 63692 5960 63726 5976
rect 63692 5368 63726 5384
rect 64710 5960 64744 5976
rect 64710 5368 64744 5384
rect 65728 5960 65762 5976
rect 65728 5368 65762 5384
rect 66746 5960 66780 5976
rect 66746 5368 66780 5384
rect 67764 5960 67798 5976
rect 67764 5368 67798 5384
rect 68782 5960 68816 5976
rect 68782 5368 68816 5384
rect 69800 5960 69834 5976
rect 69800 5368 69834 5384
rect 70818 5960 70852 5976
rect 70818 5368 70852 5384
rect 71836 5960 71870 5976
rect 71836 5368 71870 5384
rect 72854 5960 72888 5976
rect 72854 5368 72888 5384
rect 73872 5960 73906 5976
rect 73872 5368 73906 5384
rect 74890 5960 74924 5976
rect 74890 5368 74924 5384
rect 57056 5334 57116 5338
rect 54762 5300 54778 5334
rect 55334 5300 55350 5334
rect 55780 5300 55796 5334
rect 56352 5300 56368 5334
rect 56798 5300 56814 5334
rect 57370 5300 57386 5334
rect 57816 5300 57832 5334
rect 58388 5300 58404 5334
rect 58834 5300 58850 5334
rect 59406 5300 59422 5334
rect 59852 5300 59868 5334
rect 60424 5300 60440 5334
rect 60870 5300 60886 5334
rect 61442 5300 61458 5334
rect 61888 5300 61904 5334
rect 62460 5300 62476 5334
rect 62906 5300 62922 5334
rect 63478 5300 63494 5334
rect 63924 5300 63940 5334
rect 64496 5300 64512 5334
rect 64942 5300 64958 5334
rect 65514 5300 65530 5334
rect 65960 5300 65976 5334
rect 66532 5300 66548 5334
rect 66978 5300 66994 5334
rect 67550 5300 67566 5334
rect 67996 5300 68012 5334
rect 68568 5300 68584 5334
rect 69014 5300 69030 5334
rect 69586 5300 69602 5334
rect 70032 5300 70048 5334
rect 70604 5300 70620 5334
rect 71050 5300 71066 5334
rect 71622 5300 71638 5334
rect 72068 5300 72084 5334
rect 72640 5300 72656 5334
rect 73086 5300 73102 5334
rect 73658 5300 73674 5334
rect 74104 5300 74120 5334
rect 74676 5300 74692 5334
rect 41946 5274 42028 5298
rect 41946 5240 41970 5274
rect 42004 5240 42028 5274
rect 41946 5216 42028 5240
rect 42964 5274 43046 5298
rect 42964 5240 42988 5274
rect 43022 5240 43046 5274
rect 42964 5216 43046 5240
rect 43982 5274 44064 5298
rect 43982 5240 44006 5274
rect 44040 5240 44064 5274
rect 43982 5216 44064 5240
rect 45000 5274 45082 5298
rect 45000 5240 45024 5274
rect 45058 5240 45082 5274
rect 45000 5216 45082 5240
rect 46018 5274 46100 5298
rect 46018 5240 46042 5274
rect 46076 5240 46100 5274
rect 46018 5216 46100 5240
rect 47036 5274 47118 5298
rect 47036 5240 47060 5274
rect 47094 5240 47118 5274
rect 47036 5216 47118 5240
rect 48054 5274 48136 5298
rect 48054 5240 48078 5274
rect 48112 5240 48136 5274
rect 48054 5216 48136 5240
rect 49072 5274 49154 5298
rect 49072 5240 49096 5274
rect 49130 5240 49154 5274
rect 49072 5216 49154 5240
rect 50090 5274 50172 5298
rect 50090 5240 50114 5274
rect 50148 5240 50172 5274
rect 50090 5216 50172 5240
rect 51108 5274 51190 5298
rect 51108 5240 51132 5274
rect 51166 5240 51190 5274
rect 51108 5216 51190 5240
rect 52126 5274 52208 5298
rect 52126 5240 52150 5274
rect 52184 5240 52208 5274
rect 52126 5216 52208 5240
rect 55012 5074 55094 5098
rect 41674 5034 41690 5068
rect 42246 5034 42262 5068
rect 42692 5034 42708 5068
rect 43264 5034 43280 5068
rect 43710 5034 43726 5068
rect 44282 5034 44298 5068
rect 44728 5034 44744 5068
rect 45300 5034 45316 5068
rect 45746 5034 45762 5068
rect 46318 5034 46334 5068
rect 46764 5034 46780 5068
rect 47336 5034 47352 5068
rect 47782 5034 47798 5068
rect 48354 5034 48370 5068
rect 48800 5034 48816 5068
rect 49372 5034 49388 5068
rect 49818 5034 49834 5068
rect 50390 5034 50406 5068
rect 50836 5034 50852 5068
rect 51408 5034 51424 5068
rect 51854 5034 51870 5068
rect 52426 5034 52442 5068
rect 55012 5040 55036 5074
rect 55070 5040 55094 5074
rect 55012 5016 55094 5040
rect 56030 5074 56112 5098
rect 56030 5040 56054 5074
rect 56088 5040 56112 5074
rect 56030 5016 56112 5040
rect 57048 5074 57130 5098
rect 57048 5040 57072 5074
rect 57106 5040 57130 5074
rect 57048 5016 57130 5040
rect 58066 5074 58148 5098
rect 58066 5040 58090 5074
rect 58124 5040 58148 5074
rect 58066 5016 58148 5040
rect 59084 5074 59166 5098
rect 59084 5040 59108 5074
rect 59142 5040 59166 5074
rect 59084 5016 59166 5040
rect 60102 5074 60184 5098
rect 60102 5040 60126 5074
rect 60160 5040 60184 5074
rect 60102 5016 60184 5040
rect 61120 5074 61202 5098
rect 61120 5040 61144 5074
rect 61178 5040 61202 5074
rect 61120 5016 61202 5040
rect 62138 5074 62220 5098
rect 62138 5040 62162 5074
rect 62196 5040 62220 5074
rect 62138 5016 62220 5040
rect 63156 5074 63238 5098
rect 63156 5040 63180 5074
rect 63214 5040 63238 5074
rect 63156 5016 63238 5040
rect 64174 5074 64256 5098
rect 64174 5040 64198 5074
rect 64232 5040 64256 5074
rect 64174 5016 64256 5040
rect 65192 5074 65274 5098
rect 65192 5040 65216 5074
rect 65250 5040 65274 5074
rect 65192 5016 65274 5040
rect 66210 5074 66292 5098
rect 66210 5040 66234 5074
rect 66268 5040 66292 5074
rect 66210 5016 66292 5040
rect 67228 5074 67310 5098
rect 67228 5040 67252 5074
rect 67286 5040 67310 5074
rect 67228 5016 67310 5040
rect 68246 5074 68328 5098
rect 68246 5040 68270 5074
rect 68304 5040 68328 5074
rect 68246 5016 68328 5040
rect 69264 5074 69346 5098
rect 69264 5040 69288 5074
rect 69322 5040 69346 5074
rect 69264 5016 69346 5040
rect 70282 5074 70364 5098
rect 70282 5040 70306 5074
rect 70340 5040 70364 5074
rect 70282 5016 70364 5040
rect 71300 5074 71382 5098
rect 71300 5040 71324 5074
rect 71358 5040 71382 5074
rect 71300 5016 71382 5040
rect 72318 5074 72400 5098
rect 72318 5040 72342 5074
rect 72376 5040 72400 5074
rect 72318 5016 72400 5040
rect 73336 5074 73418 5098
rect 73336 5040 73360 5074
rect 73394 5040 73418 5074
rect 73336 5016 73418 5040
rect 74354 5074 74436 5098
rect 74354 5040 74378 5074
rect 74412 5040 74436 5074
rect 74354 5016 74436 5040
rect 41442 4984 41476 5000
rect 41442 4392 41476 4408
rect 42460 4984 42494 5000
rect 42460 4392 42494 4408
rect 43478 4984 43512 5000
rect 43478 4392 43512 4408
rect 44496 4984 44530 5000
rect 44496 4392 44530 4408
rect 45514 4984 45548 5000
rect 45514 4392 45548 4408
rect 46532 4984 46566 5000
rect 46532 4392 46566 4408
rect 47550 4984 47584 5000
rect 47550 4392 47584 4408
rect 48568 4984 48602 5000
rect 48568 4392 48602 4408
rect 49586 4984 49620 5000
rect 49586 4392 49620 4408
rect 50604 4984 50638 5000
rect 50604 4392 50638 4408
rect 51622 4984 51656 5000
rect 51622 4392 51656 4408
rect 52640 4984 52674 5000
rect 54762 4776 54778 4810
rect 55334 4776 55350 4810
rect 55780 4776 55796 4810
rect 56352 4776 56368 4810
rect 56798 4776 56814 4810
rect 57370 4776 57386 4810
rect 57816 4776 57832 4810
rect 58388 4776 58404 4810
rect 58834 4776 58850 4810
rect 59406 4776 59422 4810
rect 59852 4776 59868 4810
rect 60424 4776 60440 4810
rect 60870 4776 60886 4810
rect 61442 4776 61458 4810
rect 61888 4776 61904 4810
rect 62460 4776 62476 4810
rect 62906 4776 62922 4810
rect 63478 4776 63494 4810
rect 63924 4776 63940 4810
rect 64496 4776 64512 4810
rect 64942 4776 64958 4810
rect 65514 4776 65530 4810
rect 65960 4776 65976 4810
rect 66532 4776 66548 4810
rect 66978 4776 66994 4810
rect 67550 4776 67566 4810
rect 67996 4776 68012 4810
rect 68568 4776 68584 4810
rect 69014 4776 69030 4810
rect 69586 4776 69602 4810
rect 70032 4776 70048 4810
rect 70604 4776 70620 4810
rect 71050 4776 71066 4810
rect 71622 4776 71638 4810
rect 72068 4776 72084 4810
rect 72640 4776 72656 4810
rect 73086 4776 73102 4810
rect 73658 4776 73674 4810
rect 74104 4776 74120 4810
rect 74676 4776 74692 4810
rect 52640 4392 52674 4408
rect 54530 4726 54564 4742
rect 41674 4324 41690 4358
rect 42246 4324 42262 4358
rect 42692 4324 42708 4358
rect 43264 4324 43280 4358
rect 43710 4324 43726 4358
rect 44282 4324 44298 4358
rect 44728 4324 44744 4358
rect 45300 4324 45316 4358
rect 45746 4324 45762 4358
rect 46318 4324 46334 4358
rect 46764 4324 46780 4358
rect 47336 4324 47352 4358
rect 47782 4324 47798 4358
rect 48354 4324 48370 4358
rect 48800 4324 48816 4358
rect 49372 4324 49388 4358
rect 49818 4324 49834 4358
rect 50390 4324 50406 4358
rect 50836 4324 50852 4358
rect 51408 4324 51424 4358
rect 51854 4324 51870 4358
rect 52426 4324 52442 4358
rect 41924 4166 42006 4190
rect 41924 4132 41948 4166
rect 41982 4132 42006 4166
rect 41924 4108 42006 4132
rect 42942 4166 43024 4190
rect 42942 4132 42966 4166
rect 43000 4132 43024 4166
rect 42942 4108 43024 4132
rect 43960 4166 44042 4190
rect 43960 4132 43984 4166
rect 44018 4132 44042 4166
rect 43960 4108 44042 4132
rect 44978 4166 45060 4190
rect 44978 4132 45002 4166
rect 45036 4132 45060 4166
rect 44978 4108 45060 4132
rect 45996 4166 46078 4190
rect 45996 4132 46020 4166
rect 46054 4132 46078 4166
rect 45996 4108 46078 4132
rect 47014 4166 47096 4190
rect 47014 4132 47038 4166
rect 47072 4132 47096 4166
rect 47014 4108 47096 4132
rect 48032 4166 48114 4190
rect 48032 4132 48056 4166
rect 48090 4132 48114 4166
rect 48032 4108 48114 4132
rect 49050 4166 49132 4190
rect 49050 4132 49074 4166
rect 49108 4132 49132 4166
rect 49050 4108 49132 4132
rect 50068 4166 50150 4190
rect 50068 4132 50092 4166
rect 50126 4132 50150 4166
rect 50068 4108 50150 4132
rect 51086 4166 51168 4190
rect 51086 4132 51110 4166
rect 51144 4132 51168 4166
rect 51086 4108 51168 4132
rect 52104 4166 52186 4190
rect 52104 4132 52128 4166
rect 52162 4132 52186 4166
rect 54530 4134 54564 4150
rect 55548 4726 55582 4742
rect 55548 4134 55582 4150
rect 56566 4726 56600 4742
rect 56566 4134 56600 4150
rect 57584 4726 57618 4742
rect 57584 4134 57618 4150
rect 58602 4726 58636 4742
rect 58602 4134 58636 4150
rect 59620 4726 59654 4742
rect 59620 4134 59654 4150
rect 60638 4726 60672 4742
rect 60638 4134 60672 4150
rect 61656 4726 61690 4742
rect 61656 4134 61690 4150
rect 62674 4726 62708 4742
rect 62674 4134 62708 4150
rect 63692 4726 63726 4742
rect 63692 4134 63726 4150
rect 64710 4726 64744 4742
rect 64710 4134 64744 4150
rect 65728 4726 65762 4742
rect 65728 4134 65762 4150
rect 66746 4726 66780 4742
rect 66746 4134 66780 4150
rect 67764 4726 67798 4742
rect 67764 4134 67798 4150
rect 68782 4726 68816 4742
rect 68782 4134 68816 4150
rect 69800 4726 69834 4742
rect 69800 4134 69834 4150
rect 70818 4726 70852 4742
rect 70818 4134 70852 4150
rect 71836 4726 71870 4742
rect 71836 4134 71870 4150
rect 72854 4726 72888 4742
rect 72854 4134 72888 4150
rect 73872 4726 73906 4742
rect 73872 4134 73906 4150
rect 74890 4726 74924 4742
rect 74890 4134 74924 4150
rect 52104 4108 52186 4132
rect 63180 4100 63240 4102
rect 65224 4100 65284 4104
rect 68262 4100 68322 4104
rect 54762 4066 54778 4100
rect 55334 4066 55350 4100
rect 55780 4066 55796 4100
rect 56352 4066 56368 4100
rect 56798 4066 56814 4100
rect 57370 4066 57386 4100
rect 57816 4066 57832 4100
rect 58388 4066 58404 4100
rect 58834 4066 58850 4100
rect 59406 4066 59422 4100
rect 59852 4066 59868 4100
rect 60424 4066 60440 4100
rect 60870 4066 60886 4100
rect 61442 4066 61458 4100
rect 61888 4066 61904 4100
rect 62460 4066 62476 4100
rect 62906 4066 62922 4100
rect 63478 4066 63494 4100
rect 63924 4066 63940 4100
rect 64496 4066 64512 4100
rect 64942 4066 64958 4100
rect 65514 4066 65530 4100
rect 65960 4066 65976 4100
rect 66532 4066 66548 4100
rect 66978 4066 66994 4100
rect 67550 4066 67566 4100
rect 67996 4066 68012 4100
rect 68568 4066 68584 4100
rect 69014 4066 69030 4100
rect 69586 4066 69602 4100
rect 70032 4066 70048 4100
rect 70604 4066 70620 4100
rect 71050 4066 71066 4100
rect 71622 4066 71638 4100
rect 72068 4066 72084 4100
rect 72640 4066 72656 4100
rect 73086 4066 73102 4100
rect 73658 4066 73674 4100
rect 74104 4066 74120 4100
rect 74676 4066 74692 4100
rect 41674 3922 41690 3956
rect 42246 3922 42262 3956
rect 42692 3922 42708 3956
rect 43264 3922 43280 3956
rect 43710 3922 43726 3956
rect 44282 3922 44298 3956
rect 44728 3922 44744 3956
rect 45300 3922 45316 3956
rect 45746 3922 45762 3956
rect 46318 3922 46334 3956
rect 46764 3922 46780 3956
rect 47336 3922 47352 3956
rect 47782 3922 47798 3956
rect 48354 3922 48370 3956
rect 48800 3922 48816 3956
rect 49372 3922 49388 3956
rect 49818 3922 49834 3956
rect 50390 3922 50406 3956
rect 50836 3922 50852 3956
rect 51408 3922 51424 3956
rect 51854 3922 51870 3956
rect 52426 3922 52442 3956
rect 41442 3872 41476 3888
rect 41442 3280 41476 3296
rect 42460 3872 42494 3888
rect 42460 3280 42494 3296
rect 43478 3872 43512 3888
rect 43478 3280 43512 3296
rect 44496 3872 44530 3888
rect 44496 3280 44530 3296
rect 45514 3872 45548 3888
rect 45514 3280 45548 3296
rect 46532 3872 46566 3888
rect 46532 3280 46566 3296
rect 47550 3872 47584 3888
rect 47550 3280 47584 3296
rect 48568 3872 48602 3888
rect 48568 3280 48602 3296
rect 49586 3872 49620 3888
rect 49586 3280 49620 3296
rect 50604 3872 50638 3888
rect 50604 3280 50638 3296
rect 51622 3872 51656 3888
rect 51622 3280 51656 3296
rect 52640 3872 52674 3888
rect 55024 3850 55106 3874
rect 55024 3816 55048 3850
rect 55082 3816 55106 3850
rect 55024 3792 55106 3816
rect 56042 3850 56124 3874
rect 56042 3816 56066 3850
rect 56100 3816 56124 3850
rect 56042 3792 56124 3816
rect 57060 3850 57142 3874
rect 57060 3816 57084 3850
rect 57118 3816 57142 3850
rect 57060 3792 57142 3816
rect 58078 3850 58160 3874
rect 58078 3816 58102 3850
rect 58136 3816 58160 3850
rect 58078 3792 58160 3816
rect 59096 3850 59178 3874
rect 59096 3816 59120 3850
rect 59154 3816 59178 3850
rect 59096 3792 59178 3816
rect 60114 3850 60196 3874
rect 60114 3816 60138 3850
rect 60172 3816 60196 3850
rect 60114 3792 60196 3816
rect 61132 3850 61214 3874
rect 61132 3816 61156 3850
rect 61190 3816 61214 3850
rect 61132 3792 61214 3816
rect 62150 3850 62232 3874
rect 62150 3816 62174 3850
rect 62208 3816 62232 3850
rect 62150 3792 62232 3816
rect 63168 3850 63250 3874
rect 63168 3816 63192 3850
rect 63226 3816 63250 3850
rect 63168 3792 63250 3816
rect 64186 3850 64268 3874
rect 64186 3816 64210 3850
rect 64244 3816 64268 3850
rect 64186 3792 64268 3816
rect 65204 3850 65286 3874
rect 65204 3816 65228 3850
rect 65262 3816 65286 3850
rect 65204 3792 65286 3816
rect 66222 3850 66304 3874
rect 66222 3816 66246 3850
rect 66280 3816 66304 3850
rect 66222 3792 66304 3816
rect 67240 3850 67322 3874
rect 67240 3816 67264 3850
rect 67298 3816 67322 3850
rect 67240 3792 67322 3816
rect 68258 3850 68340 3874
rect 68258 3816 68282 3850
rect 68316 3816 68340 3850
rect 68258 3792 68340 3816
rect 69276 3850 69358 3874
rect 69276 3816 69300 3850
rect 69334 3816 69358 3850
rect 69276 3792 69358 3816
rect 70294 3850 70376 3874
rect 70294 3816 70318 3850
rect 70352 3816 70376 3850
rect 70294 3792 70376 3816
rect 71312 3850 71394 3874
rect 71312 3816 71336 3850
rect 71370 3816 71394 3850
rect 71312 3792 71394 3816
rect 72330 3850 72412 3874
rect 72330 3816 72354 3850
rect 72388 3816 72412 3850
rect 72330 3792 72412 3816
rect 73348 3850 73430 3874
rect 73348 3816 73372 3850
rect 73406 3816 73430 3850
rect 73348 3792 73430 3816
rect 74366 3850 74448 3874
rect 74366 3816 74390 3850
rect 74424 3816 74448 3850
rect 74366 3792 74448 3816
rect 54762 3544 54778 3578
rect 55334 3544 55350 3578
rect 55780 3544 55796 3578
rect 56352 3544 56368 3578
rect 56798 3544 56814 3578
rect 57370 3544 57386 3578
rect 57816 3544 57832 3578
rect 58388 3544 58404 3578
rect 58834 3544 58850 3578
rect 59406 3544 59422 3578
rect 59852 3544 59868 3578
rect 60424 3544 60440 3578
rect 60870 3544 60886 3578
rect 61442 3544 61458 3578
rect 61888 3544 61904 3578
rect 62460 3544 62476 3578
rect 62906 3544 62922 3578
rect 63478 3544 63494 3578
rect 63924 3544 63940 3578
rect 64496 3544 64512 3578
rect 64942 3544 64958 3578
rect 65514 3544 65530 3578
rect 65960 3544 65976 3578
rect 66532 3544 66548 3578
rect 66978 3544 66994 3578
rect 67550 3544 67566 3578
rect 67996 3544 68012 3578
rect 68568 3544 68584 3578
rect 69014 3544 69030 3578
rect 69586 3544 69602 3578
rect 70032 3544 70048 3578
rect 70604 3544 70620 3578
rect 71050 3544 71066 3578
rect 71622 3544 71638 3578
rect 72068 3544 72084 3578
rect 72640 3544 72656 3578
rect 73086 3544 73102 3578
rect 73658 3544 73674 3578
rect 74104 3544 74120 3578
rect 74676 3544 74692 3578
rect 58084 3542 58144 3544
rect 52640 3280 52674 3296
rect 54530 3494 54564 3510
rect 41674 3212 41690 3246
rect 42246 3212 42262 3246
rect 42692 3212 42708 3246
rect 43264 3212 43280 3246
rect 43710 3212 43726 3246
rect 44282 3212 44298 3246
rect 44728 3212 44744 3246
rect 45300 3212 45316 3246
rect 45746 3212 45762 3246
rect 46318 3212 46334 3246
rect 46764 3212 46780 3246
rect 47336 3212 47352 3246
rect 47782 3212 47798 3246
rect 48354 3212 48370 3246
rect 48800 3212 48816 3246
rect 49372 3212 49388 3246
rect 49818 3212 49834 3246
rect 50390 3212 50406 3246
rect 50836 3212 50852 3246
rect 51408 3212 51424 3246
rect 51854 3212 51870 3246
rect 52426 3212 52442 3246
rect 41924 3060 42006 3084
rect 41924 3026 41948 3060
rect 41982 3026 42006 3060
rect 41924 3002 42006 3026
rect 42942 3060 43024 3084
rect 42942 3026 42966 3060
rect 43000 3026 43024 3060
rect 42942 3002 43024 3026
rect 43960 3060 44042 3084
rect 43960 3026 43984 3060
rect 44018 3026 44042 3060
rect 43960 3002 44042 3026
rect 44978 3060 45060 3084
rect 44978 3026 45002 3060
rect 45036 3026 45060 3060
rect 44978 3002 45060 3026
rect 45996 3060 46078 3084
rect 45996 3026 46020 3060
rect 46054 3026 46078 3060
rect 45996 3002 46078 3026
rect 47014 3060 47096 3084
rect 47014 3026 47038 3060
rect 47072 3026 47096 3060
rect 47014 3002 47096 3026
rect 48032 3060 48114 3084
rect 48032 3026 48056 3060
rect 48090 3026 48114 3060
rect 48032 3002 48114 3026
rect 49050 3060 49132 3084
rect 49050 3026 49074 3060
rect 49108 3026 49132 3060
rect 49050 3002 49132 3026
rect 50068 3060 50150 3084
rect 50068 3026 50092 3060
rect 50126 3026 50150 3060
rect 50068 3002 50150 3026
rect 51086 3060 51168 3084
rect 51086 3026 51110 3060
rect 51144 3026 51168 3060
rect 51086 3002 51168 3026
rect 52104 3060 52186 3084
rect 52104 3026 52128 3060
rect 52162 3026 52186 3060
rect 52104 3002 52186 3026
rect 54530 2902 54564 2918
rect 55548 3494 55582 3510
rect 55548 2902 55582 2918
rect 56566 3494 56600 3510
rect 56566 2902 56600 2918
rect 57584 3494 57618 3510
rect 57584 2902 57618 2918
rect 58602 3494 58636 3510
rect 58602 2902 58636 2918
rect 59620 3494 59654 3510
rect 59620 2902 59654 2918
rect 60638 3494 60672 3510
rect 60638 2902 60672 2918
rect 61656 3494 61690 3510
rect 61656 2902 61690 2918
rect 62674 3494 62708 3510
rect 62674 2902 62708 2918
rect 63692 3494 63726 3510
rect 63692 2902 63726 2918
rect 64710 3494 64744 3510
rect 64710 2902 64744 2918
rect 65728 3494 65762 3510
rect 65728 2902 65762 2918
rect 66746 3494 66780 3510
rect 66746 2902 66780 2918
rect 67764 3494 67798 3510
rect 67764 2902 67798 2918
rect 68782 3494 68816 3510
rect 68782 2902 68816 2918
rect 69800 3494 69834 3510
rect 69800 2902 69834 2918
rect 70818 3494 70852 3510
rect 70818 2902 70852 2918
rect 71836 3494 71870 3510
rect 71836 2902 71870 2918
rect 72854 3494 72888 3510
rect 72854 2902 72888 2918
rect 73872 3494 73906 3510
rect 73872 2902 73906 2918
rect 74890 3494 74924 3510
rect 74890 2902 74924 2918
rect 62156 2868 62216 2878
rect 41674 2810 41690 2844
rect 42246 2810 42262 2844
rect 42692 2810 42708 2844
rect 43264 2810 43280 2844
rect 43710 2810 43726 2844
rect 44282 2810 44298 2844
rect 44728 2810 44744 2844
rect 45300 2810 45316 2844
rect 45746 2810 45762 2844
rect 46318 2810 46334 2844
rect 46764 2810 46780 2844
rect 47336 2810 47352 2844
rect 47782 2810 47798 2844
rect 48354 2810 48370 2844
rect 48800 2810 48816 2844
rect 49372 2810 49388 2844
rect 49818 2810 49834 2844
rect 50390 2810 50406 2844
rect 50836 2810 50852 2844
rect 51408 2810 51424 2844
rect 51854 2810 51870 2844
rect 52426 2810 52442 2844
rect 54762 2834 54778 2868
rect 55334 2834 55350 2868
rect 55780 2834 55796 2868
rect 56352 2834 56368 2868
rect 56798 2834 56814 2868
rect 57370 2834 57386 2868
rect 57816 2834 57832 2868
rect 58388 2834 58404 2868
rect 58834 2834 58850 2868
rect 59406 2834 59422 2868
rect 59852 2834 59868 2868
rect 60424 2834 60440 2868
rect 60870 2834 60886 2868
rect 61442 2834 61458 2868
rect 61888 2834 61904 2868
rect 62460 2834 62476 2868
rect 62906 2834 62922 2868
rect 63478 2834 63494 2868
rect 63924 2834 63940 2868
rect 64496 2834 64512 2868
rect 64942 2834 64958 2868
rect 65514 2834 65530 2868
rect 65960 2834 65976 2868
rect 66532 2834 66548 2868
rect 66978 2834 66994 2868
rect 67550 2834 67566 2868
rect 67996 2834 68012 2868
rect 68568 2834 68584 2868
rect 69014 2834 69030 2868
rect 69586 2834 69602 2868
rect 70032 2834 70048 2868
rect 70604 2834 70620 2868
rect 71050 2834 71066 2868
rect 71622 2834 71638 2868
rect 72068 2834 72084 2868
rect 72640 2834 72656 2868
rect 73086 2834 73102 2868
rect 73658 2834 73674 2868
rect 74104 2834 74120 2868
rect 74676 2834 74692 2868
rect 41442 2760 41476 2776
rect 41442 2168 41476 2184
rect 42460 2760 42494 2776
rect 42460 2168 42494 2184
rect 43478 2760 43512 2776
rect 43478 2168 43512 2184
rect 44496 2760 44530 2776
rect 44496 2168 44530 2184
rect 45514 2760 45548 2776
rect 45514 2168 45548 2184
rect 46532 2760 46566 2776
rect 46532 2168 46566 2184
rect 47550 2760 47584 2776
rect 47550 2168 47584 2184
rect 48568 2760 48602 2776
rect 48568 2168 48602 2184
rect 49586 2760 49620 2776
rect 49586 2168 49620 2184
rect 50604 2760 50638 2776
rect 50604 2168 50638 2184
rect 51622 2760 51656 2776
rect 51622 2168 51656 2184
rect 52640 2760 52674 2776
rect 55024 2614 55106 2638
rect 55024 2580 55048 2614
rect 55082 2580 55106 2614
rect 55024 2556 55106 2580
rect 56042 2614 56124 2638
rect 56042 2580 56066 2614
rect 56100 2580 56124 2614
rect 56042 2556 56124 2580
rect 57060 2614 57142 2638
rect 57060 2580 57084 2614
rect 57118 2580 57142 2614
rect 57060 2556 57142 2580
rect 58078 2614 58160 2638
rect 58078 2580 58102 2614
rect 58136 2580 58160 2614
rect 58078 2556 58160 2580
rect 59096 2614 59178 2638
rect 59096 2580 59120 2614
rect 59154 2580 59178 2614
rect 59096 2556 59178 2580
rect 60114 2614 60196 2638
rect 60114 2580 60138 2614
rect 60172 2580 60196 2614
rect 60114 2556 60196 2580
rect 61132 2614 61214 2638
rect 61132 2580 61156 2614
rect 61190 2580 61214 2614
rect 61132 2556 61214 2580
rect 62150 2614 62232 2638
rect 62150 2580 62174 2614
rect 62208 2580 62232 2614
rect 62150 2556 62232 2580
rect 63168 2614 63250 2638
rect 63168 2580 63192 2614
rect 63226 2580 63250 2614
rect 63168 2556 63250 2580
rect 64186 2614 64268 2638
rect 64186 2580 64210 2614
rect 64244 2580 64268 2614
rect 64186 2556 64268 2580
rect 65204 2614 65286 2638
rect 65204 2580 65228 2614
rect 65262 2580 65286 2614
rect 65204 2556 65286 2580
rect 66222 2614 66304 2638
rect 66222 2580 66246 2614
rect 66280 2580 66304 2614
rect 66222 2556 66304 2580
rect 67240 2614 67322 2638
rect 67240 2580 67264 2614
rect 67298 2580 67322 2614
rect 67240 2556 67322 2580
rect 68258 2614 68340 2638
rect 68258 2580 68282 2614
rect 68316 2580 68340 2614
rect 68258 2556 68340 2580
rect 69276 2614 69358 2638
rect 69276 2580 69300 2614
rect 69334 2580 69358 2614
rect 69276 2556 69358 2580
rect 70294 2614 70376 2638
rect 70294 2580 70318 2614
rect 70352 2580 70376 2614
rect 70294 2556 70376 2580
rect 71312 2614 71394 2638
rect 71312 2580 71336 2614
rect 71370 2580 71394 2614
rect 71312 2556 71394 2580
rect 72330 2614 72412 2638
rect 72330 2580 72354 2614
rect 72388 2580 72412 2614
rect 72330 2556 72412 2580
rect 73348 2614 73430 2638
rect 73348 2580 73372 2614
rect 73406 2580 73430 2614
rect 73348 2556 73430 2580
rect 74366 2614 74448 2638
rect 74366 2580 74390 2614
rect 74424 2580 74448 2614
rect 74366 2556 74448 2580
rect 54762 2310 54778 2344
rect 55334 2310 55350 2344
rect 55780 2310 55796 2344
rect 56352 2310 56368 2344
rect 56798 2310 56814 2344
rect 57370 2310 57386 2344
rect 57816 2310 57832 2344
rect 58388 2310 58404 2344
rect 58834 2310 58850 2344
rect 59406 2310 59422 2344
rect 59852 2310 59868 2344
rect 60424 2310 60440 2344
rect 60870 2310 60886 2344
rect 61442 2310 61458 2344
rect 61888 2310 61904 2344
rect 62460 2310 62476 2344
rect 62906 2310 62922 2344
rect 63478 2310 63494 2344
rect 63924 2310 63940 2344
rect 64496 2310 64512 2344
rect 64942 2310 64958 2344
rect 65514 2310 65530 2344
rect 65960 2310 65976 2344
rect 66532 2310 66548 2344
rect 66978 2310 66994 2344
rect 67550 2310 67566 2344
rect 67996 2310 68012 2344
rect 68568 2310 68584 2344
rect 69014 2310 69030 2344
rect 69586 2310 69602 2344
rect 70032 2310 70048 2344
rect 70604 2310 70620 2344
rect 71050 2310 71066 2344
rect 71622 2310 71638 2344
rect 72068 2310 72084 2344
rect 72640 2310 72656 2344
rect 73086 2310 73102 2344
rect 73658 2310 73674 2344
rect 74104 2310 74120 2344
rect 74676 2310 74692 2344
rect 58070 2308 58130 2310
rect 52640 2168 52674 2184
rect 54530 2260 54564 2276
rect 41674 2100 41690 2134
rect 42246 2100 42262 2134
rect 42692 2100 42708 2134
rect 43264 2100 43280 2134
rect 43710 2100 43726 2134
rect 44282 2100 44298 2134
rect 44728 2100 44744 2134
rect 45300 2100 45316 2134
rect 45746 2100 45762 2134
rect 46318 2100 46334 2134
rect 46764 2100 46780 2134
rect 47336 2100 47352 2134
rect 47782 2100 47798 2134
rect 48354 2100 48370 2134
rect 48800 2100 48816 2134
rect 49372 2100 49388 2134
rect 49818 2100 49834 2134
rect 50390 2100 50406 2134
rect 50836 2100 50852 2134
rect 51408 2100 51424 2134
rect 51854 2100 51870 2134
rect 52426 2100 52442 2134
rect 41924 1718 42006 1742
rect 41924 1684 41948 1718
rect 41982 1684 42006 1718
rect 41924 1660 42006 1684
rect 42942 1718 43024 1742
rect 42942 1684 42966 1718
rect 43000 1684 43024 1718
rect 42942 1660 43024 1684
rect 43960 1718 44042 1742
rect 43960 1684 43984 1718
rect 44018 1684 44042 1718
rect 43960 1660 44042 1684
rect 44978 1718 45060 1742
rect 44978 1684 45002 1718
rect 45036 1684 45060 1718
rect 44978 1660 45060 1684
rect 45996 1718 46078 1742
rect 45996 1684 46020 1718
rect 46054 1684 46078 1718
rect 45996 1660 46078 1684
rect 47014 1718 47096 1742
rect 47014 1684 47038 1718
rect 47072 1684 47096 1718
rect 47014 1660 47096 1684
rect 48032 1718 48114 1742
rect 48032 1684 48056 1718
rect 48090 1684 48114 1718
rect 48032 1660 48114 1684
rect 49050 1718 49132 1742
rect 49050 1684 49074 1718
rect 49108 1684 49132 1718
rect 49050 1660 49132 1684
rect 50068 1718 50150 1742
rect 50068 1684 50092 1718
rect 50126 1684 50150 1718
rect 50068 1660 50150 1684
rect 51086 1718 51168 1742
rect 51086 1684 51110 1718
rect 51144 1684 51168 1718
rect 51086 1660 51168 1684
rect 52104 1718 52186 1742
rect 52104 1684 52128 1718
rect 52162 1684 52186 1718
rect 52104 1660 52186 1684
rect 54530 1668 54564 1684
rect 55548 2260 55582 2276
rect 55548 1668 55582 1684
rect 56566 2260 56600 2276
rect 56566 1668 56600 1684
rect 57584 2260 57618 2276
rect 57584 1668 57618 1684
rect 58602 2260 58636 2276
rect 58602 1668 58636 1684
rect 59620 2260 59654 2276
rect 59620 1668 59654 1684
rect 60638 2260 60672 2276
rect 60638 1668 60672 1684
rect 61656 2260 61690 2276
rect 61656 1668 61690 1684
rect 62674 2260 62708 2276
rect 62674 1668 62708 1684
rect 63692 2260 63726 2276
rect 63692 1668 63726 1684
rect 64710 2260 64744 2276
rect 64710 1668 64744 1684
rect 65728 2260 65762 2276
rect 65728 1668 65762 1684
rect 66746 2260 66780 2276
rect 66746 1668 66780 1684
rect 67764 2260 67798 2276
rect 67764 1668 67798 1684
rect 68782 2260 68816 2276
rect 68782 1668 68816 1684
rect 69800 2260 69834 2276
rect 69800 1668 69834 1684
rect 70818 2260 70852 2276
rect 70818 1668 70852 1684
rect 71836 2260 71870 2276
rect 71836 1668 71870 1684
rect 72854 2260 72888 2276
rect 72854 1668 72888 1684
rect 73872 2260 73906 2276
rect 73872 1668 73906 1684
rect 74890 2260 74924 2276
rect 74890 1668 74924 1684
rect 56038 1634 56098 1636
rect 62150 1634 62210 1636
rect 64184 1634 64244 1636
rect 68250 1634 68310 1640
rect 72326 1634 72386 1636
rect 73342 1634 73402 1636
rect 54762 1600 54778 1634
rect 55334 1600 55350 1634
rect 55780 1600 55796 1634
rect 56352 1600 56368 1634
rect 56798 1600 56814 1634
rect 57370 1600 57386 1634
rect 57816 1600 57832 1634
rect 58388 1600 58404 1634
rect 58834 1600 58850 1634
rect 59406 1600 59422 1634
rect 59852 1600 59868 1634
rect 60424 1600 60440 1634
rect 60870 1600 60886 1634
rect 61442 1600 61458 1634
rect 61888 1600 61904 1634
rect 62460 1600 62476 1634
rect 62906 1600 62922 1634
rect 63478 1600 63494 1634
rect 63924 1600 63940 1634
rect 64496 1600 64512 1634
rect 64942 1600 64958 1634
rect 65514 1600 65530 1634
rect 65960 1600 65976 1634
rect 66532 1600 66548 1634
rect 66978 1600 66994 1634
rect 67550 1600 67566 1634
rect 67996 1600 68012 1634
rect 68568 1600 68584 1634
rect 69014 1600 69030 1634
rect 69586 1600 69602 1634
rect 70032 1600 70048 1634
rect 70604 1600 70620 1634
rect 71050 1600 71066 1634
rect 71622 1600 71638 1634
rect 72068 1600 72084 1634
rect 72640 1600 72656 1634
rect 73086 1600 73102 1634
rect 73658 1600 73674 1634
rect 74104 1600 74120 1634
rect 74676 1600 74692 1634
rect 55036 1368 55118 1392
rect 55036 1334 55060 1368
rect 55094 1334 55118 1368
rect 55036 1310 55118 1334
rect 56054 1368 56136 1392
rect 56054 1334 56078 1368
rect 56112 1334 56136 1368
rect 56054 1310 56136 1334
rect 57072 1368 57154 1392
rect 57072 1334 57096 1368
rect 57130 1334 57154 1368
rect 57072 1310 57154 1334
rect 58090 1368 58172 1392
rect 58090 1334 58114 1368
rect 58148 1334 58172 1368
rect 58090 1310 58172 1334
rect 59108 1368 59190 1392
rect 59108 1334 59132 1368
rect 59166 1334 59190 1368
rect 59108 1310 59190 1334
rect 60126 1368 60208 1392
rect 60126 1334 60150 1368
rect 60184 1334 60208 1368
rect 60126 1310 60208 1334
rect 61144 1368 61226 1392
rect 61144 1334 61168 1368
rect 61202 1334 61226 1368
rect 61144 1310 61226 1334
rect 62162 1368 62244 1392
rect 62162 1334 62186 1368
rect 62220 1334 62244 1368
rect 62162 1310 62244 1334
rect 63180 1368 63262 1392
rect 63180 1334 63204 1368
rect 63238 1334 63262 1368
rect 63180 1310 63262 1334
rect 64198 1368 64280 1392
rect 64198 1334 64222 1368
rect 64256 1334 64280 1368
rect 64198 1310 64280 1334
rect 65216 1368 65298 1392
rect 65216 1334 65240 1368
rect 65274 1334 65298 1368
rect 65216 1310 65298 1334
rect 66234 1368 66316 1392
rect 66234 1334 66258 1368
rect 66292 1334 66316 1368
rect 66234 1310 66316 1334
rect 67252 1368 67334 1392
rect 67252 1334 67276 1368
rect 67310 1334 67334 1368
rect 67252 1310 67334 1334
rect 68270 1368 68352 1392
rect 68270 1334 68294 1368
rect 68328 1334 68352 1368
rect 68270 1310 68352 1334
rect 69288 1368 69370 1392
rect 69288 1334 69312 1368
rect 69346 1334 69370 1368
rect 69288 1310 69370 1334
rect 70306 1368 70388 1392
rect 70306 1334 70330 1368
rect 70364 1334 70388 1368
rect 70306 1310 70388 1334
rect 71324 1368 71406 1392
rect 71324 1334 71348 1368
rect 71382 1334 71406 1368
rect 71324 1310 71406 1334
rect 72342 1368 72424 1392
rect 72342 1334 72366 1368
rect 72400 1334 72424 1368
rect 72342 1310 72424 1334
rect 73360 1368 73442 1392
rect 73360 1334 73384 1368
rect 73418 1334 73442 1368
rect 73360 1310 73442 1334
rect 74378 1368 74460 1392
rect 74378 1334 74402 1368
rect 74436 1334 74460 1368
rect 74378 1310 74460 1334
rect 42132 1268 42148 1302
rect 42704 1268 42720 1302
rect 43150 1268 43166 1302
rect 43722 1268 43738 1302
rect 44168 1268 44184 1302
rect 44740 1268 44756 1302
rect 45186 1268 45202 1302
rect 45758 1268 45774 1302
rect 46204 1268 46220 1302
rect 46776 1268 46792 1302
rect 47222 1268 47238 1302
rect 47794 1268 47810 1302
rect 48240 1268 48256 1302
rect 48812 1268 48828 1302
rect 49258 1268 49274 1302
rect 49830 1268 49846 1302
rect 50276 1268 50292 1302
rect 50848 1268 50864 1302
rect 51294 1268 51310 1302
rect 51866 1268 51882 1302
rect 41900 1218 41934 1234
rect 41900 626 41934 642
rect 42918 1218 42952 1234
rect 42918 626 42952 642
rect 43936 1218 43970 1234
rect 43936 626 43970 642
rect 44954 1218 44988 1234
rect 44954 626 44988 642
rect 45972 1218 46006 1234
rect 45972 626 46006 642
rect 46990 1218 47024 1234
rect 46990 626 47024 642
rect 48008 1218 48042 1234
rect 48008 626 48042 642
rect 49026 1218 49060 1234
rect 49026 626 49060 642
rect 50044 1218 50078 1234
rect 50044 626 50078 642
rect 51062 1218 51096 1234
rect 51062 626 51096 642
rect 52080 1218 52114 1234
rect 54762 1078 54778 1112
rect 55334 1078 55350 1112
rect 55780 1078 55796 1112
rect 56352 1078 56368 1112
rect 56798 1078 56814 1112
rect 57370 1078 57386 1112
rect 57816 1078 57832 1112
rect 58388 1078 58404 1112
rect 58834 1078 58850 1112
rect 59406 1078 59422 1112
rect 59852 1078 59868 1112
rect 60424 1078 60440 1112
rect 60870 1078 60886 1112
rect 61442 1078 61458 1112
rect 61888 1078 61904 1112
rect 62460 1078 62476 1112
rect 62906 1078 62922 1112
rect 63478 1078 63494 1112
rect 63924 1078 63940 1112
rect 64496 1078 64512 1112
rect 64942 1078 64958 1112
rect 65514 1078 65530 1112
rect 65960 1078 65976 1112
rect 66532 1078 66548 1112
rect 66978 1078 66994 1112
rect 67550 1078 67566 1112
rect 67996 1078 68012 1112
rect 68568 1078 68584 1112
rect 69014 1078 69030 1112
rect 69586 1078 69602 1112
rect 70032 1078 70048 1112
rect 70604 1078 70620 1112
rect 71050 1078 71066 1112
rect 71622 1078 71638 1112
rect 72068 1078 72084 1112
rect 72640 1078 72656 1112
rect 73086 1078 73102 1112
rect 73658 1078 73674 1112
rect 74104 1078 74120 1112
rect 74676 1078 74692 1112
rect 52080 626 52114 642
rect 54530 1028 54564 1044
rect 42132 558 42148 592
rect 42704 558 42720 592
rect 43150 558 43166 592
rect 43722 558 43738 592
rect 44168 558 44184 592
rect 44740 558 44756 592
rect 45186 558 45202 592
rect 45758 558 45774 592
rect 46204 558 46220 592
rect 46776 558 46792 592
rect 47222 558 47238 592
rect 47794 558 47810 592
rect 48240 558 48256 592
rect 48812 558 48828 592
rect 49258 558 49274 592
rect 49830 558 49846 592
rect 50276 558 50292 592
rect 50848 558 50864 592
rect 51294 558 51310 592
rect 51866 558 51882 592
rect 54530 436 54564 452
rect 55548 1028 55582 1044
rect 55548 436 55582 452
rect 56566 1028 56600 1044
rect 56566 436 56600 452
rect 57584 1028 57618 1044
rect 57584 436 57618 452
rect 58602 1028 58636 1044
rect 58602 436 58636 452
rect 59620 1028 59654 1044
rect 59620 436 59654 452
rect 60638 1028 60672 1044
rect 60638 436 60672 452
rect 61656 1028 61690 1044
rect 61656 436 61690 452
rect 62674 1028 62708 1044
rect 62674 436 62708 452
rect 63692 1028 63726 1044
rect 63692 436 63726 452
rect 64710 1028 64744 1044
rect 64710 436 64744 452
rect 65728 1028 65762 1044
rect 65728 436 65762 452
rect 66746 1028 66780 1044
rect 66746 436 66780 452
rect 67764 1028 67798 1044
rect 67764 436 67798 452
rect 68782 1028 68816 1044
rect 68782 436 68816 452
rect 69800 1028 69834 1044
rect 69800 436 69834 452
rect 70818 1028 70852 1044
rect 70818 436 70852 452
rect 71836 1028 71870 1044
rect 71836 436 71870 452
rect 72854 1028 72888 1044
rect 72854 436 72888 452
rect 73872 1028 73906 1044
rect 73872 436 73906 452
rect 74890 1028 74924 1044
rect 74890 436 74924 452
rect 54762 368 54778 402
rect 55334 368 55350 402
rect 55780 368 55796 402
rect 56352 368 56368 402
rect 56798 368 56814 402
rect 57370 368 57386 402
rect 57816 368 57832 402
rect 58388 368 58404 402
rect 58834 368 58850 402
rect 59406 368 59422 402
rect 59852 368 59868 402
rect 60424 368 60440 402
rect 60870 368 60886 402
rect 61442 368 61458 402
rect 61888 368 61904 402
rect 62460 368 62476 402
rect 62906 368 62922 402
rect 63478 368 63494 402
rect 63924 368 63940 402
rect 64496 368 64512 402
rect 64942 368 64958 402
rect 65514 368 65530 402
rect 65960 368 65976 402
rect 66532 368 66548 402
rect 66978 368 66994 402
rect 67550 368 67566 402
rect 67996 368 68012 402
rect 68568 368 68584 402
rect 69014 368 69030 402
rect 69586 368 69602 402
rect 70032 368 70048 402
rect 70604 368 70620 402
rect 71050 368 71066 402
rect 71622 368 71638 402
rect 72068 368 72084 402
rect 72640 368 72656 402
rect 73086 368 73102 402
rect 73658 368 73674 402
rect 74104 368 74120 402
rect 74676 368 74692 402
rect 41734 272 41816 296
rect 41734 238 41758 272
rect 41792 238 41816 272
rect 41734 214 41816 238
rect 42752 272 42834 296
rect 42752 238 42776 272
rect 42810 238 42834 272
rect 42752 214 42834 238
rect 43770 272 43852 296
rect 43770 238 43794 272
rect 43828 238 43852 272
rect 43770 214 43852 238
rect 44788 272 44870 296
rect 44788 238 44812 272
rect 44846 238 44870 272
rect 44788 214 44870 238
rect 45806 272 45888 296
rect 45806 238 45830 272
rect 45864 238 45888 272
rect 45806 214 45888 238
rect 46824 272 46906 296
rect 46824 238 46848 272
rect 46882 238 46906 272
rect 46824 214 46906 238
rect 47842 272 47924 296
rect 47842 238 47866 272
rect 47900 238 47924 272
rect 47842 214 47924 238
rect 48860 272 48942 296
rect 48860 238 48884 272
rect 48918 238 48942 272
rect 48860 214 48942 238
rect 49878 272 49960 296
rect 49878 238 49902 272
rect 49936 238 49960 272
rect 49878 214 49960 238
rect 50896 272 50978 296
rect 50896 238 50920 272
rect 50954 238 50978 272
rect 50896 214 50978 238
rect 51914 272 51996 296
rect 51914 238 51938 272
rect 51972 238 51996 272
rect 51914 214 51996 238
rect 55024 190 55106 214
rect 55024 156 55048 190
rect 55082 156 55106 190
rect 55024 132 55106 156
rect 56042 190 56124 214
rect 56042 156 56066 190
rect 56100 156 56124 190
rect 56042 132 56124 156
rect 57060 190 57142 214
rect 57060 156 57084 190
rect 57118 156 57142 190
rect 57060 132 57142 156
rect 58078 190 58160 214
rect 58078 156 58102 190
rect 58136 156 58160 190
rect 58078 132 58160 156
rect 59096 190 59178 214
rect 59096 156 59120 190
rect 59154 156 59178 190
rect 59096 132 59178 156
rect 60114 190 60196 214
rect 60114 156 60138 190
rect 60172 156 60196 190
rect 60114 132 60196 156
rect 61132 190 61214 214
rect 61132 156 61156 190
rect 61190 156 61214 190
rect 61132 132 61214 156
rect 62150 190 62232 214
rect 62150 156 62174 190
rect 62208 156 62232 190
rect 62150 132 62232 156
rect 63168 190 63250 214
rect 63168 156 63192 190
rect 63226 156 63250 190
rect 63168 132 63250 156
rect 64186 190 64268 214
rect 64186 156 64210 190
rect 64244 156 64268 190
rect 64186 132 64268 156
rect 65204 190 65286 214
rect 65204 156 65228 190
rect 65262 156 65286 190
rect 65204 132 65286 156
rect 66222 190 66304 214
rect 66222 156 66246 190
rect 66280 156 66304 190
rect 66222 132 66304 156
rect 67240 190 67322 214
rect 67240 156 67264 190
rect 67298 156 67322 190
rect 67240 132 67322 156
rect 68258 190 68340 214
rect 68258 156 68282 190
rect 68316 156 68340 190
rect 68258 132 68340 156
rect 69276 190 69358 214
rect 69276 156 69300 190
rect 69334 156 69358 190
rect 69276 132 69358 156
rect 70294 190 70376 214
rect 70294 156 70318 190
rect 70352 156 70376 190
rect 70294 132 70376 156
rect 71312 190 71394 214
rect 71312 156 71336 190
rect 71370 156 71394 190
rect 71312 132 71394 156
rect 72330 190 72412 214
rect 72330 156 72354 190
rect 72388 156 72412 190
rect 72330 132 72412 156
rect 73348 190 73430 214
rect 73348 156 73372 190
rect 73406 156 73430 190
rect 73348 132 73430 156
rect 74366 190 74448 214
rect 74366 156 74390 190
rect 74424 156 74448 190
rect 74366 132 74448 156
rect 39628 -852 39728 -690
rect 76772 -852 76872 -690
<< viali >>
rect 11428 30592 11490 30692
rect 11490 30592 35610 30692
rect 35610 30592 35672 30692
rect 11328 16642 11428 30072
rect 17732 27891 18196 27925
rect 18750 27891 19214 27925
rect 19768 27891 20232 27925
rect 20786 27891 21250 27925
rect 21804 27891 22268 27925
rect 22822 27891 23286 27925
rect 23840 27891 24304 27925
rect 24858 27891 25322 27925
rect 25876 27891 26340 27925
rect 26894 27891 27358 27925
rect 27912 27891 28376 27925
rect 28930 27891 29394 27925
rect 29948 27891 30412 27925
rect 30966 27891 31430 27925
rect 31984 27891 32448 27925
rect 33002 27891 33466 27925
rect 17438 27256 17472 27832
rect 18456 27256 18490 27832
rect 19474 27256 19508 27832
rect 20492 27256 20526 27832
rect 21510 27256 21544 27832
rect 22528 27256 22562 27832
rect 23546 27256 23580 27832
rect 24564 27256 24598 27832
rect 25582 27256 25616 27832
rect 26600 27256 26634 27832
rect 27618 27256 27652 27832
rect 28636 27256 28670 27832
rect 29654 27256 29688 27832
rect 30672 27256 30706 27832
rect 31690 27256 31724 27832
rect 32708 27256 32742 27832
rect 33726 27256 33760 27832
rect 17732 27163 18196 27197
rect 18750 27163 19214 27197
rect 19768 27163 20232 27197
rect 20786 27163 21250 27197
rect 21804 27163 22268 27197
rect 22822 27163 23286 27197
rect 23840 27163 24304 27197
rect 24858 27163 25322 27197
rect 25876 27163 26340 27197
rect 26894 27163 27358 27197
rect 27912 27163 28376 27197
rect 28930 27163 29394 27197
rect 29948 27163 30412 27197
rect 30966 27163 31430 27197
rect 31984 27163 32448 27197
rect 33002 27163 33466 27197
rect 17732 26755 18196 26789
rect 18750 26755 19214 26789
rect 19768 26755 20232 26789
rect 20786 26755 21250 26789
rect 21804 26755 22268 26789
rect 22822 26755 23286 26789
rect 23840 26755 24304 26789
rect 24858 26755 25322 26789
rect 25876 26755 26340 26789
rect 26894 26755 27358 26789
rect 27912 26755 28376 26789
rect 28930 26755 29394 26789
rect 29948 26755 30412 26789
rect 30966 26755 31430 26789
rect 31984 26755 32448 26789
rect 33002 26755 33466 26789
rect 17438 26120 17472 26696
rect 18456 26120 18490 26696
rect 19474 26120 19508 26696
rect 20492 26120 20526 26696
rect 21510 26120 21544 26696
rect 22528 26120 22562 26696
rect 23546 26120 23580 26696
rect 24564 26120 24598 26696
rect 25582 26120 25616 26696
rect 26600 26120 26634 26696
rect 27618 26120 27652 26696
rect 28636 26120 28670 26696
rect 29654 26120 29688 26696
rect 30672 26120 30706 26696
rect 31690 26120 31724 26696
rect 32708 26120 32742 26696
rect 33726 26120 33760 26696
rect 17732 26027 18196 26061
rect 18750 26027 19214 26061
rect 19768 26027 20232 26061
rect 20786 26027 21250 26061
rect 21804 26027 22268 26061
rect 22822 26027 23286 26061
rect 23840 26027 24304 26061
rect 24858 26027 25322 26061
rect 25876 26027 26340 26061
rect 26894 26027 27358 26061
rect 27912 26027 28376 26061
rect 28930 26027 29394 26061
rect 29948 26027 30412 26061
rect 30966 26027 31430 26061
rect 31984 26027 32448 26061
rect 33002 26027 33466 26061
rect 17732 25619 18196 25653
rect 18750 25619 19214 25653
rect 19768 25619 20232 25653
rect 20786 25619 21250 25653
rect 21804 25619 22268 25653
rect 22822 25619 23286 25653
rect 23840 25619 24304 25653
rect 24858 25619 25322 25653
rect 25876 25619 26340 25653
rect 26894 25619 27358 25653
rect 27912 25619 28376 25653
rect 28930 25619 29394 25653
rect 29948 25619 30412 25653
rect 30966 25619 31430 25653
rect 31984 25619 32448 25653
rect 33002 25619 33466 25653
rect 17438 24984 17472 25560
rect 18456 24984 18490 25560
rect 19474 24984 19508 25560
rect 20492 24984 20526 25560
rect 21510 24984 21544 25560
rect 22528 24984 22562 25560
rect 23546 24984 23580 25560
rect 24564 24984 24598 25560
rect 25582 24984 25616 25560
rect 26600 24984 26634 25560
rect 27618 24984 27652 25560
rect 28636 24984 28670 25560
rect 29654 24984 29688 25560
rect 30672 24984 30706 25560
rect 31690 24984 31724 25560
rect 32708 24984 32742 25560
rect 33726 24984 33760 25560
rect 17732 24891 18196 24925
rect 18750 24891 19214 24925
rect 19768 24891 20232 24925
rect 20786 24891 21250 24925
rect 21804 24891 22268 24925
rect 22822 24891 23286 24925
rect 23840 24891 24304 24925
rect 24858 24891 25322 24925
rect 25876 24891 26340 24925
rect 26894 24891 27358 24925
rect 27912 24891 28376 24925
rect 28930 24891 29394 24925
rect 29948 24891 30412 24925
rect 30966 24891 31430 24925
rect 31984 24891 32448 24925
rect 33002 24891 33466 24925
rect 18926 23981 19390 24015
rect 19944 23981 20408 24015
rect 20962 23981 21426 24015
rect 21980 23981 22444 24015
rect 22998 23981 23462 24015
rect 24016 23981 24480 24015
rect 25034 23981 25498 24015
rect 26052 23981 26516 24015
rect 27070 23981 27534 24015
rect 28088 23981 28552 24015
rect 29106 23981 29570 24015
rect 30124 23981 30588 24015
rect 31142 23981 31606 24015
rect 32160 23981 32624 24015
rect 18632 23346 18666 23922
rect 19650 23346 19684 23922
rect 20668 23346 20702 23922
rect 21686 23346 21720 23922
rect 22704 23346 22738 23922
rect 23722 23346 23756 23922
rect 24740 23346 24774 23922
rect 25758 23346 25792 23922
rect 26776 23346 26810 23922
rect 27794 23346 27828 23922
rect 28812 23346 28846 23922
rect 29830 23346 29864 23922
rect 30848 23346 30882 23922
rect 31866 23346 31900 23922
rect 32884 23346 32918 23922
rect 18926 23253 19390 23287
rect 19944 23253 20408 23287
rect 20962 23253 21426 23287
rect 21980 23253 22444 23287
rect 22998 23253 23462 23287
rect 24016 23253 24480 23287
rect 25034 23253 25498 23287
rect 26052 23253 26516 23287
rect 27070 23253 27534 23287
rect 28088 23253 28552 23287
rect 29106 23253 29570 23287
rect 30124 23253 30588 23287
rect 31142 23253 31606 23287
rect 32160 23253 32624 23287
rect 18926 22949 19390 22983
rect 19944 22949 20408 22983
rect 20962 22949 21426 22983
rect 21980 22949 22444 22983
rect 22998 22949 23462 22983
rect 24016 22949 24480 22983
rect 25034 22949 25498 22983
rect 26052 22949 26516 22983
rect 27070 22949 27534 22983
rect 28088 22949 28552 22983
rect 29106 22949 29570 22983
rect 30124 22949 30588 22983
rect 31142 22949 31606 22983
rect 32160 22949 32624 22983
rect 18632 22314 18666 22890
rect 19650 22314 19684 22890
rect 20668 22314 20702 22890
rect 21686 22314 21720 22890
rect 22704 22314 22738 22890
rect 23722 22314 23756 22890
rect 24740 22314 24774 22890
rect 25758 22314 25792 22890
rect 26776 22314 26810 22890
rect 27794 22314 27828 22890
rect 28812 22314 28846 22890
rect 29830 22314 29864 22890
rect 30848 22314 30882 22890
rect 31866 22314 31900 22890
rect 32884 22314 32918 22890
rect 18926 22221 19390 22255
rect 19944 22221 20408 22255
rect 20962 22221 21426 22255
rect 21980 22221 22444 22255
rect 22998 22221 23462 22255
rect 24016 22221 24480 22255
rect 25034 22221 25498 22255
rect 26052 22221 26516 22255
rect 27070 22221 27534 22255
rect 28088 22221 28552 22255
rect 29106 22221 29570 22255
rect 30124 22221 30588 22255
rect 31142 22221 31606 22255
rect 32160 22221 32624 22255
rect 18718 21345 19182 21379
rect 19736 21345 20200 21379
rect 20754 21345 21218 21379
rect 21772 21345 22236 21379
rect 22790 21345 23254 21379
rect 23808 21345 24272 21379
rect 24826 21345 25290 21379
rect 25844 21345 26308 21379
rect 26862 21345 27326 21379
rect 27880 21345 28344 21379
rect 28898 21345 29362 21379
rect 29916 21345 30380 21379
rect 30934 21345 31398 21379
rect 31952 21345 32416 21379
rect 32970 21345 33434 21379
rect 13414 21241 13878 21275
rect 14432 21241 14896 21275
rect 15450 21241 15914 21275
rect 16468 21241 16932 21275
rect 13120 20606 13154 21182
rect 14138 20606 14172 21182
rect 15156 20606 15190 21182
rect 16174 20606 16208 21182
rect 17192 20606 17226 21182
rect 18424 20710 18458 21286
rect 19442 20710 19476 21286
rect 20460 20710 20494 21286
rect 21478 20710 21512 21286
rect 22496 20710 22530 21286
rect 23514 20710 23548 21286
rect 24532 20710 24566 21286
rect 25550 20710 25584 21286
rect 26568 20710 26602 21286
rect 27586 20710 27620 21286
rect 28604 20710 28638 21286
rect 29622 20710 29656 21286
rect 30640 20710 30674 21286
rect 31658 20710 31692 21286
rect 32676 20710 32710 21286
rect 33694 20710 33728 21286
rect 18718 20617 19182 20651
rect 19736 20617 20200 20651
rect 20754 20617 21218 20651
rect 21772 20617 22236 20651
rect 22790 20617 23254 20651
rect 23808 20617 24272 20651
rect 24826 20617 25290 20651
rect 25844 20617 26308 20651
rect 26862 20617 27326 20651
rect 27880 20617 28344 20651
rect 28898 20617 29362 20651
rect 29916 20617 30380 20651
rect 30934 20617 31398 20651
rect 31952 20617 32416 20651
rect 32970 20617 33434 20651
rect 13414 20513 13878 20547
rect 14432 20513 14896 20547
rect 15450 20513 15914 20547
rect 16468 20513 16932 20547
rect 13414 20209 13878 20243
rect 14432 20209 14896 20243
rect 15450 20209 15914 20243
rect 16468 20209 16932 20243
rect 13120 19574 13154 20150
rect 14138 19574 14172 20150
rect 15156 19574 15190 20150
rect 16174 19574 16208 20150
rect 17192 19574 17226 20150
rect 18718 20089 19182 20123
rect 19736 20089 20200 20123
rect 20754 20089 21218 20123
rect 21772 20089 22236 20123
rect 22790 20089 23254 20123
rect 23808 20089 24272 20123
rect 24826 20089 25290 20123
rect 25844 20089 26308 20123
rect 26862 20089 27326 20123
rect 27880 20089 28344 20123
rect 28898 20089 29362 20123
rect 29916 20089 30380 20123
rect 30934 20089 31398 20123
rect 31952 20089 32416 20123
rect 32970 20089 33434 20123
rect 13414 19481 13878 19515
rect 14432 19481 14896 19515
rect 15450 19481 15914 19515
rect 16468 19481 16932 19515
rect 18424 19454 18458 20030
rect 19442 19454 19476 20030
rect 20460 19454 20494 20030
rect 21478 19454 21512 20030
rect 22496 19454 22530 20030
rect 23514 19454 23548 20030
rect 24532 19454 24566 20030
rect 25550 19454 25584 20030
rect 26568 19454 26602 20030
rect 27586 19454 27620 20030
rect 28604 19454 28638 20030
rect 29622 19454 29656 20030
rect 30640 19454 30674 20030
rect 31658 19454 31692 20030
rect 32676 19454 32710 20030
rect 33694 19454 33728 20030
rect 18718 19361 19182 19395
rect 19736 19361 20200 19395
rect 20754 19361 21218 19395
rect 21772 19361 22236 19395
rect 22790 19361 23254 19395
rect 23808 19361 24272 19395
rect 24826 19361 25290 19395
rect 25844 19361 26308 19395
rect 26862 19361 27326 19395
rect 27880 19361 28344 19395
rect 28898 19361 29362 19395
rect 29916 19361 30380 19395
rect 30934 19361 31398 19395
rect 31952 19361 32416 19395
rect 32970 19361 33434 19395
rect 13414 19177 13878 19211
rect 14432 19177 14896 19211
rect 15450 19177 15914 19211
rect 16468 19177 16932 19211
rect 13120 18542 13154 19118
rect 14138 18542 14172 19118
rect 15156 18542 15190 19118
rect 16174 18542 16208 19118
rect 17192 18542 17226 19118
rect 18718 18833 19182 18867
rect 19736 18833 20200 18867
rect 20754 18833 21218 18867
rect 21772 18833 22236 18867
rect 22790 18833 23254 18867
rect 23808 18833 24272 18867
rect 24826 18833 25290 18867
rect 25844 18833 26308 18867
rect 26862 18833 27326 18867
rect 27880 18833 28344 18867
rect 28898 18833 29362 18867
rect 29916 18833 30380 18867
rect 30934 18833 31398 18867
rect 31952 18833 32416 18867
rect 32970 18833 33434 18867
rect 13414 18449 13878 18483
rect 14432 18449 14896 18483
rect 15450 18449 15914 18483
rect 16468 18449 16932 18483
rect 18424 18198 18458 18774
rect 19442 18198 19476 18774
rect 20460 18198 20494 18774
rect 21478 18198 21512 18774
rect 22496 18198 22530 18774
rect 23514 18198 23548 18774
rect 24532 18198 24566 18774
rect 25550 18198 25584 18774
rect 26568 18198 26602 18774
rect 27586 18198 27620 18774
rect 28604 18198 28638 18774
rect 29622 18198 29656 18774
rect 30640 18198 30674 18774
rect 31658 18198 31692 18774
rect 32676 18198 32710 18774
rect 33694 18198 33728 18774
rect 13414 18145 13878 18179
rect 14432 18145 14896 18179
rect 15450 18145 15914 18179
rect 16468 18145 16932 18179
rect 18718 18105 19182 18139
rect 19736 18105 20200 18139
rect 20754 18105 21218 18139
rect 21772 18105 22236 18139
rect 22790 18105 23254 18139
rect 23808 18105 24272 18139
rect 24826 18105 25290 18139
rect 25844 18105 26308 18139
rect 26862 18105 27326 18139
rect 27880 18105 28344 18139
rect 28898 18105 29362 18139
rect 29916 18105 30380 18139
rect 30934 18105 31398 18139
rect 31952 18105 32416 18139
rect 32970 18105 33434 18139
rect 13120 17510 13154 18086
rect 14138 17510 14172 18086
rect 15156 17510 15190 18086
rect 16174 17510 16208 18086
rect 17192 17510 17226 18086
rect 18718 17577 19182 17611
rect 19736 17577 20200 17611
rect 20754 17577 21218 17611
rect 21772 17577 22236 17611
rect 22790 17577 23254 17611
rect 23808 17577 24272 17611
rect 24826 17577 25290 17611
rect 25844 17577 26308 17611
rect 26862 17577 27326 17611
rect 27880 17577 28344 17611
rect 28898 17577 29362 17611
rect 29916 17577 30380 17611
rect 30934 17577 31398 17611
rect 31952 17577 32416 17611
rect 32970 17577 33434 17611
rect 13414 17417 13878 17451
rect 14432 17417 14896 17451
rect 15450 17417 15914 17451
rect 16468 17417 16932 17451
rect 18424 16942 18458 17518
rect 19442 16942 19476 17518
rect 20460 16942 20494 17518
rect 21478 16942 21512 17518
rect 22496 16942 22530 17518
rect 23514 16942 23548 17518
rect 24532 16942 24566 17518
rect 25550 16942 25584 17518
rect 26568 16942 26602 17518
rect 27586 16942 27620 17518
rect 28604 16942 28638 17518
rect 29622 16942 29656 17518
rect 30640 16942 30674 17518
rect 31658 16942 31692 17518
rect 32676 16942 32710 17518
rect 33694 16942 33728 17518
rect 18718 16849 19182 16883
rect 19736 16849 20200 16883
rect 20754 16849 21218 16883
rect 21772 16849 22236 16883
rect 22790 16849 23254 16883
rect 23808 16849 24272 16883
rect 24826 16849 25290 16883
rect 25844 16849 26308 16883
rect 26862 16849 27326 16883
rect 27880 16849 28344 16883
rect 28898 16849 29362 16883
rect 29916 16849 30380 16883
rect 30934 16849 31398 16883
rect 31952 16849 32416 16883
rect 32970 16849 33434 16883
rect 35672 16642 35772 30072
rect 11428 16022 11490 16122
rect 11490 16022 35610 16122
rect 35610 16022 35672 16122
rect 52428 30592 52490 30692
rect 52490 30592 76610 30692
rect 76610 30592 76672 30692
rect 52328 16642 52428 30072
rect 58732 27891 59196 27925
rect 59750 27891 60214 27925
rect 60768 27891 61232 27925
rect 61786 27891 62250 27925
rect 62804 27891 63268 27925
rect 63822 27891 64286 27925
rect 64840 27891 65304 27925
rect 65858 27891 66322 27925
rect 66876 27891 67340 27925
rect 67894 27891 68358 27925
rect 68912 27891 69376 27925
rect 69930 27891 70394 27925
rect 70948 27891 71412 27925
rect 71966 27891 72430 27925
rect 72984 27891 73448 27925
rect 74002 27891 74466 27925
rect 58438 27256 58472 27832
rect 59456 27256 59490 27832
rect 60474 27256 60508 27832
rect 61492 27256 61526 27832
rect 62510 27256 62544 27832
rect 63528 27256 63562 27832
rect 64546 27256 64580 27832
rect 65564 27256 65598 27832
rect 66582 27256 66616 27832
rect 67600 27256 67634 27832
rect 68618 27256 68652 27832
rect 69636 27256 69670 27832
rect 70654 27256 70688 27832
rect 71672 27256 71706 27832
rect 72690 27256 72724 27832
rect 73708 27256 73742 27832
rect 74726 27256 74760 27832
rect 58732 27163 59196 27197
rect 59750 27163 60214 27197
rect 60768 27163 61232 27197
rect 61786 27163 62250 27197
rect 62804 27163 63268 27197
rect 63822 27163 64286 27197
rect 64840 27163 65304 27197
rect 65858 27163 66322 27197
rect 66876 27163 67340 27197
rect 67894 27163 68358 27197
rect 68912 27163 69376 27197
rect 69930 27163 70394 27197
rect 70948 27163 71412 27197
rect 71966 27163 72430 27197
rect 72984 27163 73448 27197
rect 74002 27163 74466 27197
rect 58732 26755 59196 26789
rect 59750 26755 60214 26789
rect 60768 26755 61232 26789
rect 61786 26755 62250 26789
rect 62804 26755 63268 26789
rect 63822 26755 64286 26789
rect 64840 26755 65304 26789
rect 65858 26755 66322 26789
rect 66876 26755 67340 26789
rect 67894 26755 68358 26789
rect 68912 26755 69376 26789
rect 69930 26755 70394 26789
rect 70948 26755 71412 26789
rect 71966 26755 72430 26789
rect 72984 26755 73448 26789
rect 74002 26755 74466 26789
rect 58438 26120 58472 26696
rect 59456 26120 59490 26696
rect 60474 26120 60508 26696
rect 61492 26120 61526 26696
rect 62510 26120 62544 26696
rect 63528 26120 63562 26696
rect 64546 26120 64580 26696
rect 65564 26120 65598 26696
rect 66582 26120 66616 26696
rect 67600 26120 67634 26696
rect 68618 26120 68652 26696
rect 69636 26120 69670 26696
rect 70654 26120 70688 26696
rect 71672 26120 71706 26696
rect 72690 26120 72724 26696
rect 73708 26120 73742 26696
rect 74726 26120 74760 26696
rect 58732 26027 59196 26061
rect 59750 26027 60214 26061
rect 60768 26027 61232 26061
rect 61786 26027 62250 26061
rect 62804 26027 63268 26061
rect 63822 26027 64286 26061
rect 64840 26027 65304 26061
rect 65858 26027 66322 26061
rect 66876 26027 67340 26061
rect 67894 26027 68358 26061
rect 68912 26027 69376 26061
rect 69930 26027 70394 26061
rect 70948 26027 71412 26061
rect 71966 26027 72430 26061
rect 72984 26027 73448 26061
rect 74002 26027 74466 26061
rect 58732 25619 59196 25653
rect 59750 25619 60214 25653
rect 60768 25619 61232 25653
rect 61786 25619 62250 25653
rect 62804 25619 63268 25653
rect 63822 25619 64286 25653
rect 64840 25619 65304 25653
rect 65858 25619 66322 25653
rect 66876 25619 67340 25653
rect 67894 25619 68358 25653
rect 68912 25619 69376 25653
rect 69930 25619 70394 25653
rect 70948 25619 71412 25653
rect 71966 25619 72430 25653
rect 72984 25619 73448 25653
rect 74002 25619 74466 25653
rect 58438 24984 58472 25560
rect 59456 24984 59490 25560
rect 60474 24984 60508 25560
rect 61492 24984 61526 25560
rect 62510 24984 62544 25560
rect 63528 24984 63562 25560
rect 64546 24984 64580 25560
rect 65564 24984 65598 25560
rect 66582 24984 66616 25560
rect 67600 24984 67634 25560
rect 68618 24984 68652 25560
rect 69636 24984 69670 25560
rect 70654 24984 70688 25560
rect 71672 24984 71706 25560
rect 72690 24984 72724 25560
rect 73708 24984 73742 25560
rect 74726 24984 74760 25560
rect 58732 24891 59196 24925
rect 59750 24891 60214 24925
rect 60768 24891 61232 24925
rect 61786 24891 62250 24925
rect 62804 24891 63268 24925
rect 63822 24891 64286 24925
rect 64840 24891 65304 24925
rect 65858 24891 66322 24925
rect 66876 24891 67340 24925
rect 67894 24891 68358 24925
rect 68912 24891 69376 24925
rect 69930 24891 70394 24925
rect 70948 24891 71412 24925
rect 71966 24891 72430 24925
rect 72984 24891 73448 24925
rect 74002 24891 74466 24925
rect 59926 23981 60390 24015
rect 60944 23981 61408 24015
rect 61962 23981 62426 24015
rect 62980 23981 63444 24015
rect 63998 23981 64462 24015
rect 65016 23981 65480 24015
rect 66034 23981 66498 24015
rect 67052 23981 67516 24015
rect 68070 23981 68534 24015
rect 69088 23981 69552 24015
rect 70106 23981 70570 24015
rect 71124 23981 71588 24015
rect 72142 23981 72606 24015
rect 73160 23981 73624 24015
rect 59632 23346 59666 23922
rect 60650 23346 60684 23922
rect 61668 23346 61702 23922
rect 62686 23346 62720 23922
rect 63704 23346 63738 23922
rect 64722 23346 64756 23922
rect 65740 23346 65774 23922
rect 66758 23346 66792 23922
rect 67776 23346 67810 23922
rect 68794 23346 68828 23922
rect 69812 23346 69846 23922
rect 70830 23346 70864 23922
rect 71848 23346 71882 23922
rect 72866 23346 72900 23922
rect 73884 23346 73918 23922
rect 59926 23253 60390 23287
rect 60944 23253 61408 23287
rect 61962 23253 62426 23287
rect 62980 23253 63444 23287
rect 63998 23253 64462 23287
rect 65016 23253 65480 23287
rect 66034 23253 66498 23287
rect 67052 23253 67516 23287
rect 68070 23253 68534 23287
rect 69088 23253 69552 23287
rect 70106 23253 70570 23287
rect 71124 23253 71588 23287
rect 72142 23253 72606 23287
rect 73160 23253 73624 23287
rect 59926 22949 60390 22983
rect 60944 22949 61408 22983
rect 61962 22949 62426 22983
rect 62980 22949 63444 22983
rect 63998 22949 64462 22983
rect 65016 22949 65480 22983
rect 66034 22949 66498 22983
rect 67052 22949 67516 22983
rect 68070 22949 68534 22983
rect 69088 22949 69552 22983
rect 70106 22949 70570 22983
rect 71124 22949 71588 22983
rect 72142 22949 72606 22983
rect 73160 22949 73624 22983
rect 59632 22314 59666 22890
rect 60650 22314 60684 22890
rect 61668 22314 61702 22890
rect 62686 22314 62720 22890
rect 63704 22314 63738 22890
rect 64722 22314 64756 22890
rect 65740 22314 65774 22890
rect 66758 22314 66792 22890
rect 67776 22314 67810 22890
rect 68794 22314 68828 22890
rect 69812 22314 69846 22890
rect 70830 22314 70864 22890
rect 71848 22314 71882 22890
rect 72866 22314 72900 22890
rect 73884 22314 73918 22890
rect 59926 22221 60390 22255
rect 60944 22221 61408 22255
rect 61962 22221 62426 22255
rect 62980 22221 63444 22255
rect 63998 22221 64462 22255
rect 65016 22221 65480 22255
rect 66034 22221 66498 22255
rect 67052 22221 67516 22255
rect 68070 22221 68534 22255
rect 69088 22221 69552 22255
rect 70106 22221 70570 22255
rect 71124 22221 71588 22255
rect 72142 22221 72606 22255
rect 73160 22221 73624 22255
rect 59718 21345 60182 21379
rect 60736 21345 61200 21379
rect 61754 21345 62218 21379
rect 62772 21345 63236 21379
rect 63790 21345 64254 21379
rect 64808 21345 65272 21379
rect 65826 21345 66290 21379
rect 66844 21345 67308 21379
rect 67862 21345 68326 21379
rect 68880 21345 69344 21379
rect 69898 21345 70362 21379
rect 70916 21345 71380 21379
rect 71934 21345 72398 21379
rect 72952 21345 73416 21379
rect 73970 21345 74434 21379
rect 54414 21241 54878 21275
rect 55432 21241 55896 21275
rect 56450 21241 56914 21275
rect 57468 21241 57932 21275
rect 54120 20606 54154 21182
rect 55138 20606 55172 21182
rect 56156 20606 56190 21182
rect 57174 20606 57208 21182
rect 58192 20606 58226 21182
rect 59424 20710 59458 21286
rect 60442 20710 60476 21286
rect 61460 20710 61494 21286
rect 62478 20710 62512 21286
rect 63496 20710 63530 21286
rect 64514 20710 64548 21286
rect 65532 20710 65566 21286
rect 66550 20710 66584 21286
rect 67568 20710 67602 21286
rect 68586 20710 68620 21286
rect 69604 20710 69638 21286
rect 70622 20710 70656 21286
rect 71640 20710 71674 21286
rect 72658 20710 72692 21286
rect 73676 20710 73710 21286
rect 74694 20710 74728 21286
rect 59718 20617 60182 20651
rect 60736 20617 61200 20651
rect 61754 20617 62218 20651
rect 62772 20617 63236 20651
rect 63790 20617 64254 20651
rect 64808 20617 65272 20651
rect 65826 20617 66290 20651
rect 66844 20617 67308 20651
rect 67862 20617 68326 20651
rect 68880 20617 69344 20651
rect 69898 20617 70362 20651
rect 70916 20617 71380 20651
rect 71934 20617 72398 20651
rect 72952 20617 73416 20651
rect 73970 20617 74434 20651
rect 54414 20513 54878 20547
rect 55432 20513 55896 20547
rect 56450 20513 56914 20547
rect 57468 20513 57932 20547
rect 54414 20209 54878 20243
rect 55432 20209 55896 20243
rect 56450 20209 56914 20243
rect 57468 20209 57932 20243
rect 54120 19574 54154 20150
rect 55138 19574 55172 20150
rect 56156 19574 56190 20150
rect 57174 19574 57208 20150
rect 58192 19574 58226 20150
rect 59718 20089 60182 20123
rect 60736 20089 61200 20123
rect 61754 20089 62218 20123
rect 62772 20089 63236 20123
rect 63790 20089 64254 20123
rect 64808 20089 65272 20123
rect 65826 20089 66290 20123
rect 66844 20089 67308 20123
rect 67862 20089 68326 20123
rect 68880 20089 69344 20123
rect 69898 20089 70362 20123
rect 70916 20089 71380 20123
rect 71934 20089 72398 20123
rect 72952 20089 73416 20123
rect 73970 20089 74434 20123
rect 54414 19481 54878 19515
rect 55432 19481 55896 19515
rect 56450 19481 56914 19515
rect 57468 19481 57932 19515
rect 59424 19454 59458 20030
rect 60442 19454 60476 20030
rect 61460 19454 61494 20030
rect 62478 19454 62512 20030
rect 63496 19454 63530 20030
rect 64514 19454 64548 20030
rect 65532 19454 65566 20030
rect 66550 19454 66584 20030
rect 67568 19454 67602 20030
rect 68586 19454 68620 20030
rect 69604 19454 69638 20030
rect 70622 19454 70656 20030
rect 71640 19454 71674 20030
rect 72658 19454 72692 20030
rect 73676 19454 73710 20030
rect 74694 19454 74728 20030
rect 59718 19361 60182 19395
rect 60736 19361 61200 19395
rect 61754 19361 62218 19395
rect 62772 19361 63236 19395
rect 63790 19361 64254 19395
rect 64808 19361 65272 19395
rect 65826 19361 66290 19395
rect 66844 19361 67308 19395
rect 67862 19361 68326 19395
rect 68880 19361 69344 19395
rect 69898 19361 70362 19395
rect 70916 19361 71380 19395
rect 71934 19361 72398 19395
rect 72952 19361 73416 19395
rect 73970 19361 74434 19395
rect 54414 19177 54878 19211
rect 55432 19177 55896 19211
rect 56450 19177 56914 19211
rect 57468 19177 57932 19211
rect 54120 18542 54154 19118
rect 55138 18542 55172 19118
rect 56156 18542 56190 19118
rect 57174 18542 57208 19118
rect 58192 18542 58226 19118
rect 59718 18833 60182 18867
rect 60736 18833 61200 18867
rect 61754 18833 62218 18867
rect 62772 18833 63236 18867
rect 63790 18833 64254 18867
rect 64808 18833 65272 18867
rect 65826 18833 66290 18867
rect 66844 18833 67308 18867
rect 67862 18833 68326 18867
rect 68880 18833 69344 18867
rect 69898 18833 70362 18867
rect 70916 18833 71380 18867
rect 71934 18833 72398 18867
rect 72952 18833 73416 18867
rect 73970 18833 74434 18867
rect 54414 18449 54878 18483
rect 55432 18449 55896 18483
rect 56450 18449 56914 18483
rect 57468 18449 57932 18483
rect 59424 18198 59458 18774
rect 60442 18198 60476 18774
rect 61460 18198 61494 18774
rect 62478 18198 62512 18774
rect 63496 18198 63530 18774
rect 64514 18198 64548 18774
rect 65532 18198 65566 18774
rect 66550 18198 66584 18774
rect 67568 18198 67602 18774
rect 68586 18198 68620 18774
rect 69604 18198 69638 18774
rect 70622 18198 70656 18774
rect 71640 18198 71674 18774
rect 72658 18198 72692 18774
rect 73676 18198 73710 18774
rect 74694 18198 74728 18774
rect 54414 18145 54878 18179
rect 55432 18145 55896 18179
rect 56450 18145 56914 18179
rect 57468 18145 57932 18179
rect 59718 18105 60182 18139
rect 60736 18105 61200 18139
rect 61754 18105 62218 18139
rect 62772 18105 63236 18139
rect 63790 18105 64254 18139
rect 64808 18105 65272 18139
rect 65826 18105 66290 18139
rect 66844 18105 67308 18139
rect 67862 18105 68326 18139
rect 68880 18105 69344 18139
rect 69898 18105 70362 18139
rect 70916 18105 71380 18139
rect 71934 18105 72398 18139
rect 72952 18105 73416 18139
rect 73970 18105 74434 18139
rect 54120 17510 54154 18086
rect 55138 17510 55172 18086
rect 56156 17510 56190 18086
rect 57174 17510 57208 18086
rect 58192 17510 58226 18086
rect 59718 17577 60182 17611
rect 60736 17577 61200 17611
rect 61754 17577 62218 17611
rect 62772 17577 63236 17611
rect 63790 17577 64254 17611
rect 64808 17577 65272 17611
rect 65826 17577 66290 17611
rect 66844 17577 67308 17611
rect 67862 17577 68326 17611
rect 68880 17577 69344 17611
rect 69898 17577 70362 17611
rect 70916 17577 71380 17611
rect 71934 17577 72398 17611
rect 72952 17577 73416 17611
rect 73970 17577 74434 17611
rect 54414 17417 54878 17451
rect 55432 17417 55896 17451
rect 56450 17417 56914 17451
rect 57468 17417 57932 17451
rect 59424 16942 59458 17518
rect 60442 16942 60476 17518
rect 61460 16942 61494 17518
rect 62478 16942 62512 17518
rect 63496 16942 63530 17518
rect 64514 16942 64548 17518
rect 65532 16942 65566 17518
rect 66550 16942 66584 17518
rect 67568 16942 67602 17518
rect 68586 16942 68620 17518
rect 69604 16942 69638 17518
rect 70622 16942 70656 17518
rect 71640 16942 71674 17518
rect 72658 16942 72692 17518
rect 73676 16942 73710 17518
rect 74694 16942 74728 17518
rect 59718 16849 60182 16883
rect 60736 16849 61200 16883
rect 61754 16849 62218 16883
rect 62772 16849 63236 16883
rect 63790 16849 64254 16883
rect 64808 16849 65272 16883
rect 65826 16849 66290 16883
rect 66844 16849 67308 16883
rect 67862 16849 68326 16883
rect 68880 16849 69344 16883
rect 69898 16849 70362 16883
rect 70916 16849 71380 16883
rect 71934 16849 72398 16883
rect 72952 16849 73416 16883
rect 73970 16849 74434 16883
rect 76672 16642 76772 30072
rect 52428 16022 52490 16122
rect 52490 16022 76610 16122
rect 76610 16022 76672 16122
rect -1272 15092 -1210 15192
rect -1210 15092 35710 15192
rect 35710 15092 35772 15192
rect 13826 14372 14290 14406
rect 14844 14372 15308 14406
rect 15862 14372 16326 14406
rect 16880 14372 17344 14406
rect 17898 14372 18362 14406
rect 18916 14372 19380 14406
rect 19934 14372 20398 14406
rect 20952 14372 21416 14406
rect 21970 14372 22434 14406
rect 22988 14372 23452 14406
rect 24006 14372 24470 14406
rect 25024 14372 25488 14406
rect 26042 14372 26506 14406
rect 27060 14372 27524 14406
rect 28078 14372 28542 14406
rect 29096 14372 29560 14406
rect 30114 14372 30578 14406
rect 31132 14372 31596 14406
rect 32150 14372 32614 14406
rect 33168 14372 33632 14406
rect -1372 40 -1272 14300
rect 2060 13896 2524 13930
rect 3078 13896 3542 13930
rect 4096 13896 4560 13930
rect 5114 13896 5578 13930
rect 6132 13896 6596 13930
rect 7150 13896 7614 13930
rect 8168 13896 8632 13930
rect 9186 13896 9650 13930
rect 10204 13896 10668 13930
rect 1766 13270 1800 13846
rect 2784 13270 2818 13846
rect 3802 13270 3836 13846
rect 4820 13270 4854 13846
rect 5838 13270 5872 13846
rect 6856 13270 6890 13846
rect 7874 13270 7908 13846
rect 8892 13270 8926 13846
rect 9910 13270 9944 13846
rect 10928 13270 10962 13846
rect 13532 13746 13566 14322
rect 14550 13746 14584 14322
rect 15568 13746 15602 14322
rect 16586 13746 16620 14322
rect 17604 13746 17638 14322
rect 18622 13746 18656 14322
rect 19640 13746 19674 14322
rect 20658 13746 20692 14322
rect 21676 13746 21710 14322
rect 22694 13746 22728 14322
rect 23712 13746 23746 14322
rect 24730 13746 24764 14322
rect 25748 13746 25782 14322
rect 26766 13746 26800 14322
rect 27784 13746 27818 14322
rect 28802 13746 28836 14322
rect 29820 13746 29854 14322
rect 30838 13746 30872 14322
rect 31856 13746 31890 14322
rect 32874 13746 32908 14322
rect 33892 13746 33926 14322
rect 13826 13662 14290 13696
rect 14844 13662 15308 13696
rect 15862 13662 16326 13696
rect 16880 13662 17344 13696
rect 17898 13662 18362 13696
rect 18916 13662 19380 13696
rect 19934 13662 20398 13696
rect 20952 13662 21416 13696
rect 21970 13662 22434 13696
rect 22988 13662 23452 13696
rect 24006 13662 24470 13696
rect 25024 13662 25488 13696
rect 26042 13662 26506 13696
rect 27060 13662 27524 13696
rect 28078 13662 28542 13696
rect 29096 13662 29560 13696
rect 30114 13662 30578 13696
rect 31132 13662 31596 13696
rect 32150 13662 32614 13696
rect 33168 13662 33632 13696
rect 13826 13554 14290 13588
rect 14844 13554 15308 13588
rect 15862 13554 16326 13588
rect 16880 13554 17344 13588
rect 17898 13554 18362 13588
rect 18916 13554 19380 13588
rect 19934 13554 20398 13588
rect 20952 13554 21416 13588
rect 21970 13554 22434 13588
rect 22988 13554 23452 13588
rect 24006 13554 24470 13588
rect 25024 13554 25488 13588
rect 26042 13554 26506 13588
rect 27060 13554 27524 13588
rect 28078 13554 28542 13588
rect 29096 13554 29560 13588
rect 30114 13554 30578 13588
rect 31132 13554 31596 13588
rect 32150 13554 32614 13588
rect 33168 13554 33632 13588
rect 2060 13186 2524 13220
rect 3078 13186 3542 13220
rect 2060 13078 2524 13112
rect 4096 13186 4560 13220
rect 3078 13078 3542 13112
rect 5114 13186 5578 13220
rect 4096 13078 4560 13112
rect 6132 13186 6596 13220
rect 5114 13078 5578 13112
rect 7150 13186 7614 13220
rect 6132 13078 6596 13112
rect 8168 13186 8632 13220
rect 7150 13078 7614 13112
rect 9186 13186 9650 13220
rect 8168 13078 8632 13112
rect 10204 13186 10668 13220
rect 9186 13078 9650 13112
rect 10204 13078 10668 13112
rect 1766 12452 1800 13028
rect 2784 12452 2818 13028
rect 3802 12452 3836 13028
rect 4820 12452 4854 13028
rect 5838 12452 5872 13028
rect 6856 12452 6890 13028
rect 7874 12452 7908 13028
rect 8892 12452 8926 13028
rect 9910 12452 9944 13028
rect 10928 12452 10962 13028
rect 13532 12928 13566 13504
rect 14550 12928 14584 13504
rect 15568 12928 15602 13504
rect 16586 12928 16620 13504
rect 17604 12928 17638 13504
rect 18622 12928 18656 13504
rect 19640 12928 19674 13504
rect 20658 12928 20692 13504
rect 21676 12928 21710 13504
rect 22694 12928 22728 13504
rect 23712 12928 23746 13504
rect 24730 12928 24764 13504
rect 25748 12928 25782 13504
rect 26766 12928 26800 13504
rect 27784 12928 27818 13504
rect 28802 12928 28836 13504
rect 29820 12928 29854 13504
rect 30838 12928 30872 13504
rect 31856 12928 31890 13504
rect 32874 12928 32908 13504
rect 33892 12928 33926 13504
rect 13826 12844 14290 12878
rect 14844 12844 15308 12878
rect 15862 12844 16326 12878
rect 16880 12844 17344 12878
rect 17898 12844 18362 12878
rect 18916 12844 19380 12878
rect 19934 12844 20398 12878
rect 20952 12844 21416 12878
rect 21970 12844 22434 12878
rect 22988 12844 23452 12878
rect 24006 12844 24470 12878
rect 25024 12844 25488 12878
rect 26042 12844 26506 12878
rect 27060 12844 27524 12878
rect 28078 12844 28542 12878
rect 29096 12844 29560 12878
rect 30114 12844 30578 12878
rect 31132 12844 31596 12878
rect 32150 12844 32614 12878
rect 33168 12844 33632 12878
rect 2060 12368 2524 12402
rect 3078 12368 3542 12402
rect 2060 12260 2524 12294
rect 4096 12368 4560 12402
rect 3078 12260 3542 12294
rect 5114 12368 5578 12402
rect 4096 12260 4560 12294
rect 6132 12368 6596 12402
rect 5114 12260 5578 12294
rect 7150 12368 7614 12402
rect 6132 12260 6596 12294
rect 8168 12368 8632 12402
rect 7150 12260 7614 12294
rect 9186 12368 9650 12402
rect 8168 12260 8632 12294
rect 10204 12368 10668 12402
rect 9186 12260 9650 12294
rect 10204 12260 10668 12294
rect 1766 11634 1800 12210
rect 2784 11634 2818 12210
rect 3802 11634 3836 12210
rect 4820 11634 4854 12210
rect 5838 11634 5872 12210
rect 6856 11634 6890 12210
rect 7874 11634 7908 12210
rect 8892 11634 8926 12210
rect 9910 11634 9944 12210
rect 10928 11634 10962 12210
rect 13826 12176 14290 12210
rect 14844 12176 15308 12210
rect 15862 12176 16326 12210
rect 16880 12176 17344 12210
rect 17898 12176 18362 12210
rect 18916 12176 19380 12210
rect 19934 12176 20398 12210
rect 20952 12176 21416 12210
rect 21970 12176 22434 12210
rect 22988 12176 23452 12210
rect 24006 12176 24470 12210
rect 25024 12176 25488 12210
rect 26042 12176 26506 12210
rect 27060 12176 27524 12210
rect 28078 12176 28542 12210
rect 29096 12176 29560 12210
rect 30114 12176 30578 12210
rect 31132 12176 31596 12210
rect 32150 12176 32614 12210
rect 33168 12176 33632 12210
rect 2060 11550 2524 11584
rect 3078 11550 3542 11584
rect 2060 11442 2524 11476
rect 4096 11550 4560 11584
rect 3078 11442 3542 11476
rect 5114 11550 5578 11584
rect 4096 11442 4560 11476
rect 6132 11550 6596 11584
rect 5114 11442 5578 11476
rect 7150 11550 7614 11584
rect 6132 11442 6596 11476
rect 8168 11550 8632 11584
rect 7150 11442 7614 11476
rect 9186 11550 9650 11584
rect 8168 11442 8632 11476
rect 10204 11550 10668 11584
rect 9186 11442 9650 11476
rect 13532 11550 13566 12126
rect 14550 11550 14584 12126
rect 15568 11550 15602 12126
rect 16586 11550 16620 12126
rect 17604 11550 17638 12126
rect 18622 11550 18656 12126
rect 19640 11550 19674 12126
rect 20658 11550 20692 12126
rect 21676 11550 21710 12126
rect 22694 11550 22728 12126
rect 23712 11550 23746 12126
rect 24730 11550 24764 12126
rect 25748 11550 25782 12126
rect 26766 11550 26800 12126
rect 27784 11550 27818 12126
rect 28802 11550 28836 12126
rect 29820 11550 29854 12126
rect 30838 11550 30872 12126
rect 31856 11550 31890 12126
rect 32874 11550 32908 12126
rect 33892 11550 33926 12126
rect 10204 11442 10668 11476
rect 13826 11466 14290 11500
rect 14844 11466 15308 11500
rect 15862 11466 16326 11500
rect 16880 11466 17344 11500
rect 17898 11466 18362 11500
rect 18916 11466 19380 11500
rect 19934 11466 20398 11500
rect 20952 11466 21416 11500
rect 21970 11466 22434 11500
rect 22988 11466 23452 11500
rect 24006 11466 24470 11500
rect 25024 11466 25488 11500
rect 26042 11466 26506 11500
rect 27060 11466 27524 11500
rect 28078 11466 28542 11500
rect 29096 11466 29560 11500
rect 30114 11466 30578 11500
rect 31132 11466 31596 11500
rect 32150 11466 32614 11500
rect 33168 11466 33632 11500
rect 1766 10816 1800 11392
rect 2784 10816 2818 11392
rect 3802 10816 3836 11392
rect 4820 10816 4854 11392
rect 5838 10816 5872 11392
rect 6856 10816 6890 11392
rect 7874 10816 7908 11392
rect 8892 10816 8926 11392
rect 9910 10816 9944 11392
rect 10928 10816 10962 11392
rect 13826 10944 14290 10978
rect 14844 10944 15308 10978
rect 15862 10944 16326 10978
rect 16880 10944 17344 10978
rect 17898 10944 18362 10978
rect 18916 10944 19380 10978
rect 19934 10944 20398 10978
rect 20952 10944 21416 10978
rect 21970 10944 22434 10978
rect 22988 10944 23452 10978
rect 24006 10944 24470 10978
rect 25024 10944 25488 10978
rect 26042 10944 26506 10978
rect 27060 10944 27524 10978
rect 28078 10944 28542 10978
rect 29096 10944 29560 10978
rect 30114 10944 30578 10978
rect 31132 10944 31596 10978
rect 32150 10944 32614 10978
rect 33168 10944 33632 10978
rect 2060 10732 2524 10766
rect 3078 10732 3542 10766
rect 2060 10624 2524 10658
rect 4096 10732 4560 10766
rect 3078 10624 3542 10658
rect 5114 10732 5578 10766
rect 4096 10624 4560 10658
rect 6132 10732 6596 10766
rect 5114 10624 5578 10658
rect 7150 10732 7614 10766
rect 6132 10624 6596 10658
rect 8168 10732 8632 10766
rect 7150 10624 7614 10658
rect 9186 10732 9650 10766
rect 8168 10624 8632 10658
rect 10204 10732 10668 10766
rect 9186 10624 9650 10658
rect 10204 10624 10668 10658
rect 1766 9998 1800 10574
rect 2784 9998 2818 10574
rect 3802 9998 3836 10574
rect 4820 9998 4854 10574
rect 5838 9998 5872 10574
rect 6856 9998 6890 10574
rect 7874 9998 7908 10574
rect 8892 9998 8926 10574
rect 9910 9998 9944 10574
rect 10928 9998 10962 10574
rect 13532 10318 13566 10894
rect 14550 10318 14584 10894
rect 15568 10318 15602 10894
rect 16586 10318 16620 10894
rect 17604 10318 17638 10894
rect 18622 10318 18656 10894
rect 19640 10318 19674 10894
rect 20658 10318 20692 10894
rect 21676 10318 21710 10894
rect 22694 10318 22728 10894
rect 23712 10318 23746 10894
rect 24730 10318 24764 10894
rect 25748 10318 25782 10894
rect 26766 10318 26800 10894
rect 27784 10318 27818 10894
rect 28802 10318 28836 10894
rect 29820 10318 29854 10894
rect 30838 10318 30872 10894
rect 31856 10318 31890 10894
rect 32874 10318 32908 10894
rect 33892 10318 33926 10894
rect 13826 10234 14290 10268
rect 14844 10234 15308 10268
rect 15862 10234 16326 10268
rect 16880 10234 17344 10268
rect 17898 10234 18362 10268
rect 18916 10234 19380 10268
rect 19934 10234 20398 10268
rect 20952 10234 21416 10268
rect 21970 10234 22434 10268
rect 22988 10234 23452 10268
rect 24006 10234 24470 10268
rect 25024 10234 25488 10268
rect 26042 10234 26506 10268
rect 27060 10234 27524 10268
rect 28078 10234 28542 10268
rect 29096 10234 29560 10268
rect 30114 10234 30578 10268
rect 31132 10234 31596 10268
rect 32150 10234 32614 10268
rect 33168 10234 33632 10268
rect 2060 9914 2524 9948
rect 3078 9914 3542 9948
rect 2060 9806 2524 9840
rect 4096 9914 4560 9948
rect 3078 9806 3542 9840
rect 5114 9914 5578 9948
rect 4096 9806 4560 9840
rect 6132 9914 6596 9948
rect 5114 9806 5578 9840
rect 7150 9914 7614 9948
rect 6132 9806 6596 9840
rect 8168 9914 8632 9948
rect 7150 9806 7614 9840
rect 9186 9914 9650 9948
rect 8168 9806 8632 9840
rect 10204 9914 10668 9948
rect 9186 9806 9650 9840
rect 10204 9806 10668 9840
rect 1766 9180 1800 9756
rect 2784 9180 2818 9756
rect 3802 9180 3836 9756
rect 4820 9180 4854 9756
rect 5838 9180 5872 9756
rect 6856 9180 6890 9756
rect 7874 9180 7908 9756
rect 8892 9180 8926 9756
rect 9910 9180 9944 9756
rect 10928 9180 10962 9756
rect 13824 9710 14288 9744
rect 14842 9710 15306 9744
rect 15860 9710 16324 9744
rect 16878 9710 17342 9744
rect 17896 9710 18360 9744
rect 18914 9710 19378 9744
rect 19932 9710 20396 9744
rect 20950 9710 21414 9744
rect 21968 9710 22432 9744
rect 22986 9710 23450 9744
rect 24004 9710 24468 9744
rect 25022 9710 25486 9744
rect 26040 9710 26504 9744
rect 27058 9710 27522 9744
rect 28076 9710 28540 9744
rect 29094 9710 29558 9744
rect 30112 9710 30576 9744
rect 31130 9710 31594 9744
rect 32148 9710 32612 9744
rect 33166 9710 33630 9744
rect 2060 9096 2524 9130
rect 3078 9096 3542 9130
rect 2060 8988 2524 9022
rect 4096 9096 4560 9130
rect 3078 8988 3542 9022
rect 5114 9096 5578 9130
rect 4096 8988 4560 9022
rect 6132 9096 6596 9130
rect 5114 8988 5578 9022
rect 7150 9096 7614 9130
rect 6132 8988 6596 9022
rect 8168 9096 8632 9130
rect 7150 8988 7614 9022
rect 9186 9096 9650 9130
rect 8168 8988 8632 9022
rect 10204 9096 10668 9130
rect 9186 8988 9650 9022
rect 13530 9084 13564 9660
rect 14548 9084 14582 9660
rect 15566 9084 15600 9660
rect 16584 9084 16618 9660
rect 17602 9084 17636 9660
rect 18620 9084 18654 9660
rect 19638 9084 19672 9660
rect 20656 9084 20690 9660
rect 21674 9084 21708 9660
rect 22692 9084 22726 9660
rect 23710 9084 23744 9660
rect 24728 9084 24762 9660
rect 25746 9084 25780 9660
rect 26764 9084 26798 9660
rect 27782 9084 27816 9660
rect 28800 9084 28834 9660
rect 29818 9084 29852 9660
rect 30836 9084 30870 9660
rect 31854 9084 31888 9660
rect 32872 9084 32906 9660
rect 33890 9084 33924 9660
rect 10204 8988 10668 9022
rect 13824 9000 14288 9034
rect 14842 9000 15306 9034
rect 15860 9000 16324 9034
rect 16878 9000 17342 9034
rect 17896 9000 18360 9034
rect 18914 9000 19378 9034
rect 19932 9000 20396 9034
rect 20950 9000 21414 9034
rect 21968 9000 22432 9034
rect 22986 9000 23450 9034
rect 24004 9000 24468 9034
rect 25022 9000 25486 9034
rect 26040 9000 26504 9034
rect 27058 9000 27522 9034
rect 28076 9000 28540 9034
rect 29094 9000 29558 9034
rect 30112 9000 30576 9034
rect 31130 9000 31594 9034
rect 32148 9000 32612 9034
rect 33166 9000 33630 9034
rect 1766 8362 1800 8938
rect 2784 8362 2818 8938
rect 3802 8362 3836 8938
rect 4820 8362 4854 8938
rect 5838 8362 5872 8938
rect 6856 8362 6890 8938
rect 7874 8362 7908 8938
rect 8892 8362 8926 8938
rect 9910 8362 9944 8938
rect 10928 8362 10962 8938
rect 13824 8476 14288 8510
rect 14842 8476 15306 8510
rect 15860 8476 16324 8510
rect 16878 8476 17342 8510
rect 17896 8476 18360 8510
rect 18914 8476 19378 8510
rect 19932 8476 20396 8510
rect 20950 8476 21414 8510
rect 21968 8476 22432 8510
rect 22986 8476 23450 8510
rect 24004 8476 24468 8510
rect 25022 8476 25486 8510
rect 26040 8476 26504 8510
rect 27058 8476 27522 8510
rect 28076 8476 28540 8510
rect 29094 8476 29558 8510
rect 30112 8476 30576 8510
rect 31130 8476 31594 8510
rect 32148 8476 32612 8510
rect 33166 8476 33630 8510
rect 2060 8278 2524 8312
rect 3078 8278 3542 8312
rect 2060 8170 2524 8204
rect 4096 8278 4560 8312
rect 3078 8170 3542 8204
rect 5114 8278 5578 8312
rect 4096 8170 4560 8204
rect 6132 8278 6596 8312
rect 5114 8170 5578 8204
rect 7150 8278 7614 8312
rect 6132 8170 6596 8204
rect 8168 8278 8632 8312
rect 7150 8170 7614 8204
rect 9186 8278 9650 8312
rect 8168 8170 8632 8204
rect 10204 8278 10668 8312
rect 9186 8170 9650 8204
rect 10204 8170 10668 8204
rect 1766 7544 1800 8120
rect 2784 7544 2818 8120
rect 3802 7544 3836 8120
rect 4820 7544 4854 8120
rect 5838 7544 5872 8120
rect 6856 7544 6890 8120
rect 7874 7544 7908 8120
rect 8892 7544 8926 8120
rect 9910 7544 9944 8120
rect 10928 7544 10962 8120
rect 13530 7850 13564 8426
rect 14548 7850 14582 8426
rect 15566 7850 15600 8426
rect 16584 7850 16618 8426
rect 17602 7850 17636 8426
rect 18620 7850 18654 8426
rect 19638 7850 19672 8426
rect 20656 7850 20690 8426
rect 21674 7850 21708 8426
rect 22692 7850 22726 8426
rect 23710 7850 23744 8426
rect 24728 7850 24762 8426
rect 25746 7850 25780 8426
rect 26764 7850 26798 8426
rect 27782 7850 27816 8426
rect 28800 7850 28834 8426
rect 29818 7850 29852 8426
rect 30836 7850 30870 8426
rect 31854 7850 31888 8426
rect 32872 7850 32906 8426
rect 33890 7850 33924 8426
rect 13824 7766 14288 7800
rect 14842 7766 15306 7800
rect 15860 7766 16324 7800
rect 16878 7766 17342 7800
rect 17896 7766 18360 7800
rect 18914 7766 19378 7800
rect 19932 7766 20396 7800
rect 20950 7766 21414 7800
rect 21968 7766 22432 7800
rect 22986 7766 23450 7800
rect 24004 7766 24468 7800
rect 25022 7766 25486 7800
rect 26040 7766 26504 7800
rect 27058 7766 27522 7800
rect 28076 7766 28540 7800
rect 29094 7766 29558 7800
rect 30112 7766 30576 7800
rect 31130 7766 31594 7800
rect 32148 7766 32612 7800
rect 33166 7766 33630 7800
rect 2060 7460 2524 7494
rect 3078 7460 3542 7494
rect 4096 7460 4560 7494
rect 5114 7460 5578 7494
rect 6132 7460 6596 7494
rect 7150 7460 7614 7494
rect 8168 7460 8632 7494
rect 9186 7460 9650 7494
rect 10204 7460 10668 7494
rect 13824 7244 14288 7278
rect 14842 7244 15306 7278
rect 15860 7244 16324 7278
rect 16878 7244 17342 7278
rect 17896 7244 18360 7278
rect 18914 7244 19378 7278
rect 19932 7244 20396 7278
rect 20950 7244 21414 7278
rect 21968 7244 22432 7278
rect 22986 7244 23450 7278
rect 24004 7244 24468 7278
rect 25022 7244 25486 7278
rect 26040 7244 26504 7278
rect 27058 7244 27522 7278
rect 28076 7244 28540 7278
rect 29094 7244 29558 7278
rect 30112 7244 30576 7278
rect 31130 7244 31594 7278
rect 32148 7244 32612 7278
rect 33166 7244 33630 7278
rect 13530 6618 13564 7194
rect 14548 6618 14582 7194
rect 15566 6618 15600 7194
rect 16584 6618 16618 7194
rect 17602 6618 17636 7194
rect 18620 6618 18654 7194
rect 19638 6618 19672 7194
rect 20656 6618 20690 7194
rect 21674 6618 21708 7194
rect 22692 6618 22726 7194
rect 23710 6618 23744 7194
rect 24728 6618 24762 7194
rect 25746 6618 25780 7194
rect 26764 6618 26798 7194
rect 27782 6618 27816 7194
rect 28800 6618 28834 7194
rect 29818 6618 29852 7194
rect 30836 6618 30870 7194
rect 31854 6618 31888 7194
rect 32872 6618 32906 7194
rect 33890 6618 33924 7194
rect 13824 6534 14288 6568
rect 14842 6534 15306 6568
rect 15860 6534 16324 6568
rect 16878 6534 17342 6568
rect 17896 6534 18360 6568
rect 18914 6534 19378 6568
rect 19932 6534 20396 6568
rect 20950 6534 21414 6568
rect 21968 6534 22432 6568
rect 22986 6534 23450 6568
rect 24004 6534 24468 6568
rect 25022 6534 25486 6568
rect 26040 6534 26504 6568
rect 27058 6534 27522 6568
rect 28076 6534 28540 6568
rect 29094 6534 29558 6568
rect 30112 6534 30576 6568
rect 31130 6534 31594 6568
rect 32148 6534 32612 6568
rect 33166 6534 33630 6568
rect 736 6146 1200 6180
rect 1754 6146 2218 6180
rect 2772 6146 3236 6180
rect 3790 6146 4254 6180
rect 4808 6146 5272 6180
rect 5826 6146 6290 6180
rect 6844 6146 7308 6180
rect 7862 6146 8326 6180
rect 8880 6146 9344 6180
rect 9898 6146 10362 6180
rect 10916 6146 11380 6180
rect 442 5520 476 6096
rect 1460 5520 1494 6096
rect 2478 5520 2512 6096
rect 3496 5520 3530 6096
rect 4514 5520 4548 6096
rect 5532 5520 5566 6096
rect 6550 5520 6584 6096
rect 7568 5520 7602 6096
rect 8586 5520 8620 6096
rect 9604 5520 9638 6096
rect 10622 5520 10656 6096
rect 11640 5520 11674 6096
rect 13824 6010 14288 6044
rect 14842 6010 15306 6044
rect 15860 6010 16324 6044
rect 16878 6010 17342 6044
rect 17896 6010 18360 6044
rect 18914 6010 19378 6044
rect 19932 6010 20396 6044
rect 20950 6010 21414 6044
rect 21968 6010 22432 6044
rect 22986 6010 23450 6044
rect 24004 6010 24468 6044
rect 25022 6010 25486 6044
rect 26040 6010 26504 6044
rect 27058 6010 27522 6044
rect 28076 6010 28540 6044
rect 29094 6010 29558 6044
rect 30112 6010 30576 6044
rect 31130 6010 31594 6044
rect 32148 6010 32612 6044
rect 33166 6010 33630 6044
rect 736 5436 1200 5470
rect 1754 5436 2218 5470
rect 2772 5436 3236 5470
rect 3790 5436 4254 5470
rect 4808 5436 5272 5470
rect 5826 5436 6290 5470
rect 6844 5436 7308 5470
rect 7862 5436 8326 5470
rect 8880 5436 9344 5470
rect 9898 5436 10362 5470
rect 10916 5436 11380 5470
rect 13530 5384 13564 5960
rect 14548 5384 14582 5960
rect 15566 5384 15600 5960
rect 16584 5384 16618 5960
rect 17602 5384 17636 5960
rect 18620 5384 18654 5960
rect 19638 5384 19672 5960
rect 20656 5384 20690 5960
rect 21674 5384 21708 5960
rect 22692 5384 22726 5960
rect 23710 5384 23744 5960
rect 24728 5384 24762 5960
rect 25746 5384 25780 5960
rect 26764 5384 26798 5960
rect 27782 5384 27816 5960
rect 28800 5384 28834 5960
rect 29818 5384 29852 5960
rect 30836 5384 30870 5960
rect 31854 5384 31888 5960
rect 32872 5384 32906 5960
rect 33890 5384 33924 5960
rect 13824 5300 14288 5334
rect 14842 5300 15306 5334
rect 15860 5300 16324 5334
rect 16878 5300 17342 5334
rect 17896 5300 18360 5334
rect 18914 5300 19378 5334
rect 19932 5300 20396 5334
rect 20950 5300 21414 5334
rect 21968 5300 22432 5334
rect 22986 5300 23450 5334
rect 24004 5300 24468 5334
rect 25022 5300 25486 5334
rect 26040 5300 26504 5334
rect 27058 5300 27522 5334
rect 28076 5300 28540 5334
rect 29094 5300 29558 5334
rect 30112 5300 30576 5334
rect 31130 5300 31594 5334
rect 32148 5300 32612 5334
rect 33166 5300 33630 5334
rect 736 5034 1200 5068
rect 1754 5034 2218 5068
rect 2772 5034 3236 5068
rect 3790 5034 4254 5068
rect 4808 5034 5272 5068
rect 5826 5034 6290 5068
rect 6844 5034 7308 5068
rect 7862 5034 8326 5068
rect 8880 5034 9344 5068
rect 9898 5034 10362 5068
rect 10916 5034 11380 5068
rect 442 4408 476 4984
rect 1460 4408 1494 4984
rect 2478 4408 2512 4984
rect 3496 4408 3530 4984
rect 4514 4408 4548 4984
rect 5532 4408 5566 4984
rect 6550 4408 6584 4984
rect 7568 4408 7602 4984
rect 8586 4408 8620 4984
rect 9604 4408 9638 4984
rect 10622 4408 10656 4984
rect 11640 4408 11674 4984
rect 13824 4776 14288 4810
rect 14842 4776 15306 4810
rect 15860 4776 16324 4810
rect 16878 4776 17342 4810
rect 17896 4776 18360 4810
rect 18914 4776 19378 4810
rect 19932 4776 20396 4810
rect 20950 4776 21414 4810
rect 21968 4776 22432 4810
rect 22986 4776 23450 4810
rect 24004 4776 24468 4810
rect 25022 4776 25486 4810
rect 26040 4776 26504 4810
rect 27058 4776 27522 4810
rect 28076 4776 28540 4810
rect 29094 4776 29558 4810
rect 30112 4776 30576 4810
rect 31130 4776 31594 4810
rect 32148 4776 32612 4810
rect 33166 4776 33630 4810
rect 736 4324 1200 4358
rect 1754 4324 2218 4358
rect 2772 4324 3236 4358
rect 3790 4324 4254 4358
rect 4808 4324 5272 4358
rect 5826 4324 6290 4358
rect 6844 4324 7308 4358
rect 7862 4324 8326 4358
rect 8880 4324 9344 4358
rect 9898 4324 10362 4358
rect 10916 4324 11380 4358
rect 13530 4150 13564 4726
rect 14548 4150 14582 4726
rect 15566 4150 15600 4726
rect 16584 4150 16618 4726
rect 17602 4150 17636 4726
rect 18620 4150 18654 4726
rect 19638 4150 19672 4726
rect 20656 4150 20690 4726
rect 21674 4150 21708 4726
rect 22692 4150 22726 4726
rect 23710 4150 23744 4726
rect 24728 4150 24762 4726
rect 25746 4150 25780 4726
rect 26764 4150 26798 4726
rect 27782 4150 27816 4726
rect 28800 4150 28834 4726
rect 29818 4150 29852 4726
rect 30836 4150 30870 4726
rect 31854 4150 31888 4726
rect 32872 4150 32906 4726
rect 33890 4150 33924 4726
rect 13824 4066 14288 4100
rect 14842 4066 15306 4100
rect 15860 4066 16324 4100
rect 16878 4066 17342 4100
rect 17896 4066 18360 4100
rect 18914 4066 19378 4100
rect 19932 4066 20396 4100
rect 20950 4066 21414 4100
rect 21968 4066 22432 4100
rect 22986 4066 23450 4100
rect 24004 4066 24468 4100
rect 25022 4066 25486 4100
rect 26040 4066 26504 4100
rect 27058 4066 27522 4100
rect 28076 4066 28540 4100
rect 29094 4066 29558 4100
rect 30112 4066 30576 4100
rect 31130 4066 31594 4100
rect 32148 4066 32612 4100
rect 33166 4066 33630 4100
rect 736 3922 1200 3956
rect 1754 3922 2218 3956
rect 2772 3922 3236 3956
rect 3790 3922 4254 3956
rect 4808 3922 5272 3956
rect 5826 3922 6290 3956
rect 6844 3922 7308 3956
rect 7862 3922 8326 3956
rect 8880 3922 9344 3956
rect 9898 3922 10362 3956
rect 10916 3922 11380 3956
rect 442 3296 476 3872
rect 1460 3296 1494 3872
rect 2478 3296 2512 3872
rect 3496 3296 3530 3872
rect 4514 3296 4548 3872
rect 5532 3296 5566 3872
rect 6550 3296 6584 3872
rect 7568 3296 7602 3872
rect 8586 3296 8620 3872
rect 9604 3296 9638 3872
rect 10622 3296 10656 3872
rect 11640 3296 11674 3872
rect 13824 3544 14288 3578
rect 14842 3544 15306 3578
rect 15860 3544 16324 3578
rect 16878 3544 17342 3578
rect 17896 3544 18360 3578
rect 18914 3544 19378 3578
rect 19932 3544 20396 3578
rect 20950 3544 21414 3578
rect 21968 3544 22432 3578
rect 22986 3544 23450 3578
rect 24004 3544 24468 3578
rect 25022 3544 25486 3578
rect 26040 3544 26504 3578
rect 27058 3544 27522 3578
rect 28076 3544 28540 3578
rect 29094 3544 29558 3578
rect 30112 3544 30576 3578
rect 31130 3544 31594 3578
rect 32148 3544 32612 3578
rect 33166 3544 33630 3578
rect 736 3212 1200 3246
rect 1754 3212 2218 3246
rect 2772 3212 3236 3246
rect 3790 3212 4254 3246
rect 4808 3212 5272 3246
rect 5826 3212 6290 3246
rect 6844 3212 7308 3246
rect 7862 3212 8326 3246
rect 8880 3212 9344 3246
rect 9898 3212 10362 3246
rect 10916 3212 11380 3246
rect 13530 2918 13564 3494
rect 14548 2918 14582 3494
rect 15566 2918 15600 3494
rect 16584 2918 16618 3494
rect 17602 2918 17636 3494
rect 18620 2918 18654 3494
rect 19638 2918 19672 3494
rect 20656 2918 20690 3494
rect 21674 2918 21708 3494
rect 22692 2918 22726 3494
rect 23710 2918 23744 3494
rect 24728 2918 24762 3494
rect 25746 2918 25780 3494
rect 26764 2918 26798 3494
rect 27782 2918 27816 3494
rect 28800 2918 28834 3494
rect 29818 2918 29852 3494
rect 30836 2918 30870 3494
rect 31854 2918 31888 3494
rect 32872 2918 32906 3494
rect 33890 2918 33924 3494
rect 736 2810 1200 2844
rect 1754 2810 2218 2844
rect 2772 2810 3236 2844
rect 3790 2810 4254 2844
rect 4808 2810 5272 2844
rect 5826 2810 6290 2844
rect 6844 2810 7308 2844
rect 7862 2810 8326 2844
rect 8880 2810 9344 2844
rect 9898 2810 10362 2844
rect 10916 2810 11380 2844
rect 13824 2834 14288 2868
rect 14842 2834 15306 2868
rect 15860 2834 16324 2868
rect 16878 2834 17342 2868
rect 17896 2834 18360 2868
rect 18914 2834 19378 2868
rect 19932 2834 20396 2868
rect 20950 2834 21414 2868
rect 21968 2834 22432 2868
rect 22986 2834 23450 2868
rect 24004 2834 24468 2868
rect 25022 2834 25486 2868
rect 26040 2834 26504 2868
rect 27058 2834 27522 2868
rect 28076 2834 28540 2868
rect 29094 2834 29558 2868
rect 30112 2834 30576 2868
rect 31130 2834 31594 2868
rect 32148 2834 32612 2868
rect 33166 2834 33630 2868
rect 442 2184 476 2760
rect 1460 2184 1494 2760
rect 2478 2184 2512 2760
rect 3496 2184 3530 2760
rect 4514 2184 4548 2760
rect 5532 2184 5566 2760
rect 6550 2184 6584 2760
rect 7568 2184 7602 2760
rect 8586 2184 8620 2760
rect 9604 2184 9638 2760
rect 10622 2184 10656 2760
rect 11640 2184 11674 2760
rect 13824 2310 14288 2344
rect 14842 2310 15306 2344
rect 15860 2310 16324 2344
rect 16878 2310 17342 2344
rect 17896 2310 18360 2344
rect 18914 2310 19378 2344
rect 19932 2310 20396 2344
rect 20950 2310 21414 2344
rect 21968 2310 22432 2344
rect 22986 2310 23450 2344
rect 24004 2310 24468 2344
rect 25022 2310 25486 2344
rect 26040 2310 26504 2344
rect 27058 2310 27522 2344
rect 28076 2310 28540 2344
rect 29094 2310 29558 2344
rect 30112 2310 30576 2344
rect 31130 2310 31594 2344
rect 32148 2310 32612 2344
rect 33166 2310 33630 2344
rect 736 2100 1200 2134
rect 1754 2100 2218 2134
rect 2772 2100 3236 2134
rect 3790 2100 4254 2134
rect 4808 2100 5272 2134
rect 5826 2100 6290 2134
rect 6844 2100 7308 2134
rect 7862 2100 8326 2134
rect 8880 2100 9344 2134
rect 9898 2100 10362 2134
rect 10916 2100 11380 2134
rect 13530 1684 13564 2260
rect 14548 1684 14582 2260
rect 15566 1684 15600 2260
rect 16584 1684 16618 2260
rect 17602 1684 17636 2260
rect 18620 1684 18654 2260
rect 19638 1684 19672 2260
rect 20656 1684 20690 2260
rect 21674 1684 21708 2260
rect 22692 1684 22726 2260
rect 23710 1684 23744 2260
rect 24728 1684 24762 2260
rect 25746 1684 25780 2260
rect 26764 1684 26798 2260
rect 27782 1684 27816 2260
rect 28800 1684 28834 2260
rect 29818 1684 29852 2260
rect 30836 1684 30870 2260
rect 31854 1684 31888 2260
rect 32872 1684 32906 2260
rect 33890 1684 33924 2260
rect 13824 1600 14288 1634
rect 14842 1600 15306 1634
rect 15860 1600 16324 1634
rect 16878 1600 17342 1634
rect 17896 1600 18360 1634
rect 18914 1600 19378 1634
rect 19932 1600 20396 1634
rect 20950 1600 21414 1634
rect 21968 1600 22432 1634
rect 22986 1600 23450 1634
rect 24004 1600 24468 1634
rect 25022 1600 25486 1634
rect 26040 1600 26504 1634
rect 27058 1600 27522 1634
rect 28076 1600 28540 1634
rect 29094 1600 29558 1634
rect 30112 1600 30576 1634
rect 31130 1600 31594 1634
rect 32148 1600 32612 1634
rect 33166 1600 33630 1634
rect 1194 1268 1658 1302
rect 2212 1268 2676 1302
rect 3230 1268 3694 1302
rect 4248 1268 4712 1302
rect 5266 1268 5730 1302
rect 6284 1268 6748 1302
rect 7302 1268 7766 1302
rect 8320 1268 8784 1302
rect 9338 1268 9802 1302
rect 10356 1268 10820 1302
rect 900 642 934 1218
rect 1918 642 1952 1218
rect 2936 642 2970 1218
rect 3954 642 3988 1218
rect 4972 642 5006 1218
rect 5990 642 6024 1218
rect 7008 642 7042 1218
rect 8026 642 8060 1218
rect 9044 642 9078 1218
rect 10062 642 10096 1218
rect 11080 642 11114 1218
rect 13824 1078 14288 1112
rect 14842 1078 15306 1112
rect 15860 1078 16324 1112
rect 16878 1078 17342 1112
rect 17896 1078 18360 1112
rect 18914 1078 19378 1112
rect 19932 1078 20396 1112
rect 20950 1078 21414 1112
rect 21968 1078 22432 1112
rect 22986 1078 23450 1112
rect 24004 1078 24468 1112
rect 25022 1078 25486 1112
rect 26040 1078 26504 1112
rect 27058 1078 27522 1112
rect 28076 1078 28540 1112
rect 29094 1078 29558 1112
rect 30112 1078 30576 1112
rect 31130 1078 31594 1112
rect 32148 1078 32612 1112
rect 33166 1078 33630 1112
rect 1194 558 1658 592
rect 2212 558 2676 592
rect 3230 558 3694 592
rect 4248 558 4712 592
rect 5266 558 5730 592
rect 6284 558 6748 592
rect 7302 558 7766 592
rect 8320 558 8784 592
rect 9338 558 9802 592
rect 10356 558 10820 592
rect 13530 452 13564 1028
rect 14548 452 14582 1028
rect 15566 452 15600 1028
rect 16584 452 16618 1028
rect 17602 452 17636 1028
rect 18620 452 18654 1028
rect 19638 452 19672 1028
rect 20656 452 20690 1028
rect 21674 452 21708 1028
rect 22692 452 22726 1028
rect 23710 452 23744 1028
rect 24728 452 24762 1028
rect 25746 452 25780 1028
rect 26764 452 26798 1028
rect 27782 452 27816 1028
rect 28800 452 28834 1028
rect 29818 452 29852 1028
rect 30836 452 30870 1028
rect 31854 452 31888 1028
rect 32872 452 32906 1028
rect 33890 452 33924 1028
rect -1114 362 -1092 396
rect -1092 362 -934 396
rect -934 362 -914 396
rect 13824 368 14288 402
rect 14842 368 15306 402
rect 15860 368 16324 402
rect 16878 368 17342 402
rect 17896 368 18360 402
rect 18914 368 19378 402
rect 19932 368 20396 402
rect 20950 368 21414 402
rect 21968 368 22432 402
rect 22986 368 23450 402
rect 24004 368 24468 402
rect 25022 368 25486 402
rect 26040 368 26504 402
rect 27058 368 27522 402
rect 28076 368 28540 402
rect 29094 368 29558 402
rect 30112 368 30576 402
rect 31130 368 31594 402
rect 32148 368 32612 402
rect 33166 368 33630 402
rect -1188 223 -1154 360
rect -1030 240 -996 274
rect -1188 51 -1154 223
rect -872 223 -836 358
rect -1074 84 -1040 190
rect -986 84 -952 190
rect -1188 -100 -1154 51
rect -872 51 -838 223
rect -838 51 -836 223
rect -1030 0 -996 34
rect -872 -96 -836 51
rect 35772 40 35872 14300
rect 39728 15092 39790 15192
rect 39790 15092 76710 15192
rect 76710 15092 76772 15192
rect 54826 14372 55290 14406
rect 55844 14372 56308 14406
rect 56862 14372 57326 14406
rect 57880 14372 58344 14406
rect 58898 14372 59362 14406
rect 59916 14372 60380 14406
rect 60934 14372 61398 14406
rect 61952 14372 62416 14406
rect 62970 14372 63434 14406
rect 63988 14372 64452 14406
rect 65006 14372 65470 14406
rect 66024 14372 66488 14406
rect 67042 14372 67506 14406
rect 68060 14372 68524 14406
rect 69078 14372 69542 14406
rect 70096 14372 70560 14406
rect 71114 14372 71578 14406
rect 72132 14372 72596 14406
rect 73150 14372 73614 14406
rect 74168 14372 74632 14406
rect 36818 13870 36880 13970
rect 36880 13870 38520 13970
rect 38520 13870 38582 13970
rect 36718 12593 36818 13803
rect 37014 13045 37098 13079
rect 37272 13045 37356 13079
rect 37530 13045 37614 13079
rect 37788 13045 37872 13079
rect 38046 13045 38130 13079
rect 38304 13045 38388 13079
rect 36910 12810 36944 12986
rect 37168 12810 37202 12986
rect 37426 12810 37460 12986
rect 37684 12810 37718 12986
rect 37942 12810 37976 12986
rect 38200 12810 38234 12986
rect 38458 12810 38492 12986
rect 37014 12717 37098 12751
rect 37272 12717 37356 12751
rect 37530 12717 37614 12751
rect 37788 12717 37872 12751
rect 38046 12717 38130 12751
rect 38304 12717 38388 12751
rect 38582 12593 38682 13803
rect 36818 12426 36880 12526
rect 36880 12426 38520 12526
rect 38520 12426 38582 12526
rect -1116 -136 -1092 -102
rect -1092 -136 -934 -102
rect -934 -136 -916 -102
rect -1272 -852 -1210 -752
rect -1210 -852 35710 -752
rect 35710 -852 35772 -752
rect 39628 40 39728 14300
rect 43060 13896 43524 13930
rect 44078 13896 44542 13930
rect 45096 13896 45560 13930
rect 46114 13896 46578 13930
rect 47132 13896 47596 13930
rect 48150 13896 48614 13930
rect 49168 13896 49632 13930
rect 50186 13896 50650 13930
rect 51204 13896 51668 13930
rect 42766 13270 42800 13846
rect 43784 13270 43818 13846
rect 44802 13270 44836 13846
rect 45820 13270 45854 13846
rect 46838 13270 46872 13846
rect 47856 13270 47890 13846
rect 48874 13270 48908 13846
rect 49892 13270 49926 13846
rect 50910 13270 50944 13846
rect 51928 13270 51962 13846
rect 54532 13746 54566 14322
rect 55550 13746 55584 14322
rect 56568 13746 56602 14322
rect 57586 13746 57620 14322
rect 58604 13746 58638 14322
rect 59622 13746 59656 14322
rect 60640 13746 60674 14322
rect 61658 13746 61692 14322
rect 62676 13746 62710 14322
rect 63694 13746 63728 14322
rect 64712 13746 64746 14322
rect 65730 13746 65764 14322
rect 66748 13746 66782 14322
rect 67766 13746 67800 14322
rect 68784 13746 68818 14322
rect 69802 13746 69836 14322
rect 70820 13746 70854 14322
rect 71838 13746 71872 14322
rect 72856 13746 72890 14322
rect 73874 13746 73908 14322
rect 74892 13746 74926 14322
rect 54826 13662 55290 13696
rect 55844 13662 56308 13696
rect 56862 13662 57326 13696
rect 57880 13662 58344 13696
rect 58898 13662 59362 13696
rect 59916 13662 60380 13696
rect 60934 13662 61398 13696
rect 61952 13662 62416 13696
rect 62970 13662 63434 13696
rect 63988 13662 64452 13696
rect 65006 13662 65470 13696
rect 66024 13662 66488 13696
rect 67042 13662 67506 13696
rect 68060 13662 68524 13696
rect 69078 13662 69542 13696
rect 70096 13662 70560 13696
rect 71114 13662 71578 13696
rect 72132 13662 72596 13696
rect 73150 13662 73614 13696
rect 74168 13662 74632 13696
rect 54826 13554 55290 13588
rect 55844 13554 56308 13588
rect 56862 13554 57326 13588
rect 57880 13554 58344 13588
rect 58898 13554 59362 13588
rect 59916 13554 60380 13588
rect 60934 13554 61398 13588
rect 61952 13554 62416 13588
rect 62970 13554 63434 13588
rect 63988 13554 64452 13588
rect 65006 13554 65470 13588
rect 66024 13554 66488 13588
rect 67042 13554 67506 13588
rect 68060 13554 68524 13588
rect 69078 13554 69542 13588
rect 70096 13554 70560 13588
rect 71114 13554 71578 13588
rect 72132 13554 72596 13588
rect 73150 13554 73614 13588
rect 74168 13554 74632 13588
rect 43060 13186 43524 13220
rect 44078 13186 44542 13220
rect 43060 13078 43524 13112
rect 45096 13186 45560 13220
rect 44078 13078 44542 13112
rect 46114 13186 46578 13220
rect 45096 13078 45560 13112
rect 47132 13186 47596 13220
rect 46114 13078 46578 13112
rect 48150 13186 48614 13220
rect 47132 13078 47596 13112
rect 49168 13186 49632 13220
rect 48150 13078 48614 13112
rect 50186 13186 50650 13220
rect 49168 13078 49632 13112
rect 51204 13186 51668 13220
rect 50186 13078 50650 13112
rect 51204 13078 51668 13112
rect 42766 12452 42800 13028
rect 43784 12452 43818 13028
rect 44802 12452 44836 13028
rect 45820 12452 45854 13028
rect 46838 12452 46872 13028
rect 47856 12452 47890 13028
rect 48874 12452 48908 13028
rect 49892 12452 49926 13028
rect 50910 12452 50944 13028
rect 51928 12452 51962 13028
rect 54532 12928 54566 13504
rect 55550 12928 55584 13504
rect 56568 12928 56602 13504
rect 57586 12928 57620 13504
rect 58604 12928 58638 13504
rect 59622 12928 59656 13504
rect 60640 12928 60674 13504
rect 61658 12928 61692 13504
rect 62676 12928 62710 13504
rect 63694 12928 63728 13504
rect 64712 12928 64746 13504
rect 65730 12928 65764 13504
rect 66748 12928 66782 13504
rect 67766 12928 67800 13504
rect 68784 12928 68818 13504
rect 69802 12928 69836 13504
rect 70820 12928 70854 13504
rect 71838 12928 71872 13504
rect 72856 12928 72890 13504
rect 73874 12928 73908 13504
rect 74892 12928 74926 13504
rect 54826 12844 55290 12878
rect 55844 12844 56308 12878
rect 56862 12844 57326 12878
rect 57880 12844 58344 12878
rect 58898 12844 59362 12878
rect 59916 12844 60380 12878
rect 60934 12844 61398 12878
rect 61952 12844 62416 12878
rect 62970 12844 63434 12878
rect 63988 12844 64452 12878
rect 65006 12844 65470 12878
rect 66024 12844 66488 12878
rect 67042 12844 67506 12878
rect 68060 12844 68524 12878
rect 69078 12844 69542 12878
rect 70096 12844 70560 12878
rect 71114 12844 71578 12878
rect 72132 12844 72596 12878
rect 73150 12844 73614 12878
rect 74168 12844 74632 12878
rect 43060 12368 43524 12402
rect 44078 12368 44542 12402
rect 43060 12260 43524 12294
rect 45096 12368 45560 12402
rect 44078 12260 44542 12294
rect 46114 12368 46578 12402
rect 45096 12260 45560 12294
rect 47132 12368 47596 12402
rect 46114 12260 46578 12294
rect 48150 12368 48614 12402
rect 47132 12260 47596 12294
rect 49168 12368 49632 12402
rect 48150 12260 48614 12294
rect 50186 12368 50650 12402
rect 49168 12260 49632 12294
rect 51204 12368 51668 12402
rect 50186 12260 50650 12294
rect 51204 12260 51668 12294
rect 42766 11634 42800 12210
rect 43784 11634 43818 12210
rect 44802 11634 44836 12210
rect 45820 11634 45854 12210
rect 46838 11634 46872 12210
rect 47856 11634 47890 12210
rect 48874 11634 48908 12210
rect 49892 11634 49926 12210
rect 50910 11634 50944 12210
rect 51928 11634 51962 12210
rect 54826 12176 55290 12210
rect 55844 12176 56308 12210
rect 56862 12176 57326 12210
rect 57880 12176 58344 12210
rect 58898 12176 59362 12210
rect 59916 12176 60380 12210
rect 60934 12176 61398 12210
rect 61952 12176 62416 12210
rect 62970 12176 63434 12210
rect 63988 12176 64452 12210
rect 65006 12176 65470 12210
rect 66024 12176 66488 12210
rect 67042 12176 67506 12210
rect 68060 12176 68524 12210
rect 69078 12176 69542 12210
rect 70096 12176 70560 12210
rect 71114 12176 71578 12210
rect 72132 12176 72596 12210
rect 73150 12176 73614 12210
rect 74168 12176 74632 12210
rect 43060 11550 43524 11584
rect 44078 11550 44542 11584
rect 43060 11442 43524 11476
rect 45096 11550 45560 11584
rect 44078 11442 44542 11476
rect 46114 11550 46578 11584
rect 45096 11442 45560 11476
rect 47132 11550 47596 11584
rect 46114 11442 46578 11476
rect 48150 11550 48614 11584
rect 47132 11442 47596 11476
rect 49168 11550 49632 11584
rect 48150 11442 48614 11476
rect 50186 11550 50650 11584
rect 49168 11442 49632 11476
rect 51204 11550 51668 11584
rect 50186 11442 50650 11476
rect 54532 11550 54566 12126
rect 55550 11550 55584 12126
rect 56568 11550 56602 12126
rect 57586 11550 57620 12126
rect 58604 11550 58638 12126
rect 59622 11550 59656 12126
rect 60640 11550 60674 12126
rect 61658 11550 61692 12126
rect 62676 11550 62710 12126
rect 63694 11550 63728 12126
rect 64712 11550 64746 12126
rect 65730 11550 65764 12126
rect 66748 11550 66782 12126
rect 67766 11550 67800 12126
rect 68784 11550 68818 12126
rect 69802 11550 69836 12126
rect 70820 11550 70854 12126
rect 71838 11550 71872 12126
rect 72856 11550 72890 12126
rect 73874 11550 73908 12126
rect 74892 11550 74926 12126
rect 51204 11442 51668 11476
rect 54826 11466 55290 11500
rect 55844 11466 56308 11500
rect 56862 11466 57326 11500
rect 57880 11466 58344 11500
rect 58898 11466 59362 11500
rect 59916 11466 60380 11500
rect 60934 11466 61398 11500
rect 61952 11466 62416 11500
rect 62970 11466 63434 11500
rect 63988 11466 64452 11500
rect 65006 11466 65470 11500
rect 66024 11466 66488 11500
rect 67042 11466 67506 11500
rect 68060 11466 68524 11500
rect 69078 11466 69542 11500
rect 70096 11466 70560 11500
rect 71114 11466 71578 11500
rect 72132 11466 72596 11500
rect 73150 11466 73614 11500
rect 74168 11466 74632 11500
rect 42766 10816 42800 11392
rect 43784 10816 43818 11392
rect 44802 10816 44836 11392
rect 45820 10816 45854 11392
rect 46838 10816 46872 11392
rect 47856 10816 47890 11392
rect 48874 10816 48908 11392
rect 49892 10816 49926 11392
rect 50910 10816 50944 11392
rect 51928 10816 51962 11392
rect 54826 10944 55290 10978
rect 55844 10944 56308 10978
rect 56862 10944 57326 10978
rect 57880 10944 58344 10978
rect 58898 10944 59362 10978
rect 59916 10944 60380 10978
rect 60934 10944 61398 10978
rect 61952 10944 62416 10978
rect 62970 10944 63434 10978
rect 63988 10944 64452 10978
rect 65006 10944 65470 10978
rect 66024 10944 66488 10978
rect 67042 10944 67506 10978
rect 68060 10944 68524 10978
rect 69078 10944 69542 10978
rect 70096 10944 70560 10978
rect 71114 10944 71578 10978
rect 72132 10944 72596 10978
rect 73150 10944 73614 10978
rect 74168 10944 74632 10978
rect 43060 10732 43524 10766
rect 44078 10732 44542 10766
rect 43060 10624 43524 10658
rect 45096 10732 45560 10766
rect 44078 10624 44542 10658
rect 46114 10732 46578 10766
rect 45096 10624 45560 10658
rect 47132 10732 47596 10766
rect 46114 10624 46578 10658
rect 48150 10732 48614 10766
rect 47132 10624 47596 10658
rect 49168 10732 49632 10766
rect 48150 10624 48614 10658
rect 50186 10732 50650 10766
rect 49168 10624 49632 10658
rect 51204 10732 51668 10766
rect 50186 10624 50650 10658
rect 51204 10624 51668 10658
rect 42766 9998 42800 10574
rect 43784 9998 43818 10574
rect 44802 9998 44836 10574
rect 45820 9998 45854 10574
rect 46838 9998 46872 10574
rect 47856 9998 47890 10574
rect 48874 9998 48908 10574
rect 49892 9998 49926 10574
rect 50910 9998 50944 10574
rect 51928 9998 51962 10574
rect 54532 10318 54566 10894
rect 55550 10318 55584 10894
rect 56568 10318 56602 10894
rect 57586 10318 57620 10894
rect 58604 10318 58638 10894
rect 59622 10318 59656 10894
rect 60640 10318 60674 10894
rect 61658 10318 61692 10894
rect 62676 10318 62710 10894
rect 63694 10318 63728 10894
rect 64712 10318 64746 10894
rect 65730 10318 65764 10894
rect 66748 10318 66782 10894
rect 67766 10318 67800 10894
rect 68784 10318 68818 10894
rect 69802 10318 69836 10894
rect 70820 10318 70854 10894
rect 71838 10318 71872 10894
rect 72856 10318 72890 10894
rect 73874 10318 73908 10894
rect 74892 10318 74926 10894
rect 54826 10234 55290 10268
rect 55844 10234 56308 10268
rect 56862 10234 57326 10268
rect 57880 10234 58344 10268
rect 58898 10234 59362 10268
rect 59916 10234 60380 10268
rect 60934 10234 61398 10268
rect 61952 10234 62416 10268
rect 62970 10234 63434 10268
rect 63988 10234 64452 10268
rect 65006 10234 65470 10268
rect 66024 10234 66488 10268
rect 67042 10234 67506 10268
rect 68060 10234 68524 10268
rect 69078 10234 69542 10268
rect 70096 10234 70560 10268
rect 71114 10234 71578 10268
rect 72132 10234 72596 10268
rect 73150 10234 73614 10268
rect 74168 10234 74632 10268
rect 43060 9914 43524 9948
rect 44078 9914 44542 9948
rect 43060 9806 43524 9840
rect 45096 9914 45560 9948
rect 44078 9806 44542 9840
rect 46114 9914 46578 9948
rect 45096 9806 45560 9840
rect 47132 9914 47596 9948
rect 46114 9806 46578 9840
rect 48150 9914 48614 9948
rect 47132 9806 47596 9840
rect 49168 9914 49632 9948
rect 48150 9806 48614 9840
rect 50186 9914 50650 9948
rect 49168 9806 49632 9840
rect 51204 9914 51668 9948
rect 50186 9806 50650 9840
rect 51204 9806 51668 9840
rect 42766 9180 42800 9756
rect 43784 9180 43818 9756
rect 44802 9180 44836 9756
rect 45820 9180 45854 9756
rect 46838 9180 46872 9756
rect 47856 9180 47890 9756
rect 48874 9180 48908 9756
rect 49892 9180 49926 9756
rect 50910 9180 50944 9756
rect 51928 9180 51962 9756
rect 54824 9710 55288 9744
rect 55842 9710 56306 9744
rect 56860 9710 57324 9744
rect 57878 9710 58342 9744
rect 58896 9710 59360 9744
rect 59914 9710 60378 9744
rect 60932 9710 61396 9744
rect 61950 9710 62414 9744
rect 62968 9710 63432 9744
rect 63986 9710 64450 9744
rect 65004 9710 65468 9744
rect 66022 9710 66486 9744
rect 67040 9710 67504 9744
rect 68058 9710 68522 9744
rect 69076 9710 69540 9744
rect 70094 9710 70558 9744
rect 71112 9710 71576 9744
rect 72130 9710 72594 9744
rect 73148 9710 73612 9744
rect 74166 9710 74630 9744
rect 43060 9096 43524 9130
rect 44078 9096 44542 9130
rect 43060 8988 43524 9022
rect 45096 9096 45560 9130
rect 44078 8988 44542 9022
rect 46114 9096 46578 9130
rect 45096 8988 45560 9022
rect 47132 9096 47596 9130
rect 46114 8988 46578 9022
rect 48150 9096 48614 9130
rect 47132 8988 47596 9022
rect 49168 9096 49632 9130
rect 48150 8988 48614 9022
rect 50186 9096 50650 9130
rect 49168 8988 49632 9022
rect 51204 9096 51668 9130
rect 50186 8988 50650 9022
rect 54530 9084 54564 9660
rect 55548 9084 55582 9660
rect 56566 9084 56600 9660
rect 57584 9084 57618 9660
rect 58602 9084 58636 9660
rect 59620 9084 59654 9660
rect 60638 9084 60672 9660
rect 61656 9084 61690 9660
rect 62674 9084 62708 9660
rect 63692 9084 63726 9660
rect 64710 9084 64744 9660
rect 65728 9084 65762 9660
rect 66746 9084 66780 9660
rect 67764 9084 67798 9660
rect 68782 9084 68816 9660
rect 69800 9084 69834 9660
rect 70818 9084 70852 9660
rect 71836 9084 71870 9660
rect 72854 9084 72888 9660
rect 73872 9084 73906 9660
rect 74890 9084 74924 9660
rect 51204 8988 51668 9022
rect 54824 9000 55288 9034
rect 55842 9000 56306 9034
rect 56860 9000 57324 9034
rect 57878 9000 58342 9034
rect 58896 9000 59360 9034
rect 59914 9000 60378 9034
rect 60932 9000 61396 9034
rect 61950 9000 62414 9034
rect 62968 9000 63432 9034
rect 63986 9000 64450 9034
rect 65004 9000 65468 9034
rect 66022 9000 66486 9034
rect 67040 9000 67504 9034
rect 68058 9000 68522 9034
rect 69076 9000 69540 9034
rect 70094 9000 70558 9034
rect 71112 9000 71576 9034
rect 72130 9000 72594 9034
rect 73148 9000 73612 9034
rect 74166 9000 74630 9034
rect 42766 8362 42800 8938
rect 43784 8362 43818 8938
rect 44802 8362 44836 8938
rect 45820 8362 45854 8938
rect 46838 8362 46872 8938
rect 47856 8362 47890 8938
rect 48874 8362 48908 8938
rect 49892 8362 49926 8938
rect 50910 8362 50944 8938
rect 51928 8362 51962 8938
rect 54824 8476 55288 8510
rect 55842 8476 56306 8510
rect 56860 8476 57324 8510
rect 57878 8476 58342 8510
rect 58896 8476 59360 8510
rect 59914 8476 60378 8510
rect 60932 8476 61396 8510
rect 61950 8476 62414 8510
rect 62968 8476 63432 8510
rect 63986 8476 64450 8510
rect 65004 8476 65468 8510
rect 66022 8476 66486 8510
rect 67040 8476 67504 8510
rect 68058 8476 68522 8510
rect 69076 8476 69540 8510
rect 70094 8476 70558 8510
rect 71112 8476 71576 8510
rect 72130 8476 72594 8510
rect 73148 8476 73612 8510
rect 74166 8476 74630 8510
rect 43060 8278 43524 8312
rect 44078 8278 44542 8312
rect 43060 8170 43524 8204
rect 45096 8278 45560 8312
rect 44078 8170 44542 8204
rect 46114 8278 46578 8312
rect 45096 8170 45560 8204
rect 47132 8278 47596 8312
rect 46114 8170 46578 8204
rect 48150 8278 48614 8312
rect 47132 8170 47596 8204
rect 49168 8278 49632 8312
rect 48150 8170 48614 8204
rect 50186 8278 50650 8312
rect 49168 8170 49632 8204
rect 51204 8278 51668 8312
rect 50186 8170 50650 8204
rect 51204 8170 51668 8204
rect 42766 7544 42800 8120
rect 43784 7544 43818 8120
rect 44802 7544 44836 8120
rect 45820 7544 45854 8120
rect 46838 7544 46872 8120
rect 47856 7544 47890 8120
rect 48874 7544 48908 8120
rect 49892 7544 49926 8120
rect 50910 7544 50944 8120
rect 51928 7544 51962 8120
rect 54530 7850 54564 8426
rect 55548 7850 55582 8426
rect 56566 7850 56600 8426
rect 57584 7850 57618 8426
rect 58602 7850 58636 8426
rect 59620 7850 59654 8426
rect 60638 7850 60672 8426
rect 61656 7850 61690 8426
rect 62674 7850 62708 8426
rect 63692 7850 63726 8426
rect 64710 7850 64744 8426
rect 65728 7850 65762 8426
rect 66746 7850 66780 8426
rect 67764 7850 67798 8426
rect 68782 7850 68816 8426
rect 69800 7850 69834 8426
rect 70818 7850 70852 8426
rect 71836 7850 71870 8426
rect 72854 7850 72888 8426
rect 73872 7850 73906 8426
rect 74890 7850 74924 8426
rect 54824 7766 55288 7800
rect 55842 7766 56306 7800
rect 56860 7766 57324 7800
rect 57878 7766 58342 7800
rect 58896 7766 59360 7800
rect 59914 7766 60378 7800
rect 60932 7766 61396 7800
rect 61950 7766 62414 7800
rect 62968 7766 63432 7800
rect 63986 7766 64450 7800
rect 65004 7766 65468 7800
rect 66022 7766 66486 7800
rect 67040 7766 67504 7800
rect 68058 7766 68522 7800
rect 69076 7766 69540 7800
rect 70094 7766 70558 7800
rect 71112 7766 71576 7800
rect 72130 7766 72594 7800
rect 73148 7766 73612 7800
rect 74166 7766 74630 7800
rect 43060 7460 43524 7494
rect 44078 7460 44542 7494
rect 45096 7460 45560 7494
rect 46114 7460 46578 7494
rect 47132 7460 47596 7494
rect 48150 7460 48614 7494
rect 49168 7460 49632 7494
rect 50186 7460 50650 7494
rect 51204 7460 51668 7494
rect 54824 7244 55288 7278
rect 55842 7244 56306 7278
rect 56860 7244 57324 7278
rect 57878 7244 58342 7278
rect 58896 7244 59360 7278
rect 59914 7244 60378 7278
rect 60932 7244 61396 7278
rect 61950 7244 62414 7278
rect 62968 7244 63432 7278
rect 63986 7244 64450 7278
rect 65004 7244 65468 7278
rect 66022 7244 66486 7278
rect 67040 7244 67504 7278
rect 68058 7244 68522 7278
rect 69076 7244 69540 7278
rect 70094 7244 70558 7278
rect 71112 7244 71576 7278
rect 72130 7244 72594 7278
rect 73148 7244 73612 7278
rect 74166 7244 74630 7278
rect 54530 6618 54564 7194
rect 55548 6618 55582 7194
rect 56566 6618 56600 7194
rect 57584 6618 57618 7194
rect 58602 6618 58636 7194
rect 59620 6618 59654 7194
rect 60638 6618 60672 7194
rect 61656 6618 61690 7194
rect 62674 6618 62708 7194
rect 63692 6618 63726 7194
rect 64710 6618 64744 7194
rect 65728 6618 65762 7194
rect 66746 6618 66780 7194
rect 67764 6618 67798 7194
rect 68782 6618 68816 7194
rect 69800 6618 69834 7194
rect 70818 6618 70852 7194
rect 71836 6618 71870 7194
rect 72854 6618 72888 7194
rect 73872 6618 73906 7194
rect 74890 6618 74924 7194
rect 54824 6534 55288 6568
rect 55842 6534 56306 6568
rect 56860 6534 57324 6568
rect 57878 6534 58342 6568
rect 58896 6534 59360 6568
rect 59914 6534 60378 6568
rect 60932 6534 61396 6568
rect 61950 6534 62414 6568
rect 62968 6534 63432 6568
rect 63986 6534 64450 6568
rect 65004 6534 65468 6568
rect 66022 6534 66486 6568
rect 67040 6534 67504 6568
rect 68058 6534 68522 6568
rect 69076 6534 69540 6568
rect 70094 6534 70558 6568
rect 71112 6534 71576 6568
rect 72130 6534 72594 6568
rect 73148 6534 73612 6568
rect 74166 6534 74630 6568
rect 41736 6146 42200 6180
rect 42754 6146 43218 6180
rect 43772 6146 44236 6180
rect 44790 6146 45254 6180
rect 45808 6146 46272 6180
rect 46826 6146 47290 6180
rect 47844 6146 48308 6180
rect 48862 6146 49326 6180
rect 49880 6146 50344 6180
rect 50898 6146 51362 6180
rect 51916 6146 52380 6180
rect 41442 5520 41476 6096
rect 42460 5520 42494 6096
rect 43478 5520 43512 6096
rect 44496 5520 44530 6096
rect 45514 5520 45548 6096
rect 46532 5520 46566 6096
rect 47550 5520 47584 6096
rect 48568 5520 48602 6096
rect 49586 5520 49620 6096
rect 50604 5520 50638 6096
rect 51622 5520 51656 6096
rect 52640 5520 52674 6096
rect 54824 6010 55288 6044
rect 55842 6010 56306 6044
rect 56860 6010 57324 6044
rect 57878 6010 58342 6044
rect 58896 6010 59360 6044
rect 59914 6010 60378 6044
rect 60932 6010 61396 6044
rect 61950 6010 62414 6044
rect 62968 6010 63432 6044
rect 63986 6010 64450 6044
rect 65004 6010 65468 6044
rect 66022 6010 66486 6044
rect 67040 6010 67504 6044
rect 68058 6010 68522 6044
rect 69076 6010 69540 6044
rect 70094 6010 70558 6044
rect 71112 6010 71576 6044
rect 72130 6010 72594 6044
rect 73148 6010 73612 6044
rect 74166 6010 74630 6044
rect 41736 5436 42200 5470
rect 42754 5436 43218 5470
rect 43772 5436 44236 5470
rect 44790 5436 45254 5470
rect 45808 5436 46272 5470
rect 46826 5436 47290 5470
rect 47844 5436 48308 5470
rect 48862 5436 49326 5470
rect 49880 5436 50344 5470
rect 50898 5436 51362 5470
rect 51916 5436 52380 5470
rect 54530 5384 54564 5960
rect 55548 5384 55582 5960
rect 56566 5384 56600 5960
rect 57584 5384 57618 5960
rect 58602 5384 58636 5960
rect 59620 5384 59654 5960
rect 60638 5384 60672 5960
rect 61656 5384 61690 5960
rect 62674 5384 62708 5960
rect 63692 5384 63726 5960
rect 64710 5384 64744 5960
rect 65728 5384 65762 5960
rect 66746 5384 66780 5960
rect 67764 5384 67798 5960
rect 68782 5384 68816 5960
rect 69800 5384 69834 5960
rect 70818 5384 70852 5960
rect 71836 5384 71870 5960
rect 72854 5384 72888 5960
rect 73872 5384 73906 5960
rect 74890 5384 74924 5960
rect 54824 5300 55288 5334
rect 55842 5300 56306 5334
rect 56860 5300 57324 5334
rect 57878 5300 58342 5334
rect 58896 5300 59360 5334
rect 59914 5300 60378 5334
rect 60932 5300 61396 5334
rect 61950 5300 62414 5334
rect 62968 5300 63432 5334
rect 63986 5300 64450 5334
rect 65004 5300 65468 5334
rect 66022 5300 66486 5334
rect 67040 5300 67504 5334
rect 68058 5300 68522 5334
rect 69076 5300 69540 5334
rect 70094 5300 70558 5334
rect 71112 5300 71576 5334
rect 72130 5300 72594 5334
rect 73148 5300 73612 5334
rect 74166 5300 74630 5334
rect 41736 5034 42200 5068
rect 42754 5034 43218 5068
rect 43772 5034 44236 5068
rect 44790 5034 45254 5068
rect 45808 5034 46272 5068
rect 46826 5034 47290 5068
rect 47844 5034 48308 5068
rect 48862 5034 49326 5068
rect 49880 5034 50344 5068
rect 50898 5034 51362 5068
rect 51916 5034 52380 5068
rect 41442 4408 41476 4984
rect 42460 4408 42494 4984
rect 43478 4408 43512 4984
rect 44496 4408 44530 4984
rect 45514 4408 45548 4984
rect 46532 4408 46566 4984
rect 47550 4408 47584 4984
rect 48568 4408 48602 4984
rect 49586 4408 49620 4984
rect 50604 4408 50638 4984
rect 51622 4408 51656 4984
rect 52640 4408 52674 4984
rect 54824 4776 55288 4810
rect 55842 4776 56306 4810
rect 56860 4776 57324 4810
rect 57878 4776 58342 4810
rect 58896 4776 59360 4810
rect 59914 4776 60378 4810
rect 60932 4776 61396 4810
rect 61950 4776 62414 4810
rect 62968 4776 63432 4810
rect 63986 4776 64450 4810
rect 65004 4776 65468 4810
rect 66022 4776 66486 4810
rect 67040 4776 67504 4810
rect 68058 4776 68522 4810
rect 69076 4776 69540 4810
rect 70094 4776 70558 4810
rect 71112 4776 71576 4810
rect 72130 4776 72594 4810
rect 73148 4776 73612 4810
rect 74166 4776 74630 4810
rect 41736 4324 42200 4358
rect 42754 4324 43218 4358
rect 43772 4324 44236 4358
rect 44790 4324 45254 4358
rect 45808 4324 46272 4358
rect 46826 4324 47290 4358
rect 47844 4324 48308 4358
rect 48862 4324 49326 4358
rect 49880 4324 50344 4358
rect 50898 4324 51362 4358
rect 51916 4324 52380 4358
rect 54530 4150 54564 4726
rect 55548 4150 55582 4726
rect 56566 4150 56600 4726
rect 57584 4150 57618 4726
rect 58602 4150 58636 4726
rect 59620 4150 59654 4726
rect 60638 4150 60672 4726
rect 61656 4150 61690 4726
rect 62674 4150 62708 4726
rect 63692 4150 63726 4726
rect 64710 4150 64744 4726
rect 65728 4150 65762 4726
rect 66746 4150 66780 4726
rect 67764 4150 67798 4726
rect 68782 4150 68816 4726
rect 69800 4150 69834 4726
rect 70818 4150 70852 4726
rect 71836 4150 71870 4726
rect 72854 4150 72888 4726
rect 73872 4150 73906 4726
rect 74890 4150 74924 4726
rect 54824 4066 55288 4100
rect 55842 4066 56306 4100
rect 56860 4066 57324 4100
rect 57878 4066 58342 4100
rect 58896 4066 59360 4100
rect 59914 4066 60378 4100
rect 60932 4066 61396 4100
rect 61950 4066 62414 4100
rect 62968 4066 63432 4100
rect 63986 4066 64450 4100
rect 65004 4066 65468 4100
rect 66022 4066 66486 4100
rect 67040 4066 67504 4100
rect 68058 4066 68522 4100
rect 69076 4066 69540 4100
rect 70094 4066 70558 4100
rect 71112 4066 71576 4100
rect 72130 4066 72594 4100
rect 73148 4066 73612 4100
rect 74166 4066 74630 4100
rect 41736 3922 42200 3956
rect 42754 3922 43218 3956
rect 43772 3922 44236 3956
rect 44790 3922 45254 3956
rect 45808 3922 46272 3956
rect 46826 3922 47290 3956
rect 47844 3922 48308 3956
rect 48862 3922 49326 3956
rect 49880 3922 50344 3956
rect 50898 3922 51362 3956
rect 51916 3922 52380 3956
rect 41442 3296 41476 3872
rect 42460 3296 42494 3872
rect 43478 3296 43512 3872
rect 44496 3296 44530 3872
rect 45514 3296 45548 3872
rect 46532 3296 46566 3872
rect 47550 3296 47584 3872
rect 48568 3296 48602 3872
rect 49586 3296 49620 3872
rect 50604 3296 50638 3872
rect 51622 3296 51656 3872
rect 52640 3296 52674 3872
rect 54824 3544 55288 3578
rect 55842 3544 56306 3578
rect 56860 3544 57324 3578
rect 57878 3544 58342 3578
rect 58896 3544 59360 3578
rect 59914 3544 60378 3578
rect 60932 3544 61396 3578
rect 61950 3544 62414 3578
rect 62968 3544 63432 3578
rect 63986 3544 64450 3578
rect 65004 3544 65468 3578
rect 66022 3544 66486 3578
rect 67040 3544 67504 3578
rect 68058 3544 68522 3578
rect 69076 3544 69540 3578
rect 70094 3544 70558 3578
rect 71112 3544 71576 3578
rect 72130 3544 72594 3578
rect 73148 3544 73612 3578
rect 74166 3544 74630 3578
rect 41736 3212 42200 3246
rect 42754 3212 43218 3246
rect 43772 3212 44236 3246
rect 44790 3212 45254 3246
rect 45808 3212 46272 3246
rect 46826 3212 47290 3246
rect 47844 3212 48308 3246
rect 48862 3212 49326 3246
rect 49880 3212 50344 3246
rect 50898 3212 51362 3246
rect 51916 3212 52380 3246
rect 54530 2918 54564 3494
rect 55548 2918 55582 3494
rect 56566 2918 56600 3494
rect 57584 2918 57618 3494
rect 58602 2918 58636 3494
rect 59620 2918 59654 3494
rect 60638 2918 60672 3494
rect 61656 2918 61690 3494
rect 62674 2918 62708 3494
rect 63692 2918 63726 3494
rect 64710 2918 64744 3494
rect 65728 2918 65762 3494
rect 66746 2918 66780 3494
rect 67764 2918 67798 3494
rect 68782 2918 68816 3494
rect 69800 2918 69834 3494
rect 70818 2918 70852 3494
rect 71836 2918 71870 3494
rect 72854 2918 72888 3494
rect 73872 2918 73906 3494
rect 74890 2918 74924 3494
rect 41736 2810 42200 2844
rect 42754 2810 43218 2844
rect 43772 2810 44236 2844
rect 44790 2810 45254 2844
rect 45808 2810 46272 2844
rect 46826 2810 47290 2844
rect 47844 2810 48308 2844
rect 48862 2810 49326 2844
rect 49880 2810 50344 2844
rect 50898 2810 51362 2844
rect 51916 2810 52380 2844
rect 54824 2834 55288 2868
rect 55842 2834 56306 2868
rect 56860 2834 57324 2868
rect 57878 2834 58342 2868
rect 58896 2834 59360 2868
rect 59914 2834 60378 2868
rect 60932 2834 61396 2868
rect 61950 2834 62414 2868
rect 62968 2834 63432 2868
rect 63986 2834 64450 2868
rect 65004 2834 65468 2868
rect 66022 2834 66486 2868
rect 67040 2834 67504 2868
rect 68058 2834 68522 2868
rect 69076 2834 69540 2868
rect 70094 2834 70558 2868
rect 71112 2834 71576 2868
rect 72130 2834 72594 2868
rect 73148 2834 73612 2868
rect 74166 2834 74630 2868
rect 41442 2184 41476 2760
rect 42460 2184 42494 2760
rect 43478 2184 43512 2760
rect 44496 2184 44530 2760
rect 45514 2184 45548 2760
rect 46532 2184 46566 2760
rect 47550 2184 47584 2760
rect 48568 2184 48602 2760
rect 49586 2184 49620 2760
rect 50604 2184 50638 2760
rect 51622 2184 51656 2760
rect 52640 2184 52674 2760
rect 54824 2310 55288 2344
rect 55842 2310 56306 2344
rect 56860 2310 57324 2344
rect 57878 2310 58342 2344
rect 58896 2310 59360 2344
rect 59914 2310 60378 2344
rect 60932 2310 61396 2344
rect 61950 2310 62414 2344
rect 62968 2310 63432 2344
rect 63986 2310 64450 2344
rect 65004 2310 65468 2344
rect 66022 2310 66486 2344
rect 67040 2310 67504 2344
rect 68058 2310 68522 2344
rect 69076 2310 69540 2344
rect 70094 2310 70558 2344
rect 71112 2310 71576 2344
rect 72130 2310 72594 2344
rect 73148 2310 73612 2344
rect 74166 2310 74630 2344
rect 41736 2100 42200 2134
rect 42754 2100 43218 2134
rect 43772 2100 44236 2134
rect 44790 2100 45254 2134
rect 45808 2100 46272 2134
rect 46826 2100 47290 2134
rect 47844 2100 48308 2134
rect 48862 2100 49326 2134
rect 49880 2100 50344 2134
rect 50898 2100 51362 2134
rect 51916 2100 52380 2134
rect 54530 1684 54564 2260
rect 55548 1684 55582 2260
rect 56566 1684 56600 2260
rect 57584 1684 57618 2260
rect 58602 1684 58636 2260
rect 59620 1684 59654 2260
rect 60638 1684 60672 2260
rect 61656 1684 61690 2260
rect 62674 1684 62708 2260
rect 63692 1684 63726 2260
rect 64710 1684 64744 2260
rect 65728 1684 65762 2260
rect 66746 1684 66780 2260
rect 67764 1684 67798 2260
rect 68782 1684 68816 2260
rect 69800 1684 69834 2260
rect 70818 1684 70852 2260
rect 71836 1684 71870 2260
rect 72854 1684 72888 2260
rect 73872 1684 73906 2260
rect 74890 1684 74924 2260
rect 54824 1600 55288 1634
rect 55842 1600 56306 1634
rect 56860 1600 57324 1634
rect 57878 1600 58342 1634
rect 58896 1600 59360 1634
rect 59914 1600 60378 1634
rect 60932 1600 61396 1634
rect 61950 1600 62414 1634
rect 62968 1600 63432 1634
rect 63986 1600 64450 1634
rect 65004 1600 65468 1634
rect 66022 1600 66486 1634
rect 67040 1600 67504 1634
rect 68058 1600 68522 1634
rect 69076 1600 69540 1634
rect 70094 1600 70558 1634
rect 71112 1600 71576 1634
rect 72130 1600 72594 1634
rect 73148 1600 73612 1634
rect 74166 1600 74630 1634
rect 42194 1268 42658 1302
rect 43212 1268 43676 1302
rect 44230 1268 44694 1302
rect 45248 1268 45712 1302
rect 46266 1268 46730 1302
rect 47284 1268 47748 1302
rect 48302 1268 48766 1302
rect 49320 1268 49784 1302
rect 50338 1268 50802 1302
rect 51356 1268 51820 1302
rect 41900 642 41934 1218
rect 42918 642 42952 1218
rect 43936 642 43970 1218
rect 44954 642 44988 1218
rect 45972 642 46006 1218
rect 46990 642 47024 1218
rect 48008 642 48042 1218
rect 49026 642 49060 1218
rect 50044 642 50078 1218
rect 51062 642 51096 1218
rect 52080 642 52114 1218
rect 54824 1078 55288 1112
rect 55842 1078 56306 1112
rect 56860 1078 57324 1112
rect 57878 1078 58342 1112
rect 58896 1078 59360 1112
rect 59914 1078 60378 1112
rect 60932 1078 61396 1112
rect 61950 1078 62414 1112
rect 62968 1078 63432 1112
rect 63986 1078 64450 1112
rect 65004 1078 65468 1112
rect 66022 1078 66486 1112
rect 67040 1078 67504 1112
rect 68058 1078 68522 1112
rect 69076 1078 69540 1112
rect 70094 1078 70558 1112
rect 71112 1078 71576 1112
rect 72130 1078 72594 1112
rect 73148 1078 73612 1112
rect 74166 1078 74630 1112
rect 42194 558 42658 592
rect 43212 558 43676 592
rect 44230 558 44694 592
rect 45248 558 45712 592
rect 46266 558 46730 592
rect 47284 558 47748 592
rect 48302 558 48766 592
rect 49320 558 49784 592
rect 50338 558 50802 592
rect 51356 558 51820 592
rect 54530 452 54564 1028
rect 55548 452 55582 1028
rect 56566 452 56600 1028
rect 57584 452 57618 1028
rect 58602 452 58636 1028
rect 59620 452 59654 1028
rect 60638 452 60672 1028
rect 61656 452 61690 1028
rect 62674 452 62708 1028
rect 63692 452 63726 1028
rect 64710 452 64744 1028
rect 65728 452 65762 1028
rect 66746 452 66780 1028
rect 67764 452 67798 1028
rect 68782 452 68816 1028
rect 69800 452 69834 1028
rect 70818 452 70852 1028
rect 71836 452 71870 1028
rect 72854 452 72888 1028
rect 73872 452 73906 1028
rect 74890 452 74924 1028
rect 54824 368 55288 402
rect 55842 368 56306 402
rect 56860 368 57324 402
rect 57878 368 58342 402
rect 58896 368 59360 402
rect 59914 368 60378 402
rect 60932 368 61396 402
rect 61950 368 62414 402
rect 62968 368 63432 402
rect 63986 368 64450 402
rect 65004 368 65468 402
rect 66022 368 66486 402
rect 67040 368 67504 402
rect 68058 368 68522 402
rect 69076 368 69540 402
rect 70094 368 70558 402
rect 71112 368 71576 402
rect 72130 368 72594 402
rect 73148 368 73612 402
rect 74166 368 74630 402
rect 76772 40 76872 14300
rect 39728 -852 39790 -752
rect 39790 -852 76710 -752
rect 76710 -852 76772 -752
<< metal1 >>
rect 11322 30692 35778 30698
rect 11322 30592 11428 30692
rect 35672 30592 35778 30692
rect 11322 30586 35778 30592
rect 11322 30072 11434 30586
rect 12034 30286 12044 30586
rect 35056 30286 35066 30586
rect 11322 16642 11328 30072
rect 11428 16642 11434 30072
rect 14948 30204 31828 30236
rect 14948 29990 15011 30204
rect 31796 29990 31828 30204
rect 14948 29968 14998 29990
rect 15058 29968 15434 29990
rect 15494 29968 15872 29990
rect 15932 29968 16306 29990
rect 16366 29970 31828 29990
rect 35666 30072 35778 30586
rect 16366 29968 19302 29970
rect 19462 28494 19522 29970
rect 21498 28494 21558 29970
rect 22002 28494 22062 29970
rect 22510 28494 22570 29970
rect 23022 28494 23082 29970
rect 23536 28494 23596 29970
rect 25568 28494 25628 29970
rect 27608 28494 27668 29970
rect 28098 28494 28158 29970
rect 28618 28494 28678 29970
rect 29126 28494 29186 29970
rect 29640 28494 29700 29970
rect 31676 28494 31736 29970
rect 19462 28434 31736 28494
rect 18930 28228 18936 28288
rect 18996 28228 19002 28288
rect 17424 28012 18502 28072
rect 17424 27832 17484 28012
rect 17928 27931 17988 28012
rect 17720 27925 18208 27931
rect 17720 27891 17732 27925
rect 18196 27891 18208 27925
rect 17720 27885 18208 27891
rect 17424 27792 17438 27832
rect 17432 27256 17438 27792
rect 17472 27792 17484 27832
rect 18442 27832 18502 28012
rect 18936 27931 18996 28228
rect 19462 28042 19522 28434
rect 20012 28228 20018 28288
rect 20078 28228 20084 28288
rect 20970 28228 20976 28288
rect 21036 28228 21042 28288
rect 19456 27982 19462 28042
rect 19522 27982 19528 28042
rect 18738 27925 19226 27931
rect 18738 27891 18750 27925
rect 19214 27891 19226 27925
rect 18738 27885 19226 27891
rect 18442 27806 18456 27832
rect 17472 27256 17478 27792
rect 18450 27292 18456 27806
rect 17432 27244 17478 27256
rect 18444 27256 18456 27292
rect 18490 27806 18502 27832
rect 19462 27832 19522 27982
rect 20018 27931 20078 28228
rect 20976 27931 21036 28228
rect 21498 28042 21558 28434
rect 21492 27982 21498 28042
rect 21558 27982 21564 28042
rect 19756 27925 20244 27931
rect 19756 27891 19768 27925
rect 20232 27891 20244 27925
rect 19756 27885 20244 27891
rect 20774 27925 21262 27931
rect 20774 27891 20786 27925
rect 21250 27891 21262 27925
rect 20774 27885 21262 27891
rect 20976 27882 21036 27885
rect 19462 27808 19474 27832
rect 18490 27292 18496 27806
rect 19468 27296 19474 27808
rect 18490 27256 18504 27292
rect 17720 27197 18208 27203
rect 17720 27163 17732 27197
rect 18196 27163 18208 27197
rect 17720 27157 18208 27163
rect 18444 27110 18504 27256
rect 19464 27256 19474 27296
rect 19508 27808 19522 27832
rect 20486 27832 20532 27844
rect 19508 27296 19514 27808
rect 19508 27256 19524 27296
rect 20486 27284 20492 27832
rect 18948 27203 19008 27204
rect 18738 27197 19226 27203
rect 18738 27163 18750 27197
rect 19214 27163 19226 27197
rect 18738 27157 19226 27163
rect 17274 27050 17280 27110
rect 17340 27050 17346 27110
rect 18438 27050 18444 27110
rect 18504 27050 18510 27110
rect 17144 26846 17150 26906
rect 17210 26846 17216 26906
rect 15136 24662 15142 24722
rect 15202 24662 15208 24722
rect 12964 21346 14186 21406
rect 12964 19430 13024 21346
rect 13106 21182 13166 21346
rect 13618 21281 13678 21346
rect 13402 21275 13890 21281
rect 13402 21241 13414 21275
rect 13878 21241 13890 21275
rect 13402 21235 13890 21241
rect 13106 21132 13120 21182
rect 13114 20606 13120 21132
rect 13154 21132 13166 21182
rect 14126 21182 14186 21346
rect 14420 21275 14908 21281
rect 14420 21241 14432 21275
rect 14896 21241 14908 21275
rect 14420 21235 14908 21241
rect 13154 20606 13160 21132
rect 14126 21130 14138 21182
rect 13114 20594 13160 20606
rect 14132 20606 14138 21130
rect 14172 21130 14186 21182
rect 15142 21182 15202 24662
rect 17150 24290 17210 26846
rect 17280 24436 17340 27050
rect 18438 26846 18444 26906
rect 18504 26846 18510 26906
rect 17720 26789 18208 26795
rect 17720 26755 17732 26789
rect 18196 26755 18208 26789
rect 17720 26749 18208 26755
rect 17432 26696 17478 26708
rect 17432 26156 17438 26696
rect 17426 26120 17438 26156
rect 17472 26156 17478 26696
rect 18444 26696 18504 26846
rect 18948 26795 19008 27157
rect 18738 26789 19226 26795
rect 18738 26755 18750 26789
rect 19214 26755 19226 26789
rect 18738 26749 19226 26755
rect 18948 26746 19008 26749
rect 18444 26658 18456 26696
rect 17472 26120 17486 26156
rect 18450 26150 18456 26658
rect 17426 25970 17486 26120
rect 18444 26120 18456 26150
rect 18490 26658 18504 26696
rect 19464 26696 19524 27256
rect 20480 27256 20492 27284
rect 20526 27284 20532 27832
rect 21498 27832 21558 27982
rect 22002 27931 22062 28434
rect 21792 27925 22280 27931
rect 21792 27891 21804 27925
rect 22268 27891 22280 27925
rect 21792 27885 22280 27891
rect 21498 27808 21510 27832
rect 21504 27314 21510 27808
rect 20526 27256 20540 27284
rect 19756 27197 20244 27203
rect 19756 27163 19768 27197
rect 20232 27163 20244 27197
rect 19756 27157 20244 27163
rect 20480 27006 20540 27256
rect 21488 27256 21510 27314
rect 21544 27808 21558 27832
rect 22510 27832 22570 28434
rect 23022 27931 23082 28434
rect 23536 28044 23596 28434
rect 24034 28228 24040 28288
rect 24100 28228 24106 28288
rect 25052 28228 25058 28288
rect 25118 28228 25124 28288
rect 23530 27984 23536 28044
rect 23596 27984 23602 28044
rect 22810 27925 23298 27931
rect 22810 27891 22822 27925
rect 23286 27891 23298 27925
rect 22810 27885 23298 27891
rect 21544 27314 21550 27808
rect 22510 27762 22528 27832
rect 21544 27256 21552 27314
rect 20774 27197 21262 27203
rect 20774 27163 20786 27197
rect 21250 27163 21262 27197
rect 20774 27157 21262 27163
rect 20474 26946 20480 27006
rect 20540 26946 20546 27006
rect 19756 26789 20244 26795
rect 19756 26755 19768 26789
rect 20232 26755 20244 26789
rect 19756 26749 20244 26755
rect 20774 26789 21262 26795
rect 20774 26755 20786 26789
rect 21250 26755 21262 26789
rect 20774 26749 21262 26755
rect 18490 26150 18496 26658
rect 19464 26656 19474 26696
rect 18490 26120 18504 26150
rect 19468 26146 19474 26656
rect 17720 26061 18208 26067
rect 17720 26027 17732 26061
rect 18196 26027 18208 26061
rect 17720 26021 18208 26027
rect 17938 25970 17998 26021
rect 18444 25970 18504 26120
rect 19460 26120 19474 26146
rect 19508 26656 19524 26696
rect 20486 26696 20532 26708
rect 19508 26146 19514 26656
rect 19508 26120 19520 26146
rect 20486 26140 20492 26696
rect 18930 26067 18990 26074
rect 18738 26061 19226 26067
rect 18738 26027 18750 26061
rect 19214 26027 19226 26061
rect 18738 26021 19226 26027
rect 17426 25910 18504 25970
rect 18438 25766 18498 25768
rect 17428 25706 18498 25766
rect 17428 25560 17488 25706
rect 17938 25659 17998 25706
rect 17720 25653 18208 25659
rect 17720 25619 17732 25653
rect 18196 25619 18208 25653
rect 17720 25613 18208 25619
rect 17428 25528 17438 25560
rect 17432 24984 17438 25528
rect 17472 25528 17488 25560
rect 18438 25560 18498 25706
rect 18930 25756 18990 26021
rect 18930 25659 18990 25696
rect 19460 25974 19520 26120
rect 20478 26120 20492 26140
rect 20526 26140 20532 26696
rect 21488 26696 21552 27256
rect 22522 27256 22528 27762
rect 22562 27762 22570 27832
rect 23536 27832 23596 27984
rect 24040 27931 24100 28228
rect 25058 27931 25118 28228
rect 25568 28044 25628 28434
rect 26076 28228 26082 28288
rect 26142 28228 26148 28288
rect 27088 28228 27094 28288
rect 27154 28228 27160 28288
rect 25560 27984 25566 28044
rect 25626 27984 25632 28044
rect 23828 27925 24316 27931
rect 23828 27891 23840 27925
rect 24304 27891 24316 27925
rect 23828 27885 24316 27891
rect 24846 27925 25334 27931
rect 24846 27891 24858 27925
rect 25322 27891 25334 27925
rect 24846 27885 25334 27891
rect 23536 27792 23546 27832
rect 22562 27256 22568 27762
rect 23540 27310 23546 27792
rect 22522 27244 22568 27256
rect 23524 27256 23546 27310
rect 23580 27792 23596 27832
rect 24558 27832 24604 27844
rect 23580 27310 23586 27792
rect 23580 27256 23588 27310
rect 24558 27296 24564 27832
rect 21792 27197 22280 27203
rect 21792 27163 21804 27197
rect 22268 27163 22280 27197
rect 21792 27157 22280 27163
rect 22810 27197 23298 27203
rect 22810 27163 22822 27197
rect 23286 27163 23298 27197
rect 22810 27157 23298 27163
rect 22510 26946 22516 27006
rect 22576 26946 22582 27006
rect 21792 26789 22280 26795
rect 21792 26755 21804 26789
rect 22268 26755 22280 26789
rect 21792 26749 22280 26755
rect 21488 26666 21510 26696
rect 21504 26148 21510 26666
rect 20526 26120 20538 26140
rect 19958 26067 20018 26068
rect 19756 26061 20244 26067
rect 19756 26027 19768 26061
rect 20232 26027 20244 26061
rect 19756 26021 20244 26027
rect 19958 25974 20018 26021
rect 20478 25974 20538 26120
rect 21496 26120 21510 26148
rect 21544 26666 21552 26696
rect 22516 26696 22576 26946
rect 22810 26789 23298 26795
rect 22810 26755 22822 26789
rect 23286 26755 23298 26789
rect 22810 26749 23298 26755
rect 21544 26148 21550 26666
rect 22516 26658 22528 26696
rect 22522 26156 22528 26658
rect 21544 26146 21556 26148
rect 21544 26120 21560 26146
rect 20986 26067 21046 26072
rect 20774 26061 21262 26067
rect 20774 26027 20786 26061
rect 21250 26027 21262 26061
rect 20774 26021 21262 26027
rect 20986 25974 21046 26021
rect 19460 25972 21046 25974
rect 21496 25972 21560 26120
rect 22514 26120 22528 26156
rect 22562 26658 22576 26696
rect 23524 26696 23588 27256
rect 24554 27256 24564 27296
rect 24598 27296 24604 27832
rect 25568 27832 25628 27984
rect 26082 27931 26142 28228
rect 27094 27931 27154 28228
rect 27608 28046 27668 28434
rect 27602 27986 27608 28046
rect 27668 27986 27674 28046
rect 25864 27925 26352 27931
rect 25864 27891 25876 27925
rect 26340 27891 26352 27925
rect 25864 27885 26352 27891
rect 26882 27925 27370 27931
rect 26882 27891 26894 27925
rect 27358 27891 27370 27925
rect 26882 27885 27370 27891
rect 25568 27792 25582 27832
rect 25576 27312 25582 27792
rect 24598 27256 24614 27296
rect 24042 27203 24102 27206
rect 23828 27197 24316 27203
rect 23828 27163 23840 27197
rect 24304 27163 24316 27197
rect 23828 27157 24316 27163
rect 24042 26795 24102 27157
rect 24554 27110 24614 27256
rect 25566 27256 25582 27312
rect 25616 27792 25628 27832
rect 26594 27832 26640 27844
rect 25616 27312 25622 27792
rect 25616 27256 25630 27312
rect 26594 27294 26600 27832
rect 25060 27203 25120 27212
rect 24846 27197 25334 27203
rect 24846 27163 24858 27197
rect 25322 27163 25334 27197
rect 24846 27157 25334 27163
rect 24548 27050 24554 27110
rect 24614 27050 24620 27110
rect 24544 26846 24550 26906
rect 24610 26846 24616 26906
rect 23828 26789 24316 26795
rect 23828 26755 23840 26789
rect 24304 26755 24316 26789
rect 23828 26749 24316 26755
rect 24042 26748 24102 26749
rect 23524 26662 23546 26696
rect 22562 26156 22568 26658
rect 23540 26156 23546 26662
rect 22562 26120 22578 26156
rect 21792 26061 22280 26067
rect 21792 26027 21804 26061
rect 22268 26027 22280 26061
rect 21792 26021 22280 26027
rect 19460 25914 20986 25972
rect 18738 25653 19226 25659
rect 18738 25619 18750 25653
rect 19214 25619 19226 25653
rect 18738 25613 19226 25619
rect 18438 25528 18456 25560
rect 17472 24984 17478 25528
rect 18450 25026 18456 25528
rect 17432 24972 17478 24984
rect 18438 24984 18456 25026
rect 18490 25528 18498 25560
rect 19460 25560 19520 25914
rect 21490 25912 21496 25972
rect 21556 25912 21562 25972
rect 20986 25906 21046 25912
rect 20472 25810 20478 25874
rect 20542 25810 20548 25874
rect 19962 25696 19968 25756
rect 20028 25696 20034 25756
rect 20478 25716 20542 25810
rect 19968 25659 20028 25696
rect 19756 25653 20244 25659
rect 19756 25619 19768 25653
rect 20232 25619 20244 25653
rect 19756 25613 20244 25619
rect 18490 25026 18496 25528
rect 19460 25508 19474 25560
rect 18490 24984 18502 25026
rect 19468 25020 19474 25508
rect 17720 24925 18208 24931
rect 17720 24891 17732 24925
rect 18196 24891 18208 24925
rect 17720 24885 18208 24891
rect 18438 24776 18502 24984
rect 19460 24984 19474 25020
rect 19508 25508 19520 25560
rect 20478 25560 20544 25716
rect 20974 25696 20980 25756
rect 21040 25696 21046 25756
rect 20980 25659 21040 25696
rect 20774 25653 21262 25659
rect 20774 25619 20786 25653
rect 21250 25619 21262 25653
rect 20774 25613 21262 25619
rect 20980 25612 21040 25613
rect 20478 25510 20492 25560
rect 19508 25020 19514 25508
rect 19508 24984 19520 25020
rect 20486 25008 20492 25510
rect 18738 24925 19226 24931
rect 18738 24891 18750 24925
rect 19214 24891 19226 24925
rect 18738 24885 19226 24891
rect 17994 24716 18502 24776
rect 17274 24376 17280 24436
rect 17340 24376 17346 24436
rect 17150 24230 17570 24290
rect 17510 21418 17570 24230
rect 17630 21968 17636 22028
rect 17696 21968 17702 22028
rect 16160 21350 17370 21410
rect 17504 21358 17510 21418
rect 17570 21358 17576 21418
rect 15438 21275 15926 21281
rect 15438 21241 15450 21275
rect 15914 21241 15926 21275
rect 15438 21235 15926 21241
rect 14172 20606 14178 21130
rect 14132 20594 14178 20606
rect 15142 20606 15156 21182
rect 15190 20606 15202 21182
rect 16160 21182 16220 21350
rect 16672 21281 16732 21350
rect 16456 21275 16944 21281
rect 16456 21241 16468 21275
rect 16932 21241 16944 21275
rect 16456 21235 16944 21241
rect 16160 21134 16174 21182
rect 13402 20547 13890 20553
rect 13402 20513 13414 20547
rect 13878 20513 13890 20547
rect 13402 20507 13890 20513
rect 14420 20547 14908 20553
rect 14420 20513 14432 20547
rect 14896 20513 14908 20547
rect 14420 20507 14908 20513
rect 14626 20464 14686 20507
rect 14620 20404 14626 20464
rect 14686 20404 14692 20464
rect 14728 20292 14734 20352
rect 14794 20292 14800 20352
rect 14734 20249 14794 20292
rect 13402 20243 13890 20249
rect 13402 20209 13414 20243
rect 13878 20209 13890 20243
rect 13402 20203 13890 20209
rect 14420 20243 14908 20249
rect 14420 20209 14432 20243
rect 14896 20209 14908 20243
rect 14420 20203 14908 20209
rect 13114 20150 13160 20162
rect 13114 19632 13120 20150
rect 13104 19574 13120 19632
rect 13154 19632 13160 20150
rect 14132 20150 14178 20162
rect 13154 19574 13164 19632
rect 14132 19624 14138 20150
rect 12958 19370 12964 19430
rect 13024 19370 13030 19430
rect 12838 18342 12898 18348
rect 12964 18342 13024 19370
rect 13104 19320 13164 19574
rect 14124 19574 14138 19624
rect 14172 19624 14178 20150
rect 15142 20150 15202 20606
rect 16168 20606 16174 21134
rect 16208 21134 16220 21182
rect 17178 21182 17238 21350
rect 17178 21136 17192 21182
rect 16208 20606 16214 21134
rect 16168 20594 16214 20606
rect 17186 20606 17192 21136
rect 17226 21136 17238 21182
rect 17226 20606 17232 21136
rect 17186 20594 17232 20606
rect 15438 20547 15926 20553
rect 15438 20513 15450 20547
rect 15914 20513 15926 20547
rect 15438 20507 15926 20513
rect 16456 20547 16944 20553
rect 16456 20513 16468 20547
rect 16932 20513 16944 20547
rect 16456 20507 16944 20513
rect 15518 20352 15578 20507
rect 15642 20404 15648 20464
rect 15708 20404 15714 20464
rect 15512 20292 15518 20352
rect 15578 20292 15584 20352
rect 15648 20249 15708 20404
rect 15438 20243 15926 20249
rect 15438 20209 15450 20243
rect 15914 20209 15926 20243
rect 15438 20203 15926 20209
rect 16456 20243 16944 20249
rect 16456 20209 16468 20243
rect 16932 20209 16944 20243
rect 16456 20203 16944 20209
rect 14172 19574 14184 19624
rect 13402 19515 13890 19521
rect 13402 19481 13414 19515
rect 13878 19481 13890 19515
rect 13402 19475 13890 19481
rect 13606 19320 13666 19475
rect 14124 19320 14184 19574
rect 15142 19574 15156 20150
rect 15190 19574 15202 20150
rect 16168 20150 16214 20162
rect 16168 19660 16174 20150
rect 14420 19515 14908 19521
rect 14420 19481 14432 19515
rect 14896 19481 14908 19515
rect 14420 19475 14908 19481
rect 13104 19260 14124 19320
rect 14184 19260 14190 19320
rect 13104 19118 13164 19260
rect 13606 19217 13666 19260
rect 13402 19211 13890 19217
rect 13402 19177 13414 19211
rect 13878 19177 13890 19211
rect 13402 19171 13890 19177
rect 13104 19058 13120 19118
rect 13114 18542 13120 19058
rect 13154 19058 13164 19118
rect 14124 19118 14184 19260
rect 14634 19217 14694 19475
rect 14420 19211 14908 19217
rect 14420 19177 14432 19211
rect 14896 19177 14908 19211
rect 14420 19171 14908 19177
rect 13154 18542 13160 19058
rect 14124 19054 14138 19118
rect 13114 18530 13160 18542
rect 14132 18542 14138 19054
rect 14172 19054 14184 19118
rect 15142 19118 15202 19574
rect 16158 19574 16174 19660
rect 16208 19660 16214 20150
rect 17186 20150 17232 20162
rect 16208 19574 16218 19660
rect 17186 19620 17192 20150
rect 15438 19515 15926 19521
rect 15438 19481 15450 19515
rect 15914 19481 15926 19515
rect 15438 19475 15926 19481
rect 15652 19217 15712 19475
rect 16158 19430 16218 19574
rect 17178 19574 17192 19620
rect 17226 19620 17232 20150
rect 17226 19574 17238 19620
rect 16456 19515 16944 19521
rect 16456 19481 16468 19515
rect 16932 19481 16944 19515
rect 16456 19475 16944 19481
rect 16672 19430 16732 19475
rect 17178 19430 17238 19574
rect 16152 19370 16158 19430
rect 16218 19370 17238 19430
rect 15438 19211 15926 19217
rect 15438 19177 15450 19211
rect 15914 19177 15926 19211
rect 15438 19171 15926 19177
rect 14172 18542 14178 19054
rect 14132 18530 14178 18542
rect 15142 18542 15156 19118
rect 15190 18542 15202 19118
rect 16158 19118 16218 19370
rect 16672 19217 16732 19370
rect 16456 19211 16944 19217
rect 16456 19177 16468 19211
rect 16932 19177 16944 19211
rect 16456 19171 16944 19177
rect 16158 19062 16174 19118
rect 13402 18483 13890 18489
rect 13402 18449 13414 18483
rect 13878 18449 13890 18483
rect 13402 18443 13890 18449
rect 14420 18483 14908 18489
rect 14420 18449 14432 18483
rect 14896 18449 14908 18483
rect 14420 18443 14908 18449
rect 14640 18396 14700 18443
rect 12898 18282 14188 18342
rect 14634 18336 14640 18396
rect 14700 18336 14706 18396
rect 12838 18276 12898 18282
rect 13102 18086 13162 18282
rect 13610 18185 13670 18282
rect 13402 18179 13890 18185
rect 13402 18145 13414 18179
rect 13878 18145 13890 18179
rect 13402 18139 13890 18145
rect 13102 18034 13120 18086
rect 13114 17510 13120 18034
rect 13154 18034 13162 18086
rect 14128 18086 14188 18282
rect 14740 18236 14746 18296
rect 14806 18236 14812 18296
rect 14746 18185 14806 18236
rect 14420 18179 14908 18185
rect 14420 18145 14432 18179
rect 14896 18145 14908 18179
rect 14420 18139 14908 18145
rect 14128 18038 14138 18086
rect 13154 17510 13160 18034
rect 13114 17498 13160 17510
rect 14132 17510 14138 18038
rect 14172 18038 14188 18086
rect 15142 18086 15202 18542
rect 16168 18542 16174 19062
rect 16208 19062 16218 19118
rect 17178 19118 17238 19370
rect 17310 19320 17370 21350
rect 17304 19260 17310 19320
rect 17370 19260 17376 19320
rect 17178 19082 17192 19118
rect 16208 18542 16214 19062
rect 16168 18530 16214 18542
rect 17186 18542 17192 19082
rect 17226 19082 17238 19118
rect 17226 18542 17232 19082
rect 17186 18530 17232 18542
rect 15438 18483 15926 18489
rect 15438 18449 15450 18483
rect 15914 18449 15926 18483
rect 15438 18443 15926 18449
rect 16456 18483 16944 18489
rect 16456 18449 16468 18483
rect 16932 18449 16944 18483
rect 16456 18443 16944 18449
rect 15532 18296 15592 18443
rect 15644 18336 15650 18396
rect 15710 18336 15716 18396
rect 17310 18342 17370 19260
rect 17496 19132 17502 19192
rect 17562 19132 17568 19192
rect 15526 18236 15532 18296
rect 15592 18236 15598 18296
rect 15650 18185 15710 18336
rect 16158 18282 17370 18342
rect 15438 18179 15926 18185
rect 15438 18145 15450 18179
rect 15914 18145 15926 18179
rect 15438 18139 15926 18145
rect 14172 17510 14178 18038
rect 15142 18012 15156 18086
rect 14132 17498 14178 17510
rect 15150 17510 15156 18012
rect 15190 18012 15202 18086
rect 16158 18086 16218 18282
rect 16660 18185 16720 18282
rect 16456 18179 16944 18185
rect 16456 18145 16468 18179
rect 16932 18145 16944 18179
rect 16456 18139 16944 18145
rect 16158 18056 16174 18086
rect 15190 17510 15196 18012
rect 16168 17592 16174 18056
rect 15150 17498 15196 17510
rect 16160 17510 16174 17592
rect 16208 18056 16218 18086
rect 17178 18086 17238 18282
rect 16208 17592 16214 18056
rect 17178 18018 17192 18086
rect 16208 17510 16220 17592
rect 15638 17457 15698 17461
rect 13402 17451 13890 17457
rect 13402 17417 13414 17451
rect 13878 17417 13890 17451
rect 13402 17411 13890 17417
rect 14420 17451 14908 17457
rect 14420 17417 14432 17451
rect 14896 17417 14908 17451
rect 14420 17411 14908 17417
rect 15438 17451 15926 17457
rect 15438 17417 15450 17451
rect 15914 17417 15926 17451
rect 15438 17411 15926 17417
rect 12352 17286 12412 17292
rect 14632 17286 14692 17411
rect 12412 17226 14692 17286
rect 12352 17220 12412 17226
rect 12492 17110 12552 17116
rect 15638 17112 15698 17411
rect 12552 17050 13286 17110
rect 13346 17052 15638 17110
rect 13346 17050 15698 17052
rect 12492 17044 12552 17050
rect 15638 17046 15698 17050
rect 13392 16936 13452 16942
rect 16160 16936 16220 17510
rect 17186 17510 17192 18018
rect 17226 18018 17238 18086
rect 17226 17510 17232 18018
rect 17186 17498 17232 17510
rect 16456 17451 16944 17457
rect 16456 17417 16468 17451
rect 16932 17417 16944 17451
rect 16456 17411 16944 17417
rect 13452 16876 16220 16936
rect 13392 16870 13452 16876
rect 12232 16786 12292 16792
rect 17502 16786 17562 19132
rect 17636 18040 17696 21968
rect 17746 21358 17752 21418
rect 17812 21358 17818 21418
rect 17752 19296 17812 21358
rect 17994 20454 18054 24716
rect 18438 24586 18502 24716
rect 18432 24522 18438 24586
rect 18502 24522 18508 24586
rect 18262 24436 18322 24442
rect 18262 21500 18322 24376
rect 18940 24330 19000 24885
rect 19460 24834 19520 24984
rect 20476 24984 20492 25008
rect 20526 25514 20544 25560
rect 21496 25560 21560 25912
rect 21990 25764 22050 26021
rect 22514 25874 22578 26120
rect 23530 26120 23546 26156
rect 23580 26662 23588 26696
rect 24550 26696 24610 26846
rect 25060 26795 25120 27157
rect 24846 26789 25334 26795
rect 24846 26755 24858 26789
rect 25322 26755 25334 26789
rect 24846 26749 25334 26755
rect 24550 26670 24564 26696
rect 23580 26156 23586 26662
rect 23580 26154 23590 26156
rect 23580 26120 23594 26154
rect 22810 26061 23298 26067
rect 22810 26027 22822 26061
rect 23286 26027 23298 26061
rect 22810 26021 23298 26027
rect 22348 25810 22354 25874
rect 22418 25810 22578 25874
rect 23014 25764 23074 26021
rect 23530 25972 23594 26120
rect 24558 26120 24564 26670
rect 24598 26670 24610 26696
rect 25566 26696 25630 27256
rect 26588 27256 26600 27294
rect 26634 27294 26640 27832
rect 27608 27832 27668 27986
rect 28098 27931 28158 28434
rect 28618 28046 28678 28434
rect 28612 27986 28618 28046
rect 28678 27986 28684 28046
rect 27900 27925 28388 27931
rect 27900 27891 27912 27925
rect 28376 27891 28388 27925
rect 27900 27885 28388 27891
rect 27608 27794 27618 27832
rect 27612 27296 27618 27794
rect 26634 27256 26648 27294
rect 26076 27203 26136 27209
rect 25864 27197 26352 27203
rect 25864 27163 25876 27197
rect 26340 27163 26352 27197
rect 25864 27157 26352 27163
rect 26076 26795 26136 27157
rect 26588 27110 26648 27256
rect 27604 27256 27618 27296
rect 27652 27794 27668 27832
rect 28618 27832 28678 27986
rect 29126 27931 29186 28434
rect 29640 28046 29700 28434
rect 30146 28228 30152 28288
rect 30212 28228 30218 28288
rect 31158 28228 31164 28288
rect 31224 28228 31230 28288
rect 29634 27986 29640 28046
rect 29700 27986 29706 28046
rect 28918 27925 29406 27931
rect 28918 27891 28930 27925
rect 29394 27891 29406 27925
rect 28918 27885 29406 27891
rect 29126 27882 29186 27885
rect 27652 27296 27658 27794
rect 28618 27762 28636 27832
rect 27652 27256 27668 27296
rect 27088 27203 27148 27209
rect 26882 27197 27370 27203
rect 26882 27163 26894 27197
rect 27358 27163 27370 27197
rect 26882 27157 27370 27163
rect 26582 27050 26588 27110
rect 26648 27050 26654 27110
rect 27088 26906 27148 27157
rect 26580 26846 26586 26906
rect 26646 26846 26652 26906
rect 27082 26846 27088 26906
rect 27148 26846 27154 26906
rect 25864 26789 26352 26795
rect 25864 26755 25876 26789
rect 26340 26755 26352 26789
rect 25864 26749 26352 26755
rect 26076 26746 26136 26749
rect 24598 26120 24604 26670
rect 25566 26664 25582 26696
rect 25576 26168 25582 26664
rect 24558 26108 24604 26120
rect 25568 26120 25582 26168
rect 25616 26664 25630 26696
rect 26586 26696 26646 26846
rect 27088 26795 27148 26846
rect 26882 26789 27370 26795
rect 26882 26755 26894 26789
rect 27358 26755 27370 26789
rect 26882 26749 27370 26755
rect 27088 26746 27148 26749
rect 26586 26664 26600 26696
rect 25616 26168 25622 26664
rect 25616 26166 25628 26168
rect 25616 26120 25632 26166
rect 26594 26150 26600 26664
rect 24042 26067 24102 26074
rect 23828 26061 24316 26067
rect 23828 26027 23840 26061
rect 24304 26027 24316 26061
rect 23828 26021 24316 26027
rect 24846 26061 25334 26067
rect 24846 26027 24858 26061
rect 25322 26027 25334 26061
rect 24846 26021 25334 26027
rect 23524 25912 23530 25972
rect 23590 25912 23596 25972
rect 21984 25704 21990 25764
rect 22050 25704 22056 25764
rect 23008 25704 23014 25764
rect 23074 25704 23080 25764
rect 21792 25653 22280 25659
rect 21792 25619 21804 25653
rect 22268 25619 22280 25653
rect 21792 25613 22280 25619
rect 22810 25653 23298 25659
rect 22810 25619 22822 25653
rect 23286 25619 23298 25653
rect 22810 25613 23298 25619
rect 20526 25510 20542 25514
rect 21496 25512 21510 25560
rect 20526 25008 20532 25510
rect 21504 25010 21510 25512
rect 20526 24984 20540 25008
rect 19756 24925 20244 24931
rect 19756 24891 19768 24925
rect 20232 24891 20244 24925
rect 19756 24885 20244 24891
rect 19454 24774 19460 24834
rect 19520 24774 19526 24834
rect 19982 24330 20042 24885
rect 20476 24724 20540 24984
rect 21496 24984 21510 25010
rect 21544 25512 21560 25560
rect 22522 25560 22568 25572
rect 21544 25010 21550 25512
rect 22522 25040 22528 25560
rect 21544 25008 21556 25010
rect 21544 24984 21560 25008
rect 20774 24925 21262 24931
rect 20774 24891 20786 24925
rect 21250 24891 21262 24925
rect 20774 24885 21262 24891
rect 20470 24660 20476 24724
rect 20540 24660 20546 24724
rect 20982 24330 21042 24885
rect 21496 24834 21560 24984
rect 22516 24984 22528 25040
rect 22562 25040 22568 25560
rect 23530 25560 23594 25912
rect 24042 25764 24102 26021
rect 24036 25704 24042 25764
rect 24102 25704 24108 25764
rect 24042 25659 24102 25704
rect 25070 25659 25130 26021
rect 25568 25970 25632 26120
rect 26588 26120 26600 26150
rect 26634 26664 26646 26696
rect 27604 26696 27668 27256
rect 28630 27256 28636 27762
rect 28670 27762 28678 27832
rect 29640 27832 29700 27986
rect 30152 27931 30212 28228
rect 31164 27931 31224 28228
rect 31676 28046 31736 28434
rect 32176 28228 32182 28288
rect 32242 28228 32248 28288
rect 31670 27986 31676 28046
rect 31736 27986 31742 28046
rect 29936 27925 30424 27931
rect 29936 27891 29948 27925
rect 30412 27891 30424 27925
rect 29936 27885 30424 27891
rect 30954 27925 31442 27931
rect 30954 27891 30966 27925
rect 31430 27891 31442 27925
rect 30954 27885 31442 27891
rect 29640 27804 29654 27832
rect 28670 27256 28676 27762
rect 29648 27304 29654 27804
rect 28630 27244 28676 27256
rect 29640 27256 29654 27304
rect 29688 27804 29700 27832
rect 30666 27832 30712 27844
rect 29688 27304 29694 27804
rect 29688 27256 29700 27304
rect 30666 27288 30672 27832
rect 27900 27197 28388 27203
rect 27900 27163 27912 27197
rect 28376 27163 28388 27197
rect 27900 27157 28388 27163
rect 28918 27197 29406 27203
rect 28918 27163 28930 27197
rect 29394 27163 29406 27197
rect 28918 27157 29406 27163
rect 28616 26946 28622 27006
rect 28682 26946 28688 27006
rect 28102 26846 28108 26906
rect 28168 26846 28174 26906
rect 28108 26795 28168 26846
rect 27900 26789 28388 26795
rect 27900 26755 27912 26789
rect 28376 26755 28388 26789
rect 27900 26749 28388 26755
rect 26634 26150 26640 26664
rect 27604 26648 27618 26696
rect 27612 26164 27618 26648
rect 26634 26120 26648 26150
rect 26088 26067 26148 26079
rect 25864 26061 26352 26067
rect 25864 26027 25876 26061
rect 26340 26027 26352 26061
rect 25864 26021 26352 26027
rect 25562 25910 25568 25970
rect 25628 25910 25634 25970
rect 23828 25653 24316 25659
rect 23828 25619 23840 25653
rect 24304 25619 24316 25653
rect 23828 25613 24316 25619
rect 24846 25653 25334 25659
rect 24846 25619 24858 25653
rect 25322 25619 25334 25653
rect 24846 25613 25334 25619
rect 25070 25606 25130 25613
rect 23530 25500 23546 25560
rect 22562 24984 22576 25040
rect 23540 25018 23546 25500
rect 22018 24931 22078 24934
rect 21792 24925 22280 24931
rect 21792 24891 21804 24925
rect 22268 24891 22280 24925
rect 21792 24885 22280 24891
rect 22018 24834 22078 24885
rect 22516 24834 22576 24984
rect 23530 24984 23546 25018
rect 23580 25500 23594 25560
rect 24558 25560 24604 25572
rect 23580 25018 23586 25500
rect 23580 25016 23590 25018
rect 24558 25016 24564 25560
rect 23580 24984 23594 25016
rect 22810 24925 23298 24931
rect 22810 24891 22822 24925
rect 23286 24891 23298 24925
rect 22810 24885 23298 24891
rect 21490 24774 21496 24834
rect 21556 24774 21562 24834
rect 22012 24774 22018 24834
rect 22078 24774 22084 24834
rect 22510 24774 22516 24834
rect 22576 24774 22582 24834
rect 22990 24830 23050 24885
rect 23530 24838 23594 24984
rect 24548 24984 24564 25016
rect 24598 25016 24604 25560
rect 25568 25560 25632 25910
rect 26088 25659 26148 26021
rect 26588 25872 26648 26120
rect 27604 26120 27618 26164
rect 27652 26648 27668 26696
rect 28622 26696 28682 26946
rect 29128 26846 29134 26906
rect 29194 26846 29200 26906
rect 29640 26902 29700 27256
rect 30656 27256 30672 27288
rect 30706 27288 30712 27832
rect 31676 27832 31736 27986
rect 32182 27931 32242 28228
rect 32696 27994 33776 28054
rect 31972 27925 32460 27931
rect 31972 27891 31984 27925
rect 32448 27891 32460 27925
rect 31972 27885 32460 27891
rect 31676 27800 31690 27832
rect 31684 27294 31690 27800
rect 30706 27256 30716 27288
rect 29936 27197 30424 27203
rect 29936 27163 29948 27197
rect 30412 27163 30424 27197
rect 29936 27157 30424 27163
rect 30656 27006 30716 27256
rect 31680 27256 31690 27294
rect 31724 27800 31736 27832
rect 32696 27832 32756 27994
rect 33198 27931 33258 27994
rect 32990 27925 33478 27931
rect 32990 27891 33002 27925
rect 33466 27891 33478 27925
rect 32990 27885 33478 27891
rect 32696 27802 32708 27832
rect 31724 27294 31730 27800
rect 32702 27296 32708 27802
rect 31724 27256 31740 27294
rect 30954 27197 31442 27203
rect 30954 27163 30966 27197
rect 31430 27163 31442 27197
rect 30954 27157 31442 27163
rect 30650 26946 30656 27006
rect 30716 26946 30722 27006
rect 31680 26908 31740 27256
rect 32696 27256 32708 27296
rect 32742 27802 32756 27832
rect 33716 27832 33776 27994
rect 32742 27296 32748 27802
rect 33716 27786 33726 27832
rect 32742 27256 32756 27296
rect 32160 27203 32220 27215
rect 31972 27197 32460 27203
rect 31972 27163 31984 27197
rect 32448 27163 32460 27197
rect 31972 27157 32460 27163
rect 31680 26902 31744 26908
rect 29134 26795 29194 26846
rect 29634 26842 29640 26902
rect 29700 26842 29706 26902
rect 30148 26842 30154 26902
rect 30214 26842 30220 26902
rect 30652 26842 30658 26902
rect 30718 26842 30724 26902
rect 31158 26842 31164 26902
rect 31224 26842 31230 26902
rect 31680 26842 31684 26902
rect 28918 26789 29406 26795
rect 28918 26755 28930 26789
rect 29394 26755 29406 26789
rect 28918 26749 29406 26755
rect 28622 26672 28636 26696
rect 27652 26164 27658 26648
rect 27652 26162 27664 26164
rect 27652 26120 27668 26162
rect 27088 26067 27148 26075
rect 26882 26061 27370 26067
rect 26882 26027 26894 26061
rect 27358 26027 27370 26061
rect 26882 26021 27370 26027
rect 26582 25812 26588 25872
rect 26648 25812 26654 25872
rect 27088 25659 27148 26021
rect 27604 25970 27668 26120
rect 28630 26120 28636 26672
rect 28670 26672 28682 26696
rect 29640 26696 29700 26842
rect 30154 26795 30214 26842
rect 29936 26789 30424 26795
rect 29936 26755 29948 26789
rect 30412 26755 30424 26789
rect 29936 26749 30424 26755
rect 28670 26120 28676 26672
rect 29640 26652 29654 26696
rect 29648 26156 29654 26652
rect 28630 26108 28676 26120
rect 29640 26120 29654 26156
rect 29688 26652 29700 26696
rect 30658 26696 30718 26842
rect 31164 26795 31224 26842
rect 31680 26836 31744 26842
rect 30954 26789 31442 26795
rect 30954 26755 30966 26789
rect 31430 26755 31442 26789
rect 30954 26749 31442 26755
rect 30658 26668 30672 26696
rect 29688 26156 29694 26652
rect 30666 26190 30672 26668
rect 29688 26120 29700 26156
rect 27900 26061 28388 26067
rect 27900 26027 27912 26061
rect 28376 26027 28388 26061
rect 27900 26021 28388 26027
rect 28918 26061 29406 26067
rect 28918 26027 28930 26061
rect 29394 26027 29406 26061
rect 28918 26021 29406 26027
rect 29640 25970 29700 26120
rect 30656 26120 30672 26190
rect 30706 26668 30718 26696
rect 31680 26696 31740 26836
rect 32160 26795 32220 27157
rect 32696 27110 32756 27256
rect 33720 27256 33726 27786
rect 33760 27786 33776 27832
rect 33760 27256 33766 27786
rect 33720 27244 33766 27256
rect 32990 27197 33478 27203
rect 32990 27163 33002 27197
rect 33466 27163 33478 27197
rect 32990 27157 33478 27163
rect 32690 27050 32696 27110
rect 32756 27050 32762 27110
rect 33940 27050 33946 27110
rect 34006 27050 34012 27110
rect 32700 26834 33770 26894
rect 31972 26789 32460 26795
rect 31972 26755 31984 26789
rect 32448 26755 32460 26789
rect 31972 26749 32460 26755
rect 30706 26190 30712 26668
rect 31680 26660 31690 26696
rect 30706 26120 30716 26190
rect 31684 26152 31690 26660
rect 29936 26061 30424 26067
rect 29936 26027 29948 26061
rect 30412 26027 30424 26061
rect 29936 26021 30424 26027
rect 30142 25970 30202 26021
rect 27598 25910 27604 25970
rect 27664 25910 27670 25970
rect 28098 25910 28104 25970
rect 28164 25910 28170 25970
rect 28612 25910 28618 25970
rect 28678 25910 28684 25970
rect 29136 25910 29142 25970
rect 29202 25910 29208 25970
rect 29634 25910 29640 25970
rect 29700 25910 29706 25970
rect 30136 25910 30142 25970
rect 30202 25910 30208 25970
rect 30656 25968 30716 26120
rect 31674 26120 31690 26152
rect 31724 26660 31740 26696
rect 32700 26696 32760 26834
rect 33206 26795 33266 26834
rect 32990 26789 33478 26795
rect 32990 26755 33002 26789
rect 33466 26755 33478 26789
rect 32990 26749 33478 26755
rect 32700 26668 32708 26696
rect 31724 26152 31730 26660
rect 31724 26150 31734 26152
rect 32702 26150 32708 26668
rect 31724 26120 31738 26150
rect 31164 26067 31224 26074
rect 30954 26061 31442 26067
rect 30954 26027 30966 26061
rect 31430 26027 31442 26061
rect 30954 26021 31442 26027
rect 31164 25968 31224 26021
rect 31674 25968 31738 26120
rect 32696 26120 32708 26150
rect 32742 26668 32760 26696
rect 33710 26696 33770 26834
rect 32742 26150 32748 26668
rect 33710 26662 33726 26696
rect 32742 26120 32756 26150
rect 32160 26067 32220 26073
rect 31972 26061 32460 26067
rect 31972 26027 31984 26061
rect 32448 26027 32460 26061
rect 31972 26021 32460 26027
rect 25864 25653 26352 25659
rect 25864 25619 25876 25653
rect 26340 25619 26352 25653
rect 25864 25613 26352 25619
rect 26882 25653 27370 25659
rect 26882 25619 26894 25653
rect 27358 25619 27370 25653
rect 26882 25613 27370 25619
rect 27088 25612 27148 25613
rect 25568 25520 25582 25560
rect 25576 25044 25582 25520
rect 24598 24984 24612 25016
rect 23828 24925 24316 24931
rect 23828 24891 23840 24925
rect 24304 24891 24316 24925
rect 23828 24885 24316 24891
rect 18372 24270 18378 24330
rect 18438 24270 18444 24330
rect 18934 24270 18940 24330
rect 19000 24270 19006 24330
rect 19976 24270 19982 24330
rect 20042 24270 20048 24330
rect 20976 24270 20982 24330
rect 21042 24270 21048 24330
rect 18378 21688 18438 24270
rect 22990 24232 23050 24770
rect 23498 24834 23594 24838
rect 23498 24832 23530 24834
rect 23590 24774 23596 24834
rect 23984 24774 23990 24834
rect 24050 24774 24056 24834
rect 23498 24232 23558 24772
rect 23990 24232 24050 24774
rect 24144 24330 24204 24885
rect 24548 24582 24612 24984
rect 25566 24984 25582 25044
rect 25616 25520 25632 25560
rect 26594 25560 26640 25572
rect 25616 25044 25622 25520
rect 25616 24984 25626 25044
rect 26594 25020 26600 25560
rect 24846 24925 25334 24931
rect 24846 24891 24858 24925
rect 25322 24891 25334 24925
rect 24846 24885 25334 24891
rect 24548 24512 24612 24518
rect 25034 24836 25094 24842
rect 24138 24270 24144 24330
rect 24204 24270 24210 24330
rect 25034 24232 25094 24776
rect 25154 24330 25214 24885
rect 25566 24834 25626 24984
rect 26584 24984 26600 25020
rect 26634 25020 26640 25560
rect 27604 25560 27668 25910
rect 28104 25659 28164 25910
rect 27900 25653 28388 25659
rect 27900 25619 27912 25653
rect 28376 25619 28388 25653
rect 27900 25613 28388 25619
rect 27604 25508 27618 25560
rect 27612 25026 27618 25508
rect 26634 24984 26648 25020
rect 25864 24925 26352 24931
rect 25864 24891 25876 24925
rect 26340 24891 26352 24925
rect 25864 24885 26352 24891
rect 25560 24774 25566 24834
rect 25626 24774 25632 24834
rect 26096 24330 26156 24885
rect 26584 24440 26648 24984
rect 27604 24984 27618 25026
rect 27652 25508 27668 25560
rect 28618 25560 28678 25910
rect 29142 25659 29202 25910
rect 28918 25653 29406 25659
rect 28918 25619 28930 25653
rect 29394 25619 29406 25653
rect 28918 25613 29406 25619
rect 27652 25026 27658 25508
rect 28618 25506 28636 25560
rect 28630 25430 28636 25506
rect 27652 25024 27664 25026
rect 27652 24984 27668 25024
rect 26882 24925 27370 24931
rect 26882 24891 26894 24925
rect 27358 24891 27370 24925
rect 26882 24885 27370 24891
rect 27078 24836 27138 24842
rect 27604 24836 27668 24984
rect 28622 24984 28636 25430
rect 28670 25506 28678 25560
rect 29640 25560 29700 25910
rect 30650 25908 30656 25968
rect 30716 25908 30722 25968
rect 31158 25908 31164 25968
rect 31224 25908 31230 25968
rect 31668 25908 31674 25968
rect 31734 25908 31740 25968
rect 30140 25696 30146 25756
rect 30206 25696 30212 25756
rect 31152 25696 31158 25756
rect 31218 25696 31224 25756
rect 30146 25659 30206 25696
rect 31158 25659 31218 25696
rect 29936 25653 30424 25659
rect 29936 25619 29948 25653
rect 30412 25619 30424 25653
rect 29936 25613 30424 25619
rect 30954 25653 31442 25659
rect 30954 25619 30966 25653
rect 31430 25619 31442 25653
rect 30954 25613 31442 25619
rect 29640 25506 29654 25560
rect 28670 25430 28676 25506
rect 28670 24984 28682 25430
rect 29648 25014 29654 25506
rect 28100 24931 28160 24940
rect 27900 24925 28388 24931
rect 27900 24891 27912 24925
rect 28376 24891 28388 24925
rect 27900 24885 28388 24891
rect 26578 24376 26584 24440
rect 26648 24376 26654 24440
rect 25148 24270 25154 24330
rect 25214 24270 25220 24330
rect 26090 24270 26096 24330
rect 26156 24270 26162 24330
rect 27078 24232 27138 24776
rect 27572 24832 27668 24836
rect 27572 24830 27604 24832
rect 27664 24772 27670 24832
rect 28100 24826 28160 24885
rect 28622 24836 28682 24984
rect 29640 24984 29654 25014
rect 29688 25506 29700 25560
rect 30666 25560 30712 25572
rect 29688 25014 29694 25506
rect 30666 25018 30672 25560
rect 29688 25012 29700 25014
rect 29688 24984 29704 25012
rect 29100 24931 29160 24934
rect 28918 24925 29406 24931
rect 28918 24891 28930 24925
rect 29394 24891 29406 24925
rect 28918 24885 29406 24891
rect 27572 24232 27632 24770
rect 28100 24232 28160 24766
rect 28588 24830 28682 24836
rect 28648 24828 28682 24830
rect 28588 24768 28622 24770
rect 28588 24762 28682 24768
rect 29100 24826 29160 24885
rect 29640 24830 29704 24984
rect 30656 24984 30672 25018
rect 30706 25018 30712 25560
rect 31674 25560 31738 25908
rect 32160 25756 32220 26021
rect 32696 25872 32756 26120
rect 33720 26120 33726 26662
rect 33760 26662 33770 26696
rect 33760 26120 33766 26662
rect 33720 26108 33766 26120
rect 32990 26061 33478 26067
rect 32990 26027 33002 26061
rect 33466 26027 33478 26061
rect 32990 26021 33478 26027
rect 32690 25812 32696 25872
rect 32756 25812 32762 25872
rect 32698 25758 32758 25760
rect 32154 25696 32160 25756
rect 32220 25696 32226 25756
rect 32698 25698 33770 25758
rect 32160 25659 32220 25696
rect 31972 25653 32460 25659
rect 31972 25619 31984 25653
rect 32448 25619 32460 25653
rect 31972 25613 32460 25619
rect 32160 25610 32220 25613
rect 31674 25514 31690 25560
rect 30706 24984 30720 25018
rect 31684 25014 31690 25514
rect 29936 24925 30424 24931
rect 29936 24891 29948 24925
rect 30412 24891 30424 24925
rect 29936 24885 30424 24891
rect 29634 24770 29640 24830
rect 29700 24770 29706 24830
rect 28588 24232 28648 24762
rect 29100 24232 29160 24766
rect 30656 24724 30720 24984
rect 31674 24984 31690 25014
rect 31724 25514 31738 25560
rect 32698 25560 32758 25698
rect 33202 25659 33262 25698
rect 32990 25653 33478 25659
rect 32990 25619 33002 25653
rect 33466 25619 33478 25653
rect 32990 25613 33478 25619
rect 32698 25534 32708 25560
rect 31724 25014 31730 25514
rect 32702 25072 32708 25534
rect 31724 25012 31734 25014
rect 31724 24984 31738 25012
rect 30954 24925 31442 24931
rect 30954 24891 30966 24925
rect 31430 24891 31442 24925
rect 30954 24885 31442 24891
rect 31674 24830 31738 24984
rect 32690 24984 32708 25072
rect 32742 25534 32758 25560
rect 33710 25560 33770 25698
rect 32742 25072 32748 25534
rect 33710 25510 33726 25560
rect 32742 24984 32750 25072
rect 31972 24925 32460 24931
rect 31972 24891 31984 24925
rect 32448 24891 32460 24925
rect 31972 24885 32460 24891
rect 31668 24770 31674 24830
rect 31734 24770 31740 24830
rect 30650 24660 30656 24724
rect 30720 24660 30726 24724
rect 32690 24436 32750 24984
rect 33720 24984 33726 25510
rect 33760 25510 33770 25560
rect 33760 24984 33766 25510
rect 33720 24972 33766 24984
rect 32990 24925 33478 24931
rect 32990 24891 33002 24925
rect 33466 24891 33478 24925
rect 32990 24885 33478 24891
rect 33946 24592 34006 27050
rect 33942 24586 34006 24592
rect 33942 24516 34006 24522
rect 32684 24376 32690 24436
rect 32750 24376 32756 24436
rect 20654 24172 30894 24232
rect 18486 24068 18492 24128
rect 18552 24068 18558 24128
rect 18492 22154 18552 24068
rect 18914 24015 19402 24021
rect 18914 23981 18926 24015
rect 19390 23981 19402 24015
rect 18914 23975 19402 23981
rect 19932 24015 20420 24021
rect 19932 23981 19944 24015
rect 20408 23981 20420 24015
rect 19932 23975 20420 23981
rect 18626 23922 18672 23934
rect 18626 23376 18632 23922
rect 18618 23346 18632 23376
rect 18666 23376 18672 23922
rect 19644 23922 19690 23934
rect 18666 23346 18678 23376
rect 19644 23370 19650 23922
rect 18618 23194 18678 23346
rect 19636 23346 19650 23370
rect 19684 23370 19690 23922
rect 20654 23922 20714 24172
rect 21664 24068 21670 24128
rect 21730 24068 21736 24128
rect 20950 24015 21438 24021
rect 20950 23981 20962 24015
rect 21426 23981 21438 24015
rect 20950 23975 21438 23981
rect 19684 23346 19696 23370
rect 18914 23287 19402 23293
rect 18914 23253 18926 23287
rect 19390 23253 19402 23287
rect 18914 23247 19402 23253
rect 19130 23194 19190 23247
rect 19636 23194 19696 23346
rect 20654 23346 20668 23922
rect 20702 23346 20714 23922
rect 21670 23922 21730 24068
rect 21968 24015 22456 24021
rect 21968 23981 21980 24015
rect 22444 23981 22456 24015
rect 21968 23975 22456 23981
rect 21670 23858 21686 23922
rect 19932 23287 20420 23293
rect 19932 23253 19944 23287
rect 20408 23253 20420 23287
rect 19932 23247 20420 23253
rect 18618 23192 19696 23194
rect 18618 23134 19636 23192
rect 19630 23132 19636 23134
rect 19696 23132 19702 23192
rect 20140 23084 20200 23247
rect 20134 23024 20140 23084
rect 20200 23024 20206 23084
rect 20140 22989 20200 23024
rect 18914 22983 19402 22989
rect 18914 22949 18926 22983
rect 19390 22949 19402 22983
rect 18914 22943 19402 22949
rect 19932 22983 20420 22989
rect 19932 22949 19944 22983
rect 20408 22949 20420 22983
rect 19932 22943 20420 22949
rect 18626 22890 18672 22902
rect 18626 22370 18632 22890
rect 18618 22314 18632 22370
rect 18666 22370 18672 22890
rect 19644 22890 19690 22902
rect 18666 22314 18678 22370
rect 19644 22344 19650 22890
rect 18618 22154 18678 22314
rect 19632 22314 19650 22344
rect 19684 22344 19690 22890
rect 20654 22890 20714 23346
rect 21680 23346 21686 23858
rect 21720 23858 21730 23922
rect 22692 23922 22752 24172
rect 22986 24015 23474 24021
rect 22986 23981 22998 24015
rect 23462 23981 23474 24015
rect 22986 23975 23474 23981
rect 24004 24015 24492 24021
rect 24004 23981 24016 24015
rect 24480 23981 24492 24015
rect 24004 23975 24492 23981
rect 21720 23346 21726 23858
rect 21680 23334 21726 23346
rect 22692 23346 22704 23922
rect 22738 23346 22752 23922
rect 23716 23922 23762 23934
rect 23716 23410 23722 23922
rect 21160 23293 21220 23299
rect 20950 23287 21438 23293
rect 20950 23253 20962 23287
rect 21426 23253 21438 23287
rect 20950 23247 21438 23253
rect 21968 23287 22456 23293
rect 21968 23253 21980 23287
rect 22444 23253 22456 23287
rect 21968 23247 22456 23253
rect 21160 23090 21220 23247
rect 21664 23132 21670 23192
rect 21730 23132 21736 23192
rect 21160 23084 21222 23090
rect 21160 23024 21162 23084
rect 21160 23018 21222 23024
rect 21160 22989 21220 23018
rect 20950 22983 21438 22989
rect 20950 22949 20962 22983
rect 21426 22949 21438 22983
rect 20950 22943 21438 22949
rect 19684 22314 19692 22344
rect 18914 22255 19402 22261
rect 18914 22221 18926 22255
rect 19390 22221 19402 22255
rect 18914 22215 19402 22221
rect 19120 22154 19180 22215
rect 19632 22160 19692 22314
rect 20654 22314 20668 22890
rect 20702 22314 20714 22890
rect 21670 22890 21730 23132
rect 22182 23090 22242 23247
rect 22180 23084 22242 23090
rect 22240 23024 22242 23084
rect 22180 23018 22242 23024
rect 22182 22989 22242 23018
rect 21968 22983 22456 22989
rect 21968 22949 21980 22983
rect 22444 22949 22456 22983
rect 21968 22943 22456 22949
rect 22182 22936 22242 22943
rect 21670 22844 21686 22890
rect 19932 22255 20420 22261
rect 19932 22221 19944 22255
rect 20408 22221 20420 22255
rect 19932 22215 20420 22221
rect 19626 22154 19632 22160
rect 18492 22100 19632 22154
rect 19692 22100 19698 22160
rect 18492 22094 19698 22100
rect 20138 22026 20198 22215
rect 20138 21960 20198 21966
rect 20654 21818 20714 22314
rect 21680 22314 21686 22844
rect 21720 22844 21730 22890
rect 22692 22890 22752 23346
rect 23712 23346 23722 23410
rect 23756 23410 23762 23922
rect 24730 23922 24790 24172
rect 25732 24068 25738 24128
rect 25798 24068 25804 24128
rect 25022 24015 25510 24021
rect 25022 23981 25034 24015
rect 25498 23981 25510 24015
rect 25022 23975 25510 23981
rect 23756 23346 23772 23410
rect 22986 23287 23474 23293
rect 22986 23253 22998 23287
rect 23462 23253 23474 23287
rect 22986 23247 23474 23253
rect 23202 23090 23262 23247
rect 23712 23192 23772 23346
rect 24730 23346 24740 23922
rect 24774 23346 24790 23922
rect 25738 23922 25798 24068
rect 26040 24015 26528 24021
rect 26040 23981 26052 24015
rect 26516 23981 26528 24015
rect 26040 23975 26528 23981
rect 25738 23848 25758 23922
rect 24218 23293 24278 23295
rect 24004 23287 24492 23293
rect 24004 23253 24016 23287
rect 24480 23253 24492 23287
rect 24004 23247 24492 23253
rect 23706 23132 23712 23192
rect 23772 23132 23778 23192
rect 23202 23084 23264 23090
rect 23202 23024 23204 23084
rect 23202 23018 23264 23024
rect 24218 23084 24278 23247
rect 23202 22989 23262 23018
rect 24218 22989 24278 23024
rect 22986 22983 23474 22989
rect 22986 22949 22998 22983
rect 23462 22949 23474 22983
rect 22986 22943 23474 22949
rect 24004 22983 24492 22989
rect 24004 22949 24016 22983
rect 24480 22949 24492 22983
rect 24004 22943 24492 22949
rect 21720 22314 21726 22844
rect 21680 22302 21726 22314
rect 22692 22314 22704 22890
rect 22738 22314 22752 22890
rect 23716 22890 23762 22902
rect 23716 22380 23722 22890
rect 21152 22261 21212 22264
rect 20950 22255 21438 22261
rect 20950 22221 20962 22255
rect 21426 22221 21438 22255
rect 20950 22215 21438 22221
rect 21968 22255 22456 22261
rect 21968 22221 21980 22255
rect 22444 22221 22456 22255
rect 21968 22215 22456 22221
rect 21152 22022 21212 22215
rect 22184 22030 22244 22215
rect 22184 21964 22244 21970
rect 21152 21956 21212 21962
rect 22692 21818 22752 22314
rect 23712 22314 23722 22380
rect 23756 22380 23762 22890
rect 24730 22890 24790 23346
rect 25752 23346 25758 23848
rect 25792 23346 25798 23922
rect 25752 23334 25798 23346
rect 26766 23922 26826 24172
rect 27058 24015 27546 24021
rect 27058 23981 27070 24015
rect 27534 23981 27546 24015
rect 27058 23975 27546 23981
rect 28076 24015 28564 24021
rect 28076 23981 28088 24015
rect 28552 23981 28564 24015
rect 28076 23975 28564 23981
rect 26766 23346 26776 23922
rect 26810 23346 26826 23922
rect 27788 23922 27834 23934
rect 27788 23410 27794 23922
rect 25022 23287 25510 23293
rect 25022 23253 25034 23287
rect 25498 23253 25510 23287
rect 25022 23247 25510 23253
rect 26040 23287 26528 23293
rect 26040 23253 26052 23287
rect 26516 23253 26528 23287
rect 26040 23247 26528 23253
rect 25234 23090 25294 23247
rect 25732 23132 25738 23192
rect 25798 23132 25804 23192
rect 25234 23084 25296 23090
rect 25234 23024 25236 23084
rect 25234 23018 25296 23024
rect 25234 22989 25294 23018
rect 25022 22983 25510 22989
rect 25022 22949 25034 22983
rect 25498 22949 25510 22983
rect 25022 22943 25510 22949
rect 23756 22314 23772 22380
rect 22986 22255 23474 22261
rect 22986 22221 22998 22255
rect 23462 22221 23474 22255
rect 22986 22215 23474 22221
rect 23182 22030 23242 22215
rect 23712 22160 23772 22314
rect 24730 22314 24740 22890
rect 24774 22314 24790 22890
rect 25738 22890 25798 23132
rect 26244 23090 26304 23247
rect 26244 23084 26306 23090
rect 26244 23024 26246 23084
rect 26244 23018 26306 23024
rect 26244 22989 26304 23018
rect 26040 22983 26528 22989
rect 26040 22949 26052 22983
rect 26516 22949 26528 22983
rect 26040 22943 26528 22949
rect 25738 22828 25758 22890
rect 25752 22406 25758 22828
rect 24226 22261 24286 22274
rect 24004 22255 24492 22261
rect 24004 22221 24016 22255
rect 24480 22221 24492 22255
rect 24004 22215 24492 22221
rect 23706 22100 23712 22160
rect 23772 22100 23778 22160
rect 23182 21964 23242 21970
rect 24226 22030 24286 22215
rect 24226 21964 24286 21970
rect 24730 21818 24790 22314
rect 25748 22314 25758 22406
rect 25792 22406 25798 22890
rect 26766 22890 26826 23346
rect 27780 23346 27794 23410
rect 27828 23410 27834 23922
rect 28796 23922 28856 24172
rect 29808 24068 29814 24128
rect 29874 24068 29880 24128
rect 29094 24015 29582 24021
rect 29094 23981 29106 24015
rect 29570 23981 29582 24015
rect 29094 23975 29582 23981
rect 28796 23512 28812 23922
rect 28806 23418 28812 23512
rect 27828 23346 27840 23410
rect 27266 23293 27326 23295
rect 27058 23287 27546 23293
rect 27058 23253 27070 23287
rect 27534 23253 27546 23287
rect 27058 23247 27546 23253
rect 27266 23090 27326 23247
rect 27780 23192 27840 23346
rect 28796 23346 28812 23418
rect 28846 23512 28856 23922
rect 29814 23922 29874 24068
rect 30112 24015 30600 24021
rect 30112 23981 30124 24015
rect 30588 23981 30600 24015
rect 30112 23975 30600 23981
rect 29814 23858 29830 23922
rect 28846 23418 28852 23512
rect 28846 23346 28856 23418
rect 28280 23293 28340 23295
rect 28076 23287 28564 23293
rect 28076 23253 28088 23287
rect 28552 23253 28564 23287
rect 28076 23247 28564 23253
rect 27774 23132 27780 23192
rect 27840 23132 27846 23192
rect 28280 23090 28340 23247
rect 27266 23084 27328 23090
rect 27266 23024 27268 23084
rect 27266 23018 27328 23024
rect 28280 23084 28342 23090
rect 28280 23024 28282 23084
rect 28280 23018 28342 23024
rect 27266 22989 27326 23018
rect 28280 22989 28340 23018
rect 27058 22983 27546 22989
rect 27058 22949 27070 22983
rect 27534 22949 27546 22983
rect 27058 22943 27546 22949
rect 28076 22983 28564 22989
rect 28076 22949 28088 22983
rect 28552 22949 28564 22983
rect 28076 22943 28564 22949
rect 25792 22314 25808 22406
rect 25230 22261 25290 22264
rect 25022 22255 25510 22261
rect 25022 22221 25034 22255
rect 25498 22221 25510 22255
rect 25022 22215 25510 22221
rect 25230 22026 25290 22215
rect 25230 21960 25290 21966
rect 25748 21910 25808 22314
rect 26766 22314 26776 22890
rect 26810 22314 26826 22890
rect 27788 22890 27834 22902
rect 27788 22396 27794 22890
rect 26246 22261 26306 22268
rect 26040 22255 26528 22261
rect 26040 22221 26052 22255
rect 26516 22221 26528 22255
rect 26040 22215 26528 22221
rect 26246 22026 26306 22215
rect 26246 21960 26306 21966
rect 25538 21850 25808 21910
rect 20654 21758 25030 21818
rect 25090 21758 25096 21818
rect 18378 21628 22546 21688
rect 18256 21440 18262 21500
rect 18322 21440 18328 21500
rect 19422 21440 19428 21500
rect 19488 21440 19494 21500
rect 17988 20394 17994 20454
rect 18054 20394 18060 20454
rect 17746 19236 17752 19296
rect 17812 19236 17818 19296
rect 17742 19022 17748 19082
rect 17808 19022 17814 19082
rect 17630 17980 17636 18040
rect 17696 17980 17702 18040
rect 12292 16726 17562 16786
rect 12232 16720 12292 16726
rect -3042 16188 8228 16248
rect -3042 15700 -2976 16188
rect -2748 15992 8228 16188
rect 11322 16128 11434 16642
rect 13286 16524 13346 16530
rect 17748 16524 17808 19022
rect 17994 16782 18054 20394
rect 18124 20296 18130 20356
rect 18190 20296 18196 20356
rect 17988 16722 17994 16782
rect 18054 16722 18060 16782
rect 18130 16652 18190 20296
rect 18262 17832 18322 21440
rect 18706 21379 19194 21385
rect 18706 21345 18718 21379
rect 19182 21345 19194 21379
rect 18706 21339 19194 21345
rect 18418 21286 18464 21298
rect 18418 20746 18424 21286
rect 18410 20710 18424 20746
rect 18458 20746 18464 21286
rect 19428 21286 19488 21440
rect 19724 21379 20212 21385
rect 19724 21345 19736 21379
rect 20200 21345 20212 21379
rect 19724 21339 20212 21345
rect 19428 21260 19442 21286
rect 18458 20710 18470 20746
rect 19436 20734 19442 21260
rect 18410 20552 18470 20710
rect 19426 20710 19442 20734
rect 19476 21260 19488 21286
rect 20444 21286 20504 21628
rect 21458 21440 21464 21500
rect 21524 21440 21530 21500
rect 20742 21379 21230 21385
rect 20742 21345 20754 21379
rect 21218 21345 21230 21379
rect 20742 21339 21230 21345
rect 19476 20734 19482 21260
rect 20444 21240 20460 21286
rect 20454 20734 20460 21240
rect 19476 20710 19486 20734
rect 18706 20651 19194 20657
rect 18706 20617 18718 20651
rect 19182 20617 19194 20651
rect 18706 20611 19194 20617
rect 18924 20552 18984 20611
rect 19426 20552 19486 20710
rect 20446 20710 20460 20734
rect 20494 21240 20504 21286
rect 21464 21286 21524 21440
rect 21966 21436 21972 21500
rect 22036 21436 22042 21500
rect 21972 21385 22036 21436
rect 21760 21379 22248 21385
rect 21760 21345 21772 21379
rect 22236 21345 22248 21379
rect 21760 21339 22248 21345
rect 21464 21262 21478 21286
rect 20494 20734 20500 21240
rect 20494 20710 20506 20734
rect 19724 20651 20212 20657
rect 19724 20617 19736 20651
rect 20200 20617 20212 20651
rect 19724 20611 20212 20617
rect 18410 20492 19486 20552
rect 19916 20250 19976 20611
rect 20446 20552 20506 20710
rect 21472 20710 21478 21262
rect 21512 21262 21524 21286
rect 22486 21286 22546 21628
rect 22990 21385 23050 21758
rect 22778 21379 23266 21385
rect 22778 21345 22790 21379
rect 23254 21345 23266 21379
rect 22778 21339 23266 21345
rect 21512 20710 21518 21262
rect 22486 21232 22496 21286
rect 22490 20738 22496 21232
rect 21472 20698 21518 20710
rect 22482 20710 22496 20738
rect 22530 21232 22546 21286
rect 23498 21286 23558 21758
rect 23990 21385 24050 21758
rect 25028 21385 25088 21758
rect 23796 21379 24284 21385
rect 23796 21345 23808 21379
rect 24272 21345 24284 21379
rect 23796 21339 24284 21345
rect 24814 21379 25302 21385
rect 24814 21345 24826 21379
rect 25290 21345 25302 21379
rect 24814 21339 25302 21345
rect 22530 20738 22536 21232
rect 22530 20710 22542 20738
rect 20742 20651 21230 20657
rect 20742 20617 20754 20651
rect 21218 20617 21230 20651
rect 20742 20611 21230 20617
rect 21760 20651 22248 20657
rect 21760 20617 21772 20651
rect 22236 20617 22248 20651
rect 21760 20611 22248 20617
rect 20440 20492 20446 20552
rect 20506 20492 20512 20552
rect 20954 20498 21014 20611
rect 21960 20498 22020 20611
rect 22482 20552 22542 20710
rect 23498 20710 23514 21286
rect 23548 20710 23558 21286
rect 24526 21286 24572 21298
rect 24526 20734 24532 21286
rect 22778 20651 23266 20657
rect 22778 20617 22790 20651
rect 23254 20617 23266 20651
rect 22778 20611 23266 20617
rect 22992 20556 23052 20611
rect 23498 20556 23558 20710
rect 24518 20710 24532 20734
rect 24566 20734 24572 21286
rect 25538 21286 25598 21850
rect 26766 21818 26826 22314
rect 27780 22314 27794 22396
rect 27828 22396 27834 22890
rect 28796 22890 28856 23346
rect 29824 23346 29830 23858
rect 29864 23858 29874 23922
rect 30834 23922 30894 24172
rect 33004 24068 33010 24128
rect 33070 24068 33076 24128
rect 31130 24015 31618 24021
rect 31130 23981 31142 24015
rect 31606 23981 31618 24015
rect 31130 23975 31618 23981
rect 32148 24015 32636 24021
rect 32148 23981 32160 24015
rect 32624 23981 32636 24015
rect 32148 23975 32636 23981
rect 29864 23346 29870 23858
rect 29824 23334 29870 23346
rect 30834 23346 30848 23922
rect 30882 23346 30894 23922
rect 31860 23922 31906 23934
rect 31860 23422 31866 23922
rect 29312 23293 29372 23295
rect 30322 23293 30382 23295
rect 29094 23287 29582 23293
rect 29094 23253 29106 23287
rect 29570 23253 29582 23287
rect 29094 23247 29582 23253
rect 30112 23287 30600 23293
rect 30112 23253 30124 23287
rect 30588 23253 30600 23287
rect 30112 23247 30600 23253
rect 29312 23090 29372 23247
rect 29810 23132 29816 23192
rect 29876 23132 29882 23192
rect 29312 23084 29374 23090
rect 29312 23024 29314 23084
rect 29312 23018 29374 23024
rect 29312 22989 29372 23018
rect 29094 22983 29582 22989
rect 29094 22949 29106 22983
rect 29570 22949 29582 22983
rect 29094 22943 29582 22949
rect 27828 22314 27840 22396
rect 27058 22255 27546 22261
rect 27058 22221 27070 22255
rect 27534 22221 27546 22255
rect 27058 22215 27546 22221
rect 27250 22026 27310 22215
rect 27780 22160 27840 22314
rect 28796 22314 28812 22890
rect 28846 22314 28856 22890
rect 29816 22890 29876 23132
rect 30322 23090 30382 23247
rect 30322 23084 30384 23090
rect 30322 23024 30324 23084
rect 30322 23018 30384 23024
rect 30322 22989 30382 23018
rect 30112 22983 30600 22989
rect 30112 22949 30124 22983
rect 30588 22949 30600 22983
rect 30112 22943 30600 22949
rect 29816 22822 29830 22890
rect 28076 22255 28564 22261
rect 28076 22221 28088 22255
rect 28552 22221 28564 22255
rect 28076 22215 28564 22221
rect 27774 22100 27780 22160
rect 27840 22100 27846 22160
rect 27250 21960 27310 21966
rect 28282 22030 28342 22215
rect 28282 21964 28342 21970
rect 26040 21558 26046 21622
rect 26110 21558 26116 21622
rect 26046 21500 26110 21558
rect 26766 21528 26826 21758
rect 28796 21918 28856 22314
rect 29824 22314 29830 22822
rect 29864 22822 29876 22890
rect 30834 22890 30894 23346
rect 31852 23346 31866 23422
rect 31900 23422 31906 23922
rect 32878 23922 32924 23934
rect 31900 23346 31912 23422
rect 32878 23372 32884 23922
rect 31130 23287 31618 23293
rect 31130 23253 31142 23287
rect 31606 23253 31618 23287
rect 31130 23247 31618 23253
rect 31344 23090 31404 23247
rect 31852 23194 31912 23346
rect 32868 23346 32884 23372
rect 32918 23372 32924 23922
rect 32918 23346 32928 23372
rect 32148 23287 32636 23293
rect 32148 23253 32160 23287
rect 32624 23253 32636 23287
rect 32148 23247 32636 23253
rect 32374 23194 32434 23247
rect 32868 23194 32928 23346
rect 31852 23192 32928 23194
rect 31846 23132 31852 23192
rect 31912 23134 32928 23192
rect 31912 23132 31918 23134
rect 31344 23084 31406 23090
rect 31344 23024 31346 23084
rect 31344 23018 31406 23024
rect 31344 22989 31404 23018
rect 31130 22983 31618 22989
rect 31130 22949 31142 22983
rect 31606 22949 31618 22983
rect 31130 22943 31618 22949
rect 32148 22983 32636 22989
rect 32148 22949 32160 22983
rect 32624 22949 32636 22983
rect 32148 22943 32636 22949
rect 29864 22314 29870 22822
rect 29824 22302 29870 22314
rect 30834 22314 30848 22890
rect 30882 22314 30894 22890
rect 31860 22890 31906 22902
rect 31860 22390 31866 22890
rect 29298 22261 29358 22264
rect 29094 22255 29582 22261
rect 29094 22221 29106 22255
rect 29570 22221 29582 22255
rect 29094 22215 29582 22221
rect 30112 22255 30600 22261
rect 30112 22221 30124 22255
rect 30588 22221 30600 22255
rect 30112 22215 30600 22221
rect 29298 22026 29358 22215
rect 29298 21960 29358 21966
rect 30326 22026 30386 22215
rect 30326 21960 30386 21966
rect 30834 21918 30894 22314
rect 31848 22314 31866 22390
rect 31900 22390 31906 22890
rect 32878 22890 32924 22902
rect 31900 22314 31908 22390
rect 32878 22386 32884 22890
rect 31346 22261 31406 22264
rect 31130 22255 31618 22261
rect 31130 22221 31142 22255
rect 31606 22221 31618 22255
rect 31130 22215 31618 22221
rect 31346 22026 31406 22215
rect 31848 22164 31908 22314
rect 32868 22314 32884 22386
rect 32918 22386 32924 22890
rect 32918 22314 32928 22386
rect 32148 22255 32636 22261
rect 32148 22221 32160 22255
rect 32624 22221 32636 22255
rect 32148 22215 32636 22221
rect 32336 22164 32396 22215
rect 32868 22164 32928 22314
rect 33010 22164 33070 24068
rect 31846 22160 33070 22164
rect 31842 22100 31848 22160
rect 31908 22104 33070 22160
rect 31908 22100 31914 22104
rect 33798 21968 33804 22028
rect 33864 21968 33870 22028
rect 31346 21960 31406 21966
rect 28796 21858 30894 21918
rect 28796 21528 28856 21858
rect 32658 21742 32664 21802
rect 32724 21742 32730 21802
rect 30104 21558 30110 21622
rect 30174 21558 30180 21622
rect 31128 21558 31134 21622
rect 31198 21558 31204 21622
rect 32140 21558 32146 21622
rect 32210 21558 32216 21622
rect 26042 21436 26048 21500
rect 26112 21436 26118 21500
rect 26766 21468 29160 21528
rect 30110 21504 30174 21558
rect 26046 21385 26110 21436
rect 27078 21385 27138 21468
rect 25832 21379 26320 21385
rect 25832 21345 25844 21379
rect 26308 21345 26320 21379
rect 25832 21339 26320 21345
rect 26850 21379 27338 21385
rect 26850 21345 26862 21379
rect 27326 21345 27338 21379
rect 26850 21339 27338 21345
rect 24566 20710 24578 20734
rect 23796 20651 24284 20657
rect 23796 20617 23808 20651
rect 24272 20617 24284 20651
rect 23796 20611 24284 20617
rect 24012 20556 24072 20611
rect 24518 20556 24578 20710
rect 25538 20710 25550 21286
rect 25584 20710 25598 21286
rect 26562 21286 26608 21298
rect 26562 20788 26568 21286
rect 24814 20651 25302 20657
rect 24814 20617 24826 20651
rect 25290 20617 25302 20651
rect 24814 20611 25302 20617
rect 25022 20556 25082 20611
rect 20446 20356 20506 20492
rect 20954 20438 22020 20498
rect 22476 20492 22482 20552
rect 22542 20492 22548 20552
rect 22818 20494 22824 20554
rect 22884 20494 22890 20554
rect 22992 20496 25082 20556
rect 25538 20554 25598 20710
rect 26556 20710 26568 20788
rect 26602 20788 26608 21286
rect 27572 21286 27632 21468
rect 28100 21385 28160 21468
rect 27868 21379 28356 21385
rect 27868 21345 27880 21379
rect 28344 21345 28356 21379
rect 27868 21339 28356 21345
rect 28100 21338 28160 21339
rect 26602 20710 26616 20788
rect 25832 20651 26320 20657
rect 25832 20617 25844 20651
rect 26308 20617 26320 20651
rect 25832 20611 26320 20617
rect 20440 20296 20446 20356
rect 20506 20296 20512 20356
rect 20954 20250 21014 20438
rect 21460 20298 21466 20358
rect 21526 20298 21532 20358
rect 19426 20186 19432 20246
rect 19492 20186 19498 20246
rect 19916 20190 21014 20250
rect 21466 20246 21526 20298
rect 18706 20123 19194 20129
rect 18706 20089 18718 20123
rect 19182 20089 19194 20123
rect 18706 20083 19194 20089
rect 18418 20030 18464 20042
rect 18418 19490 18424 20030
rect 18414 19454 18424 19490
rect 18458 19490 18464 20030
rect 19432 20030 19492 20186
rect 19916 20129 19976 20190
rect 20954 20129 21014 20190
rect 21460 20186 21466 20246
rect 21526 20186 21532 20246
rect 19724 20123 20212 20129
rect 19724 20089 19736 20123
rect 20200 20089 20212 20123
rect 19724 20083 20212 20089
rect 20742 20123 21230 20129
rect 20742 20089 20754 20123
rect 21218 20089 21230 20123
rect 20742 20083 21230 20089
rect 19432 20004 19442 20030
rect 18458 19454 18474 19490
rect 19436 19478 19442 20004
rect 18414 19296 18474 19454
rect 19430 19454 19442 19478
rect 19476 20004 19492 20030
rect 20454 20030 20500 20042
rect 19476 19478 19482 20004
rect 20454 19480 20460 20030
rect 19476 19454 19490 19478
rect 18706 19395 19194 19401
rect 18706 19361 18718 19395
rect 19182 19361 19194 19395
rect 18706 19355 19194 19361
rect 18928 19296 18988 19355
rect 19430 19296 19490 19454
rect 20448 19454 20460 19480
rect 20494 19480 20500 20030
rect 21466 20030 21526 20186
rect 21960 20129 22020 20438
rect 22824 20240 22884 20494
rect 22482 20180 22884 20240
rect 21760 20123 22248 20129
rect 21760 20089 21772 20123
rect 22236 20089 22248 20123
rect 21760 20083 22248 20089
rect 21466 20008 21478 20030
rect 20494 19454 20508 19480
rect 19910 19401 19970 19402
rect 19724 19395 20212 19401
rect 19724 19361 19736 19395
rect 20200 19361 20212 19395
rect 19724 19355 20212 19361
rect 18414 19236 19490 19296
rect 18414 19082 18474 19236
rect 18408 19022 18414 19082
rect 18474 19022 18480 19082
rect 18412 18912 19488 18972
rect 18412 18774 18472 18912
rect 18926 18873 18986 18912
rect 18706 18867 19194 18873
rect 18706 18833 18718 18867
rect 19182 18833 19194 18867
rect 18706 18827 19194 18833
rect 18412 18740 18424 18774
rect 18418 18198 18424 18740
rect 18458 18740 18472 18774
rect 19428 18774 19488 18912
rect 19910 18873 19970 19355
rect 20448 19192 20508 19454
rect 21472 19454 21478 20008
rect 21512 20008 21526 20030
rect 22482 20030 22542 20180
rect 22778 20123 23266 20129
rect 22778 20089 22790 20123
rect 23254 20089 23266 20123
rect 22778 20083 23266 20089
rect 21512 19454 21518 20008
rect 22482 19972 22496 20030
rect 22490 19484 22496 19972
rect 21472 19442 21518 19454
rect 22484 19454 22496 19484
rect 22530 19972 22542 20030
rect 23498 20030 23558 20496
rect 25532 20494 25538 20554
rect 25598 20494 25604 20554
rect 26556 20358 26616 20710
rect 27572 20710 27586 21286
rect 27620 20710 27632 21286
rect 26850 20651 27338 20657
rect 26850 20617 26862 20651
rect 27326 20617 27338 20651
rect 26850 20611 27338 20617
rect 27066 20556 27126 20611
rect 27572 20556 27632 20710
rect 28588 21286 28648 21468
rect 29100 21385 29160 21468
rect 29604 21440 29610 21500
rect 29670 21440 29676 21500
rect 28886 21379 29374 21385
rect 28886 21345 28898 21379
rect 29362 21345 29374 21379
rect 28886 21339 29374 21345
rect 29100 21332 29160 21339
rect 28588 20710 28604 21286
rect 28638 20710 28648 21286
rect 29610 21286 29670 21440
rect 30110 21385 30174 21440
rect 31134 21385 31198 21558
rect 31638 21440 31644 21500
rect 31704 21440 31710 21500
rect 29904 21379 30392 21385
rect 29904 21345 29916 21379
rect 30380 21345 30392 21379
rect 29904 21339 30392 21345
rect 30922 21379 31410 21385
rect 30922 21345 30934 21379
rect 31398 21345 31410 21379
rect 30922 21339 31410 21345
rect 29610 21258 29622 21286
rect 27868 20651 28356 20657
rect 27868 20617 27880 20651
rect 28344 20617 28356 20651
rect 27868 20611 28356 20617
rect 28092 20556 28152 20611
rect 28588 20556 28648 20710
rect 29616 20710 29622 21258
rect 29656 21258 29670 21286
rect 30634 21286 30680 21298
rect 29656 20710 29662 21258
rect 30634 20734 30640 21286
rect 29616 20698 29662 20710
rect 30626 20710 30640 20734
rect 30674 20734 30680 21286
rect 31644 21286 31704 21440
rect 32146 21385 32210 21558
rect 32664 21504 32724 21742
rect 32664 21444 33740 21504
rect 31940 21379 32428 21385
rect 31940 21345 31952 21379
rect 32416 21345 32428 21379
rect 31940 21339 32428 21345
rect 31644 21262 31658 21286
rect 30674 20710 30686 20734
rect 28886 20651 29374 20657
rect 28886 20617 28898 20651
rect 29362 20617 29374 20651
rect 28886 20611 29374 20617
rect 29904 20651 30392 20657
rect 29904 20617 29916 20651
rect 30380 20617 30392 20651
rect 29904 20611 30392 20617
rect 29104 20556 29164 20611
rect 27066 20496 29164 20556
rect 26550 20298 26556 20358
rect 26616 20298 26622 20358
rect 24516 20184 24522 20244
rect 24582 20184 24588 20244
rect 26550 20184 26556 20244
rect 26616 20184 26622 20244
rect 23796 20123 24284 20129
rect 23796 20089 23808 20123
rect 24272 20089 24284 20123
rect 23796 20083 24284 20089
rect 23498 19986 23514 20030
rect 22530 19484 22536 19972
rect 23508 19484 23514 19986
rect 22530 19454 22544 19484
rect 20948 19401 21008 19402
rect 21954 19401 22014 19402
rect 20742 19395 21230 19401
rect 20742 19361 20754 19395
rect 21218 19361 21230 19395
rect 20742 19355 21230 19361
rect 21760 19395 22248 19401
rect 21760 19361 21772 19395
rect 22236 19361 22248 19395
rect 21760 19355 22248 19361
rect 20448 19126 20508 19132
rect 20442 18928 20448 18988
rect 20508 18928 20514 18988
rect 19724 18867 20212 18873
rect 19724 18833 19736 18867
rect 20200 18833 20212 18867
rect 19724 18827 20212 18833
rect 19428 18752 19442 18774
rect 18458 18198 18464 18740
rect 19436 18226 19442 18752
rect 18418 18186 18464 18198
rect 19430 18198 19442 18226
rect 19476 18752 19488 18774
rect 20448 18774 20508 18928
rect 20948 18873 21008 19355
rect 21954 18873 22014 19355
rect 22484 19192 22544 19454
rect 23500 19454 23514 19484
rect 23548 19986 23558 20030
rect 24522 20030 24582 20184
rect 24814 20123 25302 20129
rect 24814 20089 24826 20123
rect 25290 20089 25302 20123
rect 24814 20083 25302 20089
rect 25832 20123 26320 20129
rect 25832 20089 25844 20123
rect 26308 20089 26320 20123
rect 25832 20083 26320 20089
rect 24522 20002 24532 20030
rect 23548 19484 23554 19986
rect 23548 19454 23560 19484
rect 22778 19395 23266 19401
rect 22778 19361 22790 19395
rect 23254 19361 23266 19395
rect 22778 19355 23266 19361
rect 23004 19300 23064 19355
rect 23500 19300 23560 19454
rect 24526 19454 24532 20002
rect 24566 20002 24582 20030
rect 25544 20030 25590 20042
rect 24566 19454 24572 20002
rect 25544 19478 25550 20030
rect 24526 19442 24572 19454
rect 25538 19454 25550 19478
rect 25584 19478 25590 20030
rect 26556 20030 26616 20184
rect 26850 20123 27338 20129
rect 26850 20089 26862 20123
rect 27326 20089 27338 20123
rect 26850 20083 27338 20089
rect 27868 20123 28356 20129
rect 27868 20089 27880 20123
rect 28344 20089 28356 20123
rect 27868 20083 28356 20089
rect 26556 20000 26568 20030
rect 26562 19482 26568 20000
rect 25584 19454 25598 19478
rect 23796 19395 24284 19401
rect 23796 19361 23808 19395
rect 24272 19361 24284 19395
rect 23796 19355 24284 19361
rect 24814 19395 25302 19401
rect 24814 19361 24826 19395
rect 25290 19361 25302 19395
rect 24814 19355 25302 19361
rect 24016 19300 24076 19355
rect 23004 19240 24076 19300
rect 22478 19132 22484 19192
rect 22544 19132 22550 19192
rect 22476 19030 22482 19090
rect 22542 19030 22548 19090
rect 22482 18988 22542 19030
rect 22476 18928 22482 18988
rect 22542 18928 22548 18988
rect 20742 18867 21230 18873
rect 20742 18833 20754 18867
rect 21218 18833 21230 18867
rect 20742 18827 21230 18833
rect 21760 18867 22248 18873
rect 21760 18833 21772 18867
rect 22236 18833 22248 18867
rect 21760 18827 22248 18833
rect 19476 18226 19482 18752
rect 20448 18750 20460 18774
rect 19476 18198 19490 18226
rect 18706 18139 19194 18145
rect 18706 18105 18718 18139
rect 19182 18105 19194 18139
rect 18706 18099 19194 18105
rect 19430 18040 19490 18198
rect 20454 18198 20460 18750
rect 20494 18750 20508 18774
rect 21472 18774 21518 18786
rect 20494 18198 20500 18750
rect 21472 18222 21478 18774
rect 20454 18186 20500 18198
rect 21466 18198 21478 18222
rect 21512 18222 21518 18774
rect 22482 18774 22542 18928
rect 22778 18867 23266 18873
rect 22778 18833 22790 18867
rect 23254 18833 23266 18867
rect 22778 18827 23266 18833
rect 22482 18746 22496 18774
rect 21512 18198 21526 18222
rect 22490 18217 22496 18746
rect 19922 18145 19982 18152
rect 20960 18145 21020 18152
rect 19724 18139 20212 18145
rect 19724 18105 19736 18139
rect 20200 18105 20212 18139
rect 19724 18099 20212 18105
rect 20742 18139 21230 18145
rect 20742 18105 20754 18139
rect 21218 18105 21230 18139
rect 20742 18099 21230 18105
rect 19424 17980 19430 18040
rect 19490 17980 19496 18040
rect 18256 17772 18262 17832
rect 18322 17772 18328 17832
rect 18412 17674 19488 17734
rect 18412 17518 18472 17674
rect 18926 17617 18986 17674
rect 18706 17611 19194 17617
rect 18706 17577 18718 17611
rect 19182 17577 19194 17611
rect 18706 17571 19194 17577
rect 18412 17480 18424 17518
rect 18418 16942 18424 17480
rect 18458 17480 18472 17518
rect 19428 17518 19488 17674
rect 19922 17617 19982 18099
rect 20438 17670 20444 17730
rect 20504 17670 20510 17730
rect 19724 17611 20212 17617
rect 19724 17577 19736 17611
rect 20200 17577 20212 17611
rect 19724 17571 20212 17577
rect 19428 17492 19442 17518
rect 18458 16942 18464 17480
rect 19436 16968 19442 17492
rect 18418 16930 18464 16942
rect 19426 16942 19442 16968
rect 19476 17492 19488 17518
rect 20444 17518 20504 17670
rect 20960 17617 21020 18099
rect 21466 18040 21526 18198
rect 22484 18198 22496 18217
rect 22530 18746 22542 18774
rect 23500 18774 23560 19240
rect 24512 19236 24518 19296
rect 24578 19236 24584 19296
rect 23796 18867 24284 18873
rect 23796 18833 23808 18867
rect 24272 18833 24284 18867
rect 23796 18827 24284 18833
rect 22530 18217 22536 18746
rect 23500 18736 23514 18774
rect 23508 18232 23514 18736
rect 22530 18198 22544 18217
rect 21966 18145 22026 18152
rect 21760 18139 22248 18145
rect 21760 18105 21772 18139
rect 22236 18105 22248 18139
rect 21760 18099 22248 18105
rect 21460 17980 21466 18040
rect 21526 17980 21532 18040
rect 21466 17932 21526 17980
rect 21460 17872 21466 17932
rect 21526 17872 21532 17932
rect 21966 17882 22026 18099
rect 22484 18048 22544 18198
rect 23498 18198 23514 18232
rect 23548 18736 23560 18774
rect 24518 18774 24578 19236
rect 25020 19134 25080 19355
rect 25538 19296 25598 19454
rect 26556 19454 26568 19482
rect 26602 20000 26616 20030
rect 27580 20030 27626 20042
rect 26602 19482 26608 20000
rect 27580 19482 27586 20030
rect 26602 19454 26616 19482
rect 26050 19401 26110 19408
rect 25832 19395 26320 19401
rect 25832 19361 25844 19395
rect 26308 19361 26320 19395
rect 25832 19355 26320 19361
rect 25532 19236 25538 19296
rect 25598 19236 25604 19296
rect 26050 19134 26110 19355
rect 25020 19074 26110 19134
rect 25020 18873 25080 19074
rect 25532 18930 25538 18990
rect 25598 18930 25604 18990
rect 24814 18867 25302 18873
rect 24814 18833 24826 18867
rect 25290 18833 25302 18867
rect 24814 18827 25302 18833
rect 25020 18822 25080 18827
rect 24518 18750 24532 18774
rect 23548 18232 23554 18736
rect 23548 18198 23558 18232
rect 24526 18228 24532 18750
rect 22778 18139 23266 18145
rect 22778 18105 22790 18139
rect 23254 18105 23266 18139
rect 22778 18099 23266 18105
rect 23002 18048 23062 18099
rect 23498 18048 23558 18198
rect 24520 18198 24532 18228
rect 24566 18750 24578 18774
rect 25538 18774 25598 18930
rect 26050 18873 26110 19074
rect 26556 18990 26616 19454
rect 27574 19454 27586 19482
rect 27620 19482 27626 20030
rect 28588 20030 28648 20496
rect 29606 20184 29612 20244
rect 29672 20184 29678 20244
rect 28886 20123 29374 20129
rect 28886 20089 28898 20123
rect 29362 20089 29374 20123
rect 28886 20083 29374 20089
rect 28588 20010 28604 20030
rect 28598 19482 28604 20010
rect 27620 19454 27634 19482
rect 27062 19401 27122 19408
rect 26850 19395 27338 19401
rect 26850 19361 26862 19395
rect 27326 19361 27338 19395
rect 26850 19355 27338 19361
rect 26550 18930 26556 18990
rect 26616 18930 26622 18990
rect 27062 18873 27122 19355
rect 27574 19296 27634 19454
rect 28588 19454 28604 19482
rect 28638 20010 28648 20030
rect 29612 20030 29672 20184
rect 30112 20129 30172 20611
rect 30626 20552 30686 20710
rect 31652 20710 31658 21262
rect 31692 21262 31704 21286
rect 32664 21286 32724 21444
rect 33178 21385 33238 21444
rect 32958 21379 33446 21385
rect 32958 21345 32970 21379
rect 33434 21345 33446 21379
rect 32958 21339 33446 21345
rect 31692 20710 31698 21262
rect 32664 21250 32676 21286
rect 32670 20738 32676 21250
rect 31652 20698 31698 20710
rect 32662 20710 32676 20738
rect 32710 21250 32724 21286
rect 33680 21286 33740 21444
rect 33680 21262 33694 21286
rect 32710 20738 32716 21250
rect 32710 20710 32722 20738
rect 32142 20657 32202 20663
rect 30922 20651 31410 20657
rect 30922 20617 30934 20651
rect 31398 20617 31410 20651
rect 30922 20611 31410 20617
rect 31940 20651 32428 20657
rect 31940 20617 31952 20651
rect 32416 20617 32428 20651
rect 31940 20611 32428 20617
rect 30620 20492 30626 20552
rect 30686 20492 30692 20552
rect 31136 20129 31196 20611
rect 31640 20184 31646 20244
rect 31706 20184 31712 20244
rect 29904 20123 30392 20129
rect 29904 20089 29916 20123
rect 30380 20089 30392 20123
rect 29904 20083 30392 20089
rect 30922 20123 31410 20129
rect 30922 20089 30934 20123
rect 31398 20089 31410 20123
rect 30922 20083 31410 20089
rect 28638 19482 28644 20010
rect 29612 20002 29622 20030
rect 28638 19454 28648 19482
rect 27868 19395 28356 19401
rect 27868 19361 27880 19395
rect 28344 19361 28356 19395
rect 27868 19355 28356 19361
rect 28092 19298 28152 19355
rect 28588 19298 28648 19454
rect 29616 19454 29622 20002
rect 29656 20002 29672 20030
rect 30634 20030 30680 20042
rect 29656 19454 29662 20002
rect 30634 19490 30640 20030
rect 29616 19442 29662 19454
rect 30624 19454 30640 19490
rect 30674 19490 30680 20030
rect 31646 20030 31706 20184
rect 32142 20129 32202 20611
rect 32662 20552 32722 20710
rect 33688 20710 33694 21262
rect 33728 21262 33740 21286
rect 33728 20710 33734 21262
rect 33688 20698 33734 20710
rect 32958 20651 33446 20657
rect 32958 20617 32970 20651
rect 33434 20617 33446 20651
rect 32958 20611 33446 20617
rect 32656 20492 32662 20552
rect 32722 20492 32728 20552
rect 32664 20190 33740 20250
rect 31940 20123 32428 20129
rect 31940 20089 31952 20123
rect 32416 20089 32428 20123
rect 31940 20083 32428 20089
rect 31646 20006 31658 20030
rect 30674 19454 30684 19490
rect 31652 19482 31658 20006
rect 30106 19401 30166 19402
rect 28886 19395 29374 19401
rect 28886 19361 28898 19395
rect 29362 19361 29374 19395
rect 28886 19355 29374 19361
rect 29904 19395 30392 19401
rect 29904 19361 29916 19395
rect 30380 19361 30392 19395
rect 29904 19355 30392 19361
rect 29104 19298 29164 19355
rect 27568 19236 27574 19296
rect 27634 19236 27640 19296
rect 28092 19238 29164 19298
rect 27566 18930 27572 18990
rect 27632 18930 27638 18990
rect 25832 18867 26320 18873
rect 25832 18833 25844 18867
rect 26308 18833 26320 18867
rect 25832 18827 26320 18833
rect 26850 18867 27338 18873
rect 26850 18833 26862 18867
rect 27326 18833 27338 18867
rect 26850 18827 27338 18833
rect 25538 18752 25550 18774
rect 24566 18228 24572 18750
rect 24566 18198 24580 18228
rect 23796 18139 24284 18145
rect 23796 18105 23808 18139
rect 24272 18105 24284 18139
rect 23796 18099 24284 18105
rect 24014 18048 24074 18099
rect 22478 17988 22484 18048
rect 22544 17988 22550 18048
rect 23002 17988 24074 18048
rect 24280 17988 24286 18048
rect 24346 17988 24352 18048
rect 24520 18042 24580 18198
rect 25544 18198 25550 18752
rect 25584 18752 25598 18774
rect 26562 18774 26608 18786
rect 25584 18198 25590 18752
rect 26562 18224 26568 18774
rect 25544 18186 25590 18198
rect 26556 18198 26568 18224
rect 26602 18224 26608 18774
rect 27572 18774 27632 18930
rect 27868 18867 28356 18873
rect 27868 18833 27880 18867
rect 28344 18833 28356 18867
rect 27868 18827 28356 18833
rect 27572 18748 27586 18774
rect 26602 18198 26616 18224
rect 24814 18139 25302 18145
rect 24814 18105 24826 18139
rect 25290 18105 25302 18139
rect 24814 18099 25302 18105
rect 25832 18139 26320 18145
rect 25832 18105 25844 18139
rect 26308 18105 26320 18139
rect 25832 18099 26320 18105
rect 21966 17822 22742 17882
rect 21966 17617 22026 17822
rect 22472 17670 22478 17730
rect 22538 17670 22544 17730
rect 22682 17718 22742 17822
rect 20742 17611 21230 17617
rect 20742 17577 20754 17611
rect 21218 17577 21230 17611
rect 20742 17571 21230 17577
rect 21760 17611 22248 17617
rect 21760 17577 21772 17611
rect 22236 17577 22248 17611
rect 21760 17571 22248 17577
rect 20444 17492 20460 17518
rect 19476 16968 19482 17492
rect 19476 16942 19486 16968
rect 18706 16883 19194 16889
rect 18706 16849 18718 16883
rect 19182 16849 19194 16883
rect 18706 16843 19194 16849
rect 19426 16782 19486 16942
rect 20454 16942 20460 17492
rect 20494 17492 20504 17518
rect 21472 17518 21518 17530
rect 20494 16942 20500 17492
rect 21472 16964 21478 17518
rect 20454 16930 20500 16942
rect 21462 16942 21478 16964
rect 21512 16964 21518 17518
rect 22478 17518 22538 17670
rect 22676 17658 22682 17718
rect 22742 17658 22748 17718
rect 22778 17611 23266 17617
rect 22778 17577 22790 17611
rect 23254 17577 23266 17611
rect 22778 17571 23266 17577
rect 22478 17488 22496 17518
rect 22490 16978 22496 17488
rect 21512 16942 21522 16964
rect 19724 16883 20212 16889
rect 19724 16849 19736 16883
rect 20200 16849 20212 16883
rect 19724 16843 20212 16849
rect 20742 16883 21230 16889
rect 20742 16849 20754 16883
rect 21218 16849 21230 16883
rect 20742 16843 21230 16849
rect 19420 16722 19426 16782
rect 19486 16722 19492 16782
rect 19934 16668 19994 16843
rect 20958 16668 21018 16843
rect 21462 16782 21522 16942
rect 22484 16942 22496 16978
rect 22530 17488 22538 17518
rect 23498 17518 23558 17988
rect 24286 17778 24346 17988
rect 24514 17982 24520 18042
rect 24580 17982 24586 18042
rect 25016 17920 25076 18099
rect 26044 17920 26104 18099
rect 26556 18042 26616 18198
rect 27580 18198 27586 18748
rect 27620 18748 27632 18774
rect 28588 18774 28648 19238
rect 29602 19132 29608 19192
rect 29668 19132 29674 19192
rect 28886 18867 29374 18873
rect 28886 18833 28898 18867
rect 29362 18833 29374 18867
rect 28886 18827 29374 18833
rect 27620 18198 27626 18748
rect 28588 18744 28604 18774
rect 28598 18230 28604 18744
rect 27580 18186 27626 18198
rect 28586 18198 28604 18230
rect 28638 18744 28648 18774
rect 29608 18774 29668 19132
rect 30106 18873 30166 19355
rect 30470 19250 30476 19310
rect 30536 19250 30542 19310
rect 30476 18990 30536 19250
rect 30624 19200 30684 19454
rect 31644 19454 31658 19482
rect 31692 20006 31706 20030
rect 32664 20030 32724 20190
rect 33178 20129 33238 20190
rect 32958 20123 33446 20129
rect 32958 20089 32970 20123
rect 33434 20089 33446 20123
rect 32958 20083 33446 20089
rect 31692 19482 31698 20006
rect 32664 19996 32676 20030
rect 32670 19494 32676 19996
rect 31692 19454 31704 19482
rect 31130 19401 31190 19402
rect 30922 19395 31410 19401
rect 30922 19361 30934 19395
rect 31398 19361 31410 19395
rect 30922 19355 31410 19361
rect 30618 19140 30624 19200
rect 30684 19140 30690 19200
rect 30470 18930 30476 18990
rect 30536 18930 30542 18990
rect 30622 18932 30628 18992
rect 30688 18932 30694 18992
rect 29904 18867 30392 18873
rect 29904 18833 29916 18867
rect 30380 18833 30392 18867
rect 29904 18827 30392 18833
rect 28638 18230 28644 18744
rect 29608 18742 29622 18774
rect 29616 18230 29622 18742
rect 28638 18198 28646 18230
rect 26850 18139 27338 18145
rect 26850 18105 26862 18139
rect 27326 18105 27338 18139
rect 26850 18099 27338 18105
rect 27868 18139 28356 18145
rect 27868 18105 27880 18139
rect 28344 18105 28356 18139
rect 27868 18099 28356 18105
rect 26550 17982 26556 18042
rect 26616 17982 26622 18042
rect 25016 17860 26104 17920
rect 26548 17872 26554 17932
rect 26614 17872 26620 17932
rect 24286 17718 25594 17778
rect 23796 17611 24284 17617
rect 23796 17577 23808 17611
rect 24272 17577 24284 17611
rect 23796 17571 24284 17577
rect 24814 17611 25302 17617
rect 24814 17577 24826 17611
rect 25290 17577 25302 17611
rect 24814 17571 25302 17577
rect 22530 16978 22536 17488
rect 23498 17460 23514 17518
rect 22530 16942 22544 16978
rect 23508 16974 23514 17460
rect 21760 16883 22248 16889
rect 21760 16849 21772 16883
rect 22236 16849 22248 16883
rect 21760 16843 22248 16849
rect 21456 16722 21462 16782
rect 21522 16722 21528 16782
rect 21964 16668 22024 16843
rect 18124 16592 18130 16652
rect 18190 16592 18196 16652
rect 19934 16608 22024 16668
rect 12484 16464 12490 16524
rect 12550 16464 13286 16524
rect 13346 16522 17808 16524
rect 13346 16464 15638 16522
rect 13286 16458 13346 16464
rect 15632 16462 15638 16464
rect 15698 16464 17808 16522
rect 15698 16462 15704 16464
rect 13166 16406 13226 16412
rect 18130 16406 18190 16592
rect 13226 16346 18190 16406
rect 13166 16340 13226 16346
rect 12720 16288 12780 16294
rect 19934 16288 19994 16608
rect 21964 16398 22024 16608
rect 22484 16512 22544 16942
rect 23498 16942 23514 16974
rect 23548 17460 23558 17518
rect 24526 17518 24572 17530
rect 23548 16974 23554 17460
rect 24526 16986 24532 17518
rect 23548 16942 23558 16974
rect 22778 16883 23266 16889
rect 22778 16849 22790 16883
rect 23254 16849 23266 16883
rect 22778 16843 23266 16849
rect 23002 16788 23062 16843
rect 23498 16788 23558 16942
rect 24520 16942 24532 16986
rect 24566 16986 24572 17518
rect 25534 17518 25594 17718
rect 26044 17718 26104 17860
rect 26044 17617 26104 17658
rect 25832 17611 26320 17617
rect 25832 17577 25844 17611
rect 26308 17577 26320 17611
rect 25832 17571 26320 17577
rect 25534 17466 25550 17518
rect 24566 16942 24580 16986
rect 23796 16883 24284 16889
rect 23796 16849 23808 16883
rect 24272 16849 24284 16883
rect 23796 16843 24284 16849
rect 24014 16788 24074 16843
rect 24520 16788 24580 16942
rect 25544 16942 25550 17466
rect 25584 17466 25594 17518
rect 26554 17518 26614 17872
rect 27060 17718 27120 18099
rect 28090 18046 28150 18099
rect 28586 18046 28646 18198
rect 29610 18198 29622 18230
rect 29656 18742 29668 18774
rect 30628 18774 30688 18932
rect 31130 18873 31190 19355
rect 31644 19090 31704 19454
rect 32664 19454 32676 19494
rect 32710 19996 32724 20030
rect 33680 20030 33740 20190
rect 33680 20008 33694 20030
rect 32710 19494 32716 19996
rect 32710 19454 32724 19494
rect 32136 19401 32196 19408
rect 31940 19395 32428 19401
rect 31940 19361 31952 19395
rect 32416 19361 32428 19395
rect 31940 19355 32428 19361
rect 31638 19030 31644 19090
rect 31704 19030 31710 19090
rect 32136 18873 32196 19355
rect 32664 19200 32724 19454
rect 33688 19454 33694 20008
rect 33728 20008 33740 20030
rect 33728 19454 33734 20008
rect 33688 19442 33734 19454
rect 32958 19395 33446 19401
rect 32958 19361 32970 19395
rect 33434 19361 33446 19395
rect 32958 19355 33446 19361
rect 33804 19200 33864 21968
rect 33946 21800 34006 24516
rect 34234 22100 34240 22160
rect 34300 22100 34306 22160
rect 33946 21734 34006 21740
rect 34082 21440 34088 21500
rect 34148 21440 34154 21500
rect 33922 20298 33928 20358
rect 33988 20298 33994 20358
rect 32658 19140 32664 19200
rect 32724 19140 32730 19200
rect 33798 19140 33804 19200
rect 33864 19140 33870 19200
rect 32656 18932 32662 18992
rect 32722 18932 32728 18992
rect 30922 18867 31410 18873
rect 30922 18833 30934 18867
rect 31398 18833 31410 18867
rect 30922 18827 31410 18833
rect 31940 18867 32428 18873
rect 31940 18833 31952 18867
rect 32416 18833 32428 18867
rect 31940 18827 32428 18833
rect 30628 18754 30640 18774
rect 29656 18230 29662 18742
rect 29656 18198 29670 18230
rect 28886 18139 29374 18145
rect 28886 18105 28898 18139
rect 29362 18105 29374 18139
rect 28886 18099 29374 18105
rect 29102 18046 29162 18099
rect 28090 17986 29162 18046
rect 29610 18044 29670 18198
rect 30634 18198 30640 18754
rect 30674 18754 30688 18774
rect 31652 18774 31698 18786
rect 30674 18198 30680 18754
rect 31652 18226 31658 18774
rect 30634 18186 30680 18198
rect 31646 18198 31658 18226
rect 31692 18226 31698 18774
rect 32662 18774 32722 18932
rect 32958 18867 33446 18873
rect 32958 18833 32970 18867
rect 33434 18833 33446 18867
rect 32958 18827 33446 18833
rect 32662 18750 32676 18774
rect 32670 18234 32676 18750
rect 31692 18198 31706 18226
rect 30118 18145 30178 18152
rect 31142 18145 31202 18152
rect 29904 18139 30392 18145
rect 29904 18105 29916 18139
rect 30380 18105 30392 18139
rect 29904 18099 30392 18105
rect 30922 18139 31410 18145
rect 30922 18105 30934 18139
rect 31398 18105 31410 18139
rect 30922 18099 31410 18105
rect 27060 17652 27120 17658
rect 26850 17611 27338 17617
rect 26850 17577 26862 17611
rect 27326 17577 27338 17611
rect 26850 17571 27338 17577
rect 27868 17611 28356 17617
rect 27868 17577 27880 17611
rect 28344 17577 28356 17611
rect 27868 17571 28356 17577
rect 25584 16942 25590 17466
rect 26554 17454 26568 17518
rect 25544 16930 25590 16942
rect 26562 16942 26568 17454
rect 26602 17454 26614 17518
rect 27580 17518 27626 17530
rect 26602 16942 26608 17454
rect 27580 16970 27586 17518
rect 26562 16930 26608 16942
rect 27572 16942 27586 16970
rect 27620 16970 27626 17518
rect 28586 17518 28646 17986
rect 29604 17984 29610 18044
rect 29670 17984 29676 18044
rect 30118 17724 30178 18099
rect 30118 17718 30180 17724
rect 30118 17658 30120 17718
rect 30626 17670 30632 17730
rect 30692 17670 30698 17730
rect 30118 17652 30180 17658
rect 30118 17617 30178 17652
rect 28886 17611 29374 17617
rect 28886 17577 28898 17611
rect 29362 17577 29374 17611
rect 28886 17571 29374 17577
rect 29904 17611 30392 17617
rect 29904 17577 29916 17611
rect 30380 17577 30392 17611
rect 29904 17571 30392 17577
rect 28586 17480 28604 17518
rect 28598 16972 28604 17480
rect 27620 16942 27632 16970
rect 24814 16883 25302 16889
rect 24814 16849 24826 16883
rect 25290 16849 25302 16883
rect 24814 16843 25302 16849
rect 25832 16883 26320 16889
rect 25832 16849 25844 16883
rect 26308 16849 26320 16883
rect 25832 16843 26320 16849
rect 26850 16883 27338 16889
rect 26850 16849 26862 16883
rect 27326 16849 27338 16883
rect 26850 16843 27338 16849
rect 25030 16788 25090 16843
rect 27056 16788 27116 16843
rect 27572 16788 27632 16942
rect 28586 16942 28604 16972
rect 28638 17480 28646 17518
rect 29616 17518 29662 17530
rect 28638 16972 28644 17480
rect 28638 16942 28646 16972
rect 29616 16968 29622 17518
rect 27868 16883 28356 16889
rect 27868 16849 27880 16883
rect 28344 16849 28356 16883
rect 27868 16843 28356 16849
rect 28090 16788 28150 16843
rect 28586 16788 28646 16942
rect 29614 16942 29622 16968
rect 29656 16968 29662 17518
rect 30632 17518 30692 17670
rect 31142 17617 31202 18099
rect 31646 18044 31706 18198
rect 32662 18198 32676 18234
rect 32710 18750 32722 18774
rect 33688 18774 33734 18786
rect 32710 18234 32716 18750
rect 32710 18198 32722 18234
rect 33688 18222 33694 18774
rect 32148 18145 32208 18158
rect 31940 18139 32428 18145
rect 31940 18105 31952 18139
rect 32416 18105 32428 18139
rect 31940 18099 32428 18105
rect 31640 17984 31646 18044
rect 31706 17984 31712 18044
rect 32148 17617 32208 18099
rect 32662 18040 32722 18198
rect 33678 18198 33694 18222
rect 33728 18222 33734 18774
rect 33728 18198 33738 18222
rect 32958 18139 33446 18145
rect 32958 18105 32970 18139
rect 33434 18105 33446 18139
rect 32958 18099 33446 18105
rect 33176 18040 33236 18099
rect 33678 18040 33738 18198
rect 32662 17980 33738 18040
rect 33804 17932 33864 19140
rect 33928 18992 33988 20298
rect 33922 18932 33928 18992
rect 33988 18932 33994 18992
rect 33798 17872 33804 17932
rect 33864 17872 33870 17932
rect 32660 17670 32666 17730
rect 32726 17670 32732 17730
rect 30922 17611 31410 17617
rect 30922 17577 30934 17611
rect 31398 17577 31410 17611
rect 30922 17571 31410 17577
rect 31940 17611 32428 17617
rect 31940 17577 31952 17611
rect 32416 17577 32428 17611
rect 31940 17571 32428 17577
rect 30632 17492 30640 17518
rect 29656 16942 29674 16968
rect 28886 16883 29374 16889
rect 28886 16849 28898 16883
rect 29362 16849 29374 16883
rect 28886 16843 29374 16849
rect 29102 16788 29162 16843
rect 23002 16728 29162 16788
rect 29614 16782 29674 16942
rect 30634 16942 30640 17492
rect 30674 17492 30692 17518
rect 31652 17518 31698 17530
rect 30674 16942 30680 17492
rect 31652 16964 31658 17518
rect 30634 16930 30680 16942
rect 31650 16942 31658 16964
rect 31692 16964 31698 17518
rect 32666 17518 32726 17670
rect 32958 17611 33446 17617
rect 32958 17577 32970 17611
rect 33434 17577 33446 17611
rect 32958 17571 33446 17577
rect 32666 17488 32676 17518
rect 32670 16980 32676 17488
rect 31692 16942 31710 16964
rect 30122 16889 30182 16896
rect 29904 16883 30392 16889
rect 29904 16849 29916 16883
rect 30380 16849 30392 16883
rect 29904 16843 30392 16849
rect 30922 16883 31410 16889
rect 30922 16849 30934 16883
rect 31398 16849 31410 16883
rect 30922 16843 31410 16849
rect 29608 16722 29614 16782
rect 29674 16722 29680 16782
rect 30122 16670 30182 16843
rect 31142 16670 31202 16843
rect 31650 16782 31710 16942
rect 32664 16942 32676 16980
rect 32710 17488 32726 17518
rect 33688 17518 33734 17530
rect 32710 16980 32716 17488
rect 32710 16942 32724 16980
rect 33688 16968 33694 17518
rect 31940 16883 32428 16889
rect 31940 16849 31952 16883
rect 32416 16849 32428 16883
rect 31940 16843 32428 16849
rect 31644 16722 31650 16782
rect 31710 16722 31716 16782
rect 32144 16670 32204 16843
rect 32664 16786 32724 16942
rect 33680 16942 33694 16968
rect 33728 16968 33734 17518
rect 33728 16942 33740 16968
rect 32958 16883 33446 16889
rect 32958 16849 32970 16883
rect 33434 16849 33446 16883
rect 32958 16843 33446 16849
rect 33178 16786 33238 16843
rect 33680 16786 33740 16942
rect 32664 16726 33740 16786
rect 30122 16610 32204 16670
rect 22478 16452 22484 16512
rect 22544 16452 22550 16512
rect 30122 16398 30182 16610
rect 34088 16512 34148 21440
rect 34240 20244 34300 22100
rect 34234 20184 34240 20244
rect 34300 20184 34306 20244
rect 35666 16642 35672 30072
rect 35772 16642 35778 30072
rect 34082 16452 34088 16512
rect 34148 16452 34154 16512
rect 21964 16338 30182 16398
rect 12780 16228 19994 16288
rect 12720 16222 12780 16228
rect 35666 16128 35778 16642
rect 52322 30692 76778 30698
rect 52322 30592 52428 30692
rect 76672 30592 76778 30692
rect 52322 30586 76778 30592
rect 52322 30072 52434 30586
rect 53034 30286 53044 30586
rect 76056 30286 76066 30586
rect 52322 16642 52328 30072
rect 52428 16642 52434 30072
rect 55948 30204 72828 30236
rect 55948 29990 56011 30204
rect 72796 29990 72828 30204
rect 55948 29968 55998 29990
rect 56058 29968 56434 29990
rect 56494 29968 56872 29990
rect 56932 29968 57306 29990
rect 57366 29970 72828 29990
rect 76666 30072 76778 30586
rect 57366 29968 60302 29970
rect 60462 28494 60522 29970
rect 62498 28494 62558 29970
rect 63002 28494 63062 29970
rect 63510 28494 63570 29970
rect 64022 28494 64082 29970
rect 64536 28494 64596 29970
rect 66568 28494 66628 29970
rect 68608 28494 68668 29970
rect 69098 28494 69158 29970
rect 69618 28494 69678 29970
rect 70126 28494 70186 29970
rect 70640 28494 70700 29970
rect 72676 28494 72736 29970
rect 60462 28434 72736 28494
rect 59930 28228 59936 28288
rect 59996 28228 60002 28288
rect 58424 28012 59502 28072
rect 58424 27832 58484 28012
rect 58928 27931 58988 28012
rect 58720 27925 59208 27931
rect 58720 27891 58732 27925
rect 59196 27891 59208 27925
rect 58720 27885 59208 27891
rect 58424 27792 58438 27832
rect 58432 27256 58438 27792
rect 58472 27792 58484 27832
rect 59442 27832 59502 28012
rect 59936 27931 59996 28228
rect 60462 28042 60522 28434
rect 61012 28228 61018 28288
rect 61078 28228 61084 28288
rect 61970 28228 61976 28288
rect 62036 28228 62042 28288
rect 60456 27982 60462 28042
rect 60522 27982 60528 28042
rect 59738 27925 60226 27931
rect 59738 27891 59750 27925
rect 60214 27891 60226 27925
rect 59738 27885 60226 27891
rect 59442 27806 59456 27832
rect 58472 27256 58478 27792
rect 59450 27292 59456 27806
rect 58432 27244 58478 27256
rect 59444 27256 59456 27292
rect 59490 27806 59502 27832
rect 60462 27832 60522 27982
rect 61018 27931 61078 28228
rect 61976 27931 62036 28228
rect 62498 28042 62558 28434
rect 62492 27982 62498 28042
rect 62558 27982 62564 28042
rect 60756 27925 61244 27931
rect 60756 27891 60768 27925
rect 61232 27891 61244 27925
rect 60756 27885 61244 27891
rect 61774 27925 62262 27931
rect 61774 27891 61786 27925
rect 62250 27891 62262 27925
rect 61774 27885 62262 27891
rect 61976 27882 62036 27885
rect 60462 27808 60474 27832
rect 59490 27292 59496 27806
rect 60468 27296 60474 27808
rect 59490 27256 59504 27292
rect 58720 27197 59208 27203
rect 58720 27163 58732 27197
rect 59196 27163 59208 27197
rect 58720 27157 59208 27163
rect 59444 27110 59504 27256
rect 60464 27256 60474 27296
rect 60508 27808 60522 27832
rect 61486 27832 61532 27844
rect 60508 27296 60514 27808
rect 60508 27256 60524 27296
rect 61486 27284 61492 27832
rect 59948 27203 60008 27204
rect 59738 27197 60226 27203
rect 59738 27163 59750 27197
rect 60214 27163 60226 27197
rect 59738 27157 60226 27163
rect 58274 27050 58280 27110
rect 58340 27050 58346 27110
rect 59438 27050 59444 27110
rect 59504 27050 59510 27110
rect 58144 26846 58150 26906
rect 58210 26846 58216 26906
rect 56136 24662 56142 24722
rect 56202 24662 56208 24722
rect 53964 21346 55186 21406
rect 53964 19430 54024 21346
rect 54106 21182 54166 21346
rect 54618 21281 54678 21346
rect 54402 21275 54890 21281
rect 54402 21241 54414 21275
rect 54878 21241 54890 21275
rect 54402 21235 54890 21241
rect 54106 21132 54120 21182
rect 54114 20606 54120 21132
rect 54154 21132 54166 21182
rect 55126 21182 55186 21346
rect 55420 21275 55908 21281
rect 55420 21241 55432 21275
rect 55896 21241 55908 21275
rect 55420 21235 55908 21241
rect 54154 20606 54160 21132
rect 55126 21130 55138 21182
rect 54114 20594 54160 20606
rect 55132 20606 55138 21130
rect 55172 21130 55186 21182
rect 56142 21182 56202 24662
rect 58150 24290 58210 26846
rect 58280 24436 58340 27050
rect 59438 26846 59444 26906
rect 59504 26846 59510 26906
rect 58720 26789 59208 26795
rect 58720 26755 58732 26789
rect 59196 26755 59208 26789
rect 58720 26749 59208 26755
rect 58432 26696 58478 26708
rect 58432 26156 58438 26696
rect 58426 26120 58438 26156
rect 58472 26156 58478 26696
rect 59444 26696 59504 26846
rect 59948 26795 60008 27157
rect 59738 26789 60226 26795
rect 59738 26755 59750 26789
rect 60214 26755 60226 26789
rect 59738 26749 60226 26755
rect 59948 26746 60008 26749
rect 59444 26658 59456 26696
rect 58472 26120 58486 26156
rect 59450 26150 59456 26658
rect 58426 25970 58486 26120
rect 59444 26120 59456 26150
rect 59490 26658 59504 26696
rect 60464 26696 60524 27256
rect 61480 27256 61492 27284
rect 61526 27284 61532 27832
rect 62498 27832 62558 27982
rect 63002 27931 63062 28434
rect 62792 27925 63280 27931
rect 62792 27891 62804 27925
rect 63268 27891 63280 27925
rect 62792 27885 63280 27891
rect 62498 27808 62510 27832
rect 62504 27314 62510 27808
rect 61526 27256 61540 27284
rect 60756 27197 61244 27203
rect 60756 27163 60768 27197
rect 61232 27163 61244 27197
rect 60756 27157 61244 27163
rect 61480 27006 61540 27256
rect 62488 27256 62510 27314
rect 62544 27808 62558 27832
rect 63510 27832 63570 28434
rect 64022 27931 64082 28434
rect 64536 28044 64596 28434
rect 65034 28228 65040 28288
rect 65100 28228 65106 28288
rect 66052 28228 66058 28288
rect 66118 28228 66124 28288
rect 64530 27984 64536 28044
rect 64596 27984 64602 28044
rect 63810 27925 64298 27931
rect 63810 27891 63822 27925
rect 64286 27891 64298 27925
rect 63810 27885 64298 27891
rect 62544 27314 62550 27808
rect 63510 27762 63528 27832
rect 62544 27256 62552 27314
rect 61774 27197 62262 27203
rect 61774 27163 61786 27197
rect 62250 27163 62262 27197
rect 61774 27157 62262 27163
rect 61474 26946 61480 27006
rect 61540 26946 61546 27006
rect 60756 26789 61244 26795
rect 60756 26755 60768 26789
rect 61232 26755 61244 26789
rect 60756 26749 61244 26755
rect 61774 26789 62262 26795
rect 61774 26755 61786 26789
rect 62250 26755 62262 26789
rect 61774 26749 62262 26755
rect 59490 26150 59496 26658
rect 60464 26656 60474 26696
rect 59490 26120 59504 26150
rect 60468 26146 60474 26656
rect 58720 26061 59208 26067
rect 58720 26027 58732 26061
rect 59196 26027 59208 26061
rect 58720 26021 59208 26027
rect 58938 25970 58998 26021
rect 59444 25970 59504 26120
rect 60460 26120 60474 26146
rect 60508 26656 60524 26696
rect 61486 26696 61532 26708
rect 60508 26146 60514 26656
rect 60508 26120 60520 26146
rect 61486 26140 61492 26696
rect 59930 26067 59990 26074
rect 59738 26061 60226 26067
rect 59738 26027 59750 26061
rect 60214 26027 60226 26061
rect 59738 26021 60226 26027
rect 58426 25910 59504 25970
rect 59438 25766 59498 25768
rect 58428 25706 59498 25766
rect 58428 25560 58488 25706
rect 58938 25659 58998 25706
rect 58720 25653 59208 25659
rect 58720 25619 58732 25653
rect 59196 25619 59208 25653
rect 58720 25613 59208 25619
rect 58428 25528 58438 25560
rect 58432 24984 58438 25528
rect 58472 25528 58488 25560
rect 59438 25560 59498 25706
rect 59930 25756 59990 26021
rect 59930 25659 59990 25696
rect 60460 25974 60520 26120
rect 61478 26120 61492 26140
rect 61526 26140 61532 26696
rect 62488 26696 62552 27256
rect 63522 27256 63528 27762
rect 63562 27762 63570 27832
rect 64536 27832 64596 27984
rect 65040 27931 65100 28228
rect 66058 27931 66118 28228
rect 66568 28044 66628 28434
rect 67076 28228 67082 28288
rect 67142 28228 67148 28288
rect 68088 28228 68094 28288
rect 68154 28228 68160 28288
rect 66560 27984 66566 28044
rect 66626 27984 66632 28044
rect 64828 27925 65316 27931
rect 64828 27891 64840 27925
rect 65304 27891 65316 27925
rect 64828 27885 65316 27891
rect 65846 27925 66334 27931
rect 65846 27891 65858 27925
rect 66322 27891 66334 27925
rect 65846 27885 66334 27891
rect 64536 27792 64546 27832
rect 63562 27256 63568 27762
rect 64540 27310 64546 27792
rect 63522 27244 63568 27256
rect 64524 27256 64546 27310
rect 64580 27792 64596 27832
rect 65558 27832 65604 27844
rect 64580 27310 64586 27792
rect 64580 27256 64588 27310
rect 65558 27296 65564 27832
rect 62792 27197 63280 27203
rect 62792 27163 62804 27197
rect 63268 27163 63280 27197
rect 62792 27157 63280 27163
rect 63810 27197 64298 27203
rect 63810 27163 63822 27197
rect 64286 27163 64298 27197
rect 63810 27157 64298 27163
rect 63510 26946 63516 27006
rect 63576 26946 63582 27006
rect 62792 26789 63280 26795
rect 62792 26755 62804 26789
rect 63268 26755 63280 26789
rect 62792 26749 63280 26755
rect 62488 26666 62510 26696
rect 62504 26148 62510 26666
rect 61526 26120 61538 26140
rect 60958 26067 61018 26068
rect 60756 26061 61244 26067
rect 60756 26027 60768 26061
rect 61232 26027 61244 26061
rect 60756 26021 61244 26027
rect 60958 25974 61018 26021
rect 61478 25974 61538 26120
rect 62496 26120 62510 26148
rect 62544 26666 62552 26696
rect 63516 26696 63576 26946
rect 63810 26789 64298 26795
rect 63810 26755 63822 26789
rect 64286 26755 64298 26789
rect 63810 26749 64298 26755
rect 62544 26148 62550 26666
rect 63516 26658 63528 26696
rect 63522 26156 63528 26658
rect 62544 26146 62556 26148
rect 62544 26120 62560 26146
rect 61986 26067 62046 26072
rect 61774 26061 62262 26067
rect 61774 26027 61786 26061
rect 62250 26027 62262 26061
rect 61774 26021 62262 26027
rect 61986 25974 62046 26021
rect 60460 25972 62046 25974
rect 62496 25972 62560 26120
rect 63514 26120 63528 26156
rect 63562 26658 63576 26696
rect 64524 26696 64588 27256
rect 65554 27256 65564 27296
rect 65598 27296 65604 27832
rect 66568 27832 66628 27984
rect 67082 27931 67142 28228
rect 68094 27931 68154 28228
rect 68608 28046 68668 28434
rect 68602 27986 68608 28046
rect 68668 27986 68674 28046
rect 66864 27925 67352 27931
rect 66864 27891 66876 27925
rect 67340 27891 67352 27925
rect 66864 27885 67352 27891
rect 67882 27925 68370 27931
rect 67882 27891 67894 27925
rect 68358 27891 68370 27925
rect 67882 27885 68370 27891
rect 66568 27792 66582 27832
rect 66576 27312 66582 27792
rect 65598 27256 65614 27296
rect 65042 27203 65102 27206
rect 64828 27197 65316 27203
rect 64828 27163 64840 27197
rect 65304 27163 65316 27197
rect 64828 27157 65316 27163
rect 65042 26795 65102 27157
rect 65554 27110 65614 27256
rect 66566 27256 66582 27312
rect 66616 27792 66628 27832
rect 67594 27832 67640 27844
rect 66616 27312 66622 27792
rect 66616 27256 66630 27312
rect 67594 27294 67600 27832
rect 66060 27203 66120 27212
rect 65846 27197 66334 27203
rect 65846 27163 65858 27197
rect 66322 27163 66334 27197
rect 65846 27157 66334 27163
rect 65548 27050 65554 27110
rect 65614 27050 65620 27110
rect 65544 26846 65550 26906
rect 65610 26846 65616 26906
rect 64828 26789 65316 26795
rect 64828 26755 64840 26789
rect 65304 26755 65316 26789
rect 64828 26749 65316 26755
rect 65042 26748 65102 26749
rect 64524 26662 64546 26696
rect 63562 26156 63568 26658
rect 64540 26156 64546 26662
rect 63562 26120 63578 26156
rect 62792 26061 63280 26067
rect 62792 26027 62804 26061
rect 63268 26027 63280 26061
rect 62792 26021 63280 26027
rect 60460 25914 61986 25972
rect 59738 25653 60226 25659
rect 59738 25619 59750 25653
rect 60214 25619 60226 25653
rect 59738 25613 60226 25619
rect 59438 25528 59456 25560
rect 58472 24984 58478 25528
rect 59450 25026 59456 25528
rect 58432 24972 58478 24984
rect 59438 24984 59456 25026
rect 59490 25528 59498 25560
rect 60460 25560 60520 25914
rect 62490 25912 62496 25972
rect 62556 25912 62562 25972
rect 61986 25906 62046 25912
rect 61472 25810 61478 25874
rect 61542 25810 61548 25874
rect 60962 25696 60968 25756
rect 61028 25696 61034 25756
rect 61478 25716 61542 25810
rect 60968 25659 61028 25696
rect 60756 25653 61244 25659
rect 60756 25619 60768 25653
rect 61232 25619 61244 25653
rect 60756 25613 61244 25619
rect 59490 25026 59496 25528
rect 60460 25508 60474 25560
rect 59490 24984 59502 25026
rect 60468 25020 60474 25508
rect 58720 24925 59208 24931
rect 58720 24891 58732 24925
rect 59196 24891 59208 24925
rect 58720 24885 59208 24891
rect 59438 24776 59502 24984
rect 60460 24984 60474 25020
rect 60508 25508 60520 25560
rect 61478 25560 61544 25716
rect 61974 25696 61980 25756
rect 62040 25696 62046 25756
rect 61980 25659 62040 25696
rect 61774 25653 62262 25659
rect 61774 25619 61786 25653
rect 62250 25619 62262 25653
rect 61774 25613 62262 25619
rect 61980 25612 62040 25613
rect 61478 25510 61492 25560
rect 60508 25020 60514 25508
rect 60508 24984 60520 25020
rect 61486 25008 61492 25510
rect 59738 24925 60226 24931
rect 59738 24891 59750 24925
rect 60214 24891 60226 24925
rect 59738 24885 60226 24891
rect 58994 24716 59502 24776
rect 58274 24376 58280 24436
rect 58340 24376 58346 24436
rect 58150 24230 58570 24290
rect 58510 21418 58570 24230
rect 58630 21968 58636 22028
rect 58696 21968 58702 22028
rect 57160 21350 58370 21410
rect 58504 21358 58510 21418
rect 58570 21358 58576 21418
rect 56438 21275 56926 21281
rect 56438 21241 56450 21275
rect 56914 21241 56926 21275
rect 56438 21235 56926 21241
rect 55172 20606 55178 21130
rect 55132 20594 55178 20606
rect 56142 20606 56156 21182
rect 56190 20606 56202 21182
rect 57160 21182 57220 21350
rect 57672 21281 57732 21350
rect 57456 21275 57944 21281
rect 57456 21241 57468 21275
rect 57932 21241 57944 21275
rect 57456 21235 57944 21241
rect 57160 21134 57174 21182
rect 54402 20547 54890 20553
rect 54402 20513 54414 20547
rect 54878 20513 54890 20547
rect 54402 20507 54890 20513
rect 55420 20547 55908 20553
rect 55420 20513 55432 20547
rect 55896 20513 55908 20547
rect 55420 20507 55908 20513
rect 55626 20464 55686 20507
rect 55620 20404 55626 20464
rect 55686 20404 55692 20464
rect 55728 20292 55734 20352
rect 55794 20292 55800 20352
rect 55734 20249 55794 20292
rect 54402 20243 54890 20249
rect 54402 20209 54414 20243
rect 54878 20209 54890 20243
rect 54402 20203 54890 20209
rect 55420 20243 55908 20249
rect 55420 20209 55432 20243
rect 55896 20209 55908 20243
rect 55420 20203 55908 20209
rect 54114 20150 54160 20162
rect 54114 19632 54120 20150
rect 54104 19574 54120 19632
rect 54154 19632 54160 20150
rect 55132 20150 55178 20162
rect 54154 19574 54164 19632
rect 55132 19624 55138 20150
rect 53958 19370 53964 19430
rect 54024 19370 54030 19430
rect 53838 18342 53898 18348
rect 53964 18342 54024 19370
rect 54104 19320 54164 19574
rect 55124 19574 55138 19624
rect 55172 19624 55178 20150
rect 56142 20150 56202 20606
rect 57168 20606 57174 21134
rect 57208 21134 57220 21182
rect 58178 21182 58238 21350
rect 58178 21136 58192 21182
rect 57208 20606 57214 21134
rect 57168 20594 57214 20606
rect 58186 20606 58192 21136
rect 58226 21136 58238 21182
rect 58226 20606 58232 21136
rect 58186 20594 58232 20606
rect 56438 20547 56926 20553
rect 56438 20513 56450 20547
rect 56914 20513 56926 20547
rect 56438 20507 56926 20513
rect 57456 20547 57944 20553
rect 57456 20513 57468 20547
rect 57932 20513 57944 20547
rect 57456 20507 57944 20513
rect 56518 20352 56578 20507
rect 56642 20404 56648 20464
rect 56708 20404 56714 20464
rect 56512 20292 56518 20352
rect 56578 20292 56584 20352
rect 56648 20249 56708 20404
rect 56438 20243 56926 20249
rect 56438 20209 56450 20243
rect 56914 20209 56926 20243
rect 56438 20203 56926 20209
rect 57456 20243 57944 20249
rect 57456 20209 57468 20243
rect 57932 20209 57944 20243
rect 57456 20203 57944 20209
rect 55172 19574 55184 19624
rect 54402 19515 54890 19521
rect 54402 19481 54414 19515
rect 54878 19481 54890 19515
rect 54402 19475 54890 19481
rect 54606 19320 54666 19475
rect 55124 19320 55184 19574
rect 56142 19574 56156 20150
rect 56190 19574 56202 20150
rect 57168 20150 57214 20162
rect 57168 19660 57174 20150
rect 55420 19515 55908 19521
rect 55420 19481 55432 19515
rect 55896 19481 55908 19515
rect 55420 19475 55908 19481
rect 54104 19260 55124 19320
rect 55184 19260 55190 19320
rect 54104 19118 54164 19260
rect 54606 19217 54666 19260
rect 54402 19211 54890 19217
rect 54402 19177 54414 19211
rect 54878 19177 54890 19211
rect 54402 19171 54890 19177
rect 54104 19058 54120 19118
rect 54114 18542 54120 19058
rect 54154 19058 54164 19118
rect 55124 19118 55184 19260
rect 55634 19217 55694 19475
rect 55420 19211 55908 19217
rect 55420 19177 55432 19211
rect 55896 19177 55908 19211
rect 55420 19171 55908 19177
rect 54154 18542 54160 19058
rect 55124 19054 55138 19118
rect 54114 18530 54160 18542
rect 55132 18542 55138 19054
rect 55172 19054 55184 19118
rect 56142 19118 56202 19574
rect 57158 19574 57174 19660
rect 57208 19660 57214 20150
rect 58186 20150 58232 20162
rect 57208 19574 57218 19660
rect 58186 19620 58192 20150
rect 56438 19515 56926 19521
rect 56438 19481 56450 19515
rect 56914 19481 56926 19515
rect 56438 19475 56926 19481
rect 56652 19217 56712 19475
rect 57158 19430 57218 19574
rect 58178 19574 58192 19620
rect 58226 19620 58232 20150
rect 58226 19574 58238 19620
rect 57456 19515 57944 19521
rect 57456 19481 57468 19515
rect 57932 19481 57944 19515
rect 57456 19475 57944 19481
rect 57672 19430 57732 19475
rect 58178 19430 58238 19574
rect 57152 19370 57158 19430
rect 57218 19370 58238 19430
rect 56438 19211 56926 19217
rect 56438 19177 56450 19211
rect 56914 19177 56926 19211
rect 56438 19171 56926 19177
rect 55172 18542 55178 19054
rect 55132 18530 55178 18542
rect 56142 18542 56156 19118
rect 56190 18542 56202 19118
rect 57158 19118 57218 19370
rect 57672 19217 57732 19370
rect 57456 19211 57944 19217
rect 57456 19177 57468 19211
rect 57932 19177 57944 19211
rect 57456 19171 57944 19177
rect 57158 19062 57174 19118
rect 54402 18483 54890 18489
rect 54402 18449 54414 18483
rect 54878 18449 54890 18483
rect 54402 18443 54890 18449
rect 55420 18483 55908 18489
rect 55420 18449 55432 18483
rect 55896 18449 55908 18483
rect 55420 18443 55908 18449
rect 55640 18396 55700 18443
rect 53898 18282 55188 18342
rect 55634 18336 55640 18396
rect 55700 18336 55706 18396
rect 53838 18276 53898 18282
rect 54102 18086 54162 18282
rect 54610 18185 54670 18282
rect 54402 18179 54890 18185
rect 54402 18145 54414 18179
rect 54878 18145 54890 18179
rect 54402 18139 54890 18145
rect 54102 18034 54120 18086
rect 54114 17510 54120 18034
rect 54154 18034 54162 18086
rect 55128 18086 55188 18282
rect 55740 18236 55746 18296
rect 55806 18236 55812 18296
rect 55746 18185 55806 18236
rect 55420 18179 55908 18185
rect 55420 18145 55432 18179
rect 55896 18145 55908 18179
rect 55420 18139 55908 18145
rect 55128 18038 55138 18086
rect 54154 17510 54160 18034
rect 54114 17498 54160 17510
rect 55132 17510 55138 18038
rect 55172 18038 55188 18086
rect 56142 18086 56202 18542
rect 57168 18542 57174 19062
rect 57208 19062 57218 19118
rect 58178 19118 58238 19370
rect 58310 19320 58370 21350
rect 58304 19260 58310 19320
rect 58370 19260 58376 19320
rect 58178 19082 58192 19118
rect 57208 18542 57214 19062
rect 57168 18530 57214 18542
rect 58186 18542 58192 19082
rect 58226 19082 58238 19118
rect 58226 18542 58232 19082
rect 58186 18530 58232 18542
rect 56438 18483 56926 18489
rect 56438 18449 56450 18483
rect 56914 18449 56926 18483
rect 56438 18443 56926 18449
rect 57456 18483 57944 18489
rect 57456 18449 57468 18483
rect 57932 18449 57944 18483
rect 57456 18443 57944 18449
rect 56532 18296 56592 18443
rect 56644 18336 56650 18396
rect 56710 18336 56716 18396
rect 58310 18342 58370 19260
rect 58496 19132 58502 19192
rect 58562 19132 58568 19192
rect 56526 18236 56532 18296
rect 56592 18236 56598 18296
rect 56650 18185 56710 18336
rect 57158 18282 58370 18342
rect 56438 18179 56926 18185
rect 56438 18145 56450 18179
rect 56914 18145 56926 18179
rect 56438 18139 56926 18145
rect 55172 17510 55178 18038
rect 56142 18012 56156 18086
rect 55132 17498 55178 17510
rect 56150 17510 56156 18012
rect 56190 18012 56202 18086
rect 57158 18086 57218 18282
rect 57660 18185 57720 18282
rect 57456 18179 57944 18185
rect 57456 18145 57468 18179
rect 57932 18145 57944 18179
rect 57456 18139 57944 18145
rect 57158 18056 57174 18086
rect 56190 17510 56196 18012
rect 57168 17592 57174 18056
rect 56150 17498 56196 17510
rect 57160 17510 57174 17592
rect 57208 18056 57218 18086
rect 58178 18086 58238 18282
rect 57208 17592 57214 18056
rect 58178 18018 58192 18086
rect 57208 17510 57220 17592
rect 56638 17457 56698 17461
rect 54402 17451 54890 17457
rect 54402 17417 54414 17451
rect 54878 17417 54890 17451
rect 54402 17411 54890 17417
rect 55420 17451 55908 17457
rect 55420 17417 55432 17451
rect 55896 17417 55908 17451
rect 55420 17411 55908 17417
rect 56438 17451 56926 17457
rect 56438 17417 56450 17451
rect 56914 17417 56926 17451
rect 56438 17411 56926 17417
rect 53352 17286 53412 17292
rect 55632 17286 55692 17411
rect 53412 17226 55692 17286
rect 53352 17220 53412 17226
rect 53492 17110 53552 17116
rect 56638 17110 56698 17411
rect 53552 17050 56698 17110
rect 53492 17044 53552 17050
rect 54392 16936 54452 16942
rect 57160 16936 57220 17510
rect 58186 17510 58192 18018
rect 58226 18018 58238 18086
rect 58226 17510 58232 18018
rect 58186 17498 58232 17510
rect 57456 17451 57944 17457
rect 57456 17417 57468 17451
rect 57932 17417 57944 17451
rect 57456 17411 57944 17417
rect 54452 16876 57220 16936
rect 54392 16870 54452 16876
rect 53232 16786 53292 16792
rect 58502 16786 58562 19132
rect 58636 18040 58696 21968
rect 58746 21358 58752 21418
rect 58812 21358 58818 21418
rect 58752 19296 58812 21358
rect 58994 20454 59054 24716
rect 59438 24586 59502 24716
rect 59432 24522 59438 24586
rect 59502 24522 59508 24586
rect 59262 24436 59322 24442
rect 59262 21500 59322 24376
rect 59940 24330 60000 24885
rect 60460 24834 60520 24984
rect 61476 24984 61492 25008
rect 61526 25514 61544 25560
rect 62496 25560 62560 25912
rect 62990 25764 63050 26021
rect 63514 25874 63578 26120
rect 64530 26120 64546 26156
rect 64580 26662 64588 26696
rect 65550 26696 65610 26846
rect 66060 26795 66120 27157
rect 65846 26789 66334 26795
rect 65846 26755 65858 26789
rect 66322 26755 66334 26789
rect 65846 26749 66334 26755
rect 65550 26670 65564 26696
rect 64580 26156 64586 26662
rect 64580 26154 64590 26156
rect 64580 26120 64594 26154
rect 63810 26061 64298 26067
rect 63810 26027 63822 26061
rect 64286 26027 64298 26061
rect 63810 26021 64298 26027
rect 63348 25810 63354 25874
rect 63418 25810 63578 25874
rect 64014 25764 64074 26021
rect 64530 25972 64594 26120
rect 65558 26120 65564 26670
rect 65598 26670 65610 26696
rect 66566 26696 66630 27256
rect 67588 27256 67600 27294
rect 67634 27294 67640 27832
rect 68608 27832 68668 27986
rect 69098 27931 69158 28434
rect 69618 28046 69678 28434
rect 69612 27986 69618 28046
rect 69678 27986 69684 28046
rect 68900 27925 69388 27931
rect 68900 27891 68912 27925
rect 69376 27891 69388 27925
rect 68900 27885 69388 27891
rect 68608 27794 68618 27832
rect 68612 27296 68618 27794
rect 67634 27256 67648 27294
rect 67076 27203 67136 27209
rect 66864 27197 67352 27203
rect 66864 27163 66876 27197
rect 67340 27163 67352 27197
rect 66864 27157 67352 27163
rect 67076 26795 67136 27157
rect 67588 27110 67648 27256
rect 68604 27256 68618 27296
rect 68652 27794 68668 27832
rect 69618 27832 69678 27986
rect 70126 27931 70186 28434
rect 70640 28046 70700 28434
rect 71146 28228 71152 28288
rect 71212 28228 71218 28288
rect 72158 28228 72164 28288
rect 72224 28228 72230 28288
rect 70634 27986 70640 28046
rect 70700 27986 70706 28046
rect 69918 27925 70406 27931
rect 69918 27891 69930 27925
rect 70394 27891 70406 27925
rect 69918 27885 70406 27891
rect 70126 27882 70186 27885
rect 68652 27296 68658 27794
rect 69618 27762 69636 27832
rect 68652 27256 68668 27296
rect 68088 27203 68148 27209
rect 67882 27197 68370 27203
rect 67882 27163 67894 27197
rect 68358 27163 68370 27197
rect 67882 27157 68370 27163
rect 67582 27050 67588 27110
rect 67648 27050 67654 27110
rect 68088 26906 68148 27157
rect 67580 26846 67586 26906
rect 67646 26846 67652 26906
rect 68082 26846 68088 26906
rect 68148 26846 68154 26906
rect 66864 26789 67352 26795
rect 66864 26755 66876 26789
rect 67340 26755 67352 26789
rect 66864 26749 67352 26755
rect 67076 26746 67136 26749
rect 65598 26120 65604 26670
rect 66566 26664 66582 26696
rect 66576 26168 66582 26664
rect 65558 26108 65604 26120
rect 66568 26120 66582 26168
rect 66616 26664 66630 26696
rect 67586 26696 67646 26846
rect 68088 26795 68148 26846
rect 67882 26789 68370 26795
rect 67882 26755 67894 26789
rect 68358 26755 68370 26789
rect 67882 26749 68370 26755
rect 68088 26746 68148 26749
rect 67586 26664 67600 26696
rect 66616 26168 66622 26664
rect 66616 26166 66628 26168
rect 66616 26120 66632 26166
rect 67594 26150 67600 26664
rect 65042 26067 65102 26074
rect 64828 26061 65316 26067
rect 64828 26027 64840 26061
rect 65304 26027 65316 26061
rect 64828 26021 65316 26027
rect 65846 26061 66334 26067
rect 65846 26027 65858 26061
rect 66322 26027 66334 26061
rect 65846 26021 66334 26027
rect 64524 25912 64530 25972
rect 64590 25912 64596 25972
rect 62984 25704 62990 25764
rect 63050 25704 63056 25764
rect 64008 25704 64014 25764
rect 64074 25704 64080 25764
rect 62792 25653 63280 25659
rect 62792 25619 62804 25653
rect 63268 25619 63280 25653
rect 62792 25613 63280 25619
rect 63810 25653 64298 25659
rect 63810 25619 63822 25653
rect 64286 25619 64298 25653
rect 63810 25613 64298 25619
rect 61526 25510 61542 25514
rect 62496 25512 62510 25560
rect 61526 25008 61532 25510
rect 62504 25010 62510 25512
rect 61526 24984 61540 25008
rect 60756 24925 61244 24931
rect 60756 24891 60768 24925
rect 61232 24891 61244 24925
rect 60756 24885 61244 24891
rect 60454 24774 60460 24834
rect 60520 24774 60526 24834
rect 60982 24330 61042 24885
rect 61476 24724 61540 24984
rect 62496 24984 62510 25010
rect 62544 25512 62560 25560
rect 63522 25560 63568 25572
rect 62544 25010 62550 25512
rect 63522 25040 63528 25560
rect 62544 25008 62556 25010
rect 62544 24984 62560 25008
rect 61774 24925 62262 24931
rect 61774 24891 61786 24925
rect 62250 24891 62262 24925
rect 61774 24885 62262 24891
rect 61470 24660 61476 24724
rect 61540 24660 61546 24724
rect 61982 24330 62042 24885
rect 62496 24834 62560 24984
rect 63516 24984 63528 25040
rect 63562 25040 63568 25560
rect 64530 25560 64594 25912
rect 65042 25764 65102 26021
rect 65036 25704 65042 25764
rect 65102 25704 65108 25764
rect 65042 25659 65102 25704
rect 66070 25659 66130 26021
rect 66568 25970 66632 26120
rect 67588 26120 67600 26150
rect 67634 26664 67646 26696
rect 68604 26696 68668 27256
rect 69630 27256 69636 27762
rect 69670 27762 69678 27832
rect 70640 27832 70700 27986
rect 71152 27931 71212 28228
rect 72164 27931 72224 28228
rect 72676 28046 72736 28434
rect 73176 28228 73182 28288
rect 73242 28228 73248 28288
rect 72670 27986 72676 28046
rect 72736 27986 72742 28046
rect 70936 27925 71424 27931
rect 70936 27891 70948 27925
rect 71412 27891 71424 27925
rect 70936 27885 71424 27891
rect 71954 27925 72442 27931
rect 71954 27891 71966 27925
rect 72430 27891 72442 27925
rect 71954 27885 72442 27891
rect 70640 27804 70654 27832
rect 69670 27256 69676 27762
rect 70648 27304 70654 27804
rect 69630 27244 69676 27256
rect 70640 27256 70654 27304
rect 70688 27804 70700 27832
rect 71666 27832 71712 27844
rect 70688 27304 70694 27804
rect 70688 27256 70700 27304
rect 71666 27288 71672 27832
rect 68900 27197 69388 27203
rect 68900 27163 68912 27197
rect 69376 27163 69388 27197
rect 68900 27157 69388 27163
rect 69918 27197 70406 27203
rect 69918 27163 69930 27197
rect 70394 27163 70406 27197
rect 69918 27157 70406 27163
rect 69616 26946 69622 27006
rect 69682 26946 69688 27006
rect 69102 26846 69108 26906
rect 69168 26846 69174 26906
rect 69108 26795 69168 26846
rect 68900 26789 69388 26795
rect 68900 26755 68912 26789
rect 69376 26755 69388 26789
rect 68900 26749 69388 26755
rect 67634 26150 67640 26664
rect 68604 26648 68618 26696
rect 68612 26164 68618 26648
rect 67634 26120 67648 26150
rect 67088 26067 67148 26079
rect 66864 26061 67352 26067
rect 66864 26027 66876 26061
rect 67340 26027 67352 26061
rect 66864 26021 67352 26027
rect 66562 25910 66568 25970
rect 66628 25910 66634 25970
rect 64828 25653 65316 25659
rect 64828 25619 64840 25653
rect 65304 25619 65316 25653
rect 64828 25613 65316 25619
rect 65846 25653 66334 25659
rect 65846 25619 65858 25653
rect 66322 25619 66334 25653
rect 65846 25613 66334 25619
rect 66070 25606 66130 25613
rect 64530 25500 64546 25560
rect 63562 24984 63576 25040
rect 64540 25018 64546 25500
rect 63018 24931 63078 24934
rect 62792 24925 63280 24931
rect 62792 24891 62804 24925
rect 63268 24891 63280 24925
rect 62792 24885 63280 24891
rect 63018 24834 63078 24885
rect 63516 24834 63576 24984
rect 64530 24984 64546 25018
rect 64580 25500 64594 25560
rect 65558 25560 65604 25572
rect 64580 25018 64586 25500
rect 64580 25016 64590 25018
rect 65558 25016 65564 25560
rect 64580 24984 64594 25016
rect 63810 24925 64298 24931
rect 63810 24891 63822 24925
rect 64286 24891 64298 24925
rect 63810 24885 64298 24891
rect 62490 24774 62496 24834
rect 62556 24774 62562 24834
rect 63012 24774 63018 24834
rect 63078 24774 63084 24834
rect 63510 24774 63516 24834
rect 63576 24774 63582 24834
rect 63990 24830 64050 24885
rect 64530 24838 64594 24984
rect 65548 24984 65564 25016
rect 65598 25016 65604 25560
rect 66568 25560 66632 25910
rect 67088 25659 67148 26021
rect 67588 25872 67648 26120
rect 68604 26120 68618 26164
rect 68652 26648 68668 26696
rect 69622 26696 69682 26946
rect 70128 26846 70134 26906
rect 70194 26846 70200 26906
rect 70640 26902 70700 27256
rect 71656 27256 71672 27288
rect 71706 27288 71712 27832
rect 72676 27832 72736 27986
rect 73182 27931 73242 28228
rect 73696 27994 74776 28054
rect 72972 27925 73460 27931
rect 72972 27891 72984 27925
rect 73448 27891 73460 27925
rect 72972 27885 73460 27891
rect 72676 27800 72690 27832
rect 72684 27294 72690 27800
rect 71706 27256 71716 27288
rect 70936 27197 71424 27203
rect 70936 27163 70948 27197
rect 71412 27163 71424 27197
rect 70936 27157 71424 27163
rect 71656 27006 71716 27256
rect 72680 27256 72690 27294
rect 72724 27800 72736 27832
rect 73696 27832 73756 27994
rect 74198 27931 74258 27994
rect 73990 27925 74478 27931
rect 73990 27891 74002 27925
rect 74466 27891 74478 27925
rect 73990 27885 74478 27891
rect 73696 27802 73708 27832
rect 72724 27294 72730 27800
rect 73702 27296 73708 27802
rect 72724 27256 72740 27294
rect 71954 27197 72442 27203
rect 71954 27163 71966 27197
rect 72430 27163 72442 27197
rect 71954 27157 72442 27163
rect 71650 26946 71656 27006
rect 71716 26946 71722 27006
rect 72680 26908 72740 27256
rect 73696 27256 73708 27296
rect 73742 27802 73756 27832
rect 74716 27832 74776 27994
rect 73742 27296 73748 27802
rect 74716 27786 74726 27832
rect 73742 27256 73756 27296
rect 73160 27203 73220 27215
rect 72972 27197 73460 27203
rect 72972 27163 72984 27197
rect 73448 27163 73460 27197
rect 72972 27157 73460 27163
rect 72680 26902 72744 26908
rect 70134 26795 70194 26846
rect 70634 26842 70640 26902
rect 70700 26842 70706 26902
rect 71148 26842 71154 26902
rect 71214 26842 71220 26902
rect 71652 26842 71658 26902
rect 71718 26842 71724 26902
rect 72158 26842 72164 26902
rect 72224 26842 72230 26902
rect 72680 26842 72684 26902
rect 69918 26789 70406 26795
rect 69918 26755 69930 26789
rect 70394 26755 70406 26789
rect 69918 26749 70406 26755
rect 69622 26672 69636 26696
rect 68652 26164 68658 26648
rect 68652 26162 68664 26164
rect 68652 26120 68668 26162
rect 68088 26067 68148 26075
rect 67882 26061 68370 26067
rect 67882 26027 67894 26061
rect 68358 26027 68370 26061
rect 67882 26021 68370 26027
rect 67582 25812 67588 25872
rect 67648 25812 67654 25872
rect 68088 25659 68148 26021
rect 68604 25970 68668 26120
rect 69630 26120 69636 26672
rect 69670 26672 69682 26696
rect 70640 26696 70700 26842
rect 71154 26795 71214 26842
rect 70936 26789 71424 26795
rect 70936 26755 70948 26789
rect 71412 26755 71424 26789
rect 70936 26749 71424 26755
rect 69670 26120 69676 26672
rect 70640 26652 70654 26696
rect 70648 26156 70654 26652
rect 69630 26108 69676 26120
rect 70640 26120 70654 26156
rect 70688 26652 70700 26696
rect 71658 26696 71718 26842
rect 72164 26795 72224 26842
rect 72680 26836 72744 26842
rect 71954 26789 72442 26795
rect 71954 26755 71966 26789
rect 72430 26755 72442 26789
rect 71954 26749 72442 26755
rect 71658 26668 71672 26696
rect 70688 26156 70694 26652
rect 71666 26190 71672 26668
rect 70688 26120 70700 26156
rect 68900 26061 69388 26067
rect 68900 26027 68912 26061
rect 69376 26027 69388 26061
rect 68900 26021 69388 26027
rect 69918 26061 70406 26067
rect 69918 26027 69930 26061
rect 70394 26027 70406 26061
rect 69918 26021 70406 26027
rect 70640 25970 70700 26120
rect 71656 26120 71672 26190
rect 71706 26668 71718 26696
rect 72680 26696 72740 26836
rect 73160 26795 73220 27157
rect 73696 27110 73756 27256
rect 74720 27256 74726 27786
rect 74760 27786 74776 27832
rect 74760 27256 74766 27786
rect 74720 27244 74766 27256
rect 73990 27197 74478 27203
rect 73990 27163 74002 27197
rect 74466 27163 74478 27197
rect 73990 27157 74478 27163
rect 73690 27050 73696 27110
rect 73756 27050 73762 27110
rect 74940 27050 74946 27110
rect 75006 27050 75012 27110
rect 73700 26834 74770 26894
rect 72972 26789 73460 26795
rect 72972 26755 72984 26789
rect 73448 26755 73460 26789
rect 72972 26749 73460 26755
rect 71706 26190 71712 26668
rect 72680 26660 72690 26696
rect 71706 26120 71716 26190
rect 72684 26152 72690 26660
rect 70936 26061 71424 26067
rect 70936 26027 70948 26061
rect 71412 26027 71424 26061
rect 70936 26021 71424 26027
rect 71142 25970 71202 26021
rect 68598 25910 68604 25970
rect 68664 25910 68670 25970
rect 69098 25910 69104 25970
rect 69164 25910 69170 25970
rect 69612 25910 69618 25970
rect 69678 25910 69684 25970
rect 70136 25910 70142 25970
rect 70202 25910 70208 25970
rect 70634 25910 70640 25970
rect 70700 25910 70706 25970
rect 71136 25910 71142 25970
rect 71202 25910 71208 25970
rect 71656 25968 71716 26120
rect 72674 26120 72690 26152
rect 72724 26660 72740 26696
rect 73700 26696 73760 26834
rect 74206 26795 74266 26834
rect 73990 26789 74478 26795
rect 73990 26755 74002 26789
rect 74466 26755 74478 26789
rect 73990 26749 74478 26755
rect 73700 26668 73708 26696
rect 72724 26152 72730 26660
rect 72724 26150 72734 26152
rect 73702 26150 73708 26668
rect 72724 26120 72738 26150
rect 72164 26067 72224 26074
rect 71954 26061 72442 26067
rect 71954 26027 71966 26061
rect 72430 26027 72442 26061
rect 71954 26021 72442 26027
rect 72164 25968 72224 26021
rect 72674 25968 72738 26120
rect 73696 26120 73708 26150
rect 73742 26668 73760 26696
rect 74710 26696 74770 26834
rect 73742 26150 73748 26668
rect 74710 26662 74726 26696
rect 73742 26120 73756 26150
rect 73160 26067 73220 26073
rect 72972 26061 73460 26067
rect 72972 26027 72984 26061
rect 73448 26027 73460 26061
rect 72972 26021 73460 26027
rect 66864 25653 67352 25659
rect 66864 25619 66876 25653
rect 67340 25619 67352 25653
rect 66864 25613 67352 25619
rect 67882 25653 68370 25659
rect 67882 25619 67894 25653
rect 68358 25619 68370 25653
rect 67882 25613 68370 25619
rect 68088 25612 68148 25613
rect 66568 25520 66582 25560
rect 66576 25044 66582 25520
rect 65598 24984 65612 25016
rect 64828 24925 65316 24931
rect 64828 24891 64840 24925
rect 65304 24891 65316 24925
rect 64828 24885 65316 24891
rect 59372 24270 59378 24330
rect 59438 24270 59444 24330
rect 59934 24270 59940 24330
rect 60000 24270 60006 24330
rect 60976 24270 60982 24330
rect 61042 24270 61048 24330
rect 61976 24270 61982 24330
rect 62042 24270 62048 24330
rect 59378 21688 59438 24270
rect 63990 24232 64050 24770
rect 64498 24834 64594 24838
rect 64498 24832 64530 24834
rect 64590 24774 64596 24834
rect 64984 24774 64990 24834
rect 65050 24774 65056 24834
rect 64498 24232 64558 24772
rect 64990 24232 65050 24774
rect 65144 24330 65204 24885
rect 65548 24582 65612 24984
rect 66566 24984 66582 25044
rect 66616 25520 66632 25560
rect 67594 25560 67640 25572
rect 66616 25044 66622 25520
rect 66616 24984 66626 25044
rect 67594 25020 67600 25560
rect 65846 24925 66334 24931
rect 65846 24891 65858 24925
rect 66322 24891 66334 24925
rect 65846 24885 66334 24891
rect 65548 24512 65612 24518
rect 66034 24836 66094 24842
rect 65138 24270 65144 24330
rect 65204 24270 65210 24330
rect 66034 24232 66094 24776
rect 66154 24330 66214 24885
rect 66566 24834 66626 24984
rect 67584 24984 67600 25020
rect 67634 25020 67640 25560
rect 68604 25560 68668 25910
rect 69104 25659 69164 25910
rect 68900 25653 69388 25659
rect 68900 25619 68912 25653
rect 69376 25619 69388 25653
rect 68900 25613 69388 25619
rect 68604 25508 68618 25560
rect 68612 25026 68618 25508
rect 67634 24984 67648 25020
rect 66864 24925 67352 24931
rect 66864 24891 66876 24925
rect 67340 24891 67352 24925
rect 66864 24885 67352 24891
rect 66560 24774 66566 24834
rect 66626 24774 66632 24834
rect 67096 24330 67156 24885
rect 67584 24440 67648 24984
rect 68604 24984 68618 25026
rect 68652 25508 68668 25560
rect 69618 25560 69678 25910
rect 70142 25659 70202 25910
rect 69918 25653 70406 25659
rect 69918 25619 69930 25653
rect 70394 25619 70406 25653
rect 69918 25613 70406 25619
rect 68652 25026 68658 25508
rect 69618 25506 69636 25560
rect 69630 25430 69636 25506
rect 68652 25024 68664 25026
rect 68652 24984 68668 25024
rect 67882 24925 68370 24931
rect 67882 24891 67894 24925
rect 68358 24891 68370 24925
rect 67882 24885 68370 24891
rect 68078 24836 68138 24842
rect 68604 24836 68668 24984
rect 69622 24984 69636 25430
rect 69670 25506 69678 25560
rect 70640 25560 70700 25910
rect 71650 25908 71656 25968
rect 71716 25908 71722 25968
rect 72158 25908 72164 25968
rect 72224 25908 72230 25968
rect 72668 25908 72674 25968
rect 72734 25908 72740 25968
rect 71140 25696 71146 25756
rect 71206 25696 71212 25756
rect 72152 25696 72158 25756
rect 72218 25696 72224 25756
rect 71146 25659 71206 25696
rect 72158 25659 72218 25696
rect 70936 25653 71424 25659
rect 70936 25619 70948 25653
rect 71412 25619 71424 25653
rect 70936 25613 71424 25619
rect 71954 25653 72442 25659
rect 71954 25619 71966 25653
rect 72430 25619 72442 25653
rect 71954 25613 72442 25619
rect 70640 25506 70654 25560
rect 69670 25430 69676 25506
rect 69670 24984 69682 25430
rect 70648 25014 70654 25506
rect 69100 24931 69160 24940
rect 68900 24925 69388 24931
rect 68900 24891 68912 24925
rect 69376 24891 69388 24925
rect 68900 24885 69388 24891
rect 67578 24376 67584 24440
rect 67648 24376 67654 24440
rect 66148 24270 66154 24330
rect 66214 24270 66220 24330
rect 67090 24270 67096 24330
rect 67156 24270 67162 24330
rect 68078 24232 68138 24776
rect 68572 24832 68668 24836
rect 68572 24830 68604 24832
rect 68664 24772 68670 24832
rect 69100 24826 69160 24885
rect 69622 24836 69682 24984
rect 70640 24984 70654 25014
rect 70688 25506 70700 25560
rect 71666 25560 71712 25572
rect 70688 25014 70694 25506
rect 71666 25018 71672 25560
rect 70688 25012 70700 25014
rect 70688 24984 70704 25012
rect 70100 24931 70160 24934
rect 69918 24925 70406 24931
rect 69918 24891 69930 24925
rect 70394 24891 70406 24925
rect 69918 24885 70406 24891
rect 68572 24232 68632 24770
rect 69100 24232 69160 24766
rect 69588 24830 69682 24836
rect 69648 24828 69682 24830
rect 69588 24768 69622 24770
rect 69588 24762 69682 24768
rect 70100 24826 70160 24885
rect 70640 24830 70704 24984
rect 71656 24984 71672 25018
rect 71706 25018 71712 25560
rect 72674 25560 72738 25908
rect 73160 25756 73220 26021
rect 73696 25872 73756 26120
rect 74720 26120 74726 26662
rect 74760 26662 74770 26696
rect 74760 26120 74766 26662
rect 74720 26108 74766 26120
rect 73990 26061 74478 26067
rect 73990 26027 74002 26061
rect 74466 26027 74478 26061
rect 73990 26021 74478 26027
rect 73690 25812 73696 25872
rect 73756 25812 73762 25872
rect 73698 25758 73758 25760
rect 73154 25696 73160 25756
rect 73220 25696 73226 25756
rect 73698 25698 74770 25758
rect 73160 25659 73220 25696
rect 72972 25653 73460 25659
rect 72972 25619 72984 25653
rect 73448 25619 73460 25653
rect 72972 25613 73460 25619
rect 73160 25610 73220 25613
rect 72674 25514 72690 25560
rect 71706 24984 71720 25018
rect 72684 25014 72690 25514
rect 70936 24925 71424 24931
rect 70936 24891 70948 24925
rect 71412 24891 71424 24925
rect 70936 24885 71424 24891
rect 70634 24770 70640 24830
rect 70700 24770 70706 24830
rect 69588 24232 69648 24762
rect 70100 24232 70160 24766
rect 71656 24724 71720 24984
rect 72674 24984 72690 25014
rect 72724 25514 72738 25560
rect 73698 25560 73758 25698
rect 74202 25659 74262 25698
rect 73990 25653 74478 25659
rect 73990 25619 74002 25653
rect 74466 25619 74478 25653
rect 73990 25613 74478 25619
rect 73698 25534 73708 25560
rect 72724 25014 72730 25514
rect 73702 25072 73708 25534
rect 72724 25012 72734 25014
rect 72724 24984 72738 25012
rect 71954 24925 72442 24931
rect 71954 24891 71966 24925
rect 72430 24891 72442 24925
rect 71954 24885 72442 24891
rect 72674 24830 72738 24984
rect 73690 24984 73708 25072
rect 73742 25534 73758 25560
rect 74710 25560 74770 25698
rect 73742 25072 73748 25534
rect 74710 25510 74726 25560
rect 73742 24984 73750 25072
rect 72972 24925 73460 24931
rect 72972 24891 72984 24925
rect 73448 24891 73460 24925
rect 72972 24885 73460 24891
rect 72668 24770 72674 24830
rect 72734 24770 72740 24830
rect 71650 24660 71656 24724
rect 71720 24660 71726 24724
rect 73690 24436 73750 24984
rect 74720 24984 74726 25510
rect 74760 25510 74770 25560
rect 74760 24984 74766 25510
rect 74720 24972 74766 24984
rect 73990 24925 74478 24931
rect 73990 24891 74002 24925
rect 74466 24891 74478 24925
rect 73990 24885 74478 24891
rect 74946 24592 75006 27050
rect 74942 24586 75006 24592
rect 74942 24516 75006 24522
rect 73684 24376 73690 24436
rect 73750 24376 73756 24436
rect 61654 24172 71894 24232
rect 59486 24068 59492 24128
rect 59552 24068 59558 24128
rect 59492 22154 59552 24068
rect 59914 24015 60402 24021
rect 59914 23981 59926 24015
rect 60390 23981 60402 24015
rect 59914 23975 60402 23981
rect 60932 24015 61420 24021
rect 60932 23981 60944 24015
rect 61408 23981 61420 24015
rect 60932 23975 61420 23981
rect 59626 23922 59672 23934
rect 59626 23376 59632 23922
rect 59618 23346 59632 23376
rect 59666 23376 59672 23922
rect 60644 23922 60690 23934
rect 59666 23346 59678 23376
rect 60644 23370 60650 23922
rect 59618 23194 59678 23346
rect 60636 23346 60650 23370
rect 60684 23370 60690 23922
rect 61654 23922 61714 24172
rect 62664 24068 62670 24128
rect 62730 24068 62736 24128
rect 61950 24015 62438 24021
rect 61950 23981 61962 24015
rect 62426 23981 62438 24015
rect 61950 23975 62438 23981
rect 60684 23346 60696 23370
rect 59914 23287 60402 23293
rect 59914 23253 59926 23287
rect 60390 23253 60402 23287
rect 59914 23247 60402 23253
rect 60130 23194 60190 23247
rect 60636 23194 60696 23346
rect 61654 23346 61668 23922
rect 61702 23346 61714 23922
rect 62670 23922 62730 24068
rect 62968 24015 63456 24021
rect 62968 23981 62980 24015
rect 63444 23981 63456 24015
rect 62968 23975 63456 23981
rect 62670 23858 62686 23922
rect 60932 23287 61420 23293
rect 60932 23253 60944 23287
rect 61408 23253 61420 23287
rect 60932 23247 61420 23253
rect 59618 23192 60696 23194
rect 59618 23134 60636 23192
rect 60630 23132 60636 23134
rect 60696 23132 60702 23192
rect 61140 23084 61200 23247
rect 61134 23024 61140 23084
rect 61200 23024 61206 23084
rect 61140 22989 61200 23024
rect 59914 22983 60402 22989
rect 59914 22949 59926 22983
rect 60390 22949 60402 22983
rect 59914 22943 60402 22949
rect 60932 22983 61420 22989
rect 60932 22949 60944 22983
rect 61408 22949 61420 22983
rect 60932 22943 61420 22949
rect 59626 22890 59672 22902
rect 59626 22370 59632 22890
rect 59618 22314 59632 22370
rect 59666 22370 59672 22890
rect 60644 22890 60690 22902
rect 59666 22314 59678 22370
rect 60644 22344 60650 22890
rect 59618 22154 59678 22314
rect 60632 22314 60650 22344
rect 60684 22344 60690 22890
rect 61654 22890 61714 23346
rect 62680 23346 62686 23858
rect 62720 23858 62730 23922
rect 63692 23922 63752 24172
rect 63986 24015 64474 24021
rect 63986 23981 63998 24015
rect 64462 23981 64474 24015
rect 63986 23975 64474 23981
rect 65004 24015 65492 24021
rect 65004 23981 65016 24015
rect 65480 23981 65492 24015
rect 65004 23975 65492 23981
rect 62720 23346 62726 23858
rect 62680 23334 62726 23346
rect 63692 23346 63704 23922
rect 63738 23346 63752 23922
rect 64716 23922 64762 23934
rect 64716 23410 64722 23922
rect 62160 23293 62220 23299
rect 61950 23287 62438 23293
rect 61950 23253 61962 23287
rect 62426 23253 62438 23287
rect 61950 23247 62438 23253
rect 62968 23287 63456 23293
rect 62968 23253 62980 23287
rect 63444 23253 63456 23287
rect 62968 23247 63456 23253
rect 62160 23090 62220 23247
rect 62664 23132 62670 23192
rect 62730 23132 62736 23192
rect 62160 23084 62222 23090
rect 62160 23024 62162 23084
rect 62160 23018 62222 23024
rect 62160 22989 62220 23018
rect 61950 22983 62438 22989
rect 61950 22949 61962 22983
rect 62426 22949 62438 22983
rect 61950 22943 62438 22949
rect 60684 22314 60692 22344
rect 59914 22255 60402 22261
rect 59914 22221 59926 22255
rect 60390 22221 60402 22255
rect 59914 22215 60402 22221
rect 60120 22154 60180 22215
rect 60632 22160 60692 22314
rect 61654 22314 61668 22890
rect 61702 22314 61714 22890
rect 62670 22890 62730 23132
rect 63182 23090 63242 23247
rect 63180 23084 63242 23090
rect 63240 23024 63242 23084
rect 63180 23018 63242 23024
rect 63182 22989 63242 23018
rect 62968 22983 63456 22989
rect 62968 22949 62980 22983
rect 63444 22949 63456 22983
rect 62968 22943 63456 22949
rect 63182 22936 63242 22943
rect 62670 22844 62686 22890
rect 60932 22255 61420 22261
rect 60932 22221 60944 22255
rect 61408 22221 61420 22255
rect 60932 22215 61420 22221
rect 60626 22154 60632 22160
rect 59492 22100 60632 22154
rect 60692 22100 60698 22160
rect 59492 22094 60698 22100
rect 61138 22026 61198 22215
rect 61138 21960 61198 21966
rect 61654 21818 61714 22314
rect 62680 22314 62686 22844
rect 62720 22844 62730 22890
rect 63692 22890 63752 23346
rect 64712 23346 64722 23410
rect 64756 23410 64762 23922
rect 65730 23922 65790 24172
rect 66732 24068 66738 24128
rect 66798 24068 66804 24128
rect 66022 24015 66510 24021
rect 66022 23981 66034 24015
rect 66498 23981 66510 24015
rect 66022 23975 66510 23981
rect 64756 23346 64772 23410
rect 63986 23287 64474 23293
rect 63986 23253 63998 23287
rect 64462 23253 64474 23287
rect 63986 23247 64474 23253
rect 64202 23090 64262 23247
rect 64712 23192 64772 23346
rect 65730 23346 65740 23922
rect 65774 23346 65790 23922
rect 66738 23922 66798 24068
rect 67040 24015 67528 24021
rect 67040 23981 67052 24015
rect 67516 23981 67528 24015
rect 67040 23975 67528 23981
rect 66738 23848 66758 23922
rect 65218 23293 65278 23295
rect 65004 23287 65492 23293
rect 65004 23253 65016 23287
rect 65480 23253 65492 23287
rect 65004 23247 65492 23253
rect 64706 23132 64712 23192
rect 64772 23132 64778 23192
rect 64202 23084 64264 23090
rect 64202 23024 64204 23084
rect 64202 23018 64264 23024
rect 65218 23084 65278 23247
rect 64202 22989 64262 23018
rect 65218 22989 65278 23024
rect 63986 22983 64474 22989
rect 63986 22949 63998 22983
rect 64462 22949 64474 22983
rect 63986 22943 64474 22949
rect 65004 22983 65492 22989
rect 65004 22949 65016 22983
rect 65480 22949 65492 22983
rect 65004 22943 65492 22949
rect 62720 22314 62726 22844
rect 62680 22302 62726 22314
rect 63692 22314 63704 22890
rect 63738 22314 63752 22890
rect 64716 22890 64762 22902
rect 64716 22380 64722 22890
rect 62152 22261 62212 22264
rect 61950 22255 62438 22261
rect 61950 22221 61962 22255
rect 62426 22221 62438 22255
rect 61950 22215 62438 22221
rect 62968 22255 63456 22261
rect 62968 22221 62980 22255
rect 63444 22221 63456 22255
rect 62968 22215 63456 22221
rect 62152 22022 62212 22215
rect 63184 22030 63244 22215
rect 63184 21964 63244 21970
rect 62152 21956 62212 21962
rect 63692 21818 63752 22314
rect 64712 22314 64722 22380
rect 64756 22380 64762 22890
rect 65730 22890 65790 23346
rect 66752 23346 66758 23848
rect 66792 23346 66798 23922
rect 66752 23334 66798 23346
rect 67766 23922 67826 24172
rect 68058 24015 68546 24021
rect 68058 23981 68070 24015
rect 68534 23981 68546 24015
rect 68058 23975 68546 23981
rect 69076 24015 69564 24021
rect 69076 23981 69088 24015
rect 69552 23981 69564 24015
rect 69076 23975 69564 23981
rect 67766 23346 67776 23922
rect 67810 23346 67826 23922
rect 68788 23922 68834 23934
rect 68788 23410 68794 23922
rect 66022 23287 66510 23293
rect 66022 23253 66034 23287
rect 66498 23253 66510 23287
rect 66022 23247 66510 23253
rect 67040 23287 67528 23293
rect 67040 23253 67052 23287
rect 67516 23253 67528 23287
rect 67040 23247 67528 23253
rect 66234 23090 66294 23247
rect 66732 23132 66738 23192
rect 66798 23132 66804 23192
rect 66234 23084 66296 23090
rect 66234 23024 66236 23084
rect 66234 23018 66296 23024
rect 66234 22989 66294 23018
rect 66022 22983 66510 22989
rect 66022 22949 66034 22983
rect 66498 22949 66510 22983
rect 66022 22943 66510 22949
rect 64756 22314 64772 22380
rect 63986 22255 64474 22261
rect 63986 22221 63998 22255
rect 64462 22221 64474 22255
rect 63986 22215 64474 22221
rect 64182 22030 64242 22215
rect 64712 22160 64772 22314
rect 65730 22314 65740 22890
rect 65774 22314 65790 22890
rect 66738 22890 66798 23132
rect 67244 23090 67304 23247
rect 67244 23084 67306 23090
rect 67244 23024 67246 23084
rect 67244 23018 67306 23024
rect 67244 22989 67304 23018
rect 67040 22983 67528 22989
rect 67040 22949 67052 22983
rect 67516 22949 67528 22983
rect 67040 22943 67528 22949
rect 66738 22828 66758 22890
rect 66752 22406 66758 22828
rect 65226 22261 65286 22274
rect 65004 22255 65492 22261
rect 65004 22221 65016 22255
rect 65480 22221 65492 22255
rect 65004 22215 65492 22221
rect 64706 22100 64712 22160
rect 64772 22100 64778 22160
rect 64182 21964 64242 21970
rect 65226 22030 65286 22215
rect 65226 21964 65286 21970
rect 65730 21818 65790 22314
rect 66748 22314 66758 22406
rect 66792 22406 66798 22890
rect 67766 22890 67826 23346
rect 68780 23346 68794 23410
rect 68828 23410 68834 23922
rect 69796 23922 69856 24172
rect 70808 24068 70814 24128
rect 70874 24068 70880 24128
rect 70094 24015 70582 24021
rect 70094 23981 70106 24015
rect 70570 23981 70582 24015
rect 70094 23975 70582 23981
rect 69796 23512 69812 23922
rect 69806 23418 69812 23512
rect 68828 23346 68840 23410
rect 68266 23293 68326 23295
rect 68058 23287 68546 23293
rect 68058 23253 68070 23287
rect 68534 23253 68546 23287
rect 68058 23247 68546 23253
rect 68266 23090 68326 23247
rect 68780 23192 68840 23346
rect 69796 23346 69812 23418
rect 69846 23512 69856 23922
rect 70814 23922 70874 24068
rect 71112 24015 71600 24021
rect 71112 23981 71124 24015
rect 71588 23981 71600 24015
rect 71112 23975 71600 23981
rect 70814 23858 70830 23922
rect 69846 23418 69852 23512
rect 69846 23346 69856 23418
rect 69280 23293 69340 23295
rect 69076 23287 69564 23293
rect 69076 23253 69088 23287
rect 69552 23253 69564 23287
rect 69076 23247 69564 23253
rect 68774 23132 68780 23192
rect 68840 23132 68846 23192
rect 69280 23090 69340 23247
rect 68266 23084 68328 23090
rect 68266 23024 68268 23084
rect 68266 23018 68328 23024
rect 69280 23084 69342 23090
rect 69280 23024 69282 23084
rect 69280 23018 69342 23024
rect 68266 22989 68326 23018
rect 69280 22989 69340 23018
rect 68058 22983 68546 22989
rect 68058 22949 68070 22983
rect 68534 22949 68546 22983
rect 68058 22943 68546 22949
rect 69076 22983 69564 22989
rect 69076 22949 69088 22983
rect 69552 22949 69564 22983
rect 69076 22943 69564 22949
rect 66792 22314 66808 22406
rect 66230 22261 66290 22264
rect 66022 22255 66510 22261
rect 66022 22221 66034 22255
rect 66498 22221 66510 22255
rect 66022 22215 66510 22221
rect 66230 22026 66290 22215
rect 66230 21960 66290 21966
rect 66748 21910 66808 22314
rect 67766 22314 67776 22890
rect 67810 22314 67826 22890
rect 68788 22890 68834 22902
rect 68788 22396 68794 22890
rect 67246 22261 67306 22268
rect 67040 22255 67528 22261
rect 67040 22221 67052 22255
rect 67516 22221 67528 22255
rect 67040 22215 67528 22221
rect 67246 22026 67306 22215
rect 67246 21960 67306 21966
rect 66538 21850 66808 21910
rect 61654 21758 66030 21818
rect 66090 21758 66096 21818
rect 59378 21628 63546 21688
rect 59256 21440 59262 21500
rect 59322 21440 59328 21500
rect 60422 21440 60428 21500
rect 60488 21440 60494 21500
rect 58988 20394 58994 20454
rect 59054 20394 59060 20454
rect 58746 19236 58752 19296
rect 58812 19236 58818 19296
rect 58742 19022 58748 19082
rect 58808 19022 58814 19082
rect 58630 17980 58636 18040
rect 58696 17980 58702 18040
rect 53292 16726 58562 16786
rect 53232 16720 53292 16726
rect 11322 16122 35778 16128
rect 11322 16022 11428 16122
rect 35672 16022 35778 16122
rect 11322 16016 35778 16022
rect 37958 16188 49228 16248
rect 8084 15700 8228 15992
rect -3042 15392 8228 15700
rect 37958 15700 38024 16188
rect 38252 15992 49228 16188
rect 52322 16128 52434 16642
rect 54286 16524 54346 16530
rect 58748 16524 58808 19022
rect 58994 16782 59054 20394
rect 59124 20296 59130 20356
rect 59190 20296 59196 20356
rect 58988 16722 58994 16782
rect 59054 16722 59060 16782
rect 59130 16652 59190 20296
rect 59262 17832 59322 21440
rect 59706 21379 60194 21385
rect 59706 21345 59718 21379
rect 60182 21345 60194 21379
rect 59706 21339 60194 21345
rect 59418 21286 59464 21298
rect 59418 20746 59424 21286
rect 59410 20710 59424 20746
rect 59458 20746 59464 21286
rect 60428 21286 60488 21440
rect 60724 21379 61212 21385
rect 60724 21345 60736 21379
rect 61200 21345 61212 21379
rect 60724 21339 61212 21345
rect 60428 21260 60442 21286
rect 59458 20710 59470 20746
rect 60436 20734 60442 21260
rect 59410 20552 59470 20710
rect 60426 20710 60442 20734
rect 60476 21260 60488 21286
rect 61444 21286 61504 21628
rect 62458 21440 62464 21500
rect 62524 21440 62530 21500
rect 61742 21379 62230 21385
rect 61742 21345 61754 21379
rect 62218 21345 62230 21379
rect 61742 21339 62230 21345
rect 60476 20734 60482 21260
rect 61444 21240 61460 21286
rect 61454 20734 61460 21240
rect 60476 20710 60486 20734
rect 59706 20651 60194 20657
rect 59706 20617 59718 20651
rect 60182 20617 60194 20651
rect 59706 20611 60194 20617
rect 59924 20552 59984 20611
rect 60426 20552 60486 20710
rect 61446 20710 61460 20734
rect 61494 21240 61504 21286
rect 62464 21286 62524 21440
rect 62966 21436 62972 21500
rect 63036 21436 63042 21500
rect 62972 21385 63036 21436
rect 62760 21379 63248 21385
rect 62760 21345 62772 21379
rect 63236 21345 63248 21379
rect 62760 21339 63248 21345
rect 62464 21262 62478 21286
rect 61494 20734 61500 21240
rect 61494 20710 61506 20734
rect 60724 20651 61212 20657
rect 60724 20617 60736 20651
rect 61200 20617 61212 20651
rect 60724 20611 61212 20617
rect 59410 20492 60486 20552
rect 60916 20250 60976 20611
rect 61446 20552 61506 20710
rect 62472 20710 62478 21262
rect 62512 21262 62524 21286
rect 63486 21286 63546 21628
rect 63990 21385 64050 21758
rect 63778 21379 64266 21385
rect 63778 21345 63790 21379
rect 64254 21345 64266 21379
rect 63778 21339 64266 21345
rect 62512 20710 62518 21262
rect 63486 21232 63496 21286
rect 63490 20738 63496 21232
rect 62472 20698 62518 20710
rect 63482 20710 63496 20738
rect 63530 21232 63546 21286
rect 64498 21286 64558 21758
rect 64990 21385 65050 21758
rect 66028 21385 66088 21758
rect 64796 21379 65284 21385
rect 64796 21345 64808 21379
rect 65272 21345 65284 21379
rect 64796 21339 65284 21345
rect 65814 21379 66302 21385
rect 65814 21345 65826 21379
rect 66290 21345 66302 21379
rect 65814 21339 66302 21345
rect 63530 20738 63536 21232
rect 63530 20710 63542 20738
rect 61742 20651 62230 20657
rect 61742 20617 61754 20651
rect 62218 20617 62230 20651
rect 61742 20611 62230 20617
rect 62760 20651 63248 20657
rect 62760 20617 62772 20651
rect 63236 20617 63248 20651
rect 62760 20611 63248 20617
rect 61440 20492 61446 20552
rect 61506 20492 61512 20552
rect 61954 20498 62014 20611
rect 62960 20498 63020 20611
rect 63482 20552 63542 20710
rect 64498 20710 64514 21286
rect 64548 20710 64558 21286
rect 65526 21286 65572 21298
rect 65526 20734 65532 21286
rect 63778 20651 64266 20657
rect 63778 20617 63790 20651
rect 64254 20617 64266 20651
rect 63778 20611 64266 20617
rect 63992 20556 64052 20611
rect 64498 20556 64558 20710
rect 65518 20710 65532 20734
rect 65566 20734 65572 21286
rect 66538 21286 66598 21850
rect 67766 21818 67826 22314
rect 68780 22314 68794 22396
rect 68828 22396 68834 22890
rect 69796 22890 69856 23346
rect 70824 23346 70830 23858
rect 70864 23858 70874 23922
rect 71834 23922 71894 24172
rect 74004 24068 74010 24128
rect 74070 24068 74076 24128
rect 72130 24015 72618 24021
rect 72130 23981 72142 24015
rect 72606 23981 72618 24015
rect 72130 23975 72618 23981
rect 73148 24015 73636 24021
rect 73148 23981 73160 24015
rect 73624 23981 73636 24015
rect 73148 23975 73636 23981
rect 70864 23346 70870 23858
rect 70824 23334 70870 23346
rect 71834 23346 71848 23922
rect 71882 23346 71894 23922
rect 72860 23922 72906 23934
rect 72860 23422 72866 23922
rect 70312 23293 70372 23295
rect 71322 23293 71382 23295
rect 70094 23287 70582 23293
rect 70094 23253 70106 23287
rect 70570 23253 70582 23287
rect 70094 23247 70582 23253
rect 71112 23287 71600 23293
rect 71112 23253 71124 23287
rect 71588 23253 71600 23287
rect 71112 23247 71600 23253
rect 70312 23090 70372 23247
rect 70810 23132 70816 23192
rect 70876 23132 70882 23192
rect 70312 23084 70374 23090
rect 70312 23024 70314 23084
rect 70312 23018 70374 23024
rect 70312 22989 70372 23018
rect 70094 22983 70582 22989
rect 70094 22949 70106 22983
rect 70570 22949 70582 22983
rect 70094 22943 70582 22949
rect 68828 22314 68840 22396
rect 68058 22255 68546 22261
rect 68058 22221 68070 22255
rect 68534 22221 68546 22255
rect 68058 22215 68546 22221
rect 68250 22026 68310 22215
rect 68780 22160 68840 22314
rect 69796 22314 69812 22890
rect 69846 22314 69856 22890
rect 70816 22890 70876 23132
rect 71322 23090 71382 23247
rect 71322 23084 71384 23090
rect 71322 23024 71324 23084
rect 71322 23018 71384 23024
rect 71322 22989 71382 23018
rect 71112 22983 71600 22989
rect 71112 22949 71124 22983
rect 71588 22949 71600 22983
rect 71112 22943 71600 22949
rect 70816 22822 70830 22890
rect 69076 22255 69564 22261
rect 69076 22221 69088 22255
rect 69552 22221 69564 22255
rect 69076 22215 69564 22221
rect 68774 22100 68780 22160
rect 68840 22100 68846 22160
rect 68250 21960 68310 21966
rect 69282 22030 69342 22215
rect 69282 21964 69342 21970
rect 67040 21558 67046 21622
rect 67110 21558 67116 21622
rect 67046 21500 67110 21558
rect 67766 21528 67826 21758
rect 69796 21918 69856 22314
rect 70824 22314 70830 22822
rect 70864 22822 70876 22890
rect 71834 22890 71894 23346
rect 72852 23346 72866 23422
rect 72900 23422 72906 23922
rect 73878 23922 73924 23934
rect 72900 23346 72912 23422
rect 73878 23372 73884 23922
rect 72130 23287 72618 23293
rect 72130 23253 72142 23287
rect 72606 23253 72618 23287
rect 72130 23247 72618 23253
rect 72344 23090 72404 23247
rect 72852 23194 72912 23346
rect 73868 23346 73884 23372
rect 73918 23372 73924 23922
rect 73918 23346 73928 23372
rect 73148 23287 73636 23293
rect 73148 23253 73160 23287
rect 73624 23253 73636 23287
rect 73148 23247 73636 23253
rect 73374 23194 73434 23247
rect 73868 23194 73928 23346
rect 72852 23192 73928 23194
rect 72846 23132 72852 23192
rect 72912 23134 73928 23192
rect 72912 23132 72918 23134
rect 72344 23084 72406 23090
rect 72344 23024 72346 23084
rect 72344 23018 72406 23024
rect 72344 22989 72404 23018
rect 72130 22983 72618 22989
rect 72130 22949 72142 22983
rect 72606 22949 72618 22983
rect 72130 22943 72618 22949
rect 73148 22983 73636 22989
rect 73148 22949 73160 22983
rect 73624 22949 73636 22983
rect 73148 22943 73636 22949
rect 70864 22314 70870 22822
rect 70824 22302 70870 22314
rect 71834 22314 71848 22890
rect 71882 22314 71894 22890
rect 72860 22890 72906 22902
rect 72860 22390 72866 22890
rect 70298 22261 70358 22264
rect 70094 22255 70582 22261
rect 70094 22221 70106 22255
rect 70570 22221 70582 22255
rect 70094 22215 70582 22221
rect 71112 22255 71600 22261
rect 71112 22221 71124 22255
rect 71588 22221 71600 22255
rect 71112 22215 71600 22221
rect 70298 22026 70358 22215
rect 70298 21960 70358 21966
rect 71326 22026 71386 22215
rect 71326 21960 71386 21966
rect 71834 21918 71894 22314
rect 72848 22314 72866 22390
rect 72900 22390 72906 22890
rect 73878 22890 73924 22902
rect 72900 22314 72908 22390
rect 73878 22386 73884 22890
rect 72346 22261 72406 22264
rect 72130 22255 72618 22261
rect 72130 22221 72142 22255
rect 72606 22221 72618 22255
rect 72130 22215 72618 22221
rect 72346 22026 72406 22215
rect 72848 22164 72908 22314
rect 73868 22314 73884 22386
rect 73918 22386 73924 22890
rect 73918 22314 73928 22386
rect 73148 22255 73636 22261
rect 73148 22221 73160 22255
rect 73624 22221 73636 22255
rect 73148 22215 73636 22221
rect 73336 22164 73396 22215
rect 73868 22164 73928 22314
rect 74010 22164 74070 24068
rect 72846 22160 74070 22164
rect 72842 22100 72848 22160
rect 72908 22104 74070 22160
rect 72908 22100 72914 22104
rect 74798 21968 74804 22028
rect 74864 21968 74870 22028
rect 72346 21960 72406 21966
rect 69796 21858 71894 21918
rect 69796 21528 69856 21858
rect 73658 21742 73664 21802
rect 73724 21742 73730 21802
rect 71104 21558 71110 21622
rect 71174 21558 71180 21622
rect 72128 21558 72134 21622
rect 72198 21558 72204 21622
rect 73140 21558 73146 21622
rect 73210 21558 73216 21622
rect 67042 21436 67048 21500
rect 67112 21436 67118 21500
rect 67766 21468 70160 21528
rect 71110 21504 71174 21558
rect 67046 21385 67110 21436
rect 68078 21385 68138 21468
rect 66832 21379 67320 21385
rect 66832 21345 66844 21379
rect 67308 21345 67320 21379
rect 66832 21339 67320 21345
rect 67850 21379 68338 21385
rect 67850 21345 67862 21379
rect 68326 21345 68338 21379
rect 67850 21339 68338 21345
rect 65566 20710 65578 20734
rect 64796 20651 65284 20657
rect 64796 20617 64808 20651
rect 65272 20617 65284 20651
rect 64796 20611 65284 20617
rect 65012 20556 65072 20611
rect 65518 20556 65578 20710
rect 66538 20710 66550 21286
rect 66584 20710 66598 21286
rect 67562 21286 67608 21298
rect 67562 20788 67568 21286
rect 65814 20651 66302 20657
rect 65814 20617 65826 20651
rect 66290 20617 66302 20651
rect 65814 20611 66302 20617
rect 66022 20556 66082 20611
rect 61446 20356 61506 20492
rect 61954 20438 63020 20498
rect 63476 20492 63482 20552
rect 63542 20492 63548 20552
rect 63818 20494 63824 20554
rect 63884 20494 63890 20554
rect 63992 20496 66082 20556
rect 66538 20554 66598 20710
rect 67556 20710 67568 20788
rect 67602 20788 67608 21286
rect 68572 21286 68632 21468
rect 69100 21385 69160 21468
rect 68868 21379 69356 21385
rect 68868 21345 68880 21379
rect 69344 21345 69356 21379
rect 68868 21339 69356 21345
rect 69100 21338 69160 21339
rect 67602 20710 67616 20788
rect 66832 20651 67320 20657
rect 66832 20617 66844 20651
rect 67308 20617 67320 20651
rect 66832 20611 67320 20617
rect 61440 20296 61446 20356
rect 61506 20296 61512 20356
rect 61954 20250 62014 20438
rect 62460 20298 62466 20358
rect 62526 20298 62532 20358
rect 60426 20186 60432 20246
rect 60492 20186 60498 20246
rect 60916 20190 62014 20250
rect 62466 20246 62526 20298
rect 59706 20123 60194 20129
rect 59706 20089 59718 20123
rect 60182 20089 60194 20123
rect 59706 20083 60194 20089
rect 59418 20030 59464 20042
rect 59418 19490 59424 20030
rect 59414 19454 59424 19490
rect 59458 19490 59464 20030
rect 60432 20030 60492 20186
rect 60916 20129 60976 20190
rect 61954 20129 62014 20190
rect 62460 20186 62466 20246
rect 62526 20186 62532 20246
rect 60724 20123 61212 20129
rect 60724 20089 60736 20123
rect 61200 20089 61212 20123
rect 60724 20083 61212 20089
rect 61742 20123 62230 20129
rect 61742 20089 61754 20123
rect 62218 20089 62230 20123
rect 61742 20083 62230 20089
rect 60432 20004 60442 20030
rect 59458 19454 59474 19490
rect 60436 19478 60442 20004
rect 59414 19296 59474 19454
rect 60430 19454 60442 19478
rect 60476 20004 60492 20030
rect 61454 20030 61500 20042
rect 60476 19478 60482 20004
rect 61454 19480 61460 20030
rect 60476 19454 60490 19478
rect 59706 19395 60194 19401
rect 59706 19361 59718 19395
rect 60182 19361 60194 19395
rect 59706 19355 60194 19361
rect 59928 19296 59988 19355
rect 60430 19296 60490 19454
rect 61448 19454 61460 19480
rect 61494 19480 61500 20030
rect 62466 20030 62526 20186
rect 62960 20129 63020 20438
rect 63824 20240 63884 20494
rect 63482 20180 63884 20240
rect 62760 20123 63248 20129
rect 62760 20089 62772 20123
rect 63236 20089 63248 20123
rect 62760 20083 63248 20089
rect 62466 20008 62478 20030
rect 61494 19454 61508 19480
rect 60910 19401 60970 19402
rect 60724 19395 61212 19401
rect 60724 19361 60736 19395
rect 61200 19361 61212 19395
rect 60724 19355 61212 19361
rect 59414 19236 60490 19296
rect 59414 19082 59474 19236
rect 59408 19022 59414 19082
rect 59474 19022 59480 19082
rect 59412 18912 60488 18972
rect 59412 18774 59472 18912
rect 59926 18873 59986 18912
rect 59706 18867 60194 18873
rect 59706 18833 59718 18867
rect 60182 18833 60194 18867
rect 59706 18827 60194 18833
rect 59412 18740 59424 18774
rect 59418 18198 59424 18740
rect 59458 18740 59472 18774
rect 60428 18774 60488 18912
rect 60910 18873 60970 19355
rect 61448 19192 61508 19454
rect 62472 19454 62478 20008
rect 62512 20008 62526 20030
rect 63482 20030 63542 20180
rect 63778 20123 64266 20129
rect 63778 20089 63790 20123
rect 64254 20089 64266 20123
rect 63778 20083 64266 20089
rect 62512 19454 62518 20008
rect 63482 19972 63496 20030
rect 63490 19484 63496 19972
rect 62472 19442 62518 19454
rect 63484 19454 63496 19484
rect 63530 19972 63542 20030
rect 64498 20030 64558 20496
rect 66532 20494 66538 20554
rect 66598 20494 66604 20554
rect 67556 20358 67616 20710
rect 68572 20710 68586 21286
rect 68620 20710 68632 21286
rect 67850 20651 68338 20657
rect 67850 20617 67862 20651
rect 68326 20617 68338 20651
rect 67850 20611 68338 20617
rect 68066 20556 68126 20611
rect 68572 20556 68632 20710
rect 69588 21286 69648 21468
rect 70100 21385 70160 21468
rect 70604 21440 70610 21500
rect 70670 21440 70676 21500
rect 69886 21379 70374 21385
rect 69886 21345 69898 21379
rect 70362 21345 70374 21379
rect 69886 21339 70374 21345
rect 70100 21332 70160 21339
rect 69588 20710 69604 21286
rect 69638 20710 69648 21286
rect 70610 21286 70670 21440
rect 71110 21385 71174 21440
rect 72134 21385 72198 21558
rect 72638 21440 72644 21500
rect 72704 21440 72710 21500
rect 70904 21379 71392 21385
rect 70904 21345 70916 21379
rect 71380 21345 71392 21379
rect 70904 21339 71392 21345
rect 71922 21379 72410 21385
rect 71922 21345 71934 21379
rect 72398 21345 72410 21379
rect 71922 21339 72410 21345
rect 70610 21258 70622 21286
rect 68868 20651 69356 20657
rect 68868 20617 68880 20651
rect 69344 20617 69356 20651
rect 68868 20611 69356 20617
rect 69092 20556 69152 20611
rect 69588 20556 69648 20710
rect 70616 20710 70622 21258
rect 70656 21258 70670 21286
rect 71634 21286 71680 21298
rect 70656 20710 70662 21258
rect 71634 20734 71640 21286
rect 70616 20698 70662 20710
rect 71626 20710 71640 20734
rect 71674 20734 71680 21286
rect 72644 21286 72704 21440
rect 73146 21385 73210 21558
rect 73664 21504 73724 21742
rect 73664 21444 74740 21504
rect 72940 21379 73428 21385
rect 72940 21345 72952 21379
rect 73416 21345 73428 21379
rect 72940 21339 73428 21345
rect 72644 21262 72658 21286
rect 71674 20710 71686 20734
rect 69886 20651 70374 20657
rect 69886 20617 69898 20651
rect 70362 20617 70374 20651
rect 69886 20611 70374 20617
rect 70904 20651 71392 20657
rect 70904 20617 70916 20651
rect 71380 20617 71392 20651
rect 70904 20611 71392 20617
rect 70104 20556 70164 20611
rect 68066 20496 70164 20556
rect 67550 20298 67556 20358
rect 67616 20298 67622 20358
rect 65516 20184 65522 20244
rect 65582 20184 65588 20244
rect 67550 20184 67556 20244
rect 67616 20184 67622 20244
rect 64796 20123 65284 20129
rect 64796 20089 64808 20123
rect 65272 20089 65284 20123
rect 64796 20083 65284 20089
rect 64498 19986 64514 20030
rect 63530 19484 63536 19972
rect 64508 19484 64514 19986
rect 63530 19454 63544 19484
rect 61948 19401 62008 19402
rect 62954 19401 63014 19402
rect 61742 19395 62230 19401
rect 61742 19361 61754 19395
rect 62218 19361 62230 19395
rect 61742 19355 62230 19361
rect 62760 19395 63248 19401
rect 62760 19361 62772 19395
rect 63236 19361 63248 19395
rect 62760 19355 63248 19361
rect 61448 19126 61508 19132
rect 61442 18928 61448 18988
rect 61508 18928 61514 18988
rect 60724 18867 61212 18873
rect 60724 18833 60736 18867
rect 61200 18833 61212 18867
rect 60724 18827 61212 18833
rect 60428 18752 60442 18774
rect 59458 18198 59464 18740
rect 60436 18226 60442 18752
rect 59418 18186 59464 18198
rect 60430 18198 60442 18226
rect 60476 18752 60488 18774
rect 61448 18774 61508 18928
rect 61948 18873 62008 19355
rect 62954 18873 63014 19355
rect 63484 19192 63544 19454
rect 64500 19454 64514 19484
rect 64548 19986 64558 20030
rect 65522 20030 65582 20184
rect 65814 20123 66302 20129
rect 65814 20089 65826 20123
rect 66290 20089 66302 20123
rect 65814 20083 66302 20089
rect 66832 20123 67320 20129
rect 66832 20089 66844 20123
rect 67308 20089 67320 20123
rect 66832 20083 67320 20089
rect 65522 20002 65532 20030
rect 64548 19484 64554 19986
rect 64548 19454 64560 19484
rect 63778 19395 64266 19401
rect 63778 19361 63790 19395
rect 64254 19361 64266 19395
rect 63778 19355 64266 19361
rect 64004 19300 64064 19355
rect 64500 19300 64560 19454
rect 65526 19454 65532 20002
rect 65566 20002 65582 20030
rect 66544 20030 66590 20042
rect 65566 19454 65572 20002
rect 66544 19478 66550 20030
rect 65526 19442 65572 19454
rect 66538 19454 66550 19478
rect 66584 19478 66590 20030
rect 67556 20030 67616 20184
rect 67850 20123 68338 20129
rect 67850 20089 67862 20123
rect 68326 20089 68338 20123
rect 67850 20083 68338 20089
rect 68868 20123 69356 20129
rect 68868 20089 68880 20123
rect 69344 20089 69356 20123
rect 68868 20083 69356 20089
rect 67556 20000 67568 20030
rect 67562 19482 67568 20000
rect 66584 19454 66598 19478
rect 64796 19395 65284 19401
rect 64796 19361 64808 19395
rect 65272 19361 65284 19395
rect 64796 19355 65284 19361
rect 65814 19395 66302 19401
rect 65814 19361 65826 19395
rect 66290 19361 66302 19395
rect 65814 19355 66302 19361
rect 65016 19300 65076 19355
rect 64004 19240 65076 19300
rect 63478 19132 63484 19192
rect 63544 19132 63550 19192
rect 63476 19030 63482 19090
rect 63542 19030 63548 19090
rect 63482 18988 63542 19030
rect 63476 18928 63482 18988
rect 63542 18928 63548 18988
rect 61742 18867 62230 18873
rect 61742 18833 61754 18867
rect 62218 18833 62230 18867
rect 61742 18827 62230 18833
rect 62760 18867 63248 18873
rect 62760 18833 62772 18867
rect 63236 18833 63248 18867
rect 62760 18827 63248 18833
rect 60476 18226 60482 18752
rect 61448 18750 61460 18774
rect 60476 18198 60490 18226
rect 59706 18139 60194 18145
rect 59706 18105 59718 18139
rect 60182 18105 60194 18139
rect 59706 18099 60194 18105
rect 60430 18040 60490 18198
rect 61454 18198 61460 18750
rect 61494 18750 61508 18774
rect 62472 18774 62518 18786
rect 61494 18198 61500 18750
rect 62472 18222 62478 18774
rect 61454 18186 61500 18198
rect 62466 18198 62478 18222
rect 62512 18222 62518 18774
rect 63482 18774 63542 18928
rect 63778 18867 64266 18873
rect 63778 18833 63790 18867
rect 64254 18833 64266 18867
rect 63778 18827 64266 18833
rect 63482 18746 63496 18774
rect 62512 18198 62526 18222
rect 63490 18217 63496 18746
rect 60922 18145 60982 18152
rect 61960 18145 62020 18152
rect 60724 18139 61212 18145
rect 60724 18105 60736 18139
rect 61200 18105 61212 18139
rect 60724 18099 61212 18105
rect 61742 18139 62230 18145
rect 61742 18105 61754 18139
rect 62218 18105 62230 18139
rect 61742 18099 62230 18105
rect 60424 17980 60430 18040
rect 60490 17980 60496 18040
rect 59256 17772 59262 17832
rect 59322 17772 59328 17832
rect 59412 17674 60488 17734
rect 59412 17518 59472 17674
rect 59926 17617 59986 17674
rect 59706 17611 60194 17617
rect 59706 17577 59718 17611
rect 60182 17577 60194 17611
rect 59706 17571 60194 17577
rect 59412 17480 59424 17518
rect 59418 16942 59424 17480
rect 59458 17480 59472 17518
rect 60428 17518 60488 17674
rect 60922 17617 60982 18099
rect 61438 17670 61444 17730
rect 61504 17670 61510 17730
rect 60724 17611 61212 17617
rect 60724 17577 60736 17611
rect 61200 17577 61212 17611
rect 60724 17571 61212 17577
rect 60428 17492 60442 17518
rect 59458 16942 59464 17480
rect 60436 16968 60442 17492
rect 59418 16930 59464 16942
rect 60426 16942 60442 16968
rect 60476 17492 60488 17518
rect 61444 17518 61504 17670
rect 61960 17617 62020 18099
rect 62466 18040 62526 18198
rect 63484 18198 63496 18217
rect 63530 18746 63542 18774
rect 64500 18774 64560 19240
rect 65512 19236 65518 19296
rect 65578 19236 65584 19296
rect 64796 18867 65284 18873
rect 64796 18833 64808 18867
rect 65272 18833 65284 18867
rect 64796 18827 65284 18833
rect 63530 18217 63536 18746
rect 64500 18736 64514 18774
rect 64508 18232 64514 18736
rect 63530 18198 63544 18217
rect 62966 18145 63026 18152
rect 62760 18139 63248 18145
rect 62760 18105 62772 18139
rect 63236 18105 63248 18139
rect 62760 18099 63248 18105
rect 62460 17980 62466 18040
rect 62526 17980 62532 18040
rect 62466 17932 62526 17980
rect 62460 17872 62466 17932
rect 62526 17872 62532 17932
rect 62966 17882 63026 18099
rect 63484 18048 63544 18198
rect 64498 18198 64514 18232
rect 64548 18736 64560 18774
rect 65518 18774 65578 19236
rect 66020 19134 66080 19355
rect 66538 19296 66598 19454
rect 67556 19454 67568 19482
rect 67602 20000 67616 20030
rect 68580 20030 68626 20042
rect 67602 19482 67608 20000
rect 68580 19482 68586 20030
rect 67602 19454 67616 19482
rect 67050 19401 67110 19408
rect 66832 19395 67320 19401
rect 66832 19361 66844 19395
rect 67308 19361 67320 19395
rect 66832 19355 67320 19361
rect 66532 19236 66538 19296
rect 66598 19236 66604 19296
rect 67050 19134 67110 19355
rect 66020 19074 67110 19134
rect 66020 18873 66080 19074
rect 66532 18930 66538 18990
rect 66598 18930 66604 18990
rect 65814 18867 66302 18873
rect 65814 18833 65826 18867
rect 66290 18833 66302 18867
rect 65814 18827 66302 18833
rect 66020 18822 66080 18827
rect 65518 18750 65532 18774
rect 64548 18232 64554 18736
rect 64548 18198 64558 18232
rect 65526 18228 65532 18750
rect 63778 18139 64266 18145
rect 63778 18105 63790 18139
rect 64254 18105 64266 18139
rect 63778 18099 64266 18105
rect 64002 18048 64062 18099
rect 64498 18048 64558 18198
rect 65520 18198 65532 18228
rect 65566 18750 65578 18774
rect 66538 18774 66598 18930
rect 67050 18873 67110 19074
rect 67556 18990 67616 19454
rect 68574 19454 68586 19482
rect 68620 19482 68626 20030
rect 69588 20030 69648 20496
rect 70606 20184 70612 20244
rect 70672 20184 70678 20244
rect 69886 20123 70374 20129
rect 69886 20089 69898 20123
rect 70362 20089 70374 20123
rect 69886 20083 70374 20089
rect 69588 20010 69604 20030
rect 69598 19482 69604 20010
rect 68620 19454 68634 19482
rect 68062 19401 68122 19408
rect 67850 19395 68338 19401
rect 67850 19361 67862 19395
rect 68326 19361 68338 19395
rect 67850 19355 68338 19361
rect 67550 18930 67556 18990
rect 67616 18930 67622 18990
rect 68062 18873 68122 19355
rect 68574 19296 68634 19454
rect 69588 19454 69604 19482
rect 69638 20010 69648 20030
rect 70612 20030 70672 20184
rect 71112 20129 71172 20611
rect 71626 20552 71686 20710
rect 72652 20710 72658 21262
rect 72692 21262 72704 21286
rect 73664 21286 73724 21444
rect 74178 21385 74238 21444
rect 73958 21379 74446 21385
rect 73958 21345 73970 21379
rect 74434 21345 74446 21379
rect 73958 21339 74446 21345
rect 72692 20710 72698 21262
rect 73664 21250 73676 21286
rect 73670 20738 73676 21250
rect 72652 20698 72698 20710
rect 73662 20710 73676 20738
rect 73710 21250 73724 21286
rect 74680 21286 74740 21444
rect 74680 21262 74694 21286
rect 73710 20738 73716 21250
rect 73710 20710 73722 20738
rect 73142 20657 73202 20663
rect 71922 20651 72410 20657
rect 71922 20617 71934 20651
rect 72398 20617 72410 20651
rect 71922 20611 72410 20617
rect 72940 20651 73428 20657
rect 72940 20617 72952 20651
rect 73416 20617 73428 20651
rect 72940 20611 73428 20617
rect 71620 20492 71626 20552
rect 71686 20492 71692 20552
rect 72136 20129 72196 20611
rect 72640 20184 72646 20244
rect 72706 20184 72712 20244
rect 70904 20123 71392 20129
rect 70904 20089 70916 20123
rect 71380 20089 71392 20123
rect 70904 20083 71392 20089
rect 71922 20123 72410 20129
rect 71922 20089 71934 20123
rect 72398 20089 72410 20123
rect 71922 20083 72410 20089
rect 69638 19482 69644 20010
rect 70612 20002 70622 20030
rect 69638 19454 69648 19482
rect 68868 19395 69356 19401
rect 68868 19361 68880 19395
rect 69344 19361 69356 19395
rect 68868 19355 69356 19361
rect 69092 19298 69152 19355
rect 69588 19298 69648 19454
rect 70616 19454 70622 20002
rect 70656 20002 70672 20030
rect 71634 20030 71680 20042
rect 70656 19454 70662 20002
rect 71634 19490 71640 20030
rect 70616 19442 70662 19454
rect 71624 19454 71640 19490
rect 71674 19490 71680 20030
rect 72646 20030 72706 20184
rect 73142 20129 73202 20611
rect 73662 20552 73722 20710
rect 74688 20710 74694 21262
rect 74728 21262 74740 21286
rect 74728 20710 74734 21262
rect 74688 20698 74734 20710
rect 73958 20651 74446 20657
rect 73958 20617 73970 20651
rect 74434 20617 74446 20651
rect 73958 20611 74446 20617
rect 73656 20492 73662 20552
rect 73722 20492 73728 20552
rect 73664 20190 74740 20250
rect 72940 20123 73428 20129
rect 72940 20089 72952 20123
rect 73416 20089 73428 20123
rect 72940 20083 73428 20089
rect 72646 20006 72658 20030
rect 71674 19454 71684 19490
rect 72652 19482 72658 20006
rect 71106 19401 71166 19402
rect 69886 19395 70374 19401
rect 69886 19361 69898 19395
rect 70362 19361 70374 19395
rect 69886 19355 70374 19361
rect 70904 19395 71392 19401
rect 70904 19361 70916 19395
rect 71380 19361 71392 19395
rect 70904 19355 71392 19361
rect 70104 19298 70164 19355
rect 68568 19236 68574 19296
rect 68634 19236 68640 19296
rect 69092 19238 70164 19298
rect 68566 18930 68572 18990
rect 68632 18930 68638 18990
rect 66832 18867 67320 18873
rect 66832 18833 66844 18867
rect 67308 18833 67320 18867
rect 66832 18827 67320 18833
rect 67850 18867 68338 18873
rect 67850 18833 67862 18867
rect 68326 18833 68338 18867
rect 67850 18827 68338 18833
rect 66538 18752 66550 18774
rect 65566 18228 65572 18750
rect 65566 18198 65580 18228
rect 64796 18139 65284 18145
rect 64796 18105 64808 18139
rect 65272 18105 65284 18139
rect 64796 18099 65284 18105
rect 65014 18048 65074 18099
rect 63478 17988 63484 18048
rect 63544 17988 63550 18048
rect 64002 17988 65074 18048
rect 65280 17988 65286 18048
rect 65346 17988 65352 18048
rect 65520 18042 65580 18198
rect 66544 18198 66550 18752
rect 66584 18752 66598 18774
rect 67562 18774 67608 18786
rect 66584 18198 66590 18752
rect 67562 18224 67568 18774
rect 66544 18186 66590 18198
rect 67556 18198 67568 18224
rect 67602 18224 67608 18774
rect 68572 18774 68632 18930
rect 68868 18867 69356 18873
rect 68868 18833 68880 18867
rect 69344 18833 69356 18867
rect 68868 18827 69356 18833
rect 68572 18748 68586 18774
rect 67602 18198 67616 18224
rect 65814 18139 66302 18145
rect 65814 18105 65826 18139
rect 66290 18105 66302 18139
rect 65814 18099 66302 18105
rect 66832 18139 67320 18145
rect 66832 18105 66844 18139
rect 67308 18105 67320 18139
rect 66832 18099 67320 18105
rect 62966 17822 63742 17882
rect 62966 17617 63026 17822
rect 63472 17670 63478 17730
rect 63538 17670 63544 17730
rect 63682 17718 63742 17822
rect 61742 17611 62230 17617
rect 61742 17577 61754 17611
rect 62218 17577 62230 17611
rect 61742 17571 62230 17577
rect 62760 17611 63248 17617
rect 62760 17577 62772 17611
rect 63236 17577 63248 17611
rect 62760 17571 63248 17577
rect 61444 17492 61460 17518
rect 60476 16968 60482 17492
rect 60476 16942 60486 16968
rect 59706 16883 60194 16889
rect 59706 16849 59718 16883
rect 60182 16849 60194 16883
rect 59706 16843 60194 16849
rect 60426 16782 60486 16942
rect 61454 16942 61460 17492
rect 61494 17492 61504 17518
rect 62472 17518 62518 17530
rect 61494 16942 61500 17492
rect 62472 16964 62478 17518
rect 61454 16930 61500 16942
rect 62462 16942 62478 16964
rect 62512 16964 62518 17518
rect 63478 17518 63538 17670
rect 63676 17658 63682 17718
rect 63742 17658 63748 17718
rect 63778 17611 64266 17617
rect 63778 17577 63790 17611
rect 64254 17577 64266 17611
rect 63778 17571 64266 17577
rect 63478 17488 63496 17518
rect 63490 16978 63496 17488
rect 62512 16942 62522 16964
rect 60724 16883 61212 16889
rect 60724 16849 60736 16883
rect 61200 16849 61212 16883
rect 60724 16843 61212 16849
rect 61742 16883 62230 16889
rect 61742 16849 61754 16883
rect 62218 16849 62230 16883
rect 61742 16843 62230 16849
rect 60420 16722 60426 16782
rect 60486 16722 60492 16782
rect 60934 16668 60994 16843
rect 61958 16668 62018 16843
rect 62462 16782 62522 16942
rect 63484 16942 63496 16978
rect 63530 17488 63538 17518
rect 64498 17518 64558 17988
rect 65286 17778 65346 17988
rect 65514 17982 65520 18042
rect 65580 17982 65586 18042
rect 66016 17920 66076 18099
rect 67044 17920 67104 18099
rect 67556 18042 67616 18198
rect 68580 18198 68586 18748
rect 68620 18748 68632 18774
rect 69588 18774 69648 19238
rect 70602 19132 70608 19192
rect 70668 19132 70674 19192
rect 69886 18867 70374 18873
rect 69886 18833 69898 18867
rect 70362 18833 70374 18867
rect 69886 18827 70374 18833
rect 68620 18198 68626 18748
rect 69588 18744 69604 18774
rect 69598 18230 69604 18744
rect 68580 18186 68626 18198
rect 69586 18198 69604 18230
rect 69638 18744 69648 18774
rect 70608 18774 70668 19132
rect 71106 18873 71166 19355
rect 71470 19250 71476 19310
rect 71536 19250 71542 19310
rect 71476 18990 71536 19250
rect 71624 19200 71684 19454
rect 72644 19454 72658 19482
rect 72692 20006 72706 20030
rect 73664 20030 73724 20190
rect 74178 20129 74238 20190
rect 73958 20123 74446 20129
rect 73958 20089 73970 20123
rect 74434 20089 74446 20123
rect 73958 20083 74446 20089
rect 72692 19482 72698 20006
rect 73664 19996 73676 20030
rect 73670 19494 73676 19996
rect 72692 19454 72704 19482
rect 72130 19401 72190 19402
rect 71922 19395 72410 19401
rect 71922 19361 71934 19395
rect 72398 19361 72410 19395
rect 71922 19355 72410 19361
rect 71618 19140 71624 19200
rect 71684 19140 71690 19200
rect 71470 18930 71476 18990
rect 71536 18930 71542 18990
rect 71622 18932 71628 18992
rect 71688 18932 71694 18992
rect 70904 18867 71392 18873
rect 70904 18833 70916 18867
rect 71380 18833 71392 18867
rect 70904 18827 71392 18833
rect 69638 18230 69644 18744
rect 70608 18742 70622 18774
rect 70616 18230 70622 18742
rect 69638 18198 69646 18230
rect 67850 18139 68338 18145
rect 67850 18105 67862 18139
rect 68326 18105 68338 18139
rect 67850 18099 68338 18105
rect 68868 18139 69356 18145
rect 68868 18105 68880 18139
rect 69344 18105 69356 18139
rect 68868 18099 69356 18105
rect 67550 17982 67556 18042
rect 67616 17982 67622 18042
rect 66016 17860 67104 17920
rect 67548 17872 67554 17932
rect 67614 17872 67620 17932
rect 65286 17718 66594 17778
rect 64796 17611 65284 17617
rect 64796 17577 64808 17611
rect 65272 17577 65284 17611
rect 64796 17571 65284 17577
rect 65814 17611 66302 17617
rect 65814 17577 65826 17611
rect 66290 17577 66302 17611
rect 65814 17571 66302 17577
rect 63530 16978 63536 17488
rect 64498 17460 64514 17518
rect 63530 16942 63544 16978
rect 64508 16974 64514 17460
rect 62760 16883 63248 16889
rect 62760 16849 62772 16883
rect 63236 16849 63248 16883
rect 62760 16843 63248 16849
rect 62456 16722 62462 16782
rect 62522 16722 62528 16782
rect 62964 16668 63024 16843
rect 59124 16592 59130 16652
rect 59190 16592 59196 16652
rect 60934 16608 63024 16668
rect 54282 16464 54286 16524
rect 54346 16464 58808 16524
rect 54286 16458 54346 16464
rect 54166 16406 54226 16412
rect 59130 16406 59190 16592
rect 54226 16346 59190 16406
rect 54166 16340 54226 16346
rect 53720 16288 53780 16294
rect 60934 16288 60994 16608
rect 62964 16398 63024 16608
rect 63484 16512 63544 16942
rect 64498 16942 64514 16974
rect 64548 17460 64558 17518
rect 65526 17518 65572 17530
rect 64548 16974 64554 17460
rect 65526 16986 65532 17518
rect 64548 16942 64558 16974
rect 63778 16883 64266 16889
rect 63778 16849 63790 16883
rect 64254 16849 64266 16883
rect 63778 16843 64266 16849
rect 64002 16788 64062 16843
rect 64498 16788 64558 16942
rect 65520 16942 65532 16986
rect 65566 16986 65572 17518
rect 66534 17518 66594 17718
rect 67044 17718 67104 17860
rect 67044 17617 67104 17658
rect 66832 17611 67320 17617
rect 66832 17577 66844 17611
rect 67308 17577 67320 17611
rect 66832 17571 67320 17577
rect 66534 17466 66550 17518
rect 65566 16942 65580 16986
rect 64796 16883 65284 16889
rect 64796 16849 64808 16883
rect 65272 16849 65284 16883
rect 64796 16843 65284 16849
rect 65014 16788 65074 16843
rect 65520 16788 65580 16942
rect 66544 16942 66550 17466
rect 66584 17466 66594 17518
rect 67554 17518 67614 17872
rect 68060 17718 68120 18099
rect 69090 18046 69150 18099
rect 69586 18046 69646 18198
rect 70610 18198 70622 18230
rect 70656 18742 70668 18774
rect 71628 18774 71688 18932
rect 72130 18873 72190 19355
rect 72644 19090 72704 19454
rect 73664 19454 73676 19494
rect 73710 19996 73724 20030
rect 74680 20030 74740 20190
rect 74680 20008 74694 20030
rect 73710 19494 73716 19996
rect 73710 19454 73724 19494
rect 73136 19401 73196 19408
rect 72940 19395 73428 19401
rect 72940 19361 72952 19395
rect 73416 19361 73428 19395
rect 72940 19355 73428 19361
rect 72638 19030 72644 19090
rect 72704 19030 72710 19090
rect 73136 18873 73196 19355
rect 73664 19200 73724 19454
rect 74688 19454 74694 20008
rect 74728 20008 74740 20030
rect 74728 19454 74734 20008
rect 74688 19442 74734 19454
rect 73958 19395 74446 19401
rect 73958 19361 73970 19395
rect 74434 19361 74446 19395
rect 73958 19355 74446 19361
rect 74804 19200 74864 21968
rect 74946 21800 75006 24516
rect 75234 22100 75240 22160
rect 75300 22100 75306 22160
rect 74946 21734 75006 21740
rect 75082 21440 75088 21500
rect 75148 21440 75154 21500
rect 74922 20298 74928 20358
rect 74988 20298 74994 20358
rect 73658 19140 73664 19200
rect 73724 19140 73730 19200
rect 74798 19140 74804 19200
rect 74864 19140 74870 19200
rect 73656 18932 73662 18992
rect 73722 18932 73728 18992
rect 71922 18867 72410 18873
rect 71922 18833 71934 18867
rect 72398 18833 72410 18867
rect 71922 18827 72410 18833
rect 72940 18867 73428 18873
rect 72940 18833 72952 18867
rect 73416 18833 73428 18867
rect 72940 18827 73428 18833
rect 71628 18754 71640 18774
rect 70656 18230 70662 18742
rect 70656 18198 70670 18230
rect 69886 18139 70374 18145
rect 69886 18105 69898 18139
rect 70362 18105 70374 18139
rect 69886 18099 70374 18105
rect 70102 18046 70162 18099
rect 69090 17986 70162 18046
rect 70610 18044 70670 18198
rect 71634 18198 71640 18754
rect 71674 18754 71688 18774
rect 72652 18774 72698 18786
rect 71674 18198 71680 18754
rect 72652 18226 72658 18774
rect 71634 18186 71680 18198
rect 72646 18198 72658 18226
rect 72692 18226 72698 18774
rect 73662 18774 73722 18932
rect 73958 18867 74446 18873
rect 73958 18833 73970 18867
rect 74434 18833 74446 18867
rect 73958 18827 74446 18833
rect 73662 18750 73676 18774
rect 73670 18234 73676 18750
rect 72692 18198 72706 18226
rect 71118 18145 71178 18152
rect 72142 18145 72202 18152
rect 70904 18139 71392 18145
rect 70904 18105 70916 18139
rect 71380 18105 71392 18139
rect 70904 18099 71392 18105
rect 71922 18139 72410 18145
rect 71922 18105 71934 18139
rect 72398 18105 72410 18139
rect 71922 18099 72410 18105
rect 68060 17652 68120 17658
rect 67850 17611 68338 17617
rect 67850 17577 67862 17611
rect 68326 17577 68338 17611
rect 67850 17571 68338 17577
rect 68868 17611 69356 17617
rect 68868 17577 68880 17611
rect 69344 17577 69356 17611
rect 68868 17571 69356 17577
rect 66584 16942 66590 17466
rect 67554 17454 67568 17518
rect 66544 16930 66590 16942
rect 67562 16942 67568 17454
rect 67602 17454 67614 17518
rect 68580 17518 68626 17530
rect 67602 16942 67608 17454
rect 68580 16970 68586 17518
rect 67562 16930 67608 16942
rect 68572 16942 68586 16970
rect 68620 16970 68626 17518
rect 69586 17518 69646 17986
rect 70604 17984 70610 18044
rect 70670 17984 70676 18044
rect 71118 17724 71178 18099
rect 71118 17718 71180 17724
rect 71118 17658 71120 17718
rect 71626 17670 71632 17730
rect 71692 17670 71698 17730
rect 71118 17652 71180 17658
rect 71118 17617 71178 17652
rect 69886 17611 70374 17617
rect 69886 17577 69898 17611
rect 70362 17577 70374 17611
rect 69886 17571 70374 17577
rect 70904 17611 71392 17617
rect 70904 17577 70916 17611
rect 71380 17577 71392 17611
rect 70904 17571 71392 17577
rect 69586 17480 69604 17518
rect 69598 16972 69604 17480
rect 68620 16942 68632 16970
rect 65814 16883 66302 16889
rect 65814 16849 65826 16883
rect 66290 16849 66302 16883
rect 65814 16843 66302 16849
rect 66832 16883 67320 16889
rect 66832 16849 66844 16883
rect 67308 16849 67320 16883
rect 66832 16843 67320 16849
rect 67850 16883 68338 16889
rect 67850 16849 67862 16883
rect 68326 16849 68338 16883
rect 67850 16843 68338 16849
rect 66030 16788 66090 16843
rect 68056 16788 68116 16843
rect 68572 16788 68632 16942
rect 69586 16942 69604 16972
rect 69638 17480 69646 17518
rect 70616 17518 70662 17530
rect 69638 16972 69644 17480
rect 69638 16942 69646 16972
rect 70616 16968 70622 17518
rect 68868 16883 69356 16889
rect 68868 16849 68880 16883
rect 69344 16849 69356 16883
rect 68868 16843 69356 16849
rect 69090 16788 69150 16843
rect 69586 16788 69646 16942
rect 70614 16942 70622 16968
rect 70656 16968 70662 17518
rect 71632 17518 71692 17670
rect 72142 17617 72202 18099
rect 72646 18044 72706 18198
rect 73662 18198 73676 18234
rect 73710 18750 73722 18774
rect 74688 18774 74734 18786
rect 73710 18234 73716 18750
rect 73710 18198 73722 18234
rect 74688 18222 74694 18774
rect 73148 18145 73208 18158
rect 72940 18139 73428 18145
rect 72940 18105 72952 18139
rect 73416 18105 73428 18139
rect 72940 18099 73428 18105
rect 72640 17984 72646 18044
rect 72706 17984 72712 18044
rect 73148 17617 73208 18099
rect 73662 18040 73722 18198
rect 74678 18198 74694 18222
rect 74728 18222 74734 18774
rect 74728 18198 74738 18222
rect 73958 18139 74446 18145
rect 73958 18105 73970 18139
rect 74434 18105 74446 18139
rect 73958 18099 74446 18105
rect 74176 18040 74236 18099
rect 74678 18040 74738 18198
rect 73662 17980 74738 18040
rect 74804 17932 74864 19140
rect 74928 18992 74988 20298
rect 74922 18932 74928 18992
rect 74988 18932 74994 18992
rect 74798 17872 74804 17932
rect 74864 17872 74870 17932
rect 73660 17670 73666 17730
rect 73726 17670 73732 17730
rect 71922 17611 72410 17617
rect 71922 17577 71934 17611
rect 72398 17577 72410 17611
rect 71922 17571 72410 17577
rect 72940 17611 73428 17617
rect 72940 17577 72952 17611
rect 73416 17577 73428 17611
rect 72940 17571 73428 17577
rect 71632 17492 71640 17518
rect 70656 16942 70674 16968
rect 69886 16883 70374 16889
rect 69886 16849 69898 16883
rect 70362 16849 70374 16883
rect 69886 16843 70374 16849
rect 70102 16788 70162 16843
rect 64002 16728 70162 16788
rect 70614 16782 70674 16942
rect 71634 16942 71640 17492
rect 71674 17492 71692 17518
rect 72652 17518 72698 17530
rect 71674 16942 71680 17492
rect 72652 16964 72658 17518
rect 71634 16930 71680 16942
rect 72650 16942 72658 16964
rect 72692 16964 72698 17518
rect 73666 17518 73726 17670
rect 73958 17611 74446 17617
rect 73958 17577 73970 17611
rect 74434 17577 74446 17611
rect 73958 17571 74446 17577
rect 73666 17488 73676 17518
rect 73670 16980 73676 17488
rect 72692 16942 72710 16964
rect 71122 16889 71182 16896
rect 70904 16883 71392 16889
rect 70904 16849 70916 16883
rect 71380 16849 71392 16883
rect 70904 16843 71392 16849
rect 71922 16883 72410 16889
rect 71922 16849 71934 16883
rect 72398 16849 72410 16883
rect 71922 16843 72410 16849
rect 70608 16722 70614 16782
rect 70674 16722 70680 16782
rect 71122 16670 71182 16843
rect 72142 16670 72202 16843
rect 72650 16782 72710 16942
rect 73664 16942 73676 16980
rect 73710 17488 73726 17518
rect 74688 17518 74734 17530
rect 73710 16980 73716 17488
rect 73710 16942 73724 16980
rect 74688 16968 74694 17518
rect 72940 16883 73428 16889
rect 72940 16849 72952 16883
rect 73416 16849 73428 16883
rect 72940 16843 73428 16849
rect 72644 16722 72650 16782
rect 72710 16722 72716 16782
rect 73144 16670 73204 16843
rect 73664 16786 73724 16942
rect 74680 16942 74694 16968
rect 74728 16968 74734 17518
rect 74728 16942 74740 16968
rect 73958 16883 74446 16889
rect 73958 16849 73970 16883
rect 74434 16849 74446 16883
rect 73958 16843 74446 16849
rect 74178 16786 74238 16843
rect 74680 16786 74740 16942
rect 73664 16726 74740 16786
rect 71122 16610 73204 16670
rect 63478 16452 63484 16512
rect 63544 16452 63550 16512
rect 71122 16398 71182 16610
rect 75088 16512 75148 21440
rect 75240 20244 75300 22100
rect 75234 20184 75240 20244
rect 75300 20184 75306 20244
rect 76666 16642 76672 30072
rect 76772 16642 76778 30072
rect 75082 16452 75088 16512
rect 75148 16452 75154 16512
rect 62964 16338 71182 16398
rect 53780 16228 60994 16288
rect 53720 16222 53780 16228
rect 76666 16128 76778 16642
rect 52322 16122 76778 16128
rect 52322 16022 52428 16122
rect 76672 16022 76778 16122
rect 52322 16016 76778 16022
rect 49084 15700 49228 15992
rect 37958 15392 49228 15700
rect -3042 15198 9310 15392
rect 37958 15198 50310 15392
rect -3042 15192 35878 15198
rect -3042 15092 -1272 15192
rect 35772 15092 35878 15192
rect -3042 15086 35878 15092
rect -3042 15070 9308 15086
rect -1378 14548 -1266 15070
rect 12838 15012 12898 15018
rect 13160 14962 13166 15022
rect 13226 14962 13232 15022
rect 13286 15014 13346 15020
rect 12226 14816 12232 14876
rect 12292 14816 12298 14876
rect 12346 14818 12352 14878
rect 12412 14818 12418 14878
rect 12486 14836 12492 14896
rect 12552 14836 12558 14896
rect 12714 14852 12720 14912
rect 12780 14852 12786 14912
rect 12094 14688 12100 14748
rect 12160 14688 12166 14748
rect -3432 14300 -1262 14548
rect -3432 13782 -2276 14300
rect -1748 13782 -1372 14300
rect -3432 13306 -1372 13782
rect -3432 1924 -3342 13306
rect -2908 1924 -1372 13306
rect -3432 1842 -1372 1924
rect -1378 40 -1372 1842
rect -1272 1842 -1262 14300
rect 9382 14090 9388 14150
rect 9448 14090 9454 14150
rect 9388 14046 9448 14090
rect 1754 13986 9448 14046
rect 1754 13846 1814 13986
rect 2264 13936 2324 13986
rect 2048 13930 2536 13936
rect 2048 13896 2060 13930
rect 2524 13896 2536 13930
rect 2048 13890 2536 13896
rect 1754 13816 1766 13846
rect 1760 13288 1766 13816
rect 1750 13270 1766 13288
rect 1800 13816 1814 13846
rect 2770 13846 2830 13986
rect 3272 13936 3332 13986
rect 4300 13936 4360 13986
rect 3066 13930 3554 13936
rect 3066 13896 3078 13930
rect 3542 13896 3554 13930
rect 3066 13890 3554 13896
rect 4084 13930 4572 13936
rect 4084 13896 4096 13930
rect 4560 13896 4572 13930
rect 4084 13890 4572 13896
rect 2770 13822 2784 13846
rect 1800 13288 1806 13816
rect 2778 13292 2784 13822
rect 1800 13270 1810 13288
rect 1750 13028 1810 13270
rect 2770 13270 2784 13292
rect 2818 13822 2830 13846
rect 3796 13846 3842 13858
rect 2818 13292 2824 13822
rect 3796 13294 3802 13846
rect 2818 13270 2830 13292
rect 2048 13220 2536 13226
rect 2048 13186 2060 13220
rect 2524 13186 2536 13220
rect 2048 13180 2536 13186
rect 2264 13118 2324 13180
rect 2048 13112 2536 13118
rect 2048 13078 2060 13112
rect 2524 13078 2536 13112
rect 2048 13072 2536 13078
rect 1750 12998 1766 13028
rect 1760 12474 1766 12998
rect 1752 12452 1766 12474
rect 1800 12998 1810 13028
rect 2770 13028 2830 13270
rect 3790 13270 3802 13294
rect 3836 13294 3842 13846
rect 4808 13846 4868 13986
rect 5314 13936 5374 13986
rect 6328 13936 6388 13986
rect 5102 13930 5590 13936
rect 5102 13896 5114 13930
rect 5578 13896 5590 13930
rect 5102 13890 5590 13896
rect 6120 13930 6608 13936
rect 6120 13896 6132 13930
rect 6596 13896 6608 13930
rect 6120 13890 6608 13896
rect 4808 13808 4820 13846
rect 3836 13270 3850 13294
rect 4814 13290 4820 13808
rect 3066 13220 3554 13226
rect 3066 13186 3078 13220
rect 3542 13186 3554 13220
rect 3066 13180 3554 13186
rect 3268 13118 3328 13180
rect 3066 13112 3554 13118
rect 3066 13078 3078 13112
rect 3542 13078 3554 13112
rect 3066 13072 3554 13078
rect 2770 13002 2784 13028
rect 1800 12474 1806 12998
rect 2778 12478 2784 13002
rect 1800 12452 1812 12474
rect 1752 12210 1812 12452
rect 2772 12452 2784 12478
rect 2818 13002 2830 13028
rect 3790 13028 3850 13270
rect 4808 13270 4820 13290
rect 4854 13808 4868 13846
rect 5832 13846 5878 13858
rect 6844 13846 6904 13986
rect 7360 13936 7420 13986
rect 8366 13936 8426 13986
rect 7138 13930 7626 13936
rect 7138 13896 7150 13930
rect 7614 13896 7626 13930
rect 7138 13890 7626 13896
rect 8156 13930 8644 13936
rect 8156 13896 8168 13930
rect 8632 13896 8644 13930
rect 8156 13890 8644 13896
rect 4854 13290 4860 13808
rect 5832 13298 5838 13846
rect 4854 13270 4868 13290
rect 4084 13220 4572 13226
rect 4084 13186 4096 13220
rect 4560 13186 4572 13220
rect 4084 13180 4572 13186
rect 4298 13118 4358 13180
rect 4084 13112 4572 13118
rect 4084 13078 4096 13112
rect 4560 13078 4572 13112
rect 4084 13072 4572 13078
rect 3790 13004 3802 13028
rect 2818 12478 2824 13002
rect 3796 12480 3802 13004
rect 2818 12452 2832 12478
rect 2048 12402 2536 12408
rect 2048 12368 2060 12402
rect 2524 12368 2536 12402
rect 2048 12362 2536 12368
rect 2264 12300 2324 12362
rect 2048 12294 2536 12300
rect 2048 12260 2060 12294
rect 2524 12260 2536 12294
rect 2048 12254 2536 12260
rect 1752 12184 1766 12210
rect 1760 11646 1766 12184
rect 1752 11634 1766 11646
rect 1800 12184 1812 12210
rect 2772 12210 2832 12452
rect 3792 12452 3802 12480
rect 3836 13004 3850 13028
rect 4808 13028 4868 13270
rect 5828 13270 5838 13298
rect 5872 13298 5878 13846
rect 6842 13812 6856 13846
rect 6844 13800 6856 13812
rect 5872 13270 5888 13298
rect 6850 13290 6856 13800
rect 5102 13220 5590 13226
rect 5102 13186 5114 13220
rect 5578 13186 5590 13220
rect 5102 13180 5590 13186
rect 5300 13118 5360 13180
rect 5102 13112 5590 13118
rect 5102 13078 5114 13112
rect 5578 13078 5590 13112
rect 5102 13072 5590 13078
rect 3836 12480 3842 13004
rect 4808 13000 4820 13028
rect 3836 12452 3852 12480
rect 4814 12476 4820 13000
rect 3066 12402 3554 12408
rect 3066 12368 3078 12402
rect 3542 12368 3554 12402
rect 3066 12362 3554 12368
rect 3280 12300 3340 12362
rect 3066 12294 3554 12300
rect 3066 12260 3078 12294
rect 3542 12260 3554 12294
rect 3066 12254 3554 12260
rect 2772 12188 2784 12210
rect 1800 11646 1806 12184
rect 2778 11650 2784 12188
rect 1800 11634 1812 11646
rect 1752 11392 1812 11634
rect 2772 11634 2784 11650
rect 2818 12188 2832 12210
rect 3792 12210 3852 12452
rect 4810 12452 4820 12476
rect 4854 13000 4868 13028
rect 5828 13028 5888 13270
rect 6840 13270 6856 13290
rect 6890 13800 6904 13846
rect 7868 13846 7914 13858
rect 6890 13290 6896 13800
rect 7868 13290 7874 13846
rect 6890 13270 6900 13290
rect 6120 13220 6608 13226
rect 6120 13186 6132 13220
rect 6596 13186 6608 13220
rect 6120 13180 6608 13186
rect 6330 13118 6390 13180
rect 6120 13112 6608 13118
rect 6120 13078 6132 13112
rect 6596 13078 6608 13112
rect 6120 13072 6608 13078
rect 5828 13008 5838 13028
rect 4854 12476 4860 13000
rect 5832 12484 5838 13008
rect 4854 12452 4870 12476
rect 4084 12402 4572 12408
rect 4084 12368 4096 12402
rect 4560 12368 4572 12402
rect 4084 12362 4572 12368
rect 4298 12300 4358 12362
rect 4084 12294 4572 12300
rect 4084 12260 4096 12294
rect 4560 12260 4572 12294
rect 4084 12254 4572 12260
rect 3792 12190 3802 12210
rect 2818 11650 2824 12188
rect 3796 11652 3802 12190
rect 2818 11634 2832 11650
rect 2048 11584 2536 11590
rect 2048 11550 2060 11584
rect 2524 11550 2536 11584
rect 2048 11544 2536 11550
rect 2258 11482 2318 11544
rect 2048 11476 2536 11482
rect 2048 11442 2060 11476
rect 2524 11442 2536 11476
rect 2048 11436 2536 11442
rect 1752 11356 1766 11392
rect 1760 10834 1766 11356
rect 1752 10816 1766 10834
rect 1800 11356 1812 11392
rect 2772 11392 2832 11634
rect 3792 11634 3802 11652
rect 3836 12190 3852 12210
rect 4810 12210 4870 12452
rect 5830 12452 5838 12484
rect 5872 13008 5888 13028
rect 6840 13028 6900 13270
rect 7862 13270 7874 13290
rect 7908 13290 7914 13846
rect 8878 13846 8938 13986
rect 9388 13936 9448 13986
rect 10908 13956 10914 14016
rect 10974 13956 10980 14016
rect 9174 13930 9662 13936
rect 9174 13896 9186 13930
rect 9650 13896 9662 13930
rect 9174 13890 9662 13896
rect 10192 13930 10680 13936
rect 10192 13896 10204 13930
rect 10668 13896 10680 13930
rect 10192 13890 10680 13896
rect 8878 13810 8892 13846
rect 8886 13290 8892 13810
rect 7908 13270 7922 13290
rect 7138 13220 7626 13226
rect 7138 13186 7150 13220
rect 7614 13186 7626 13220
rect 7138 13180 7626 13186
rect 7346 13118 7406 13180
rect 7138 13112 7626 13118
rect 7138 13078 7150 13112
rect 7614 13078 7626 13112
rect 7138 13072 7626 13078
rect 5872 12484 5878 13008
rect 6840 13000 6856 13028
rect 5872 12452 5890 12484
rect 6850 12476 6856 13000
rect 5102 12402 5590 12408
rect 5102 12368 5114 12402
rect 5578 12368 5590 12402
rect 5102 12362 5590 12368
rect 5300 12300 5360 12362
rect 5102 12294 5590 12300
rect 5102 12260 5114 12294
rect 5578 12260 5590 12294
rect 5102 12254 5590 12260
rect 3836 11652 3842 12190
rect 4810 12186 4820 12210
rect 3836 11634 3852 11652
rect 4814 11648 4820 12186
rect 3066 11584 3554 11590
rect 3066 11550 3078 11584
rect 3542 11550 3554 11584
rect 3066 11544 3554 11550
rect 3280 11482 3340 11544
rect 3066 11476 3554 11482
rect 3066 11442 3078 11476
rect 3542 11442 3554 11476
rect 3066 11436 3554 11442
rect 2772 11360 2784 11392
rect 1800 10834 1806 11356
rect 2778 10838 2784 11360
rect 1800 10816 1812 10834
rect 1752 10574 1812 10816
rect 2772 10816 2784 10838
rect 2818 11360 2832 11392
rect 3792 11392 3852 11634
rect 4810 11634 4820 11648
rect 4854 12186 4870 12210
rect 5830 12210 5890 12452
rect 6842 12452 6856 12476
rect 6890 13000 6900 13028
rect 7862 13028 7922 13270
rect 8882 13270 8892 13290
rect 8926 13810 8938 13846
rect 9904 13846 9950 13858
rect 8926 13290 8932 13810
rect 9904 13294 9910 13846
rect 8926 13270 8942 13290
rect 8156 13220 8644 13226
rect 8156 13186 8168 13220
rect 8632 13186 8644 13220
rect 8156 13180 8644 13186
rect 8368 13118 8428 13180
rect 8156 13112 8644 13118
rect 8156 13078 8168 13112
rect 8632 13078 8644 13112
rect 8156 13072 8644 13078
rect 7862 13000 7874 13028
rect 6890 12476 6896 13000
rect 7868 12476 7874 13000
rect 6890 12452 6902 12476
rect 6120 12402 6608 12408
rect 6120 12368 6132 12402
rect 6596 12368 6608 12402
rect 6120 12362 6608 12368
rect 6330 12300 6390 12362
rect 6120 12294 6608 12300
rect 6120 12260 6132 12294
rect 6596 12260 6608 12294
rect 6120 12254 6608 12260
rect 5830 12194 5838 12210
rect 4854 11648 4860 12186
rect 5832 11656 5838 12194
rect 4854 11634 4870 11648
rect 4084 11584 4572 11590
rect 4084 11550 4096 11584
rect 4560 11550 4572 11584
rect 4084 11544 4572 11550
rect 4292 11482 4352 11544
rect 4084 11476 4572 11482
rect 4084 11442 4096 11476
rect 4560 11442 4572 11476
rect 4084 11436 4572 11442
rect 3792 11362 3802 11392
rect 2818 10838 2824 11360
rect 3796 10840 3802 11362
rect 2818 10816 2832 10838
rect 2048 10766 2536 10772
rect 2048 10732 2060 10766
rect 2524 10732 2536 10766
rect 2048 10726 2536 10732
rect 2256 10664 2316 10726
rect 2048 10658 2536 10664
rect 2048 10624 2060 10658
rect 2524 10624 2536 10658
rect 2048 10618 2536 10624
rect 1752 10544 1766 10574
rect 1760 10014 1766 10544
rect 1752 9998 1766 10014
rect 1800 10544 1812 10574
rect 2772 10574 2832 10816
rect 3792 10816 3802 10840
rect 3836 11362 3852 11392
rect 4810 11392 4870 11634
rect 5830 11634 5838 11656
rect 5872 12194 5890 12210
rect 6842 12210 6902 12452
rect 7864 12452 7874 12476
rect 7908 13000 7922 13028
rect 8882 13028 8942 13270
rect 9898 13270 9910 13294
rect 9944 13294 9950 13846
rect 10914 13846 10974 13956
rect 10914 13810 10928 13846
rect 9944 13270 9958 13294
rect 10922 13290 10928 13810
rect 9174 13220 9662 13226
rect 9174 13186 9186 13220
rect 9650 13186 9662 13220
rect 9174 13180 9662 13186
rect 9380 13118 9440 13180
rect 9174 13112 9662 13118
rect 9174 13078 9186 13112
rect 9650 13078 9662 13112
rect 9174 13072 9662 13078
rect 8882 13000 8892 13028
rect 7908 12476 7914 13000
rect 8886 12476 8892 13000
rect 7908 12452 7924 12476
rect 7138 12402 7626 12408
rect 7138 12368 7150 12402
rect 7614 12368 7626 12402
rect 7138 12362 7626 12368
rect 7346 12300 7406 12362
rect 7138 12294 7626 12300
rect 7138 12260 7150 12294
rect 7614 12260 7626 12294
rect 7138 12254 7626 12260
rect 5872 11656 5878 12194
rect 6842 12186 6856 12210
rect 5872 11634 5890 11656
rect 6850 11648 6856 12186
rect 5102 11584 5590 11590
rect 5102 11550 5114 11584
rect 5578 11550 5590 11584
rect 5102 11544 5590 11550
rect 5294 11482 5354 11544
rect 5102 11476 5590 11482
rect 5102 11442 5114 11476
rect 5578 11442 5590 11476
rect 5102 11436 5590 11442
rect 3836 10840 3842 11362
rect 4810 11358 4820 11392
rect 3836 10816 3852 10840
rect 4814 10836 4820 11358
rect 3066 10766 3554 10772
rect 3066 10732 3078 10766
rect 3542 10732 3554 10766
rect 3066 10726 3554 10732
rect 3274 10664 3334 10726
rect 3066 10658 3554 10664
rect 3066 10624 3078 10658
rect 3542 10624 3554 10658
rect 3066 10618 3554 10624
rect 2772 10548 2784 10574
rect 1800 10014 1806 10544
rect 2778 10018 2784 10548
rect 1800 9998 1812 10014
rect 1752 9756 1812 9998
rect 2772 9998 2784 10018
rect 2818 10548 2832 10574
rect 3792 10574 3852 10816
rect 4810 10816 4820 10836
rect 4854 11358 4870 11392
rect 5830 11392 5890 11634
rect 6842 11634 6856 11648
rect 6890 12186 6902 12210
rect 7864 12210 7924 12452
rect 8884 12452 8892 12476
rect 8926 13000 8942 13028
rect 9898 13028 9958 13270
rect 10920 13270 10928 13290
rect 10962 13810 10974 13846
rect 10962 13290 10968 13810
rect 10962 13270 10980 13290
rect 10192 13220 10680 13226
rect 10192 13186 10204 13220
rect 10668 13186 10680 13220
rect 10192 13180 10680 13186
rect 10400 13118 10460 13180
rect 10192 13112 10680 13118
rect 10192 13078 10204 13112
rect 10668 13078 10680 13112
rect 10192 13072 10680 13078
rect 9898 13004 9910 13028
rect 8926 12476 8932 13000
rect 9904 12480 9910 13004
rect 8926 12452 8944 12476
rect 8156 12402 8644 12408
rect 8156 12368 8168 12402
rect 8632 12368 8644 12402
rect 8156 12362 8644 12368
rect 8368 12300 8428 12362
rect 8156 12294 8644 12300
rect 8156 12260 8168 12294
rect 8632 12260 8644 12294
rect 8156 12254 8644 12260
rect 7864 12186 7874 12210
rect 6890 11648 6896 12186
rect 7868 11648 7874 12186
rect 6890 11634 6902 11648
rect 6120 11584 6608 11590
rect 6120 11550 6132 11584
rect 6596 11550 6608 11584
rect 6120 11544 6608 11550
rect 6324 11482 6384 11544
rect 6120 11476 6608 11482
rect 6120 11442 6132 11476
rect 6596 11442 6608 11476
rect 6120 11436 6608 11442
rect 5830 11366 5838 11392
rect 4854 10836 4860 11358
rect 5832 10844 5838 11366
rect 4854 10816 4870 10836
rect 4084 10766 4572 10772
rect 4084 10732 4096 10766
rect 4560 10732 4572 10766
rect 4084 10726 4572 10732
rect 4290 10664 4350 10726
rect 4084 10658 4572 10664
rect 4084 10624 4096 10658
rect 4560 10624 4572 10658
rect 4084 10618 4572 10624
rect 3792 10550 3802 10574
rect 2818 10018 2824 10548
rect 3796 10020 3802 10550
rect 2818 9998 2832 10018
rect 2048 9948 2536 9954
rect 2048 9914 2060 9948
rect 2524 9914 2536 9948
rect 2048 9908 2536 9914
rect 2258 9846 2318 9908
rect 2048 9840 2536 9846
rect 2048 9806 2060 9840
rect 2524 9806 2536 9840
rect 2048 9800 2536 9806
rect 1752 9724 1766 9756
rect 1760 9202 1766 9724
rect 1752 9180 1766 9202
rect 1800 9724 1812 9756
rect 2772 9756 2832 9998
rect 3792 9998 3802 10020
rect 3836 10550 3852 10574
rect 4810 10574 4870 10816
rect 5830 10816 5838 10844
rect 5872 11366 5890 11392
rect 6842 11392 6902 11634
rect 7864 11634 7874 11648
rect 7908 12186 7924 12210
rect 8884 12210 8944 12452
rect 9900 12452 9910 12480
rect 9944 13004 9958 13028
rect 10920 13028 10980 13270
rect 9944 12480 9950 13004
rect 10920 13000 10928 13028
rect 9944 12452 9960 12480
rect 9174 12402 9662 12408
rect 9174 12368 9186 12402
rect 9650 12368 9662 12402
rect 9174 12362 9662 12368
rect 9380 12300 9440 12362
rect 9174 12294 9662 12300
rect 9174 12260 9186 12294
rect 9650 12260 9662 12294
rect 9174 12254 9662 12260
rect 8884 12186 8892 12210
rect 7908 11648 7914 12186
rect 8886 11648 8892 12186
rect 7908 11634 7924 11648
rect 7138 11584 7626 11590
rect 7138 11550 7150 11584
rect 7614 11550 7626 11584
rect 7138 11544 7626 11550
rect 7340 11482 7400 11544
rect 7138 11476 7626 11482
rect 7138 11442 7150 11476
rect 7614 11442 7626 11476
rect 7138 11436 7626 11442
rect 5872 10844 5878 11366
rect 6842 11358 6856 11392
rect 5872 10816 5890 10844
rect 6850 10836 6856 11358
rect 5102 10766 5590 10772
rect 5102 10732 5114 10766
rect 5578 10732 5590 10766
rect 5102 10726 5590 10732
rect 5292 10664 5352 10726
rect 5102 10658 5590 10664
rect 5102 10624 5114 10658
rect 5578 10624 5590 10658
rect 5102 10618 5590 10624
rect 3836 10020 3842 10550
rect 4810 10546 4820 10574
rect 3836 9998 3852 10020
rect 4814 10016 4820 10546
rect 3066 9948 3554 9954
rect 3066 9914 3078 9948
rect 3542 9914 3554 9948
rect 3066 9908 3554 9914
rect 3272 9846 3332 9908
rect 3066 9840 3554 9846
rect 3066 9806 3078 9840
rect 3542 9806 3554 9840
rect 3066 9800 3554 9806
rect 2772 9728 2784 9756
rect 1800 9202 1806 9724
rect 2778 9206 2784 9728
rect 1800 9180 1812 9202
rect 1752 8938 1812 9180
rect 2772 9180 2784 9206
rect 2818 9728 2832 9756
rect 3792 9756 3852 9998
rect 4810 9998 4820 10016
rect 4854 10546 4870 10574
rect 5830 10574 5890 10816
rect 6842 10816 6856 10836
rect 6890 11358 6902 11392
rect 7864 11392 7924 11634
rect 8884 11634 8892 11648
rect 8926 12186 8944 12210
rect 9900 12210 9960 12452
rect 10922 12452 10928 13000
rect 10962 13000 10980 13028
rect 10962 12476 10968 13000
rect 10962 12452 10982 12476
rect 10192 12402 10680 12408
rect 10192 12368 10204 12402
rect 10668 12368 10680 12402
rect 10192 12362 10680 12368
rect 10400 12300 10460 12362
rect 10192 12294 10680 12300
rect 10192 12260 10204 12294
rect 10668 12260 10680 12294
rect 10192 12254 10680 12260
rect 9900 12190 9910 12210
rect 8926 11648 8932 12186
rect 9904 11652 9910 12190
rect 8926 11634 8944 11648
rect 8156 11584 8644 11590
rect 8156 11550 8168 11584
rect 8632 11550 8644 11584
rect 8156 11544 8644 11550
rect 8362 11482 8422 11544
rect 8156 11476 8644 11482
rect 8156 11442 8168 11476
rect 8632 11442 8644 11476
rect 8156 11436 8644 11442
rect 7864 11358 7874 11392
rect 6890 10836 6896 11358
rect 7868 10836 7874 11358
rect 6890 10816 6902 10836
rect 6120 10766 6608 10772
rect 6120 10732 6132 10766
rect 6596 10732 6608 10766
rect 6120 10726 6608 10732
rect 6322 10664 6382 10726
rect 6120 10658 6608 10664
rect 6120 10624 6132 10658
rect 6596 10624 6608 10658
rect 6120 10618 6608 10624
rect 5830 10554 5838 10574
rect 4854 10016 4860 10546
rect 5832 10024 5838 10554
rect 4854 9998 4870 10016
rect 4084 9948 4572 9954
rect 4084 9914 4096 9948
rect 4560 9914 4572 9948
rect 4084 9908 4572 9914
rect 4292 9846 4352 9908
rect 4084 9840 4572 9846
rect 4084 9806 4096 9840
rect 4560 9806 4572 9840
rect 4084 9800 4572 9806
rect 3792 9730 3802 9756
rect 2818 9206 2824 9728
rect 3796 9208 3802 9730
rect 2818 9180 2832 9206
rect 2048 9130 2536 9136
rect 2048 9096 2060 9130
rect 2524 9096 2536 9130
rect 2048 9090 2536 9096
rect 2260 9028 2320 9090
rect 2048 9022 2536 9028
rect 2048 8988 2060 9022
rect 2524 8988 2536 9022
rect 2048 8982 2536 8988
rect 1752 8912 1766 8938
rect 1760 8384 1766 8912
rect 1752 8362 1766 8384
rect 1800 8912 1812 8938
rect 2772 8938 2832 9180
rect 3792 9180 3802 9208
rect 3836 9730 3852 9756
rect 4810 9756 4870 9998
rect 5830 9998 5838 10024
rect 5872 10554 5890 10574
rect 6842 10574 6902 10816
rect 7864 10816 7874 10836
rect 7908 11358 7924 11392
rect 8884 11392 8944 11634
rect 9900 11634 9910 11652
rect 9944 12190 9960 12210
rect 10922 12210 10982 12452
rect 9944 11652 9950 12190
rect 9944 11634 9960 11652
rect 9174 11584 9662 11590
rect 9174 11550 9186 11584
rect 9650 11550 9662 11584
rect 9174 11544 9662 11550
rect 9374 11482 9434 11544
rect 9174 11476 9662 11482
rect 9174 11442 9186 11476
rect 9650 11442 9662 11476
rect 9174 11436 9662 11442
rect 8884 11358 8892 11392
rect 7908 10836 7914 11358
rect 8886 10836 8892 11358
rect 7908 10816 7924 10836
rect 7138 10766 7626 10772
rect 7138 10732 7150 10766
rect 7614 10732 7626 10766
rect 7138 10726 7626 10732
rect 7338 10664 7398 10726
rect 7138 10658 7626 10664
rect 7138 10624 7150 10658
rect 7614 10624 7626 10658
rect 7138 10618 7626 10624
rect 5872 10024 5878 10554
rect 6842 10546 6856 10574
rect 5872 9998 5890 10024
rect 6850 10016 6856 10546
rect 5102 9948 5590 9954
rect 5102 9914 5114 9948
rect 5578 9914 5590 9948
rect 5102 9908 5590 9914
rect 5294 9846 5354 9908
rect 5102 9840 5590 9846
rect 5102 9806 5114 9840
rect 5578 9806 5590 9840
rect 5102 9800 5590 9806
rect 3836 9208 3842 9730
rect 4810 9726 4820 9756
rect 3836 9180 3852 9208
rect 4814 9204 4820 9726
rect 3066 9130 3554 9136
rect 3066 9096 3078 9130
rect 3542 9096 3554 9130
rect 3066 9090 3554 9096
rect 3274 9028 3334 9090
rect 3066 9022 3554 9028
rect 3066 8988 3078 9022
rect 3542 8988 3554 9022
rect 3066 8982 3554 8988
rect 2772 8916 2784 8938
rect 1800 8384 1806 8912
rect 2778 8388 2784 8916
rect 1800 8362 1812 8384
rect 1752 8120 1812 8362
rect 2772 8362 2784 8388
rect 2818 8916 2832 8938
rect 3792 8938 3852 9180
rect 4810 9180 4820 9204
rect 4854 9726 4870 9756
rect 5830 9756 5890 9998
rect 6842 9998 6856 10016
rect 6890 10546 6902 10574
rect 7864 10574 7924 10816
rect 8884 10816 8892 10836
rect 8926 11358 8944 11392
rect 9900 11392 9960 11634
rect 10922 11634 10928 12210
rect 10962 12186 10982 12210
rect 10962 11648 10968 12186
rect 10962 11634 10982 11648
rect 10192 11584 10680 11590
rect 10192 11550 10204 11584
rect 10668 11550 10680 11584
rect 10192 11544 10680 11550
rect 10394 11482 10454 11544
rect 10192 11476 10680 11482
rect 10192 11442 10204 11476
rect 10668 11442 10680 11476
rect 10192 11436 10680 11442
rect 9900 11362 9910 11392
rect 8926 10836 8932 11358
rect 9904 10840 9910 11362
rect 8926 10816 8944 10836
rect 8156 10766 8644 10772
rect 8156 10732 8168 10766
rect 8632 10732 8644 10766
rect 8156 10726 8644 10732
rect 8360 10664 8420 10726
rect 8156 10658 8644 10664
rect 8156 10624 8168 10658
rect 8632 10624 8644 10658
rect 8156 10618 8644 10624
rect 7864 10546 7874 10574
rect 6890 10016 6896 10546
rect 7868 10016 7874 10546
rect 6890 9998 6902 10016
rect 6120 9948 6608 9954
rect 6120 9914 6132 9948
rect 6596 9914 6608 9948
rect 6120 9908 6608 9914
rect 6324 9846 6384 9908
rect 6120 9840 6608 9846
rect 6120 9806 6132 9840
rect 6596 9806 6608 9840
rect 6120 9800 6608 9806
rect 5830 9734 5838 9756
rect 4854 9204 4860 9726
rect 5832 9212 5838 9734
rect 4854 9180 4870 9204
rect 4084 9130 4572 9136
rect 4084 9096 4096 9130
rect 4560 9096 4572 9130
rect 4084 9090 4572 9096
rect 4294 9028 4354 9090
rect 4084 9022 4572 9028
rect 4084 8988 4096 9022
rect 4560 8988 4572 9022
rect 4084 8982 4572 8988
rect 3792 8918 3802 8938
rect 2818 8388 2824 8916
rect 3796 8390 3802 8918
rect 2818 8362 2832 8388
rect 2048 8312 2536 8318
rect 2048 8278 2060 8312
rect 2524 8278 2536 8312
rect 2048 8272 2536 8278
rect 2262 8210 2322 8272
rect 2048 8204 2536 8210
rect 2048 8170 2060 8204
rect 2524 8170 2536 8204
rect 2048 8164 2536 8170
rect 1752 8094 1766 8120
rect 1760 7544 1766 8094
rect 1800 8094 1812 8120
rect 2772 8120 2832 8362
rect 3792 8362 3802 8390
rect 3836 8918 3852 8938
rect 4810 8938 4870 9180
rect 5830 9180 5838 9212
rect 5872 9734 5890 9756
rect 6842 9756 6902 9998
rect 7864 9998 7874 10016
rect 7908 10546 7924 10574
rect 8884 10574 8944 10816
rect 9900 10816 9910 10840
rect 9944 11362 9960 11392
rect 10922 11392 10982 11634
rect 9944 10840 9950 11362
rect 9944 10816 9960 10840
rect 9174 10766 9662 10772
rect 9174 10732 9186 10766
rect 9650 10732 9662 10766
rect 9174 10726 9662 10732
rect 9372 10664 9432 10726
rect 9174 10658 9662 10664
rect 9174 10624 9186 10658
rect 9650 10624 9662 10658
rect 9174 10618 9662 10624
rect 8884 10546 8892 10574
rect 7908 10016 7914 10546
rect 8886 10016 8892 10546
rect 7908 9998 7924 10016
rect 7138 9948 7626 9954
rect 7138 9914 7150 9948
rect 7614 9914 7626 9948
rect 7138 9908 7626 9914
rect 7340 9846 7400 9908
rect 7138 9840 7626 9846
rect 7138 9806 7150 9840
rect 7614 9806 7626 9840
rect 7138 9800 7626 9806
rect 5872 9212 5878 9734
rect 6842 9726 6856 9756
rect 5872 9180 5890 9212
rect 6850 9204 6856 9726
rect 5102 9130 5590 9136
rect 5102 9096 5114 9130
rect 5578 9096 5590 9130
rect 5102 9090 5590 9096
rect 5296 9028 5356 9090
rect 5102 9022 5590 9028
rect 5102 8988 5114 9022
rect 5578 8988 5590 9022
rect 5102 8982 5590 8988
rect 3836 8390 3842 8918
rect 4810 8914 4820 8938
rect 3836 8362 3852 8390
rect 4814 8386 4820 8914
rect 3066 8312 3554 8318
rect 3066 8278 3078 8312
rect 3542 8278 3554 8312
rect 3066 8272 3554 8278
rect 3276 8210 3336 8272
rect 3066 8204 3554 8210
rect 3066 8170 3078 8204
rect 3542 8170 3554 8204
rect 3066 8164 3554 8170
rect 2772 8098 2784 8120
rect 1800 7544 1806 8094
rect 1760 7532 1806 7544
rect 2778 7544 2784 8098
rect 2818 8098 2832 8120
rect 3792 8120 3852 8362
rect 4810 8362 4820 8386
rect 4854 8914 4870 8938
rect 5830 8938 5890 9180
rect 6842 9180 6856 9204
rect 6890 9726 6902 9756
rect 7864 9756 7924 9998
rect 8884 9998 8892 10016
rect 8926 10546 8944 10574
rect 9900 10574 9960 10816
rect 10922 10816 10928 11392
rect 10962 11358 10982 11392
rect 10962 10836 10968 11358
rect 10962 10816 10982 10836
rect 10192 10766 10680 10772
rect 10192 10732 10204 10766
rect 10668 10732 10680 10766
rect 10192 10726 10680 10732
rect 10392 10664 10452 10726
rect 10192 10658 10680 10664
rect 10192 10624 10204 10658
rect 10668 10624 10680 10658
rect 10192 10618 10680 10624
rect 9900 10550 9910 10574
rect 8926 10016 8932 10546
rect 9904 10020 9910 10550
rect 8926 9998 8944 10016
rect 8156 9948 8644 9954
rect 8156 9914 8168 9948
rect 8632 9914 8644 9948
rect 8156 9908 8644 9914
rect 8362 9846 8422 9908
rect 8156 9840 8644 9846
rect 8156 9806 8168 9840
rect 8632 9806 8644 9840
rect 8156 9800 8644 9806
rect 7864 9726 7874 9756
rect 6890 9204 6896 9726
rect 7868 9204 7874 9726
rect 6890 9180 6902 9204
rect 6120 9130 6608 9136
rect 6120 9096 6132 9130
rect 6596 9096 6608 9130
rect 6120 9090 6608 9096
rect 6326 9028 6386 9090
rect 6120 9022 6608 9028
rect 6120 8988 6132 9022
rect 6596 8988 6608 9022
rect 6120 8982 6608 8988
rect 5830 8922 5838 8938
rect 4854 8386 4860 8914
rect 5832 8394 5838 8922
rect 4854 8362 4870 8386
rect 4084 8312 4572 8318
rect 4084 8278 4096 8312
rect 4560 8278 4572 8312
rect 4084 8272 4572 8278
rect 4296 8210 4356 8272
rect 4084 8204 4572 8210
rect 4084 8170 4096 8204
rect 4560 8170 4572 8204
rect 4084 8164 4572 8170
rect 3792 8100 3802 8120
rect 2818 7544 2824 8098
rect 3796 7590 3802 8100
rect 2778 7532 2824 7544
rect 3786 7544 3802 7590
rect 3836 8100 3852 8120
rect 4810 8120 4870 8362
rect 5830 8362 5838 8394
rect 5872 8922 5890 8938
rect 6842 8938 6902 9180
rect 7864 9180 7874 9204
rect 7908 9726 7924 9756
rect 8884 9756 8944 9998
rect 9900 9998 9910 10020
rect 9944 10550 9960 10574
rect 10922 10574 10982 10816
rect 9944 10020 9950 10550
rect 9944 9998 9960 10020
rect 9174 9948 9662 9954
rect 9174 9914 9186 9948
rect 9650 9914 9662 9948
rect 9174 9908 9662 9914
rect 9374 9846 9434 9908
rect 9174 9840 9662 9846
rect 9174 9806 9186 9840
rect 9650 9806 9662 9840
rect 9174 9800 9662 9806
rect 8884 9726 8892 9756
rect 7908 9204 7914 9726
rect 8886 9204 8892 9726
rect 7908 9180 7924 9204
rect 7138 9130 7626 9136
rect 7138 9096 7150 9130
rect 7614 9096 7626 9130
rect 7138 9090 7626 9096
rect 7342 9028 7402 9090
rect 7138 9022 7626 9028
rect 7138 8988 7150 9022
rect 7614 8988 7626 9022
rect 7138 8982 7626 8988
rect 5872 8394 5878 8922
rect 6842 8914 6856 8938
rect 5872 8362 5890 8394
rect 6850 8386 6856 8914
rect 5102 8312 5590 8318
rect 5102 8278 5114 8312
rect 5578 8278 5590 8312
rect 5102 8272 5590 8278
rect 5298 8210 5358 8272
rect 5102 8204 5590 8210
rect 5102 8170 5114 8204
rect 5578 8170 5590 8204
rect 5102 8164 5590 8170
rect 3836 7590 3842 8100
rect 4810 8096 4820 8120
rect 3836 7544 3846 7590
rect 2048 7494 2536 7500
rect 2048 7460 2060 7494
rect 2524 7460 2536 7494
rect 2048 7454 2536 7460
rect 3066 7494 3554 7500
rect 3066 7460 3078 7494
rect 3542 7460 3554 7494
rect 3066 7454 3554 7460
rect 3786 7370 3846 7544
rect 4814 7544 4820 8096
rect 4854 8096 4870 8120
rect 5830 8120 5890 8362
rect 6842 8362 6856 8386
rect 6890 8914 6902 8938
rect 7864 8938 7924 9180
rect 8884 9180 8892 9204
rect 8926 9726 8944 9756
rect 9900 9756 9960 9998
rect 10922 9998 10928 10574
rect 10962 10546 10982 10574
rect 10962 10016 10968 10546
rect 10962 9998 10982 10016
rect 10192 9948 10680 9954
rect 10192 9914 10204 9948
rect 10668 9914 10680 9948
rect 10192 9908 10680 9914
rect 10394 9846 10454 9908
rect 10192 9840 10680 9846
rect 10192 9806 10204 9840
rect 10668 9806 10680 9840
rect 10192 9800 10680 9806
rect 9900 9730 9910 9756
rect 8926 9204 8932 9726
rect 9904 9208 9910 9730
rect 8926 9180 8944 9204
rect 8156 9130 8644 9136
rect 8156 9096 8168 9130
rect 8632 9096 8644 9130
rect 8156 9090 8644 9096
rect 8364 9028 8424 9090
rect 8156 9022 8644 9028
rect 8156 8988 8168 9022
rect 8632 8988 8644 9022
rect 8156 8982 8644 8988
rect 7864 8914 7874 8938
rect 6890 8386 6896 8914
rect 7868 8386 7874 8914
rect 6890 8362 6902 8386
rect 6120 8312 6608 8318
rect 6120 8278 6132 8312
rect 6596 8278 6608 8312
rect 6120 8272 6608 8278
rect 6328 8210 6388 8272
rect 6120 8204 6608 8210
rect 6120 8170 6132 8204
rect 6596 8170 6608 8204
rect 6120 8164 6608 8170
rect 5830 8104 5838 8120
rect 4854 7544 4860 8096
rect 5832 7592 5838 8104
rect 4814 7532 4860 7544
rect 5824 7544 5838 7592
rect 5872 8104 5890 8120
rect 6842 8120 6902 8362
rect 7864 8362 7874 8386
rect 7908 8914 7924 8938
rect 8884 8938 8944 9180
rect 9900 9180 9910 9208
rect 9944 9730 9960 9756
rect 10922 9756 10982 9998
rect 9944 9208 9950 9730
rect 9944 9180 9960 9208
rect 9174 9130 9662 9136
rect 9174 9096 9186 9130
rect 9650 9096 9662 9130
rect 9174 9090 9662 9096
rect 9376 9028 9436 9090
rect 9174 9022 9662 9028
rect 9174 8988 9186 9022
rect 9650 8988 9662 9022
rect 9174 8982 9662 8988
rect 8884 8914 8892 8938
rect 7908 8386 7914 8914
rect 8886 8386 8892 8914
rect 7908 8362 7924 8386
rect 7138 8312 7626 8318
rect 7138 8278 7150 8312
rect 7614 8278 7626 8312
rect 7138 8272 7626 8278
rect 7344 8210 7404 8272
rect 7138 8204 7626 8210
rect 7138 8170 7150 8204
rect 7614 8170 7626 8204
rect 7138 8164 7626 8170
rect 5872 7592 5878 8104
rect 6842 8096 6856 8120
rect 5872 7544 5884 7592
rect 4084 7494 4572 7500
rect 4084 7460 4096 7494
rect 4560 7460 4572 7494
rect 4084 7454 4572 7460
rect 5102 7494 5590 7500
rect 5102 7460 5114 7494
rect 5578 7460 5590 7494
rect 5102 7454 5590 7460
rect 5824 7370 5884 7544
rect 6850 7544 6856 8096
rect 6890 8096 6902 8120
rect 7864 8120 7924 8362
rect 8884 8362 8892 8386
rect 8926 8914 8944 8938
rect 9900 8938 9960 9180
rect 10922 9180 10928 9756
rect 10962 9726 10982 9756
rect 10962 9204 10968 9726
rect 10962 9180 10982 9204
rect 10192 9130 10680 9136
rect 10192 9096 10204 9130
rect 10668 9096 10680 9130
rect 10192 9090 10680 9096
rect 10396 9028 10456 9090
rect 10192 9022 10680 9028
rect 10192 8988 10204 9022
rect 10668 8988 10680 9022
rect 10192 8982 10680 8988
rect 9900 8918 9910 8938
rect 8926 8386 8932 8914
rect 9904 8390 9910 8918
rect 8926 8362 8944 8386
rect 8156 8312 8644 8318
rect 8156 8278 8168 8312
rect 8632 8278 8644 8312
rect 8156 8272 8644 8278
rect 8366 8210 8426 8272
rect 8156 8204 8644 8210
rect 8156 8170 8168 8204
rect 8632 8170 8644 8204
rect 8156 8164 8644 8170
rect 7864 8096 7874 8120
rect 6890 7544 6896 8096
rect 7868 7588 7874 8096
rect 6850 7532 6896 7544
rect 7860 7544 7874 7588
rect 7908 8096 7924 8120
rect 8884 8120 8944 8362
rect 9900 8362 9910 8390
rect 9944 8918 9960 8938
rect 10922 8938 10982 9180
rect 9944 8390 9950 8918
rect 9944 8362 9960 8390
rect 9174 8312 9662 8318
rect 9174 8278 9186 8312
rect 9650 8278 9662 8312
rect 9174 8272 9662 8278
rect 9378 8210 9438 8272
rect 9174 8204 9662 8210
rect 9174 8170 9186 8204
rect 9650 8170 9662 8204
rect 9174 8164 9662 8170
rect 8884 8096 8892 8120
rect 7908 7588 7914 8096
rect 7908 7544 7920 7588
rect 6120 7494 6608 7500
rect 6120 7460 6132 7494
rect 6596 7460 6608 7494
rect 6120 7454 6608 7460
rect 7138 7494 7626 7500
rect 7138 7460 7150 7494
rect 7614 7460 7626 7494
rect 7138 7454 7626 7460
rect 7860 7370 7920 7544
rect 8886 7544 8892 8096
rect 8926 8096 8944 8120
rect 9900 8120 9960 8362
rect 10922 8362 10928 8938
rect 10962 8914 10982 8938
rect 10962 8386 10968 8914
rect 10962 8362 10982 8386
rect 10192 8312 10680 8318
rect 10192 8278 10204 8312
rect 10668 8278 10680 8312
rect 10192 8272 10680 8278
rect 10398 8210 10458 8272
rect 10192 8204 10680 8210
rect 10192 8170 10204 8204
rect 10668 8170 10680 8204
rect 10192 8164 10680 8170
rect 9900 8100 9910 8120
rect 8926 7544 8932 8096
rect 9904 7586 9910 8100
rect 8886 7532 8932 7544
rect 9896 7544 9910 7586
rect 9944 8100 9960 8120
rect 10922 8120 10982 8362
rect 9944 7586 9950 8100
rect 10922 7598 10928 8120
rect 9944 7544 9956 7586
rect 8156 7494 8644 7500
rect 8156 7460 8168 7494
rect 8632 7460 8644 7494
rect 8156 7454 8644 7460
rect 9174 7494 9662 7500
rect 9174 7460 9186 7494
rect 9650 7460 9662 7494
rect 9174 7454 9662 7460
rect 9896 7370 9956 7544
rect 10916 7544 10928 7598
rect 10962 8096 10982 8120
rect 10962 7598 10968 8096
rect 10962 7544 10976 7598
rect 12100 7548 12160 14688
rect 10192 7494 10680 7500
rect 10192 7460 10204 7494
rect 10668 7460 10680 7494
rect 10192 7454 10680 7460
rect 10410 7370 10470 7454
rect 10916 7370 10976 7544
rect 12094 7488 12100 7548
rect 12160 7488 12166 7548
rect 3786 7310 12080 7370
rect 7546 6562 7552 6622
rect 7612 6562 7618 6622
rect 1442 6476 1502 6482
rect 5516 6416 5522 6476
rect 5582 6416 5588 6476
rect 282 6288 288 6348
rect 348 6288 354 6348
rect 288 4116 348 6288
rect 1442 6284 1502 6416
rect 2960 6288 2966 6348
rect 3026 6288 3032 6348
rect 3992 6288 3998 6348
rect 4058 6288 4064 6348
rect 426 6224 1502 6284
rect 426 6096 486 6224
rect 934 6186 994 6224
rect 724 6180 1212 6186
rect 724 6146 736 6180
rect 1200 6146 1212 6180
rect 724 6140 1212 6146
rect 426 6050 442 6096
rect 436 5520 442 6050
rect 476 6050 486 6096
rect 1442 6096 1502 6224
rect 2966 6186 3026 6288
rect 3998 6186 4058 6288
rect 1742 6180 2230 6186
rect 1742 6146 1754 6180
rect 2218 6146 2230 6180
rect 1742 6140 2230 6146
rect 2760 6180 3248 6186
rect 2760 6146 2772 6180
rect 3236 6146 3248 6180
rect 2760 6140 3248 6146
rect 3778 6180 4266 6186
rect 3778 6146 3790 6180
rect 4254 6146 4266 6180
rect 3778 6140 4266 6146
rect 4796 6180 5284 6186
rect 4796 6146 4808 6180
rect 5272 6146 5284 6180
rect 4796 6140 5284 6146
rect 1442 6056 1460 6096
rect 476 5520 482 6050
rect 436 5508 482 5520
rect 1454 5520 1460 6056
rect 1494 6056 1502 6096
rect 2472 6096 2518 6108
rect 1494 5520 1500 6056
rect 2472 5584 2478 6096
rect 1454 5508 1500 5520
rect 2464 5520 2478 5584
rect 2512 5584 2518 6096
rect 3490 6096 3536 6108
rect 2512 5520 2524 5584
rect 3490 5566 3496 6096
rect 724 5470 1212 5476
rect 724 5436 736 5470
rect 1200 5436 1212 5470
rect 724 5430 1212 5436
rect 1742 5470 2230 5476
rect 1742 5436 1754 5470
rect 2218 5436 2230 5470
rect 1742 5430 2230 5436
rect 1946 5386 2006 5430
rect 1940 5326 1946 5386
rect 2006 5326 2012 5386
rect 1440 5222 1446 5282
rect 1506 5222 1512 5282
rect 1446 5180 1506 5222
rect 426 5120 1506 5180
rect 426 4984 486 5120
rect 930 5074 990 5120
rect 724 5068 1212 5074
rect 724 5034 736 5068
rect 1200 5034 1212 5068
rect 724 5028 1212 5034
rect 426 4938 442 4984
rect 436 4408 442 4938
rect 476 4938 486 4984
rect 1446 4984 1506 5120
rect 2464 5178 2524 5520
rect 3482 5520 3496 5566
rect 3530 5566 3536 6096
rect 4508 6096 4554 6108
rect 4508 5582 4514 6096
rect 3530 5520 3542 5566
rect 2760 5470 3248 5476
rect 2760 5436 2772 5470
rect 3236 5436 3248 5470
rect 2760 5430 3248 5436
rect 2964 5326 2970 5386
rect 3030 5326 3036 5386
rect 1742 5068 2230 5074
rect 1742 5034 1754 5068
rect 2218 5034 2230 5068
rect 1742 5028 2230 5034
rect 476 4408 482 4938
rect 436 4396 482 4408
rect 1446 4408 1460 4984
rect 1494 4408 1506 4984
rect 724 4358 1212 4364
rect 724 4324 736 4358
rect 1200 4324 1212 4358
rect 724 4318 1212 4324
rect 282 4056 288 4116
rect 348 4056 354 4116
rect 288 1990 348 4056
rect 724 3956 1212 3962
rect 724 3922 736 3956
rect 1200 3922 1212 3956
rect 724 3916 1212 3922
rect 436 3872 482 3884
rect 436 3330 442 3872
rect 430 3296 442 3330
rect 476 3330 482 3872
rect 1446 3872 1506 4408
rect 2464 4984 2524 5118
rect 2970 5074 3030 5326
rect 3482 5282 3542 5520
rect 4500 5520 4514 5582
rect 4548 5582 4554 6096
rect 5522 6096 5582 6416
rect 7052 6288 7058 6348
rect 7118 6288 7124 6348
rect 7058 6186 7118 6288
rect 5814 6180 6302 6186
rect 5814 6146 5826 6180
rect 6290 6146 6302 6180
rect 5814 6140 6302 6146
rect 6832 6180 7320 6186
rect 6832 6146 6844 6180
rect 7308 6146 7320 6180
rect 6832 6140 7320 6146
rect 5522 6032 5532 6096
rect 4548 5520 4560 5582
rect 3778 5470 4266 5476
rect 3778 5436 3790 5470
rect 4254 5436 4266 5470
rect 3778 5430 4266 5436
rect 3996 5326 4002 5386
rect 4062 5326 4068 5386
rect 3476 5222 3482 5282
rect 3542 5222 3548 5282
rect 4002 5074 4062 5326
rect 4500 5178 4560 5520
rect 5526 5520 5532 6032
rect 5566 6032 5582 6096
rect 6544 6096 6590 6108
rect 5566 5520 5572 6032
rect 6544 5592 6550 6096
rect 5526 5508 5572 5520
rect 6532 5520 6550 5592
rect 6584 5592 6590 6096
rect 7552 6096 7612 6562
rect 9576 6416 9582 6476
rect 9642 6416 9648 6476
rect 11760 6416 11766 6476
rect 11826 6416 11832 6476
rect 8048 6288 8054 6348
rect 8114 6288 8120 6348
rect 8054 6186 8114 6288
rect 7850 6180 8338 6186
rect 7850 6146 7862 6180
rect 8326 6146 8338 6180
rect 7850 6140 8338 6146
rect 8868 6180 9356 6186
rect 8868 6146 8880 6180
rect 9344 6146 9356 6180
rect 8868 6140 9356 6146
rect 8054 6138 8114 6140
rect 9582 6108 9642 6416
rect 9886 6180 10374 6186
rect 9886 6146 9898 6180
rect 10362 6146 10374 6180
rect 9886 6140 10374 6146
rect 10904 6180 11392 6186
rect 10904 6146 10916 6180
rect 11380 6146 11392 6180
rect 10904 6140 11392 6146
rect 6584 5520 6592 5592
rect 4796 5470 5284 5476
rect 4796 5436 4808 5470
rect 5272 5436 5284 5470
rect 4796 5430 5284 5436
rect 5814 5470 6302 5476
rect 5814 5436 5826 5470
rect 6290 5436 6302 5470
rect 5814 5430 6302 5436
rect 5002 5386 5062 5430
rect 6022 5386 6082 5430
rect 4996 5326 5002 5386
rect 5062 5326 5068 5386
rect 6016 5326 6022 5386
rect 6082 5326 6088 5386
rect 5512 5222 5518 5282
rect 5578 5222 5584 5282
rect 2760 5068 3248 5074
rect 2760 5034 2772 5068
rect 3236 5034 3248 5068
rect 2760 5028 3248 5034
rect 3778 5068 4266 5074
rect 3778 5034 3790 5068
rect 4254 5034 4266 5068
rect 3778 5028 4266 5034
rect 2464 4408 2478 4984
rect 2512 4408 2524 4984
rect 3490 4984 3536 4996
rect 3490 4446 3496 4984
rect 1742 4358 2230 4364
rect 1742 4324 1754 4358
rect 2218 4324 2230 4358
rect 1742 4318 2230 4324
rect 1938 4116 1998 4318
rect 1932 4056 1938 4116
rect 1998 4056 2004 4116
rect 1938 3962 1998 4056
rect 1742 3956 2230 3962
rect 1742 3922 1754 3956
rect 2218 3922 2230 3956
rect 1742 3916 2230 3922
rect 1446 3800 1460 3872
rect 476 3296 490 3330
rect 1454 3326 1460 3800
rect 430 3164 490 3296
rect 1450 3296 1460 3326
rect 1494 3800 1506 3872
rect 2464 3872 2524 4408
rect 3476 4408 3496 4446
rect 3530 4408 3536 4984
rect 2760 4358 3248 4364
rect 2760 4324 2772 4358
rect 3236 4324 3248 4358
rect 2760 4318 3248 4324
rect 3476 4236 3536 4408
rect 4500 4984 4560 5118
rect 4796 5068 5284 5074
rect 4796 5034 4808 5068
rect 5272 5034 5284 5068
rect 4796 5028 5284 5034
rect 4500 4408 4514 4984
rect 4548 4408 4560 4984
rect 3778 4358 4266 4364
rect 3778 4324 3790 4358
rect 4254 4324 4266 4358
rect 3778 4318 4266 4324
rect 3470 4176 3476 4236
rect 3536 4176 3542 4236
rect 2760 3956 3248 3962
rect 2760 3922 2772 3956
rect 3236 3922 3248 3956
rect 2760 3916 3248 3922
rect 1494 3326 1500 3800
rect 1494 3296 1510 3326
rect 724 3246 1212 3252
rect 724 3212 736 3246
rect 1200 3212 1212 3246
rect 724 3206 1212 3212
rect 922 3164 982 3206
rect 1450 3164 1510 3296
rect 2464 3296 2478 3872
rect 2512 3296 2524 3872
rect 3476 3872 3536 4176
rect 3778 3956 4266 3962
rect 3778 3922 3790 3956
rect 4254 3922 4266 3956
rect 3778 3916 4266 3922
rect 3476 3802 3496 3872
rect 1742 3246 2230 3252
rect 1742 3212 1754 3246
rect 2218 3212 2230 3246
rect 1742 3206 2230 3212
rect 430 3104 1510 3164
rect 1450 3064 1510 3104
rect 2464 3172 2524 3296
rect 3490 3296 3496 3802
rect 3530 3296 3536 3872
rect 3490 3284 3536 3296
rect 4500 3872 4560 4408
rect 5518 4984 5578 5222
rect 6532 5178 6592 5520
rect 7552 5520 7568 6096
rect 7602 5520 7612 6096
rect 8580 6096 8626 6108
rect 8580 5582 8586 6096
rect 6832 5470 7320 5476
rect 6832 5436 6844 5470
rect 7308 5436 7320 5470
rect 6832 5430 7320 5436
rect 7036 5326 7042 5386
rect 7102 5326 7108 5386
rect 6526 5118 6532 5178
rect 6592 5118 6598 5178
rect 5814 5068 6302 5074
rect 5814 5034 5826 5068
rect 6290 5034 6302 5068
rect 5814 5028 6302 5034
rect 5518 4408 5532 4984
rect 5566 4408 5578 4984
rect 4796 4358 5284 4364
rect 4796 4324 4808 4358
rect 5272 4324 5284 4358
rect 4796 4318 5284 4324
rect 5008 4116 5068 4318
rect 5002 4056 5008 4116
rect 5068 4056 5074 4116
rect 5008 3962 5068 4056
rect 4796 3956 5284 3962
rect 4796 3922 4808 3956
rect 5272 3922 5284 3956
rect 4796 3916 5284 3922
rect 4500 3296 4514 3872
rect 4548 3296 4560 3872
rect 5518 3872 5578 4408
rect 6532 4984 6592 5118
rect 7042 5074 7102 5326
rect 7552 5282 7612 5520
rect 8566 5520 8586 5582
rect 8620 5520 8626 6096
rect 9582 6096 9644 6108
rect 9582 6064 9604 6096
rect 7850 5470 8338 5476
rect 7850 5436 7862 5470
rect 8326 5436 8338 5470
rect 7850 5430 8338 5436
rect 8052 5386 8112 5392
rect 7546 5222 7552 5282
rect 7612 5222 7618 5282
rect 8052 5074 8112 5326
rect 8566 5178 8626 5520
rect 9598 5520 9604 6064
rect 9638 5520 9644 6096
rect 10616 6096 10662 6108
rect 10616 5554 10622 6096
rect 9598 5508 9644 5520
rect 10610 5520 10622 5554
rect 10656 5554 10662 6096
rect 11634 6096 11680 6108
rect 11634 5574 11640 6096
rect 10656 5520 10670 5554
rect 8868 5470 9356 5476
rect 8868 5436 8880 5470
rect 9344 5436 9356 5470
rect 8868 5430 9356 5436
rect 9886 5470 10374 5476
rect 9886 5436 9898 5470
rect 10362 5436 10374 5470
rect 9886 5430 10374 5436
rect 9066 5386 9126 5430
rect 10084 5386 10144 5430
rect 9060 5326 9066 5386
rect 9126 5326 9132 5386
rect 10084 5320 10144 5326
rect 10610 5292 10670 5520
rect 11626 5520 11640 5574
rect 11674 5574 11680 6096
rect 11674 5520 11686 5574
rect 10904 5470 11392 5476
rect 10904 5436 10916 5470
rect 11380 5436 11392 5470
rect 10904 5430 11392 5436
rect 11114 5292 11174 5430
rect 11626 5292 11686 5520
rect 9582 5222 9588 5282
rect 9648 5222 9654 5282
rect 10610 5232 11686 5292
rect 6832 5068 7320 5074
rect 6832 5034 6844 5068
rect 7308 5034 7320 5068
rect 6832 5028 7320 5034
rect 7850 5068 8338 5074
rect 7850 5034 7862 5068
rect 8326 5034 8338 5068
rect 7850 5028 8338 5034
rect 6532 4408 6550 4984
rect 6584 4408 6592 4984
rect 7562 4984 7608 4996
rect 7562 4464 7568 4984
rect 5814 4358 6302 4364
rect 5814 4324 5826 4358
rect 6290 4324 6302 4358
rect 5814 4318 6302 4324
rect 6016 4116 6076 4318
rect 6010 4056 6016 4116
rect 6076 4056 6082 4116
rect 6016 3962 6076 4056
rect 5814 3956 6302 3962
rect 5814 3922 5826 3956
rect 6290 3922 6302 3956
rect 5814 3916 6302 3922
rect 5518 3766 5532 3872
rect 5526 3358 5532 3766
rect 2760 3246 3248 3252
rect 2760 3212 2772 3246
rect 3236 3212 3248 3246
rect 2760 3206 3248 3212
rect 3778 3246 4266 3252
rect 3778 3212 3790 3246
rect 4254 3212 4266 3246
rect 3778 3206 4266 3212
rect 1444 3004 1450 3064
rect 1510 3004 1516 3064
rect 1938 2892 1944 2952
rect 2004 2892 2010 2952
rect 1944 2850 2004 2892
rect 724 2844 1212 2850
rect 724 2810 736 2844
rect 1200 2810 1212 2844
rect 724 2804 1212 2810
rect 1742 2844 2230 2850
rect 1742 2810 1754 2844
rect 2218 2810 2230 2844
rect 1742 2804 2230 2810
rect 436 2760 482 2772
rect 436 2226 442 2760
rect 426 2184 442 2226
rect 476 2226 482 2760
rect 1454 2760 1500 2772
rect 476 2184 486 2226
rect 1454 2220 1460 2760
rect 426 2040 486 2184
rect 1444 2184 1460 2220
rect 1494 2220 1500 2760
rect 2464 2760 2524 3112
rect 2968 2952 3028 3206
rect 3480 3004 3486 3064
rect 3546 3004 3552 3064
rect 2962 2892 2968 2952
rect 3028 2892 3034 2952
rect 2760 2844 3248 2850
rect 2760 2810 2772 2844
rect 3236 2810 3248 2844
rect 2760 2804 3248 2810
rect 2464 2658 2478 2760
rect 1494 2184 1504 2220
rect 724 2134 1212 2140
rect 724 2100 736 2134
rect 1200 2100 1212 2134
rect 724 2094 1212 2100
rect 930 2040 990 2094
rect 1444 2040 1504 2184
rect 2472 2184 2478 2658
rect 2512 2658 2524 2760
rect 3486 2760 3546 3004
rect 4000 2952 4060 3206
rect 4500 3172 4560 3296
rect 5522 3296 5532 3358
rect 5566 3766 5578 3872
rect 6532 3872 6592 4408
rect 7552 4408 7568 4464
rect 7602 4464 7608 4984
rect 8566 4984 8626 5118
rect 8868 5068 9356 5074
rect 8868 5034 8880 5068
rect 9344 5034 9356 5068
rect 8868 5028 9356 5034
rect 7602 4408 7612 4464
rect 6832 4358 7320 4364
rect 6832 4324 6844 4358
rect 7308 4324 7320 4358
rect 6832 4318 7320 4324
rect 7552 4236 7612 4408
rect 8566 4408 8586 4984
rect 8620 4408 8626 4984
rect 7850 4358 8338 4364
rect 7850 4324 7862 4358
rect 8326 4324 8338 4358
rect 7850 4318 8338 4324
rect 7546 4176 7552 4236
rect 7612 4176 7618 4236
rect 6832 3956 7320 3962
rect 6832 3922 6844 3956
rect 7308 3922 7320 3956
rect 6832 3916 7320 3922
rect 5566 3358 5572 3766
rect 5566 3296 5582 3358
rect 4796 3246 5284 3252
rect 4796 3212 4808 3246
rect 5272 3212 5284 3246
rect 4796 3206 5284 3212
rect 3994 2892 4000 2952
rect 4060 2892 4066 2952
rect 3778 2844 4266 2850
rect 3778 2810 3790 2844
rect 4254 2810 4266 2844
rect 3778 2804 4266 2810
rect 3486 2720 3496 2760
rect 2512 2184 2518 2658
rect 2472 2172 2518 2184
rect 3490 2184 3496 2720
rect 3530 2720 3546 2760
rect 4500 2760 4560 3112
rect 5522 3064 5582 3296
rect 6532 3296 6550 3872
rect 6584 3296 6592 3872
rect 7552 3872 7612 4176
rect 7850 3956 8338 3962
rect 7850 3922 7862 3956
rect 8326 3922 8338 3956
rect 7850 3916 8338 3922
rect 7552 3830 7568 3872
rect 5814 3246 6302 3252
rect 5814 3212 5826 3246
rect 6290 3212 6302 3246
rect 5814 3206 6302 3212
rect 6532 3172 6592 3296
rect 7562 3296 7568 3830
rect 7602 3830 7612 3872
rect 8566 3872 8626 4408
rect 9588 4984 9648 5222
rect 10610 5178 10670 5232
rect 9886 5068 10374 5074
rect 9886 5034 9898 5068
rect 10362 5034 10374 5068
rect 9886 5028 10374 5034
rect 9588 4408 9604 4984
rect 9638 4408 9648 4984
rect 8868 4358 9356 4364
rect 8868 4324 8880 4358
rect 9344 4324 9356 4358
rect 8868 4318 9356 4324
rect 9078 4116 9138 4318
rect 9072 4056 9078 4116
rect 9138 4056 9144 4116
rect 9078 3962 9138 4056
rect 8868 3956 9356 3962
rect 8868 3922 8880 3956
rect 9344 3922 9356 3956
rect 8868 3916 9356 3922
rect 7602 3296 7608 3830
rect 7562 3284 7608 3296
rect 8566 3296 8586 3872
rect 8620 3296 8626 3872
rect 9588 3872 9648 4408
rect 10610 4984 10670 5118
rect 11114 5074 11174 5232
rect 10904 5068 11392 5074
rect 10904 5034 10916 5068
rect 11380 5034 11392 5068
rect 10904 5028 11392 5034
rect 10610 4408 10622 4984
rect 10656 4408 10670 4984
rect 9886 4358 10374 4364
rect 9886 4324 9898 4358
rect 10362 4324 10374 4358
rect 9886 4318 10374 4324
rect 10104 4116 10164 4318
rect 10610 4172 10670 4408
rect 11626 4984 11686 5232
rect 11626 4408 11640 4984
rect 11674 4408 11686 4984
rect 10904 4358 11392 4364
rect 10904 4324 10916 4358
rect 11380 4324 11392 4358
rect 10904 4318 11392 4324
rect 11110 4172 11170 4318
rect 11626 4172 11686 4408
rect 11766 4236 11826 6416
rect 11880 5326 11886 5386
rect 11946 5326 11952 5386
rect 11886 4730 11946 5326
rect 11882 4670 11888 4730
rect 11948 4670 11954 4730
rect 11760 4176 11766 4236
rect 11826 4176 11832 4236
rect 10098 4056 10104 4116
rect 10164 4056 10170 4116
rect 10610 4112 11686 4172
rect 10104 3962 10164 4056
rect 9886 3956 10374 3962
rect 9886 3922 9898 3956
rect 10362 3922 10374 3956
rect 9886 3916 10374 3922
rect 9588 3816 9604 3872
rect 9598 3342 9604 3816
rect 6832 3246 7320 3252
rect 6832 3212 6844 3246
rect 7308 3212 7320 3246
rect 6832 3206 7320 3212
rect 7850 3246 8338 3252
rect 7850 3212 7862 3246
rect 8326 3212 8338 3246
rect 7850 3206 8338 3212
rect 5516 3004 5522 3064
rect 5582 3004 5588 3064
rect 4994 2892 5000 2952
rect 5060 2892 5066 2952
rect 6014 2892 6020 2952
rect 6080 2892 6086 2952
rect 5000 2850 5060 2892
rect 6020 2850 6080 2892
rect 4796 2844 5284 2850
rect 4796 2810 4808 2844
rect 5272 2810 5284 2844
rect 4796 2804 5284 2810
rect 5814 2844 6302 2850
rect 5814 2810 5826 2844
rect 6290 2810 6302 2844
rect 5814 2804 6302 2810
rect 4500 2722 4514 2760
rect 3530 2184 3536 2720
rect 3490 2172 3536 2184
rect 4508 2184 4514 2722
rect 4548 2722 4560 2760
rect 5526 2760 5572 2772
rect 4548 2184 4554 2722
rect 5526 2244 5532 2760
rect 4508 2172 4554 2184
rect 5524 2184 5532 2244
rect 5566 2244 5572 2760
rect 6532 2760 6592 3112
rect 7040 2952 7100 3206
rect 7550 3004 7556 3064
rect 7616 3004 7622 3064
rect 7034 2892 7040 2952
rect 7100 2892 7106 2952
rect 6832 2844 7320 2850
rect 6832 2810 6844 2844
rect 7308 2810 7320 2844
rect 6832 2804 7320 2810
rect 6532 2700 6550 2760
rect 5566 2184 5584 2244
rect 1742 2134 2230 2140
rect 1742 2100 1754 2134
rect 2218 2100 2230 2134
rect 1742 2094 2230 2100
rect 2760 2134 3248 2140
rect 2760 2100 2772 2134
rect 3236 2100 3248 2134
rect 2760 2094 3248 2100
rect 3778 2134 4266 2140
rect 3778 2100 3790 2134
rect 4254 2100 4266 2134
rect 3778 2094 4266 2100
rect 4796 2134 5284 2140
rect 4796 2100 4808 2134
rect 5272 2100 5284 2134
rect 4796 2094 5284 2100
rect 282 1930 288 1990
rect 348 1930 354 1990
rect 426 1980 1504 2040
rect 2958 1990 3018 2094
rect 3990 1990 4050 2094
rect 1444 1860 1504 1980
rect 2952 1930 2958 1990
rect 3018 1930 3024 1990
rect 3984 1930 3990 1990
rect 4050 1930 4056 1990
rect 5524 1860 5584 2184
rect 6544 2184 6550 2700
rect 6584 2700 6592 2760
rect 7556 2760 7616 3004
rect 8050 2952 8110 3206
rect 8050 2886 8110 2892
rect 8566 3172 8626 3296
rect 9592 3296 9604 3342
rect 9638 3816 9648 3872
rect 10610 3872 10670 4112
rect 11110 3962 11170 4112
rect 10904 3956 11392 3962
rect 10904 3922 10916 3956
rect 11380 3922 11392 3956
rect 10904 3916 11392 3922
rect 9638 3342 9644 3816
rect 9638 3296 9652 3342
rect 8868 3246 9356 3252
rect 8868 3212 8880 3246
rect 9344 3212 9356 3246
rect 8868 3206 9356 3212
rect 7850 2844 8338 2850
rect 7850 2810 7862 2844
rect 8326 2810 8338 2844
rect 7850 2804 8338 2810
rect 7556 2714 7568 2760
rect 6584 2184 6590 2700
rect 6544 2172 6590 2184
rect 7562 2184 7568 2714
rect 7602 2714 7616 2760
rect 8566 2760 8626 3112
rect 9592 3064 9652 3296
rect 10610 3296 10622 3872
rect 10656 3296 10670 3872
rect 9886 3246 10374 3252
rect 9886 3212 9898 3246
rect 10362 3212 10374 3246
rect 9886 3206 10374 3212
rect 10610 3172 10670 3296
rect 11626 3872 11686 4112
rect 11626 3296 11640 3872
rect 11674 3296 11686 3872
rect 10904 3246 11392 3252
rect 10904 3212 10916 3246
rect 11380 3212 11392 3246
rect 10904 3206 11392 3212
rect 10604 3112 10610 3172
rect 10670 3112 10676 3172
rect 9586 3004 9592 3064
rect 9652 3004 9658 3064
rect 10610 3060 10670 3112
rect 11118 3060 11178 3206
rect 11626 3060 11686 3296
rect 10610 3000 11686 3060
rect 10082 2952 10142 2958
rect 9058 2892 9064 2952
rect 9124 2892 9130 2952
rect 9064 2850 9124 2892
rect 10082 2850 10142 2892
rect 8868 2844 9356 2850
rect 8868 2810 8880 2844
rect 9344 2810 9356 2844
rect 8868 2804 9356 2810
rect 9886 2844 10374 2850
rect 9886 2810 9898 2844
rect 10362 2810 10374 2844
rect 9886 2804 10374 2810
rect 8566 2718 8586 2760
rect 7602 2184 7608 2714
rect 7562 2172 7608 2184
rect 8580 2184 8586 2718
rect 8620 2184 8626 2760
rect 9598 2760 9644 2772
rect 9598 2212 9604 2760
rect 8580 2172 8626 2184
rect 9584 2184 9604 2212
rect 9638 2184 9644 2760
rect 10610 2760 10670 3000
rect 11118 2850 11178 3000
rect 10904 2844 11392 2850
rect 10904 2810 10916 2844
rect 11380 2810 11392 2844
rect 10904 2804 11392 2810
rect 10610 2696 10622 2760
rect 5814 2134 6302 2140
rect 5814 2100 5826 2134
rect 6290 2100 6302 2134
rect 5814 2094 6302 2100
rect 6832 2134 7320 2140
rect 6832 2100 6844 2134
rect 7308 2100 7320 2134
rect 6832 2094 7320 2100
rect 7850 2134 8338 2140
rect 7850 2100 7862 2134
rect 8326 2100 8338 2134
rect 7850 2094 8338 2100
rect 8868 2134 9356 2140
rect 8868 2100 8880 2134
rect 9344 2100 9356 2134
rect 8868 2094 9356 2100
rect 7050 1990 7110 2094
rect 8046 1990 8106 2094
rect 7044 1930 7050 1990
rect 7110 1930 7116 1990
rect 8040 1930 8046 1990
rect 8106 1930 8112 1990
rect 9584 1860 9644 2184
rect 10616 2184 10622 2696
rect 10656 2696 10670 2760
rect 11626 2760 11686 3000
rect 11626 2718 11640 2760
rect 10656 2184 10662 2696
rect 10616 2172 10662 2184
rect 11634 2184 11640 2718
rect 11674 2718 11686 2760
rect 11674 2184 11680 2718
rect 11634 2172 11680 2184
rect 9886 2134 10374 2140
rect 9886 2100 9898 2134
rect 10362 2100 10374 2134
rect 9886 2094 10374 2100
rect 10904 2134 11392 2140
rect 10904 2100 10916 2134
rect 11380 2100 11392 2134
rect 10904 2094 11392 2100
rect 11766 1860 11826 4176
rect 11886 2952 11946 4670
rect 11880 2892 11886 2952
rect 11946 2892 11952 2952
rect -1272 414 -1266 1842
rect 5518 1800 5524 1860
rect 5584 1800 5590 1860
rect 9578 1800 9584 1860
rect 9644 1800 9650 1860
rect 11760 1800 11766 1860
rect 11826 1800 11832 1860
rect 1444 1794 1504 1800
rect 886 1394 11122 1454
rect 886 1218 946 1394
rect 1386 1308 1446 1394
rect 1182 1302 1670 1308
rect 1182 1268 1194 1302
rect 1658 1268 1670 1302
rect 1182 1262 1670 1268
rect 886 1184 900 1218
rect 894 642 900 1184
rect 934 1184 946 1218
rect 1908 1218 1968 1394
rect 2406 1308 2466 1394
rect 3440 1308 3500 1394
rect 4462 1308 4522 1394
rect 5452 1308 5512 1394
rect 2200 1302 2688 1308
rect 2200 1268 2212 1302
rect 2676 1268 2688 1302
rect 2200 1262 2688 1268
rect 3218 1302 3706 1308
rect 3218 1268 3230 1302
rect 3694 1268 3706 1302
rect 3218 1262 3706 1268
rect 4236 1302 4724 1308
rect 4236 1268 4248 1302
rect 4712 1268 4724 1302
rect 4236 1262 4724 1268
rect 5254 1302 5742 1308
rect 5254 1268 5266 1302
rect 5730 1268 5742 1302
rect 5254 1262 5742 1268
rect 934 642 940 1184
rect 1908 1174 1918 1218
rect 894 630 940 642
rect 1912 642 1918 1174
rect 1952 1174 1968 1218
rect 2930 1218 2976 1230
rect 1952 642 1958 1174
rect 2930 700 2936 1218
rect 1912 630 1958 642
rect 2922 642 2936 700
rect 2970 700 2976 1218
rect 3948 1218 3994 1230
rect 2970 642 2982 700
rect 3948 676 3954 1218
rect 1182 592 1670 598
rect 1182 558 1194 592
rect 1658 558 1670 592
rect 1182 552 1670 558
rect 2200 592 2688 598
rect 2200 558 2212 592
rect 2676 558 2688 592
rect 2200 552 2688 558
rect 2922 494 2982 642
rect 3940 642 3954 676
rect 3988 676 3994 1218
rect 4966 1218 5012 1230
rect 4966 688 4972 1218
rect 3988 642 4000 676
rect 3218 592 3706 598
rect 3218 558 3230 592
rect 3694 558 3706 592
rect 3218 552 3706 558
rect 2916 434 2922 494
rect 2982 434 2988 494
rect -1272 396 -810 414
rect -1272 362 -1114 396
rect -914 362 -810 396
rect -1272 360 -810 362
rect -1272 40 -1188 360
rect -1378 -76 -1188 40
rect -1154 358 -810 360
rect -1154 344 -872 358
rect -1154 164 -1132 344
rect -1052 232 -1046 292
rect -986 232 -980 292
rect -1080 190 -1034 202
rect -1080 164 -1074 190
rect -1154 104 -1074 164
rect -1154 -68 -1132 104
rect -1080 84 -1074 104
rect -1040 84 -1034 190
rect -992 190 -946 202
rect -992 172 -986 190
rect -998 166 -986 172
rect -952 172 -946 190
rect -952 166 -938 172
rect -1004 106 -998 166
rect -938 106 -932 166
rect -998 100 -986 106
rect -1080 72 -1034 84
rect -992 84 -986 100
rect -952 100 -938 106
rect -952 84 -946 100
rect -992 72 -946 84
rect -1052 -18 -1046 42
rect -986 -18 -980 42
rect -894 -68 -872 344
rect -1154 -76 -872 -68
rect -836 -68 -810 358
rect 2922 -60 2982 434
rect 3940 382 4000 642
rect 4960 642 4972 688
rect 5006 688 5012 1218
rect 5976 1218 6036 1394
rect 6486 1308 6546 1394
rect 7476 1308 7536 1394
rect 8508 1308 8568 1394
rect 9512 1308 9572 1394
rect 6272 1302 6760 1308
rect 6272 1268 6284 1302
rect 6748 1268 6760 1302
rect 6272 1262 6760 1268
rect 7290 1302 7778 1308
rect 7290 1268 7302 1302
rect 7766 1268 7778 1302
rect 7290 1262 7778 1268
rect 8308 1302 8796 1308
rect 8308 1268 8320 1302
rect 8784 1268 8796 1302
rect 8308 1262 8796 1268
rect 9326 1302 9814 1308
rect 9326 1268 9338 1302
rect 9802 1268 9814 1302
rect 9326 1262 9814 1268
rect 6486 1260 6546 1262
rect 8508 1260 8568 1262
rect 5976 1176 5990 1218
rect 5006 642 5020 688
rect 4236 592 4724 598
rect 4236 558 4248 592
rect 4712 558 4724 592
rect 4236 552 4724 558
rect 4960 494 5020 642
rect 5984 642 5990 1176
rect 6024 1176 6036 1218
rect 7002 1218 7048 1230
rect 6024 642 6030 1176
rect 7002 688 7008 1218
rect 5984 630 6030 642
rect 6996 642 7008 688
rect 7042 688 7048 1218
rect 8020 1218 8066 1230
rect 7042 642 7056 688
rect 8020 680 8026 1218
rect 5254 592 5742 598
rect 5254 558 5266 592
rect 5730 558 5742 592
rect 5254 552 5742 558
rect 6272 592 6760 598
rect 6272 558 6284 592
rect 6748 558 6760 592
rect 6272 552 6760 558
rect 6996 494 7056 642
rect 8014 642 8026 680
rect 8060 680 8066 1218
rect 9038 1218 9084 1230
rect 8060 642 8074 680
rect 9038 674 9044 1218
rect 7290 592 7778 598
rect 7290 558 7302 592
rect 7766 558 7778 592
rect 7290 552 7778 558
rect 4954 434 4960 494
rect 5020 434 5026 494
rect 6990 434 6996 494
rect 7056 434 7062 494
rect 3934 322 3940 382
rect 4000 322 4006 382
rect 4960 -60 5020 434
rect 6996 -60 7056 434
rect 8014 382 8074 642
rect 9032 642 9044 674
rect 9078 674 9084 1218
rect 10052 1218 10112 1394
rect 10532 1308 10592 1394
rect 10344 1302 10832 1308
rect 10344 1268 10356 1302
rect 10820 1268 10832 1302
rect 10344 1262 10832 1268
rect 10052 1150 10062 1218
rect 9078 642 9092 674
rect 8308 592 8796 598
rect 8308 558 8320 592
rect 8784 558 8796 592
rect 8308 552 8796 558
rect 9032 494 9092 642
rect 10056 642 10062 1150
rect 10096 1150 10112 1218
rect 11062 1218 11122 1394
rect 11062 1178 11080 1218
rect 10096 642 10102 1150
rect 10056 630 10102 642
rect 11074 642 11080 1178
rect 11114 1178 11122 1218
rect 11114 642 11120 1178
rect 11074 630 11120 642
rect 9326 592 9814 598
rect 9326 558 9338 592
rect 9802 558 9814 592
rect 9326 552 9814 558
rect 10344 592 10832 598
rect 10344 558 10356 592
rect 10820 558 10832 592
rect 10344 552 10832 558
rect 9026 434 9032 494
rect 9092 434 9098 494
rect 8008 322 8014 382
rect 8074 322 8080 382
rect 9032 -60 9092 434
rect 12020 382 12080 7310
rect 12232 6476 12292 14816
rect 12226 6416 12232 6476
rect 12292 6416 12298 6476
rect 12352 6348 12412 14818
rect 12492 12066 12552 14836
rect 12604 14698 12610 14758
rect 12670 14698 12676 14758
rect 12492 9974 12552 12006
rect 12492 8732 12552 9914
rect 12492 7496 12552 8672
rect 12610 8630 12670 14698
rect 12720 14016 12780 14852
rect 12714 13956 12720 14016
rect 12780 13956 12786 14016
rect 12838 11096 12898 14952
rect 13166 14150 13226 14962
rect 13160 14090 13166 14150
rect 13226 14090 13232 14150
rect 12956 12732 12962 12792
rect 13022 12732 13028 12792
rect 12836 11090 12898 11096
rect 12896 11030 12898 11090
rect 12836 11024 12898 11030
rect 12604 8570 12610 8630
rect 12670 8570 12676 8630
rect 12492 6970 12552 7436
rect 12486 6910 12492 6970
rect 12552 6910 12558 6970
rect 12346 6288 12352 6348
rect 12412 6288 12418 6348
rect 12492 5386 12552 6910
rect 12486 5326 12492 5386
rect 12552 5326 12558 5386
rect 12838 5028 12898 11024
rect 12962 10096 13022 12732
rect 13168 12396 13174 12456
rect 13234 12396 13240 12456
rect 13064 11136 13070 11196
rect 13130 11136 13136 11196
rect 12956 10036 12962 10096
rect 13022 10036 13028 10096
rect 13070 5178 13130 11136
rect 13174 9860 13234 12396
rect 13286 12066 13346 14954
rect 13392 14878 13452 14884
rect 13392 12334 13452 14818
rect 24198 14522 24204 14528
rect 13518 14468 24204 14522
rect 24264 14522 24270 14528
rect 29302 14522 29308 14528
rect 24264 14468 29308 14522
rect 29368 14522 29374 14528
rect 33368 14522 33428 14528
rect 29368 14468 33368 14522
rect 13518 14462 33368 14468
rect 33428 14462 33940 14522
rect 13518 14322 13578 14462
rect 14040 14412 14100 14462
rect 15050 14412 15110 14462
rect 13814 14406 14302 14412
rect 13814 14372 13826 14406
rect 14290 14372 14302 14406
rect 13814 14366 14302 14372
rect 14832 14406 15320 14412
rect 14832 14372 14844 14406
rect 15308 14372 15320 14406
rect 14832 14366 15320 14372
rect 15050 14360 15110 14366
rect 13518 13746 13532 14322
rect 13566 13746 13578 14322
rect 14544 14322 14590 14334
rect 14544 13780 14550 14322
rect 13518 13504 13578 13746
rect 14536 13746 14550 13780
rect 14584 13780 14590 14322
rect 15556 14322 15616 14462
rect 16080 14412 16140 14462
rect 17092 14412 17152 14462
rect 15850 14406 16338 14412
rect 15850 14372 15862 14406
rect 16326 14372 16338 14406
rect 15850 14366 16338 14372
rect 16868 14406 17356 14412
rect 16868 14372 16880 14406
rect 17344 14372 17356 14406
rect 16868 14366 17356 14372
rect 17092 14360 17152 14366
rect 14584 13746 14596 13780
rect 13814 13696 14302 13702
rect 13814 13662 13826 13696
rect 14290 13662 14302 13696
rect 13814 13656 14302 13662
rect 14030 13594 14090 13656
rect 13814 13588 14302 13594
rect 13814 13554 13826 13588
rect 14290 13554 14302 13588
rect 13814 13548 14302 13554
rect 14030 13542 14090 13548
rect 13518 12928 13532 13504
rect 13566 12928 13578 13504
rect 13518 12456 13578 12928
rect 14536 13504 14596 13746
rect 15556 13746 15568 14322
rect 15602 13746 15616 14322
rect 16580 14322 16626 14334
rect 16580 13792 16586 14322
rect 15036 13702 15096 13704
rect 14832 13696 15320 13702
rect 14832 13662 14844 13696
rect 15308 13662 15320 13696
rect 14832 13656 15320 13662
rect 15036 13594 15096 13656
rect 14832 13588 15320 13594
rect 14832 13554 14844 13588
rect 15308 13554 15320 13588
rect 14832 13548 15320 13554
rect 14536 12928 14550 13504
rect 14584 12928 14596 13504
rect 15556 13504 15616 13746
rect 16570 13746 16586 13792
rect 16620 13792 16626 14322
rect 17588 14322 17648 14462
rect 18104 14412 18164 14462
rect 19104 14412 19164 14462
rect 17886 14406 18374 14412
rect 17886 14372 17898 14406
rect 18362 14372 18374 14406
rect 17886 14366 18374 14372
rect 18904 14406 19392 14412
rect 18904 14372 18916 14406
rect 19380 14372 19392 14406
rect 18904 14366 19392 14372
rect 16620 13746 16630 13792
rect 16048 13702 16108 13710
rect 15850 13696 16338 13702
rect 15850 13662 15862 13696
rect 16326 13662 16338 13696
rect 15850 13656 16338 13662
rect 16048 13594 16108 13656
rect 15850 13588 16338 13594
rect 15850 13554 15862 13588
rect 16326 13554 16338 13588
rect 15850 13548 16338 13554
rect 15556 13446 15568 13504
rect 13814 12878 14302 12884
rect 13814 12844 13826 12878
rect 14290 12844 14302 12878
rect 13814 12838 14302 12844
rect 14536 12792 14596 12928
rect 15562 12928 15568 13446
rect 15602 13446 15616 13504
rect 16570 13504 16630 13746
rect 17588 13746 17604 14322
rect 17638 13746 17648 14322
rect 18616 14322 18662 14334
rect 18616 13786 18622 14322
rect 16868 13696 17356 13702
rect 16868 13662 16880 13696
rect 17344 13662 17356 13696
rect 16868 13656 17356 13662
rect 17070 13594 17130 13656
rect 16868 13588 17356 13594
rect 16868 13554 16880 13588
rect 17344 13554 17356 13588
rect 16868 13548 17356 13554
rect 17070 13542 17130 13548
rect 15602 12928 15608 13446
rect 15562 12916 15608 12928
rect 16570 12928 16586 13504
rect 16620 12928 16630 13504
rect 17588 13504 17648 13746
rect 18606 13746 18622 13786
rect 18656 13786 18662 14322
rect 19626 14322 19686 14462
rect 20138 14412 20198 14462
rect 21150 14412 21210 14462
rect 19922 14406 20410 14412
rect 19922 14372 19934 14406
rect 20398 14372 20410 14406
rect 19922 14366 20410 14372
rect 20940 14406 21428 14412
rect 20940 14372 20952 14406
rect 21416 14372 21428 14406
rect 20940 14366 21428 14372
rect 18656 13746 18666 13786
rect 17886 13696 18374 13702
rect 17886 13662 17898 13696
rect 18362 13662 18374 13696
rect 17886 13656 18374 13662
rect 18082 13594 18142 13656
rect 17886 13588 18374 13594
rect 17886 13554 17898 13588
rect 18362 13554 18374 13588
rect 17886 13548 18374 13554
rect 18082 13542 18142 13548
rect 17588 13442 17604 13504
rect 14832 12878 15320 12884
rect 14832 12844 14844 12878
rect 15308 12844 15320 12878
rect 14832 12838 15320 12844
rect 15850 12878 16338 12884
rect 15850 12844 15862 12878
rect 16326 12844 16338 12878
rect 15850 12838 16338 12844
rect 16570 12790 16630 12928
rect 17598 12928 17604 13442
rect 17638 13442 17648 13504
rect 18606 13504 18666 13746
rect 19626 13746 19640 14322
rect 19674 13746 19686 14322
rect 20652 14322 20698 14334
rect 20652 13786 20658 14322
rect 18904 13696 19392 13702
rect 18904 13662 18916 13696
rect 19380 13662 19392 13696
rect 18904 13656 19392 13662
rect 19112 13594 19172 13656
rect 18904 13588 19392 13594
rect 18904 13554 18916 13588
rect 19380 13554 19392 13588
rect 18904 13548 19392 13554
rect 19112 13542 19172 13548
rect 17638 12928 17644 13442
rect 17598 12916 17644 12928
rect 18606 12928 18622 13504
rect 18656 12928 18666 13504
rect 19626 13504 19686 13746
rect 20644 13746 20658 13786
rect 20692 13786 20698 14322
rect 21662 14322 21722 14462
rect 22174 14412 22234 14462
rect 23186 14412 23246 14462
rect 21958 14406 22446 14412
rect 21958 14372 21970 14406
rect 22434 14372 22446 14406
rect 21958 14366 22446 14372
rect 22976 14406 23464 14412
rect 22976 14372 22988 14406
rect 23452 14372 23464 14406
rect 22976 14366 23464 14372
rect 20692 13746 20704 13786
rect 20118 13702 20178 13704
rect 19922 13696 20410 13702
rect 19922 13662 19934 13696
rect 20398 13662 20410 13696
rect 19922 13656 20410 13662
rect 20118 13594 20178 13656
rect 19922 13588 20410 13594
rect 19922 13554 19934 13588
rect 20398 13554 20410 13588
rect 19922 13548 20410 13554
rect 19626 13462 19640 13504
rect 16868 12878 17356 12884
rect 16868 12844 16880 12878
rect 17344 12844 17356 12878
rect 16868 12838 17356 12844
rect 17886 12878 18374 12884
rect 17886 12844 17898 12878
rect 18362 12844 18374 12878
rect 17886 12838 18374 12844
rect 18606 12790 18666 12928
rect 19634 12928 19640 13462
rect 19674 13462 19686 13504
rect 20644 13504 20704 13746
rect 21662 13746 21676 14322
rect 21710 13746 21722 14322
rect 22688 14322 22734 14334
rect 22688 13792 22694 14322
rect 21140 13702 21200 13704
rect 20940 13696 21428 13702
rect 20940 13662 20952 13696
rect 21416 13662 21428 13696
rect 20940 13656 21428 13662
rect 21140 13594 21200 13656
rect 20940 13588 21428 13594
rect 20940 13554 20952 13588
rect 21416 13554 21428 13588
rect 20940 13548 21428 13554
rect 19674 12928 19680 13462
rect 19634 12916 19680 12928
rect 20644 12928 20658 13504
rect 20692 12928 20704 13504
rect 21662 13504 21722 13746
rect 22682 13746 22694 13792
rect 22728 13792 22734 14322
rect 23694 14322 23754 14462
rect 24208 14412 24268 14462
rect 25220 14412 25280 14462
rect 23994 14406 24482 14412
rect 23994 14372 24006 14406
rect 24470 14372 24482 14406
rect 23994 14366 24482 14372
rect 25012 14406 25500 14412
rect 25012 14372 25024 14406
rect 25488 14372 25500 14406
rect 25012 14366 25500 14372
rect 25220 14360 25280 14366
rect 22728 13746 22742 13792
rect 21958 13696 22446 13702
rect 21958 13662 21970 13696
rect 22434 13662 22446 13696
rect 21958 13656 22446 13662
rect 22164 13594 22224 13656
rect 21958 13588 22446 13594
rect 21958 13554 21970 13588
rect 22434 13554 22446 13588
rect 21958 13548 22446 13554
rect 22164 13542 22224 13548
rect 21662 13454 21676 13504
rect 18904 12878 19392 12884
rect 18904 12844 18916 12878
rect 19380 12844 19392 12878
rect 18904 12838 19392 12844
rect 19922 12878 20410 12884
rect 19922 12844 19934 12878
rect 20398 12844 20410 12878
rect 19922 12838 20410 12844
rect 20644 12790 20704 12928
rect 21670 12928 21676 13454
rect 21710 13454 21722 13504
rect 22682 13504 22742 13746
rect 23694 13746 23712 14322
rect 23746 13746 23754 14322
rect 24724 14322 24770 14334
rect 24724 13792 24730 14322
rect 23170 13702 23230 13704
rect 22976 13696 23464 13702
rect 22976 13662 22988 13696
rect 23452 13662 23464 13696
rect 22976 13656 23464 13662
rect 23170 13594 23230 13656
rect 22976 13588 23464 13594
rect 22976 13554 22988 13588
rect 23452 13554 23464 13588
rect 22976 13548 23464 13554
rect 21710 12928 21716 13454
rect 21670 12916 21716 12928
rect 22682 12928 22694 13504
rect 22728 12928 22742 13504
rect 23694 13504 23754 13746
rect 24716 13746 24730 13792
rect 24764 13792 24770 14322
rect 25732 14322 25792 14462
rect 26244 14412 26304 14462
rect 27262 14412 27322 14462
rect 26030 14406 26518 14412
rect 26030 14372 26042 14406
rect 26506 14372 26518 14406
rect 26030 14366 26518 14372
rect 27048 14406 27536 14412
rect 27048 14372 27060 14406
rect 27524 14372 27536 14406
rect 27048 14366 27536 14372
rect 26244 14360 26304 14366
rect 24764 13746 24776 13792
rect 24194 13702 24254 13710
rect 23994 13696 24482 13702
rect 23994 13662 24006 13696
rect 24470 13662 24482 13696
rect 23994 13656 24482 13662
rect 24194 13594 24254 13656
rect 23994 13588 24482 13594
rect 23994 13554 24006 13588
rect 24470 13554 24482 13588
rect 23994 13548 24482 13554
rect 23694 13456 23712 13504
rect 20940 12878 21428 12884
rect 20940 12844 20952 12878
rect 21416 12844 21428 12878
rect 20940 12838 21428 12844
rect 21958 12878 22446 12884
rect 21958 12844 21970 12878
rect 22434 12844 22446 12878
rect 21958 12838 22446 12844
rect 22682 12790 22742 12928
rect 23706 12928 23712 13456
rect 23746 13456 23754 13504
rect 24716 13504 24776 13746
rect 25732 13746 25748 14322
rect 25782 13746 25792 14322
rect 26760 14322 26806 14334
rect 26760 13792 26766 14322
rect 25216 13702 25276 13704
rect 25012 13696 25500 13702
rect 25012 13662 25024 13696
rect 25488 13662 25500 13696
rect 25012 13656 25500 13662
rect 25216 13594 25276 13656
rect 25012 13588 25500 13594
rect 25012 13554 25024 13588
rect 25488 13554 25500 13588
rect 25012 13548 25500 13554
rect 23746 12928 23752 13456
rect 23706 12916 23752 12928
rect 24716 12928 24730 13504
rect 24764 12928 24776 13504
rect 25732 13504 25792 13746
rect 26752 13746 26766 13792
rect 26800 13792 26806 14322
rect 27768 14322 27828 14462
rect 28284 14412 28344 14462
rect 29308 14412 29368 14462
rect 28066 14406 28554 14412
rect 28066 14372 28078 14406
rect 28542 14372 28554 14406
rect 28066 14366 28554 14372
rect 29084 14406 29572 14412
rect 29084 14372 29096 14406
rect 29560 14372 29572 14406
rect 29084 14366 29572 14372
rect 26800 13746 26812 13792
rect 26228 13702 26288 13704
rect 26030 13696 26518 13702
rect 26030 13662 26042 13696
rect 26506 13662 26518 13696
rect 26030 13656 26518 13662
rect 26228 13594 26288 13656
rect 26030 13588 26518 13594
rect 26030 13554 26042 13588
rect 26506 13554 26518 13588
rect 26030 13548 26518 13554
rect 25732 13454 25748 13504
rect 22976 12878 23464 12884
rect 22976 12844 22988 12878
rect 23452 12844 23464 12878
rect 22976 12838 23464 12844
rect 23994 12878 24482 12884
rect 23994 12844 24006 12878
rect 24470 12844 24482 12878
rect 23994 12838 24482 12844
rect 24716 12790 24776 12928
rect 25742 12928 25748 13454
rect 25782 13454 25792 13504
rect 26752 13504 26812 13746
rect 27768 13746 27784 14322
rect 27818 13746 27828 14322
rect 28796 14322 28842 14334
rect 28796 13816 28802 14322
rect 27048 13696 27536 13702
rect 27048 13662 27060 13696
rect 27524 13662 27536 13696
rect 27048 13656 27536 13662
rect 27240 13594 27300 13656
rect 27048 13588 27536 13594
rect 27048 13554 27060 13588
rect 27524 13554 27536 13588
rect 27048 13548 27536 13554
rect 27240 13542 27300 13548
rect 25782 12928 25788 13454
rect 25742 12916 25788 12928
rect 26752 12928 26766 13504
rect 26800 12928 26812 13504
rect 27768 13504 27828 13746
rect 28790 13746 28802 13816
rect 28836 13816 28842 14322
rect 29804 14322 29864 14462
rect 30326 14412 30386 14462
rect 31338 14412 31398 14462
rect 30102 14406 30590 14412
rect 30102 14372 30114 14406
rect 30578 14372 30590 14406
rect 30102 14366 30590 14372
rect 31120 14406 31608 14412
rect 31120 14372 31132 14406
rect 31596 14372 31608 14406
rect 31120 14366 31608 14372
rect 28836 13746 28850 13816
rect 28264 13702 28324 13710
rect 28066 13696 28554 13702
rect 28066 13662 28078 13696
rect 28542 13662 28554 13696
rect 28066 13656 28554 13662
rect 28264 13594 28324 13656
rect 28066 13588 28554 13594
rect 28066 13554 28078 13588
rect 28542 13554 28554 13588
rect 28066 13548 28554 13554
rect 27768 13480 27784 13504
rect 25012 12878 25500 12884
rect 25012 12844 25024 12878
rect 25488 12844 25500 12878
rect 25012 12838 25500 12844
rect 26030 12878 26518 12884
rect 26030 12844 26042 12878
rect 26506 12844 26518 12878
rect 26030 12838 26518 12844
rect 26752 12790 26812 12928
rect 27778 12928 27784 13480
rect 27818 13480 27828 13504
rect 28790 13504 28850 13746
rect 29804 13746 29820 14322
rect 29854 13746 29864 14322
rect 30832 14322 30878 14334
rect 30832 13856 30838 14322
rect 29084 13696 29572 13702
rect 29084 13662 29096 13696
rect 29560 13662 29572 13696
rect 29084 13656 29572 13662
rect 29286 13594 29346 13656
rect 29084 13588 29572 13594
rect 29084 13554 29096 13588
rect 29560 13554 29572 13588
rect 29084 13548 29572 13554
rect 29286 13536 29346 13548
rect 27818 12928 27824 13480
rect 27778 12916 27824 12928
rect 28790 12928 28802 13504
rect 28836 12928 28850 13504
rect 29804 13504 29864 13746
rect 30824 13746 30838 13856
rect 30872 13856 30878 14322
rect 31842 14322 31902 14462
rect 32348 14412 32408 14462
rect 33366 14456 33428 14462
rect 33366 14412 33426 14456
rect 32138 14406 32626 14412
rect 32138 14372 32150 14406
rect 32614 14372 32626 14406
rect 32138 14366 32626 14372
rect 33156 14406 33644 14412
rect 33156 14372 33168 14406
rect 33632 14372 33644 14406
rect 33156 14366 33644 14372
rect 30872 13746 30884 13856
rect 30304 13702 30364 13704
rect 30102 13696 30590 13702
rect 30102 13662 30114 13696
rect 30578 13662 30590 13696
rect 30102 13656 30590 13662
rect 30304 13594 30364 13656
rect 30102 13588 30590 13594
rect 30102 13554 30114 13588
rect 30578 13554 30590 13588
rect 30102 13548 30590 13554
rect 29804 13462 29820 13504
rect 27048 12878 27536 12884
rect 27048 12844 27060 12878
rect 27524 12844 27536 12878
rect 27048 12838 27536 12844
rect 28066 12878 28554 12884
rect 28066 12844 28078 12878
rect 28542 12844 28554 12878
rect 28066 12838 28554 12844
rect 28790 12790 28850 12928
rect 29814 12928 29820 13462
rect 29854 13462 29864 13504
rect 30824 13504 30884 13746
rect 31842 13746 31856 14322
rect 31890 13746 31902 14322
rect 32868 14322 32914 14334
rect 32868 13806 32874 14322
rect 31334 13702 31394 13716
rect 31120 13696 31608 13702
rect 31120 13662 31132 13696
rect 31596 13662 31608 13696
rect 31120 13656 31608 13662
rect 31334 13594 31394 13656
rect 31120 13588 31608 13594
rect 31120 13554 31132 13588
rect 31596 13554 31608 13588
rect 31120 13548 31608 13554
rect 29854 12928 29860 13462
rect 29814 12916 29860 12928
rect 30824 12928 30838 13504
rect 30872 12928 30884 13504
rect 31842 13504 31902 13746
rect 32860 13746 32874 13806
rect 32908 13806 32914 14322
rect 33880 14322 33940 14462
rect 32908 13746 32920 13806
rect 32346 13702 32406 13716
rect 32138 13696 32626 13702
rect 32138 13662 32150 13696
rect 32614 13662 32626 13696
rect 32138 13656 32626 13662
rect 32346 13594 32406 13656
rect 32138 13588 32626 13594
rect 32138 13554 32150 13588
rect 32614 13554 32626 13588
rect 32138 13548 32626 13554
rect 31842 13462 31856 13504
rect 29084 12878 29572 12884
rect 29084 12844 29096 12878
rect 29560 12844 29572 12878
rect 29084 12838 29572 12844
rect 30102 12878 30590 12884
rect 30102 12844 30114 12878
rect 30578 12844 30590 12878
rect 30102 12838 30590 12844
rect 30824 12790 30884 12928
rect 31850 12928 31856 13462
rect 31890 13462 31902 13504
rect 32860 13504 32920 13746
rect 33880 13746 33892 14322
rect 33926 13746 33940 14322
rect 33156 13696 33644 13702
rect 33156 13662 33168 13696
rect 33632 13662 33644 13696
rect 33156 13656 33644 13662
rect 33346 13594 33406 13656
rect 33880 13654 33940 13746
rect 35766 14300 35878 15086
rect 37958 15192 76878 15198
rect 37958 15092 39728 15192
rect 76772 15092 76878 15192
rect 37958 15086 76878 15092
rect 37958 15070 50308 15086
rect 33880 13594 34660 13654
rect 33156 13588 33644 13594
rect 33156 13554 33168 13588
rect 33632 13554 33644 13588
rect 33156 13548 33644 13554
rect 33346 13542 33406 13548
rect 31890 12928 31896 13462
rect 31850 12916 31896 12928
rect 32860 12928 32874 13504
rect 32908 12928 32920 13504
rect 33880 13504 33940 13594
rect 33880 13454 33892 13504
rect 31120 12878 31608 12884
rect 31120 12844 31132 12878
rect 31596 12844 31608 12878
rect 31120 12838 31608 12844
rect 32138 12878 32626 12884
rect 32138 12844 32150 12878
rect 32614 12844 32626 12878
rect 32138 12838 32626 12844
rect 32860 12790 32920 12928
rect 33886 12928 33892 13454
rect 33926 13454 33940 13504
rect 33926 12928 33932 13454
rect 33886 12916 33932 12928
rect 33156 12878 33644 12884
rect 33156 12844 33168 12878
rect 33632 12844 33644 12878
rect 33156 12838 33644 12844
rect 14596 12732 34538 12790
rect 14536 12730 34538 12732
rect 14536 12726 14596 12730
rect 15544 12516 15550 12576
rect 15610 12516 15616 12576
rect 17584 12516 17590 12576
rect 17650 12516 17656 12576
rect 19624 12516 19630 12576
rect 19690 12516 19696 12576
rect 21654 12516 21660 12576
rect 21720 12516 21726 12576
rect 23694 12516 23700 12576
rect 23760 12516 23766 12576
rect 25726 12516 25732 12576
rect 25792 12516 25798 12576
rect 27766 12516 27772 12576
rect 27832 12516 27838 12576
rect 29802 12516 29808 12576
rect 29868 12516 29874 12576
rect 31836 12516 31842 12576
rect 31902 12516 31908 12576
rect 13512 12396 13518 12456
rect 13578 12396 13584 12456
rect 15036 12390 15042 12450
rect 15102 12390 15108 12450
rect 13386 12274 13392 12334
rect 13452 12274 13458 12334
rect 13280 12006 13286 12066
rect 13346 12006 13352 12066
rect 13286 9974 13346 12006
rect 13392 10200 13452 12274
rect 15042 12216 15102 12390
rect 13814 12210 14302 12216
rect 13814 12176 13826 12210
rect 14290 12176 14302 12210
rect 13814 12170 14302 12176
rect 14832 12210 15320 12216
rect 14832 12176 14844 12210
rect 15308 12176 15320 12210
rect 14832 12170 15320 12176
rect 13526 12126 13572 12138
rect 14544 12126 14590 12138
rect 15550 12126 15610 12516
rect 16056 12450 16116 12456
rect 16056 12216 16116 12390
rect 17078 12450 17138 12456
rect 17078 12216 17138 12390
rect 15850 12210 16338 12216
rect 15850 12176 15862 12210
rect 16326 12176 16338 12210
rect 15850 12170 16338 12176
rect 16868 12210 17356 12216
rect 16868 12176 16880 12210
rect 17344 12176 17356 12210
rect 16868 12170 17356 12176
rect 16580 12126 16626 12138
rect 13518 12092 13532 12126
rect 13526 11600 13532 12092
rect 13518 11550 13532 11600
rect 13566 12092 13578 12126
rect 13566 11600 13572 12092
rect 14536 12078 14550 12126
rect 13566 11550 13578 11600
rect 14544 11586 14550 12078
rect 13518 11412 13578 11550
rect 14536 11550 14550 11586
rect 14584 12078 14596 12126
rect 14584 11586 14590 12078
rect 15550 12058 15568 12126
rect 15562 11614 15568 12058
rect 14584 11550 14596 11586
rect 13814 11500 14302 11506
rect 13814 11466 13826 11500
rect 14290 11466 14302 11500
rect 13814 11460 14302 11466
rect 14020 11412 14080 11460
rect 14536 11412 14596 11550
rect 15554 11550 15568 11614
rect 15602 12094 15614 12126
rect 15602 12058 15610 12094
rect 15602 11614 15608 12058
rect 15602 11550 15614 11614
rect 16580 11596 16586 12126
rect 16576 11578 16586 11596
rect 16574 11550 16586 11578
rect 16620 11596 16626 12126
rect 17590 12126 17650 12516
rect 18092 12450 18152 12456
rect 18090 12390 18092 12396
rect 19118 12450 19178 12456
rect 18090 12384 18152 12390
rect 19116 12390 19118 12396
rect 19116 12384 19178 12390
rect 18090 12216 18150 12384
rect 18600 12274 18606 12334
rect 18666 12274 18672 12334
rect 17886 12210 18374 12216
rect 17886 12176 17898 12210
rect 18362 12176 18374 12210
rect 17886 12170 18374 12176
rect 17590 12072 17604 12126
rect 17598 11622 17604 12072
rect 17594 11598 17604 11622
rect 16620 11550 16636 11596
rect 17592 11550 17604 11598
rect 17638 12072 17650 12126
rect 18606 12126 18666 12274
rect 19116 12216 19176 12384
rect 18904 12210 19392 12216
rect 18904 12176 18916 12210
rect 19380 12176 19392 12210
rect 18904 12170 19392 12176
rect 18606 12084 18622 12126
rect 17638 11622 17644 12072
rect 18616 11626 18622 12084
rect 17638 11550 17654 11622
rect 18606 11550 18622 11626
rect 18656 12084 18666 12126
rect 19630 12126 19690 12516
rect 20130 12450 20190 12456
rect 20130 12216 20190 12390
rect 21166 12450 21226 12456
rect 21166 12216 21226 12390
rect 19922 12210 20410 12216
rect 19922 12176 19934 12210
rect 20398 12176 20410 12210
rect 19922 12170 20410 12176
rect 20940 12210 21428 12216
rect 20940 12176 20952 12210
rect 21416 12176 21428 12210
rect 20940 12170 21428 12176
rect 20652 12126 20698 12138
rect 21660 12126 21720 12516
rect 22172 12450 22232 12456
rect 23180 12390 23186 12450
rect 23246 12390 23252 12450
rect 22172 12216 22232 12390
rect 23186 12216 23246 12390
rect 21958 12210 22446 12216
rect 21958 12176 21970 12210
rect 22434 12176 22446 12210
rect 21958 12170 22446 12176
rect 22976 12210 23464 12216
rect 22976 12176 22988 12210
rect 23452 12176 23464 12210
rect 22976 12170 23464 12176
rect 18656 11626 18662 12084
rect 19630 12052 19640 12126
rect 18656 11610 18666 11626
rect 18656 11550 18670 11610
rect 19634 11606 19640 12052
rect 19626 11550 19640 11606
rect 19674 12052 19690 12126
rect 20646 12076 20658 12126
rect 19674 11606 19680 12052
rect 20652 11614 20658 12076
rect 19674 11550 19686 11606
rect 20646 11586 20658 11614
rect 20644 11550 20658 11586
rect 20692 12076 20706 12126
rect 20692 11614 20698 12076
rect 21660 12058 21676 12126
rect 21670 11626 21676 12058
rect 20692 11550 20706 11614
rect 14832 11500 15320 11506
rect 14832 11466 14844 11500
rect 15308 11466 15320 11500
rect 14832 11460 15320 11466
rect 13518 11352 14596 11412
rect 14536 11196 14596 11352
rect 15046 11302 15106 11460
rect 15554 11412 15614 11550
rect 15850 11500 16338 11506
rect 15850 11466 15862 11500
rect 16326 11466 16338 11500
rect 15850 11460 16338 11466
rect 15548 11352 15554 11412
rect 15614 11352 15620 11412
rect 15040 11242 15046 11302
rect 15106 11242 15112 11302
rect 14530 11136 14536 11196
rect 14596 11136 14602 11196
rect 13516 11030 13522 11090
rect 13582 11030 13588 11090
rect 14014 11030 14020 11090
rect 14080 11030 14086 11090
rect 14526 11030 14532 11090
rect 14592 11030 14598 11090
rect 13522 10894 13582 11030
rect 14020 10984 14080 11030
rect 13814 10978 14302 10984
rect 13814 10944 13826 10978
rect 14290 10944 14302 10978
rect 13814 10938 14302 10944
rect 13522 10854 13532 10894
rect 13526 10318 13532 10854
rect 13566 10854 13582 10894
rect 14532 10894 14592 11030
rect 15046 10984 15106 11242
rect 14832 10978 15320 10984
rect 14832 10944 14844 10978
rect 15308 10944 15320 10978
rect 14832 10938 15320 10944
rect 13566 10318 13572 10854
rect 14532 10848 14550 10894
rect 13526 10306 13572 10318
rect 14544 10318 14550 10848
rect 14584 10848 14592 10894
rect 15554 10894 15614 11352
rect 16068 11302 16128 11460
rect 16062 11242 16068 11302
rect 16128 11242 16134 11302
rect 16068 10984 16128 11242
rect 16576 11196 16636 11550
rect 16868 11500 17356 11506
rect 16868 11466 16880 11500
rect 17344 11466 17356 11500
rect 16868 11460 17356 11466
rect 17082 11302 17142 11460
rect 17594 11412 17654 11550
rect 18616 11538 18662 11550
rect 17886 11500 18374 11506
rect 17886 11466 17898 11500
rect 18362 11466 18374 11500
rect 17886 11460 18374 11466
rect 18904 11500 19392 11506
rect 18904 11466 18916 11500
rect 19380 11466 19392 11500
rect 18904 11460 19392 11466
rect 17588 11352 17594 11412
rect 17654 11352 17660 11412
rect 17076 11242 17082 11302
rect 17142 11242 17148 11302
rect 16570 11136 16576 11196
rect 16636 11136 16642 11196
rect 17082 10984 17142 11242
rect 15850 10978 16338 10984
rect 15850 10944 15862 10978
rect 16326 10944 16338 10978
rect 15850 10938 16338 10944
rect 16868 10978 17356 10984
rect 16868 10944 16880 10978
rect 17344 10944 17356 10978
rect 16868 10938 17356 10944
rect 16580 10894 16626 10906
rect 17594 10894 17654 11352
rect 18096 11302 18156 11460
rect 19114 11302 19174 11460
rect 19626 11412 19686 11550
rect 19922 11500 20410 11506
rect 19922 11466 19934 11500
rect 20398 11466 20410 11500
rect 19922 11460 20410 11466
rect 19620 11352 19626 11412
rect 19686 11352 19692 11412
rect 18090 11242 18096 11302
rect 18156 11242 18162 11302
rect 19108 11242 19114 11302
rect 19174 11242 19180 11302
rect 18096 10984 18156 11242
rect 18600 11136 18606 11196
rect 18666 11136 18672 11196
rect 17886 10978 18374 10984
rect 17886 10944 17898 10978
rect 18362 10944 18374 10978
rect 17886 10938 18374 10944
rect 15554 10856 15568 10894
rect 14584 10318 14590 10848
rect 15562 10376 15568 10856
rect 14544 10306 14590 10318
rect 15548 10318 15568 10376
rect 15602 10856 15614 10894
rect 15602 10318 15608 10856
rect 16574 10842 16586 10894
rect 16580 10338 16586 10842
rect 13814 10268 14302 10274
rect 13814 10234 13826 10268
rect 14290 10234 14302 10268
rect 13814 10228 14302 10234
rect 14832 10268 15320 10274
rect 14832 10234 14844 10268
rect 15308 10234 15320 10268
rect 14832 10228 15320 10234
rect 13386 10140 13392 10200
rect 13452 10140 13458 10200
rect 15548 10096 15608 10318
rect 16570 10318 16586 10338
rect 16620 10842 16634 10894
rect 16620 10338 16626 10842
rect 17592 10830 17604 10894
rect 17598 10382 17604 10830
rect 16620 10318 16630 10338
rect 15850 10268 16338 10274
rect 15850 10234 15862 10268
rect 16326 10234 16338 10268
rect 15850 10228 16338 10234
rect 13510 10036 13516 10096
rect 13576 10036 13582 10096
rect 15030 10036 15036 10096
rect 15096 10036 15102 10096
rect 15542 10036 15548 10096
rect 15608 10036 15614 10096
rect 13280 9914 13286 9974
rect 13346 9914 13352 9974
rect 13168 9800 13174 9860
rect 13234 9800 13240 9860
rect 13286 8732 13346 9914
rect 13516 9660 13576 10036
rect 14016 9800 14022 9860
rect 14082 9800 14088 9860
rect 14022 9750 14082 9800
rect 15036 9750 15096 10036
rect 15548 9802 15554 9862
rect 15614 9802 15620 9862
rect 13812 9744 14300 9750
rect 13812 9710 13824 9744
rect 14288 9710 14300 9744
rect 13812 9704 14300 9710
rect 14830 9744 15318 9750
rect 14830 9710 14842 9744
rect 15306 9710 15318 9744
rect 14830 9704 15318 9710
rect 14542 9660 14588 9672
rect 15554 9660 15614 9802
rect 16052 9750 16112 10228
rect 16570 10200 16630 10318
rect 17584 10318 17604 10382
rect 17638 10860 17654 10894
rect 18606 10894 18666 11136
rect 19114 10984 19174 11242
rect 18904 10978 19392 10984
rect 18904 10944 18916 10978
rect 19380 10944 19392 10978
rect 18904 10938 19392 10944
rect 19626 10894 19686 11352
rect 20140 11302 20200 11460
rect 20646 11342 20706 11550
rect 21658 11550 21676 11626
rect 21710 12058 21720 12126
rect 22688 12126 22734 12138
rect 21710 11626 21716 12058
rect 21710 11550 21718 11626
rect 22688 11612 22694 12126
rect 22682 11610 22694 11612
rect 20940 11500 21428 11506
rect 20940 11466 20952 11500
rect 21416 11466 21428 11500
rect 20940 11460 21428 11466
rect 20134 11242 20140 11302
rect 20200 11242 20206 11302
rect 20646 11282 20872 11342
rect 21160 11302 21220 11460
rect 21658 11412 21718 11550
rect 22680 11550 22694 11610
rect 22728 11612 22734 12126
rect 23700 12126 23760 12516
rect 24202 12450 24262 12456
rect 24202 12216 24262 12390
rect 25210 12450 25270 12456
rect 25270 12390 25272 12396
rect 25210 12384 25272 12390
rect 25212 12216 25272 12384
rect 23994 12210 24482 12216
rect 23994 12176 24006 12210
rect 24470 12176 24482 12210
rect 23994 12170 24482 12176
rect 25012 12210 25500 12216
rect 25012 12176 25024 12210
rect 25488 12176 25500 12210
rect 25012 12170 25500 12176
rect 24724 12126 24770 12138
rect 25732 12126 25792 12516
rect 26226 12450 26286 12456
rect 27250 12450 27310 12456
rect 26286 12390 26288 12396
rect 26226 12384 26288 12390
rect 26228 12216 26288 12384
rect 27250 12216 27310 12390
rect 26030 12210 26518 12216
rect 26030 12176 26042 12210
rect 26506 12176 26518 12210
rect 26030 12170 26518 12176
rect 27048 12210 27536 12216
rect 27048 12176 27060 12210
rect 27524 12176 27536 12210
rect 27048 12170 27536 12176
rect 26760 12126 26806 12138
rect 27772 12126 27832 12516
rect 28272 12450 28332 12456
rect 29294 12450 29354 12456
rect 28272 12216 28332 12390
rect 29292 12390 29294 12396
rect 29292 12384 29354 12390
rect 28788 12274 28794 12334
rect 28854 12274 28860 12334
rect 28066 12210 28554 12216
rect 28066 12176 28078 12210
rect 28542 12176 28554 12210
rect 28066 12170 28554 12176
rect 23700 12058 23712 12126
rect 23706 11616 23712 12058
rect 22728 11550 22742 11612
rect 23694 11550 23712 11616
rect 23746 12058 23760 12126
rect 24714 12092 24730 12126
rect 23746 11616 23752 12058
rect 23746 11550 23754 11616
rect 24724 11598 24730 12092
rect 21958 11500 22446 11506
rect 21958 11466 21970 11500
rect 22434 11466 22446 11500
rect 21958 11460 22446 11466
rect 21652 11352 21658 11412
rect 21718 11352 21724 11412
rect 20140 10984 20200 11242
rect 20640 11136 20646 11196
rect 20706 11136 20712 11196
rect 19922 10978 20410 10984
rect 19922 10944 19934 10978
rect 20398 10944 20410 10978
rect 19922 10938 20410 10944
rect 20646 10894 20706 11136
rect 20812 11090 20872 11282
rect 21154 11242 21160 11302
rect 21220 11242 21226 11302
rect 20806 11030 20812 11090
rect 20872 11030 20878 11090
rect 21160 10984 21220 11242
rect 20940 10978 21428 10984
rect 20940 10944 20952 10978
rect 21416 10944 21428 10978
rect 20940 10938 21428 10944
rect 17638 10830 17652 10860
rect 18606 10850 18622 10894
rect 17638 10318 17644 10830
rect 16868 10268 17356 10274
rect 16868 10234 16880 10268
rect 17344 10234 17356 10268
rect 16868 10228 17356 10234
rect 16564 10140 16570 10200
rect 16630 10140 16636 10200
rect 16566 10036 16572 10096
rect 16632 10036 16638 10096
rect 15848 9744 16336 9750
rect 15848 9710 15860 9744
rect 16324 9710 16336 9744
rect 15848 9704 16336 9710
rect 13516 9604 13530 9660
rect 13524 9084 13530 9604
rect 13564 9604 13576 9660
rect 14536 9628 14548 9660
rect 13564 9084 13570 9604
rect 14542 9128 14548 9628
rect 13524 9072 13570 9084
rect 14536 9084 14548 9128
rect 14582 9628 14596 9660
rect 15554 9634 15566 9660
rect 14582 9128 14588 9628
rect 14582 9084 14596 9128
rect 13812 9034 14300 9040
rect 13812 9000 13824 9034
rect 14288 9000 14300 9034
rect 13812 8994 14300 9000
rect 14536 8932 14596 9084
rect 15560 9084 15566 9634
rect 15600 9634 15614 9660
rect 16572 9660 16632 10036
rect 17072 9750 17132 10228
rect 17584 10096 17644 10318
rect 18616 10318 18622 10850
rect 18656 10860 18668 10894
rect 18656 10850 18666 10860
rect 19626 10852 19640 10894
rect 18656 10318 18662 10850
rect 19634 10360 19640 10852
rect 19626 10318 19640 10360
rect 19674 10852 19686 10894
rect 19674 10360 19680 10852
rect 20642 10832 20658 10894
rect 19674 10318 19686 10360
rect 20652 10318 20658 10832
rect 20692 10854 20706 10894
rect 21658 10894 21718 11352
rect 22180 11302 22240 11460
rect 22174 11242 22180 11302
rect 22240 11242 22246 11302
rect 22180 10984 22240 11242
rect 22680 11196 22740 11550
rect 22976 11500 23464 11506
rect 22976 11466 22988 11500
rect 23452 11466 23464 11500
rect 22976 11460 23464 11466
rect 23182 11302 23242 11460
rect 23694 11412 23754 11550
rect 24716 11550 24730 11598
rect 24764 12092 24774 12126
rect 24764 11598 24770 12092
rect 25732 12072 25748 12126
rect 25742 11610 25748 12072
rect 24764 11550 24776 11598
rect 23994 11500 24482 11506
rect 23994 11466 24006 11500
rect 24470 11466 24482 11500
rect 23994 11460 24482 11466
rect 23688 11352 23694 11412
rect 23754 11352 23760 11412
rect 23176 11242 23182 11302
rect 23242 11242 23248 11302
rect 22674 11136 22680 11196
rect 22740 11136 22746 11196
rect 22674 11030 22680 11090
rect 22740 11030 22746 11090
rect 21958 10978 22446 10984
rect 21958 10944 21970 10978
rect 22434 10944 22446 10978
rect 21958 10938 22446 10944
rect 22680 10894 22740 11030
rect 23182 10984 23242 11242
rect 22976 10978 23464 10984
rect 22976 10944 22988 10978
rect 23452 10944 23464 10978
rect 22976 10938 23464 10944
rect 23694 10894 23754 11352
rect 24208 11302 24268 11460
rect 24202 11242 24208 11302
rect 24268 11242 24274 11302
rect 24208 10984 24268 11242
rect 24716 11196 24776 11550
rect 25730 11550 25748 11610
rect 25782 12072 25792 12126
rect 26752 12086 26766 12126
rect 25782 11610 25788 12072
rect 26760 11616 26766 12086
rect 25782 11550 25790 11610
rect 26756 11590 26766 11616
rect 25012 11500 25500 11506
rect 25012 11466 25024 11500
rect 25488 11466 25500 11500
rect 25012 11460 25500 11466
rect 25226 11302 25286 11460
rect 25730 11412 25790 11550
rect 26754 11550 26766 11590
rect 26800 12086 26812 12126
rect 26800 11616 26806 12086
rect 27772 12072 27784 12126
rect 26800 11550 26816 11616
rect 27778 11600 27784 12072
rect 27768 11550 27784 11600
rect 27818 12072 27832 12126
rect 28794 12126 28854 12274
rect 29292 12216 29352 12384
rect 29084 12210 29572 12216
rect 29084 12176 29096 12210
rect 29560 12176 29572 12210
rect 29084 12170 29572 12176
rect 27818 11600 27824 12072
rect 28794 12062 28802 12126
rect 28796 11606 28802 12062
rect 27818 11550 27828 11600
rect 28788 11550 28802 11606
rect 28836 12062 28854 12126
rect 29808 12126 29868 12516
rect 30312 12450 30372 12456
rect 31326 12450 31386 12456
rect 30372 12390 30374 12396
rect 30312 12384 30374 12390
rect 31386 12390 31388 12396
rect 31326 12384 31388 12390
rect 30314 12216 30374 12384
rect 31328 12216 31388 12384
rect 30102 12210 30590 12216
rect 30102 12176 30114 12210
rect 30578 12176 30590 12210
rect 30102 12170 30590 12176
rect 31120 12210 31608 12216
rect 31120 12176 31132 12210
rect 31596 12176 31608 12210
rect 31120 12170 31608 12176
rect 30832 12126 30878 12138
rect 31842 12126 31902 12516
rect 32350 12450 32410 12456
rect 32348 12390 32350 12396
rect 32348 12384 32410 12390
rect 32348 12216 32408 12384
rect 32860 12274 32866 12334
rect 32926 12274 32932 12334
rect 33992 12274 33998 12334
rect 34058 12274 34064 12334
rect 32138 12210 32626 12216
rect 32138 12176 32150 12210
rect 32614 12176 32626 12210
rect 32138 12170 32626 12176
rect 32866 12126 32926 12274
rect 33156 12210 33644 12216
rect 33156 12176 33168 12210
rect 33632 12176 33644 12210
rect 33156 12170 33644 12176
rect 29808 12066 29820 12126
rect 28836 11606 28842 12062
rect 28836 11604 28848 11606
rect 28836 11550 28850 11604
rect 29814 11586 29820 12066
rect 29806 11550 29820 11586
rect 29854 12066 29868 12126
rect 30824 12086 30838 12126
rect 29854 11586 29860 12066
rect 30832 11606 30838 12086
rect 29854 11550 29866 11586
rect 26030 11500 26518 11506
rect 26030 11466 26042 11500
rect 26506 11466 26518 11500
rect 26030 11460 26518 11466
rect 25724 11352 25730 11412
rect 25790 11352 25796 11412
rect 25220 11242 25226 11302
rect 25286 11242 25292 11302
rect 24710 11136 24716 11196
rect 24776 11136 24782 11196
rect 24712 11030 24718 11090
rect 24778 11030 24784 11090
rect 23994 10978 24482 10984
rect 23994 10944 24006 10978
rect 24470 10944 24482 10978
rect 23994 10938 24482 10944
rect 24718 10894 24778 11030
rect 25226 10984 25286 11242
rect 25012 10978 25500 10984
rect 25012 10944 25024 10978
rect 25488 10944 25500 10978
rect 25012 10938 25500 10944
rect 25730 10894 25790 11352
rect 26234 11302 26294 11460
rect 26754 11334 26814 11550
rect 27246 11506 27306 11508
rect 27048 11500 27536 11506
rect 27048 11466 27060 11500
rect 27524 11466 27536 11500
rect 27048 11460 27536 11466
rect 26228 11242 26234 11302
rect 26294 11242 26300 11302
rect 26598 11274 26814 11334
rect 27246 11302 27306 11460
rect 27768 11412 27828 11550
rect 28796 11538 28842 11550
rect 28278 11506 28338 11508
rect 28066 11500 28554 11506
rect 28066 11466 28078 11500
rect 28542 11466 28554 11500
rect 28066 11460 28554 11466
rect 29084 11500 29572 11506
rect 29084 11466 29096 11500
rect 29560 11466 29572 11500
rect 29084 11460 29572 11466
rect 27762 11352 27768 11412
rect 27828 11352 27834 11412
rect 26234 10984 26294 11242
rect 26598 11090 26658 11274
rect 27240 11242 27246 11302
rect 27306 11242 27312 11302
rect 26746 11136 26752 11196
rect 26812 11136 26818 11196
rect 26592 11030 26598 11090
rect 26658 11030 26664 11090
rect 26030 10978 26518 10984
rect 26030 10944 26042 10978
rect 26506 10944 26518 10978
rect 26030 10938 26518 10944
rect 20692 10832 20702 10854
rect 21658 10838 21676 10894
rect 20692 10318 20698 10832
rect 21670 10360 21676 10838
rect 18616 10306 18662 10318
rect 19634 10306 19680 10318
rect 20652 10306 20698 10318
rect 21662 10318 21676 10360
rect 21710 10838 21718 10894
rect 22678 10842 22694 10894
rect 21710 10360 21716 10838
rect 21710 10318 21722 10360
rect 17886 10268 18374 10274
rect 17886 10234 17898 10268
rect 18362 10234 18374 10268
rect 17886 10228 18374 10234
rect 18904 10268 19392 10274
rect 18904 10234 18916 10268
rect 19380 10234 19392 10268
rect 18904 10228 19392 10234
rect 19922 10268 20410 10274
rect 19922 10234 19934 10268
rect 20398 10234 20410 10268
rect 19922 10228 20410 10234
rect 20940 10268 21428 10274
rect 20940 10234 20952 10268
rect 21416 10234 21428 10268
rect 20940 10228 21428 10234
rect 17578 10036 17584 10096
rect 17644 10036 17650 10096
rect 17584 9802 17590 9862
rect 17650 9802 17656 9862
rect 16866 9744 17354 9750
rect 16866 9710 16878 9744
rect 17342 9710 17354 9744
rect 16866 9704 17354 9710
rect 15600 9084 15606 9634
rect 16572 9628 16584 9660
rect 16578 9124 16584 9628
rect 15560 9072 15606 9084
rect 16570 9084 16584 9124
rect 16618 9628 16632 9660
rect 17590 9660 17650 9802
rect 18084 9750 18144 10228
rect 18598 10036 18604 10096
rect 18664 10036 18670 10096
rect 17884 9744 18372 9750
rect 17884 9710 17896 9744
rect 18360 9710 18372 9744
rect 17884 9704 18372 9710
rect 17590 9630 17602 9660
rect 16618 9124 16624 9628
rect 16618 9084 16630 9124
rect 14830 9034 15318 9040
rect 14830 9000 14842 9034
rect 15306 9000 15318 9034
rect 14830 8994 15318 9000
rect 15848 9034 16336 9040
rect 15848 9000 15860 9034
rect 16324 9000 16336 9034
rect 15848 8994 16336 9000
rect 13392 8872 13398 8932
rect 13458 8872 13464 8932
rect 14530 8872 14536 8932
rect 14596 8872 14602 8932
rect 13280 8672 13286 8732
rect 13346 8672 13352 8732
rect 13174 8570 13180 8630
rect 13240 8570 13246 8630
rect 13064 5118 13070 5178
rect 13130 5118 13136 5178
rect 13180 5140 13240 8570
rect 13286 7496 13346 8672
rect 13280 7436 13286 7496
rect 13346 7436 13352 7496
rect 13286 6976 13346 7436
rect 13286 6970 13350 6976
rect 13286 6910 13290 6970
rect 13286 6904 13350 6910
rect 13286 5386 13346 6904
rect 13398 6158 13458 8872
rect 14528 8672 14534 8732
rect 14594 8672 14600 8732
rect 14534 8628 14594 8672
rect 13518 8568 14594 8628
rect 13518 8566 14082 8568
rect 13518 8426 13578 8566
rect 14022 8516 14082 8566
rect 13812 8510 14300 8516
rect 13812 8476 13824 8510
rect 14288 8476 14300 8510
rect 13812 8470 14300 8476
rect 13518 8394 13530 8426
rect 13524 7850 13530 8394
rect 13564 8394 13578 8426
rect 14534 8426 14594 8568
rect 15038 8516 15098 8994
rect 15546 8792 15552 8852
rect 15612 8792 15618 8852
rect 14830 8510 15318 8516
rect 14830 8476 14842 8510
rect 15306 8476 15318 8510
rect 14830 8470 15318 8476
rect 13564 7850 13570 8394
rect 14534 8390 14548 8426
rect 13524 7838 13570 7850
rect 14542 7850 14548 8390
rect 14582 8390 14594 8426
rect 15552 8426 15612 8792
rect 16066 8738 16126 8994
rect 16570 8956 16630 9084
rect 17596 9084 17602 9630
rect 17636 9630 17650 9660
rect 18604 9660 18664 10036
rect 19110 9750 19170 10228
rect 19620 10140 19626 10200
rect 19686 10140 19692 10200
rect 18902 9744 19390 9750
rect 18902 9710 18914 9744
rect 19378 9710 19390 9744
rect 18902 9704 19390 9710
rect 17636 9084 17642 9630
rect 18604 9616 18620 9660
rect 18614 9134 18620 9616
rect 17596 9072 17642 9084
rect 18606 9084 18620 9134
rect 18654 9616 18664 9660
rect 19626 9660 19686 10140
rect 21662 10096 21722 10318
rect 22688 10318 22694 10842
rect 22728 10850 22742 10894
rect 22728 10842 22738 10850
rect 23694 10846 23712 10894
rect 22728 10318 22734 10842
rect 23706 10366 23712 10846
rect 22688 10306 22734 10318
rect 23700 10318 23712 10366
rect 23746 10846 23754 10894
rect 24714 10854 24730 10894
rect 23746 10366 23752 10846
rect 23746 10318 23760 10366
rect 21958 10268 22446 10274
rect 21958 10234 21970 10268
rect 22434 10234 22446 10268
rect 21958 10228 22446 10234
rect 22976 10268 23464 10274
rect 22976 10234 22988 10268
rect 23452 10234 23464 10268
rect 22976 10228 23464 10234
rect 23700 10096 23760 10318
rect 24724 10318 24730 10854
rect 24764 10856 24780 10894
rect 24764 10854 24778 10856
rect 24764 10318 24770 10854
rect 25730 10848 25748 10894
rect 25742 10372 25748 10848
rect 25730 10318 25748 10372
rect 25782 10848 25790 10894
rect 26752 10894 26812 11136
rect 27246 10984 27306 11242
rect 27048 10978 27536 10984
rect 27048 10944 27060 10978
rect 27524 10944 27536 10978
rect 27048 10938 27536 10944
rect 27768 10894 27828 11352
rect 28278 11302 28338 11460
rect 29292 11302 29352 11460
rect 29806 11412 29866 11550
rect 30822 11550 30838 11606
rect 30872 12086 30884 12126
rect 30872 11606 30878 12086
rect 30872 11550 30882 11606
rect 30102 11500 30590 11506
rect 30102 11466 30114 11500
rect 30578 11466 30590 11500
rect 30102 11460 30590 11466
rect 29800 11352 29806 11412
rect 29866 11352 29872 11412
rect 28272 11242 28278 11302
rect 28338 11242 28344 11302
rect 29286 11242 29292 11302
rect 29352 11242 29358 11302
rect 28278 10984 28338 11242
rect 28786 11136 28792 11196
rect 28852 11136 28858 11196
rect 28066 10978 28554 10984
rect 28066 10944 28078 10978
rect 28542 10944 28554 10978
rect 28066 10938 28554 10944
rect 28792 10894 28852 11136
rect 29292 10984 29352 11242
rect 29084 10978 29572 10984
rect 29084 10944 29096 10978
rect 29560 10944 29572 10978
rect 29084 10938 29572 10944
rect 25782 10372 25788 10848
rect 26752 10842 26766 10894
rect 25782 10318 25790 10372
rect 26760 10318 26766 10842
rect 26800 10852 26816 10894
rect 26800 10842 26812 10852
rect 26800 10318 26806 10842
rect 24724 10306 24770 10318
rect 25742 10306 25788 10318
rect 26760 10306 26806 10318
rect 27768 10318 27784 10894
rect 27818 10318 27828 10894
rect 28788 10852 28802 10894
rect 28792 10832 28802 10852
rect 23994 10268 24482 10274
rect 23994 10234 24006 10268
rect 24470 10234 24482 10268
rect 23994 10228 24482 10234
rect 25012 10268 25500 10274
rect 25012 10234 25024 10268
rect 25488 10234 25500 10268
rect 25012 10228 25500 10234
rect 26030 10268 26518 10274
rect 26030 10234 26042 10268
rect 26506 10234 26518 10268
rect 26030 10228 26518 10234
rect 27048 10268 27536 10274
rect 27048 10234 27060 10268
rect 27524 10234 27536 10268
rect 27048 10228 27536 10234
rect 25726 10140 25732 10200
rect 25792 10140 25798 10200
rect 21656 10036 21662 10096
rect 21722 10036 21728 10096
rect 23694 10036 23700 10096
rect 23760 10036 23766 10096
rect 20640 9914 20646 9974
rect 20706 9914 20712 9974
rect 22674 9914 22680 9974
rect 22740 9914 22746 9974
rect 24704 9914 24710 9974
rect 24770 9914 24776 9974
rect 19920 9744 20408 9750
rect 19920 9710 19932 9744
rect 20396 9710 20408 9744
rect 19920 9704 20408 9710
rect 18654 9134 18660 9616
rect 19626 9598 19638 9660
rect 18654 9084 18666 9134
rect 19632 9120 19638 9598
rect 16866 9034 17354 9040
rect 16866 9000 16878 9034
rect 17342 9000 17354 9034
rect 16866 8994 17354 9000
rect 17884 9034 18372 9040
rect 17884 9000 17896 9034
rect 18360 9000 18372 9034
rect 17884 8994 18372 9000
rect 16564 8896 16570 8956
rect 16630 8896 16636 8956
rect 16060 8678 16066 8738
rect 16126 8678 16132 8738
rect 16066 8516 16126 8678
rect 15848 8510 16336 8516
rect 15848 8476 15860 8510
rect 16324 8476 16336 8510
rect 15848 8470 16336 8476
rect 14582 7850 14588 8390
rect 15552 8384 15566 8426
rect 15560 7908 15566 8384
rect 14542 7838 14588 7850
rect 15554 7850 15566 7908
rect 15600 8384 15612 8426
rect 16570 8426 16630 8896
rect 17068 8744 17128 8994
rect 17586 8792 17592 8852
rect 17652 8792 17658 8852
rect 17068 8738 17130 8744
rect 17068 8678 17070 8738
rect 17068 8672 17130 8678
rect 17068 8516 17128 8672
rect 16866 8510 17354 8516
rect 16866 8476 16878 8510
rect 17342 8476 17354 8510
rect 16866 8470 17354 8476
rect 15600 7908 15606 8384
rect 16570 8382 16584 8426
rect 15600 7850 15614 7908
rect 16578 7898 16584 8382
rect 13812 7800 14300 7806
rect 13812 7766 13824 7800
rect 14288 7766 14300 7800
rect 13812 7760 14300 7766
rect 14830 7800 15318 7806
rect 14830 7766 14842 7800
rect 15306 7766 15318 7800
rect 14830 7760 15318 7766
rect 14528 7640 14534 7700
rect 14594 7640 14600 7700
rect 13812 7278 14300 7284
rect 13812 7244 13824 7278
rect 14288 7244 14300 7278
rect 13812 7238 14300 7244
rect 13524 7194 13570 7206
rect 13524 6664 13530 7194
rect 13514 6618 13530 6664
rect 13564 6664 13570 7194
rect 14534 7194 14594 7640
rect 15040 7598 15100 7760
rect 15034 7538 15040 7598
rect 15100 7538 15106 7598
rect 15554 7396 15614 7850
rect 16572 7850 16584 7898
rect 16618 8382 16630 8426
rect 17592 8426 17652 8792
rect 18084 8744 18144 8994
rect 18606 8956 18666 9084
rect 19624 9084 19638 9120
rect 19672 9598 19686 9660
rect 20646 9660 20706 9914
rect 20938 9744 21426 9750
rect 20938 9710 20950 9744
rect 21414 9710 21426 9744
rect 20938 9704 21426 9710
rect 21956 9744 22444 9750
rect 21956 9710 21968 9744
rect 22432 9710 22444 9744
rect 21956 9704 22444 9710
rect 20646 9604 20656 9660
rect 19672 9120 19678 9598
rect 19672 9084 19684 9120
rect 18902 9034 19390 9040
rect 18902 9000 18914 9034
rect 19378 9000 19390 9034
rect 18902 8994 19390 9000
rect 18600 8896 18606 8956
rect 18666 8896 18672 8956
rect 18082 8738 18144 8744
rect 18142 8678 18144 8738
rect 18082 8672 18144 8678
rect 18084 8516 18144 8672
rect 17884 8510 18372 8516
rect 17884 8476 17896 8510
rect 18360 8476 18372 8510
rect 17884 8470 18372 8476
rect 17592 8384 17602 8426
rect 16618 7898 16624 8382
rect 16618 7850 16632 7898
rect 15848 7800 16336 7806
rect 15848 7766 15860 7800
rect 16324 7766 16336 7800
rect 15848 7760 16336 7766
rect 16572 7700 16632 7850
rect 17596 7850 17602 8384
rect 17636 8384 17652 8426
rect 18606 8426 18666 8896
rect 19102 8738 19162 8994
rect 19624 8852 19684 9084
rect 20650 9084 20656 9604
rect 20690 9604 20706 9660
rect 21668 9660 21714 9672
rect 20690 9084 20696 9604
rect 21668 9114 21674 9660
rect 20650 9072 20696 9084
rect 21658 9084 21674 9114
rect 21708 9114 21714 9660
rect 22680 9660 22740 9914
rect 22974 9744 23462 9750
rect 22974 9710 22986 9744
rect 23450 9710 23462 9744
rect 22974 9704 23462 9710
rect 23992 9744 24480 9750
rect 23992 9710 24004 9744
rect 24468 9710 24480 9744
rect 23992 9704 24480 9710
rect 22680 9610 22692 9660
rect 21708 9084 21718 9114
rect 19920 9034 20408 9040
rect 19920 9000 19932 9034
rect 20396 9000 20408 9034
rect 19920 8994 20408 9000
rect 20938 9034 21426 9040
rect 20938 9000 20950 9034
rect 21414 9000 21426 9034
rect 20938 8994 21426 9000
rect 19618 8792 19624 8852
rect 19684 8792 19690 8852
rect 20114 8796 20174 8994
rect 21156 8796 21216 8994
rect 21658 8852 21718 9084
rect 22686 9084 22692 9610
rect 22726 9610 22740 9660
rect 23704 9660 23750 9672
rect 22726 9084 22732 9610
rect 23704 9126 23710 9660
rect 22686 9072 22732 9084
rect 23698 9084 23710 9126
rect 23744 9126 23750 9660
rect 24710 9660 24770 9914
rect 25010 9744 25498 9750
rect 25010 9710 25022 9744
rect 25486 9710 25498 9744
rect 25010 9704 25498 9710
rect 24710 9616 24728 9660
rect 23744 9084 23758 9126
rect 21956 9034 22444 9040
rect 21956 9000 21968 9034
rect 22432 9000 22444 9034
rect 21956 8994 22444 9000
rect 22974 9034 23462 9040
rect 22974 9000 22986 9034
rect 23450 9000 23462 9034
rect 22974 8994 23462 9000
rect 19618 8680 19624 8740
rect 19684 8680 19690 8740
rect 20114 8736 21216 8796
rect 21652 8792 21658 8852
rect 21718 8792 21724 8852
rect 19102 8516 19162 8678
rect 18902 8510 19390 8516
rect 18902 8476 18914 8510
rect 19378 8476 19390 8510
rect 18902 8470 19390 8476
rect 17636 7850 17642 8384
rect 18606 8378 18620 8426
rect 18614 7900 18620 8378
rect 17596 7838 17642 7850
rect 18608 7850 18620 7900
rect 18654 8378 18666 8426
rect 19624 8426 19684 8680
rect 20114 8516 20174 8736
rect 20636 8570 20642 8630
rect 20702 8570 20708 8630
rect 19920 8510 20408 8516
rect 19920 8476 19932 8510
rect 20396 8476 20408 8510
rect 19920 8470 20408 8476
rect 18654 7900 18660 8378
rect 19624 8368 19638 8426
rect 18654 7850 18668 7900
rect 16866 7800 17354 7806
rect 16866 7766 16878 7800
rect 17342 7766 17354 7800
rect 16866 7760 17354 7766
rect 17884 7800 18372 7806
rect 17884 7766 17896 7800
rect 18360 7766 18372 7800
rect 17884 7760 18372 7766
rect 16566 7640 16572 7700
rect 16632 7640 16638 7700
rect 16564 7436 16570 7496
rect 16630 7436 16636 7496
rect 17078 7490 17138 7760
rect 18100 7490 18160 7760
rect 18608 7700 18668 7850
rect 19632 7850 19638 8368
rect 19672 8368 19684 8426
rect 20642 8426 20702 8570
rect 21156 8516 21216 8736
rect 21654 8680 21660 8740
rect 21720 8680 21726 8740
rect 20938 8510 21426 8516
rect 20938 8476 20950 8510
rect 21414 8476 21426 8510
rect 20938 8470 21426 8476
rect 20642 8380 20656 8426
rect 19672 7850 19678 8368
rect 19632 7838 19678 7850
rect 20650 7850 20656 8380
rect 20690 8380 20702 8426
rect 21660 8426 21720 8680
rect 22156 8516 22216 8994
rect 22670 8570 22676 8630
rect 22736 8570 22742 8630
rect 21956 8510 22444 8516
rect 21956 8476 21968 8510
rect 22432 8476 22444 8510
rect 21956 8470 22444 8476
rect 20690 7850 20696 8380
rect 21660 8358 21674 8426
rect 20650 7838 20696 7850
rect 21668 7850 21674 8358
rect 21708 8358 21720 8426
rect 22676 8426 22736 8570
rect 23190 8516 23250 8994
rect 23698 8852 23758 9084
rect 24722 9084 24728 9616
rect 24762 9616 24770 9660
rect 25732 9660 25792 10140
rect 26254 9750 26314 10228
rect 26744 10036 26750 10096
rect 26810 10036 26816 10096
rect 26028 9744 26516 9750
rect 26028 9710 26040 9744
rect 26504 9710 26516 9744
rect 26028 9704 26516 9710
rect 24762 9084 24768 9616
rect 25732 9608 25746 9660
rect 25740 9136 25746 9608
rect 24722 9072 24768 9084
rect 25732 9084 25746 9136
rect 25780 9608 25792 9660
rect 26750 9660 26810 10036
rect 27256 9750 27316 10228
rect 27768 10096 27828 10318
rect 28796 10318 28802 10832
rect 28836 10832 28852 10894
rect 29806 10894 29866 11352
rect 30310 11302 30370 11460
rect 30304 11242 30310 11302
rect 30370 11242 30376 11302
rect 30310 10984 30370 11242
rect 30822 11196 30882 11550
rect 31842 11550 31856 12126
rect 31890 12094 31904 12126
rect 32862 12098 32874 12126
rect 31890 11550 31902 12094
rect 32866 12062 32874 12098
rect 32868 11610 32874 12062
rect 31120 11500 31608 11506
rect 31120 11466 31132 11500
rect 31596 11466 31608 11500
rect 31120 11460 31608 11466
rect 31334 11302 31394 11460
rect 31842 11412 31902 11550
rect 32862 11550 32874 11610
rect 32908 12062 32926 12126
rect 33886 12126 33932 12138
rect 32908 11610 32914 12062
rect 32908 11550 32922 11610
rect 33886 11598 33892 12126
rect 32138 11500 32626 11506
rect 32138 11466 32150 11500
rect 32614 11466 32626 11500
rect 32138 11460 32626 11466
rect 31836 11352 31842 11412
rect 31902 11352 31908 11412
rect 31328 11242 31334 11302
rect 31394 11242 31400 11302
rect 30816 11136 30822 11196
rect 30882 11136 30888 11196
rect 30816 11032 30822 11092
rect 30882 11032 30888 11092
rect 30102 10978 30590 10984
rect 30102 10944 30114 10978
rect 30578 10944 30590 10978
rect 30102 10938 30590 10944
rect 30302 10926 30362 10938
rect 30822 10894 30882 11032
rect 31334 10984 31394 11242
rect 31120 10978 31608 10984
rect 31120 10944 31132 10978
rect 31596 10944 31608 10978
rect 31120 10938 31608 10944
rect 29806 10836 29820 10894
rect 28836 10318 28842 10832
rect 29814 10366 29820 10836
rect 28796 10306 28842 10318
rect 29804 10318 29820 10366
rect 29854 10836 29866 10894
rect 30820 10848 30838 10894
rect 29854 10366 29860 10836
rect 30822 10820 30838 10848
rect 30832 10372 30838 10820
rect 29854 10318 29864 10366
rect 28066 10268 28554 10274
rect 28066 10234 28078 10268
rect 28542 10234 28554 10268
rect 28066 10228 28554 10234
rect 29084 10268 29572 10274
rect 29084 10234 29096 10268
rect 29560 10234 29572 10268
rect 29084 10228 29572 10234
rect 27762 10036 27768 10096
rect 27828 10036 27834 10096
rect 28268 9750 28328 10228
rect 28782 10036 28788 10096
rect 28848 10036 28854 10096
rect 27046 9744 27534 9750
rect 27046 9710 27058 9744
rect 27522 9710 27534 9744
rect 27046 9704 27534 9710
rect 28064 9744 28552 9750
rect 28064 9710 28076 9744
rect 28540 9710 28552 9744
rect 28064 9704 28552 9710
rect 26750 9612 26764 9660
rect 25780 9136 25786 9608
rect 25780 9084 25792 9136
rect 26758 9116 26764 9612
rect 23992 9034 24480 9040
rect 23992 9000 24004 9034
rect 24468 9000 24480 9034
rect 23992 8994 24480 9000
rect 25010 9034 25498 9040
rect 25010 9000 25022 9034
rect 25486 9000 25498 9034
rect 25010 8994 25498 9000
rect 23692 8792 23698 8852
rect 23758 8792 23764 8852
rect 24212 8796 24272 8994
rect 25220 8796 25280 8994
rect 25732 8852 25792 9084
rect 26750 9084 26764 9116
rect 26798 9612 26810 9660
rect 27776 9660 27822 9672
rect 26798 9116 26804 9612
rect 27776 9120 27782 9660
rect 26798 9084 26810 9116
rect 26028 9034 26516 9040
rect 26028 9000 26040 9034
rect 26504 9000 26516 9034
rect 26028 8994 26516 9000
rect 23690 8680 23696 8740
rect 23756 8680 23762 8740
rect 24212 8736 25280 8796
rect 25726 8792 25732 8852
rect 25792 8792 25798 8852
rect 25922 8788 25928 8848
rect 25988 8788 25994 8848
rect 22974 8510 23462 8516
rect 22974 8476 22986 8510
rect 23450 8476 23462 8510
rect 22974 8470 23462 8476
rect 22676 8378 22692 8426
rect 21708 7850 21714 8358
rect 21668 7838 21714 7850
rect 22686 7850 22692 8378
rect 22726 8378 22736 8426
rect 23696 8426 23756 8680
rect 24212 8516 24272 8736
rect 24710 8570 24716 8630
rect 24776 8570 24782 8630
rect 23992 8510 24480 8516
rect 23992 8476 24004 8510
rect 24468 8476 24480 8510
rect 23992 8470 24480 8476
rect 22726 7850 22732 8378
rect 23696 8376 23710 8426
rect 22686 7838 22732 7850
rect 23704 7850 23710 8376
rect 23744 8376 23756 8426
rect 24716 8426 24776 8570
rect 25220 8516 25280 8736
rect 25726 8680 25732 8740
rect 25792 8680 25798 8740
rect 25010 8510 25498 8516
rect 25010 8476 25022 8510
rect 25486 8476 25498 8510
rect 25010 8470 25498 8476
rect 24716 8388 24728 8426
rect 23744 7850 23750 8376
rect 24722 7896 24728 8388
rect 23704 7838 23750 7850
rect 24716 7850 24728 7896
rect 24762 8388 24776 8426
rect 25732 8426 25792 8680
rect 25928 8630 25988 8788
rect 26222 8632 26282 8994
rect 26750 8956 26810 9084
rect 27766 9084 27782 9120
rect 27816 9120 27822 9660
rect 28788 9660 28848 10036
rect 29302 9750 29362 10228
rect 29804 10096 29864 10318
rect 30826 10318 30838 10372
rect 30872 10820 30882 10894
rect 31842 10894 31902 11352
rect 32354 11302 32414 11460
rect 32862 11402 32922 11550
rect 33878 11550 33892 11598
rect 33926 11598 33932 12126
rect 33926 11550 33938 11598
rect 33156 11500 33644 11506
rect 33156 11466 33168 11500
rect 33632 11466 33644 11500
rect 33156 11460 33644 11466
rect 33372 11402 33432 11460
rect 33878 11402 33938 11550
rect 33998 11402 34058 12274
rect 32862 11342 34058 11402
rect 32348 11242 32354 11302
rect 32414 11242 32420 11302
rect 32354 10984 32414 11242
rect 32856 11136 32862 11196
rect 32922 11136 32928 11196
rect 32862 11094 32922 11136
rect 32862 11034 33940 11094
rect 33998 11092 34058 11342
rect 32138 10978 32626 10984
rect 32138 10944 32150 10978
rect 32614 10944 32626 10978
rect 32138 10938 32626 10944
rect 31842 10868 31856 10894
rect 30872 10372 30878 10820
rect 31850 10376 31856 10868
rect 30872 10318 30886 10372
rect 30102 10268 30590 10274
rect 30102 10234 30114 10268
rect 30578 10234 30590 10268
rect 30102 10228 30590 10234
rect 30826 10200 30886 10318
rect 31840 10318 31856 10376
rect 31890 10868 31902 10894
rect 32862 10894 32922 11034
rect 33348 10984 33408 11034
rect 33156 10978 33644 10984
rect 33156 10944 33168 10978
rect 33632 10944 33644 10978
rect 33156 10938 33644 10944
rect 33880 10894 33940 11034
rect 33992 11032 33998 11092
rect 34058 11032 34064 11092
rect 31890 10376 31896 10868
rect 32862 10838 32874 10894
rect 31890 10318 31900 10376
rect 31120 10268 31608 10274
rect 31120 10234 31132 10268
rect 31596 10234 31608 10268
rect 31120 10228 31608 10234
rect 30820 10140 30826 10200
rect 30886 10140 30892 10200
rect 31840 10096 31900 10318
rect 32868 10318 32874 10838
rect 32908 10838 32922 10894
rect 33876 10858 33892 10894
rect 33880 10852 33892 10858
rect 32908 10318 32914 10838
rect 33886 10362 33892 10852
rect 32868 10306 32914 10318
rect 33882 10318 33892 10362
rect 33926 10852 33940 10894
rect 33926 10362 33932 10852
rect 33926 10318 33942 10362
rect 32138 10268 32626 10274
rect 32138 10234 32150 10268
rect 32614 10234 32626 10268
rect 32138 10228 32626 10234
rect 33156 10268 33644 10274
rect 33156 10234 33168 10268
rect 33632 10234 33644 10268
rect 33156 10228 33644 10234
rect 29798 10036 29804 10096
rect 29864 10036 29870 10096
rect 31834 10036 31840 10096
rect 31900 10036 31906 10096
rect 32330 9750 32390 10228
rect 33882 10192 33942 10318
rect 33882 10132 34172 10192
rect 33368 9826 33936 9886
rect 33368 9750 33428 9826
rect 29082 9744 29570 9750
rect 29082 9710 29094 9744
rect 29558 9710 29570 9744
rect 29082 9704 29570 9710
rect 30100 9744 30588 9750
rect 30100 9710 30112 9744
rect 30576 9710 30588 9744
rect 30100 9704 30588 9710
rect 31118 9744 31606 9750
rect 31118 9710 31130 9744
rect 31594 9710 31606 9744
rect 31118 9704 31606 9710
rect 32136 9744 32624 9750
rect 32136 9710 32148 9744
rect 32612 9710 32624 9744
rect 32136 9704 32624 9710
rect 33154 9744 33642 9750
rect 33154 9710 33166 9744
rect 33630 9710 33642 9744
rect 33154 9704 33642 9710
rect 28788 9602 28800 9660
rect 28794 9130 28800 9602
rect 27816 9084 27826 9120
rect 27046 9034 27534 9040
rect 27046 9000 27058 9034
rect 27522 9000 27534 9034
rect 27046 8994 27534 9000
rect 26744 8896 26750 8956
rect 26810 8896 26816 8956
rect 25922 8570 25928 8630
rect 25988 8570 25994 8630
rect 26216 8572 26222 8632
rect 26282 8572 26288 8632
rect 26222 8516 26282 8572
rect 26028 8510 26516 8516
rect 26028 8476 26040 8510
rect 26504 8476 26516 8510
rect 26028 8470 26516 8476
rect 24762 7896 24768 8388
rect 25732 8382 25746 8426
rect 24762 7850 24776 7896
rect 18902 7800 19390 7806
rect 18902 7766 18914 7800
rect 19378 7766 19390 7800
rect 18902 7760 19390 7766
rect 19920 7800 20408 7806
rect 19920 7766 19932 7800
rect 20396 7766 20408 7800
rect 19920 7760 20408 7766
rect 20938 7800 21426 7806
rect 20938 7766 20950 7800
rect 21414 7766 21426 7800
rect 20938 7760 21426 7766
rect 21956 7800 22444 7806
rect 21956 7766 21968 7800
rect 22432 7766 22444 7800
rect 21956 7760 22444 7766
rect 22974 7800 23462 7806
rect 22974 7766 22986 7800
rect 23450 7766 23462 7800
rect 22974 7760 23462 7766
rect 23992 7800 24480 7806
rect 23992 7766 24004 7800
rect 24468 7766 24480 7800
rect 23992 7760 24480 7766
rect 18602 7640 18608 7700
rect 18668 7640 18674 7700
rect 15548 7336 15554 7396
rect 15614 7336 15620 7396
rect 14830 7278 15318 7284
rect 14830 7244 14842 7278
rect 15306 7244 15318 7278
rect 14830 7238 15318 7244
rect 14534 7156 14548 7194
rect 13564 6618 13574 6664
rect 14542 6660 14548 7156
rect 13514 6456 13574 6618
rect 14532 6618 14548 6660
rect 14582 7156 14594 7194
rect 15554 7194 15614 7336
rect 15848 7278 16336 7284
rect 15848 7244 15860 7278
rect 16324 7244 16336 7278
rect 15848 7238 16336 7244
rect 14582 6660 14588 7156
rect 15554 7154 15566 7194
rect 14582 6618 14592 6660
rect 13812 6568 14300 6574
rect 13812 6534 13824 6568
rect 14288 6534 14300 6568
rect 13812 6528 14300 6534
rect 14026 6456 14086 6528
rect 14532 6456 14592 6618
rect 15560 6618 15566 7154
rect 15600 7154 15614 7194
rect 16570 7194 16630 7436
rect 17072 7430 17078 7490
rect 17138 7430 17144 7490
rect 18094 7430 18100 7490
rect 18160 7430 18166 7490
rect 17582 7336 17588 7396
rect 17648 7336 17654 7396
rect 16866 7278 17354 7284
rect 16866 7244 16878 7278
rect 17342 7244 17354 7278
rect 16866 7238 17354 7244
rect 15600 6618 15606 7154
rect 16570 7142 16584 7194
rect 15560 6606 15606 6618
rect 16578 6618 16584 7142
rect 16618 7142 16630 7194
rect 17588 7194 17648 7336
rect 18100 7284 18160 7430
rect 17884 7278 18372 7284
rect 17884 7244 17896 7278
rect 18360 7244 18372 7278
rect 17884 7238 18372 7244
rect 17588 7150 17602 7194
rect 16618 6618 16624 7142
rect 17596 6654 17602 7150
rect 16578 6606 16624 6618
rect 17588 6618 17602 6654
rect 17636 7150 17648 7194
rect 18608 7194 18668 7640
rect 19114 7490 19174 7760
rect 20132 7598 20192 7760
rect 21152 7710 21212 7760
rect 22152 7710 22212 7760
rect 23190 7710 23250 7760
rect 24218 7710 24278 7760
rect 20634 7640 20640 7700
rect 20700 7640 20706 7700
rect 21152 7650 24278 7710
rect 20126 7538 20132 7598
rect 20192 7538 20198 7598
rect 19108 7430 19114 7490
rect 19174 7430 19180 7490
rect 20126 7430 20132 7490
rect 20192 7430 20198 7490
rect 19114 7284 19174 7430
rect 19618 7336 19624 7396
rect 19684 7336 19690 7396
rect 18902 7278 19390 7284
rect 18902 7244 18914 7278
rect 19378 7244 19390 7278
rect 18902 7238 19390 7244
rect 17636 6654 17642 7150
rect 17636 6618 17648 6654
rect 14830 6568 15318 6574
rect 14830 6534 14842 6568
rect 15306 6534 15318 6568
rect 14830 6528 15318 6534
rect 15848 6568 16336 6574
rect 15848 6534 15860 6568
rect 16324 6534 16336 6568
rect 15848 6528 16336 6534
rect 16866 6568 17354 6574
rect 16866 6534 16878 6568
rect 17342 6534 17354 6568
rect 16866 6528 17354 6534
rect 15036 6472 15096 6528
rect 13514 6396 14592 6456
rect 15030 6412 15036 6472
rect 15096 6412 15102 6472
rect 15940 6412 15946 6472
rect 16006 6412 16012 6472
rect 15030 6196 15036 6256
rect 15096 6196 15102 6256
rect 15036 6190 15098 6196
rect 13398 6152 13460 6158
rect 13398 6092 13400 6152
rect 13398 6086 13460 6092
rect 13282 5326 13288 5386
rect 13348 5326 13354 5386
rect 12832 4968 12838 5028
rect 12898 4968 12904 5028
rect 13070 1442 13130 5118
rect 13174 5080 13180 5140
rect 13240 5080 13246 5140
rect 13180 2650 13240 5080
rect 13286 4730 13346 5326
rect 13280 4670 13286 4730
rect 13346 4670 13352 4730
rect 13286 2776 13346 4670
rect 13398 3908 13458 6086
rect 15038 6050 15098 6190
rect 15946 6050 16006 6412
rect 16074 6256 16134 6528
rect 16942 6412 16948 6472
rect 17008 6412 17014 6472
rect 16074 6190 16134 6196
rect 16948 6050 17008 6412
rect 17088 6256 17148 6528
rect 17588 6370 17648 6618
rect 18608 6618 18620 7194
rect 18654 6618 18668 7194
rect 19624 7194 19684 7336
rect 20132 7284 20192 7430
rect 19920 7278 20408 7284
rect 19920 7244 19932 7278
rect 20396 7244 20408 7278
rect 19920 7238 20408 7244
rect 19624 7158 19638 7194
rect 17884 6568 18372 6574
rect 17884 6534 17896 6568
rect 18360 6534 18372 6568
rect 17884 6528 18372 6534
rect 18100 6472 18160 6528
rect 18094 6412 18100 6472
rect 18160 6412 18166 6472
rect 17582 6310 17588 6370
rect 17648 6310 17654 6370
rect 17082 6196 17088 6256
rect 17148 6196 17154 6256
rect 18100 6050 18160 6412
rect 13812 6044 14300 6050
rect 13812 6010 13824 6044
rect 14288 6010 14300 6044
rect 13812 6004 14300 6010
rect 14830 6044 15318 6050
rect 14830 6010 14842 6044
rect 15306 6010 15318 6044
rect 14830 6004 15318 6010
rect 15848 6044 16336 6050
rect 15848 6010 15860 6044
rect 16324 6010 16336 6044
rect 15848 6004 16336 6010
rect 16866 6044 17354 6050
rect 16866 6010 16878 6044
rect 17342 6010 17354 6044
rect 16866 6004 17354 6010
rect 17884 6044 18372 6050
rect 17884 6010 17896 6044
rect 18360 6010 18372 6044
rect 17884 6004 18372 6010
rect 13524 5960 13570 5972
rect 13524 5422 13530 5960
rect 13518 5384 13530 5422
rect 13564 5422 13570 5960
rect 14542 5960 14588 5972
rect 14542 5422 14548 5960
rect 13564 5384 13578 5422
rect 13518 5254 13578 5384
rect 14536 5384 14548 5422
rect 14582 5422 14588 5960
rect 15560 5960 15606 5972
rect 15560 5434 15566 5960
rect 14582 5384 14596 5422
rect 13812 5334 14300 5340
rect 13812 5300 13824 5334
rect 14288 5300 14300 5334
rect 13812 5294 14300 5300
rect 14016 5254 14076 5294
rect 14536 5254 14596 5384
rect 15552 5384 15566 5434
rect 15600 5434 15606 5960
rect 16578 5960 16624 5972
rect 16578 5442 16584 5960
rect 15600 5384 15612 5434
rect 14830 5334 15318 5340
rect 14830 5300 14842 5334
rect 15306 5300 15318 5334
rect 14830 5294 15318 5300
rect 13518 5194 14596 5254
rect 14536 5140 14596 5194
rect 15028 5184 15034 5244
rect 15094 5184 15100 5244
rect 14530 5080 14536 5140
rect 14596 5080 14602 5140
rect 14526 4870 14532 4930
rect 14592 4870 14598 4930
rect 13812 4810 14300 4816
rect 13812 4776 13824 4810
rect 14288 4776 14300 4810
rect 13812 4770 14300 4776
rect 13524 4726 13570 4738
rect 13524 4184 13530 4726
rect 13514 4150 13530 4184
rect 13564 4184 13570 4726
rect 14532 4726 14592 4870
rect 15034 4816 15094 5184
rect 15552 5028 15612 5384
rect 16570 5384 16584 5442
rect 16618 5442 16624 5960
rect 17596 5960 17642 5972
rect 16618 5384 16630 5442
rect 17596 5430 17602 5960
rect 15848 5334 16336 5340
rect 15848 5300 15860 5334
rect 16324 5300 16336 5334
rect 15848 5294 16336 5300
rect 16042 5244 16102 5294
rect 16036 5184 16042 5244
rect 16102 5184 16108 5244
rect 15546 4968 15552 5028
rect 15612 4968 15618 5028
rect 16570 4930 16630 5384
rect 17590 5384 17602 5430
rect 17636 5430 17642 5960
rect 18608 5960 18668 6618
rect 19632 6618 19638 7158
rect 19672 7158 19684 7194
rect 20640 7194 20700 7640
rect 21146 7430 21152 7490
rect 21212 7430 21218 7490
rect 24218 7474 24278 7650
rect 24716 7584 24776 7850
rect 25740 7850 25746 8382
rect 25780 8382 25792 8426
rect 26750 8426 26810 8896
rect 27252 8638 27312 8994
rect 27766 8740 27826 9084
rect 28786 9084 28800 9130
rect 28834 9602 28848 9660
rect 29812 9660 29858 9672
rect 28834 9130 28840 9602
rect 29812 9140 29818 9660
rect 28834 9084 28846 9130
rect 28064 9034 28552 9040
rect 28064 9000 28076 9034
rect 28540 9000 28552 9034
rect 28064 8994 28552 9000
rect 27760 8680 27766 8740
rect 27826 8680 27832 8740
rect 27250 8632 27312 8638
rect 27310 8572 27312 8632
rect 27250 8566 27312 8572
rect 27762 8566 27768 8626
rect 27828 8566 27834 8626
rect 27252 8516 27312 8566
rect 27046 8510 27534 8516
rect 27046 8476 27058 8510
rect 27522 8476 27534 8510
rect 27046 8470 27534 8476
rect 26750 8382 26764 8426
rect 25780 7850 25786 8382
rect 25740 7838 25786 7850
rect 26758 7850 26764 8382
rect 26798 8382 26810 8426
rect 27768 8426 27828 8566
rect 28276 8516 28336 8994
rect 28786 8956 28846 9084
rect 29804 9084 29818 9140
rect 29852 9140 29858 9660
rect 30830 9660 30876 9672
rect 29852 9084 29864 9140
rect 30830 9128 30836 9660
rect 29082 9034 29570 9040
rect 29082 9000 29094 9034
rect 29558 9000 29570 9034
rect 29082 8994 29570 9000
rect 28780 8896 28786 8956
rect 28846 8896 28852 8956
rect 28064 8510 28552 8516
rect 28064 8476 28076 8510
rect 28540 8476 28552 8510
rect 28064 8470 28552 8476
rect 27768 8396 27782 8426
rect 26798 7850 26804 8382
rect 27776 7890 27782 8396
rect 26758 7838 26804 7850
rect 27768 7850 27782 7890
rect 27816 8396 27828 8426
rect 28786 8426 28846 8896
rect 29302 8516 29362 8994
rect 29804 8740 29864 9084
rect 30820 9084 30836 9128
rect 30870 9128 30876 9660
rect 31848 9660 31894 9672
rect 31848 9128 31854 9660
rect 30870 9084 30880 9128
rect 30100 9034 30588 9040
rect 30100 9000 30112 9034
rect 30576 9000 30588 9034
rect 30100 8994 30588 9000
rect 29798 8680 29804 8740
rect 29864 8680 29870 8740
rect 30310 8690 30370 8994
rect 30820 8848 30880 9084
rect 31844 9084 31854 9128
rect 31888 9128 31894 9660
rect 32866 9660 32912 9672
rect 32866 9134 32872 9660
rect 31888 9084 31904 9128
rect 31118 9034 31606 9040
rect 31118 9000 31130 9034
rect 31594 9000 31606 9034
rect 31118 8994 31606 9000
rect 31326 8850 31386 8994
rect 30814 8788 30820 8848
rect 30880 8788 30886 8848
rect 31324 8844 31386 8850
rect 31384 8784 31386 8844
rect 31324 8778 31386 8784
rect 31326 8690 31386 8778
rect 31844 8740 31904 9084
rect 32860 9084 32872 9134
rect 32906 9134 32912 9660
rect 33876 9660 33936 9826
rect 33978 9802 33984 9862
rect 34044 9802 34050 9862
rect 34112 9844 34172 10132
rect 33876 9632 33890 9660
rect 33884 9142 33890 9632
rect 32906 9084 32920 9134
rect 32136 9034 32624 9040
rect 32136 9000 32148 9034
rect 32612 9000 32624 9034
rect 32136 8994 32624 9000
rect 30310 8630 31386 8690
rect 31838 8680 31844 8740
rect 31904 8680 31910 8740
rect 29798 8566 29804 8626
rect 29864 8566 29870 8626
rect 29082 8510 29570 8516
rect 29082 8476 29094 8510
rect 29558 8476 29570 8510
rect 29082 8470 29570 8476
rect 27816 7890 27822 8396
rect 28786 8386 28800 8426
rect 27816 7850 27828 7890
rect 28794 7884 28800 8386
rect 25010 7800 25498 7806
rect 25010 7766 25022 7800
rect 25486 7766 25498 7800
rect 25010 7760 25498 7766
rect 26028 7800 26516 7806
rect 26028 7766 26040 7800
rect 26504 7766 26516 7800
rect 26028 7760 26516 7766
rect 27046 7800 27534 7806
rect 27046 7766 27058 7800
rect 27522 7766 27534 7800
rect 27046 7760 27534 7766
rect 25222 7712 25282 7760
rect 24710 7524 24716 7584
rect 24776 7524 24782 7584
rect 25222 7474 25282 7652
rect 21152 7284 21212 7430
rect 24218 7414 25282 7474
rect 26746 7326 26752 7386
rect 26812 7326 26818 7386
rect 20938 7278 21426 7284
rect 20938 7244 20950 7278
rect 21414 7244 21426 7278
rect 20938 7238 21426 7244
rect 21956 7278 22444 7284
rect 21956 7244 21968 7278
rect 22432 7244 22444 7278
rect 21956 7238 22444 7244
rect 22974 7278 23462 7284
rect 22974 7244 22986 7278
rect 23450 7244 23462 7278
rect 22974 7238 23462 7244
rect 23992 7278 24480 7284
rect 23992 7244 24004 7278
rect 24468 7244 24480 7278
rect 23992 7238 24480 7244
rect 25010 7278 25498 7284
rect 25010 7244 25022 7278
rect 25486 7244 25498 7278
rect 25010 7238 25498 7244
rect 26028 7278 26516 7284
rect 26028 7244 26040 7278
rect 26504 7244 26516 7278
rect 26028 7238 26516 7244
rect 19672 6618 19678 7158
rect 20640 7156 20656 7194
rect 19632 6606 19678 6618
rect 20650 6618 20656 7156
rect 20690 7156 20700 7194
rect 21668 7194 21714 7206
rect 20690 6618 20696 7156
rect 21668 6660 21674 7194
rect 20650 6606 20696 6618
rect 21660 6618 21674 6660
rect 21708 6660 21714 7194
rect 22686 7194 22732 7206
rect 21708 6618 21720 6660
rect 22686 6656 22692 7194
rect 18902 6568 19390 6574
rect 18902 6534 18914 6568
rect 19378 6534 19390 6568
rect 18902 6528 19390 6534
rect 19920 6568 20408 6574
rect 19920 6534 19932 6568
rect 20396 6534 20408 6568
rect 19920 6528 20408 6534
rect 20938 6568 21426 6574
rect 20938 6534 20950 6568
rect 21414 6534 21426 6568
rect 20938 6528 21426 6534
rect 19110 6472 19170 6528
rect 20116 6472 20176 6528
rect 21160 6472 21220 6528
rect 21660 6478 21720 6618
rect 22680 6618 22692 6656
rect 22726 6656 22732 7194
rect 23704 7194 23750 7206
rect 22726 6618 22740 6656
rect 23704 6650 23710 7194
rect 21956 6568 22444 6574
rect 21956 6534 21968 6568
rect 22432 6534 22444 6568
rect 21956 6528 22444 6534
rect 19104 6412 19110 6472
rect 19170 6412 19176 6472
rect 20110 6412 20116 6472
rect 20176 6412 20182 6472
rect 21154 6412 21160 6472
rect 21220 6412 21226 6472
rect 21654 6418 21660 6478
rect 21720 6418 21726 6478
rect 19110 6050 19170 6412
rect 20108 6196 20114 6256
rect 20174 6196 20180 6256
rect 21148 6196 21154 6256
rect 21214 6196 21220 6256
rect 20114 6050 20174 6196
rect 20632 6092 20638 6152
rect 20698 6092 20704 6152
rect 18902 6044 19390 6050
rect 18902 6010 18914 6044
rect 19378 6010 19390 6044
rect 18902 6004 19390 6010
rect 19920 6044 20408 6050
rect 19920 6010 19932 6044
rect 20396 6010 20408 6044
rect 19920 6004 20408 6010
rect 18608 5878 18620 5960
rect 18614 5430 18620 5878
rect 17636 5384 17650 5430
rect 16866 5334 17354 5340
rect 16866 5300 16878 5334
rect 17342 5300 17354 5334
rect 16866 5294 17354 5300
rect 17056 5244 17116 5294
rect 17050 5184 17056 5244
rect 17116 5184 17122 5244
rect 17590 5028 17650 5384
rect 18610 5384 18620 5430
rect 18654 5878 18668 5960
rect 19632 5960 19678 5972
rect 18654 5430 18660 5878
rect 18654 5384 18670 5430
rect 19632 5428 19638 5960
rect 17884 5334 18372 5340
rect 17884 5300 17896 5334
rect 18360 5300 18372 5334
rect 17884 5294 18372 5300
rect 18094 5244 18154 5294
rect 18088 5184 18094 5244
rect 18154 5184 18160 5244
rect 17584 4968 17590 5028
rect 17650 4968 17656 5028
rect 16564 4870 16570 4930
rect 16630 4870 16636 4930
rect 18094 4816 18154 5184
rect 18610 4930 18670 5384
rect 19628 5384 19638 5428
rect 19672 5428 19678 5960
rect 20638 5960 20698 6092
rect 21154 6050 21214 6196
rect 20938 6044 21426 6050
rect 20938 6010 20950 6044
rect 21414 6010 21426 6044
rect 20938 6004 21426 6010
rect 20638 5896 20656 5960
rect 19672 5384 19688 5428
rect 18902 5334 19390 5340
rect 18902 5300 18914 5334
rect 19378 5300 19390 5334
rect 18902 5294 19390 5300
rect 19112 5244 19172 5294
rect 19628 5250 19688 5384
rect 20650 5384 20656 5896
rect 20690 5896 20698 5960
rect 21660 5960 21720 6418
rect 22168 6256 22228 6528
rect 22162 6196 22168 6256
rect 22228 6196 22234 6256
rect 22168 6050 22228 6196
rect 22680 6152 22740 6618
rect 23696 6618 23710 6650
rect 23744 6650 23750 7194
rect 24722 7194 24768 7206
rect 24722 6652 24728 7194
rect 23744 6618 23756 6650
rect 22974 6568 23462 6574
rect 22974 6534 22986 6568
rect 23450 6534 23462 6568
rect 22974 6528 23462 6534
rect 23176 6256 23236 6528
rect 23696 6478 23756 6618
rect 24718 6618 24728 6652
rect 24762 6652 24768 7194
rect 25740 7194 25786 7206
rect 24762 6618 24778 6652
rect 25740 6650 25746 7194
rect 23992 6568 24480 6574
rect 23992 6534 24004 6568
rect 24468 6534 24480 6568
rect 23992 6528 24480 6534
rect 23690 6418 23696 6478
rect 23756 6418 23762 6478
rect 24220 6256 24280 6528
rect 23170 6196 23176 6256
rect 23236 6196 23242 6256
rect 24214 6196 24220 6256
rect 24280 6196 24286 6256
rect 22674 6092 22680 6152
rect 22740 6092 22746 6152
rect 21956 6044 22444 6050
rect 21956 6010 21968 6044
rect 22432 6010 22444 6044
rect 21956 6004 22444 6010
rect 21660 5924 21674 5960
rect 20690 5384 20696 5896
rect 21668 5442 21674 5924
rect 20650 5372 20696 5384
rect 21664 5384 21674 5442
rect 21708 5924 21720 5960
rect 22680 5960 22740 6092
rect 23176 6050 23236 6196
rect 24220 6050 24280 6196
rect 24718 6152 24778 6618
rect 25732 6618 25746 6650
rect 25780 6650 25786 7194
rect 26752 7194 26812 7326
rect 27046 7278 27534 7284
rect 27046 7244 27058 7278
rect 27522 7244 27534 7278
rect 27046 7238 27534 7244
rect 25780 6618 25792 6650
rect 25010 6568 25498 6574
rect 25010 6534 25022 6568
rect 25486 6534 25498 6568
rect 25010 6528 25498 6534
rect 25210 6256 25270 6528
rect 25732 6478 25792 6618
rect 26752 6618 26764 7194
rect 26798 6618 26812 7194
rect 27768 7194 27828 7850
rect 28788 7850 28800 7884
rect 28834 8386 28846 8426
rect 29804 8426 29864 8566
rect 30310 8516 30370 8630
rect 31326 8516 31386 8630
rect 31836 8566 31842 8626
rect 31902 8566 31908 8626
rect 30100 8510 30588 8516
rect 30100 8476 30112 8510
rect 30576 8476 30588 8510
rect 30100 8470 30588 8476
rect 31118 8510 31606 8516
rect 31118 8476 31130 8510
rect 31594 8476 31606 8510
rect 31118 8470 31606 8476
rect 28834 7884 28840 8386
rect 29804 8384 29818 8426
rect 28834 7850 28848 7884
rect 28064 7800 28552 7806
rect 28064 7766 28076 7800
rect 28540 7766 28552 7800
rect 28064 7760 28552 7766
rect 28264 7490 28324 7760
rect 28258 7430 28264 7490
rect 28324 7430 28330 7490
rect 28264 7284 28324 7430
rect 28064 7278 28552 7284
rect 28064 7244 28076 7278
rect 28540 7244 28552 7278
rect 28064 7238 28552 7244
rect 27768 7154 27782 7194
rect 27776 6650 27782 7154
rect 26028 6568 26516 6574
rect 26028 6534 26040 6568
rect 26504 6534 26516 6568
rect 26028 6528 26516 6534
rect 25726 6418 25732 6478
rect 25792 6418 25798 6478
rect 26228 6256 26288 6528
rect 25204 6196 25210 6256
rect 25270 6196 25276 6256
rect 26222 6196 26228 6256
rect 26288 6196 26294 6256
rect 24712 6092 24718 6152
rect 24778 6092 24784 6152
rect 22974 6044 23462 6050
rect 22974 6010 22986 6044
rect 23450 6010 23462 6044
rect 22974 6004 23462 6010
rect 23992 6044 24480 6050
rect 23992 6010 24004 6044
rect 24468 6010 24480 6044
rect 23992 6004 24480 6010
rect 21708 5442 21714 5924
rect 22680 5922 22692 5960
rect 21708 5384 21724 5442
rect 19920 5334 20408 5340
rect 19920 5300 19932 5334
rect 20396 5300 20408 5334
rect 19920 5294 20408 5300
rect 20938 5334 21426 5340
rect 20938 5300 20950 5334
rect 21414 5300 21426 5334
rect 20938 5294 21426 5300
rect 21664 5250 21724 5384
rect 22686 5384 22692 5922
rect 22726 5922 22740 5960
rect 23704 5960 23750 5972
rect 22726 5384 22732 5922
rect 23704 5434 23710 5960
rect 22686 5372 22732 5384
rect 23696 5384 23710 5434
rect 23744 5434 23750 5960
rect 24718 5960 24778 6092
rect 25210 6050 25270 6196
rect 26752 6152 26812 6618
rect 27770 6618 27782 6650
rect 27816 7154 27828 7194
rect 28788 7194 28848 7850
rect 29812 7850 29818 8384
rect 29852 8384 29864 8426
rect 30830 8426 30876 8438
rect 29852 7850 29858 8384
rect 30830 7908 30836 8426
rect 29812 7838 29858 7850
rect 30822 7850 30836 7908
rect 30870 7908 30876 8426
rect 31842 8426 31902 8566
rect 32344 8516 32404 8994
rect 32860 8956 32920 9084
rect 33878 9084 33890 9142
rect 33924 9632 33936 9660
rect 33924 9142 33930 9632
rect 33924 9084 33938 9142
rect 33154 9034 33642 9040
rect 33154 9000 33166 9034
rect 33630 9000 33642 9034
rect 33154 8994 33642 9000
rect 33878 8974 33938 9084
rect 32854 8896 32860 8956
rect 32920 8896 32926 8956
rect 33872 8914 33878 8974
rect 33938 8914 33944 8974
rect 32860 8678 32920 8896
rect 32860 8618 33934 8678
rect 33984 8626 34044 9802
rect 34106 9784 34112 9844
rect 34172 9784 34178 9844
rect 34478 8844 34538 12730
rect 34472 8784 34478 8844
rect 34538 8784 34544 8844
rect 34222 8680 34228 8740
rect 34288 8680 34294 8740
rect 32136 8510 32624 8516
rect 32136 8476 32148 8510
rect 32612 8476 32624 8510
rect 32136 8470 32624 8476
rect 31842 8384 31854 8426
rect 30870 7850 30882 7908
rect 29294 7806 29354 7808
rect 29082 7800 29570 7806
rect 29082 7766 29094 7800
rect 29558 7766 29570 7800
rect 29082 7760 29570 7766
rect 30100 7800 30588 7806
rect 30100 7766 30112 7800
rect 30576 7766 30588 7800
rect 30100 7760 30588 7766
rect 29294 7490 29354 7760
rect 30316 7712 30376 7760
rect 30310 7652 30316 7712
rect 30376 7652 30382 7712
rect 30448 7656 30454 7716
rect 30514 7656 30520 7716
rect 30454 7490 30514 7656
rect 30822 7490 30882 7850
rect 31848 7850 31854 8384
rect 31888 8384 31902 8426
rect 32860 8426 32920 8618
rect 33364 8516 33424 8618
rect 33154 8510 33642 8516
rect 33154 8476 33166 8510
rect 33630 8476 33642 8510
rect 33154 8470 33642 8476
rect 32860 8392 32872 8426
rect 31888 7850 31894 8384
rect 32866 7890 32872 8392
rect 31848 7838 31894 7850
rect 32860 7850 32872 7890
rect 32906 8392 32920 8426
rect 33874 8426 33934 8618
rect 33978 8566 33984 8626
rect 34044 8566 34050 8626
rect 33874 8402 33890 8426
rect 32906 7890 32912 8392
rect 32906 7850 32920 7890
rect 31118 7800 31606 7806
rect 31118 7766 31130 7800
rect 31594 7766 31606 7800
rect 31118 7760 31606 7766
rect 32136 7800 32624 7806
rect 32136 7766 32148 7800
rect 32612 7766 32624 7800
rect 32136 7760 32624 7766
rect 32342 7716 32402 7760
rect 31330 7656 31336 7716
rect 31396 7656 31402 7716
rect 32336 7656 32342 7716
rect 32402 7656 32408 7716
rect 32860 7712 32920 7850
rect 33884 7850 33890 8402
rect 33924 8402 33934 8426
rect 33924 7850 33930 8402
rect 33884 7838 33930 7850
rect 33154 7800 33642 7806
rect 33154 7766 33166 7800
rect 33630 7766 33642 7800
rect 33154 7760 33642 7766
rect 29288 7430 29294 7490
rect 29354 7430 29360 7490
rect 30448 7430 30454 7490
rect 30514 7430 30520 7490
rect 30816 7430 30822 7490
rect 30882 7430 30888 7490
rect 29294 7284 29354 7430
rect 30454 7284 30514 7430
rect 30822 7386 30882 7430
rect 30816 7326 30822 7386
rect 30882 7326 30888 7386
rect 31336 7284 31396 7656
rect 32854 7652 32860 7712
rect 32920 7652 32926 7712
rect 32854 7524 32860 7584
rect 32920 7524 32926 7584
rect 31832 7328 31838 7388
rect 31898 7328 31904 7388
rect 29082 7278 29570 7284
rect 29082 7244 29094 7278
rect 29558 7244 29570 7278
rect 29082 7238 29570 7244
rect 30100 7278 30588 7284
rect 30100 7244 30112 7278
rect 30576 7244 30588 7278
rect 30100 7238 30588 7244
rect 31118 7278 31606 7284
rect 31118 7244 31130 7278
rect 31594 7244 31606 7278
rect 31118 7238 31606 7244
rect 31336 7236 31396 7238
rect 27816 6650 27822 7154
rect 28788 7148 28800 7194
rect 28794 6662 28800 7148
rect 27816 6618 27830 6650
rect 27046 6568 27534 6574
rect 27046 6534 27058 6568
rect 27522 6534 27534 6568
rect 27046 6528 27534 6534
rect 27262 6256 27322 6528
rect 27770 6478 27830 6618
rect 28786 6618 28800 6662
rect 28834 7148 28848 7194
rect 29812 7194 29858 7206
rect 28834 6662 28840 7148
rect 28834 6618 28846 6662
rect 29812 6658 29818 7194
rect 28064 6568 28552 6574
rect 28064 6534 28076 6568
rect 28540 6534 28552 6568
rect 28064 6528 28552 6534
rect 27764 6418 27770 6478
rect 27830 6418 27836 6478
rect 27756 6310 27762 6370
rect 27822 6310 27828 6370
rect 27256 6196 27262 6256
rect 27322 6196 27328 6256
rect 26746 6092 26752 6152
rect 26812 6092 26818 6152
rect 27258 6088 27264 6148
rect 27324 6088 27330 6148
rect 27264 6050 27324 6088
rect 25010 6044 25498 6050
rect 25010 6010 25022 6044
rect 25486 6010 25498 6044
rect 25010 6004 25498 6010
rect 26028 6044 26516 6050
rect 26028 6010 26040 6044
rect 26504 6010 26516 6044
rect 26028 6004 26516 6010
rect 27046 6044 27534 6050
rect 27046 6010 27058 6044
rect 27522 6010 27534 6044
rect 27046 6004 27534 6010
rect 24718 5924 24728 5960
rect 23744 5384 23756 5434
rect 21956 5334 22444 5340
rect 21956 5300 21968 5334
rect 22432 5300 22444 5334
rect 21956 5294 22444 5300
rect 22974 5334 23462 5340
rect 22974 5300 22986 5334
rect 23450 5300 23462 5334
rect 22974 5294 23462 5300
rect 23696 5250 23756 5384
rect 24722 5384 24728 5924
rect 24762 5924 24778 5960
rect 25740 5960 25786 5972
rect 24762 5384 24768 5924
rect 25740 5446 25746 5960
rect 24722 5372 24768 5384
rect 25730 5384 25746 5446
rect 25780 5446 25786 5960
rect 26758 5960 26804 5972
rect 25780 5384 25790 5446
rect 26758 5426 26764 5960
rect 23992 5334 24480 5340
rect 23992 5300 24004 5334
rect 24468 5300 24480 5334
rect 23992 5294 24480 5300
rect 25010 5334 25498 5340
rect 25010 5300 25022 5334
rect 25486 5300 25498 5334
rect 25010 5294 25498 5300
rect 25730 5250 25790 5384
rect 26752 5384 26764 5426
rect 26798 5426 26804 5960
rect 27762 5960 27822 6310
rect 28286 6148 28346 6528
rect 28786 6154 28846 6618
rect 29806 6618 29818 6658
rect 29852 6658 29858 7194
rect 30830 7194 30876 7206
rect 30830 6662 30836 7194
rect 29852 6618 29866 6658
rect 29082 6568 29570 6574
rect 29082 6534 29094 6568
rect 29558 6534 29570 6568
rect 29082 6528 29570 6534
rect 28280 6088 28286 6148
rect 28346 6088 28352 6148
rect 28780 6094 28786 6154
rect 28846 6094 28852 6154
rect 28286 6050 28346 6088
rect 28064 6044 28552 6050
rect 28064 6010 28076 6044
rect 28540 6010 28552 6044
rect 28064 6004 28552 6010
rect 27762 5924 27782 5960
rect 26798 5384 26812 5426
rect 26028 5334 26516 5340
rect 26028 5300 26040 5334
rect 26504 5300 26516 5334
rect 26028 5294 26516 5300
rect 19106 5184 19112 5244
rect 19172 5184 19178 5244
rect 19622 5190 19628 5250
rect 19688 5190 19694 5250
rect 23690 5190 23696 5250
rect 23756 5190 23762 5250
rect 25724 5190 25730 5250
rect 25790 5190 25796 5250
rect 18604 4870 18610 4930
rect 18670 4870 18676 4930
rect 14830 4810 15318 4816
rect 14830 4776 14842 4810
rect 15306 4776 15318 4810
rect 14830 4770 15318 4776
rect 15848 4810 16336 4816
rect 15848 4776 15860 4810
rect 16324 4776 16336 4810
rect 15848 4770 16336 4776
rect 16866 4810 17354 4816
rect 16866 4776 16878 4810
rect 17342 4776 17354 4810
rect 16866 4770 17354 4776
rect 17884 4810 18372 4816
rect 17884 4776 17896 4810
rect 18360 4776 18372 4810
rect 17884 4770 18372 4776
rect 14532 4672 14548 4726
rect 13564 4150 13574 4184
rect 14542 4180 14548 4672
rect 13514 4018 13574 4150
rect 14538 4150 14548 4180
rect 14582 4672 14592 4726
rect 15560 4726 15606 4738
rect 14582 4180 14588 4672
rect 15560 4196 15566 4726
rect 14582 4150 14598 4180
rect 13812 4100 14300 4106
rect 13812 4066 13824 4100
rect 14288 4066 14300 4100
rect 13812 4060 14300 4066
rect 14034 4018 14094 4060
rect 14538 4018 14598 4150
rect 15552 4150 15566 4196
rect 15600 4196 15606 4726
rect 16578 4726 16624 4738
rect 15600 4150 15612 4196
rect 16578 4180 16584 4726
rect 14830 4100 15318 4106
rect 14830 4066 14842 4100
rect 15306 4066 15318 4100
rect 14830 4060 15318 4066
rect 13514 3958 14598 4018
rect 13392 3848 13398 3908
rect 13458 3848 13464 3908
rect 14538 3812 14598 3958
rect 13514 3752 14598 3812
rect 13514 3494 13574 3752
rect 14026 3584 14086 3752
rect 14538 3692 14598 3752
rect 14532 3632 14538 3692
rect 14598 3632 14604 3692
rect 13812 3578 14300 3584
rect 13812 3544 13824 3578
rect 14288 3544 14300 3578
rect 13812 3538 14300 3544
rect 13514 3458 13530 3494
rect 13524 2918 13530 3458
rect 13564 3458 13574 3494
rect 14538 3494 14598 3632
rect 15030 3584 15090 4060
rect 15552 4006 15612 4150
rect 16570 4150 16584 4180
rect 16618 4180 16624 4726
rect 17596 4726 17642 4738
rect 17596 4192 17602 4726
rect 16618 4150 16630 4180
rect 15848 4100 16336 4106
rect 15848 4066 15860 4100
rect 16324 4066 16336 4100
rect 15848 4060 16336 4066
rect 15546 3946 15552 4006
rect 15612 3946 15618 4006
rect 15550 3752 15556 3812
rect 15616 3752 15622 3812
rect 14830 3578 15318 3584
rect 14830 3544 14842 3578
rect 15306 3544 15318 3578
rect 14830 3538 15318 3544
rect 13564 2918 13570 3458
rect 14538 3454 14548 3494
rect 13524 2906 13570 2918
rect 14542 2918 14548 3454
rect 14582 3454 14598 3494
rect 15556 3494 15616 3752
rect 16050 3748 16110 4060
rect 16570 3908 16630 4150
rect 17588 4150 17602 4192
rect 17636 4192 17642 4726
rect 18610 4726 18670 4870
rect 19112 4816 19172 5184
rect 18902 4810 19390 4816
rect 18902 4776 18914 4810
rect 19378 4776 19390 4810
rect 18902 4770 19390 4776
rect 18610 4696 18620 4726
rect 18614 4214 18620 4696
rect 17636 4150 17648 4192
rect 16866 4100 17354 4106
rect 16866 4066 16878 4100
rect 17342 4066 17354 4100
rect 16866 4060 17354 4066
rect 16564 3848 16570 3908
rect 16630 3848 16636 3908
rect 17084 3748 17144 4060
rect 17588 4006 17648 4150
rect 18606 4150 18620 4214
rect 18654 4696 18670 4726
rect 19628 4726 19688 5190
rect 21664 5184 21724 5190
rect 22674 5080 22680 5140
rect 22740 5080 22746 5140
rect 24710 5080 24716 5140
rect 24776 5080 24782 5140
rect 21656 4968 21662 5028
rect 21722 4968 21728 5028
rect 20640 4870 20646 4930
rect 20706 4870 20712 4930
rect 19920 4810 20408 4816
rect 19920 4776 19932 4810
rect 20396 4776 20408 4810
rect 19920 4770 20408 4776
rect 18654 4214 18660 4696
rect 19628 4684 19638 4726
rect 18654 4150 18666 4214
rect 19632 4190 19638 4684
rect 17884 4100 18372 4106
rect 17884 4066 17896 4100
rect 18360 4066 18372 4100
rect 17884 4060 18372 4066
rect 17582 3946 17588 4006
rect 17648 3946 17654 4006
rect 18094 3908 18154 4060
rect 18088 3848 18094 3908
rect 18154 3848 18160 3908
rect 17586 3752 17592 3812
rect 17652 3752 17658 3812
rect 16050 3688 17144 3748
rect 16050 3584 16110 3688
rect 17084 3584 17144 3688
rect 15848 3578 16336 3584
rect 15848 3544 15860 3578
rect 16324 3544 16336 3578
rect 15848 3538 16336 3544
rect 16866 3578 17354 3584
rect 16866 3544 16878 3578
rect 17342 3544 17354 3578
rect 16866 3538 17354 3544
rect 14582 2918 14588 3454
rect 15556 3450 15566 3494
rect 14542 2906 14588 2918
rect 15560 2918 15566 3450
rect 15600 3450 15616 3494
rect 16578 3494 16624 3506
rect 15600 2918 15606 3450
rect 16578 2960 16584 3494
rect 15560 2906 15606 2918
rect 16570 2918 16584 2960
rect 16618 2960 16624 3494
rect 17592 3494 17652 3752
rect 18094 3584 18154 3848
rect 18606 3692 18666 4150
rect 19626 4150 19638 4190
rect 19672 4684 19688 4726
rect 20646 4726 20706 4870
rect 20938 4810 21426 4816
rect 20938 4776 20950 4810
rect 21414 4776 21426 4810
rect 20938 4770 21426 4776
rect 20646 4690 20656 4726
rect 19672 4190 19678 4684
rect 19672 4150 19686 4190
rect 20650 4184 20656 4690
rect 18902 4100 19390 4106
rect 18902 4066 18914 4100
rect 19378 4066 19390 4100
rect 18902 4060 19390 4066
rect 19116 3908 19176 4060
rect 19626 4006 19686 4150
rect 20640 4150 20656 4184
rect 20690 4690 20706 4726
rect 21662 4726 21722 4968
rect 21956 4810 22444 4816
rect 21956 4776 21968 4810
rect 22432 4776 22444 4810
rect 21956 4770 22444 4776
rect 21662 4700 21674 4726
rect 20690 4184 20696 4690
rect 21668 4206 21674 4700
rect 20690 4150 20700 4184
rect 19920 4100 20408 4106
rect 19920 4066 19932 4100
rect 20396 4066 20408 4100
rect 19920 4060 20408 4066
rect 19620 3946 19626 4006
rect 19686 3946 19692 4006
rect 20140 3914 20200 4060
rect 18600 3632 18606 3692
rect 18666 3632 18672 3692
rect 17884 3578 18372 3584
rect 17884 3544 17896 3578
rect 18360 3544 18372 3578
rect 17884 3538 18372 3544
rect 17592 3442 17602 3494
rect 16618 2918 16630 2960
rect 13812 2868 14300 2874
rect 13812 2834 13824 2868
rect 14288 2834 14300 2868
rect 13812 2828 14300 2834
rect 14830 2868 15318 2874
rect 14830 2834 14842 2868
rect 15306 2834 15318 2868
rect 14830 2828 15318 2834
rect 15848 2868 16336 2874
rect 15848 2834 15860 2868
rect 16324 2834 16336 2868
rect 15848 2828 16336 2834
rect 13280 2716 13286 2776
rect 13346 2716 13352 2776
rect 13174 2590 13180 2650
rect 13240 2590 13246 2650
rect 13514 2410 14594 2470
rect 13514 2260 13574 2410
rect 14022 2350 14082 2410
rect 13812 2344 14300 2350
rect 13812 2310 13824 2344
rect 14288 2310 14300 2344
rect 13812 2304 14300 2310
rect 13514 2204 13530 2260
rect 13524 1684 13530 2204
rect 13564 2204 13574 2260
rect 14534 2260 14594 2410
rect 15032 2350 15092 2828
rect 16570 2650 16630 2918
rect 17596 2918 17602 3442
rect 17636 3442 17652 3494
rect 18606 3494 18666 3632
rect 19116 3584 19176 3848
rect 20138 3908 20200 3914
rect 20198 3848 20200 3908
rect 20138 3842 20200 3848
rect 19614 3752 19620 3812
rect 19680 3752 19686 3812
rect 18902 3578 19390 3584
rect 18902 3544 18914 3578
rect 19378 3544 19390 3578
rect 18902 3538 19390 3544
rect 18606 3454 18620 3494
rect 17636 2918 17642 3442
rect 18614 2972 18620 3454
rect 17596 2906 17642 2918
rect 18608 2918 18620 2972
rect 18654 3454 18666 3494
rect 19620 3494 19680 3752
rect 20140 3584 20200 3842
rect 20640 3692 20700 4150
rect 21658 4150 21674 4206
rect 21708 4700 21722 4726
rect 22680 4726 22740 5080
rect 22974 4810 23462 4816
rect 22974 4776 22986 4810
rect 23450 4776 23462 4810
rect 22974 4770 23462 4776
rect 23992 4810 24480 4816
rect 23992 4776 24004 4810
rect 24468 4776 24480 4810
rect 23992 4770 24480 4776
rect 21708 4206 21714 4700
rect 22680 4694 22692 4726
rect 21708 4150 21718 4206
rect 20938 4100 21426 4106
rect 20938 4066 20950 4100
rect 21414 4066 21426 4100
rect 20938 4060 21426 4066
rect 21142 3908 21202 4060
rect 21488 4026 21548 4032
rect 21658 4026 21718 4150
rect 22686 4150 22692 4694
rect 22726 4694 22740 4726
rect 23704 4726 23750 4738
rect 22726 4150 22732 4694
rect 23704 4220 23710 4726
rect 22686 4138 22732 4150
rect 23700 4150 23710 4220
rect 23744 4220 23750 4726
rect 24716 4726 24776 5080
rect 26258 5042 26318 5294
rect 26752 5252 26812 5384
rect 27776 5384 27782 5924
rect 27816 5384 27822 5960
rect 28786 5960 28846 6094
rect 29264 6050 29324 6528
rect 29806 6478 29866 6618
rect 30820 6618 30836 6662
rect 30870 6662 30876 7194
rect 31838 7194 31898 7328
rect 32136 7278 32624 7284
rect 32136 7244 32148 7278
rect 32612 7244 32624 7278
rect 32136 7238 32624 7244
rect 31838 7144 31854 7194
rect 30870 6618 30880 6662
rect 31848 6646 31854 7144
rect 30100 6568 30588 6574
rect 30100 6534 30112 6568
rect 30576 6534 30588 6568
rect 30100 6528 30588 6534
rect 29800 6418 29806 6478
rect 29866 6418 29872 6478
rect 29796 6310 29802 6370
rect 29862 6310 29868 6370
rect 29082 6044 29570 6050
rect 29082 6010 29094 6044
rect 29558 6010 29570 6044
rect 29082 6004 29570 6010
rect 28786 5866 28800 5960
rect 28794 5426 28800 5866
rect 27776 5372 27822 5384
rect 28786 5384 28800 5426
rect 28834 5866 28846 5960
rect 29802 5960 29862 6310
rect 30288 6196 30294 6256
rect 30354 6196 30360 6256
rect 30294 6050 30354 6196
rect 30820 6154 30880 6618
rect 31844 6618 31854 6646
rect 31888 7144 31898 7194
rect 32860 7194 32920 7524
rect 33154 7278 33642 7284
rect 33154 7244 33166 7278
rect 33630 7244 33642 7278
rect 33154 7238 33642 7244
rect 31888 6646 31894 7144
rect 32860 7142 32872 7194
rect 32866 6646 32872 7142
rect 31888 6618 31904 6646
rect 31118 6568 31606 6574
rect 31118 6534 31130 6568
rect 31594 6534 31606 6568
rect 31118 6528 31606 6534
rect 31844 6478 31904 6618
rect 32860 6618 32872 6646
rect 32906 7142 32920 7194
rect 33884 7194 33930 7206
rect 32906 6646 32912 7142
rect 33884 6652 33890 7194
rect 32906 6618 32920 6646
rect 32136 6568 32624 6574
rect 32136 6534 32148 6568
rect 32612 6534 32624 6568
rect 32136 6528 32624 6534
rect 31838 6418 31844 6478
rect 31904 6418 31910 6478
rect 31834 6310 31840 6370
rect 31900 6310 31906 6370
rect 31326 6196 31332 6256
rect 31392 6196 31398 6256
rect 30814 6094 30820 6154
rect 30880 6094 30886 6154
rect 31332 6050 31392 6196
rect 30100 6044 30588 6050
rect 30100 6010 30112 6044
rect 30576 6010 30588 6044
rect 30100 6004 30588 6010
rect 31118 6044 31606 6050
rect 31118 6010 31130 6044
rect 31594 6010 31606 6044
rect 31118 6004 31606 6010
rect 29802 5894 29818 5960
rect 28834 5426 28840 5866
rect 28834 5384 28846 5426
rect 27046 5334 27534 5340
rect 27046 5300 27058 5334
rect 27522 5300 27534 5334
rect 27046 5294 27534 5300
rect 28064 5334 28552 5340
rect 28064 5300 28076 5334
rect 28540 5300 28552 5334
rect 28064 5294 28552 5300
rect 26746 5192 26752 5252
rect 26812 5192 26818 5252
rect 27100 5192 27106 5252
rect 27166 5192 27172 5252
rect 26742 5080 26748 5140
rect 26808 5080 26814 5140
rect 26252 4982 26258 5042
rect 26318 4982 26324 5042
rect 25010 4810 25498 4816
rect 25010 4776 25022 4810
rect 25486 4776 25498 4810
rect 25010 4770 25498 4776
rect 26028 4810 26516 4816
rect 26028 4776 26040 4810
rect 26504 4776 26516 4810
rect 26028 4770 26516 4776
rect 24716 4688 24728 4726
rect 23744 4150 23760 4220
rect 21956 4100 22444 4106
rect 21956 4066 21968 4100
rect 22432 4066 22444 4100
rect 21956 4060 22444 4066
rect 22974 4100 23462 4106
rect 22974 4066 22986 4100
rect 23450 4066 23462 4100
rect 22974 4060 23462 4066
rect 21652 3966 21658 4026
rect 21718 3966 21724 4026
rect 21136 3848 21142 3908
rect 21202 3848 21208 3908
rect 20634 3632 20640 3692
rect 20700 3632 20706 3692
rect 19920 3578 20408 3584
rect 19920 3544 19932 3578
rect 20396 3544 20408 3578
rect 19920 3538 20408 3544
rect 18654 2972 18660 3454
rect 19620 3434 19638 3494
rect 18654 2918 18668 2972
rect 16866 2868 17354 2874
rect 16866 2834 16878 2868
rect 17342 2834 17354 2868
rect 16866 2828 17354 2834
rect 17884 2868 18372 2874
rect 17884 2834 17896 2868
rect 18360 2834 18372 2868
rect 17884 2828 18372 2834
rect 17090 2662 17150 2828
rect 16564 2590 16570 2650
rect 16630 2590 16636 2650
rect 17084 2602 17090 2662
rect 17150 2602 17156 2662
rect 15546 2488 15552 2548
rect 15612 2488 15618 2548
rect 17582 2488 17588 2548
rect 17648 2488 17654 2548
rect 14830 2344 15318 2350
rect 14830 2310 14842 2344
rect 15306 2310 15318 2344
rect 14830 2304 15318 2310
rect 13564 1684 13570 2204
rect 13524 1672 13570 1684
rect 14534 1684 14548 2260
rect 14582 1684 14594 2260
rect 15552 2260 15612 2488
rect 16564 2384 16570 2444
rect 16630 2384 16636 2444
rect 15848 2344 16336 2350
rect 15848 2310 15860 2344
rect 16324 2310 16336 2344
rect 15848 2304 16336 2310
rect 15552 2200 15566 2260
rect 15560 1720 15566 2200
rect 13812 1634 14300 1640
rect 13812 1600 13824 1634
rect 14288 1600 14300 1634
rect 13812 1594 14300 1600
rect 13392 1486 13398 1546
rect 13458 1486 13464 1546
rect 13064 1382 13070 1442
rect 13130 1382 13136 1442
rect 13398 1216 13458 1486
rect 14534 1442 14594 1684
rect 15554 1684 15566 1720
rect 15600 2200 15612 2260
rect 16570 2260 16630 2384
rect 16866 2344 17354 2350
rect 16866 2310 16878 2344
rect 17342 2310 17354 2344
rect 16866 2304 17354 2310
rect 16570 2206 16584 2260
rect 15600 1720 15606 2200
rect 16578 1724 16584 2206
rect 15600 1684 15614 1720
rect 14830 1634 15318 1640
rect 14830 1600 14842 1634
rect 15306 1600 15318 1634
rect 14830 1594 15318 1600
rect 14528 1382 14534 1442
rect 14594 1382 14600 1442
rect 15042 1336 15102 1594
rect 15036 1276 15042 1336
rect 15102 1276 15108 1336
rect 13398 1156 14598 1216
rect 12014 322 12020 382
rect 12080 322 12086 382
rect 13398 304 13458 1156
rect 13518 1028 13578 1156
rect 14004 1118 14064 1156
rect 13812 1112 14300 1118
rect 13812 1078 13824 1112
rect 14288 1078 14300 1112
rect 13812 1072 14300 1078
rect 13518 956 13530 1028
rect 13524 452 13530 956
rect 13564 956 13578 1028
rect 14538 1028 14598 1156
rect 15042 1118 15102 1276
rect 15554 1226 15614 1684
rect 16568 1684 16584 1724
rect 16618 2206 16630 2260
rect 17588 2260 17648 2488
rect 18090 2350 18150 2828
rect 18608 2548 18668 2918
rect 19632 2918 19638 3434
rect 19672 3434 19680 3494
rect 20640 3494 20700 3632
rect 21142 3584 21202 3848
rect 21488 3812 21548 3966
rect 21482 3752 21488 3812
rect 21548 3752 21554 3812
rect 21658 3758 21664 3818
rect 21724 3758 21730 3818
rect 20938 3578 21426 3584
rect 20938 3544 20950 3578
rect 21414 3544 21426 3578
rect 20938 3538 21426 3544
rect 20640 3454 20656 3494
rect 19672 2918 19678 3434
rect 20650 2984 20656 3454
rect 19632 2906 19678 2918
rect 20644 2918 20656 2984
rect 20690 3454 20700 3494
rect 21664 3494 21724 3758
rect 22180 3756 22240 4060
rect 23194 3920 23254 4060
rect 23700 4026 23760 4150
rect 24722 4150 24728 4688
rect 24762 4688 24776 4726
rect 25740 4726 25786 4738
rect 24762 4150 24768 4688
rect 25740 4220 25746 4726
rect 24722 4138 24768 4150
rect 25732 4150 25746 4220
rect 25780 4220 25786 4726
rect 26748 4726 26808 5080
rect 27106 4934 27166 5192
rect 27296 5042 27356 5294
rect 28272 5042 28332 5294
rect 27290 4982 27296 5042
rect 27356 4982 27362 5042
rect 28266 4982 28272 5042
rect 28332 4982 28338 5042
rect 28786 4930 28846 5384
rect 29812 5384 29818 5894
rect 29852 5894 29862 5960
rect 30830 5960 30876 5972
rect 29852 5384 29858 5894
rect 30830 5428 30836 5960
rect 29812 5372 29858 5384
rect 30824 5384 30836 5428
rect 30870 5428 30876 5960
rect 31840 5960 31900 6310
rect 32358 6256 32418 6528
rect 32860 6436 32920 6618
rect 33874 6618 33890 6652
rect 33924 6652 33930 7194
rect 33924 6618 33934 6652
rect 33154 6568 33642 6574
rect 33154 6534 33166 6568
rect 33630 6534 33642 6568
rect 33154 6528 33642 6534
rect 33368 6436 33428 6528
rect 33874 6436 33934 6618
rect 32860 6376 33934 6436
rect 32352 6196 32358 6256
rect 32418 6196 32424 6256
rect 32856 6094 32862 6154
rect 32922 6094 32928 6154
rect 32136 6044 32624 6050
rect 32136 6010 32148 6044
rect 32612 6010 32624 6044
rect 32136 6004 32624 6010
rect 31840 5908 31854 5960
rect 31848 5434 31854 5908
rect 30870 5384 30884 5428
rect 29082 5334 29570 5340
rect 29082 5300 29094 5334
rect 29558 5300 29570 5334
rect 29082 5294 29570 5300
rect 30100 5334 30588 5340
rect 30100 5300 30112 5334
rect 30576 5300 30588 5334
rect 30100 5294 30588 5300
rect 29288 5042 29348 5294
rect 30824 5252 30884 5384
rect 31842 5384 31854 5434
rect 31888 5908 31900 5960
rect 32862 5960 32922 6094
rect 33154 6044 33642 6050
rect 33154 6010 33166 6044
rect 33630 6010 33642 6044
rect 33154 6004 33642 6010
rect 32862 5926 32872 5960
rect 31888 5434 31894 5908
rect 31888 5384 31902 5434
rect 32866 5428 32872 5926
rect 31118 5334 31606 5340
rect 31118 5300 31130 5334
rect 31594 5300 31606 5334
rect 31118 5294 31606 5300
rect 30818 5192 30824 5252
rect 30884 5192 30890 5252
rect 29282 4982 29288 5042
rect 29348 4982 29354 5042
rect 31308 4982 31314 5042
rect 31374 4982 31380 5042
rect 27106 4868 27166 4874
rect 28780 4870 28786 4930
rect 28846 4870 28852 4930
rect 30816 4870 30822 4930
rect 30882 4870 30888 4930
rect 27046 4810 27534 4816
rect 27046 4776 27058 4810
rect 27522 4776 27534 4810
rect 27046 4770 27534 4776
rect 28064 4810 28552 4816
rect 28064 4776 28076 4810
rect 28540 4776 28552 4810
rect 28064 4770 28552 4776
rect 26748 4684 26764 4726
rect 25780 4150 25792 4220
rect 23992 4100 24480 4106
rect 23992 4066 24004 4100
rect 24468 4066 24480 4100
rect 23992 4060 24480 4066
rect 25010 4100 25498 4106
rect 25010 4066 25022 4100
rect 25486 4066 25498 4100
rect 25010 4060 25498 4066
rect 23694 3966 23700 4026
rect 23760 3966 23766 4026
rect 24216 3920 24276 4060
rect 25230 3920 25290 4060
rect 25732 4026 25792 4150
rect 26758 4150 26764 4684
rect 26798 4684 26808 4726
rect 27776 4726 27822 4738
rect 26798 4150 26804 4684
rect 27776 4186 27782 4726
rect 26758 4138 26804 4150
rect 27772 4150 27782 4186
rect 27816 4186 27822 4726
rect 28786 4726 28846 4870
rect 29082 4810 29570 4816
rect 29082 4776 29094 4810
rect 29558 4776 29570 4810
rect 29082 4770 29570 4776
rect 30100 4810 30588 4816
rect 30100 4776 30112 4810
rect 30576 4776 30588 4810
rect 30100 4770 30588 4776
rect 28786 4688 28800 4726
rect 28794 4202 28800 4688
rect 27816 4150 27832 4186
rect 26028 4100 26516 4106
rect 26028 4066 26040 4100
rect 26504 4066 26516 4100
rect 26028 4060 26516 4066
rect 27046 4100 27534 4106
rect 27046 4066 27058 4100
rect 27522 4066 27534 4100
rect 27046 4060 27534 4066
rect 25726 3966 25732 4026
rect 25792 3966 25798 4026
rect 26232 4020 26292 4060
rect 27258 4020 27318 4060
rect 27772 4026 27832 4150
rect 28790 4150 28800 4202
rect 28834 4688 28846 4726
rect 29812 4726 29858 4738
rect 28834 4202 28840 4688
rect 28834 4150 28850 4202
rect 29812 4194 29818 4726
rect 28064 4100 28552 4106
rect 28064 4066 28076 4100
rect 28540 4066 28552 4100
rect 28064 4060 28552 4066
rect 26232 3960 27318 4020
rect 27766 3966 27772 4026
rect 27832 3966 27838 4026
rect 26232 3920 26292 3960
rect 23194 3860 26292 3920
rect 26744 3868 26750 3928
rect 26810 3868 26816 3928
rect 23194 3756 23254 3860
rect 23686 3758 23692 3818
rect 23752 3758 23758 3818
rect 22180 3696 23254 3756
rect 22180 3584 22240 3696
rect 23194 3584 23254 3696
rect 21956 3578 22444 3584
rect 21956 3544 21968 3578
rect 22432 3544 22444 3578
rect 21956 3538 22444 3544
rect 22974 3578 23462 3584
rect 22974 3544 22986 3578
rect 23450 3544 23462 3578
rect 22974 3538 23462 3544
rect 20690 2984 20696 3454
rect 21664 3450 21674 3494
rect 20690 2918 20704 2984
rect 21668 2976 21674 3450
rect 18902 2868 19390 2874
rect 18902 2834 18914 2868
rect 19378 2834 19390 2868
rect 18902 2828 19390 2834
rect 19920 2868 20408 2874
rect 19920 2834 19932 2868
rect 20396 2834 20408 2868
rect 19920 2828 20408 2834
rect 18602 2488 18608 2548
rect 18668 2488 18674 2548
rect 19112 2350 19172 2828
rect 19618 2488 19624 2548
rect 19684 2488 19690 2548
rect 17884 2344 18372 2350
rect 17884 2310 17896 2344
rect 18360 2310 18372 2344
rect 17884 2304 18372 2310
rect 18902 2344 19390 2350
rect 18902 2310 18914 2344
rect 19378 2310 19390 2344
rect 18902 2304 19390 2310
rect 17588 2210 17602 2260
rect 16618 1724 16624 2206
rect 16618 1684 16628 1724
rect 17596 1708 17602 2210
rect 15848 1634 16336 1640
rect 15848 1600 15860 1634
rect 16324 1600 16336 1634
rect 15848 1594 16336 1600
rect 16062 1336 16122 1594
rect 16568 1546 16628 1684
rect 17590 1684 17602 1708
rect 17636 2210 17648 2260
rect 18614 2260 18660 2272
rect 17636 1708 17642 2210
rect 17636 1684 17650 1708
rect 18614 1698 18620 2260
rect 16866 1634 17354 1640
rect 16866 1600 16878 1634
rect 17342 1600 17354 1634
rect 16866 1594 17354 1600
rect 16562 1486 16568 1546
rect 16628 1486 16634 1546
rect 16568 1382 16574 1442
rect 16634 1382 16640 1442
rect 16056 1276 16062 1336
rect 16122 1276 16128 1336
rect 15548 1166 15554 1226
rect 15614 1166 15620 1226
rect 14830 1112 15318 1118
rect 14830 1078 14842 1112
rect 15306 1078 15318 1112
rect 14830 1072 15318 1078
rect 13564 452 13570 956
rect 14538 952 14548 1028
rect 14542 500 14548 952
rect 13524 440 13570 452
rect 14534 452 14548 500
rect 14582 952 14598 1028
rect 15554 1028 15614 1166
rect 16062 1118 16122 1276
rect 15848 1112 16336 1118
rect 15848 1078 15860 1112
rect 16324 1078 16336 1112
rect 15848 1072 16336 1078
rect 14582 500 14588 952
rect 14582 452 14594 500
rect 13812 402 14300 408
rect 13812 368 13824 402
rect 14288 368 14300 402
rect 13812 362 14300 368
rect 14534 304 14594 452
rect 15554 452 15566 1028
rect 15600 452 15614 1028
rect 16574 1028 16634 1382
rect 17086 1336 17146 1594
rect 17080 1276 17086 1336
rect 17146 1276 17152 1336
rect 17086 1118 17146 1276
rect 17590 1226 17650 1684
rect 18604 1684 18620 1698
rect 18654 1698 18660 2260
rect 19624 2260 19684 2488
rect 20124 2350 20184 2828
rect 20644 2548 20704 2918
rect 21656 2918 21674 2976
rect 21708 3450 21724 3494
rect 22686 3494 22732 3506
rect 21708 2976 21714 3450
rect 21708 2918 21716 2976
rect 22686 2970 22692 3494
rect 20938 2868 21426 2874
rect 20938 2834 20950 2868
rect 21414 2834 21426 2868
rect 20938 2828 21426 2834
rect 20638 2488 20644 2548
rect 20704 2488 20710 2548
rect 21154 2350 21214 2828
rect 21656 2716 21716 2918
rect 22674 2918 22692 2970
rect 22726 2970 22732 3494
rect 23692 3494 23752 3758
rect 24216 3584 24276 3860
rect 25230 3584 25290 3860
rect 25730 3758 25736 3818
rect 25796 3758 25802 3818
rect 23992 3578 24480 3584
rect 23992 3544 24004 3578
rect 24468 3544 24480 3578
rect 23992 3538 24480 3544
rect 25010 3578 25498 3584
rect 25010 3544 25022 3578
rect 25486 3544 25498 3578
rect 25010 3538 25498 3544
rect 23692 3450 23710 3494
rect 22726 2918 22734 2970
rect 21956 2868 22444 2874
rect 21956 2834 21968 2868
rect 22432 2834 22444 2868
rect 21956 2828 22444 2834
rect 21506 2656 21716 2716
rect 22170 2662 22230 2828
rect 22674 2776 22734 2918
rect 23704 2918 23710 3450
rect 23744 3450 23752 3494
rect 24722 3494 24768 3506
rect 23744 2918 23750 3450
rect 24722 2970 24728 3494
rect 23704 2906 23750 2918
rect 24716 2918 24728 2970
rect 24762 2970 24768 3494
rect 25736 3494 25796 3758
rect 26232 3584 26292 3860
rect 26028 3578 26516 3584
rect 26028 3544 26040 3578
rect 26504 3544 26516 3578
rect 26028 3538 26516 3544
rect 25736 3446 25746 3494
rect 24762 2918 24776 2970
rect 22974 2868 23462 2874
rect 22974 2834 22986 2868
rect 23450 2834 23462 2868
rect 22974 2828 23462 2834
rect 23992 2868 24480 2874
rect 23992 2834 24004 2868
rect 24468 2834 24480 2868
rect 23992 2828 24480 2834
rect 24716 2776 24776 2918
rect 25740 2918 25746 3446
rect 25780 3446 25796 3494
rect 26750 3494 26810 3868
rect 27258 3584 27318 3960
rect 27758 3758 27764 3818
rect 27824 3758 27830 3818
rect 27046 3578 27534 3584
rect 27046 3544 27058 3578
rect 27522 3544 27534 3578
rect 27046 3538 27534 3544
rect 26750 3458 26764 3494
rect 25780 2918 25786 3446
rect 26758 2962 26764 3458
rect 25740 2906 25786 2918
rect 26752 2918 26764 2962
rect 26798 3458 26810 3494
rect 27764 3494 27824 3758
rect 28278 3584 28338 4060
rect 28790 3692 28850 4150
rect 29802 4150 29818 4194
rect 29852 4194 29858 4726
rect 30822 4726 30882 4870
rect 31314 4816 31374 4982
rect 31118 4810 31606 4816
rect 31118 4776 31130 4810
rect 31594 4776 31606 4810
rect 31118 4770 31606 4776
rect 30822 4668 30836 4726
rect 29852 4150 29862 4194
rect 30830 4190 30836 4668
rect 29082 4100 29570 4106
rect 29082 4066 29094 4100
rect 29558 4066 29570 4100
rect 29082 4060 29570 4066
rect 28784 3632 28790 3692
rect 28850 3632 28856 3692
rect 28064 3578 28552 3584
rect 28064 3544 28076 3578
rect 28540 3544 28552 3578
rect 28064 3538 28552 3544
rect 26798 2962 26804 3458
rect 27764 3446 27782 3494
rect 26798 2918 26812 2962
rect 27776 2958 27782 3446
rect 25010 2868 25498 2874
rect 25010 2834 25022 2868
rect 25486 2834 25498 2868
rect 25010 2828 25498 2834
rect 26028 2868 26516 2874
rect 26028 2834 26040 2868
rect 26504 2834 26516 2868
rect 26028 2828 26516 2834
rect 26752 2776 26812 2918
rect 27766 2918 27782 2958
rect 27816 3446 27824 3494
rect 28790 3494 28850 3632
rect 29294 3584 29354 4060
rect 29802 3818 29862 4150
rect 30820 4150 30836 4190
rect 30870 4668 30882 4726
rect 31842 4726 31902 5384
rect 32858 5384 32872 5428
rect 32906 5926 32922 5960
rect 33884 5960 33930 5972
rect 32906 5428 32912 5926
rect 32906 5384 32918 5428
rect 33884 5414 33890 5960
rect 32136 5334 32624 5340
rect 32136 5300 32148 5334
rect 32612 5300 32624 5334
rect 32136 5294 32624 5300
rect 32344 5042 32404 5294
rect 32858 5202 32918 5384
rect 33874 5384 33890 5414
rect 33924 5414 33930 5960
rect 33924 5384 33934 5414
rect 33154 5334 33642 5340
rect 33154 5300 33166 5334
rect 33630 5300 33642 5334
rect 33154 5294 33642 5300
rect 33364 5202 33424 5294
rect 33874 5202 33934 5384
rect 32858 5142 33934 5202
rect 32338 4982 32344 5042
rect 32404 4982 32410 5042
rect 32858 4930 32918 5142
rect 32852 4870 32858 4930
rect 32918 4870 32924 4930
rect 32136 4810 32624 4816
rect 32136 4776 32148 4810
rect 32612 4776 32624 4810
rect 32136 4770 32624 4776
rect 33154 4810 33642 4816
rect 33154 4776 33166 4810
rect 33630 4776 33642 4810
rect 33154 4770 33642 4776
rect 31842 4684 31854 4726
rect 30870 4190 30876 4668
rect 31848 4204 31854 4684
rect 30870 4150 30880 4190
rect 30100 4100 30588 4106
rect 30100 4066 30112 4100
rect 30576 4066 30588 4100
rect 30100 4060 30588 4066
rect 29796 3758 29802 3818
rect 29862 3758 29868 3818
rect 30328 3584 30388 4060
rect 30820 3692 30880 4150
rect 31842 4150 31854 4204
rect 31888 4684 31902 4726
rect 32866 4726 32912 4738
rect 31888 4204 31894 4684
rect 31888 4150 31902 4204
rect 32866 4196 32872 4726
rect 31118 4100 31606 4106
rect 31118 4066 31130 4100
rect 31594 4066 31606 4100
rect 31118 4060 31606 4066
rect 31346 3694 31406 4060
rect 31842 3818 31902 4150
rect 32856 4150 32872 4196
rect 32906 4196 32912 4726
rect 33884 4726 33930 4738
rect 32906 4150 32916 4196
rect 33884 4178 33890 4726
rect 32136 4100 32624 4106
rect 32136 4066 32148 4100
rect 32612 4066 32624 4100
rect 32136 4060 32624 4066
rect 32360 3822 32420 4060
rect 32856 4024 32916 4150
rect 33876 4150 33890 4178
rect 33924 4178 33930 4726
rect 33924 4150 33936 4178
rect 33154 4100 33642 4106
rect 33154 4066 33166 4100
rect 33630 4066 33642 4100
rect 33154 4060 33642 4066
rect 33362 4026 33422 4060
rect 33876 4026 33936 4150
rect 33362 4024 33936 4026
rect 32856 3964 33936 4024
rect 32856 3928 32916 3964
rect 32850 3868 32856 3928
rect 32916 3868 32922 3928
rect 31836 3758 31842 3818
rect 31902 3758 31908 3818
rect 32354 3762 32360 3822
rect 32420 3762 32426 3822
rect 33866 3762 33872 3822
rect 33932 3762 33938 3822
rect 30814 3632 30820 3692
rect 30880 3632 30886 3692
rect 29082 3578 29570 3584
rect 29082 3544 29094 3578
rect 29558 3544 29570 3578
rect 29082 3538 29570 3544
rect 30100 3578 30588 3584
rect 30100 3544 30112 3578
rect 30576 3544 30588 3578
rect 30100 3538 30588 3544
rect 28790 3448 28800 3494
rect 27816 2958 27822 3446
rect 28794 2978 28800 3448
rect 27816 2918 27826 2958
rect 27046 2868 27534 2874
rect 27046 2834 27058 2868
rect 27522 2834 27534 2868
rect 27046 2828 27534 2834
rect 22668 2716 22674 2776
rect 22734 2716 22740 2776
rect 24710 2716 24716 2776
rect 24776 2716 24782 2776
rect 26746 2716 26752 2776
rect 26812 2716 26818 2776
rect 27258 2666 27318 2828
rect 27766 2768 27826 2918
rect 28788 2918 28800 2978
rect 28834 3448 28850 3494
rect 29812 3494 29858 3506
rect 28834 2978 28840 3448
rect 28834 2918 28848 2978
rect 29812 2962 29818 3494
rect 28064 2868 28552 2874
rect 28064 2834 28076 2868
rect 28540 2834 28552 2868
rect 28064 2828 28552 2834
rect 27766 2708 27972 2768
rect 21506 2444 21566 2656
rect 22164 2602 22170 2662
rect 22230 2602 22236 2662
rect 27252 2606 27258 2666
rect 27318 2606 27324 2666
rect 21656 2488 21662 2548
rect 21722 2488 21728 2548
rect 23686 2488 23692 2548
rect 23752 2488 23758 2548
rect 25724 2488 25730 2548
rect 25790 2488 25796 2548
rect 27760 2488 27766 2548
rect 27826 2488 27832 2548
rect 21500 2384 21506 2444
rect 21566 2384 21572 2444
rect 19920 2344 20408 2350
rect 19920 2310 19932 2344
rect 20396 2310 20408 2344
rect 19920 2304 20408 2310
rect 20938 2344 21426 2350
rect 20938 2310 20950 2344
rect 21414 2310 21426 2344
rect 20938 2304 21426 2310
rect 19624 1778 19638 2260
rect 19632 1704 19638 1778
rect 18654 1684 18664 1698
rect 17884 1634 18372 1640
rect 17884 1600 17896 1634
rect 18360 1600 18372 1634
rect 17884 1594 18372 1600
rect 18104 1336 18164 1594
rect 18604 1442 18664 1684
rect 19628 1684 19638 1704
rect 19672 1778 19684 2260
rect 20650 2260 20696 2272
rect 19672 1704 19678 1778
rect 20650 1710 20656 2260
rect 19672 1684 19688 1704
rect 18902 1634 19390 1640
rect 18902 1600 18914 1634
rect 19378 1600 19390 1634
rect 18902 1594 19390 1600
rect 18598 1382 18604 1442
rect 18664 1382 18670 1442
rect 19118 1336 19178 1594
rect 18098 1276 18104 1336
rect 18164 1276 18170 1336
rect 19112 1276 19118 1336
rect 19178 1276 19184 1336
rect 17584 1166 17590 1226
rect 17650 1166 17656 1226
rect 16866 1112 17354 1118
rect 16866 1078 16878 1112
rect 17342 1078 17354 1112
rect 16866 1072 17354 1078
rect 16574 1014 16584 1028
rect 14830 402 15318 408
rect 14830 368 14842 402
rect 15306 368 15318 402
rect 14830 362 15318 368
rect 13392 244 13398 304
rect 13458 244 13464 304
rect 14528 244 14534 304
rect 14594 244 14600 304
rect 15046 196 15106 362
rect 15040 136 15046 196
rect 15106 136 15112 196
rect 15554 -60 15614 452
rect 16578 452 16584 1014
rect 16618 1014 16634 1028
rect 17590 1028 17650 1166
rect 18104 1118 18164 1276
rect 19118 1118 19178 1276
rect 19628 1226 19688 1684
rect 20644 1684 20656 1710
rect 20690 1710 20696 2260
rect 21662 2260 21722 2488
rect 21956 2344 22444 2350
rect 21956 2310 21968 2344
rect 22432 2310 22444 2344
rect 21956 2304 22444 2310
rect 22974 2344 23462 2350
rect 22974 2310 22986 2344
rect 23450 2310 23462 2344
rect 22974 2304 23462 2310
rect 22686 2260 22732 2272
rect 23692 2260 23752 2488
rect 23992 2344 24480 2350
rect 23992 2310 24004 2344
rect 24468 2310 24480 2344
rect 23992 2304 24480 2310
rect 25010 2344 25498 2350
rect 25010 2310 25022 2344
rect 25486 2310 25498 2344
rect 25010 2304 25498 2310
rect 24722 2260 24768 2272
rect 25730 2260 25790 2488
rect 26028 2344 26516 2350
rect 26028 2310 26040 2344
rect 26504 2310 26516 2344
rect 26028 2304 26516 2310
rect 27046 2344 27534 2350
rect 27046 2310 27058 2344
rect 27522 2310 27534 2344
rect 27046 2304 27534 2310
rect 21662 2204 21674 2260
rect 20690 1684 20704 1710
rect 21668 1708 21674 2204
rect 19920 1634 20408 1640
rect 19920 1600 19932 1634
rect 20396 1600 20408 1634
rect 19920 1594 20408 1600
rect 20150 1336 20210 1594
rect 20644 1442 20704 1684
rect 21666 1684 21674 1708
rect 21708 2204 21722 2260
rect 22680 2224 22692 2260
rect 21708 1708 21714 2204
rect 22686 1736 22692 2224
rect 21708 1684 21726 1708
rect 20938 1634 21426 1640
rect 20938 1600 20950 1634
rect 21414 1600 21426 1634
rect 20938 1594 21426 1600
rect 20792 1488 20798 1548
rect 20858 1488 20864 1548
rect 20638 1382 20644 1442
rect 20704 1382 20710 1442
rect 20144 1276 20150 1336
rect 20210 1276 20216 1336
rect 20798 1304 20858 1488
rect 21162 1336 21222 1594
rect 19622 1166 19628 1226
rect 19688 1166 19694 1226
rect 17884 1112 18372 1118
rect 17884 1078 17896 1112
rect 18360 1078 18372 1112
rect 17884 1072 18372 1078
rect 18902 1112 19390 1118
rect 18902 1078 18914 1112
rect 19378 1078 19390 1112
rect 18902 1072 19390 1078
rect 16618 452 16624 1014
rect 16578 440 16624 452
rect 17590 452 17602 1028
rect 17636 452 17650 1028
rect 18614 1028 18660 1040
rect 18614 494 18620 1028
rect 15848 402 16336 408
rect 15848 368 15860 402
rect 16324 368 16336 402
rect 15848 362 16336 368
rect 16866 402 17354 408
rect 16866 368 16878 402
rect 17342 368 17354 402
rect 16866 362 17354 368
rect 16060 196 16120 362
rect 16060 130 16120 136
rect 17082 196 17142 362
rect 17082 130 17142 136
rect 17590 -60 17650 452
rect 18604 452 18620 494
rect 18654 494 18660 1028
rect 19628 1028 19688 1166
rect 20150 1118 20210 1276
rect 20642 1244 20858 1304
rect 21156 1276 21162 1336
rect 21222 1276 21228 1336
rect 19920 1112 20408 1118
rect 19920 1078 19932 1112
rect 20396 1078 20408 1112
rect 19920 1072 20408 1078
rect 18654 452 18664 494
rect 17884 402 18372 408
rect 17884 368 17896 402
rect 18360 368 18372 402
rect 17884 362 18372 368
rect 18094 202 18154 362
rect 18604 304 18664 452
rect 19628 452 19638 1028
rect 19672 452 19688 1028
rect 20642 1028 20702 1244
rect 21162 1118 21222 1276
rect 21666 1226 21726 1684
rect 22676 1684 22692 1736
rect 22726 2224 22740 2260
rect 22726 1736 22732 2224
rect 23692 2210 23710 2260
rect 22726 1684 22736 1736
rect 23704 1714 23710 2210
rect 21956 1634 22444 1640
rect 21956 1600 21968 1634
rect 22432 1600 22444 1634
rect 21956 1594 22444 1600
rect 22170 1336 22230 1594
rect 22676 1548 22736 1684
rect 23702 1684 23710 1714
rect 23744 2210 23752 2260
rect 24716 2228 24728 2260
rect 23744 1714 23750 2210
rect 24722 1724 24728 2228
rect 23744 1684 23762 1714
rect 22974 1634 23462 1640
rect 22974 1600 22986 1634
rect 23450 1600 23462 1634
rect 22974 1594 23462 1600
rect 22670 1488 22676 1548
rect 22736 1488 22742 1548
rect 22674 1382 22680 1442
rect 22740 1382 22746 1442
rect 22164 1276 22170 1336
rect 22230 1276 22236 1336
rect 21660 1166 21666 1226
rect 21726 1166 21732 1226
rect 20938 1112 21426 1118
rect 20938 1078 20950 1112
rect 21414 1078 21426 1112
rect 20938 1072 21426 1078
rect 20642 1002 20656 1028
rect 18902 402 19390 408
rect 18902 368 18914 402
rect 19378 368 19390 402
rect 18902 362 19390 368
rect 18598 244 18604 304
rect 18664 244 18670 304
rect 19120 202 19180 362
rect 18094 196 18156 202
rect 18094 190 18096 196
rect 19120 196 19182 202
rect 19120 190 19122 196
rect 18096 130 18156 136
rect 19122 130 19182 136
rect 19628 -60 19688 452
rect 20650 452 20656 1002
rect 20690 1002 20702 1028
rect 21666 1028 21726 1166
rect 22170 1118 22230 1276
rect 21956 1112 22444 1118
rect 21956 1078 21968 1112
rect 22432 1078 22444 1112
rect 21956 1072 22444 1078
rect 20690 452 20696 1002
rect 20650 440 20696 452
rect 21666 452 21674 1028
rect 21708 452 21726 1028
rect 22680 1028 22740 1382
rect 23188 1336 23248 1594
rect 23182 1276 23188 1336
rect 23248 1276 23254 1336
rect 23188 1118 23248 1276
rect 23702 1226 23762 1684
rect 24714 1684 24728 1724
rect 24762 2228 24776 2260
rect 24762 1724 24768 2228
rect 25730 2216 25746 2260
rect 24762 1684 24774 1724
rect 25740 1708 25746 2216
rect 23992 1634 24480 1640
rect 23992 1600 24004 1634
rect 24468 1600 24480 1634
rect 23992 1594 24480 1600
rect 24214 1336 24274 1594
rect 24714 1548 24774 1684
rect 25738 1684 25746 1708
rect 25780 2216 25790 2260
rect 26758 2260 26804 2272
rect 25780 1708 25786 2216
rect 26758 1730 26764 2260
rect 25780 1684 25798 1708
rect 25010 1634 25498 1640
rect 25010 1600 25022 1634
rect 25486 1600 25498 1634
rect 25010 1594 25498 1600
rect 24708 1488 24714 1548
rect 24774 1488 24780 1548
rect 24710 1382 24716 1442
rect 24776 1382 24782 1442
rect 24208 1276 24214 1336
rect 24274 1276 24280 1336
rect 23696 1166 23702 1226
rect 23762 1166 23768 1226
rect 22974 1112 23462 1118
rect 22974 1078 22986 1112
rect 23450 1078 23462 1112
rect 22974 1072 23462 1078
rect 22680 1002 22692 1028
rect 19920 402 20408 408
rect 19920 368 19932 402
rect 20396 368 20408 402
rect 19920 362 20408 368
rect 20938 402 21426 408
rect 20938 368 20950 402
rect 21414 368 21426 402
rect 20938 362 21426 368
rect 20134 196 20194 362
rect 20134 130 20194 136
rect 21170 196 21230 362
rect 21170 130 21230 136
rect 21666 -60 21726 452
rect 22686 452 22692 1002
rect 22726 1002 22740 1028
rect 23702 1028 23762 1166
rect 24214 1118 24274 1276
rect 23992 1112 24480 1118
rect 23992 1078 24004 1112
rect 24468 1078 24480 1112
rect 23992 1072 24480 1078
rect 22726 452 22732 1002
rect 22686 440 22732 452
rect 23702 452 23710 1028
rect 23744 452 23762 1028
rect 24716 1028 24776 1382
rect 25216 1336 25276 1594
rect 25210 1276 25216 1336
rect 25276 1276 25282 1336
rect 25216 1118 25276 1276
rect 25738 1226 25798 1684
rect 26750 1684 26764 1730
rect 26798 1730 26804 2260
rect 27766 2260 27826 2488
rect 27912 2444 27972 2708
rect 27906 2384 27912 2444
rect 27972 2384 27978 2444
rect 28276 2350 28336 2828
rect 28788 2548 28848 2918
rect 29806 2918 29818 2962
rect 29852 2962 29858 3494
rect 30820 3494 30880 3632
rect 31346 3584 31406 3634
rect 32360 3584 32420 3762
rect 32854 3634 32860 3694
rect 32920 3634 32926 3694
rect 31118 3578 31606 3584
rect 31118 3544 31130 3578
rect 31594 3544 31606 3578
rect 31118 3538 31606 3544
rect 32136 3578 32624 3584
rect 32136 3544 32148 3578
rect 32612 3544 32624 3578
rect 32136 3538 32624 3544
rect 30820 3448 30836 3494
rect 30830 2966 30836 3448
rect 29852 2918 29866 2962
rect 29082 2868 29570 2874
rect 29082 2834 29094 2868
rect 29558 2834 29570 2868
rect 29082 2828 29570 2834
rect 28782 2488 28788 2548
rect 28848 2488 28854 2548
rect 29296 2350 29356 2828
rect 29806 2776 29866 2918
rect 30822 2918 30836 2966
rect 30870 3448 30880 3494
rect 31848 3494 31894 3506
rect 32860 3494 32920 3634
rect 33154 3578 33642 3584
rect 33154 3544 33166 3578
rect 33630 3544 33642 3578
rect 33154 3538 33642 3544
rect 30870 2966 30876 3448
rect 30870 2918 30882 2966
rect 31848 2962 31854 3494
rect 30100 2868 30588 2874
rect 30100 2834 30112 2868
rect 30576 2834 30588 2868
rect 30100 2828 30588 2834
rect 29800 2716 29806 2776
rect 29866 2716 29872 2776
rect 29802 2488 29808 2548
rect 29868 2488 29874 2548
rect 28064 2344 28552 2350
rect 28064 2310 28076 2344
rect 28540 2310 28552 2344
rect 28064 2304 28552 2310
rect 29082 2344 29570 2350
rect 29082 2310 29094 2344
rect 29558 2310 29570 2344
rect 29082 2304 29570 2310
rect 27766 2216 27782 2260
rect 26798 1684 26810 1730
rect 27776 1710 27782 2216
rect 26028 1634 26516 1640
rect 26028 1600 26040 1634
rect 26504 1600 26516 1634
rect 26028 1594 26516 1600
rect 26236 1336 26296 1594
rect 26578 1488 26584 1548
rect 26644 1488 26650 1548
rect 26230 1276 26236 1336
rect 26296 1276 26302 1336
rect 26584 1296 26644 1488
rect 26750 1442 26810 1684
rect 27770 1684 27782 1710
rect 27816 2216 27826 2260
rect 28794 2260 28840 2272
rect 27816 1710 27822 2216
rect 28794 1724 28800 2260
rect 27816 1684 27830 1710
rect 27046 1634 27534 1640
rect 27046 1600 27058 1634
rect 27522 1600 27534 1634
rect 27046 1594 27534 1600
rect 26744 1382 26750 1442
rect 26810 1382 26816 1442
rect 27256 1336 27316 1594
rect 25732 1166 25738 1226
rect 25798 1166 25804 1226
rect 25010 1112 25498 1118
rect 25010 1078 25022 1112
rect 25486 1078 25498 1112
rect 25010 1072 25498 1078
rect 24716 992 24728 1028
rect 21956 402 22444 408
rect 21956 368 21968 402
rect 22432 368 22444 402
rect 21956 362 22444 368
rect 22974 402 23462 408
rect 22974 368 22986 402
rect 23450 368 23462 402
rect 22974 362 23462 368
rect 22176 196 22236 362
rect 23190 196 23250 362
rect 23184 136 23190 196
rect 23250 136 23256 196
rect 22176 130 22236 136
rect 23702 -60 23762 452
rect 24722 452 24728 992
rect 24762 992 24776 1028
rect 25738 1028 25798 1166
rect 26236 1118 26296 1276
rect 26584 1236 26810 1296
rect 27250 1276 27256 1336
rect 27316 1276 27322 1336
rect 26028 1112 26516 1118
rect 26028 1078 26040 1112
rect 26504 1078 26516 1112
rect 26028 1072 26516 1078
rect 24762 452 24768 992
rect 24722 440 24768 452
rect 25738 452 25746 1028
rect 25780 452 25798 1028
rect 26750 1028 26810 1236
rect 27256 1118 27316 1276
rect 27770 1226 27830 1684
rect 28790 1684 28800 1724
rect 28834 1724 28840 2260
rect 29808 2260 29868 2488
rect 30310 2350 30370 2828
rect 30822 2548 30882 2918
rect 31838 2918 31854 2962
rect 31888 2962 31894 3494
rect 32858 3460 32872 3494
rect 32860 3450 32872 3460
rect 31888 2918 31898 2962
rect 31118 2868 31606 2874
rect 31118 2834 31130 2868
rect 31594 2834 31606 2868
rect 31118 2828 31606 2834
rect 30816 2488 30822 2548
rect 30882 2488 30888 2548
rect 30816 2384 30822 2444
rect 30882 2384 30888 2444
rect 30100 2344 30588 2350
rect 30100 2310 30112 2344
rect 30576 2310 30588 2344
rect 30100 2304 30588 2310
rect 30318 2300 30378 2304
rect 29808 2194 29818 2260
rect 29812 1730 29818 2194
rect 28834 1684 28850 1724
rect 28064 1634 28552 1640
rect 28064 1600 28076 1634
rect 28540 1600 28552 1634
rect 28064 1594 28552 1600
rect 28282 1336 28342 1594
rect 28790 1442 28850 1684
rect 29802 1684 29818 1730
rect 29852 2194 29868 2260
rect 30822 2260 30882 2384
rect 31346 2350 31406 2828
rect 31838 2776 31898 2918
rect 32866 2918 32872 3450
rect 32906 3450 32920 3494
rect 33872 3494 33932 3762
rect 32906 2918 32912 3450
rect 33872 3440 33890 3494
rect 32866 2906 32912 2918
rect 33884 2918 33890 3440
rect 33924 3456 33936 3494
rect 33924 3440 33932 3456
rect 33924 2918 33930 3440
rect 33884 2906 33930 2918
rect 32136 2868 32624 2874
rect 32136 2834 32148 2868
rect 32612 2834 32624 2868
rect 32136 2828 32624 2834
rect 33154 2868 33642 2874
rect 33154 2834 33166 2868
rect 33630 2834 33642 2868
rect 33154 2828 33642 2834
rect 31832 2716 31838 2776
rect 31898 2716 31904 2776
rect 32358 2666 32418 2828
rect 33366 2666 33426 2828
rect 33984 2776 34044 8566
rect 34106 7652 34112 7712
rect 34172 7652 34178 7712
rect 34112 6154 34172 7652
rect 34228 7388 34288 8680
rect 34344 7430 34350 7490
rect 34410 7430 34416 7490
rect 34222 7328 34228 7388
rect 34288 7328 34294 7388
rect 34106 6094 34112 6154
rect 34172 6094 34178 6154
rect 34102 5192 34108 5252
rect 34168 5192 34174 5252
rect 34108 3928 34168 5192
rect 34228 4026 34288 7328
rect 34222 3966 34228 4026
rect 34288 3966 34294 4026
rect 34102 3868 34108 3928
rect 34168 3868 34174 3928
rect 33978 2716 33984 2776
rect 34044 2716 34050 2776
rect 32352 2606 32358 2666
rect 32418 2606 32424 2666
rect 33360 2606 33366 2666
rect 33426 2606 33432 2666
rect 34228 2550 34288 3966
rect 34350 3694 34410 7430
rect 34478 6262 34538 8784
rect 34476 6256 34538 6262
rect 34536 6196 34538 6256
rect 34476 6190 34538 6196
rect 34478 3822 34538 6190
rect 34472 3762 34478 3822
rect 34538 3762 34544 3822
rect 34344 3634 34350 3694
rect 34410 3634 34416 3694
rect 34600 2666 34660 13594
rect 34706 9784 34712 9844
rect 34772 9784 34778 9844
rect 34594 2606 34600 2666
rect 34660 2606 34666 2666
rect 31838 2488 31844 2548
rect 31904 2488 31910 2548
rect 32860 2490 34288 2550
rect 31118 2344 31606 2350
rect 31118 2310 31130 2344
rect 31594 2310 31606 2344
rect 31118 2304 31606 2310
rect 30822 2214 30836 2260
rect 29852 1730 29858 2194
rect 29852 1684 29862 1730
rect 29082 1634 29570 1640
rect 29082 1600 29094 1634
rect 29558 1600 29570 1634
rect 29082 1594 29570 1600
rect 28784 1382 28790 1442
rect 28850 1382 28856 1442
rect 29300 1336 29360 1594
rect 28276 1276 28282 1336
rect 28342 1276 28348 1336
rect 29294 1276 29300 1336
rect 29360 1276 29366 1336
rect 27764 1166 27770 1226
rect 27830 1166 27836 1226
rect 27046 1112 27534 1118
rect 27046 1078 27058 1112
rect 27522 1078 27534 1112
rect 27046 1072 27534 1078
rect 26750 992 26764 1028
rect 23992 402 24480 408
rect 23992 368 24004 402
rect 24468 368 24480 402
rect 23992 362 24480 368
rect 25010 402 25498 408
rect 25010 368 25022 402
rect 25486 368 25498 402
rect 25010 362 25498 368
rect 24206 196 24266 362
rect 25216 202 25276 362
rect 24206 130 24266 136
rect 25214 196 25276 202
rect 25274 190 25276 196
rect 25214 130 25274 136
rect 25738 -60 25798 452
rect 26758 452 26764 992
rect 26798 992 26810 1028
rect 27770 1028 27830 1166
rect 28282 1118 28342 1276
rect 29300 1118 29360 1276
rect 29802 1226 29862 1684
rect 30830 1684 30836 2214
rect 30870 2214 30882 2260
rect 31844 2260 31904 2488
rect 32136 2344 32624 2350
rect 32136 2310 32148 2344
rect 32612 2310 32624 2344
rect 32136 2304 32624 2310
rect 30870 1684 30876 2214
rect 31844 2200 31854 2260
rect 31848 1708 31854 2200
rect 30830 1672 30876 1684
rect 31842 1684 31854 1708
rect 31888 2200 31904 2260
rect 32860 2260 32920 2490
rect 33358 2350 33418 2490
rect 33154 2344 33642 2350
rect 33154 2310 33166 2344
rect 33630 2310 33642 2344
rect 33154 2304 33642 2310
rect 31888 1708 31894 2200
rect 31888 1684 31902 1708
rect 30100 1634 30588 1640
rect 30100 1600 30112 1634
rect 30576 1600 30588 1634
rect 30100 1594 30588 1600
rect 31118 1634 31606 1640
rect 31118 1600 31130 1634
rect 31594 1600 31606 1634
rect 31118 1594 31606 1600
rect 30314 1336 30374 1594
rect 30814 1382 30820 1442
rect 30880 1382 30886 1442
rect 30308 1276 30314 1336
rect 30374 1276 30380 1336
rect 29796 1166 29802 1226
rect 29862 1166 29868 1226
rect 28064 1112 28552 1118
rect 28064 1078 28076 1112
rect 28540 1078 28552 1112
rect 28064 1072 28552 1078
rect 29082 1112 29570 1118
rect 29082 1078 29094 1112
rect 29558 1078 29570 1112
rect 29082 1072 29570 1078
rect 26798 452 26804 992
rect 26758 440 26804 452
rect 27770 452 27782 1028
rect 27816 452 27830 1028
rect 28794 1028 28840 1040
rect 28794 504 28800 1028
rect 27254 408 27314 410
rect 26028 402 26516 408
rect 26028 368 26040 402
rect 26504 368 26516 402
rect 26028 362 26516 368
rect 27046 402 27534 408
rect 27046 368 27058 402
rect 27522 368 27534 402
rect 27046 362 27534 368
rect 26232 202 26292 362
rect 26230 196 26292 202
rect 26290 190 26292 196
rect 27254 196 27314 362
rect 26230 130 26290 136
rect 27254 130 27314 136
rect 27770 -60 27830 452
rect 28784 452 28800 504
rect 28834 504 28840 1028
rect 29802 1028 29862 1166
rect 30314 1118 30374 1276
rect 30100 1112 30588 1118
rect 30100 1078 30112 1112
rect 30576 1078 30588 1112
rect 30100 1072 30588 1078
rect 28834 452 28844 504
rect 28064 402 28552 408
rect 28064 368 28076 402
rect 28540 368 28552 402
rect 28064 362 28552 368
rect 28276 196 28336 362
rect 28784 304 28844 452
rect 29802 452 29818 1028
rect 29852 452 29862 1028
rect 30820 1028 30880 1382
rect 31328 1336 31388 1594
rect 31322 1276 31328 1336
rect 31388 1276 31394 1336
rect 31328 1118 31388 1276
rect 31842 1226 31902 1684
rect 32860 1684 32872 2260
rect 32906 1684 32920 2260
rect 33874 2260 33934 2490
rect 33998 2384 34004 2444
rect 34064 2384 34070 2444
rect 33874 2206 33890 2260
rect 32136 1634 32624 1640
rect 32136 1600 32148 1634
rect 32612 1600 32624 1634
rect 32136 1594 32624 1600
rect 32350 1336 32410 1594
rect 32860 1548 32920 1684
rect 33884 1684 33890 2206
rect 33924 2206 33934 2260
rect 33924 1684 33930 2206
rect 33884 1672 33930 1684
rect 33154 1634 33642 1640
rect 33154 1600 33166 1634
rect 33630 1600 33642 1634
rect 33154 1594 33642 1600
rect 32854 1488 32860 1548
rect 32920 1488 32926 1548
rect 32854 1382 32860 1442
rect 32920 1382 32926 1442
rect 32344 1276 32350 1336
rect 32410 1276 32416 1336
rect 31836 1166 31842 1226
rect 31902 1166 31908 1226
rect 31118 1112 31606 1118
rect 31118 1078 31130 1112
rect 31594 1078 31606 1112
rect 31118 1072 31606 1078
rect 30820 984 30836 1028
rect 29082 402 29570 408
rect 29082 368 29094 402
rect 29558 368 29570 402
rect 29082 362 29570 368
rect 28778 244 28784 304
rect 28844 244 28850 304
rect 29296 202 29356 362
rect 29296 196 29358 202
rect 29296 190 29298 196
rect 28276 130 28336 136
rect 29298 130 29358 136
rect 29802 -60 29862 452
rect 30830 452 30836 984
rect 30870 984 30880 1028
rect 31842 1028 31902 1166
rect 32350 1118 32410 1276
rect 32860 1226 32920 1382
rect 32860 1166 33938 1226
rect 32136 1112 32624 1118
rect 32136 1078 32148 1112
rect 32612 1078 32624 1112
rect 32136 1072 32624 1078
rect 30870 452 30876 984
rect 30830 440 30876 452
rect 31842 452 31854 1028
rect 31888 452 31902 1028
rect 32860 1028 32920 1166
rect 33376 1118 33436 1166
rect 33154 1112 33642 1118
rect 33154 1078 33166 1112
rect 33630 1078 33642 1112
rect 33154 1072 33642 1078
rect 32860 1020 32872 1028
rect 30318 408 30378 410
rect 30100 402 30588 408
rect 30100 368 30112 402
rect 30576 368 30588 402
rect 30100 362 30588 368
rect 31118 402 31606 408
rect 31118 368 31130 402
rect 31594 368 31606 402
rect 31118 362 31606 368
rect 30318 202 30378 362
rect 31332 202 31392 362
rect 30316 196 30378 202
rect 30376 190 30378 196
rect 31330 196 31392 202
rect 30316 130 30376 136
rect 31390 190 31392 196
rect 31330 130 31390 136
rect 31842 -60 31902 452
rect 32866 452 32872 1020
rect 32906 1020 32920 1028
rect 33878 1028 33938 1166
rect 32906 452 32912 1020
rect 33878 1010 33890 1028
rect 32866 440 32912 452
rect 33884 452 33890 1010
rect 33924 1010 33938 1028
rect 33924 452 33930 1010
rect 33884 440 33930 452
rect 32352 408 32412 410
rect 32136 402 32624 408
rect 32136 368 32148 402
rect 32612 368 32624 402
rect 32136 362 32624 368
rect 33154 402 33642 408
rect 33154 368 33166 402
rect 33630 368 33642 402
rect 33154 362 33642 368
rect 32352 202 32412 362
rect 34004 304 34064 2384
rect 34712 1442 34772 9784
rect 34706 1382 34712 1442
rect 34772 1382 34778 1442
rect 33998 244 34004 304
rect 34064 244 34070 304
rect 32352 196 32414 202
rect 32352 190 32354 196
rect 32354 130 32414 136
rect 35766 40 35772 14300
rect 35872 40 35878 14300
rect 39622 14300 39734 15070
rect 53838 15012 53898 15018
rect 54160 14962 54166 15022
rect 54226 14962 54232 15022
rect 54286 15014 54346 15020
rect 53226 14816 53232 14876
rect 53292 14816 53298 14876
rect 53346 14818 53352 14878
rect 53412 14818 53418 14878
rect 53486 14836 53492 14896
rect 53552 14836 53558 14896
rect 53714 14852 53720 14912
rect 53780 14852 53786 14912
rect 53094 14688 53100 14748
rect 53160 14688 53166 14748
rect 36712 13970 38688 13976
rect 36712 13870 36818 13970
rect 38582 13870 38688 13970
rect 36712 13864 38688 13870
rect 36712 13803 36824 13864
rect 36712 12593 36718 13803
rect 36818 12593 36824 13803
rect 37424 13564 37434 13864
rect 37966 13564 37976 13864
rect 38576 13803 38688 13864
rect 36890 13396 38514 13426
rect 36890 13300 36928 13396
rect 38480 13300 38514 13396
rect 36890 13272 38514 13300
rect 36900 13130 37084 13272
rect 36900 12986 36960 13130
rect 37024 13085 37084 13130
rect 37002 13079 37110 13085
rect 37002 13045 37014 13079
rect 37098 13045 37110 13079
rect 37002 13039 37110 13045
rect 37260 13079 37368 13085
rect 37260 13045 37272 13079
rect 37356 13045 37368 13079
rect 37260 13039 37368 13045
rect 36900 12810 36910 12986
rect 36944 12810 36960 12986
rect 37162 12986 37208 12998
rect 37162 12876 37168 12986
rect 36900 12658 36960 12810
rect 37156 12810 37168 12876
rect 37202 12876 37208 12986
rect 37414 12986 37474 13272
rect 37666 13134 37672 13194
rect 37732 13134 37738 13194
rect 37518 13079 37626 13085
rect 37518 13045 37530 13079
rect 37614 13045 37626 13079
rect 37518 13039 37626 13045
rect 37414 12936 37426 12986
rect 37202 12810 37216 12876
rect 37002 12751 37110 12757
rect 37002 12717 37014 12751
rect 37098 12717 37110 12751
rect 37002 12711 37110 12717
rect 37028 12658 37088 12711
rect 37156 12660 37216 12810
rect 37420 12810 37426 12936
rect 37460 12936 37474 12986
rect 37672 12986 37732 13134
rect 37776 13079 37884 13085
rect 37776 13045 37788 13079
rect 37872 13045 37884 13079
rect 37776 13039 37884 13045
rect 37460 12810 37466 12936
rect 37420 12798 37466 12810
rect 37672 12810 37684 12986
rect 37718 12810 37732 12986
rect 37930 12986 37990 13272
rect 38316 13135 38502 13272
rect 38316 13085 38376 13135
rect 38034 13079 38142 13085
rect 38034 13045 38046 13079
rect 38130 13045 38142 13079
rect 38034 13039 38142 13045
rect 38292 13079 38400 13085
rect 38292 13045 38304 13079
rect 38388 13045 38400 13079
rect 38292 13039 38400 13045
rect 37930 12938 37942 12986
rect 37260 12751 37368 12757
rect 37260 12717 37272 12751
rect 37356 12717 37368 12751
rect 37260 12711 37368 12717
rect 37518 12751 37626 12757
rect 37518 12717 37530 12751
rect 37614 12717 37626 12751
rect 37518 12711 37626 12717
rect 37284 12662 37344 12711
rect 37540 12662 37600 12711
rect 37672 12662 37732 12810
rect 37936 12810 37942 12938
rect 37976 12938 37990 12986
rect 38194 12986 38240 12998
rect 37976 12810 37982 12938
rect 38194 12844 38200 12986
rect 37936 12798 37982 12810
rect 38186 12810 38200 12844
rect 38234 12844 38240 12986
rect 38442 12986 38502 13135
rect 38234 12810 38246 12844
rect 37776 12751 37884 12757
rect 37776 12717 37788 12751
rect 37872 12717 37884 12751
rect 37776 12711 37884 12717
rect 38034 12751 38142 12757
rect 38034 12717 38046 12751
rect 38130 12717 38142 12751
rect 38034 12711 38142 12717
rect 37802 12662 37862 12711
rect 38058 12662 38118 12711
rect 36900 12598 37088 12658
rect 37150 12600 37156 12660
rect 37216 12600 37222 12660
rect 37284 12602 38118 12662
rect 38186 12660 38246 12810
rect 38442 12810 38458 12986
rect 38492 12810 38502 12986
rect 38292 12751 38400 12757
rect 38292 12717 38304 12751
rect 38388 12717 38400 12751
rect 38292 12711 38400 12717
rect 38314 12660 38374 12711
rect 38442 12660 38502 12810
rect 38180 12600 38186 12660
rect 38246 12600 38252 12660
rect 38314 12600 38502 12660
rect 36712 12532 36824 12593
rect 38576 12593 38582 13803
rect 38682 12593 38688 13803
rect 38576 12532 38688 12593
rect 36712 12526 38688 12532
rect 36712 12426 36818 12526
rect 38582 12426 38688 12526
rect 36712 12420 38688 12426
rect -836 -76 -808 -68
rect -1378 -142 -1198 -76
rect -814 -142 -808 -76
rect -1378 -152 -808 -142
rect 2832 -106 2982 -60
rect 3028 -106 6202 -60
rect 6262 -106 12654 -60
rect 12714 -106 34756 -60
rect 34816 -106 34918 -60
rect -1378 -154 -1140 -152
rect -894 -154 -810 -152
rect -1378 -746 -1266 -154
rect 2832 -260 2878 -106
rect 34878 -260 34918 -106
rect 2832 -306 34918 -260
rect -666 -746 -656 -446
rect 35156 -746 35166 -446
rect 35766 -746 35878 40
rect -1378 -752 35878 -746
rect -1378 -852 -1272 -752
rect 35772 -852 35878 -752
rect -1378 -858 35878 -852
rect 39622 40 39628 14300
rect 39728 40 39734 14300
rect 50382 14090 50388 14150
rect 50448 14090 50454 14150
rect 50388 14046 50448 14090
rect 42754 13986 50448 14046
rect 42754 13846 42814 13986
rect 43264 13936 43324 13986
rect 43048 13930 43536 13936
rect 43048 13896 43060 13930
rect 43524 13896 43536 13930
rect 43048 13890 43536 13896
rect 42754 13816 42766 13846
rect 42760 13288 42766 13816
rect 42750 13270 42766 13288
rect 42800 13816 42814 13846
rect 43770 13846 43830 13986
rect 44272 13936 44332 13986
rect 45300 13936 45360 13986
rect 44066 13930 44554 13936
rect 44066 13896 44078 13930
rect 44542 13896 44554 13930
rect 44066 13890 44554 13896
rect 45084 13930 45572 13936
rect 45084 13896 45096 13930
rect 45560 13896 45572 13930
rect 45084 13890 45572 13896
rect 43770 13822 43784 13846
rect 42800 13288 42806 13816
rect 43778 13292 43784 13822
rect 42800 13270 42810 13288
rect 42750 13028 42810 13270
rect 43770 13270 43784 13292
rect 43818 13822 43830 13846
rect 44796 13846 44842 13858
rect 43818 13292 43824 13822
rect 44796 13294 44802 13846
rect 43818 13270 43830 13292
rect 43048 13220 43536 13226
rect 43048 13186 43060 13220
rect 43524 13186 43536 13220
rect 43048 13180 43536 13186
rect 43264 13118 43324 13180
rect 43048 13112 43536 13118
rect 43048 13078 43060 13112
rect 43524 13078 43536 13112
rect 43048 13072 43536 13078
rect 42750 12998 42766 13028
rect 42760 12474 42766 12998
rect 42752 12452 42766 12474
rect 42800 12998 42810 13028
rect 43770 13028 43830 13270
rect 44790 13270 44802 13294
rect 44836 13294 44842 13846
rect 45808 13846 45868 13986
rect 46314 13936 46374 13986
rect 47328 13936 47388 13986
rect 46102 13930 46590 13936
rect 46102 13896 46114 13930
rect 46578 13896 46590 13930
rect 46102 13890 46590 13896
rect 47120 13930 47608 13936
rect 47120 13896 47132 13930
rect 47596 13896 47608 13930
rect 47120 13890 47608 13896
rect 45808 13808 45820 13846
rect 44836 13270 44850 13294
rect 45814 13290 45820 13808
rect 44066 13220 44554 13226
rect 44066 13186 44078 13220
rect 44542 13186 44554 13220
rect 44066 13180 44554 13186
rect 44268 13118 44328 13180
rect 44066 13112 44554 13118
rect 44066 13078 44078 13112
rect 44542 13078 44554 13112
rect 44066 13072 44554 13078
rect 43770 13002 43784 13028
rect 42800 12474 42806 12998
rect 43778 12478 43784 13002
rect 42800 12452 42812 12474
rect 42752 12210 42812 12452
rect 43772 12452 43784 12478
rect 43818 13002 43830 13028
rect 44790 13028 44850 13270
rect 45808 13270 45820 13290
rect 45854 13808 45868 13846
rect 46832 13846 46878 13858
rect 47844 13846 47904 13986
rect 48360 13936 48420 13986
rect 49366 13936 49426 13986
rect 48138 13930 48626 13936
rect 48138 13896 48150 13930
rect 48614 13896 48626 13930
rect 48138 13890 48626 13896
rect 49156 13930 49644 13936
rect 49156 13896 49168 13930
rect 49632 13896 49644 13930
rect 49156 13890 49644 13896
rect 45854 13290 45860 13808
rect 46832 13298 46838 13846
rect 45854 13270 45868 13290
rect 45084 13220 45572 13226
rect 45084 13186 45096 13220
rect 45560 13186 45572 13220
rect 45084 13180 45572 13186
rect 45298 13118 45358 13180
rect 45084 13112 45572 13118
rect 45084 13078 45096 13112
rect 45560 13078 45572 13112
rect 45084 13072 45572 13078
rect 44790 13004 44802 13028
rect 43818 12478 43824 13002
rect 44796 12480 44802 13004
rect 43818 12452 43832 12478
rect 43048 12402 43536 12408
rect 43048 12368 43060 12402
rect 43524 12368 43536 12402
rect 43048 12362 43536 12368
rect 43264 12300 43324 12362
rect 43048 12294 43536 12300
rect 43048 12260 43060 12294
rect 43524 12260 43536 12294
rect 43048 12254 43536 12260
rect 42752 12184 42766 12210
rect 42760 11646 42766 12184
rect 42752 11634 42766 11646
rect 42800 12184 42812 12210
rect 43772 12210 43832 12452
rect 44792 12452 44802 12480
rect 44836 13004 44850 13028
rect 45808 13028 45868 13270
rect 46828 13270 46838 13298
rect 46872 13298 46878 13846
rect 47842 13812 47856 13846
rect 47844 13800 47856 13812
rect 46872 13270 46888 13298
rect 47850 13290 47856 13800
rect 46102 13220 46590 13226
rect 46102 13186 46114 13220
rect 46578 13186 46590 13220
rect 46102 13180 46590 13186
rect 46300 13118 46360 13180
rect 46102 13112 46590 13118
rect 46102 13078 46114 13112
rect 46578 13078 46590 13112
rect 46102 13072 46590 13078
rect 44836 12480 44842 13004
rect 45808 13000 45820 13028
rect 44836 12452 44852 12480
rect 45814 12476 45820 13000
rect 44066 12402 44554 12408
rect 44066 12368 44078 12402
rect 44542 12368 44554 12402
rect 44066 12362 44554 12368
rect 44280 12300 44340 12362
rect 44066 12294 44554 12300
rect 44066 12260 44078 12294
rect 44542 12260 44554 12294
rect 44066 12254 44554 12260
rect 43772 12188 43784 12210
rect 42800 11646 42806 12184
rect 43778 11650 43784 12188
rect 42800 11634 42812 11646
rect 42752 11392 42812 11634
rect 43772 11634 43784 11650
rect 43818 12188 43832 12210
rect 44792 12210 44852 12452
rect 45810 12452 45820 12476
rect 45854 13000 45868 13028
rect 46828 13028 46888 13270
rect 47840 13270 47856 13290
rect 47890 13800 47904 13846
rect 48868 13846 48914 13858
rect 47890 13290 47896 13800
rect 48868 13290 48874 13846
rect 47890 13270 47900 13290
rect 47120 13220 47608 13226
rect 47120 13186 47132 13220
rect 47596 13186 47608 13220
rect 47120 13180 47608 13186
rect 47330 13118 47390 13180
rect 47120 13112 47608 13118
rect 47120 13078 47132 13112
rect 47596 13078 47608 13112
rect 47120 13072 47608 13078
rect 46828 13008 46838 13028
rect 45854 12476 45860 13000
rect 46832 12484 46838 13008
rect 45854 12452 45870 12476
rect 45084 12402 45572 12408
rect 45084 12368 45096 12402
rect 45560 12368 45572 12402
rect 45084 12362 45572 12368
rect 45298 12300 45358 12362
rect 45084 12294 45572 12300
rect 45084 12260 45096 12294
rect 45560 12260 45572 12294
rect 45084 12254 45572 12260
rect 44792 12190 44802 12210
rect 43818 11650 43824 12188
rect 44796 11652 44802 12190
rect 43818 11634 43832 11650
rect 43048 11584 43536 11590
rect 43048 11550 43060 11584
rect 43524 11550 43536 11584
rect 43048 11544 43536 11550
rect 43258 11482 43318 11544
rect 43048 11476 43536 11482
rect 43048 11442 43060 11476
rect 43524 11442 43536 11476
rect 43048 11436 43536 11442
rect 42752 11356 42766 11392
rect 42760 10834 42766 11356
rect 42752 10816 42766 10834
rect 42800 11356 42812 11392
rect 43772 11392 43832 11634
rect 44792 11634 44802 11652
rect 44836 12190 44852 12210
rect 45810 12210 45870 12452
rect 46830 12452 46838 12484
rect 46872 13008 46888 13028
rect 47840 13028 47900 13270
rect 48862 13270 48874 13290
rect 48908 13290 48914 13846
rect 49878 13846 49938 13986
rect 50388 13936 50448 13986
rect 51908 13956 51914 14016
rect 51974 13956 51980 14016
rect 50174 13930 50662 13936
rect 50174 13896 50186 13930
rect 50650 13896 50662 13930
rect 50174 13890 50662 13896
rect 51192 13930 51680 13936
rect 51192 13896 51204 13930
rect 51668 13896 51680 13930
rect 51192 13890 51680 13896
rect 49878 13810 49892 13846
rect 49886 13290 49892 13810
rect 48908 13270 48922 13290
rect 48138 13220 48626 13226
rect 48138 13186 48150 13220
rect 48614 13186 48626 13220
rect 48138 13180 48626 13186
rect 48346 13118 48406 13180
rect 48138 13112 48626 13118
rect 48138 13078 48150 13112
rect 48614 13078 48626 13112
rect 48138 13072 48626 13078
rect 46872 12484 46878 13008
rect 47840 13000 47856 13028
rect 46872 12452 46890 12484
rect 47850 12476 47856 13000
rect 46102 12402 46590 12408
rect 46102 12368 46114 12402
rect 46578 12368 46590 12402
rect 46102 12362 46590 12368
rect 46300 12300 46360 12362
rect 46102 12294 46590 12300
rect 46102 12260 46114 12294
rect 46578 12260 46590 12294
rect 46102 12254 46590 12260
rect 44836 11652 44842 12190
rect 45810 12186 45820 12210
rect 44836 11634 44852 11652
rect 45814 11648 45820 12186
rect 44066 11584 44554 11590
rect 44066 11550 44078 11584
rect 44542 11550 44554 11584
rect 44066 11544 44554 11550
rect 44280 11482 44340 11544
rect 44066 11476 44554 11482
rect 44066 11442 44078 11476
rect 44542 11442 44554 11476
rect 44066 11436 44554 11442
rect 43772 11360 43784 11392
rect 42800 10834 42806 11356
rect 43778 10838 43784 11360
rect 42800 10816 42812 10834
rect 42752 10574 42812 10816
rect 43772 10816 43784 10838
rect 43818 11360 43832 11392
rect 44792 11392 44852 11634
rect 45810 11634 45820 11648
rect 45854 12186 45870 12210
rect 46830 12210 46890 12452
rect 47842 12452 47856 12476
rect 47890 13000 47900 13028
rect 48862 13028 48922 13270
rect 49882 13270 49892 13290
rect 49926 13810 49938 13846
rect 50904 13846 50950 13858
rect 49926 13290 49932 13810
rect 50904 13294 50910 13846
rect 49926 13270 49942 13290
rect 49156 13220 49644 13226
rect 49156 13186 49168 13220
rect 49632 13186 49644 13220
rect 49156 13180 49644 13186
rect 49368 13118 49428 13180
rect 49156 13112 49644 13118
rect 49156 13078 49168 13112
rect 49632 13078 49644 13112
rect 49156 13072 49644 13078
rect 48862 13000 48874 13028
rect 47890 12476 47896 13000
rect 48868 12476 48874 13000
rect 47890 12452 47902 12476
rect 47120 12402 47608 12408
rect 47120 12368 47132 12402
rect 47596 12368 47608 12402
rect 47120 12362 47608 12368
rect 47330 12300 47390 12362
rect 47120 12294 47608 12300
rect 47120 12260 47132 12294
rect 47596 12260 47608 12294
rect 47120 12254 47608 12260
rect 46830 12194 46838 12210
rect 45854 11648 45860 12186
rect 46832 11656 46838 12194
rect 45854 11634 45870 11648
rect 45084 11584 45572 11590
rect 45084 11550 45096 11584
rect 45560 11550 45572 11584
rect 45084 11544 45572 11550
rect 45292 11482 45352 11544
rect 45084 11476 45572 11482
rect 45084 11442 45096 11476
rect 45560 11442 45572 11476
rect 45084 11436 45572 11442
rect 44792 11362 44802 11392
rect 43818 10838 43824 11360
rect 44796 10840 44802 11362
rect 43818 10816 43832 10838
rect 43048 10766 43536 10772
rect 43048 10732 43060 10766
rect 43524 10732 43536 10766
rect 43048 10726 43536 10732
rect 43256 10664 43316 10726
rect 43048 10658 43536 10664
rect 43048 10624 43060 10658
rect 43524 10624 43536 10658
rect 43048 10618 43536 10624
rect 42752 10544 42766 10574
rect 42760 10014 42766 10544
rect 42752 9998 42766 10014
rect 42800 10544 42812 10574
rect 43772 10574 43832 10816
rect 44792 10816 44802 10840
rect 44836 11362 44852 11392
rect 45810 11392 45870 11634
rect 46830 11634 46838 11656
rect 46872 12194 46890 12210
rect 47842 12210 47902 12452
rect 48864 12452 48874 12476
rect 48908 13000 48922 13028
rect 49882 13028 49942 13270
rect 50898 13270 50910 13294
rect 50944 13294 50950 13846
rect 51914 13846 51974 13956
rect 51914 13810 51928 13846
rect 50944 13270 50958 13294
rect 51922 13290 51928 13810
rect 50174 13220 50662 13226
rect 50174 13186 50186 13220
rect 50650 13186 50662 13220
rect 50174 13180 50662 13186
rect 50380 13118 50440 13180
rect 50174 13112 50662 13118
rect 50174 13078 50186 13112
rect 50650 13078 50662 13112
rect 50174 13072 50662 13078
rect 49882 13000 49892 13028
rect 48908 12476 48914 13000
rect 49886 12476 49892 13000
rect 48908 12452 48924 12476
rect 48138 12402 48626 12408
rect 48138 12368 48150 12402
rect 48614 12368 48626 12402
rect 48138 12362 48626 12368
rect 48346 12300 48406 12362
rect 48138 12294 48626 12300
rect 48138 12260 48150 12294
rect 48614 12260 48626 12294
rect 48138 12254 48626 12260
rect 46872 11656 46878 12194
rect 47842 12186 47856 12210
rect 46872 11634 46890 11656
rect 47850 11648 47856 12186
rect 46102 11584 46590 11590
rect 46102 11550 46114 11584
rect 46578 11550 46590 11584
rect 46102 11544 46590 11550
rect 46294 11482 46354 11544
rect 46102 11476 46590 11482
rect 46102 11442 46114 11476
rect 46578 11442 46590 11476
rect 46102 11436 46590 11442
rect 44836 10840 44842 11362
rect 45810 11358 45820 11392
rect 44836 10816 44852 10840
rect 45814 10836 45820 11358
rect 44066 10766 44554 10772
rect 44066 10732 44078 10766
rect 44542 10732 44554 10766
rect 44066 10726 44554 10732
rect 44274 10664 44334 10726
rect 44066 10658 44554 10664
rect 44066 10624 44078 10658
rect 44542 10624 44554 10658
rect 44066 10618 44554 10624
rect 43772 10548 43784 10574
rect 42800 10014 42806 10544
rect 43778 10018 43784 10548
rect 42800 9998 42812 10014
rect 42752 9756 42812 9998
rect 43772 9998 43784 10018
rect 43818 10548 43832 10574
rect 44792 10574 44852 10816
rect 45810 10816 45820 10836
rect 45854 11358 45870 11392
rect 46830 11392 46890 11634
rect 47842 11634 47856 11648
rect 47890 12186 47902 12210
rect 48864 12210 48924 12452
rect 49884 12452 49892 12476
rect 49926 13000 49942 13028
rect 50898 13028 50958 13270
rect 51920 13270 51928 13290
rect 51962 13810 51974 13846
rect 51962 13290 51968 13810
rect 51962 13270 51980 13290
rect 51192 13220 51680 13226
rect 51192 13186 51204 13220
rect 51668 13186 51680 13220
rect 51192 13180 51680 13186
rect 51400 13118 51460 13180
rect 51192 13112 51680 13118
rect 51192 13078 51204 13112
rect 51668 13078 51680 13112
rect 51192 13072 51680 13078
rect 50898 13004 50910 13028
rect 49926 12476 49932 13000
rect 50904 12480 50910 13004
rect 49926 12452 49944 12476
rect 49156 12402 49644 12408
rect 49156 12368 49168 12402
rect 49632 12368 49644 12402
rect 49156 12362 49644 12368
rect 49368 12300 49428 12362
rect 49156 12294 49644 12300
rect 49156 12260 49168 12294
rect 49632 12260 49644 12294
rect 49156 12254 49644 12260
rect 48864 12186 48874 12210
rect 47890 11648 47896 12186
rect 48868 11648 48874 12186
rect 47890 11634 47902 11648
rect 47120 11584 47608 11590
rect 47120 11550 47132 11584
rect 47596 11550 47608 11584
rect 47120 11544 47608 11550
rect 47324 11482 47384 11544
rect 47120 11476 47608 11482
rect 47120 11442 47132 11476
rect 47596 11442 47608 11476
rect 47120 11436 47608 11442
rect 46830 11366 46838 11392
rect 45854 10836 45860 11358
rect 46832 10844 46838 11366
rect 45854 10816 45870 10836
rect 45084 10766 45572 10772
rect 45084 10732 45096 10766
rect 45560 10732 45572 10766
rect 45084 10726 45572 10732
rect 45290 10664 45350 10726
rect 45084 10658 45572 10664
rect 45084 10624 45096 10658
rect 45560 10624 45572 10658
rect 45084 10618 45572 10624
rect 44792 10550 44802 10574
rect 43818 10018 43824 10548
rect 44796 10020 44802 10550
rect 43818 9998 43832 10018
rect 43048 9948 43536 9954
rect 43048 9914 43060 9948
rect 43524 9914 43536 9948
rect 43048 9908 43536 9914
rect 43258 9846 43318 9908
rect 43048 9840 43536 9846
rect 43048 9806 43060 9840
rect 43524 9806 43536 9840
rect 43048 9800 43536 9806
rect 42752 9724 42766 9756
rect 42760 9202 42766 9724
rect 42752 9180 42766 9202
rect 42800 9724 42812 9756
rect 43772 9756 43832 9998
rect 44792 9998 44802 10020
rect 44836 10550 44852 10574
rect 45810 10574 45870 10816
rect 46830 10816 46838 10844
rect 46872 11366 46890 11392
rect 47842 11392 47902 11634
rect 48864 11634 48874 11648
rect 48908 12186 48924 12210
rect 49884 12210 49944 12452
rect 50900 12452 50910 12480
rect 50944 13004 50958 13028
rect 51920 13028 51980 13270
rect 50944 12480 50950 13004
rect 51920 13000 51928 13028
rect 50944 12452 50960 12480
rect 50174 12402 50662 12408
rect 50174 12368 50186 12402
rect 50650 12368 50662 12402
rect 50174 12362 50662 12368
rect 50380 12300 50440 12362
rect 50174 12294 50662 12300
rect 50174 12260 50186 12294
rect 50650 12260 50662 12294
rect 50174 12254 50662 12260
rect 49884 12186 49892 12210
rect 48908 11648 48914 12186
rect 49886 11648 49892 12186
rect 48908 11634 48924 11648
rect 48138 11584 48626 11590
rect 48138 11550 48150 11584
rect 48614 11550 48626 11584
rect 48138 11544 48626 11550
rect 48340 11482 48400 11544
rect 48138 11476 48626 11482
rect 48138 11442 48150 11476
rect 48614 11442 48626 11476
rect 48138 11436 48626 11442
rect 46872 10844 46878 11366
rect 47842 11358 47856 11392
rect 46872 10816 46890 10844
rect 47850 10836 47856 11358
rect 46102 10766 46590 10772
rect 46102 10732 46114 10766
rect 46578 10732 46590 10766
rect 46102 10726 46590 10732
rect 46292 10664 46352 10726
rect 46102 10658 46590 10664
rect 46102 10624 46114 10658
rect 46578 10624 46590 10658
rect 46102 10618 46590 10624
rect 44836 10020 44842 10550
rect 45810 10546 45820 10574
rect 44836 9998 44852 10020
rect 45814 10016 45820 10546
rect 44066 9948 44554 9954
rect 44066 9914 44078 9948
rect 44542 9914 44554 9948
rect 44066 9908 44554 9914
rect 44272 9846 44332 9908
rect 44066 9840 44554 9846
rect 44066 9806 44078 9840
rect 44542 9806 44554 9840
rect 44066 9800 44554 9806
rect 43772 9728 43784 9756
rect 42800 9202 42806 9724
rect 43778 9206 43784 9728
rect 42800 9180 42812 9202
rect 42752 8938 42812 9180
rect 43772 9180 43784 9206
rect 43818 9728 43832 9756
rect 44792 9756 44852 9998
rect 45810 9998 45820 10016
rect 45854 10546 45870 10574
rect 46830 10574 46890 10816
rect 47842 10816 47856 10836
rect 47890 11358 47902 11392
rect 48864 11392 48924 11634
rect 49884 11634 49892 11648
rect 49926 12186 49944 12210
rect 50900 12210 50960 12452
rect 51922 12452 51928 13000
rect 51962 13000 51980 13028
rect 51962 12476 51968 13000
rect 51962 12452 51982 12476
rect 51192 12402 51680 12408
rect 51192 12368 51204 12402
rect 51668 12368 51680 12402
rect 51192 12362 51680 12368
rect 51400 12300 51460 12362
rect 51192 12294 51680 12300
rect 51192 12260 51204 12294
rect 51668 12260 51680 12294
rect 51192 12254 51680 12260
rect 50900 12190 50910 12210
rect 49926 11648 49932 12186
rect 50904 11652 50910 12190
rect 49926 11634 49944 11648
rect 49156 11584 49644 11590
rect 49156 11550 49168 11584
rect 49632 11550 49644 11584
rect 49156 11544 49644 11550
rect 49362 11482 49422 11544
rect 49156 11476 49644 11482
rect 49156 11442 49168 11476
rect 49632 11442 49644 11476
rect 49156 11436 49644 11442
rect 48864 11358 48874 11392
rect 47890 10836 47896 11358
rect 48868 10836 48874 11358
rect 47890 10816 47902 10836
rect 47120 10766 47608 10772
rect 47120 10732 47132 10766
rect 47596 10732 47608 10766
rect 47120 10726 47608 10732
rect 47322 10664 47382 10726
rect 47120 10658 47608 10664
rect 47120 10624 47132 10658
rect 47596 10624 47608 10658
rect 47120 10618 47608 10624
rect 46830 10554 46838 10574
rect 45854 10016 45860 10546
rect 46832 10024 46838 10554
rect 45854 9998 45870 10016
rect 45084 9948 45572 9954
rect 45084 9914 45096 9948
rect 45560 9914 45572 9948
rect 45084 9908 45572 9914
rect 45292 9846 45352 9908
rect 45084 9840 45572 9846
rect 45084 9806 45096 9840
rect 45560 9806 45572 9840
rect 45084 9800 45572 9806
rect 44792 9730 44802 9756
rect 43818 9206 43824 9728
rect 44796 9208 44802 9730
rect 43818 9180 43832 9206
rect 43048 9130 43536 9136
rect 43048 9096 43060 9130
rect 43524 9096 43536 9130
rect 43048 9090 43536 9096
rect 43260 9028 43320 9090
rect 43048 9022 43536 9028
rect 43048 8988 43060 9022
rect 43524 8988 43536 9022
rect 43048 8982 43536 8988
rect 42752 8912 42766 8938
rect 42760 8384 42766 8912
rect 42752 8362 42766 8384
rect 42800 8912 42812 8938
rect 43772 8938 43832 9180
rect 44792 9180 44802 9208
rect 44836 9730 44852 9756
rect 45810 9756 45870 9998
rect 46830 9998 46838 10024
rect 46872 10554 46890 10574
rect 47842 10574 47902 10816
rect 48864 10816 48874 10836
rect 48908 11358 48924 11392
rect 49884 11392 49944 11634
rect 50900 11634 50910 11652
rect 50944 12190 50960 12210
rect 51922 12210 51982 12452
rect 50944 11652 50950 12190
rect 50944 11634 50960 11652
rect 50174 11584 50662 11590
rect 50174 11550 50186 11584
rect 50650 11550 50662 11584
rect 50174 11544 50662 11550
rect 50374 11482 50434 11544
rect 50174 11476 50662 11482
rect 50174 11442 50186 11476
rect 50650 11442 50662 11476
rect 50174 11436 50662 11442
rect 49884 11358 49892 11392
rect 48908 10836 48914 11358
rect 49886 10836 49892 11358
rect 48908 10816 48924 10836
rect 48138 10766 48626 10772
rect 48138 10732 48150 10766
rect 48614 10732 48626 10766
rect 48138 10726 48626 10732
rect 48338 10664 48398 10726
rect 48138 10658 48626 10664
rect 48138 10624 48150 10658
rect 48614 10624 48626 10658
rect 48138 10618 48626 10624
rect 46872 10024 46878 10554
rect 47842 10546 47856 10574
rect 46872 9998 46890 10024
rect 47850 10016 47856 10546
rect 46102 9948 46590 9954
rect 46102 9914 46114 9948
rect 46578 9914 46590 9948
rect 46102 9908 46590 9914
rect 46294 9846 46354 9908
rect 46102 9840 46590 9846
rect 46102 9806 46114 9840
rect 46578 9806 46590 9840
rect 46102 9800 46590 9806
rect 44836 9208 44842 9730
rect 45810 9726 45820 9756
rect 44836 9180 44852 9208
rect 45814 9204 45820 9726
rect 44066 9130 44554 9136
rect 44066 9096 44078 9130
rect 44542 9096 44554 9130
rect 44066 9090 44554 9096
rect 44274 9028 44334 9090
rect 44066 9022 44554 9028
rect 44066 8988 44078 9022
rect 44542 8988 44554 9022
rect 44066 8982 44554 8988
rect 43772 8916 43784 8938
rect 42800 8384 42806 8912
rect 43778 8388 43784 8916
rect 42800 8362 42812 8384
rect 42752 8120 42812 8362
rect 43772 8362 43784 8388
rect 43818 8916 43832 8938
rect 44792 8938 44852 9180
rect 45810 9180 45820 9204
rect 45854 9726 45870 9756
rect 46830 9756 46890 9998
rect 47842 9998 47856 10016
rect 47890 10546 47902 10574
rect 48864 10574 48924 10816
rect 49884 10816 49892 10836
rect 49926 11358 49944 11392
rect 50900 11392 50960 11634
rect 51922 11634 51928 12210
rect 51962 12186 51982 12210
rect 51962 11648 51968 12186
rect 51962 11634 51982 11648
rect 51192 11584 51680 11590
rect 51192 11550 51204 11584
rect 51668 11550 51680 11584
rect 51192 11544 51680 11550
rect 51394 11482 51454 11544
rect 51192 11476 51680 11482
rect 51192 11442 51204 11476
rect 51668 11442 51680 11476
rect 51192 11436 51680 11442
rect 50900 11362 50910 11392
rect 49926 10836 49932 11358
rect 50904 10840 50910 11362
rect 49926 10816 49944 10836
rect 49156 10766 49644 10772
rect 49156 10732 49168 10766
rect 49632 10732 49644 10766
rect 49156 10726 49644 10732
rect 49360 10664 49420 10726
rect 49156 10658 49644 10664
rect 49156 10624 49168 10658
rect 49632 10624 49644 10658
rect 49156 10618 49644 10624
rect 48864 10546 48874 10574
rect 47890 10016 47896 10546
rect 48868 10016 48874 10546
rect 47890 9998 47902 10016
rect 47120 9948 47608 9954
rect 47120 9914 47132 9948
rect 47596 9914 47608 9948
rect 47120 9908 47608 9914
rect 47324 9846 47384 9908
rect 47120 9840 47608 9846
rect 47120 9806 47132 9840
rect 47596 9806 47608 9840
rect 47120 9800 47608 9806
rect 46830 9734 46838 9756
rect 45854 9204 45860 9726
rect 46832 9212 46838 9734
rect 45854 9180 45870 9204
rect 45084 9130 45572 9136
rect 45084 9096 45096 9130
rect 45560 9096 45572 9130
rect 45084 9090 45572 9096
rect 45294 9028 45354 9090
rect 45084 9022 45572 9028
rect 45084 8988 45096 9022
rect 45560 8988 45572 9022
rect 45084 8982 45572 8988
rect 44792 8918 44802 8938
rect 43818 8388 43824 8916
rect 44796 8390 44802 8918
rect 43818 8362 43832 8388
rect 43048 8312 43536 8318
rect 43048 8278 43060 8312
rect 43524 8278 43536 8312
rect 43048 8272 43536 8278
rect 43262 8210 43322 8272
rect 43048 8204 43536 8210
rect 43048 8170 43060 8204
rect 43524 8170 43536 8204
rect 43048 8164 43536 8170
rect 42752 8094 42766 8120
rect 42760 7544 42766 8094
rect 42800 8094 42812 8120
rect 43772 8120 43832 8362
rect 44792 8362 44802 8390
rect 44836 8918 44852 8938
rect 45810 8938 45870 9180
rect 46830 9180 46838 9212
rect 46872 9734 46890 9756
rect 47842 9756 47902 9998
rect 48864 9998 48874 10016
rect 48908 10546 48924 10574
rect 49884 10574 49944 10816
rect 50900 10816 50910 10840
rect 50944 11362 50960 11392
rect 51922 11392 51982 11634
rect 50944 10840 50950 11362
rect 50944 10816 50960 10840
rect 50174 10766 50662 10772
rect 50174 10732 50186 10766
rect 50650 10732 50662 10766
rect 50174 10726 50662 10732
rect 50372 10664 50432 10726
rect 50174 10658 50662 10664
rect 50174 10624 50186 10658
rect 50650 10624 50662 10658
rect 50174 10618 50662 10624
rect 49884 10546 49892 10574
rect 48908 10016 48914 10546
rect 49886 10016 49892 10546
rect 48908 9998 48924 10016
rect 48138 9948 48626 9954
rect 48138 9914 48150 9948
rect 48614 9914 48626 9948
rect 48138 9908 48626 9914
rect 48340 9846 48400 9908
rect 48138 9840 48626 9846
rect 48138 9806 48150 9840
rect 48614 9806 48626 9840
rect 48138 9800 48626 9806
rect 46872 9212 46878 9734
rect 47842 9726 47856 9756
rect 46872 9180 46890 9212
rect 47850 9204 47856 9726
rect 46102 9130 46590 9136
rect 46102 9096 46114 9130
rect 46578 9096 46590 9130
rect 46102 9090 46590 9096
rect 46296 9028 46356 9090
rect 46102 9022 46590 9028
rect 46102 8988 46114 9022
rect 46578 8988 46590 9022
rect 46102 8982 46590 8988
rect 44836 8390 44842 8918
rect 45810 8914 45820 8938
rect 44836 8362 44852 8390
rect 45814 8386 45820 8914
rect 44066 8312 44554 8318
rect 44066 8278 44078 8312
rect 44542 8278 44554 8312
rect 44066 8272 44554 8278
rect 44276 8210 44336 8272
rect 44066 8204 44554 8210
rect 44066 8170 44078 8204
rect 44542 8170 44554 8204
rect 44066 8164 44554 8170
rect 43772 8098 43784 8120
rect 42800 7544 42806 8094
rect 42760 7532 42806 7544
rect 43778 7544 43784 8098
rect 43818 8098 43832 8120
rect 44792 8120 44852 8362
rect 45810 8362 45820 8386
rect 45854 8914 45870 8938
rect 46830 8938 46890 9180
rect 47842 9180 47856 9204
rect 47890 9726 47902 9756
rect 48864 9756 48924 9998
rect 49884 9998 49892 10016
rect 49926 10546 49944 10574
rect 50900 10574 50960 10816
rect 51922 10816 51928 11392
rect 51962 11358 51982 11392
rect 51962 10836 51968 11358
rect 51962 10816 51982 10836
rect 51192 10766 51680 10772
rect 51192 10732 51204 10766
rect 51668 10732 51680 10766
rect 51192 10726 51680 10732
rect 51392 10664 51452 10726
rect 51192 10658 51680 10664
rect 51192 10624 51204 10658
rect 51668 10624 51680 10658
rect 51192 10618 51680 10624
rect 50900 10550 50910 10574
rect 49926 10016 49932 10546
rect 50904 10020 50910 10550
rect 49926 9998 49944 10016
rect 49156 9948 49644 9954
rect 49156 9914 49168 9948
rect 49632 9914 49644 9948
rect 49156 9908 49644 9914
rect 49362 9846 49422 9908
rect 49156 9840 49644 9846
rect 49156 9806 49168 9840
rect 49632 9806 49644 9840
rect 49156 9800 49644 9806
rect 48864 9726 48874 9756
rect 47890 9204 47896 9726
rect 48868 9204 48874 9726
rect 47890 9180 47902 9204
rect 47120 9130 47608 9136
rect 47120 9096 47132 9130
rect 47596 9096 47608 9130
rect 47120 9090 47608 9096
rect 47326 9028 47386 9090
rect 47120 9022 47608 9028
rect 47120 8988 47132 9022
rect 47596 8988 47608 9022
rect 47120 8982 47608 8988
rect 46830 8922 46838 8938
rect 45854 8386 45860 8914
rect 46832 8394 46838 8922
rect 45854 8362 45870 8386
rect 45084 8312 45572 8318
rect 45084 8278 45096 8312
rect 45560 8278 45572 8312
rect 45084 8272 45572 8278
rect 45296 8210 45356 8272
rect 45084 8204 45572 8210
rect 45084 8170 45096 8204
rect 45560 8170 45572 8204
rect 45084 8164 45572 8170
rect 44792 8100 44802 8120
rect 43818 7544 43824 8098
rect 44796 7590 44802 8100
rect 43778 7532 43824 7544
rect 44786 7544 44802 7590
rect 44836 8100 44852 8120
rect 45810 8120 45870 8362
rect 46830 8362 46838 8394
rect 46872 8922 46890 8938
rect 47842 8938 47902 9180
rect 48864 9180 48874 9204
rect 48908 9726 48924 9756
rect 49884 9756 49944 9998
rect 50900 9998 50910 10020
rect 50944 10550 50960 10574
rect 51922 10574 51982 10816
rect 50944 10020 50950 10550
rect 50944 9998 50960 10020
rect 50174 9948 50662 9954
rect 50174 9914 50186 9948
rect 50650 9914 50662 9948
rect 50174 9908 50662 9914
rect 50374 9846 50434 9908
rect 50174 9840 50662 9846
rect 50174 9806 50186 9840
rect 50650 9806 50662 9840
rect 50174 9800 50662 9806
rect 49884 9726 49892 9756
rect 48908 9204 48914 9726
rect 49886 9204 49892 9726
rect 48908 9180 48924 9204
rect 48138 9130 48626 9136
rect 48138 9096 48150 9130
rect 48614 9096 48626 9130
rect 48138 9090 48626 9096
rect 48342 9028 48402 9090
rect 48138 9022 48626 9028
rect 48138 8988 48150 9022
rect 48614 8988 48626 9022
rect 48138 8982 48626 8988
rect 46872 8394 46878 8922
rect 47842 8914 47856 8938
rect 46872 8362 46890 8394
rect 47850 8386 47856 8914
rect 46102 8312 46590 8318
rect 46102 8278 46114 8312
rect 46578 8278 46590 8312
rect 46102 8272 46590 8278
rect 46298 8210 46358 8272
rect 46102 8204 46590 8210
rect 46102 8170 46114 8204
rect 46578 8170 46590 8204
rect 46102 8164 46590 8170
rect 44836 7590 44842 8100
rect 45810 8096 45820 8120
rect 44836 7544 44846 7590
rect 43048 7494 43536 7500
rect 43048 7460 43060 7494
rect 43524 7460 43536 7494
rect 43048 7454 43536 7460
rect 44066 7494 44554 7500
rect 44066 7460 44078 7494
rect 44542 7460 44554 7494
rect 44066 7454 44554 7460
rect 44786 7370 44846 7544
rect 45814 7544 45820 8096
rect 45854 8096 45870 8120
rect 46830 8120 46890 8362
rect 47842 8362 47856 8386
rect 47890 8914 47902 8938
rect 48864 8938 48924 9180
rect 49884 9180 49892 9204
rect 49926 9726 49944 9756
rect 50900 9756 50960 9998
rect 51922 9998 51928 10574
rect 51962 10546 51982 10574
rect 51962 10016 51968 10546
rect 51962 9998 51982 10016
rect 51192 9948 51680 9954
rect 51192 9914 51204 9948
rect 51668 9914 51680 9948
rect 51192 9908 51680 9914
rect 51394 9846 51454 9908
rect 51192 9840 51680 9846
rect 51192 9806 51204 9840
rect 51668 9806 51680 9840
rect 51192 9800 51680 9806
rect 50900 9730 50910 9756
rect 49926 9204 49932 9726
rect 50904 9208 50910 9730
rect 49926 9180 49944 9204
rect 49156 9130 49644 9136
rect 49156 9096 49168 9130
rect 49632 9096 49644 9130
rect 49156 9090 49644 9096
rect 49364 9028 49424 9090
rect 49156 9022 49644 9028
rect 49156 8988 49168 9022
rect 49632 8988 49644 9022
rect 49156 8982 49644 8988
rect 48864 8914 48874 8938
rect 47890 8386 47896 8914
rect 48868 8386 48874 8914
rect 47890 8362 47902 8386
rect 47120 8312 47608 8318
rect 47120 8278 47132 8312
rect 47596 8278 47608 8312
rect 47120 8272 47608 8278
rect 47328 8210 47388 8272
rect 47120 8204 47608 8210
rect 47120 8170 47132 8204
rect 47596 8170 47608 8204
rect 47120 8164 47608 8170
rect 46830 8104 46838 8120
rect 45854 7544 45860 8096
rect 46832 7592 46838 8104
rect 45814 7532 45860 7544
rect 46824 7544 46838 7592
rect 46872 8104 46890 8120
rect 47842 8120 47902 8362
rect 48864 8362 48874 8386
rect 48908 8914 48924 8938
rect 49884 8938 49944 9180
rect 50900 9180 50910 9208
rect 50944 9730 50960 9756
rect 51922 9756 51982 9998
rect 50944 9208 50950 9730
rect 50944 9180 50960 9208
rect 50174 9130 50662 9136
rect 50174 9096 50186 9130
rect 50650 9096 50662 9130
rect 50174 9090 50662 9096
rect 50376 9028 50436 9090
rect 50174 9022 50662 9028
rect 50174 8988 50186 9022
rect 50650 8988 50662 9022
rect 50174 8982 50662 8988
rect 49884 8914 49892 8938
rect 48908 8386 48914 8914
rect 49886 8386 49892 8914
rect 48908 8362 48924 8386
rect 48138 8312 48626 8318
rect 48138 8278 48150 8312
rect 48614 8278 48626 8312
rect 48138 8272 48626 8278
rect 48344 8210 48404 8272
rect 48138 8204 48626 8210
rect 48138 8170 48150 8204
rect 48614 8170 48626 8204
rect 48138 8164 48626 8170
rect 46872 7592 46878 8104
rect 47842 8096 47856 8120
rect 46872 7544 46884 7592
rect 45084 7494 45572 7500
rect 45084 7460 45096 7494
rect 45560 7460 45572 7494
rect 45084 7454 45572 7460
rect 46102 7494 46590 7500
rect 46102 7460 46114 7494
rect 46578 7460 46590 7494
rect 46102 7454 46590 7460
rect 46824 7370 46884 7544
rect 47850 7544 47856 8096
rect 47890 8096 47902 8120
rect 48864 8120 48924 8362
rect 49884 8362 49892 8386
rect 49926 8914 49944 8938
rect 50900 8938 50960 9180
rect 51922 9180 51928 9756
rect 51962 9726 51982 9756
rect 51962 9204 51968 9726
rect 51962 9180 51982 9204
rect 51192 9130 51680 9136
rect 51192 9096 51204 9130
rect 51668 9096 51680 9130
rect 51192 9090 51680 9096
rect 51396 9028 51456 9090
rect 51192 9022 51680 9028
rect 51192 8988 51204 9022
rect 51668 8988 51680 9022
rect 51192 8982 51680 8988
rect 50900 8918 50910 8938
rect 49926 8386 49932 8914
rect 50904 8390 50910 8918
rect 49926 8362 49944 8386
rect 49156 8312 49644 8318
rect 49156 8278 49168 8312
rect 49632 8278 49644 8312
rect 49156 8272 49644 8278
rect 49366 8210 49426 8272
rect 49156 8204 49644 8210
rect 49156 8170 49168 8204
rect 49632 8170 49644 8204
rect 49156 8164 49644 8170
rect 48864 8096 48874 8120
rect 47890 7544 47896 8096
rect 48868 7588 48874 8096
rect 47850 7532 47896 7544
rect 48860 7544 48874 7588
rect 48908 8096 48924 8120
rect 49884 8120 49944 8362
rect 50900 8362 50910 8390
rect 50944 8918 50960 8938
rect 51922 8938 51982 9180
rect 50944 8390 50950 8918
rect 50944 8362 50960 8390
rect 50174 8312 50662 8318
rect 50174 8278 50186 8312
rect 50650 8278 50662 8312
rect 50174 8272 50662 8278
rect 50378 8210 50438 8272
rect 50174 8204 50662 8210
rect 50174 8170 50186 8204
rect 50650 8170 50662 8204
rect 50174 8164 50662 8170
rect 49884 8096 49892 8120
rect 48908 7588 48914 8096
rect 48908 7544 48920 7588
rect 47120 7494 47608 7500
rect 47120 7460 47132 7494
rect 47596 7460 47608 7494
rect 47120 7454 47608 7460
rect 48138 7494 48626 7500
rect 48138 7460 48150 7494
rect 48614 7460 48626 7494
rect 48138 7454 48626 7460
rect 48860 7370 48920 7544
rect 49886 7544 49892 8096
rect 49926 8096 49944 8120
rect 50900 8120 50960 8362
rect 51922 8362 51928 8938
rect 51962 8914 51982 8938
rect 51962 8386 51968 8914
rect 51962 8362 51982 8386
rect 51192 8312 51680 8318
rect 51192 8278 51204 8312
rect 51668 8278 51680 8312
rect 51192 8272 51680 8278
rect 51398 8210 51458 8272
rect 51192 8204 51680 8210
rect 51192 8170 51204 8204
rect 51668 8170 51680 8204
rect 51192 8164 51680 8170
rect 50900 8100 50910 8120
rect 49926 7544 49932 8096
rect 50904 7586 50910 8100
rect 49886 7532 49932 7544
rect 50896 7544 50910 7586
rect 50944 8100 50960 8120
rect 51922 8120 51982 8362
rect 50944 7586 50950 8100
rect 51922 7598 51928 8120
rect 50944 7544 50956 7586
rect 49156 7494 49644 7500
rect 49156 7460 49168 7494
rect 49632 7460 49644 7494
rect 49156 7454 49644 7460
rect 50174 7494 50662 7500
rect 50174 7460 50186 7494
rect 50650 7460 50662 7494
rect 50174 7454 50662 7460
rect 50896 7370 50956 7544
rect 51916 7544 51928 7598
rect 51962 8096 51982 8120
rect 51962 7598 51968 8096
rect 51962 7544 51976 7598
rect 53100 7548 53160 14688
rect 51192 7494 51680 7500
rect 51192 7460 51204 7494
rect 51668 7460 51680 7494
rect 51192 7454 51680 7460
rect 51410 7370 51470 7454
rect 51916 7370 51976 7544
rect 53094 7488 53100 7548
rect 53160 7488 53166 7548
rect 44786 7310 53080 7370
rect 48546 6562 48552 6622
rect 48612 6562 48618 6622
rect 42442 6476 42502 6482
rect 46516 6416 46522 6476
rect 46582 6416 46588 6476
rect 41282 6288 41288 6348
rect 41348 6288 41354 6348
rect 41288 5252 41348 6288
rect 42442 6284 42502 6416
rect 43960 6288 43966 6348
rect 44026 6288 44032 6348
rect 44992 6288 44998 6348
rect 45058 6288 45064 6348
rect 41426 6224 42502 6284
rect 41426 6096 41486 6224
rect 41934 6186 41994 6224
rect 41724 6180 42212 6186
rect 41724 6146 41736 6180
rect 42200 6146 42212 6180
rect 41724 6140 42212 6146
rect 41426 6050 41442 6096
rect 41436 5520 41442 6050
rect 41476 6050 41486 6096
rect 42442 6096 42502 6224
rect 43966 6186 44026 6288
rect 44998 6186 45058 6288
rect 42742 6180 43230 6186
rect 42742 6146 42754 6180
rect 43218 6146 43230 6180
rect 42742 6140 43230 6146
rect 43760 6180 44248 6186
rect 43760 6146 43772 6180
rect 44236 6146 44248 6180
rect 43760 6140 44248 6146
rect 44778 6180 45266 6186
rect 44778 6146 44790 6180
rect 45254 6146 45266 6180
rect 44778 6140 45266 6146
rect 45796 6180 46284 6186
rect 45796 6146 45808 6180
rect 46272 6146 46284 6180
rect 45796 6140 46284 6146
rect 42442 6056 42460 6096
rect 41476 5520 41482 6050
rect 41436 5508 41482 5520
rect 42454 5520 42460 6056
rect 42494 6056 42502 6096
rect 43472 6096 43518 6108
rect 42494 5520 42500 6056
rect 43472 5584 43478 6096
rect 42454 5508 42500 5520
rect 43464 5520 43478 5584
rect 43512 5584 43518 6096
rect 44490 6096 44536 6108
rect 43512 5520 43524 5584
rect 44490 5566 44496 6096
rect 41724 5470 42212 5476
rect 41724 5436 41736 5470
rect 42200 5436 42212 5470
rect 41724 5430 42212 5436
rect 42742 5470 43230 5476
rect 42742 5436 42754 5470
rect 43218 5436 43230 5470
rect 42742 5430 43230 5436
rect 42946 5386 43006 5430
rect 42940 5326 42946 5386
rect 43006 5326 43012 5386
rect 42440 5222 42446 5282
rect 42506 5222 42512 5282
rect 41288 4116 41348 5192
rect 42446 5180 42506 5222
rect 41426 5120 42506 5180
rect 41426 4984 41486 5120
rect 41930 5074 41990 5120
rect 41724 5068 42212 5074
rect 41724 5034 41736 5068
rect 42200 5034 42212 5068
rect 41724 5028 42212 5034
rect 41426 4938 41442 4984
rect 41436 4408 41442 4938
rect 41476 4938 41486 4984
rect 42446 4984 42506 5120
rect 43464 5178 43524 5520
rect 44482 5520 44496 5566
rect 44530 5566 44536 6096
rect 45508 6096 45554 6108
rect 45508 5582 45514 6096
rect 44530 5520 44542 5566
rect 43760 5470 44248 5476
rect 43760 5436 43772 5470
rect 44236 5436 44248 5470
rect 43760 5430 44248 5436
rect 43964 5326 43970 5386
rect 44030 5326 44036 5386
rect 42742 5068 43230 5074
rect 42742 5034 42754 5068
rect 43218 5034 43230 5068
rect 42742 5028 43230 5034
rect 41476 4408 41482 4938
rect 41436 4396 41482 4408
rect 42446 4408 42460 4984
rect 42494 4408 42506 4984
rect 41724 4358 42212 4364
rect 41724 4324 41736 4358
rect 42200 4324 42212 4358
rect 41724 4318 42212 4324
rect 41282 4056 41288 4116
rect 41348 4056 41354 4116
rect 41288 1990 41348 4056
rect 41724 3956 42212 3962
rect 41724 3922 41736 3956
rect 42200 3922 42212 3956
rect 41724 3916 42212 3922
rect 41436 3872 41482 3884
rect 41436 3330 41442 3872
rect 41430 3296 41442 3330
rect 41476 3330 41482 3872
rect 42446 3872 42506 4408
rect 43464 4984 43524 5118
rect 43970 5074 44030 5326
rect 44482 5282 44542 5520
rect 45500 5520 45514 5582
rect 45548 5582 45554 6096
rect 46522 6096 46582 6416
rect 48052 6288 48058 6348
rect 48118 6288 48124 6348
rect 48058 6186 48118 6288
rect 46814 6180 47302 6186
rect 46814 6146 46826 6180
rect 47290 6146 47302 6180
rect 46814 6140 47302 6146
rect 47832 6180 48320 6186
rect 47832 6146 47844 6180
rect 48308 6146 48320 6180
rect 47832 6140 48320 6146
rect 46522 6032 46532 6096
rect 45548 5520 45560 5582
rect 44778 5470 45266 5476
rect 44778 5436 44790 5470
rect 45254 5436 45266 5470
rect 44778 5430 45266 5436
rect 44996 5326 45002 5386
rect 45062 5326 45068 5386
rect 44476 5222 44482 5282
rect 44542 5222 44548 5282
rect 45002 5074 45062 5326
rect 45500 5178 45560 5520
rect 46526 5520 46532 6032
rect 46566 6032 46582 6096
rect 47544 6096 47590 6108
rect 46566 5520 46572 6032
rect 47544 5592 47550 6096
rect 46526 5508 46572 5520
rect 47532 5520 47550 5592
rect 47584 5592 47590 6096
rect 48552 6096 48612 6562
rect 50576 6416 50582 6476
rect 50642 6416 50648 6476
rect 52760 6416 52766 6476
rect 52826 6416 52832 6476
rect 49048 6288 49054 6348
rect 49114 6288 49120 6348
rect 49054 6186 49114 6288
rect 48850 6180 49338 6186
rect 48850 6146 48862 6180
rect 49326 6146 49338 6180
rect 48850 6140 49338 6146
rect 49868 6180 50356 6186
rect 49868 6146 49880 6180
rect 50344 6146 50356 6180
rect 49868 6140 50356 6146
rect 49054 6138 49114 6140
rect 50582 6108 50642 6416
rect 50886 6180 51374 6186
rect 50886 6146 50898 6180
rect 51362 6146 51374 6180
rect 50886 6140 51374 6146
rect 51904 6180 52392 6186
rect 51904 6146 51916 6180
rect 52380 6146 52392 6180
rect 51904 6140 52392 6146
rect 47584 5520 47592 5592
rect 45796 5470 46284 5476
rect 45796 5436 45808 5470
rect 46272 5436 46284 5470
rect 45796 5430 46284 5436
rect 46814 5470 47302 5476
rect 46814 5436 46826 5470
rect 47290 5436 47302 5470
rect 46814 5430 47302 5436
rect 46002 5386 46062 5430
rect 47022 5386 47082 5430
rect 45996 5326 46002 5386
rect 46062 5326 46068 5386
rect 47016 5326 47022 5386
rect 47082 5326 47088 5386
rect 46512 5222 46518 5282
rect 46578 5222 46584 5282
rect 43760 5068 44248 5074
rect 43760 5034 43772 5068
rect 44236 5034 44248 5068
rect 43760 5028 44248 5034
rect 44778 5068 45266 5074
rect 44778 5034 44790 5068
rect 45254 5034 45266 5068
rect 44778 5028 45266 5034
rect 43464 4408 43478 4984
rect 43512 4408 43524 4984
rect 44490 4984 44536 4996
rect 44490 4446 44496 4984
rect 42742 4358 43230 4364
rect 42742 4324 42754 4358
rect 43218 4324 43230 4358
rect 42742 4318 43230 4324
rect 42938 4116 42998 4318
rect 42932 4056 42938 4116
rect 42998 4056 43004 4116
rect 42938 3962 42998 4056
rect 42742 3956 43230 3962
rect 42742 3922 42754 3956
rect 43218 3922 43230 3956
rect 42742 3916 43230 3922
rect 42446 3800 42460 3872
rect 41476 3296 41490 3330
rect 42454 3326 42460 3800
rect 41430 3164 41490 3296
rect 42450 3296 42460 3326
rect 42494 3800 42506 3872
rect 43464 3872 43524 4408
rect 44476 4408 44496 4446
rect 44530 4408 44536 4984
rect 43760 4358 44248 4364
rect 43760 4324 43772 4358
rect 44236 4324 44248 4358
rect 43760 4318 44248 4324
rect 44476 4236 44536 4408
rect 45500 4984 45560 5118
rect 45796 5068 46284 5074
rect 45796 5034 45808 5068
rect 46272 5034 46284 5068
rect 45796 5028 46284 5034
rect 45500 4408 45514 4984
rect 45548 4408 45560 4984
rect 44778 4358 45266 4364
rect 44778 4324 44790 4358
rect 45254 4324 45266 4358
rect 44778 4318 45266 4324
rect 44470 4176 44476 4236
rect 44536 4176 44542 4236
rect 43760 3956 44248 3962
rect 43760 3922 43772 3956
rect 44236 3922 44248 3956
rect 43760 3916 44248 3922
rect 42494 3326 42500 3800
rect 42494 3296 42510 3326
rect 41724 3246 42212 3252
rect 41724 3212 41736 3246
rect 42200 3212 42212 3246
rect 41724 3206 42212 3212
rect 41922 3164 41982 3206
rect 42450 3164 42510 3296
rect 43464 3296 43478 3872
rect 43512 3296 43524 3872
rect 44476 3872 44536 4176
rect 44778 3956 45266 3962
rect 44778 3922 44790 3956
rect 45254 3922 45266 3956
rect 44778 3916 45266 3922
rect 44476 3802 44496 3872
rect 42742 3246 43230 3252
rect 42742 3212 42754 3246
rect 43218 3212 43230 3246
rect 42742 3206 43230 3212
rect 41430 3104 42510 3164
rect 42450 3064 42510 3104
rect 43464 3172 43524 3296
rect 44490 3296 44496 3802
rect 44530 3296 44536 3872
rect 44490 3284 44536 3296
rect 45500 3872 45560 4408
rect 46518 4984 46578 5222
rect 47532 5178 47592 5520
rect 48552 5520 48568 6096
rect 48602 5520 48612 6096
rect 49580 6096 49626 6108
rect 49580 5582 49586 6096
rect 47832 5470 48320 5476
rect 47832 5436 47844 5470
rect 48308 5436 48320 5470
rect 47832 5430 48320 5436
rect 48036 5326 48042 5386
rect 48102 5326 48108 5386
rect 47526 5118 47532 5178
rect 47592 5118 47598 5178
rect 46814 5068 47302 5074
rect 46814 5034 46826 5068
rect 47290 5034 47302 5068
rect 46814 5028 47302 5034
rect 46518 4408 46532 4984
rect 46566 4408 46578 4984
rect 45796 4358 46284 4364
rect 45796 4324 45808 4358
rect 46272 4324 46284 4358
rect 45796 4318 46284 4324
rect 46008 4116 46068 4318
rect 46002 4056 46008 4116
rect 46068 4056 46074 4116
rect 46008 3962 46068 4056
rect 45796 3956 46284 3962
rect 45796 3922 45808 3956
rect 46272 3922 46284 3956
rect 45796 3916 46284 3922
rect 45500 3296 45514 3872
rect 45548 3296 45560 3872
rect 46518 3872 46578 4408
rect 47532 4984 47592 5118
rect 48042 5074 48102 5326
rect 48552 5282 48612 5520
rect 49566 5520 49586 5582
rect 49620 5520 49626 6096
rect 50582 6096 50644 6108
rect 50582 6064 50604 6096
rect 48850 5470 49338 5476
rect 48850 5436 48862 5470
rect 49326 5436 49338 5470
rect 48850 5430 49338 5436
rect 49052 5386 49112 5392
rect 48546 5222 48552 5282
rect 48612 5222 48618 5282
rect 49052 5074 49112 5326
rect 49566 5178 49626 5520
rect 50598 5520 50604 6064
rect 50638 5520 50644 6096
rect 51616 6096 51662 6108
rect 51616 5554 51622 6096
rect 50598 5508 50644 5520
rect 51610 5520 51622 5554
rect 51656 5554 51662 6096
rect 52634 6096 52680 6108
rect 52634 5574 52640 6096
rect 51656 5520 51670 5554
rect 49868 5470 50356 5476
rect 49868 5436 49880 5470
rect 50344 5436 50356 5470
rect 49868 5430 50356 5436
rect 50886 5470 51374 5476
rect 50886 5436 50898 5470
rect 51362 5436 51374 5470
rect 50886 5430 51374 5436
rect 50066 5386 50126 5430
rect 51084 5386 51144 5430
rect 50060 5326 50066 5386
rect 50126 5326 50132 5386
rect 51084 5320 51144 5326
rect 51610 5292 51670 5520
rect 52626 5520 52640 5574
rect 52674 5574 52680 6096
rect 52674 5520 52686 5574
rect 51904 5470 52392 5476
rect 51904 5436 51916 5470
rect 52380 5436 52392 5470
rect 51904 5430 52392 5436
rect 52114 5292 52174 5430
rect 52626 5292 52686 5520
rect 50582 5222 50588 5282
rect 50648 5222 50654 5282
rect 51610 5232 52686 5292
rect 47832 5068 48320 5074
rect 47832 5034 47844 5068
rect 48308 5034 48320 5068
rect 47832 5028 48320 5034
rect 48850 5068 49338 5074
rect 48850 5034 48862 5068
rect 49326 5034 49338 5068
rect 48850 5028 49338 5034
rect 47532 4408 47550 4984
rect 47584 4408 47592 4984
rect 48562 4984 48608 4996
rect 48562 4464 48568 4984
rect 46814 4358 47302 4364
rect 46814 4324 46826 4358
rect 47290 4324 47302 4358
rect 46814 4318 47302 4324
rect 47016 4116 47076 4318
rect 47010 4056 47016 4116
rect 47076 4056 47082 4116
rect 47016 3962 47076 4056
rect 46814 3956 47302 3962
rect 46814 3922 46826 3956
rect 47290 3922 47302 3956
rect 46814 3916 47302 3922
rect 46518 3766 46532 3872
rect 46526 3358 46532 3766
rect 43760 3246 44248 3252
rect 43760 3212 43772 3246
rect 44236 3212 44248 3246
rect 43760 3206 44248 3212
rect 44778 3246 45266 3252
rect 44778 3212 44790 3246
rect 45254 3212 45266 3246
rect 44778 3206 45266 3212
rect 42444 3004 42450 3064
rect 42510 3004 42516 3064
rect 42938 2892 42944 2952
rect 43004 2892 43010 2952
rect 42944 2850 43004 2892
rect 41724 2844 42212 2850
rect 41724 2810 41736 2844
rect 42200 2810 42212 2844
rect 41724 2804 42212 2810
rect 42742 2844 43230 2850
rect 42742 2810 42754 2844
rect 43218 2810 43230 2844
rect 42742 2804 43230 2810
rect 41436 2760 41482 2772
rect 41436 2226 41442 2760
rect 41426 2184 41442 2226
rect 41476 2226 41482 2760
rect 42454 2760 42500 2772
rect 41476 2184 41486 2226
rect 42454 2220 42460 2760
rect 41426 2040 41486 2184
rect 42444 2184 42460 2220
rect 42494 2220 42500 2760
rect 43464 2760 43524 3112
rect 43968 2952 44028 3206
rect 44480 3004 44486 3064
rect 44546 3004 44552 3064
rect 43962 2892 43968 2952
rect 44028 2892 44034 2952
rect 43760 2844 44248 2850
rect 43760 2810 43772 2844
rect 44236 2810 44248 2844
rect 43760 2804 44248 2810
rect 43464 2658 43478 2760
rect 42494 2184 42504 2220
rect 41724 2134 42212 2140
rect 41724 2100 41736 2134
rect 42200 2100 42212 2134
rect 41724 2094 42212 2100
rect 41930 2040 41990 2094
rect 42444 2040 42504 2184
rect 43472 2184 43478 2658
rect 43512 2658 43524 2760
rect 44486 2760 44546 3004
rect 45000 2952 45060 3206
rect 45500 3172 45560 3296
rect 46522 3296 46532 3358
rect 46566 3766 46578 3872
rect 47532 3872 47592 4408
rect 48552 4408 48568 4464
rect 48602 4464 48608 4984
rect 49566 4984 49626 5118
rect 49868 5068 50356 5074
rect 49868 5034 49880 5068
rect 50344 5034 50356 5068
rect 49868 5028 50356 5034
rect 48602 4408 48612 4464
rect 47832 4358 48320 4364
rect 47832 4324 47844 4358
rect 48308 4324 48320 4358
rect 47832 4318 48320 4324
rect 48552 4236 48612 4408
rect 49566 4408 49586 4984
rect 49620 4408 49626 4984
rect 48850 4358 49338 4364
rect 48850 4324 48862 4358
rect 49326 4324 49338 4358
rect 48850 4318 49338 4324
rect 48546 4176 48552 4236
rect 48612 4176 48618 4236
rect 47832 3956 48320 3962
rect 47832 3922 47844 3956
rect 48308 3922 48320 3956
rect 47832 3916 48320 3922
rect 46566 3358 46572 3766
rect 46566 3296 46582 3358
rect 45796 3246 46284 3252
rect 45796 3212 45808 3246
rect 46272 3212 46284 3246
rect 45796 3206 46284 3212
rect 44994 2892 45000 2952
rect 45060 2892 45066 2952
rect 44778 2844 45266 2850
rect 44778 2810 44790 2844
rect 45254 2810 45266 2844
rect 44778 2804 45266 2810
rect 44486 2720 44496 2760
rect 43512 2184 43518 2658
rect 43472 2172 43518 2184
rect 44490 2184 44496 2720
rect 44530 2720 44546 2760
rect 45500 2760 45560 3112
rect 46522 3064 46582 3296
rect 47532 3296 47550 3872
rect 47584 3296 47592 3872
rect 48552 3872 48612 4176
rect 48850 3956 49338 3962
rect 48850 3922 48862 3956
rect 49326 3922 49338 3956
rect 48850 3916 49338 3922
rect 48552 3830 48568 3872
rect 46814 3246 47302 3252
rect 46814 3212 46826 3246
rect 47290 3212 47302 3246
rect 46814 3206 47302 3212
rect 47532 3172 47592 3296
rect 48562 3296 48568 3830
rect 48602 3830 48612 3872
rect 49566 3872 49626 4408
rect 50588 4984 50648 5222
rect 51610 5178 51670 5232
rect 50886 5068 51374 5074
rect 50886 5034 50898 5068
rect 51362 5034 51374 5068
rect 50886 5028 51374 5034
rect 50588 4408 50604 4984
rect 50638 4408 50648 4984
rect 49868 4358 50356 4364
rect 49868 4324 49880 4358
rect 50344 4324 50356 4358
rect 49868 4318 50356 4324
rect 50078 4116 50138 4318
rect 50072 4056 50078 4116
rect 50138 4056 50144 4116
rect 50078 3962 50138 4056
rect 49868 3956 50356 3962
rect 49868 3922 49880 3956
rect 50344 3922 50356 3956
rect 49868 3916 50356 3922
rect 48602 3296 48608 3830
rect 48562 3284 48608 3296
rect 49566 3296 49586 3872
rect 49620 3296 49626 3872
rect 50588 3872 50648 4408
rect 51610 4984 51670 5118
rect 52114 5074 52174 5232
rect 51904 5068 52392 5074
rect 51904 5034 51916 5068
rect 52380 5034 52392 5068
rect 51904 5028 52392 5034
rect 51610 4408 51622 4984
rect 51656 4408 51670 4984
rect 50886 4358 51374 4364
rect 50886 4324 50898 4358
rect 51362 4324 51374 4358
rect 50886 4318 51374 4324
rect 51104 4116 51164 4318
rect 51610 4172 51670 4408
rect 52626 4984 52686 5232
rect 52626 4408 52640 4984
rect 52674 4408 52686 4984
rect 51904 4358 52392 4364
rect 51904 4324 51916 4358
rect 52380 4324 52392 4358
rect 51904 4318 52392 4324
rect 52110 4172 52170 4318
rect 52626 4172 52686 4408
rect 52766 4236 52826 6416
rect 52880 5326 52886 5386
rect 52946 5326 52952 5386
rect 52760 4176 52766 4236
rect 52826 4176 52832 4236
rect 51098 4056 51104 4116
rect 51164 4056 51170 4116
rect 51610 4112 52686 4172
rect 51104 3962 51164 4056
rect 50886 3956 51374 3962
rect 50886 3922 50898 3956
rect 51362 3922 51374 3956
rect 50886 3916 51374 3922
rect 50588 3816 50604 3872
rect 50598 3342 50604 3816
rect 47832 3246 48320 3252
rect 47832 3212 47844 3246
rect 48308 3212 48320 3246
rect 47832 3206 48320 3212
rect 48850 3246 49338 3252
rect 48850 3212 48862 3246
rect 49326 3212 49338 3246
rect 48850 3206 49338 3212
rect 46516 3004 46522 3064
rect 46582 3004 46588 3064
rect 45994 2892 46000 2952
rect 46060 2892 46066 2952
rect 47014 2892 47020 2952
rect 47080 2892 47086 2952
rect 46000 2850 46060 2892
rect 47020 2850 47080 2892
rect 45796 2844 46284 2850
rect 45796 2810 45808 2844
rect 46272 2810 46284 2844
rect 45796 2804 46284 2810
rect 46814 2844 47302 2850
rect 46814 2810 46826 2844
rect 47290 2810 47302 2844
rect 46814 2804 47302 2810
rect 45500 2722 45514 2760
rect 44530 2184 44536 2720
rect 44490 2172 44536 2184
rect 45508 2184 45514 2722
rect 45548 2722 45560 2760
rect 46526 2760 46572 2772
rect 45548 2184 45554 2722
rect 46526 2244 46532 2760
rect 45508 2172 45554 2184
rect 46524 2184 46532 2244
rect 46566 2244 46572 2760
rect 47532 2760 47592 3112
rect 48040 2952 48100 3206
rect 48550 3004 48556 3064
rect 48616 3004 48622 3064
rect 48034 2892 48040 2952
rect 48100 2892 48106 2952
rect 47832 2844 48320 2850
rect 47832 2810 47844 2844
rect 48308 2810 48320 2844
rect 47832 2804 48320 2810
rect 47532 2700 47550 2760
rect 46566 2184 46584 2244
rect 42742 2134 43230 2140
rect 42742 2100 42754 2134
rect 43218 2100 43230 2134
rect 42742 2094 43230 2100
rect 43760 2134 44248 2140
rect 43760 2100 43772 2134
rect 44236 2100 44248 2134
rect 43760 2094 44248 2100
rect 44778 2134 45266 2140
rect 44778 2100 44790 2134
rect 45254 2100 45266 2134
rect 44778 2094 45266 2100
rect 45796 2134 46284 2140
rect 45796 2100 45808 2134
rect 46272 2100 46284 2134
rect 45796 2094 46284 2100
rect 41282 1930 41288 1990
rect 41348 1930 41354 1990
rect 41426 1980 42504 2040
rect 43958 1990 44018 2094
rect 44990 1990 45050 2094
rect 42444 1860 42504 1980
rect 43952 1930 43958 1990
rect 44018 1930 44024 1990
rect 44984 1930 44990 1990
rect 45050 1930 45056 1990
rect 46524 1860 46584 2184
rect 47544 2184 47550 2700
rect 47584 2700 47592 2760
rect 48556 2760 48616 3004
rect 49050 2952 49110 3206
rect 49050 2886 49110 2892
rect 49566 3172 49626 3296
rect 50592 3296 50604 3342
rect 50638 3816 50648 3872
rect 51610 3872 51670 4112
rect 52110 3962 52170 4112
rect 51904 3956 52392 3962
rect 51904 3922 51916 3956
rect 52380 3922 52392 3956
rect 51904 3916 52392 3922
rect 50638 3342 50644 3816
rect 50638 3296 50652 3342
rect 49868 3246 50356 3252
rect 49868 3212 49880 3246
rect 50344 3212 50356 3246
rect 49868 3206 50356 3212
rect 48850 2844 49338 2850
rect 48850 2810 48862 2844
rect 49326 2810 49338 2844
rect 48850 2804 49338 2810
rect 48556 2714 48568 2760
rect 47584 2184 47590 2700
rect 47544 2172 47590 2184
rect 48562 2184 48568 2714
rect 48602 2714 48616 2760
rect 49566 2760 49626 3112
rect 50592 3064 50652 3296
rect 51610 3296 51622 3872
rect 51656 3296 51670 3872
rect 50886 3246 51374 3252
rect 50886 3212 50898 3246
rect 51362 3212 51374 3246
rect 50886 3206 51374 3212
rect 51610 3172 51670 3296
rect 52626 3872 52686 4112
rect 52626 3296 52640 3872
rect 52674 3296 52686 3872
rect 51904 3246 52392 3252
rect 51904 3212 51916 3246
rect 52380 3212 52392 3246
rect 51904 3206 52392 3212
rect 51604 3112 51610 3172
rect 51670 3112 51676 3172
rect 50586 3004 50592 3064
rect 50652 3004 50658 3064
rect 51610 3060 51670 3112
rect 52118 3060 52178 3206
rect 52626 3060 52686 3296
rect 51610 3000 52686 3060
rect 51082 2952 51142 2958
rect 50058 2892 50064 2952
rect 50124 2892 50130 2952
rect 50064 2850 50124 2892
rect 51082 2850 51142 2892
rect 49868 2844 50356 2850
rect 49868 2810 49880 2844
rect 50344 2810 50356 2844
rect 49868 2804 50356 2810
rect 50886 2844 51374 2850
rect 50886 2810 50898 2844
rect 51362 2810 51374 2844
rect 50886 2804 51374 2810
rect 49566 2718 49586 2760
rect 48602 2184 48608 2714
rect 48562 2172 48608 2184
rect 49580 2184 49586 2718
rect 49620 2184 49626 2760
rect 50598 2760 50644 2772
rect 50598 2212 50604 2760
rect 49580 2172 49626 2184
rect 50584 2184 50604 2212
rect 50638 2184 50644 2760
rect 51610 2760 51670 3000
rect 52118 2850 52178 3000
rect 51904 2844 52392 2850
rect 51904 2810 51916 2844
rect 52380 2810 52392 2844
rect 51904 2804 52392 2810
rect 51610 2696 51622 2760
rect 46814 2134 47302 2140
rect 46814 2100 46826 2134
rect 47290 2100 47302 2134
rect 46814 2094 47302 2100
rect 47832 2134 48320 2140
rect 47832 2100 47844 2134
rect 48308 2100 48320 2134
rect 47832 2094 48320 2100
rect 48850 2134 49338 2140
rect 48850 2100 48862 2134
rect 49326 2100 49338 2134
rect 48850 2094 49338 2100
rect 49868 2134 50356 2140
rect 49868 2100 49880 2134
rect 50344 2100 50356 2134
rect 49868 2094 50356 2100
rect 48050 1990 48110 2094
rect 49046 1990 49106 2094
rect 48044 1930 48050 1990
rect 48110 1930 48116 1990
rect 49040 1930 49046 1990
rect 49106 1930 49112 1990
rect 50584 1860 50644 2184
rect 51616 2184 51622 2696
rect 51656 2696 51670 2760
rect 52626 2760 52686 3000
rect 52626 2718 52640 2760
rect 51656 2184 51662 2696
rect 51616 2172 51662 2184
rect 52634 2184 52640 2718
rect 52674 2718 52686 2760
rect 52674 2184 52680 2718
rect 52634 2172 52680 2184
rect 50886 2134 51374 2140
rect 50886 2100 50898 2134
rect 51362 2100 51374 2134
rect 50886 2094 51374 2100
rect 51904 2134 52392 2140
rect 51904 2100 51916 2134
rect 52380 2100 52392 2134
rect 51904 2094 52392 2100
rect 52766 1860 52826 4176
rect 52886 2952 52946 5326
rect 52880 2892 52886 2952
rect 52946 2892 52952 2952
rect 46518 1800 46524 1860
rect 46584 1800 46590 1860
rect 50578 1800 50584 1860
rect 50644 1800 50650 1860
rect 52760 1800 52766 1860
rect 52826 1800 52832 1860
rect 42444 1794 42504 1800
rect 41886 1394 52122 1454
rect 41886 1218 41946 1394
rect 42386 1308 42446 1394
rect 42182 1302 42670 1308
rect 42182 1268 42194 1302
rect 42658 1268 42670 1302
rect 42182 1262 42670 1268
rect 41886 1184 41900 1218
rect 41894 642 41900 1184
rect 41934 1184 41946 1218
rect 42908 1218 42968 1394
rect 43406 1308 43466 1394
rect 44440 1308 44500 1394
rect 45462 1308 45522 1394
rect 46452 1308 46512 1394
rect 43200 1302 43688 1308
rect 43200 1268 43212 1302
rect 43676 1268 43688 1302
rect 43200 1262 43688 1268
rect 44218 1302 44706 1308
rect 44218 1268 44230 1302
rect 44694 1268 44706 1302
rect 44218 1262 44706 1268
rect 45236 1302 45724 1308
rect 45236 1268 45248 1302
rect 45712 1268 45724 1302
rect 45236 1262 45724 1268
rect 46254 1302 46742 1308
rect 46254 1268 46266 1302
rect 46730 1268 46742 1302
rect 46254 1262 46742 1268
rect 41934 642 41940 1184
rect 42908 1174 42918 1218
rect 41894 630 41940 642
rect 42912 642 42918 1174
rect 42952 1174 42968 1218
rect 43930 1218 43976 1230
rect 42952 642 42958 1174
rect 43930 700 43936 1218
rect 42912 630 42958 642
rect 43922 642 43936 700
rect 43970 700 43976 1218
rect 44948 1218 44994 1230
rect 43970 642 43982 700
rect 44948 676 44954 1218
rect 42182 592 42670 598
rect 42182 558 42194 592
rect 42658 558 42670 592
rect 42182 552 42670 558
rect 43200 592 43688 598
rect 43200 558 43212 592
rect 43676 558 43688 592
rect 43200 552 43688 558
rect 43922 494 43982 642
rect 44940 642 44954 676
rect 44988 676 44994 1218
rect 45966 1218 46012 1230
rect 45966 688 45972 1218
rect 44988 642 45000 676
rect 44218 592 44706 598
rect 44218 558 44230 592
rect 44694 558 44706 592
rect 44218 552 44706 558
rect 43916 434 43922 494
rect 43982 434 43988 494
rect 39622 -746 39734 40
rect 43922 -60 43982 434
rect 44940 382 45000 642
rect 45960 642 45972 688
rect 46006 688 46012 1218
rect 46976 1218 47036 1394
rect 47486 1308 47546 1394
rect 48476 1308 48536 1394
rect 49508 1308 49568 1394
rect 50512 1308 50572 1394
rect 47272 1302 47760 1308
rect 47272 1268 47284 1302
rect 47748 1268 47760 1302
rect 47272 1262 47760 1268
rect 48290 1302 48778 1308
rect 48290 1268 48302 1302
rect 48766 1268 48778 1302
rect 48290 1262 48778 1268
rect 49308 1302 49796 1308
rect 49308 1268 49320 1302
rect 49784 1268 49796 1302
rect 49308 1262 49796 1268
rect 50326 1302 50814 1308
rect 50326 1268 50338 1302
rect 50802 1268 50814 1302
rect 50326 1262 50814 1268
rect 47486 1260 47546 1262
rect 49508 1260 49568 1262
rect 46976 1176 46990 1218
rect 46006 642 46020 688
rect 45236 592 45724 598
rect 45236 558 45248 592
rect 45712 558 45724 592
rect 45236 552 45724 558
rect 45960 494 46020 642
rect 46984 642 46990 1176
rect 47024 1176 47036 1218
rect 48002 1218 48048 1230
rect 47024 642 47030 1176
rect 48002 688 48008 1218
rect 46984 630 47030 642
rect 47996 642 48008 688
rect 48042 688 48048 1218
rect 49020 1218 49066 1230
rect 48042 642 48056 688
rect 49020 680 49026 1218
rect 46254 592 46742 598
rect 46254 558 46266 592
rect 46730 558 46742 592
rect 46254 552 46742 558
rect 47272 592 47760 598
rect 47272 558 47284 592
rect 47748 558 47760 592
rect 47272 552 47760 558
rect 47996 494 48056 642
rect 49014 642 49026 680
rect 49060 680 49066 1218
rect 50038 1218 50084 1230
rect 49060 642 49074 680
rect 50038 674 50044 1218
rect 48290 592 48778 598
rect 48290 558 48302 592
rect 48766 558 48778 592
rect 48290 552 48778 558
rect 45954 434 45960 494
rect 46020 434 46026 494
rect 47990 434 47996 494
rect 48056 434 48062 494
rect 44934 322 44940 382
rect 45000 322 45006 382
rect 45960 -60 46020 434
rect 47996 -60 48056 434
rect 49014 382 49074 642
rect 50032 642 50044 674
rect 50078 674 50084 1218
rect 51052 1218 51112 1394
rect 51532 1308 51592 1394
rect 51344 1302 51832 1308
rect 51344 1268 51356 1302
rect 51820 1268 51832 1302
rect 51344 1262 51832 1268
rect 51052 1150 51062 1218
rect 50078 642 50092 674
rect 49308 592 49796 598
rect 49308 558 49320 592
rect 49784 558 49796 592
rect 49308 552 49796 558
rect 50032 494 50092 642
rect 51056 642 51062 1150
rect 51096 1150 51112 1218
rect 52062 1218 52122 1394
rect 52062 1178 52080 1218
rect 51096 642 51102 1150
rect 51056 630 51102 642
rect 52074 642 52080 1178
rect 52114 1178 52122 1218
rect 52114 642 52120 1178
rect 52074 630 52120 642
rect 50326 592 50814 598
rect 50326 558 50338 592
rect 50802 558 50814 592
rect 50326 552 50814 558
rect 51344 592 51832 598
rect 51344 558 51356 592
rect 51820 558 51832 592
rect 51344 552 51832 558
rect 50026 434 50032 494
rect 50092 434 50098 494
rect 49008 322 49014 382
rect 49074 322 49080 382
rect 50032 -60 50092 434
rect 53020 382 53080 7310
rect 53232 6476 53292 14816
rect 53226 6416 53232 6476
rect 53292 6416 53298 6476
rect 53352 6348 53412 14818
rect 53346 6288 53352 6348
rect 53412 6288 53418 6348
rect 53492 5386 53552 14836
rect 53604 14698 53610 14758
rect 53670 14698 53676 14758
rect 53610 8630 53670 14698
rect 53720 14016 53780 14852
rect 53714 13956 53720 14016
rect 53780 13956 53786 14016
rect 53838 11096 53898 14952
rect 54166 14150 54226 14962
rect 54160 14090 54166 14150
rect 54226 14090 54232 14150
rect 53956 12732 53962 12792
rect 54022 12732 54028 12792
rect 53836 11090 53898 11096
rect 53896 11030 53898 11090
rect 53836 11024 53898 11030
rect 53604 8570 53610 8630
rect 53670 8570 53676 8630
rect 53486 5326 53492 5386
rect 53552 5326 53558 5386
rect 53838 5028 53898 11024
rect 53962 10096 54022 12732
rect 54168 12396 54174 12456
rect 54234 12396 54240 12456
rect 54064 11136 54070 11196
rect 54130 11136 54136 11196
rect 53956 10036 53962 10096
rect 54022 10036 54028 10096
rect 54070 5178 54130 11136
rect 54174 9860 54234 12396
rect 54286 9974 54346 14954
rect 54392 14878 54452 14884
rect 54392 12334 54452 14818
rect 65198 14522 65204 14528
rect 54518 14468 65204 14522
rect 65264 14522 65270 14528
rect 70302 14522 70308 14528
rect 65264 14468 70308 14522
rect 70368 14522 70374 14528
rect 74368 14522 74428 14528
rect 70368 14468 74368 14522
rect 54518 14462 74368 14468
rect 74428 14462 74940 14522
rect 54518 14322 54578 14462
rect 55040 14412 55100 14462
rect 56050 14412 56110 14462
rect 54814 14406 55302 14412
rect 54814 14372 54826 14406
rect 55290 14372 55302 14406
rect 54814 14366 55302 14372
rect 55832 14406 56320 14412
rect 55832 14372 55844 14406
rect 56308 14372 56320 14406
rect 55832 14366 56320 14372
rect 56050 14360 56110 14366
rect 54518 13746 54532 14322
rect 54566 13746 54578 14322
rect 55544 14322 55590 14334
rect 55544 13780 55550 14322
rect 54518 13504 54578 13746
rect 55536 13746 55550 13780
rect 55584 13780 55590 14322
rect 56556 14322 56616 14462
rect 57080 14412 57140 14462
rect 58092 14412 58152 14462
rect 56850 14406 57338 14412
rect 56850 14372 56862 14406
rect 57326 14372 57338 14406
rect 56850 14366 57338 14372
rect 57868 14406 58356 14412
rect 57868 14372 57880 14406
rect 58344 14372 58356 14406
rect 57868 14366 58356 14372
rect 58092 14360 58152 14366
rect 55584 13746 55596 13780
rect 54814 13696 55302 13702
rect 54814 13662 54826 13696
rect 55290 13662 55302 13696
rect 54814 13656 55302 13662
rect 55030 13594 55090 13656
rect 54814 13588 55302 13594
rect 54814 13554 54826 13588
rect 55290 13554 55302 13588
rect 54814 13548 55302 13554
rect 55030 13542 55090 13548
rect 54518 12928 54532 13504
rect 54566 12928 54578 13504
rect 54518 12456 54578 12928
rect 55536 13504 55596 13746
rect 56556 13746 56568 14322
rect 56602 13746 56616 14322
rect 57580 14322 57626 14334
rect 57580 13792 57586 14322
rect 56036 13702 56096 13704
rect 55832 13696 56320 13702
rect 55832 13662 55844 13696
rect 56308 13662 56320 13696
rect 55832 13656 56320 13662
rect 56036 13594 56096 13656
rect 55832 13588 56320 13594
rect 55832 13554 55844 13588
rect 56308 13554 56320 13588
rect 55832 13548 56320 13554
rect 55536 12928 55550 13504
rect 55584 12928 55596 13504
rect 56556 13504 56616 13746
rect 57570 13746 57586 13792
rect 57620 13792 57626 14322
rect 58588 14322 58648 14462
rect 59104 14412 59164 14462
rect 60104 14412 60164 14462
rect 58886 14406 59374 14412
rect 58886 14372 58898 14406
rect 59362 14372 59374 14406
rect 58886 14366 59374 14372
rect 59904 14406 60392 14412
rect 59904 14372 59916 14406
rect 60380 14372 60392 14406
rect 59904 14366 60392 14372
rect 57620 13746 57630 13792
rect 57048 13702 57108 13710
rect 56850 13696 57338 13702
rect 56850 13662 56862 13696
rect 57326 13662 57338 13696
rect 56850 13656 57338 13662
rect 57048 13594 57108 13656
rect 56850 13588 57338 13594
rect 56850 13554 56862 13588
rect 57326 13554 57338 13588
rect 56850 13548 57338 13554
rect 56556 13446 56568 13504
rect 54814 12878 55302 12884
rect 54814 12844 54826 12878
rect 55290 12844 55302 12878
rect 54814 12838 55302 12844
rect 55536 12792 55596 12928
rect 56562 12928 56568 13446
rect 56602 13446 56616 13504
rect 57570 13504 57630 13746
rect 58588 13746 58604 14322
rect 58638 13746 58648 14322
rect 59616 14322 59662 14334
rect 59616 13786 59622 14322
rect 57868 13696 58356 13702
rect 57868 13662 57880 13696
rect 58344 13662 58356 13696
rect 57868 13656 58356 13662
rect 58070 13594 58130 13656
rect 57868 13588 58356 13594
rect 57868 13554 57880 13588
rect 58344 13554 58356 13588
rect 57868 13548 58356 13554
rect 58070 13542 58130 13548
rect 56602 12928 56608 13446
rect 56562 12916 56608 12928
rect 57570 12928 57586 13504
rect 57620 12928 57630 13504
rect 58588 13504 58648 13746
rect 59606 13746 59622 13786
rect 59656 13786 59662 14322
rect 60626 14322 60686 14462
rect 61138 14412 61198 14462
rect 62150 14412 62210 14462
rect 60922 14406 61410 14412
rect 60922 14372 60934 14406
rect 61398 14372 61410 14406
rect 60922 14366 61410 14372
rect 61940 14406 62428 14412
rect 61940 14372 61952 14406
rect 62416 14372 62428 14406
rect 61940 14366 62428 14372
rect 59656 13746 59666 13786
rect 58886 13696 59374 13702
rect 58886 13662 58898 13696
rect 59362 13662 59374 13696
rect 58886 13656 59374 13662
rect 59082 13594 59142 13656
rect 58886 13588 59374 13594
rect 58886 13554 58898 13588
rect 59362 13554 59374 13588
rect 58886 13548 59374 13554
rect 59082 13542 59142 13548
rect 58588 13442 58604 13504
rect 55832 12878 56320 12884
rect 55832 12844 55844 12878
rect 56308 12844 56320 12878
rect 55832 12838 56320 12844
rect 56850 12878 57338 12884
rect 56850 12844 56862 12878
rect 57326 12844 57338 12878
rect 56850 12838 57338 12844
rect 57570 12790 57630 12928
rect 58598 12928 58604 13442
rect 58638 13442 58648 13504
rect 59606 13504 59666 13746
rect 60626 13746 60640 14322
rect 60674 13746 60686 14322
rect 61652 14322 61698 14334
rect 61652 13786 61658 14322
rect 59904 13696 60392 13702
rect 59904 13662 59916 13696
rect 60380 13662 60392 13696
rect 59904 13656 60392 13662
rect 60112 13594 60172 13656
rect 59904 13588 60392 13594
rect 59904 13554 59916 13588
rect 60380 13554 60392 13588
rect 59904 13548 60392 13554
rect 60112 13542 60172 13548
rect 58638 12928 58644 13442
rect 58598 12916 58644 12928
rect 59606 12928 59622 13504
rect 59656 12928 59666 13504
rect 60626 13504 60686 13746
rect 61644 13746 61658 13786
rect 61692 13786 61698 14322
rect 62662 14322 62722 14462
rect 63174 14412 63234 14462
rect 64186 14412 64246 14462
rect 62958 14406 63446 14412
rect 62958 14372 62970 14406
rect 63434 14372 63446 14406
rect 62958 14366 63446 14372
rect 63976 14406 64464 14412
rect 63976 14372 63988 14406
rect 64452 14372 64464 14406
rect 63976 14366 64464 14372
rect 61692 13746 61704 13786
rect 61118 13702 61178 13704
rect 60922 13696 61410 13702
rect 60922 13662 60934 13696
rect 61398 13662 61410 13696
rect 60922 13656 61410 13662
rect 61118 13594 61178 13656
rect 60922 13588 61410 13594
rect 60922 13554 60934 13588
rect 61398 13554 61410 13588
rect 60922 13548 61410 13554
rect 60626 13462 60640 13504
rect 57868 12878 58356 12884
rect 57868 12844 57880 12878
rect 58344 12844 58356 12878
rect 57868 12838 58356 12844
rect 58886 12878 59374 12884
rect 58886 12844 58898 12878
rect 59362 12844 59374 12878
rect 58886 12838 59374 12844
rect 59606 12790 59666 12928
rect 60634 12928 60640 13462
rect 60674 13462 60686 13504
rect 61644 13504 61704 13746
rect 62662 13746 62676 14322
rect 62710 13746 62722 14322
rect 63688 14322 63734 14334
rect 63688 13792 63694 14322
rect 62140 13702 62200 13704
rect 61940 13696 62428 13702
rect 61940 13662 61952 13696
rect 62416 13662 62428 13696
rect 61940 13656 62428 13662
rect 62140 13594 62200 13656
rect 61940 13588 62428 13594
rect 61940 13554 61952 13588
rect 62416 13554 62428 13588
rect 61940 13548 62428 13554
rect 60674 12928 60680 13462
rect 60634 12916 60680 12928
rect 61644 12928 61658 13504
rect 61692 12928 61704 13504
rect 62662 13504 62722 13746
rect 63682 13746 63694 13792
rect 63728 13792 63734 14322
rect 64694 14322 64754 14462
rect 65208 14412 65268 14462
rect 66220 14412 66280 14462
rect 64994 14406 65482 14412
rect 64994 14372 65006 14406
rect 65470 14372 65482 14406
rect 64994 14366 65482 14372
rect 66012 14406 66500 14412
rect 66012 14372 66024 14406
rect 66488 14372 66500 14406
rect 66012 14366 66500 14372
rect 66220 14360 66280 14366
rect 63728 13746 63742 13792
rect 62958 13696 63446 13702
rect 62958 13662 62970 13696
rect 63434 13662 63446 13696
rect 62958 13656 63446 13662
rect 63164 13594 63224 13656
rect 62958 13588 63446 13594
rect 62958 13554 62970 13588
rect 63434 13554 63446 13588
rect 62958 13548 63446 13554
rect 63164 13542 63224 13548
rect 62662 13454 62676 13504
rect 59904 12878 60392 12884
rect 59904 12844 59916 12878
rect 60380 12844 60392 12878
rect 59904 12838 60392 12844
rect 60922 12878 61410 12884
rect 60922 12844 60934 12878
rect 61398 12844 61410 12878
rect 60922 12838 61410 12844
rect 61644 12790 61704 12928
rect 62670 12928 62676 13454
rect 62710 13454 62722 13504
rect 63682 13504 63742 13746
rect 64694 13746 64712 14322
rect 64746 13746 64754 14322
rect 65724 14322 65770 14334
rect 65724 13792 65730 14322
rect 64170 13702 64230 13704
rect 63976 13696 64464 13702
rect 63976 13662 63988 13696
rect 64452 13662 64464 13696
rect 63976 13656 64464 13662
rect 64170 13594 64230 13656
rect 63976 13588 64464 13594
rect 63976 13554 63988 13588
rect 64452 13554 64464 13588
rect 63976 13548 64464 13554
rect 62710 12928 62716 13454
rect 62670 12916 62716 12928
rect 63682 12928 63694 13504
rect 63728 12928 63742 13504
rect 64694 13504 64754 13746
rect 65716 13746 65730 13792
rect 65764 13792 65770 14322
rect 66732 14322 66792 14462
rect 67244 14412 67304 14462
rect 68262 14412 68322 14462
rect 67030 14406 67518 14412
rect 67030 14372 67042 14406
rect 67506 14372 67518 14406
rect 67030 14366 67518 14372
rect 68048 14406 68536 14412
rect 68048 14372 68060 14406
rect 68524 14372 68536 14406
rect 68048 14366 68536 14372
rect 67244 14360 67304 14366
rect 65764 13746 65776 13792
rect 65194 13702 65254 13710
rect 64994 13696 65482 13702
rect 64994 13662 65006 13696
rect 65470 13662 65482 13696
rect 64994 13656 65482 13662
rect 65194 13594 65254 13656
rect 64994 13588 65482 13594
rect 64994 13554 65006 13588
rect 65470 13554 65482 13588
rect 64994 13548 65482 13554
rect 64694 13456 64712 13504
rect 61940 12878 62428 12884
rect 61940 12844 61952 12878
rect 62416 12844 62428 12878
rect 61940 12838 62428 12844
rect 62958 12878 63446 12884
rect 62958 12844 62970 12878
rect 63434 12844 63446 12878
rect 62958 12838 63446 12844
rect 63682 12790 63742 12928
rect 64706 12928 64712 13456
rect 64746 13456 64754 13504
rect 65716 13504 65776 13746
rect 66732 13746 66748 14322
rect 66782 13746 66792 14322
rect 67760 14322 67806 14334
rect 67760 13792 67766 14322
rect 66216 13702 66276 13704
rect 66012 13696 66500 13702
rect 66012 13662 66024 13696
rect 66488 13662 66500 13696
rect 66012 13656 66500 13662
rect 66216 13594 66276 13656
rect 66012 13588 66500 13594
rect 66012 13554 66024 13588
rect 66488 13554 66500 13588
rect 66012 13548 66500 13554
rect 64746 12928 64752 13456
rect 64706 12916 64752 12928
rect 65716 12928 65730 13504
rect 65764 12928 65776 13504
rect 66732 13504 66792 13746
rect 67752 13746 67766 13792
rect 67800 13792 67806 14322
rect 68768 14322 68828 14462
rect 69284 14412 69344 14462
rect 70308 14412 70368 14462
rect 69066 14406 69554 14412
rect 69066 14372 69078 14406
rect 69542 14372 69554 14406
rect 69066 14366 69554 14372
rect 70084 14406 70572 14412
rect 70084 14372 70096 14406
rect 70560 14372 70572 14406
rect 70084 14366 70572 14372
rect 67800 13746 67812 13792
rect 67228 13702 67288 13704
rect 67030 13696 67518 13702
rect 67030 13662 67042 13696
rect 67506 13662 67518 13696
rect 67030 13656 67518 13662
rect 67228 13594 67288 13656
rect 67030 13588 67518 13594
rect 67030 13554 67042 13588
rect 67506 13554 67518 13588
rect 67030 13548 67518 13554
rect 66732 13454 66748 13504
rect 63976 12878 64464 12884
rect 63976 12844 63988 12878
rect 64452 12844 64464 12878
rect 63976 12838 64464 12844
rect 64994 12878 65482 12884
rect 64994 12844 65006 12878
rect 65470 12844 65482 12878
rect 64994 12838 65482 12844
rect 65716 12790 65776 12928
rect 66742 12928 66748 13454
rect 66782 13454 66792 13504
rect 67752 13504 67812 13746
rect 68768 13746 68784 14322
rect 68818 13746 68828 14322
rect 69796 14322 69842 14334
rect 69796 13816 69802 14322
rect 68048 13696 68536 13702
rect 68048 13662 68060 13696
rect 68524 13662 68536 13696
rect 68048 13656 68536 13662
rect 68240 13594 68300 13656
rect 68048 13588 68536 13594
rect 68048 13554 68060 13588
rect 68524 13554 68536 13588
rect 68048 13548 68536 13554
rect 68240 13542 68300 13548
rect 66782 12928 66788 13454
rect 66742 12916 66788 12928
rect 67752 12928 67766 13504
rect 67800 12928 67812 13504
rect 68768 13504 68828 13746
rect 69790 13746 69802 13816
rect 69836 13816 69842 14322
rect 70804 14322 70864 14462
rect 71326 14412 71386 14462
rect 72338 14412 72398 14462
rect 71102 14406 71590 14412
rect 71102 14372 71114 14406
rect 71578 14372 71590 14406
rect 71102 14366 71590 14372
rect 72120 14406 72608 14412
rect 72120 14372 72132 14406
rect 72596 14372 72608 14406
rect 72120 14366 72608 14372
rect 69836 13746 69850 13816
rect 69264 13702 69324 13710
rect 69066 13696 69554 13702
rect 69066 13662 69078 13696
rect 69542 13662 69554 13696
rect 69066 13656 69554 13662
rect 69264 13594 69324 13656
rect 69066 13588 69554 13594
rect 69066 13554 69078 13588
rect 69542 13554 69554 13588
rect 69066 13548 69554 13554
rect 68768 13480 68784 13504
rect 66012 12878 66500 12884
rect 66012 12844 66024 12878
rect 66488 12844 66500 12878
rect 66012 12838 66500 12844
rect 67030 12878 67518 12884
rect 67030 12844 67042 12878
rect 67506 12844 67518 12878
rect 67030 12838 67518 12844
rect 67752 12790 67812 12928
rect 68778 12928 68784 13480
rect 68818 13480 68828 13504
rect 69790 13504 69850 13746
rect 70804 13746 70820 14322
rect 70854 13746 70864 14322
rect 71832 14322 71878 14334
rect 71832 13856 71838 14322
rect 70084 13696 70572 13702
rect 70084 13662 70096 13696
rect 70560 13662 70572 13696
rect 70084 13656 70572 13662
rect 70286 13594 70346 13656
rect 70084 13588 70572 13594
rect 70084 13554 70096 13588
rect 70560 13554 70572 13588
rect 70084 13548 70572 13554
rect 70286 13536 70346 13548
rect 68818 12928 68824 13480
rect 68778 12916 68824 12928
rect 69790 12928 69802 13504
rect 69836 12928 69850 13504
rect 70804 13504 70864 13746
rect 71824 13746 71838 13856
rect 71872 13856 71878 14322
rect 72842 14322 72902 14462
rect 73348 14412 73408 14462
rect 74366 14456 74428 14462
rect 74366 14412 74426 14456
rect 73138 14406 73626 14412
rect 73138 14372 73150 14406
rect 73614 14372 73626 14406
rect 73138 14366 73626 14372
rect 74156 14406 74644 14412
rect 74156 14372 74168 14406
rect 74632 14372 74644 14406
rect 74156 14366 74644 14372
rect 71872 13746 71884 13856
rect 71304 13702 71364 13704
rect 71102 13696 71590 13702
rect 71102 13662 71114 13696
rect 71578 13662 71590 13696
rect 71102 13656 71590 13662
rect 71304 13594 71364 13656
rect 71102 13588 71590 13594
rect 71102 13554 71114 13588
rect 71578 13554 71590 13588
rect 71102 13548 71590 13554
rect 70804 13462 70820 13504
rect 68048 12878 68536 12884
rect 68048 12844 68060 12878
rect 68524 12844 68536 12878
rect 68048 12838 68536 12844
rect 69066 12878 69554 12884
rect 69066 12844 69078 12878
rect 69542 12844 69554 12878
rect 69066 12838 69554 12844
rect 69790 12790 69850 12928
rect 70814 12928 70820 13462
rect 70854 13462 70864 13504
rect 71824 13504 71884 13746
rect 72842 13746 72856 14322
rect 72890 13746 72902 14322
rect 73868 14322 73914 14334
rect 73868 13806 73874 14322
rect 72334 13702 72394 13716
rect 72120 13696 72608 13702
rect 72120 13662 72132 13696
rect 72596 13662 72608 13696
rect 72120 13656 72608 13662
rect 72334 13594 72394 13656
rect 72120 13588 72608 13594
rect 72120 13554 72132 13588
rect 72596 13554 72608 13588
rect 72120 13548 72608 13554
rect 70854 12928 70860 13462
rect 70814 12916 70860 12928
rect 71824 12928 71838 13504
rect 71872 12928 71884 13504
rect 72842 13504 72902 13746
rect 73860 13746 73874 13806
rect 73908 13806 73914 14322
rect 74880 14322 74940 14462
rect 73908 13746 73920 13806
rect 73346 13702 73406 13716
rect 73138 13696 73626 13702
rect 73138 13662 73150 13696
rect 73614 13662 73626 13696
rect 73138 13656 73626 13662
rect 73346 13594 73406 13656
rect 73138 13588 73626 13594
rect 73138 13554 73150 13588
rect 73614 13554 73626 13588
rect 73138 13548 73626 13554
rect 72842 13462 72856 13504
rect 70084 12878 70572 12884
rect 70084 12844 70096 12878
rect 70560 12844 70572 12878
rect 70084 12838 70572 12844
rect 71102 12878 71590 12884
rect 71102 12844 71114 12878
rect 71578 12844 71590 12878
rect 71102 12838 71590 12844
rect 71824 12790 71884 12928
rect 72850 12928 72856 13462
rect 72890 13462 72902 13504
rect 73860 13504 73920 13746
rect 74880 13746 74892 14322
rect 74926 13746 74940 14322
rect 74156 13696 74644 13702
rect 74156 13662 74168 13696
rect 74632 13662 74644 13696
rect 74156 13656 74644 13662
rect 74346 13594 74406 13656
rect 74880 13654 74940 13746
rect 76766 14300 76878 15086
rect 74880 13594 75660 13654
rect 74156 13588 74644 13594
rect 74156 13554 74168 13588
rect 74632 13554 74644 13588
rect 74156 13548 74644 13554
rect 74346 13542 74406 13548
rect 72890 12928 72896 13462
rect 72850 12916 72896 12928
rect 73860 12928 73874 13504
rect 73908 12928 73920 13504
rect 74880 13504 74940 13594
rect 74880 13454 74892 13504
rect 72120 12878 72608 12884
rect 72120 12844 72132 12878
rect 72596 12844 72608 12878
rect 72120 12838 72608 12844
rect 73138 12878 73626 12884
rect 73138 12844 73150 12878
rect 73614 12844 73626 12878
rect 73138 12838 73626 12844
rect 73860 12790 73920 12928
rect 74886 12928 74892 13454
rect 74926 13454 74940 13504
rect 74926 12928 74932 13454
rect 74886 12916 74932 12928
rect 74156 12878 74644 12884
rect 74156 12844 74168 12878
rect 74632 12844 74644 12878
rect 74156 12838 74644 12844
rect 55596 12732 75538 12790
rect 55536 12730 75538 12732
rect 55536 12726 55596 12730
rect 56544 12516 56550 12576
rect 56610 12516 56616 12576
rect 58584 12516 58590 12576
rect 58650 12516 58656 12576
rect 60624 12516 60630 12576
rect 60690 12516 60696 12576
rect 62654 12516 62660 12576
rect 62720 12516 62726 12576
rect 64694 12516 64700 12576
rect 64760 12516 64766 12576
rect 66726 12516 66732 12576
rect 66792 12516 66798 12576
rect 68766 12516 68772 12576
rect 68832 12516 68838 12576
rect 70802 12516 70808 12576
rect 70868 12516 70874 12576
rect 72836 12516 72842 12576
rect 72902 12516 72908 12576
rect 54512 12396 54518 12456
rect 54578 12396 54584 12456
rect 56036 12390 56042 12450
rect 56102 12390 56108 12450
rect 54386 12274 54392 12334
rect 54452 12274 54458 12334
rect 54392 10200 54452 12274
rect 56042 12216 56102 12390
rect 54814 12210 55302 12216
rect 54814 12176 54826 12210
rect 55290 12176 55302 12210
rect 54814 12170 55302 12176
rect 55832 12210 56320 12216
rect 55832 12176 55844 12210
rect 56308 12176 56320 12210
rect 55832 12170 56320 12176
rect 54526 12126 54572 12138
rect 55544 12126 55590 12138
rect 56550 12126 56610 12516
rect 57056 12450 57116 12456
rect 57056 12216 57116 12390
rect 58078 12450 58138 12456
rect 58078 12216 58138 12390
rect 56850 12210 57338 12216
rect 56850 12176 56862 12210
rect 57326 12176 57338 12210
rect 56850 12170 57338 12176
rect 57868 12210 58356 12216
rect 57868 12176 57880 12210
rect 58344 12176 58356 12210
rect 57868 12170 58356 12176
rect 57580 12126 57626 12138
rect 54518 12092 54532 12126
rect 54526 11600 54532 12092
rect 54518 11550 54532 11600
rect 54566 12092 54578 12126
rect 54566 11600 54572 12092
rect 55536 12078 55550 12126
rect 54566 11550 54578 11600
rect 55544 11586 55550 12078
rect 54518 11412 54578 11550
rect 55536 11550 55550 11586
rect 55584 12078 55596 12126
rect 55584 11586 55590 12078
rect 56550 12058 56568 12126
rect 56562 11614 56568 12058
rect 55584 11550 55596 11586
rect 54814 11500 55302 11506
rect 54814 11466 54826 11500
rect 55290 11466 55302 11500
rect 54814 11460 55302 11466
rect 55020 11412 55080 11460
rect 55536 11412 55596 11550
rect 56554 11550 56568 11614
rect 56602 12094 56614 12126
rect 56602 12058 56610 12094
rect 56602 11614 56608 12058
rect 56602 11550 56614 11614
rect 57580 11596 57586 12126
rect 57576 11578 57586 11596
rect 57574 11550 57586 11578
rect 57620 11596 57626 12126
rect 58590 12126 58650 12516
rect 59092 12450 59152 12456
rect 59090 12390 59092 12396
rect 60118 12450 60178 12456
rect 59090 12384 59152 12390
rect 60116 12390 60118 12396
rect 60116 12384 60178 12390
rect 59090 12216 59150 12384
rect 59600 12274 59606 12334
rect 59666 12274 59672 12334
rect 58886 12210 59374 12216
rect 58886 12176 58898 12210
rect 59362 12176 59374 12210
rect 58886 12170 59374 12176
rect 58590 12072 58604 12126
rect 58598 11622 58604 12072
rect 58594 11598 58604 11622
rect 57620 11550 57636 11596
rect 58592 11550 58604 11598
rect 58638 12072 58650 12126
rect 59606 12126 59666 12274
rect 60116 12216 60176 12384
rect 59904 12210 60392 12216
rect 59904 12176 59916 12210
rect 60380 12176 60392 12210
rect 59904 12170 60392 12176
rect 59606 12084 59622 12126
rect 58638 11622 58644 12072
rect 59616 11626 59622 12084
rect 58638 11550 58654 11622
rect 59606 11550 59622 11626
rect 59656 12084 59666 12126
rect 60630 12126 60690 12516
rect 61130 12450 61190 12456
rect 61130 12216 61190 12390
rect 62166 12450 62226 12456
rect 62166 12216 62226 12390
rect 60922 12210 61410 12216
rect 60922 12176 60934 12210
rect 61398 12176 61410 12210
rect 60922 12170 61410 12176
rect 61940 12210 62428 12216
rect 61940 12176 61952 12210
rect 62416 12176 62428 12210
rect 61940 12170 62428 12176
rect 61652 12126 61698 12138
rect 62660 12126 62720 12516
rect 63172 12450 63232 12456
rect 64180 12390 64186 12450
rect 64246 12390 64252 12450
rect 63172 12216 63232 12390
rect 64186 12216 64246 12390
rect 62958 12210 63446 12216
rect 62958 12176 62970 12210
rect 63434 12176 63446 12210
rect 62958 12170 63446 12176
rect 63976 12210 64464 12216
rect 63976 12176 63988 12210
rect 64452 12176 64464 12210
rect 63976 12170 64464 12176
rect 59656 11626 59662 12084
rect 60630 12052 60640 12126
rect 59656 11610 59666 11626
rect 59656 11550 59670 11610
rect 60634 11606 60640 12052
rect 60626 11550 60640 11606
rect 60674 12052 60690 12126
rect 61646 12076 61658 12126
rect 60674 11606 60680 12052
rect 61652 11614 61658 12076
rect 60674 11550 60686 11606
rect 61646 11586 61658 11614
rect 61644 11550 61658 11586
rect 61692 12076 61706 12126
rect 61692 11614 61698 12076
rect 62660 12058 62676 12126
rect 62670 11626 62676 12058
rect 61692 11550 61706 11614
rect 55832 11500 56320 11506
rect 55832 11466 55844 11500
rect 56308 11466 56320 11500
rect 55832 11460 56320 11466
rect 54518 11352 55596 11412
rect 55536 11196 55596 11352
rect 56046 11302 56106 11460
rect 56554 11412 56614 11550
rect 56850 11500 57338 11506
rect 56850 11466 56862 11500
rect 57326 11466 57338 11500
rect 56850 11460 57338 11466
rect 56548 11352 56554 11412
rect 56614 11352 56620 11412
rect 56040 11242 56046 11302
rect 56106 11242 56112 11302
rect 55530 11136 55536 11196
rect 55596 11136 55602 11196
rect 54516 11030 54522 11090
rect 54582 11030 54588 11090
rect 55014 11030 55020 11090
rect 55080 11030 55086 11090
rect 55526 11030 55532 11090
rect 55592 11030 55598 11090
rect 54522 10894 54582 11030
rect 55020 10984 55080 11030
rect 54814 10978 55302 10984
rect 54814 10944 54826 10978
rect 55290 10944 55302 10978
rect 54814 10938 55302 10944
rect 54522 10854 54532 10894
rect 54526 10318 54532 10854
rect 54566 10854 54582 10894
rect 55532 10894 55592 11030
rect 56046 10984 56106 11242
rect 55832 10978 56320 10984
rect 55832 10944 55844 10978
rect 56308 10944 56320 10978
rect 55832 10938 56320 10944
rect 54566 10318 54572 10854
rect 55532 10848 55550 10894
rect 54526 10306 54572 10318
rect 55544 10318 55550 10848
rect 55584 10848 55592 10894
rect 56554 10894 56614 11352
rect 57068 11302 57128 11460
rect 57062 11242 57068 11302
rect 57128 11242 57134 11302
rect 57068 10984 57128 11242
rect 57576 11196 57636 11550
rect 57868 11500 58356 11506
rect 57868 11466 57880 11500
rect 58344 11466 58356 11500
rect 57868 11460 58356 11466
rect 58082 11302 58142 11460
rect 58594 11412 58654 11550
rect 59616 11538 59662 11550
rect 58886 11500 59374 11506
rect 58886 11466 58898 11500
rect 59362 11466 59374 11500
rect 58886 11460 59374 11466
rect 59904 11500 60392 11506
rect 59904 11466 59916 11500
rect 60380 11466 60392 11500
rect 59904 11460 60392 11466
rect 58588 11352 58594 11412
rect 58654 11352 58660 11412
rect 58076 11242 58082 11302
rect 58142 11242 58148 11302
rect 57570 11136 57576 11196
rect 57636 11136 57642 11196
rect 58082 10984 58142 11242
rect 56850 10978 57338 10984
rect 56850 10944 56862 10978
rect 57326 10944 57338 10978
rect 56850 10938 57338 10944
rect 57868 10978 58356 10984
rect 57868 10944 57880 10978
rect 58344 10944 58356 10978
rect 57868 10938 58356 10944
rect 57580 10894 57626 10906
rect 58594 10894 58654 11352
rect 59096 11302 59156 11460
rect 60114 11302 60174 11460
rect 60626 11412 60686 11550
rect 60922 11500 61410 11506
rect 60922 11466 60934 11500
rect 61398 11466 61410 11500
rect 60922 11460 61410 11466
rect 60620 11352 60626 11412
rect 60686 11352 60692 11412
rect 59090 11242 59096 11302
rect 59156 11242 59162 11302
rect 60108 11242 60114 11302
rect 60174 11242 60180 11302
rect 59096 10984 59156 11242
rect 59600 11136 59606 11196
rect 59666 11136 59672 11196
rect 58886 10978 59374 10984
rect 58886 10944 58898 10978
rect 59362 10944 59374 10978
rect 58886 10938 59374 10944
rect 56554 10856 56568 10894
rect 55584 10318 55590 10848
rect 56562 10376 56568 10856
rect 55544 10306 55590 10318
rect 56548 10318 56568 10376
rect 56602 10856 56614 10894
rect 56602 10318 56608 10856
rect 57574 10842 57586 10894
rect 57580 10338 57586 10842
rect 54814 10268 55302 10274
rect 54814 10234 54826 10268
rect 55290 10234 55302 10268
rect 54814 10228 55302 10234
rect 55832 10268 56320 10274
rect 55832 10234 55844 10268
rect 56308 10234 56320 10268
rect 55832 10228 56320 10234
rect 54386 10140 54392 10200
rect 54452 10140 54458 10200
rect 56548 10096 56608 10318
rect 57570 10318 57586 10338
rect 57620 10842 57634 10894
rect 57620 10338 57626 10842
rect 58592 10830 58604 10894
rect 58598 10382 58604 10830
rect 57620 10318 57630 10338
rect 56850 10268 57338 10274
rect 56850 10234 56862 10268
rect 57326 10234 57338 10268
rect 56850 10228 57338 10234
rect 54510 10036 54516 10096
rect 54576 10036 54582 10096
rect 56030 10036 56036 10096
rect 56096 10036 56102 10096
rect 56542 10036 56548 10096
rect 56608 10036 56614 10096
rect 54280 9914 54286 9974
rect 54346 9914 54352 9974
rect 54168 9800 54174 9860
rect 54234 9800 54240 9860
rect 54286 8732 54346 9914
rect 54516 9660 54576 10036
rect 55016 9800 55022 9860
rect 55082 9800 55088 9860
rect 55022 9750 55082 9800
rect 56036 9750 56096 10036
rect 56548 9802 56554 9862
rect 56614 9802 56620 9862
rect 54812 9744 55300 9750
rect 54812 9710 54824 9744
rect 55288 9710 55300 9744
rect 54812 9704 55300 9710
rect 55830 9744 56318 9750
rect 55830 9710 55842 9744
rect 56306 9710 56318 9744
rect 55830 9704 56318 9710
rect 55542 9660 55588 9672
rect 56554 9660 56614 9802
rect 57052 9750 57112 10228
rect 57570 10200 57630 10318
rect 58584 10318 58604 10382
rect 58638 10860 58654 10894
rect 59606 10894 59666 11136
rect 60114 10984 60174 11242
rect 59904 10978 60392 10984
rect 59904 10944 59916 10978
rect 60380 10944 60392 10978
rect 59904 10938 60392 10944
rect 60626 10894 60686 11352
rect 61140 11302 61200 11460
rect 61646 11342 61706 11550
rect 62658 11550 62676 11626
rect 62710 12058 62720 12126
rect 63688 12126 63734 12138
rect 62710 11626 62716 12058
rect 62710 11550 62718 11626
rect 63688 11612 63694 12126
rect 63682 11610 63694 11612
rect 61940 11500 62428 11506
rect 61940 11466 61952 11500
rect 62416 11466 62428 11500
rect 61940 11460 62428 11466
rect 61134 11242 61140 11302
rect 61200 11242 61206 11302
rect 61646 11282 61872 11342
rect 62160 11302 62220 11460
rect 62658 11412 62718 11550
rect 63680 11550 63694 11610
rect 63728 11612 63734 12126
rect 64700 12126 64760 12516
rect 65202 12450 65262 12456
rect 65202 12216 65262 12390
rect 66210 12450 66270 12456
rect 66270 12390 66272 12396
rect 66210 12384 66272 12390
rect 66212 12216 66272 12384
rect 64994 12210 65482 12216
rect 64994 12176 65006 12210
rect 65470 12176 65482 12210
rect 64994 12170 65482 12176
rect 66012 12210 66500 12216
rect 66012 12176 66024 12210
rect 66488 12176 66500 12210
rect 66012 12170 66500 12176
rect 65724 12126 65770 12138
rect 66732 12126 66792 12516
rect 67226 12450 67286 12456
rect 68250 12450 68310 12456
rect 67286 12390 67288 12396
rect 67226 12384 67288 12390
rect 67228 12216 67288 12384
rect 68250 12216 68310 12390
rect 67030 12210 67518 12216
rect 67030 12176 67042 12210
rect 67506 12176 67518 12210
rect 67030 12170 67518 12176
rect 68048 12210 68536 12216
rect 68048 12176 68060 12210
rect 68524 12176 68536 12210
rect 68048 12170 68536 12176
rect 67760 12126 67806 12138
rect 68772 12126 68832 12516
rect 69272 12450 69332 12456
rect 70294 12450 70354 12456
rect 69272 12216 69332 12390
rect 70292 12390 70294 12396
rect 70292 12384 70354 12390
rect 69788 12274 69794 12334
rect 69854 12274 69860 12334
rect 69066 12210 69554 12216
rect 69066 12176 69078 12210
rect 69542 12176 69554 12210
rect 69066 12170 69554 12176
rect 64700 12058 64712 12126
rect 64706 11616 64712 12058
rect 63728 11550 63742 11612
rect 64694 11550 64712 11616
rect 64746 12058 64760 12126
rect 65714 12092 65730 12126
rect 64746 11616 64752 12058
rect 64746 11550 64754 11616
rect 65724 11598 65730 12092
rect 62958 11500 63446 11506
rect 62958 11466 62970 11500
rect 63434 11466 63446 11500
rect 62958 11460 63446 11466
rect 62652 11352 62658 11412
rect 62718 11352 62724 11412
rect 61140 10984 61200 11242
rect 61640 11136 61646 11196
rect 61706 11136 61712 11196
rect 60922 10978 61410 10984
rect 60922 10944 60934 10978
rect 61398 10944 61410 10978
rect 60922 10938 61410 10944
rect 61646 10894 61706 11136
rect 61812 11090 61872 11282
rect 62154 11242 62160 11302
rect 62220 11242 62226 11302
rect 61806 11030 61812 11090
rect 61872 11030 61878 11090
rect 62160 10984 62220 11242
rect 61940 10978 62428 10984
rect 61940 10944 61952 10978
rect 62416 10944 62428 10978
rect 61940 10938 62428 10944
rect 58638 10830 58652 10860
rect 59606 10850 59622 10894
rect 58638 10318 58644 10830
rect 57868 10268 58356 10274
rect 57868 10234 57880 10268
rect 58344 10234 58356 10268
rect 57868 10228 58356 10234
rect 57564 10140 57570 10200
rect 57630 10140 57636 10200
rect 57566 10036 57572 10096
rect 57632 10036 57638 10096
rect 56848 9744 57336 9750
rect 56848 9710 56860 9744
rect 57324 9710 57336 9744
rect 56848 9704 57336 9710
rect 54516 9604 54530 9660
rect 54524 9084 54530 9604
rect 54564 9604 54576 9660
rect 55536 9628 55548 9660
rect 54564 9084 54570 9604
rect 55542 9128 55548 9628
rect 54524 9072 54570 9084
rect 55536 9084 55548 9128
rect 55582 9628 55596 9660
rect 56554 9634 56566 9660
rect 55582 9128 55588 9628
rect 55582 9084 55596 9128
rect 54812 9034 55300 9040
rect 54812 9000 54824 9034
rect 55288 9000 55300 9034
rect 54812 8994 55300 9000
rect 55536 8932 55596 9084
rect 56560 9084 56566 9634
rect 56600 9634 56614 9660
rect 57572 9660 57632 10036
rect 58072 9750 58132 10228
rect 58584 10096 58644 10318
rect 59616 10318 59622 10850
rect 59656 10860 59668 10894
rect 59656 10850 59666 10860
rect 60626 10852 60640 10894
rect 59656 10318 59662 10850
rect 60634 10360 60640 10852
rect 60626 10318 60640 10360
rect 60674 10852 60686 10894
rect 60674 10360 60680 10852
rect 61642 10832 61658 10894
rect 60674 10318 60686 10360
rect 61652 10318 61658 10832
rect 61692 10854 61706 10894
rect 62658 10894 62718 11352
rect 63180 11302 63240 11460
rect 63174 11242 63180 11302
rect 63240 11242 63246 11302
rect 63180 10984 63240 11242
rect 63680 11196 63740 11550
rect 63976 11500 64464 11506
rect 63976 11466 63988 11500
rect 64452 11466 64464 11500
rect 63976 11460 64464 11466
rect 64182 11302 64242 11460
rect 64694 11412 64754 11550
rect 65716 11550 65730 11598
rect 65764 12092 65774 12126
rect 65764 11598 65770 12092
rect 66732 12072 66748 12126
rect 66742 11610 66748 12072
rect 65764 11550 65776 11598
rect 64994 11500 65482 11506
rect 64994 11466 65006 11500
rect 65470 11466 65482 11500
rect 64994 11460 65482 11466
rect 64688 11352 64694 11412
rect 64754 11352 64760 11412
rect 64176 11242 64182 11302
rect 64242 11242 64248 11302
rect 63674 11136 63680 11196
rect 63740 11136 63746 11196
rect 63674 11030 63680 11090
rect 63740 11030 63746 11090
rect 62958 10978 63446 10984
rect 62958 10944 62970 10978
rect 63434 10944 63446 10978
rect 62958 10938 63446 10944
rect 63680 10894 63740 11030
rect 64182 10984 64242 11242
rect 63976 10978 64464 10984
rect 63976 10944 63988 10978
rect 64452 10944 64464 10978
rect 63976 10938 64464 10944
rect 64694 10894 64754 11352
rect 65208 11302 65268 11460
rect 65202 11242 65208 11302
rect 65268 11242 65274 11302
rect 65208 10984 65268 11242
rect 65716 11196 65776 11550
rect 66730 11550 66748 11610
rect 66782 12072 66792 12126
rect 67752 12086 67766 12126
rect 66782 11610 66788 12072
rect 67760 11616 67766 12086
rect 66782 11550 66790 11610
rect 67756 11590 67766 11616
rect 66012 11500 66500 11506
rect 66012 11466 66024 11500
rect 66488 11466 66500 11500
rect 66012 11460 66500 11466
rect 66226 11302 66286 11460
rect 66730 11412 66790 11550
rect 67754 11550 67766 11590
rect 67800 12086 67812 12126
rect 67800 11616 67806 12086
rect 68772 12072 68784 12126
rect 67800 11550 67816 11616
rect 68778 11600 68784 12072
rect 68768 11550 68784 11600
rect 68818 12072 68832 12126
rect 69794 12126 69854 12274
rect 70292 12216 70352 12384
rect 70084 12210 70572 12216
rect 70084 12176 70096 12210
rect 70560 12176 70572 12210
rect 70084 12170 70572 12176
rect 68818 11600 68824 12072
rect 69794 12062 69802 12126
rect 69796 11606 69802 12062
rect 68818 11550 68828 11600
rect 69788 11550 69802 11606
rect 69836 12062 69854 12126
rect 70808 12126 70868 12516
rect 71312 12450 71372 12456
rect 72326 12450 72386 12456
rect 71372 12390 71374 12396
rect 71312 12384 71374 12390
rect 72386 12390 72388 12396
rect 72326 12384 72388 12390
rect 71314 12216 71374 12384
rect 72328 12216 72388 12384
rect 71102 12210 71590 12216
rect 71102 12176 71114 12210
rect 71578 12176 71590 12210
rect 71102 12170 71590 12176
rect 72120 12210 72608 12216
rect 72120 12176 72132 12210
rect 72596 12176 72608 12210
rect 72120 12170 72608 12176
rect 71832 12126 71878 12138
rect 72842 12126 72902 12516
rect 73350 12450 73410 12456
rect 73348 12390 73350 12396
rect 73348 12384 73410 12390
rect 73348 12216 73408 12384
rect 73860 12274 73866 12334
rect 73926 12274 73932 12334
rect 74992 12274 74998 12334
rect 75058 12274 75064 12334
rect 73138 12210 73626 12216
rect 73138 12176 73150 12210
rect 73614 12176 73626 12210
rect 73138 12170 73626 12176
rect 73866 12126 73926 12274
rect 74156 12210 74644 12216
rect 74156 12176 74168 12210
rect 74632 12176 74644 12210
rect 74156 12170 74644 12176
rect 70808 12066 70820 12126
rect 69836 11606 69842 12062
rect 69836 11604 69848 11606
rect 69836 11550 69850 11604
rect 70814 11586 70820 12066
rect 70806 11550 70820 11586
rect 70854 12066 70868 12126
rect 71824 12086 71838 12126
rect 70854 11586 70860 12066
rect 71832 11606 71838 12086
rect 70854 11550 70866 11586
rect 67030 11500 67518 11506
rect 67030 11466 67042 11500
rect 67506 11466 67518 11500
rect 67030 11460 67518 11466
rect 66724 11352 66730 11412
rect 66790 11352 66796 11412
rect 66220 11242 66226 11302
rect 66286 11242 66292 11302
rect 65710 11136 65716 11196
rect 65776 11136 65782 11196
rect 65712 11030 65718 11090
rect 65778 11030 65784 11090
rect 64994 10978 65482 10984
rect 64994 10944 65006 10978
rect 65470 10944 65482 10978
rect 64994 10938 65482 10944
rect 65718 10894 65778 11030
rect 66226 10984 66286 11242
rect 66012 10978 66500 10984
rect 66012 10944 66024 10978
rect 66488 10944 66500 10978
rect 66012 10938 66500 10944
rect 66730 10894 66790 11352
rect 67234 11302 67294 11460
rect 67754 11334 67814 11550
rect 68246 11506 68306 11508
rect 68048 11500 68536 11506
rect 68048 11466 68060 11500
rect 68524 11466 68536 11500
rect 68048 11460 68536 11466
rect 67228 11242 67234 11302
rect 67294 11242 67300 11302
rect 67598 11274 67814 11334
rect 68246 11302 68306 11460
rect 68768 11412 68828 11550
rect 69796 11538 69842 11550
rect 69278 11506 69338 11508
rect 69066 11500 69554 11506
rect 69066 11466 69078 11500
rect 69542 11466 69554 11500
rect 69066 11460 69554 11466
rect 70084 11500 70572 11506
rect 70084 11466 70096 11500
rect 70560 11466 70572 11500
rect 70084 11460 70572 11466
rect 68762 11352 68768 11412
rect 68828 11352 68834 11412
rect 67234 10984 67294 11242
rect 67598 11090 67658 11274
rect 68240 11242 68246 11302
rect 68306 11242 68312 11302
rect 67746 11136 67752 11196
rect 67812 11136 67818 11196
rect 67592 11030 67598 11090
rect 67658 11030 67664 11090
rect 67030 10978 67518 10984
rect 67030 10944 67042 10978
rect 67506 10944 67518 10978
rect 67030 10938 67518 10944
rect 61692 10832 61702 10854
rect 62658 10838 62676 10894
rect 61692 10318 61698 10832
rect 62670 10360 62676 10838
rect 59616 10306 59662 10318
rect 60634 10306 60680 10318
rect 61652 10306 61698 10318
rect 62662 10318 62676 10360
rect 62710 10838 62718 10894
rect 63678 10842 63694 10894
rect 62710 10360 62716 10838
rect 62710 10318 62722 10360
rect 58886 10268 59374 10274
rect 58886 10234 58898 10268
rect 59362 10234 59374 10268
rect 58886 10228 59374 10234
rect 59904 10268 60392 10274
rect 59904 10234 59916 10268
rect 60380 10234 60392 10268
rect 59904 10228 60392 10234
rect 60922 10268 61410 10274
rect 60922 10234 60934 10268
rect 61398 10234 61410 10268
rect 60922 10228 61410 10234
rect 61940 10268 62428 10274
rect 61940 10234 61952 10268
rect 62416 10234 62428 10268
rect 61940 10228 62428 10234
rect 58578 10036 58584 10096
rect 58644 10036 58650 10096
rect 58584 9802 58590 9862
rect 58650 9802 58656 9862
rect 57866 9744 58354 9750
rect 57866 9710 57878 9744
rect 58342 9710 58354 9744
rect 57866 9704 58354 9710
rect 56600 9084 56606 9634
rect 57572 9628 57584 9660
rect 57578 9124 57584 9628
rect 56560 9072 56606 9084
rect 57570 9084 57584 9124
rect 57618 9628 57632 9660
rect 58590 9660 58650 9802
rect 59084 9750 59144 10228
rect 59598 10036 59604 10096
rect 59664 10036 59670 10096
rect 58884 9744 59372 9750
rect 58884 9710 58896 9744
rect 59360 9710 59372 9744
rect 58884 9704 59372 9710
rect 58590 9630 58602 9660
rect 57618 9124 57624 9628
rect 57618 9084 57630 9124
rect 55830 9034 56318 9040
rect 55830 9000 55842 9034
rect 56306 9000 56318 9034
rect 55830 8994 56318 9000
rect 56848 9034 57336 9040
rect 56848 9000 56860 9034
rect 57324 9000 57336 9034
rect 56848 8994 57336 9000
rect 54392 8872 54398 8932
rect 54458 8872 54464 8932
rect 55530 8872 55536 8932
rect 55596 8872 55602 8932
rect 54280 8672 54286 8732
rect 54346 8672 54352 8732
rect 54174 8570 54180 8630
rect 54240 8570 54246 8630
rect 54064 5118 54070 5178
rect 54130 5118 54136 5178
rect 54180 5140 54240 8570
rect 54286 7496 54346 8672
rect 54280 7436 54286 7496
rect 54346 7436 54352 7496
rect 53832 4968 53838 5028
rect 53898 4968 53904 5028
rect 54070 1442 54130 5118
rect 54174 5080 54180 5140
rect 54240 5080 54246 5140
rect 54180 2650 54240 5080
rect 54286 2776 54346 7436
rect 54398 6158 54458 8872
rect 55528 8672 55534 8732
rect 55594 8672 55600 8732
rect 55534 8628 55594 8672
rect 54518 8568 55594 8628
rect 54518 8566 55082 8568
rect 54518 8426 54578 8566
rect 55022 8516 55082 8566
rect 54812 8510 55300 8516
rect 54812 8476 54824 8510
rect 55288 8476 55300 8510
rect 54812 8470 55300 8476
rect 54518 8394 54530 8426
rect 54524 7850 54530 8394
rect 54564 8394 54578 8426
rect 55534 8426 55594 8568
rect 56038 8516 56098 8994
rect 56546 8792 56552 8852
rect 56612 8792 56618 8852
rect 55830 8510 56318 8516
rect 55830 8476 55842 8510
rect 56306 8476 56318 8510
rect 55830 8470 56318 8476
rect 54564 7850 54570 8394
rect 55534 8390 55548 8426
rect 54524 7838 54570 7850
rect 55542 7850 55548 8390
rect 55582 8390 55594 8426
rect 56552 8426 56612 8792
rect 57066 8738 57126 8994
rect 57570 8956 57630 9084
rect 58596 9084 58602 9630
rect 58636 9630 58650 9660
rect 59604 9660 59664 10036
rect 60110 9750 60170 10228
rect 60620 10140 60626 10200
rect 60686 10140 60692 10200
rect 59902 9744 60390 9750
rect 59902 9710 59914 9744
rect 60378 9710 60390 9744
rect 59902 9704 60390 9710
rect 58636 9084 58642 9630
rect 59604 9616 59620 9660
rect 59614 9134 59620 9616
rect 58596 9072 58642 9084
rect 59606 9084 59620 9134
rect 59654 9616 59664 9660
rect 60626 9660 60686 10140
rect 62662 10096 62722 10318
rect 63688 10318 63694 10842
rect 63728 10850 63742 10894
rect 63728 10842 63738 10850
rect 64694 10846 64712 10894
rect 63728 10318 63734 10842
rect 64706 10366 64712 10846
rect 63688 10306 63734 10318
rect 64700 10318 64712 10366
rect 64746 10846 64754 10894
rect 65714 10854 65730 10894
rect 64746 10366 64752 10846
rect 64746 10318 64760 10366
rect 62958 10268 63446 10274
rect 62958 10234 62970 10268
rect 63434 10234 63446 10268
rect 62958 10228 63446 10234
rect 63976 10268 64464 10274
rect 63976 10234 63988 10268
rect 64452 10234 64464 10268
rect 63976 10228 64464 10234
rect 64700 10096 64760 10318
rect 65724 10318 65730 10854
rect 65764 10856 65780 10894
rect 65764 10854 65778 10856
rect 65764 10318 65770 10854
rect 66730 10848 66748 10894
rect 66742 10372 66748 10848
rect 66730 10318 66748 10372
rect 66782 10848 66790 10894
rect 67752 10894 67812 11136
rect 68246 10984 68306 11242
rect 68048 10978 68536 10984
rect 68048 10944 68060 10978
rect 68524 10944 68536 10978
rect 68048 10938 68536 10944
rect 68768 10894 68828 11352
rect 69278 11302 69338 11460
rect 70292 11302 70352 11460
rect 70806 11412 70866 11550
rect 71822 11550 71838 11606
rect 71872 12086 71884 12126
rect 71872 11606 71878 12086
rect 71872 11550 71882 11606
rect 71102 11500 71590 11506
rect 71102 11466 71114 11500
rect 71578 11466 71590 11500
rect 71102 11460 71590 11466
rect 70800 11352 70806 11412
rect 70866 11352 70872 11412
rect 69272 11242 69278 11302
rect 69338 11242 69344 11302
rect 70286 11242 70292 11302
rect 70352 11242 70358 11302
rect 69278 10984 69338 11242
rect 69786 11136 69792 11196
rect 69852 11136 69858 11196
rect 69066 10978 69554 10984
rect 69066 10944 69078 10978
rect 69542 10944 69554 10978
rect 69066 10938 69554 10944
rect 69792 10894 69852 11136
rect 70292 10984 70352 11242
rect 70084 10978 70572 10984
rect 70084 10944 70096 10978
rect 70560 10944 70572 10978
rect 70084 10938 70572 10944
rect 66782 10372 66788 10848
rect 67752 10842 67766 10894
rect 66782 10318 66790 10372
rect 67760 10318 67766 10842
rect 67800 10852 67816 10894
rect 67800 10842 67812 10852
rect 67800 10318 67806 10842
rect 65724 10306 65770 10318
rect 66742 10306 66788 10318
rect 67760 10306 67806 10318
rect 68768 10318 68784 10894
rect 68818 10318 68828 10894
rect 69788 10852 69802 10894
rect 69792 10832 69802 10852
rect 64994 10268 65482 10274
rect 64994 10234 65006 10268
rect 65470 10234 65482 10268
rect 64994 10228 65482 10234
rect 66012 10268 66500 10274
rect 66012 10234 66024 10268
rect 66488 10234 66500 10268
rect 66012 10228 66500 10234
rect 67030 10268 67518 10274
rect 67030 10234 67042 10268
rect 67506 10234 67518 10268
rect 67030 10228 67518 10234
rect 68048 10268 68536 10274
rect 68048 10234 68060 10268
rect 68524 10234 68536 10268
rect 68048 10228 68536 10234
rect 66726 10140 66732 10200
rect 66792 10140 66798 10200
rect 62656 10036 62662 10096
rect 62722 10036 62728 10096
rect 64694 10036 64700 10096
rect 64760 10036 64766 10096
rect 61640 9914 61646 9974
rect 61706 9914 61712 9974
rect 63674 9914 63680 9974
rect 63740 9914 63746 9974
rect 65704 9914 65710 9974
rect 65770 9914 65776 9974
rect 60920 9744 61408 9750
rect 60920 9710 60932 9744
rect 61396 9710 61408 9744
rect 60920 9704 61408 9710
rect 59654 9134 59660 9616
rect 60626 9598 60638 9660
rect 59654 9084 59666 9134
rect 60632 9120 60638 9598
rect 57866 9034 58354 9040
rect 57866 9000 57878 9034
rect 58342 9000 58354 9034
rect 57866 8994 58354 9000
rect 58884 9034 59372 9040
rect 58884 9000 58896 9034
rect 59360 9000 59372 9034
rect 58884 8994 59372 9000
rect 57564 8896 57570 8956
rect 57630 8896 57636 8956
rect 57060 8678 57066 8738
rect 57126 8678 57132 8738
rect 57066 8516 57126 8678
rect 56848 8510 57336 8516
rect 56848 8476 56860 8510
rect 57324 8476 57336 8510
rect 56848 8470 57336 8476
rect 55582 7850 55588 8390
rect 56552 8384 56566 8426
rect 56560 7908 56566 8384
rect 55542 7838 55588 7850
rect 56554 7850 56566 7908
rect 56600 8384 56612 8426
rect 57570 8426 57630 8896
rect 58068 8744 58128 8994
rect 58586 8792 58592 8852
rect 58652 8792 58658 8852
rect 58068 8738 58130 8744
rect 58068 8678 58070 8738
rect 58068 8672 58130 8678
rect 58068 8516 58128 8672
rect 57866 8510 58354 8516
rect 57866 8476 57878 8510
rect 58342 8476 58354 8510
rect 57866 8470 58354 8476
rect 56600 7908 56606 8384
rect 57570 8382 57584 8426
rect 56600 7850 56614 7908
rect 57578 7898 57584 8382
rect 54812 7800 55300 7806
rect 54812 7766 54824 7800
rect 55288 7766 55300 7800
rect 54812 7760 55300 7766
rect 55830 7800 56318 7806
rect 55830 7766 55842 7800
rect 56306 7766 56318 7800
rect 55830 7760 56318 7766
rect 55528 7640 55534 7700
rect 55594 7640 55600 7700
rect 54812 7278 55300 7284
rect 54812 7244 54824 7278
rect 55288 7244 55300 7278
rect 54812 7238 55300 7244
rect 54524 7194 54570 7206
rect 54524 6664 54530 7194
rect 54514 6618 54530 6664
rect 54564 6664 54570 7194
rect 55534 7194 55594 7640
rect 56040 7598 56100 7760
rect 56034 7538 56040 7598
rect 56100 7538 56106 7598
rect 56554 7396 56614 7850
rect 57572 7850 57584 7898
rect 57618 8382 57630 8426
rect 58592 8426 58652 8792
rect 59084 8744 59144 8994
rect 59606 8956 59666 9084
rect 60624 9084 60638 9120
rect 60672 9598 60686 9660
rect 61646 9660 61706 9914
rect 61938 9744 62426 9750
rect 61938 9710 61950 9744
rect 62414 9710 62426 9744
rect 61938 9704 62426 9710
rect 62956 9744 63444 9750
rect 62956 9710 62968 9744
rect 63432 9710 63444 9744
rect 62956 9704 63444 9710
rect 61646 9604 61656 9660
rect 60672 9120 60678 9598
rect 60672 9084 60684 9120
rect 59902 9034 60390 9040
rect 59902 9000 59914 9034
rect 60378 9000 60390 9034
rect 59902 8994 60390 9000
rect 59600 8896 59606 8956
rect 59666 8896 59672 8956
rect 59082 8738 59144 8744
rect 59142 8678 59144 8738
rect 59082 8672 59144 8678
rect 59084 8516 59144 8672
rect 58884 8510 59372 8516
rect 58884 8476 58896 8510
rect 59360 8476 59372 8510
rect 58884 8470 59372 8476
rect 58592 8384 58602 8426
rect 57618 7898 57624 8382
rect 57618 7850 57632 7898
rect 56848 7800 57336 7806
rect 56848 7766 56860 7800
rect 57324 7766 57336 7800
rect 56848 7760 57336 7766
rect 57572 7700 57632 7850
rect 58596 7850 58602 8384
rect 58636 8384 58652 8426
rect 59606 8426 59666 8896
rect 60102 8738 60162 8994
rect 60624 8852 60684 9084
rect 61650 9084 61656 9604
rect 61690 9604 61706 9660
rect 62668 9660 62714 9672
rect 61690 9084 61696 9604
rect 62668 9114 62674 9660
rect 61650 9072 61696 9084
rect 62658 9084 62674 9114
rect 62708 9114 62714 9660
rect 63680 9660 63740 9914
rect 63974 9744 64462 9750
rect 63974 9710 63986 9744
rect 64450 9710 64462 9744
rect 63974 9704 64462 9710
rect 64992 9744 65480 9750
rect 64992 9710 65004 9744
rect 65468 9710 65480 9744
rect 64992 9704 65480 9710
rect 63680 9610 63692 9660
rect 62708 9084 62718 9114
rect 60920 9034 61408 9040
rect 60920 9000 60932 9034
rect 61396 9000 61408 9034
rect 60920 8994 61408 9000
rect 61938 9034 62426 9040
rect 61938 9000 61950 9034
rect 62414 9000 62426 9034
rect 61938 8994 62426 9000
rect 60618 8792 60624 8852
rect 60684 8792 60690 8852
rect 61114 8796 61174 8994
rect 62156 8796 62216 8994
rect 62658 8852 62718 9084
rect 63686 9084 63692 9610
rect 63726 9610 63740 9660
rect 64704 9660 64750 9672
rect 63726 9084 63732 9610
rect 64704 9126 64710 9660
rect 63686 9072 63732 9084
rect 64698 9084 64710 9126
rect 64744 9126 64750 9660
rect 65710 9660 65770 9914
rect 66010 9744 66498 9750
rect 66010 9710 66022 9744
rect 66486 9710 66498 9744
rect 66010 9704 66498 9710
rect 65710 9616 65728 9660
rect 64744 9084 64758 9126
rect 62956 9034 63444 9040
rect 62956 9000 62968 9034
rect 63432 9000 63444 9034
rect 62956 8994 63444 9000
rect 63974 9034 64462 9040
rect 63974 9000 63986 9034
rect 64450 9000 64462 9034
rect 63974 8994 64462 9000
rect 60618 8680 60624 8740
rect 60684 8680 60690 8740
rect 61114 8736 62216 8796
rect 62652 8792 62658 8852
rect 62718 8792 62724 8852
rect 60102 8516 60162 8678
rect 59902 8510 60390 8516
rect 59902 8476 59914 8510
rect 60378 8476 60390 8510
rect 59902 8470 60390 8476
rect 58636 7850 58642 8384
rect 59606 8378 59620 8426
rect 59614 7900 59620 8378
rect 58596 7838 58642 7850
rect 59608 7850 59620 7900
rect 59654 8378 59666 8426
rect 60624 8426 60684 8680
rect 61114 8516 61174 8736
rect 61636 8570 61642 8630
rect 61702 8570 61708 8630
rect 60920 8510 61408 8516
rect 60920 8476 60932 8510
rect 61396 8476 61408 8510
rect 60920 8470 61408 8476
rect 59654 7900 59660 8378
rect 60624 8368 60638 8426
rect 59654 7850 59668 7900
rect 57866 7800 58354 7806
rect 57866 7766 57878 7800
rect 58342 7766 58354 7800
rect 57866 7760 58354 7766
rect 58884 7800 59372 7806
rect 58884 7766 58896 7800
rect 59360 7766 59372 7800
rect 58884 7760 59372 7766
rect 57566 7640 57572 7700
rect 57632 7640 57638 7700
rect 57564 7436 57570 7496
rect 57630 7436 57636 7496
rect 58078 7490 58138 7760
rect 59100 7490 59160 7760
rect 59608 7700 59668 7850
rect 60632 7850 60638 8368
rect 60672 8368 60684 8426
rect 61642 8426 61702 8570
rect 62156 8516 62216 8736
rect 62654 8680 62660 8740
rect 62720 8680 62726 8740
rect 61938 8510 62426 8516
rect 61938 8476 61950 8510
rect 62414 8476 62426 8510
rect 61938 8470 62426 8476
rect 61642 8380 61656 8426
rect 60672 7850 60678 8368
rect 60632 7838 60678 7850
rect 61650 7850 61656 8380
rect 61690 8380 61702 8426
rect 62660 8426 62720 8680
rect 63156 8516 63216 8994
rect 63670 8570 63676 8630
rect 63736 8570 63742 8630
rect 62956 8510 63444 8516
rect 62956 8476 62968 8510
rect 63432 8476 63444 8510
rect 62956 8470 63444 8476
rect 61690 7850 61696 8380
rect 62660 8358 62674 8426
rect 61650 7838 61696 7850
rect 62668 7850 62674 8358
rect 62708 8358 62720 8426
rect 63676 8426 63736 8570
rect 64190 8516 64250 8994
rect 64698 8852 64758 9084
rect 65722 9084 65728 9616
rect 65762 9616 65770 9660
rect 66732 9660 66792 10140
rect 67254 9750 67314 10228
rect 67744 10036 67750 10096
rect 67810 10036 67816 10096
rect 67028 9744 67516 9750
rect 67028 9710 67040 9744
rect 67504 9710 67516 9744
rect 67028 9704 67516 9710
rect 65762 9084 65768 9616
rect 66732 9608 66746 9660
rect 66740 9136 66746 9608
rect 65722 9072 65768 9084
rect 66732 9084 66746 9136
rect 66780 9608 66792 9660
rect 67750 9660 67810 10036
rect 68256 9750 68316 10228
rect 68768 10096 68828 10318
rect 69796 10318 69802 10832
rect 69836 10832 69852 10894
rect 70806 10894 70866 11352
rect 71310 11302 71370 11460
rect 71304 11242 71310 11302
rect 71370 11242 71376 11302
rect 71310 10984 71370 11242
rect 71822 11196 71882 11550
rect 72842 11550 72856 12126
rect 72890 12094 72904 12126
rect 73862 12098 73874 12126
rect 72890 11550 72902 12094
rect 73866 12062 73874 12098
rect 73868 11610 73874 12062
rect 72120 11500 72608 11506
rect 72120 11466 72132 11500
rect 72596 11466 72608 11500
rect 72120 11460 72608 11466
rect 72334 11302 72394 11460
rect 72842 11412 72902 11550
rect 73862 11550 73874 11610
rect 73908 12062 73926 12126
rect 74886 12126 74932 12138
rect 73908 11610 73914 12062
rect 73908 11550 73922 11610
rect 74886 11598 74892 12126
rect 73138 11500 73626 11506
rect 73138 11466 73150 11500
rect 73614 11466 73626 11500
rect 73138 11460 73626 11466
rect 72836 11352 72842 11412
rect 72902 11352 72908 11412
rect 72328 11242 72334 11302
rect 72394 11242 72400 11302
rect 71816 11136 71822 11196
rect 71882 11136 71888 11196
rect 71816 11032 71822 11092
rect 71882 11032 71888 11092
rect 71102 10978 71590 10984
rect 71102 10944 71114 10978
rect 71578 10944 71590 10978
rect 71102 10938 71590 10944
rect 71302 10926 71362 10938
rect 71822 10894 71882 11032
rect 72334 10984 72394 11242
rect 72120 10978 72608 10984
rect 72120 10944 72132 10978
rect 72596 10944 72608 10978
rect 72120 10938 72608 10944
rect 70806 10836 70820 10894
rect 69836 10318 69842 10832
rect 70814 10366 70820 10836
rect 69796 10306 69842 10318
rect 70804 10318 70820 10366
rect 70854 10836 70866 10894
rect 71820 10848 71838 10894
rect 70854 10366 70860 10836
rect 71822 10820 71838 10848
rect 71832 10372 71838 10820
rect 70854 10318 70864 10366
rect 69066 10268 69554 10274
rect 69066 10234 69078 10268
rect 69542 10234 69554 10268
rect 69066 10228 69554 10234
rect 70084 10268 70572 10274
rect 70084 10234 70096 10268
rect 70560 10234 70572 10268
rect 70084 10228 70572 10234
rect 68762 10036 68768 10096
rect 68828 10036 68834 10096
rect 69268 9750 69328 10228
rect 69782 10036 69788 10096
rect 69848 10036 69854 10096
rect 68046 9744 68534 9750
rect 68046 9710 68058 9744
rect 68522 9710 68534 9744
rect 68046 9704 68534 9710
rect 69064 9744 69552 9750
rect 69064 9710 69076 9744
rect 69540 9710 69552 9744
rect 69064 9704 69552 9710
rect 67750 9612 67764 9660
rect 66780 9136 66786 9608
rect 66780 9084 66792 9136
rect 67758 9116 67764 9612
rect 64992 9034 65480 9040
rect 64992 9000 65004 9034
rect 65468 9000 65480 9034
rect 64992 8994 65480 9000
rect 66010 9034 66498 9040
rect 66010 9000 66022 9034
rect 66486 9000 66498 9034
rect 66010 8994 66498 9000
rect 64692 8792 64698 8852
rect 64758 8792 64764 8852
rect 65212 8796 65272 8994
rect 66220 8796 66280 8994
rect 66732 8852 66792 9084
rect 67750 9084 67764 9116
rect 67798 9612 67810 9660
rect 68776 9660 68822 9672
rect 67798 9116 67804 9612
rect 68776 9120 68782 9660
rect 67798 9084 67810 9116
rect 67028 9034 67516 9040
rect 67028 9000 67040 9034
rect 67504 9000 67516 9034
rect 67028 8994 67516 9000
rect 64690 8680 64696 8740
rect 64756 8680 64762 8740
rect 65212 8736 66280 8796
rect 66726 8792 66732 8852
rect 66792 8792 66798 8852
rect 66922 8788 66928 8848
rect 66988 8788 66994 8848
rect 63974 8510 64462 8516
rect 63974 8476 63986 8510
rect 64450 8476 64462 8510
rect 63974 8470 64462 8476
rect 63676 8378 63692 8426
rect 62708 7850 62714 8358
rect 62668 7838 62714 7850
rect 63686 7850 63692 8378
rect 63726 8378 63736 8426
rect 64696 8426 64756 8680
rect 65212 8516 65272 8736
rect 65710 8570 65716 8630
rect 65776 8570 65782 8630
rect 64992 8510 65480 8516
rect 64992 8476 65004 8510
rect 65468 8476 65480 8510
rect 64992 8470 65480 8476
rect 63726 7850 63732 8378
rect 64696 8376 64710 8426
rect 63686 7838 63732 7850
rect 64704 7850 64710 8376
rect 64744 8376 64756 8426
rect 65716 8426 65776 8570
rect 66220 8516 66280 8736
rect 66726 8680 66732 8740
rect 66792 8680 66798 8740
rect 66010 8510 66498 8516
rect 66010 8476 66022 8510
rect 66486 8476 66498 8510
rect 66010 8470 66498 8476
rect 65716 8388 65728 8426
rect 64744 7850 64750 8376
rect 65722 7896 65728 8388
rect 64704 7838 64750 7850
rect 65716 7850 65728 7896
rect 65762 8388 65776 8426
rect 66732 8426 66792 8680
rect 66928 8630 66988 8788
rect 67222 8632 67282 8994
rect 67750 8956 67810 9084
rect 68766 9084 68782 9120
rect 68816 9120 68822 9660
rect 69788 9660 69848 10036
rect 70302 9750 70362 10228
rect 70804 10096 70864 10318
rect 71826 10318 71838 10372
rect 71872 10820 71882 10894
rect 72842 10894 72902 11352
rect 73354 11302 73414 11460
rect 73862 11402 73922 11550
rect 74878 11550 74892 11598
rect 74926 11598 74932 12126
rect 74926 11550 74938 11598
rect 74156 11500 74644 11506
rect 74156 11466 74168 11500
rect 74632 11466 74644 11500
rect 74156 11460 74644 11466
rect 74372 11402 74432 11460
rect 74878 11402 74938 11550
rect 74998 11402 75058 12274
rect 73862 11342 75058 11402
rect 73348 11242 73354 11302
rect 73414 11242 73420 11302
rect 73354 10984 73414 11242
rect 73856 11136 73862 11196
rect 73922 11136 73928 11196
rect 73862 11094 73922 11136
rect 73862 11034 74940 11094
rect 74998 11092 75058 11342
rect 73138 10978 73626 10984
rect 73138 10944 73150 10978
rect 73614 10944 73626 10978
rect 73138 10938 73626 10944
rect 72842 10868 72856 10894
rect 71872 10372 71878 10820
rect 72850 10376 72856 10868
rect 71872 10318 71886 10372
rect 71102 10268 71590 10274
rect 71102 10234 71114 10268
rect 71578 10234 71590 10268
rect 71102 10228 71590 10234
rect 71826 10200 71886 10318
rect 72840 10318 72856 10376
rect 72890 10868 72902 10894
rect 73862 10894 73922 11034
rect 74348 10984 74408 11034
rect 74156 10978 74644 10984
rect 74156 10944 74168 10978
rect 74632 10944 74644 10978
rect 74156 10938 74644 10944
rect 74880 10894 74940 11034
rect 74992 11032 74998 11092
rect 75058 11032 75064 11092
rect 72890 10376 72896 10868
rect 73862 10838 73874 10894
rect 72890 10318 72900 10376
rect 72120 10268 72608 10274
rect 72120 10234 72132 10268
rect 72596 10234 72608 10268
rect 72120 10228 72608 10234
rect 71820 10140 71826 10200
rect 71886 10140 71892 10200
rect 72840 10096 72900 10318
rect 73868 10318 73874 10838
rect 73908 10838 73922 10894
rect 74876 10858 74892 10894
rect 74880 10852 74892 10858
rect 73908 10318 73914 10838
rect 74886 10362 74892 10852
rect 73868 10306 73914 10318
rect 74882 10318 74892 10362
rect 74926 10852 74940 10894
rect 74926 10362 74932 10852
rect 74926 10318 74942 10362
rect 73138 10268 73626 10274
rect 73138 10234 73150 10268
rect 73614 10234 73626 10268
rect 73138 10228 73626 10234
rect 74156 10268 74644 10274
rect 74156 10234 74168 10268
rect 74632 10234 74644 10268
rect 74156 10228 74644 10234
rect 70798 10036 70804 10096
rect 70864 10036 70870 10096
rect 72834 10036 72840 10096
rect 72900 10036 72906 10096
rect 73330 9750 73390 10228
rect 74882 10192 74942 10318
rect 74882 10132 75172 10192
rect 74368 9826 74936 9886
rect 74368 9750 74428 9826
rect 70082 9744 70570 9750
rect 70082 9710 70094 9744
rect 70558 9710 70570 9744
rect 70082 9704 70570 9710
rect 71100 9744 71588 9750
rect 71100 9710 71112 9744
rect 71576 9710 71588 9744
rect 71100 9704 71588 9710
rect 72118 9744 72606 9750
rect 72118 9710 72130 9744
rect 72594 9710 72606 9744
rect 72118 9704 72606 9710
rect 73136 9744 73624 9750
rect 73136 9710 73148 9744
rect 73612 9710 73624 9744
rect 73136 9704 73624 9710
rect 74154 9744 74642 9750
rect 74154 9710 74166 9744
rect 74630 9710 74642 9744
rect 74154 9704 74642 9710
rect 69788 9602 69800 9660
rect 69794 9130 69800 9602
rect 68816 9084 68826 9120
rect 68046 9034 68534 9040
rect 68046 9000 68058 9034
rect 68522 9000 68534 9034
rect 68046 8994 68534 9000
rect 67744 8896 67750 8956
rect 67810 8896 67816 8956
rect 66922 8570 66928 8630
rect 66988 8570 66994 8630
rect 67216 8572 67222 8632
rect 67282 8572 67288 8632
rect 67222 8516 67282 8572
rect 67028 8510 67516 8516
rect 67028 8476 67040 8510
rect 67504 8476 67516 8510
rect 67028 8470 67516 8476
rect 65762 7896 65768 8388
rect 66732 8382 66746 8426
rect 65762 7850 65776 7896
rect 59902 7800 60390 7806
rect 59902 7766 59914 7800
rect 60378 7766 60390 7800
rect 59902 7760 60390 7766
rect 60920 7800 61408 7806
rect 60920 7766 60932 7800
rect 61396 7766 61408 7800
rect 60920 7760 61408 7766
rect 61938 7800 62426 7806
rect 61938 7766 61950 7800
rect 62414 7766 62426 7800
rect 61938 7760 62426 7766
rect 62956 7800 63444 7806
rect 62956 7766 62968 7800
rect 63432 7766 63444 7800
rect 62956 7760 63444 7766
rect 63974 7800 64462 7806
rect 63974 7766 63986 7800
rect 64450 7766 64462 7800
rect 63974 7760 64462 7766
rect 64992 7800 65480 7806
rect 64992 7766 65004 7800
rect 65468 7766 65480 7800
rect 64992 7760 65480 7766
rect 59602 7640 59608 7700
rect 59668 7640 59674 7700
rect 56548 7336 56554 7396
rect 56614 7336 56620 7396
rect 55830 7278 56318 7284
rect 55830 7244 55842 7278
rect 56306 7244 56318 7278
rect 55830 7238 56318 7244
rect 55534 7156 55548 7194
rect 54564 6618 54574 6664
rect 55542 6660 55548 7156
rect 54514 6456 54574 6618
rect 55532 6618 55548 6660
rect 55582 7156 55594 7194
rect 56554 7194 56614 7336
rect 56848 7278 57336 7284
rect 56848 7244 56860 7278
rect 57324 7244 57336 7278
rect 56848 7238 57336 7244
rect 55582 6660 55588 7156
rect 56554 7154 56566 7194
rect 55582 6618 55592 6660
rect 54812 6568 55300 6574
rect 54812 6534 54824 6568
rect 55288 6534 55300 6568
rect 54812 6528 55300 6534
rect 55026 6456 55086 6528
rect 55532 6456 55592 6618
rect 56560 6618 56566 7154
rect 56600 7154 56614 7194
rect 57570 7194 57630 7436
rect 58072 7430 58078 7490
rect 58138 7430 58144 7490
rect 59094 7430 59100 7490
rect 59160 7430 59166 7490
rect 58582 7336 58588 7396
rect 58648 7336 58654 7396
rect 57866 7278 58354 7284
rect 57866 7244 57878 7278
rect 58342 7244 58354 7278
rect 57866 7238 58354 7244
rect 56600 6618 56606 7154
rect 57570 7142 57584 7194
rect 56560 6606 56606 6618
rect 57578 6618 57584 7142
rect 57618 7142 57630 7194
rect 58588 7194 58648 7336
rect 59100 7284 59160 7430
rect 58884 7278 59372 7284
rect 58884 7244 58896 7278
rect 59360 7244 59372 7278
rect 58884 7238 59372 7244
rect 58588 7150 58602 7194
rect 57618 6618 57624 7142
rect 58596 6654 58602 7150
rect 57578 6606 57624 6618
rect 58588 6618 58602 6654
rect 58636 7150 58648 7194
rect 59608 7194 59668 7640
rect 60114 7490 60174 7760
rect 61132 7598 61192 7760
rect 62152 7710 62212 7760
rect 63152 7710 63212 7760
rect 64190 7710 64250 7760
rect 65218 7710 65278 7760
rect 61634 7640 61640 7700
rect 61700 7640 61706 7700
rect 62152 7650 65278 7710
rect 61126 7538 61132 7598
rect 61192 7538 61198 7598
rect 60108 7430 60114 7490
rect 60174 7430 60180 7490
rect 61126 7430 61132 7490
rect 61192 7430 61198 7490
rect 60114 7284 60174 7430
rect 60618 7336 60624 7396
rect 60684 7336 60690 7396
rect 59902 7278 60390 7284
rect 59902 7244 59914 7278
rect 60378 7244 60390 7278
rect 59902 7238 60390 7244
rect 58636 6654 58642 7150
rect 58636 6618 58648 6654
rect 55830 6568 56318 6574
rect 55830 6534 55842 6568
rect 56306 6534 56318 6568
rect 55830 6528 56318 6534
rect 56848 6568 57336 6574
rect 56848 6534 56860 6568
rect 57324 6534 57336 6568
rect 56848 6528 57336 6534
rect 57866 6568 58354 6574
rect 57866 6534 57878 6568
rect 58342 6534 58354 6568
rect 57866 6528 58354 6534
rect 56036 6472 56096 6528
rect 54514 6396 55592 6456
rect 56030 6412 56036 6472
rect 56096 6412 56102 6472
rect 56940 6412 56946 6472
rect 57006 6412 57012 6472
rect 56030 6196 56036 6256
rect 56096 6196 56102 6256
rect 56036 6190 56098 6196
rect 54398 6152 54460 6158
rect 54398 6092 54400 6152
rect 54398 6086 54460 6092
rect 54398 3908 54458 6086
rect 56038 6050 56098 6190
rect 56946 6050 57006 6412
rect 57074 6256 57134 6528
rect 57942 6412 57948 6472
rect 58008 6412 58014 6472
rect 57074 6190 57134 6196
rect 57948 6050 58008 6412
rect 58088 6256 58148 6528
rect 58588 6370 58648 6618
rect 59608 6618 59620 7194
rect 59654 6618 59668 7194
rect 60624 7194 60684 7336
rect 61132 7284 61192 7430
rect 60920 7278 61408 7284
rect 60920 7244 60932 7278
rect 61396 7244 61408 7278
rect 60920 7238 61408 7244
rect 60624 7158 60638 7194
rect 58884 6568 59372 6574
rect 58884 6534 58896 6568
rect 59360 6534 59372 6568
rect 58884 6528 59372 6534
rect 59100 6472 59160 6528
rect 59094 6412 59100 6472
rect 59160 6412 59166 6472
rect 58582 6310 58588 6370
rect 58648 6310 58654 6370
rect 58082 6196 58088 6256
rect 58148 6196 58154 6256
rect 59100 6050 59160 6412
rect 54812 6044 55300 6050
rect 54812 6010 54824 6044
rect 55288 6010 55300 6044
rect 54812 6004 55300 6010
rect 55830 6044 56318 6050
rect 55830 6010 55842 6044
rect 56306 6010 56318 6044
rect 55830 6004 56318 6010
rect 56848 6044 57336 6050
rect 56848 6010 56860 6044
rect 57324 6010 57336 6044
rect 56848 6004 57336 6010
rect 57866 6044 58354 6050
rect 57866 6010 57878 6044
rect 58342 6010 58354 6044
rect 57866 6004 58354 6010
rect 58884 6044 59372 6050
rect 58884 6010 58896 6044
rect 59360 6010 59372 6044
rect 58884 6004 59372 6010
rect 54524 5960 54570 5972
rect 54524 5422 54530 5960
rect 54518 5384 54530 5422
rect 54564 5422 54570 5960
rect 55542 5960 55588 5972
rect 55542 5422 55548 5960
rect 54564 5384 54578 5422
rect 54518 5254 54578 5384
rect 55536 5384 55548 5422
rect 55582 5422 55588 5960
rect 56560 5960 56606 5972
rect 56560 5434 56566 5960
rect 55582 5384 55596 5422
rect 54812 5334 55300 5340
rect 54812 5300 54824 5334
rect 55288 5300 55300 5334
rect 54812 5294 55300 5300
rect 55016 5254 55076 5294
rect 55536 5254 55596 5384
rect 56552 5384 56566 5434
rect 56600 5434 56606 5960
rect 57578 5960 57624 5972
rect 57578 5442 57584 5960
rect 56600 5384 56612 5434
rect 55830 5334 56318 5340
rect 55830 5300 55842 5334
rect 56306 5300 56318 5334
rect 55830 5294 56318 5300
rect 54518 5194 55596 5254
rect 55536 5140 55596 5194
rect 56028 5184 56034 5244
rect 56094 5184 56100 5244
rect 55530 5080 55536 5140
rect 55596 5080 55602 5140
rect 55526 4870 55532 4930
rect 55592 4870 55598 4930
rect 54812 4810 55300 4816
rect 54812 4776 54824 4810
rect 55288 4776 55300 4810
rect 54812 4770 55300 4776
rect 54524 4726 54570 4738
rect 54524 4184 54530 4726
rect 54514 4150 54530 4184
rect 54564 4184 54570 4726
rect 55532 4726 55592 4870
rect 56034 4816 56094 5184
rect 56552 5028 56612 5384
rect 57570 5384 57584 5442
rect 57618 5442 57624 5960
rect 58596 5960 58642 5972
rect 57618 5384 57630 5442
rect 58596 5430 58602 5960
rect 56848 5334 57336 5340
rect 56848 5300 56860 5334
rect 57324 5300 57336 5334
rect 56848 5294 57336 5300
rect 57042 5244 57102 5294
rect 57036 5184 57042 5244
rect 57102 5184 57108 5244
rect 56546 4968 56552 5028
rect 56612 4968 56618 5028
rect 57570 4930 57630 5384
rect 58590 5384 58602 5430
rect 58636 5430 58642 5960
rect 59608 5960 59668 6618
rect 60632 6618 60638 7158
rect 60672 7158 60684 7194
rect 61640 7194 61700 7640
rect 62146 7430 62152 7490
rect 62212 7430 62218 7490
rect 65218 7474 65278 7650
rect 65716 7584 65776 7850
rect 66740 7850 66746 8382
rect 66780 8382 66792 8426
rect 67750 8426 67810 8896
rect 68252 8638 68312 8994
rect 68766 8740 68826 9084
rect 69786 9084 69800 9130
rect 69834 9602 69848 9660
rect 70812 9660 70858 9672
rect 69834 9130 69840 9602
rect 70812 9140 70818 9660
rect 69834 9084 69846 9130
rect 69064 9034 69552 9040
rect 69064 9000 69076 9034
rect 69540 9000 69552 9034
rect 69064 8994 69552 9000
rect 68760 8680 68766 8740
rect 68826 8680 68832 8740
rect 68250 8632 68312 8638
rect 68310 8572 68312 8632
rect 68250 8566 68312 8572
rect 68762 8566 68768 8626
rect 68828 8566 68834 8626
rect 68252 8516 68312 8566
rect 68046 8510 68534 8516
rect 68046 8476 68058 8510
rect 68522 8476 68534 8510
rect 68046 8470 68534 8476
rect 67750 8382 67764 8426
rect 66780 7850 66786 8382
rect 66740 7838 66786 7850
rect 67758 7850 67764 8382
rect 67798 8382 67810 8426
rect 68768 8426 68828 8566
rect 69276 8516 69336 8994
rect 69786 8956 69846 9084
rect 70804 9084 70818 9140
rect 70852 9140 70858 9660
rect 71830 9660 71876 9672
rect 70852 9084 70864 9140
rect 71830 9128 71836 9660
rect 70082 9034 70570 9040
rect 70082 9000 70094 9034
rect 70558 9000 70570 9034
rect 70082 8994 70570 9000
rect 69780 8896 69786 8956
rect 69846 8896 69852 8956
rect 69064 8510 69552 8516
rect 69064 8476 69076 8510
rect 69540 8476 69552 8510
rect 69064 8470 69552 8476
rect 68768 8396 68782 8426
rect 67798 7850 67804 8382
rect 68776 7890 68782 8396
rect 67758 7838 67804 7850
rect 68768 7850 68782 7890
rect 68816 8396 68828 8426
rect 69786 8426 69846 8896
rect 70302 8516 70362 8994
rect 70804 8740 70864 9084
rect 71820 9084 71836 9128
rect 71870 9128 71876 9660
rect 72848 9660 72894 9672
rect 72848 9128 72854 9660
rect 71870 9084 71880 9128
rect 71100 9034 71588 9040
rect 71100 9000 71112 9034
rect 71576 9000 71588 9034
rect 71100 8994 71588 9000
rect 70798 8680 70804 8740
rect 70864 8680 70870 8740
rect 71310 8690 71370 8994
rect 71820 8848 71880 9084
rect 72844 9084 72854 9128
rect 72888 9128 72894 9660
rect 73866 9660 73912 9672
rect 73866 9134 73872 9660
rect 72888 9084 72904 9128
rect 72118 9034 72606 9040
rect 72118 9000 72130 9034
rect 72594 9000 72606 9034
rect 72118 8994 72606 9000
rect 72326 8850 72386 8994
rect 71814 8788 71820 8848
rect 71880 8788 71886 8848
rect 72324 8844 72386 8850
rect 72384 8784 72386 8844
rect 72324 8778 72386 8784
rect 72326 8690 72386 8778
rect 72844 8740 72904 9084
rect 73860 9084 73872 9134
rect 73906 9134 73912 9660
rect 74876 9660 74936 9826
rect 74978 9802 74984 9862
rect 75044 9802 75050 9862
rect 75112 9844 75172 10132
rect 74876 9632 74890 9660
rect 74884 9142 74890 9632
rect 73906 9084 73920 9134
rect 73136 9034 73624 9040
rect 73136 9000 73148 9034
rect 73612 9000 73624 9034
rect 73136 8994 73624 9000
rect 71310 8630 72386 8690
rect 72838 8680 72844 8740
rect 72904 8680 72910 8740
rect 70798 8566 70804 8626
rect 70864 8566 70870 8626
rect 70082 8510 70570 8516
rect 70082 8476 70094 8510
rect 70558 8476 70570 8510
rect 70082 8470 70570 8476
rect 68816 7890 68822 8396
rect 69786 8386 69800 8426
rect 68816 7850 68828 7890
rect 69794 7884 69800 8386
rect 66010 7800 66498 7806
rect 66010 7766 66022 7800
rect 66486 7766 66498 7800
rect 66010 7760 66498 7766
rect 67028 7800 67516 7806
rect 67028 7766 67040 7800
rect 67504 7766 67516 7800
rect 67028 7760 67516 7766
rect 68046 7800 68534 7806
rect 68046 7766 68058 7800
rect 68522 7766 68534 7800
rect 68046 7760 68534 7766
rect 66222 7712 66282 7760
rect 65710 7524 65716 7584
rect 65776 7524 65782 7584
rect 66222 7474 66282 7652
rect 62152 7284 62212 7430
rect 65218 7414 66282 7474
rect 67746 7326 67752 7386
rect 67812 7326 67818 7386
rect 61938 7278 62426 7284
rect 61938 7244 61950 7278
rect 62414 7244 62426 7278
rect 61938 7238 62426 7244
rect 62956 7278 63444 7284
rect 62956 7244 62968 7278
rect 63432 7244 63444 7278
rect 62956 7238 63444 7244
rect 63974 7278 64462 7284
rect 63974 7244 63986 7278
rect 64450 7244 64462 7278
rect 63974 7238 64462 7244
rect 64992 7278 65480 7284
rect 64992 7244 65004 7278
rect 65468 7244 65480 7278
rect 64992 7238 65480 7244
rect 66010 7278 66498 7284
rect 66010 7244 66022 7278
rect 66486 7244 66498 7278
rect 66010 7238 66498 7244
rect 67028 7278 67516 7284
rect 67028 7244 67040 7278
rect 67504 7244 67516 7278
rect 67028 7238 67516 7244
rect 60672 6618 60678 7158
rect 61640 7156 61656 7194
rect 60632 6606 60678 6618
rect 61650 6618 61656 7156
rect 61690 7156 61700 7194
rect 62668 7194 62714 7206
rect 61690 6618 61696 7156
rect 62668 6660 62674 7194
rect 61650 6606 61696 6618
rect 62660 6618 62674 6660
rect 62708 6660 62714 7194
rect 63686 7194 63732 7206
rect 62708 6618 62720 6660
rect 63686 6656 63692 7194
rect 59902 6568 60390 6574
rect 59902 6534 59914 6568
rect 60378 6534 60390 6568
rect 59902 6528 60390 6534
rect 60920 6568 61408 6574
rect 60920 6534 60932 6568
rect 61396 6534 61408 6568
rect 60920 6528 61408 6534
rect 61938 6568 62426 6574
rect 61938 6534 61950 6568
rect 62414 6534 62426 6568
rect 61938 6528 62426 6534
rect 60110 6472 60170 6528
rect 61116 6472 61176 6528
rect 62160 6472 62220 6528
rect 62660 6478 62720 6618
rect 63680 6618 63692 6656
rect 63726 6656 63732 7194
rect 64704 7194 64750 7206
rect 63726 6618 63740 6656
rect 64704 6650 64710 7194
rect 62956 6568 63444 6574
rect 62956 6534 62968 6568
rect 63432 6534 63444 6568
rect 62956 6528 63444 6534
rect 60104 6412 60110 6472
rect 60170 6412 60176 6472
rect 61110 6412 61116 6472
rect 61176 6412 61182 6472
rect 62154 6412 62160 6472
rect 62220 6412 62226 6472
rect 62654 6418 62660 6478
rect 62720 6418 62726 6478
rect 60110 6050 60170 6412
rect 61108 6196 61114 6256
rect 61174 6196 61180 6256
rect 62148 6196 62154 6256
rect 62214 6196 62220 6256
rect 61114 6050 61174 6196
rect 61632 6092 61638 6152
rect 61698 6092 61704 6152
rect 59902 6044 60390 6050
rect 59902 6010 59914 6044
rect 60378 6010 60390 6044
rect 59902 6004 60390 6010
rect 60920 6044 61408 6050
rect 60920 6010 60932 6044
rect 61396 6010 61408 6044
rect 60920 6004 61408 6010
rect 59608 5878 59620 5960
rect 59614 5430 59620 5878
rect 58636 5384 58650 5430
rect 57866 5334 58354 5340
rect 57866 5300 57878 5334
rect 58342 5300 58354 5334
rect 57866 5294 58354 5300
rect 58056 5244 58116 5294
rect 58050 5184 58056 5244
rect 58116 5184 58122 5244
rect 58590 5028 58650 5384
rect 59610 5384 59620 5430
rect 59654 5878 59668 5960
rect 60632 5960 60678 5972
rect 59654 5430 59660 5878
rect 59654 5384 59670 5430
rect 60632 5428 60638 5960
rect 58884 5334 59372 5340
rect 58884 5300 58896 5334
rect 59360 5300 59372 5334
rect 58884 5294 59372 5300
rect 59094 5244 59154 5294
rect 59088 5184 59094 5244
rect 59154 5184 59160 5244
rect 58584 4968 58590 5028
rect 58650 4968 58656 5028
rect 57564 4870 57570 4930
rect 57630 4870 57636 4930
rect 59094 4816 59154 5184
rect 59610 4930 59670 5384
rect 60628 5384 60638 5428
rect 60672 5428 60678 5960
rect 61638 5960 61698 6092
rect 62154 6050 62214 6196
rect 61938 6044 62426 6050
rect 61938 6010 61950 6044
rect 62414 6010 62426 6044
rect 61938 6004 62426 6010
rect 61638 5896 61656 5960
rect 60672 5384 60688 5428
rect 59902 5334 60390 5340
rect 59902 5300 59914 5334
rect 60378 5300 60390 5334
rect 59902 5294 60390 5300
rect 60112 5244 60172 5294
rect 60628 5250 60688 5384
rect 61650 5384 61656 5896
rect 61690 5896 61698 5960
rect 62660 5960 62720 6418
rect 63168 6256 63228 6528
rect 63162 6196 63168 6256
rect 63228 6196 63234 6256
rect 63168 6050 63228 6196
rect 63680 6152 63740 6618
rect 64696 6618 64710 6650
rect 64744 6650 64750 7194
rect 65722 7194 65768 7206
rect 65722 6652 65728 7194
rect 64744 6618 64756 6650
rect 63974 6568 64462 6574
rect 63974 6534 63986 6568
rect 64450 6534 64462 6568
rect 63974 6528 64462 6534
rect 64176 6256 64236 6528
rect 64696 6478 64756 6618
rect 65718 6618 65728 6652
rect 65762 6652 65768 7194
rect 66740 7194 66786 7206
rect 65762 6618 65778 6652
rect 66740 6650 66746 7194
rect 64992 6568 65480 6574
rect 64992 6534 65004 6568
rect 65468 6534 65480 6568
rect 64992 6528 65480 6534
rect 64690 6418 64696 6478
rect 64756 6418 64762 6478
rect 65220 6256 65280 6528
rect 64170 6196 64176 6256
rect 64236 6196 64242 6256
rect 65214 6196 65220 6256
rect 65280 6196 65286 6256
rect 63674 6092 63680 6152
rect 63740 6092 63746 6152
rect 62956 6044 63444 6050
rect 62956 6010 62968 6044
rect 63432 6010 63444 6044
rect 62956 6004 63444 6010
rect 62660 5924 62674 5960
rect 61690 5384 61696 5896
rect 62668 5442 62674 5924
rect 61650 5372 61696 5384
rect 62664 5384 62674 5442
rect 62708 5924 62720 5960
rect 63680 5960 63740 6092
rect 64176 6050 64236 6196
rect 65220 6050 65280 6196
rect 65718 6152 65778 6618
rect 66732 6618 66746 6650
rect 66780 6650 66786 7194
rect 67752 7194 67812 7326
rect 68046 7278 68534 7284
rect 68046 7244 68058 7278
rect 68522 7244 68534 7278
rect 68046 7238 68534 7244
rect 66780 6618 66792 6650
rect 66010 6568 66498 6574
rect 66010 6534 66022 6568
rect 66486 6534 66498 6568
rect 66010 6528 66498 6534
rect 66210 6256 66270 6528
rect 66732 6478 66792 6618
rect 67752 6618 67764 7194
rect 67798 6618 67812 7194
rect 68768 7194 68828 7850
rect 69788 7850 69800 7884
rect 69834 8386 69846 8426
rect 70804 8426 70864 8566
rect 71310 8516 71370 8630
rect 72326 8516 72386 8630
rect 72836 8566 72842 8626
rect 72902 8566 72908 8626
rect 71100 8510 71588 8516
rect 71100 8476 71112 8510
rect 71576 8476 71588 8510
rect 71100 8470 71588 8476
rect 72118 8510 72606 8516
rect 72118 8476 72130 8510
rect 72594 8476 72606 8510
rect 72118 8470 72606 8476
rect 69834 7884 69840 8386
rect 70804 8384 70818 8426
rect 69834 7850 69848 7884
rect 69064 7800 69552 7806
rect 69064 7766 69076 7800
rect 69540 7766 69552 7800
rect 69064 7760 69552 7766
rect 69264 7490 69324 7760
rect 69258 7430 69264 7490
rect 69324 7430 69330 7490
rect 69264 7284 69324 7430
rect 69064 7278 69552 7284
rect 69064 7244 69076 7278
rect 69540 7244 69552 7278
rect 69064 7238 69552 7244
rect 68768 7154 68782 7194
rect 68776 6650 68782 7154
rect 67028 6568 67516 6574
rect 67028 6534 67040 6568
rect 67504 6534 67516 6568
rect 67028 6528 67516 6534
rect 66726 6418 66732 6478
rect 66792 6418 66798 6478
rect 67228 6256 67288 6528
rect 66204 6196 66210 6256
rect 66270 6196 66276 6256
rect 67222 6196 67228 6256
rect 67288 6196 67294 6256
rect 65712 6092 65718 6152
rect 65778 6092 65784 6152
rect 63974 6044 64462 6050
rect 63974 6010 63986 6044
rect 64450 6010 64462 6044
rect 63974 6004 64462 6010
rect 64992 6044 65480 6050
rect 64992 6010 65004 6044
rect 65468 6010 65480 6044
rect 64992 6004 65480 6010
rect 62708 5442 62714 5924
rect 63680 5922 63692 5960
rect 62708 5384 62724 5442
rect 60920 5334 61408 5340
rect 60920 5300 60932 5334
rect 61396 5300 61408 5334
rect 60920 5294 61408 5300
rect 61938 5334 62426 5340
rect 61938 5300 61950 5334
rect 62414 5300 62426 5334
rect 61938 5294 62426 5300
rect 62664 5250 62724 5384
rect 63686 5384 63692 5922
rect 63726 5922 63740 5960
rect 64704 5960 64750 5972
rect 63726 5384 63732 5922
rect 64704 5434 64710 5960
rect 63686 5372 63732 5384
rect 64696 5384 64710 5434
rect 64744 5434 64750 5960
rect 65718 5960 65778 6092
rect 66210 6050 66270 6196
rect 67752 6152 67812 6618
rect 68770 6618 68782 6650
rect 68816 7154 68828 7194
rect 69788 7194 69848 7850
rect 70812 7850 70818 8384
rect 70852 8384 70864 8426
rect 71830 8426 71876 8438
rect 70852 7850 70858 8384
rect 71830 7908 71836 8426
rect 70812 7838 70858 7850
rect 71822 7850 71836 7908
rect 71870 7908 71876 8426
rect 72842 8426 72902 8566
rect 73344 8516 73404 8994
rect 73860 8956 73920 9084
rect 74878 9084 74890 9142
rect 74924 9632 74936 9660
rect 74924 9142 74930 9632
rect 74924 9084 74938 9142
rect 74154 9034 74642 9040
rect 74154 9000 74166 9034
rect 74630 9000 74642 9034
rect 74154 8994 74642 9000
rect 74878 8974 74938 9084
rect 73854 8896 73860 8956
rect 73920 8896 73926 8956
rect 74872 8914 74878 8974
rect 74938 8914 74944 8974
rect 73860 8678 73920 8896
rect 73860 8618 74934 8678
rect 74984 8626 75044 9802
rect 75106 9784 75112 9844
rect 75172 9784 75178 9844
rect 75478 8844 75538 12730
rect 75472 8784 75478 8844
rect 75538 8784 75544 8844
rect 75222 8680 75228 8740
rect 75288 8680 75294 8740
rect 73136 8510 73624 8516
rect 73136 8476 73148 8510
rect 73612 8476 73624 8510
rect 73136 8470 73624 8476
rect 72842 8384 72854 8426
rect 71870 7850 71882 7908
rect 70294 7806 70354 7808
rect 70082 7800 70570 7806
rect 70082 7766 70094 7800
rect 70558 7766 70570 7800
rect 70082 7760 70570 7766
rect 71100 7800 71588 7806
rect 71100 7766 71112 7800
rect 71576 7766 71588 7800
rect 71100 7760 71588 7766
rect 70294 7490 70354 7760
rect 71316 7712 71376 7760
rect 71310 7652 71316 7712
rect 71376 7652 71382 7712
rect 71448 7656 71454 7716
rect 71514 7656 71520 7716
rect 71454 7490 71514 7656
rect 71822 7490 71882 7850
rect 72848 7850 72854 8384
rect 72888 8384 72902 8426
rect 73860 8426 73920 8618
rect 74364 8516 74424 8618
rect 74154 8510 74642 8516
rect 74154 8476 74166 8510
rect 74630 8476 74642 8510
rect 74154 8470 74642 8476
rect 73860 8392 73872 8426
rect 72888 7850 72894 8384
rect 73866 7890 73872 8392
rect 72848 7838 72894 7850
rect 73860 7850 73872 7890
rect 73906 8392 73920 8426
rect 74874 8426 74934 8618
rect 74978 8566 74984 8626
rect 75044 8566 75050 8626
rect 74874 8402 74890 8426
rect 73906 7890 73912 8392
rect 73906 7850 73920 7890
rect 72118 7800 72606 7806
rect 72118 7766 72130 7800
rect 72594 7766 72606 7800
rect 72118 7760 72606 7766
rect 73136 7800 73624 7806
rect 73136 7766 73148 7800
rect 73612 7766 73624 7800
rect 73136 7760 73624 7766
rect 73342 7716 73402 7760
rect 72330 7656 72336 7716
rect 72396 7656 72402 7716
rect 73336 7656 73342 7716
rect 73402 7656 73408 7716
rect 73860 7712 73920 7850
rect 74884 7850 74890 8402
rect 74924 8402 74934 8426
rect 74924 7850 74930 8402
rect 74884 7838 74930 7850
rect 74154 7800 74642 7806
rect 74154 7766 74166 7800
rect 74630 7766 74642 7800
rect 74154 7760 74642 7766
rect 70288 7430 70294 7490
rect 70354 7430 70360 7490
rect 71448 7430 71454 7490
rect 71514 7430 71520 7490
rect 71816 7430 71822 7490
rect 71882 7430 71888 7490
rect 70294 7284 70354 7430
rect 71454 7284 71514 7430
rect 71822 7386 71882 7430
rect 71816 7326 71822 7386
rect 71882 7326 71888 7386
rect 72336 7284 72396 7656
rect 73854 7652 73860 7712
rect 73920 7652 73926 7712
rect 73854 7524 73860 7584
rect 73920 7524 73926 7584
rect 72832 7328 72838 7388
rect 72898 7328 72904 7388
rect 70082 7278 70570 7284
rect 70082 7244 70094 7278
rect 70558 7244 70570 7278
rect 70082 7238 70570 7244
rect 71100 7278 71588 7284
rect 71100 7244 71112 7278
rect 71576 7244 71588 7278
rect 71100 7238 71588 7244
rect 72118 7278 72606 7284
rect 72118 7244 72130 7278
rect 72594 7244 72606 7278
rect 72118 7238 72606 7244
rect 72336 7236 72396 7238
rect 68816 6650 68822 7154
rect 69788 7148 69800 7194
rect 69794 6662 69800 7148
rect 68816 6618 68830 6650
rect 68046 6568 68534 6574
rect 68046 6534 68058 6568
rect 68522 6534 68534 6568
rect 68046 6528 68534 6534
rect 68262 6256 68322 6528
rect 68770 6478 68830 6618
rect 69786 6618 69800 6662
rect 69834 7148 69848 7194
rect 70812 7194 70858 7206
rect 69834 6662 69840 7148
rect 69834 6618 69846 6662
rect 70812 6658 70818 7194
rect 69064 6568 69552 6574
rect 69064 6534 69076 6568
rect 69540 6534 69552 6568
rect 69064 6528 69552 6534
rect 68764 6418 68770 6478
rect 68830 6418 68836 6478
rect 68756 6310 68762 6370
rect 68822 6310 68828 6370
rect 68256 6196 68262 6256
rect 68322 6196 68328 6256
rect 67746 6092 67752 6152
rect 67812 6092 67818 6152
rect 68258 6088 68264 6148
rect 68324 6088 68330 6148
rect 68264 6050 68324 6088
rect 66010 6044 66498 6050
rect 66010 6010 66022 6044
rect 66486 6010 66498 6044
rect 66010 6004 66498 6010
rect 67028 6044 67516 6050
rect 67028 6010 67040 6044
rect 67504 6010 67516 6044
rect 67028 6004 67516 6010
rect 68046 6044 68534 6050
rect 68046 6010 68058 6044
rect 68522 6010 68534 6044
rect 68046 6004 68534 6010
rect 65718 5924 65728 5960
rect 64744 5384 64756 5434
rect 62956 5334 63444 5340
rect 62956 5300 62968 5334
rect 63432 5300 63444 5334
rect 62956 5294 63444 5300
rect 63974 5334 64462 5340
rect 63974 5300 63986 5334
rect 64450 5300 64462 5334
rect 63974 5294 64462 5300
rect 64696 5250 64756 5384
rect 65722 5384 65728 5924
rect 65762 5924 65778 5960
rect 66740 5960 66786 5972
rect 65762 5384 65768 5924
rect 66740 5446 66746 5960
rect 65722 5372 65768 5384
rect 66730 5384 66746 5446
rect 66780 5446 66786 5960
rect 67758 5960 67804 5972
rect 66780 5384 66790 5446
rect 67758 5426 67764 5960
rect 64992 5334 65480 5340
rect 64992 5300 65004 5334
rect 65468 5300 65480 5334
rect 64992 5294 65480 5300
rect 66010 5334 66498 5340
rect 66010 5300 66022 5334
rect 66486 5300 66498 5334
rect 66010 5294 66498 5300
rect 66730 5250 66790 5384
rect 67752 5384 67764 5426
rect 67798 5426 67804 5960
rect 68762 5960 68822 6310
rect 69286 6148 69346 6528
rect 69786 6154 69846 6618
rect 70806 6618 70818 6658
rect 70852 6658 70858 7194
rect 71830 7194 71876 7206
rect 71830 6662 71836 7194
rect 70852 6618 70866 6658
rect 70082 6568 70570 6574
rect 70082 6534 70094 6568
rect 70558 6534 70570 6568
rect 70082 6528 70570 6534
rect 69280 6088 69286 6148
rect 69346 6088 69352 6148
rect 69780 6094 69786 6154
rect 69846 6094 69852 6154
rect 69286 6050 69346 6088
rect 69064 6044 69552 6050
rect 69064 6010 69076 6044
rect 69540 6010 69552 6044
rect 69064 6004 69552 6010
rect 68762 5924 68782 5960
rect 67798 5384 67812 5426
rect 67028 5334 67516 5340
rect 67028 5300 67040 5334
rect 67504 5300 67516 5334
rect 67028 5294 67516 5300
rect 60106 5184 60112 5244
rect 60172 5184 60178 5244
rect 60622 5190 60628 5250
rect 60688 5190 60694 5250
rect 64690 5190 64696 5250
rect 64756 5190 64762 5250
rect 66724 5190 66730 5250
rect 66790 5190 66796 5250
rect 59604 4870 59610 4930
rect 59670 4870 59676 4930
rect 55830 4810 56318 4816
rect 55830 4776 55842 4810
rect 56306 4776 56318 4810
rect 55830 4770 56318 4776
rect 56848 4810 57336 4816
rect 56848 4776 56860 4810
rect 57324 4776 57336 4810
rect 56848 4770 57336 4776
rect 57866 4810 58354 4816
rect 57866 4776 57878 4810
rect 58342 4776 58354 4810
rect 57866 4770 58354 4776
rect 58884 4810 59372 4816
rect 58884 4776 58896 4810
rect 59360 4776 59372 4810
rect 58884 4770 59372 4776
rect 55532 4672 55548 4726
rect 54564 4150 54574 4184
rect 55542 4180 55548 4672
rect 54514 4018 54574 4150
rect 55538 4150 55548 4180
rect 55582 4672 55592 4726
rect 56560 4726 56606 4738
rect 55582 4180 55588 4672
rect 56560 4196 56566 4726
rect 55582 4150 55598 4180
rect 54812 4100 55300 4106
rect 54812 4066 54824 4100
rect 55288 4066 55300 4100
rect 54812 4060 55300 4066
rect 55034 4018 55094 4060
rect 55538 4018 55598 4150
rect 56552 4150 56566 4196
rect 56600 4196 56606 4726
rect 57578 4726 57624 4738
rect 56600 4150 56612 4196
rect 57578 4180 57584 4726
rect 55830 4100 56318 4106
rect 55830 4066 55842 4100
rect 56306 4066 56318 4100
rect 55830 4060 56318 4066
rect 54514 3958 55598 4018
rect 54392 3848 54398 3908
rect 54458 3848 54464 3908
rect 55538 3812 55598 3958
rect 54514 3752 55598 3812
rect 54514 3494 54574 3752
rect 55026 3584 55086 3752
rect 55538 3692 55598 3752
rect 55532 3632 55538 3692
rect 55598 3632 55604 3692
rect 54812 3578 55300 3584
rect 54812 3544 54824 3578
rect 55288 3544 55300 3578
rect 54812 3538 55300 3544
rect 54514 3458 54530 3494
rect 54524 2918 54530 3458
rect 54564 3458 54574 3494
rect 55538 3494 55598 3632
rect 56030 3584 56090 4060
rect 56552 4006 56612 4150
rect 57570 4150 57584 4180
rect 57618 4180 57624 4726
rect 58596 4726 58642 4738
rect 58596 4192 58602 4726
rect 57618 4150 57630 4180
rect 56848 4100 57336 4106
rect 56848 4066 56860 4100
rect 57324 4066 57336 4100
rect 56848 4060 57336 4066
rect 56546 3946 56552 4006
rect 56612 3946 56618 4006
rect 56550 3752 56556 3812
rect 56616 3752 56622 3812
rect 55830 3578 56318 3584
rect 55830 3544 55842 3578
rect 56306 3544 56318 3578
rect 55830 3538 56318 3544
rect 54564 2918 54570 3458
rect 55538 3454 55548 3494
rect 54524 2906 54570 2918
rect 55542 2918 55548 3454
rect 55582 3454 55598 3494
rect 56556 3494 56616 3752
rect 57050 3748 57110 4060
rect 57570 3908 57630 4150
rect 58588 4150 58602 4192
rect 58636 4192 58642 4726
rect 59610 4726 59670 4870
rect 60112 4816 60172 5184
rect 59902 4810 60390 4816
rect 59902 4776 59914 4810
rect 60378 4776 60390 4810
rect 59902 4770 60390 4776
rect 59610 4696 59620 4726
rect 59614 4214 59620 4696
rect 58636 4150 58648 4192
rect 57866 4100 58354 4106
rect 57866 4066 57878 4100
rect 58342 4066 58354 4100
rect 57866 4060 58354 4066
rect 57564 3848 57570 3908
rect 57630 3848 57636 3908
rect 58084 3748 58144 4060
rect 58588 4006 58648 4150
rect 59606 4150 59620 4214
rect 59654 4696 59670 4726
rect 60628 4726 60688 5190
rect 62664 5184 62724 5190
rect 63674 5080 63680 5140
rect 63740 5080 63746 5140
rect 65710 5080 65716 5140
rect 65776 5080 65782 5140
rect 62656 4968 62662 5028
rect 62722 4968 62728 5028
rect 61640 4870 61646 4930
rect 61706 4870 61712 4930
rect 60920 4810 61408 4816
rect 60920 4776 60932 4810
rect 61396 4776 61408 4810
rect 60920 4770 61408 4776
rect 59654 4214 59660 4696
rect 60628 4684 60638 4726
rect 59654 4150 59666 4214
rect 60632 4190 60638 4684
rect 58884 4100 59372 4106
rect 58884 4066 58896 4100
rect 59360 4066 59372 4100
rect 58884 4060 59372 4066
rect 58582 3946 58588 4006
rect 58648 3946 58654 4006
rect 59094 3908 59154 4060
rect 59088 3848 59094 3908
rect 59154 3848 59160 3908
rect 58586 3752 58592 3812
rect 58652 3752 58658 3812
rect 57050 3688 58144 3748
rect 57050 3584 57110 3688
rect 58084 3584 58144 3688
rect 56848 3578 57336 3584
rect 56848 3544 56860 3578
rect 57324 3544 57336 3578
rect 56848 3538 57336 3544
rect 57866 3578 58354 3584
rect 57866 3544 57878 3578
rect 58342 3544 58354 3578
rect 57866 3538 58354 3544
rect 55582 2918 55588 3454
rect 56556 3450 56566 3494
rect 55542 2906 55588 2918
rect 56560 2918 56566 3450
rect 56600 3450 56616 3494
rect 57578 3494 57624 3506
rect 56600 2918 56606 3450
rect 57578 2960 57584 3494
rect 56560 2906 56606 2918
rect 57570 2918 57584 2960
rect 57618 2960 57624 3494
rect 58592 3494 58652 3752
rect 59094 3584 59154 3848
rect 59606 3692 59666 4150
rect 60626 4150 60638 4190
rect 60672 4684 60688 4726
rect 61646 4726 61706 4870
rect 61938 4810 62426 4816
rect 61938 4776 61950 4810
rect 62414 4776 62426 4810
rect 61938 4770 62426 4776
rect 61646 4690 61656 4726
rect 60672 4190 60678 4684
rect 60672 4150 60686 4190
rect 61650 4184 61656 4690
rect 59902 4100 60390 4106
rect 59902 4066 59914 4100
rect 60378 4066 60390 4100
rect 59902 4060 60390 4066
rect 60116 3908 60176 4060
rect 60626 4006 60686 4150
rect 61640 4150 61656 4184
rect 61690 4690 61706 4726
rect 62662 4726 62722 4968
rect 62956 4810 63444 4816
rect 62956 4776 62968 4810
rect 63432 4776 63444 4810
rect 62956 4770 63444 4776
rect 62662 4700 62674 4726
rect 61690 4184 61696 4690
rect 62668 4206 62674 4700
rect 61690 4150 61700 4184
rect 60920 4100 61408 4106
rect 60920 4066 60932 4100
rect 61396 4066 61408 4100
rect 60920 4060 61408 4066
rect 60620 3946 60626 4006
rect 60686 3946 60692 4006
rect 61140 3914 61200 4060
rect 59600 3632 59606 3692
rect 59666 3632 59672 3692
rect 58884 3578 59372 3584
rect 58884 3544 58896 3578
rect 59360 3544 59372 3578
rect 58884 3538 59372 3544
rect 58592 3442 58602 3494
rect 57618 2918 57630 2960
rect 54812 2868 55300 2874
rect 54812 2834 54824 2868
rect 55288 2834 55300 2868
rect 54812 2828 55300 2834
rect 55830 2868 56318 2874
rect 55830 2834 55842 2868
rect 56306 2834 56318 2868
rect 55830 2828 56318 2834
rect 56848 2868 57336 2874
rect 56848 2834 56860 2868
rect 57324 2834 57336 2868
rect 56848 2828 57336 2834
rect 54280 2716 54286 2776
rect 54346 2716 54352 2776
rect 54174 2590 54180 2650
rect 54240 2590 54246 2650
rect 54514 2410 55594 2470
rect 54514 2260 54574 2410
rect 55022 2350 55082 2410
rect 54812 2344 55300 2350
rect 54812 2310 54824 2344
rect 55288 2310 55300 2344
rect 54812 2304 55300 2310
rect 54514 2204 54530 2260
rect 54524 1684 54530 2204
rect 54564 2204 54574 2260
rect 55534 2260 55594 2410
rect 56032 2350 56092 2828
rect 57570 2650 57630 2918
rect 58596 2918 58602 3442
rect 58636 3442 58652 3494
rect 59606 3494 59666 3632
rect 60116 3584 60176 3848
rect 61138 3908 61200 3914
rect 61198 3848 61200 3908
rect 61138 3842 61200 3848
rect 60614 3752 60620 3812
rect 60680 3752 60686 3812
rect 59902 3578 60390 3584
rect 59902 3544 59914 3578
rect 60378 3544 60390 3578
rect 59902 3538 60390 3544
rect 59606 3454 59620 3494
rect 58636 2918 58642 3442
rect 59614 2972 59620 3454
rect 58596 2906 58642 2918
rect 59608 2918 59620 2972
rect 59654 3454 59666 3494
rect 60620 3494 60680 3752
rect 61140 3584 61200 3842
rect 61640 3692 61700 4150
rect 62658 4150 62674 4206
rect 62708 4700 62722 4726
rect 63680 4726 63740 5080
rect 63974 4810 64462 4816
rect 63974 4776 63986 4810
rect 64450 4776 64462 4810
rect 63974 4770 64462 4776
rect 64992 4810 65480 4816
rect 64992 4776 65004 4810
rect 65468 4776 65480 4810
rect 64992 4770 65480 4776
rect 62708 4206 62714 4700
rect 63680 4694 63692 4726
rect 62708 4150 62718 4206
rect 61938 4100 62426 4106
rect 61938 4066 61950 4100
rect 62414 4066 62426 4100
rect 61938 4060 62426 4066
rect 62142 3908 62202 4060
rect 62488 4026 62548 4032
rect 62658 4026 62718 4150
rect 63686 4150 63692 4694
rect 63726 4694 63740 4726
rect 64704 4726 64750 4738
rect 63726 4150 63732 4694
rect 64704 4220 64710 4726
rect 63686 4138 63732 4150
rect 64700 4150 64710 4220
rect 64744 4220 64750 4726
rect 65716 4726 65776 5080
rect 67258 5042 67318 5294
rect 67752 5252 67812 5384
rect 68776 5384 68782 5924
rect 68816 5384 68822 5960
rect 69786 5960 69846 6094
rect 70264 6050 70324 6528
rect 70806 6478 70866 6618
rect 71820 6618 71836 6662
rect 71870 6662 71876 7194
rect 72838 7194 72898 7328
rect 73136 7278 73624 7284
rect 73136 7244 73148 7278
rect 73612 7244 73624 7278
rect 73136 7238 73624 7244
rect 72838 7144 72854 7194
rect 71870 6618 71880 6662
rect 72848 6646 72854 7144
rect 71100 6568 71588 6574
rect 71100 6534 71112 6568
rect 71576 6534 71588 6568
rect 71100 6528 71588 6534
rect 70800 6418 70806 6478
rect 70866 6418 70872 6478
rect 70796 6310 70802 6370
rect 70862 6310 70868 6370
rect 70082 6044 70570 6050
rect 70082 6010 70094 6044
rect 70558 6010 70570 6044
rect 70082 6004 70570 6010
rect 69786 5866 69800 5960
rect 69794 5426 69800 5866
rect 68776 5372 68822 5384
rect 69786 5384 69800 5426
rect 69834 5866 69846 5960
rect 70802 5960 70862 6310
rect 71288 6196 71294 6256
rect 71354 6196 71360 6256
rect 71294 6050 71354 6196
rect 71820 6154 71880 6618
rect 72844 6618 72854 6646
rect 72888 7144 72898 7194
rect 73860 7194 73920 7524
rect 74154 7278 74642 7284
rect 74154 7244 74166 7278
rect 74630 7244 74642 7278
rect 74154 7238 74642 7244
rect 72888 6646 72894 7144
rect 73860 7142 73872 7194
rect 73866 6646 73872 7142
rect 72888 6618 72904 6646
rect 72118 6568 72606 6574
rect 72118 6534 72130 6568
rect 72594 6534 72606 6568
rect 72118 6528 72606 6534
rect 72844 6478 72904 6618
rect 73860 6618 73872 6646
rect 73906 7142 73920 7194
rect 74884 7194 74930 7206
rect 73906 6646 73912 7142
rect 74884 6652 74890 7194
rect 73906 6618 73920 6646
rect 73136 6568 73624 6574
rect 73136 6534 73148 6568
rect 73612 6534 73624 6568
rect 73136 6528 73624 6534
rect 72838 6418 72844 6478
rect 72904 6418 72910 6478
rect 72834 6310 72840 6370
rect 72900 6310 72906 6370
rect 72326 6196 72332 6256
rect 72392 6196 72398 6256
rect 71814 6094 71820 6154
rect 71880 6094 71886 6154
rect 72332 6050 72392 6196
rect 71100 6044 71588 6050
rect 71100 6010 71112 6044
rect 71576 6010 71588 6044
rect 71100 6004 71588 6010
rect 72118 6044 72606 6050
rect 72118 6010 72130 6044
rect 72594 6010 72606 6044
rect 72118 6004 72606 6010
rect 70802 5894 70818 5960
rect 69834 5426 69840 5866
rect 69834 5384 69846 5426
rect 68046 5334 68534 5340
rect 68046 5300 68058 5334
rect 68522 5300 68534 5334
rect 68046 5294 68534 5300
rect 69064 5334 69552 5340
rect 69064 5300 69076 5334
rect 69540 5300 69552 5334
rect 69064 5294 69552 5300
rect 67746 5192 67752 5252
rect 67812 5192 67818 5252
rect 68100 5192 68106 5252
rect 68166 5192 68172 5252
rect 67742 5080 67748 5140
rect 67808 5080 67814 5140
rect 67252 4982 67258 5042
rect 67318 4982 67324 5042
rect 66010 4810 66498 4816
rect 66010 4776 66022 4810
rect 66486 4776 66498 4810
rect 66010 4770 66498 4776
rect 67028 4810 67516 4816
rect 67028 4776 67040 4810
rect 67504 4776 67516 4810
rect 67028 4770 67516 4776
rect 65716 4688 65728 4726
rect 64744 4150 64760 4220
rect 62956 4100 63444 4106
rect 62956 4066 62968 4100
rect 63432 4066 63444 4100
rect 62956 4060 63444 4066
rect 63974 4100 64462 4106
rect 63974 4066 63986 4100
rect 64450 4066 64462 4100
rect 63974 4060 64462 4066
rect 62652 3966 62658 4026
rect 62718 3966 62724 4026
rect 62136 3848 62142 3908
rect 62202 3848 62208 3908
rect 61634 3632 61640 3692
rect 61700 3632 61706 3692
rect 60920 3578 61408 3584
rect 60920 3544 60932 3578
rect 61396 3544 61408 3578
rect 60920 3538 61408 3544
rect 59654 2972 59660 3454
rect 60620 3434 60638 3494
rect 59654 2918 59668 2972
rect 57866 2868 58354 2874
rect 57866 2834 57878 2868
rect 58342 2834 58354 2868
rect 57866 2828 58354 2834
rect 58884 2868 59372 2874
rect 58884 2834 58896 2868
rect 59360 2834 59372 2868
rect 58884 2828 59372 2834
rect 58090 2662 58150 2828
rect 57564 2590 57570 2650
rect 57630 2590 57636 2650
rect 58084 2602 58090 2662
rect 58150 2602 58156 2662
rect 56546 2488 56552 2548
rect 56612 2488 56618 2548
rect 58582 2488 58588 2548
rect 58648 2488 58654 2548
rect 55830 2344 56318 2350
rect 55830 2310 55842 2344
rect 56306 2310 56318 2344
rect 55830 2304 56318 2310
rect 54564 1684 54570 2204
rect 54524 1672 54570 1684
rect 55534 1684 55548 2260
rect 55582 1684 55594 2260
rect 56552 2260 56612 2488
rect 57564 2384 57570 2444
rect 57630 2384 57636 2444
rect 56848 2344 57336 2350
rect 56848 2310 56860 2344
rect 57324 2310 57336 2344
rect 56848 2304 57336 2310
rect 56552 2200 56566 2260
rect 56560 1720 56566 2200
rect 54812 1634 55300 1640
rect 54812 1600 54824 1634
rect 55288 1600 55300 1634
rect 54812 1594 55300 1600
rect 54392 1486 54398 1546
rect 54458 1486 54464 1546
rect 54064 1382 54070 1442
rect 54130 1382 54136 1442
rect 54398 1216 54458 1486
rect 55534 1442 55594 1684
rect 56554 1684 56566 1720
rect 56600 2200 56612 2260
rect 57570 2260 57630 2384
rect 57866 2344 58354 2350
rect 57866 2310 57878 2344
rect 58342 2310 58354 2344
rect 57866 2304 58354 2310
rect 57570 2206 57584 2260
rect 56600 1720 56606 2200
rect 57578 1724 57584 2206
rect 56600 1684 56614 1720
rect 55830 1634 56318 1640
rect 55830 1600 55842 1634
rect 56306 1600 56318 1634
rect 55830 1594 56318 1600
rect 55528 1382 55534 1442
rect 55594 1382 55600 1442
rect 56042 1336 56102 1594
rect 56036 1276 56042 1336
rect 56102 1276 56108 1336
rect 54398 1156 55598 1216
rect 53014 322 53020 382
rect 53080 322 53086 382
rect 54398 304 54458 1156
rect 54518 1028 54578 1156
rect 55004 1118 55064 1156
rect 54812 1112 55300 1118
rect 54812 1078 54824 1112
rect 55288 1078 55300 1112
rect 54812 1072 55300 1078
rect 54518 956 54530 1028
rect 54524 452 54530 956
rect 54564 956 54578 1028
rect 55538 1028 55598 1156
rect 56042 1118 56102 1276
rect 56554 1226 56614 1684
rect 57568 1684 57584 1724
rect 57618 2206 57630 2260
rect 58588 2260 58648 2488
rect 59090 2350 59150 2828
rect 59608 2548 59668 2918
rect 60632 2918 60638 3434
rect 60672 3434 60680 3494
rect 61640 3494 61700 3632
rect 62142 3584 62202 3848
rect 62488 3812 62548 3966
rect 62482 3752 62488 3812
rect 62548 3752 62554 3812
rect 62658 3758 62664 3818
rect 62724 3758 62730 3818
rect 61938 3578 62426 3584
rect 61938 3544 61950 3578
rect 62414 3544 62426 3578
rect 61938 3538 62426 3544
rect 61640 3454 61656 3494
rect 60672 2918 60678 3434
rect 61650 2984 61656 3454
rect 60632 2906 60678 2918
rect 61644 2918 61656 2984
rect 61690 3454 61700 3494
rect 62664 3494 62724 3758
rect 63180 3756 63240 4060
rect 64194 3920 64254 4060
rect 64700 4026 64760 4150
rect 65722 4150 65728 4688
rect 65762 4688 65776 4726
rect 66740 4726 66786 4738
rect 65762 4150 65768 4688
rect 66740 4220 66746 4726
rect 65722 4138 65768 4150
rect 66732 4150 66746 4220
rect 66780 4220 66786 4726
rect 67748 4726 67808 5080
rect 68106 4934 68166 5192
rect 68296 5042 68356 5294
rect 69272 5042 69332 5294
rect 68290 4982 68296 5042
rect 68356 4982 68362 5042
rect 69266 4982 69272 5042
rect 69332 4982 69338 5042
rect 69786 4930 69846 5384
rect 70812 5384 70818 5894
rect 70852 5894 70862 5960
rect 71830 5960 71876 5972
rect 70852 5384 70858 5894
rect 71830 5428 71836 5960
rect 70812 5372 70858 5384
rect 71824 5384 71836 5428
rect 71870 5428 71876 5960
rect 72840 5960 72900 6310
rect 73358 6256 73418 6528
rect 73860 6436 73920 6618
rect 74874 6618 74890 6652
rect 74924 6652 74930 7194
rect 74924 6618 74934 6652
rect 74154 6568 74642 6574
rect 74154 6534 74166 6568
rect 74630 6534 74642 6568
rect 74154 6528 74642 6534
rect 74368 6436 74428 6528
rect 74874 6436 74934 6618
rect 73860 6376 74934 6436
rect 73352 6196 73358 6256
rect 73418 6196 73424 6256
rect 73856 6094 73862 6154
rect 73922 6094 73928 6154
rect 73136 6044 73624 6050
rect 73136 6010 73148 6044
rect 73612 6010 73624 6044
rect 73136 6004 73624 6010
rect 72840 5908 72854 5960
rect 72848 5434 72854 5908
rect 71870 5384 71884 5428
rect 70082 5334 70570 5340
rect 70082 5300 70094 5334
rect 70558 5300 70570 5334
rect 70082 5294 70570 5300
rect 71100 5334 71588 5340
rect 71100 5300 71112 5334
rect 71576 5300 71588 5334
rect 71100 5294 71588 5300
rect 70288 5042 70348 5294
rect 71824 5252 71884 5384
rect 72842 5384 72854 5434
rect 72888 5908 72900 5960
rect 73862 5960 73922 6094
rect 74154 6044 74642 6050
rect 74154 6010 74166 6044
rect 74630 6010 74642 6044
rect 74154 6004 74642 6010
rect 73862 5926 73872 5960
rect 72888 5434 72894 5908
rect 72888 5384 72902 5434
rect 73866 5428 73872 5926
rect 72118 5334 72606 5340
rect 72118 5300 72130 5334
rect 72594 5300 72606 5334
rect 72118 5294 72606 5300
rect 71818 5192 71824 5252
rect 71884 5192 71890 5252
rect 70282 4982 70288 5042
rect 70348 4982 70354 5042
rect 72308 4982 72314 5042
rect 72374 4982 72380 5042
rect 68106 4868 68166 4874
rect 69780 4870 69786 4930
rect 69846 4870 69852 4930
rect 71816 4870 71822 4930
rect 71882 4870 71888 4930
rect 68046 4810 68534 4816
rect 68046 4776 68058 4810
rect 68522 4776 68534 4810
rect 68046 4770 68534 4776
rect 69064 4810 69552 4816
rect 69064 4776 69076 4810
rect 69540 4776 69552 4810
rect 69064 4770 69552 4776
rect 67748 4684 67764 4726
rect 66780 4150 66792 4220
rect 64992 4100 65480 4106
rect 64992 4066 65004 4100
rect 65468 4066 65480 4100
rect 64992 4060 65480 4066
rect 66010 4100 66498 4106
rect 66010 4066 66022 4100
rect 66486 4066 66498 4100
rect 66010 4060 66498 4066
rect 64694 3966 64700 4026
rect 64760 3966 64766 4026
rect 65216 3920 65276 4060
rect 66230 3920 66290 4060
rect 66732 4026 66792 4150
rect 67758 4150 67764 4684
rect 67798 4684 67808 4726
rect 68776 4726 68822 4738
rect 67798 4150 67804 4684
rect 68776 4186 68782 4726
rect 67758 4138 67804 4150
rect 68772 4150 68782 4186
rect 68816 4186 68822 4726
rect 69786 4726 69846 4870
rect 70082 4810 70570 4816
rect 70082 4776 70094 4810
rect 70558 4776 70570 4810
rect 70082 4770 70570 4776
rect 71100 4810 71588 4816
rect 71100 4776 71112 4810
rect 71576 4776 71588 4810
rect 71100 4770 71588 4776
rect 69786 4688 69800 4726
rect 69794 4202 69800 4688
rect 68816 4150 68832 4186
rect 67028 4100 67516 4106
rect 67028 4066 67040 4100
rect 67504 4066 67516 4100
rect 67028 4060 67516 4066
rect 68046 4100 68534 4106
rect 68046 4066 68058 4100
rect 68522 4066 68534 4100
rect 68046 4060 68534 4066
rect 66726 3966 66732 4026
rect 66792 3966 66798 4026
rect 67232 4020 67292 4060
rect 68258 4020 68318 4060
rect 68772 4026 68832 4150
rect 69790 4150 69800 4202
rect 69834 4688 69846 4726
rect 70812 4726 70858 4738
rect 69834 4202 69840 4688
rect 69834 4150 69850 4202
rect 70812 4194 70818 4726
rect 69064 4100 69552 4106
rect 69064 4066 69076 4100
rect 69540 4066 69552 4100
rect 69064 4060 69552 4066
rect 67232 3960 68318 4020
rect 68766 3966 68772 4026
rect 68832 3966 68838 4026
rect 67232 3920 67292 3960
rect 64194 3860 67292 3920
rect 67744 3868 67750 3928
rect 67810 3868 67816 3928
rect 64194 3756 64254 3860
rect 64686 3758 64692 3818
rect 64752 3758 64758 3818
rect 63180 3696 64254 3756
rect 63180 3584 63240 3696
rect 64194 3584 64254 3696
rect 62956 3578 63444 3584
rect 62956 3544 62968 3578
rect 63432 3544 63444 3578
rect 62956 3538 63444 3544
rect 63974 3578 64462 3584
rect 63974 3544 63986 3578
rect 64450 3544 64462 3578
rect 63974 3538 64462 3544
rect 61690 2984 61696 3454
rect 62664 3450 62674 3494
rect 61690 2918 61704 2984
rect 62668 2976 62674 3450
rect 59902 2868 60390 2874
rect 59902 2834 59914 2868
rect 60378 2834 60390 2868
rect 59902 2828 60390 2834
rect 60920 2868 61408 2874
rect 60920 2834 60932 2868
rect 61396 2834 61408 2868
rect 60920 2828 61408 2834
rect 59602 2488 59608 2548
rect 59668 2488 59674 2548
rect 60112 2350 60172 2828
rect 60618 2488 60624 2548
rect 60684 2488 60690 2548
rect 58884 2344 59372 2350
rect 58884 2310 58896 2344
rect 59360 2310 59372 2344
rect 58884 2304 59372 2310
rect 59902 2344 60390 2350
rect 59902 2310 59914 2344
rect 60378 2310 60390 2344
rect 59902 2304 60390 2310
rect 58588 2210 58602 2260
rect 57618 1724 57624 2206
rect 57618 1684 57628 1724
rect 58596 1708 58602 2210
rect 56848 1634 57336 1640
rect 56848 1600 56860 1634
rect 57324 1600 57336 1634
rect 56848 1594 57336 1600
rect 57062 1336 57122 1594
rect 57568 1546 57628 1684
rect 58590 1684 58602 1708
rect 58636 2210 58648 2260
rect 59614 2260 59660 2272
rect 58636 1708 58642 2210
rect 58636 1684 58650 1708
rect 59614 1698 59620 2260
rect 57866 1634 58354 1640
rect 57866 1600 57878 1634
rect 58342 1600 58354 1634
rect 57866 1594 58354 1600
rect 57562 1486 57568 1546
rect 57628 1486 57634 1546
rect 57568 1382 57574 1442
rect 57634 1382 57640 1442
rect 57056 1276 57062 1336
rect 57122 1276 57128 1336
rect 56548 1166 56554 1226
rect 56614 1166 56620 1226
rect 55830 1112 56318 1118
rect 55830 1078 55842 1112
rect 56306 1078 56318 1112
rect 55830 1072 56318 1078
rect 54564 452 54570 956
rect 55538 952 55548 1028
rect 55542 500 55548 952
rect 54524 440 54570 452
rect 55534 452 55548 500
rect 55582 952 55598 1028
rect 56554 1028 56614 1166
rect 57062 1118 57122 1276
rect 56848 1112 57336 1118
rect 56848 1078 56860 1112
rect 57324 1078 57336 1112
rect 56848 1072 57336 1078
rect 55582 500 55588 952
rect 55582 452 55594 500
rect 54812 402 55300 408
rect 54812 368 54824 402
rect 55288 368 55300 402
rect 54812 362 55300 368
rect 55534 304 55594 452
rect 56554 452 56566 1028
rect 56600 452 56614 1028
rect 57574 1028 57634 1382
rect 58086 1336 58146 1594
rect 58080 1276 58086 1336
rect 58146 1276 58152 1336
rect 58086 1118 58146 1276
rect 58590 1226 58650 1684
rect 59604 1684 59620 1698
rect 59654 1698 59660 2260
rect 60624 2260 60684 2488
rect 61124 2350 61184 2828
rect 61644 2548 61704 2918
rect 62656 2918 62674 2976
rect 62708 3450 62724 3494
rect 63686 3494 63732 3506
rect 62708 2976 62714 3450
rect 62708 2918 62716 2976
rect 63686 2970 63692 3494
rect 61938 2868 62426 2874
rect 61938 2834 61950 2868
rect 62414 2834 62426 2868
rect 61938 2828 62426 2834
rect 61638 2488 61644 2548
rect 61704 2488 61710 2548
rect 62154 2350 62214 2828
rect 62656 2716 62716 2918
rect 63674 2918 63692 2970
rect 63726 2970 63732 3494
rect 64692 3494 64752 3758
rect 65216 3584 65276 3860
rect 66230 3584 66290 3860
rect 66730 3758 66736 3818
rect 66796 3758 66802 3818
rect 64992 3578 65480 3584
rect 64992 3544 65004 3578
rect 65468 3544 65480 3578
rect 64992 3538 65480 3544
rect 66010 3578 66498 3584
rect 66010 3544 66022 3578
rect 66486 3544 66498 3578
rect 66010 3538 66498 3544
rect 64692 3450 64710 3494
rect 63726 2918 63734 2970
rect 62956 2868 63444 2874
rect 62956 2834 62968 2868
rect 63432 2834 63444 2868
rect 62956 2828 63444 2834
rect 62506 2656 62716 2716
rect 63170 2662 63230 2828
rect 63674 2776 63734 2918
rect 64704 2918 64710 3450
rect 64744 3450 64752 3494
rect 65722 3494 65768 3506
rect 64744 2918 64750 3450
rect 65722 2970 65728 3494
rect 64704 2906 64750 2918
rect 65716 2918 65728 2970
rect 65762 2970 65768 3494
rect 66736 3494 66796 3758
rect 67232 3584 67292 3860
rect 67028 3578 67516 3584
rect 67028 3544 67040 3578
rect 67504 3544 67516 3578
rect 67028 3538 67516 3544
rect 66736 3446 66746 3494
rect 65762 2918 65776 2970
rect 63974 2868 64462 2874
rect 63974 2834 63986 2868
rect 64450 2834 64462 2868
rect 63974 2828 64462 2834
rect 64992 2868 65480 2874
rect 64992 2834 65004 2868
rect 65468 2834 65480 2868
rect 64992 2828 65480 2834
rect 65716 2776 65776 2918
rect 66740 2918 66746 3446
rect 66780 3446 66796 3494
rect 67750 3494 67810 3868
rect 68258 3584 68318 3960
rect 68758 3758 68764 3818
rect 68824 3758 68830 3818
rect 68046 3578 68534 3584
rect 68046 3544 68058 3578
rect 68522 3544 68534 3578
rect 68046 3538 68534 3544
rect 67750 3458 67764 3494
rect 66780 2918 66786 3446
rect 67758 2962 67764 3458
rect 66740 2906 66786 2918
rect 67752 2918 67764 2962
rect 67798 3458 67810 3494
rect 68764 3494 68824 3758
rect 69278 3584 69338 4060
rect 69790 3692 69850 4150
rect 70802 4150 70818 4194
rect 70852 4194 70858 4726
rect 71822 4726 71882 4870
rect 72314 4816 72374 4982
rect 72118 4810 72606 4816
rect 72118 4776 72130 4810
rect 72594 4776 72606 4810
rect 72118 4770 72606 4776
rect 71822 4668 71836 4726
rect 70852 4150 70862 4194
rect 71830 4190 71836 4668
rect 70082 4100 70570 4106
rect 70082 4066 70094 4100
rect 70558 4066 70570 4100
rect 70082 4060 70570 4066
rect 69784 3632 69790 3692
rect 69850 3632 69856 3692
rect 69064 3578 69552 3584
rect 69064 3544 69076 3578
rect 69540 3544 69552 3578
rect 69064 3538 69552 3544
rect 67798 2962 67804 3458
rect 68764 3446 68782 3494
rect 67798 2918 67812 2962
rect 68776 2958 68782 3446
rect 66010 2868 66498 2874
rect 66010 2834 66022 2868
rect 66486 2834 66498 2868
rect 66010 2828 66498 2834
rect 67028 2868 67516 2874
rect 67028 2834 67040 2868
rect 67504 2834 67516 2868
rect 67028 2828 67516 2834
rect 67752 2776 67812 2918
rect 68766 2918 68782 2958
rect 68816 3446 68824 3494
rect 69790 3494 69850 3632
rect 70294 3584 70354 4060
rect 70802 3818 70862 4150
rect 71820 4150 71836 4190
rect 71870 4668 71882 4726
rect 72842 4726 72902 5384
rect 73858 5384 73872 5428
rect 73906 5926 73922 5960
rect 74884 5960 74930 5972
rect 73906 5428 73912 5926
rect 73906 5384 73918 5428
rect 74884 5414 74890 5960
rect 73136 5334 73624 5340
rect 73136 5300 73148 5334
rect 73612 5300 73624 5334
rect 73136 5294 73624 5300
rect 73344 5042 73404 5294
rect 73858 5202 73918 5384
rect 74874 5384 74890 5414
rect 74924 5414 74930 5960
rect 74924 5384 74934 5414
rect 74154 5334 74642 5340
rect 74154 5300 74166 5334
rect 74630 5300 74642 5334
rect 74154 5294 74642 5300
rect 74364 5202 74424 5294
rect 74874 5202 74934 5384
rect 73858 5142 74934 5202
rect 73338 4982 73344 5042
rect 73404 4982 73410 5042
rect 73858 4930 73918 5142
rect 73852 4870 73858 4930
rect 73918 4870 73924 4930
rect 73136 4810 73624 4816
rect 73136 4776 73148 4810
rect 73612 4776 73624 4810
rect 73136 4770 73624 4776
rect 74154 4810 74642 4816
rect 74154 4776 74166 4810
rect 74630 4776 74642 4810
rect 74154 4770 74642 4776
rect 72842 4684 72854 4726
rect 71870 4190 71876 4668
rect 72848 4204 72854 4684
rect 71870 4150 71880 4190
rect 71100 4100 71588 4106
rect 71100 4066 71112 4100
rect 71576 4066 71588 4100
rect 71100 4060 71588 4066
rect 70796 3758 70802 3818
rect 70862 3758 70868 3818
rect 71328 3584 71388 4060
rect 71820 3692 71880 4150
rect 72842 4150 72854 4204
rect 72888 4684 72902 4726
rect 73866 4726 73912 4738
rect 72888 4204 72894 4684
rect 72888 4150 72902 4204
rect 73866 4196 73872 4726
rect 72118 4100 72606 4106
rect 72118 4066 72130 4100
rect 72594 4066 72606 4100
rect 72118 4060 72606 4066
rect 72346 3694 72406 4060
rect 72842 3818 72902 4150
rect 73856 4150 73872 4196
rect 73906 4196 73912 4726
rect 74884 4726 74930 4738
rect 73906 4150 73916 4196
rect 74884 4178 74890 4726
rect 73136 4100 73624 4106
rect 73136 4066 73148 4100
rect 73612 4066 73624 4100
rect 73136 4060 73624 4066
rect 73360 3822 73420 4060
rect 73856 4024 73916 4150
rect 74876 4150 74890 4178
rect 74924 4178 74930 4726
rect 74924 4150 74936 4178
rect 74154 4100 74642 4106
rect 74154 4066 74166 4100
rect 74630 4066 74642 4100
rect 74154 4060 74642 4066
rect 74362 4026 74422 4060
rect 74876 4026 74936 4150
rect 74362 4024 74936 4026
rect 73856 3964 74936 4024
rect 73856 3928 73916 3964
rect 73850 3868 73856 3928
rect 73916 3868 73922 3928
rect 72836 3758 72842 3818
rect 72902 3758 72908 3818
rect 73354 3762 73360 3822
rect 73420 3762 73426 3822
rect 74866 3762 74872 3822
rect 74932 3762 74938 3822
rect 71814 3632 71820 3692
rect 71880 3632 71886 3692
rect 70082 3578 70570 3584
rect 70082 3544 70094 3578
rect 70558 3544 70570 3578
rect 70082 3538 70570 3544
rect 71100 3578 71588 3584
rect 71100 3544 71112 3578
rect 71576 3544 71588 3578
rect 71100 3538 71588 3544
rect 69790 3448 69800 3494
rect 68816 2958 68822 3446
rect 69794 2978 69800 3448
rect 68816 2918 68826 2958
rect 68046 2868 68534 2874
rect 68046 2834 68058 2868
rect 68522 2834 68534 2868
rect 68046 2828 68534 2834
rect 63668 2716 63674 2776
rect 63734 2716 63740 2776
rect 65710 2716 65716 2776
rect 65776 2716 65782 2776
rect 67746 2716 67752 2776
rect 67812 2716 67818 2776
rect 68258 2666 68318 2828
rect 68766 2768 68826 2918
rect 69788 2918 69800 2978
rect 69834 3448 69850 3494
rect 70812 3494 70858 3506
rect 69834 2978 69840 3448
rect 69834 2918 69848 2978
rect 70812 2962 70818 3494
rect 69064 2868 69552 2874
rect 69064 2834 69076 2868
rect 69540 2834 69552 2868
rect 69064 2828 69552 2834
rect 68766 2708 68972 2768
rect 62506 2444 62566 2656
rect 63164 2602 63170 2662
rect 63230 2602 63236 2662
rect 68252 2606 68258 2666
rect 68318 2606 68324 2666
rect 62656 2488 62662 2548
rect 62722 2488 62728 2548
rect 64686 2488 64692 2548
rect 64752 2488 64758 2548
rect 66724 2488 66730 2548
rect 66790 2488 66796 2548
rect 68760 2488 68766 2548
rect 68826 2488 68832 2548
rect 62500 2384 62506 2444
rect 62566 2384 62572 2444
rect 60920 2344 61408 2350
rect 60920 2310 60932 2344
rect 61396 2310 61408 2344
rect 60920 2304 61408 2310
rect 61938 2344 62426 2350
rect 61938 2310 61950 2344
rect 62414 2310 62426 2344
rect 61938 2304 62426 2310
rect 60624 1778 60638 2260
rect 60632 1704 60638 1778
rect 59654 1684 59664 1698
rect 58884 1634 59372 1640
rect 58884 1600 58896 1634
rect 59360 1600 59372 1634
rect 58884 1594 59372 1600
rect 59104 1336 59164 1594
rect 59604 1442 59664 1684
rect 60628 1684 60638 1704
rect 60672 1778 60684 2260
rect 61650 2260 61696 2272
rect 60672 1704 60678 1778
rect 61650 1710 61656 2260
rect 60672 1684 60688 1704
rect 59902 1634 60390 1640
rect 59902 1600 59914 1634
rect 60378 1600 60390 1634
rect 59902 1594 60390 1600
rect 59598 1382 59604 1442
rect 59664 1382 59670 1442
rect 60118 1336 60178 1594
rect 59098 1276 59104 1336
rect 59164 1276 59170 1336
rect 60112 1276 60118 1336
rect 60178 1276 60184 1336
rect 58584 1166 58590 1226
rect 58650 1166 58656 1226
rect 57866 1112 58354 1118
rect 57866 1078 57878 1112
rect 58342 1078 58354 1112
rect 57866 1072 58354 1078
rect 57574 1014 57584 1028
rect 55830 402 56318 408
rect 55830 368 55842 402
rect 56306 368 56318 402
rect 55830 362 56318 368
rect 54392 244 54398 304
rect 54458 244 54464 304
rect 55528 244 55534 304
rect 55594 244 55600 304
rect 56046 196 56106 362
rect 56040 136 56046 196
rect 56106 136 56112 196
rect 56554 -60 56614 452
rect 57578 452 57584 1014
rect 57618 1014 57634 1028
rect 58590 1028 58650 1166
rect 59104 1118 59164 1276
rect 60118 1118 60178 1276
rect 60628 1226 60688 1684
rect 61644 1684 61656 1710
rect 61690 1710 61696 2260
rect 62662 2260 62722 2488
rect 62956 2344 63444 2350
rect 62956 2310 62968 2344
rect 63432 2310 63444 2344
rect 62956 2304 63444 2310
rect 63974 2344 64462 2350
rect 63974 2310 63986 2344
rect 64450 2310 64462 2344
rect 63974 2304 64462 2310
rect 63686 2260 63732 2272
rect 64692 2260 64752 2488
rect 64992 2344 65480 2350
rect 64992 2310 65004 2344
rect 65468 2310 65480 2344
rect 64992 2304 65480 2310
rect 66010 2344 66498 2350
rect 66010 2310 66022 2344
rect 66486 2310 66498 2344
rect 66010 2304 66498 2310
rect 65722 2260 65768 2272
rect 66730 2260 66790 2488
rect 67028 2344 67516 2350
rect 67028 2310 67040 2344
rect 67504 2310 67516 2344
rect 67028 2304 67516 2310
rect 68046 2344 68534 2350
rect 68046 2310 68058 2344
rect 68522 2310 68534 2344
rect 68046 2304 68534 2310
rect 62662 2204 62674 2260
rect 61690 1684 61704 1710
rect 62668 1708 62674 2204
rect 60920 1634 61408 1640
rect 60920 1600 60932 1634
rect 61396 1600 61408 1634
rect 60920 1594 61408 1600
rect 61150 1336 61210 1594
rect 61644 1442 61704 1684
rect 62666 1684 62674 1708
rect 62708 2204 62722 2260
rect 63680 2224 63692 2260
rect 62708 1708 62714 2204
rect 63686 1736 63692 2224
rect 62708 1684 62726 1708
rect 61938 1634 62426 1640
rect 61938 1600 61950 1634
rect 62414 1600 62426 1634
rect 61938 1594 62426 1600
rect 61792 1488 61798 1548
rect 61858 1488 61864 1548
rect 61638 1382 61644 1442
rect 61704 1382 61710 1442
rect 61144 1276 61150 1336
rect 61210 1276 61216 1336
rect 61798 1304 61858 1488
rect 62162 1336 62222 1594
rect 60622 1166 60628 1226
rect 60688 1166 60694 1226
rect 58884 1112 59372 1118
rect 58884 1078 58896 1112
rect 59360 1078 59372 1112
rect 58884 1072 59372 1078
rect 59902 1112 60390 1118
rect 59902 1078 59914 1112
rect 60378 1078 60390 1112
rect 59902 1072 60390 1078
rect 57618 452 57624 1014
rect 57578 440 57624 452
rect 58590 452 58602 1028
rect 58636 452 58650 1028
rect 59614 1028 59660 1040
rect 59614 494 59620 1028
rect 56848 402 57336 408
rect 56848 368 56860 402
rect 57324 368 57336 402
rect 56848 362 57336 368
rect 57866 402 58354 408
rect 57866 368 57878 402
rect 58342 368 58354 402
rect 57866 362 58354 368
rect 57060 196 57120 362
rect 57060 130 57120 136
rect 58082 196 58142 362
rect 58082 130 58142 136
rect 58590 -60 58650 452
rect 59604 452 59620 494
rect 59654 494 59660 1028
rect 60628 1028 60688 1166
rect 61150 1118 61210 1276
rect 61642 1244 61858 1304
rect 62156 1276 62162 1336
rect 62222 1276 62228 1336
rect 60920 1112 61408 1118
rect 60920 1078 60932 1112
rect 61396 1078 61408 1112
rect 60920 1072 61408 1078
rect 59654 452 59664 494
rect 58884 402 59372 408
rect 58884 368 58896 402
rect 59360 368 59372 402
rect 58884 362 59372 368
rect 59094 202 59154 362
rect 59604 304 59664 452
rect 60628 452 60638 1028
rect 60672 452 60688 1028
rect 61642 1028 61702 1244
rect 62162 1118 62222 1276
rect 62666 1226 62726 1684
rect 63676 1684 63692 1736
rect 63726 2224 63740 2260
rect 63726 1736 63732 2224
rect 64692 2210 64710 2260
rect 63726 1684 63736 1736
rect 64704 1714 64710 2210
rect 62956 1634 63444 1640
rect 62956 1600 62968 1634
rect 63432 1600 63444 1634
rect 62956 1594 63444 1600
rect 63170 1336 63230 1594
rect 63676 1548 63736 1684
rect 64702 1684 64710 1714
rect 64744 2210 64752 2260
rect 65716 2228 65728 2260
rect 64744 1714 64750 2210
rect 65722 1724 65728 2228
rect 64744 1684 64762 1714
rect 63974 1634 64462 1640
rect 63974 1600 63986 1634
rect 64450 1600 64462 1634
rect 63974 1594 64462 1600
rect 63670 1488 63676 1548
rect 63736 1488 63742 1548
rect 63674 1382 63680 1442
rect 63740 1382 63746 1442
rect 63164 1276 63170 1336
rect 63230 1276 63236 1336
rect 62660 1166 62666 1226
rect 62726 1166 62732 1226
rect 61938 1112 62426 1118
rect 61938 1078 61950 1112
rect 62414 1078 62426 1112
rect 61938 1072 62426 1078
rect 61642 1002 61656 1028
rect 59902 402 60390 408
rect 59902 368 59914 402
rect 60378 368 60390 402
rect 59902 362 60390 368
rect 59598 244 59604 304
rect 59664 244 59670 304
rect 60120 202 60180 362
rect 59094 196 59156 202
rect 59094 190 59096 196
rect 60120 196 60182 202
rect 60120 190 60122 196
rect 59096 130 59156 136
rect 60122 130 60182 136
rect 60628 -60 60688 452
rect 61650 452 61656 1002
rect 61690 1002 61702 1028
rect 62666 1028 62726 1166
rect 63170 1118 63230 1276
rect 62956 1112 63444 1118
rect 62956 1078 62968 1112
rect 63432 1078 63444 1112
rect 62956 1072 63444 1078
rect 61690 452 61696 1002
rect 61650 440 61696 452
rect 62666 452 62674 1028
rect 62708 452 62726 1028
rect 63680 1028 63740 1382
rect 64188 1336 64248 1594
rect 64182 1276 64188 1336
rect 64248 1276 64254 1336
rect 64188 1118 64248 1276
rect 64702 1226 64762 1684
rect 65714 1684 65728 1724
rect 65762 2228 65776 2260
rect 65762 1724 65768 2228
rect 66730 2216 66746 2260
rect 65762 1684 65774 1724
rect 66740 1708 66746 2216
rect 64992 1634 65480 1640
rect 64992 1600 65004 1634
rect 65468 1600 65480 1634
rect 64992 1594 65480 1600
rect 65214 1336 65274 1594
rect 65714 1548 65774 1684
rect 66738 1684 66746 1708
rect 66780 2216 66790 2260
rect 67758 2260 67804 2272
rect 66780 1708 66786 2216
rect 67758 1730 67764 2260
rect 66780 1684 66798 1708
rect 66010 1634 66498 1640
rect 66010 1600 66022 1634
rect 66486 1600 66498 1634
rect 66010 1594 66498 1600
rect 65708 1488 65714 1548
rect 65774 1488 65780 1548
rect 65710 1382 65716 1442
rect 65776 1382 65782 1442
rect 65208 1276 65214 1336
rect 65274 1276 65280 1336
rect 64696 1166 64702 1226
rect 64762 1166 64768 1226
rect 63974 1112 64462 1118
rect 63974 1078 63986 1112
rect 64450 1078 64462 1112
rect 63974 1072 64462 1078
rect 63680 1002 63692 1028
rect 60920 402 61408 408
rect 60920 368 60932 402
rect 61396 368 61408 402
rect 60920 362 61408 368
rect 61938 402 62426 408
rect 61938 368 61950 402
rect 62414 368 62426 402
rect 61938 362 62426 368
rect 61134 196 61194 362
rect 61134 130 61194 136
rect 62170 196 62230 362
rect 62170 130 62230 136
rect 62666 -60 62726 452
rect 63686 452 63692 1002
rect 63726 1002 63740 1028
rect 64702 1028 64762 1166
rect 65214 1118 65274 1276
rect 64992 1112 65480 1118
rect 64992 1078 65004 1112
rect 65468 1078 65480 1112
rect 64992 1072 65480 1078
rect 63726 452 63732 1002
rect 63686 440 63732 452
rect 64702 452 64710 1028
rect 64744 452 64762 1028
rect 65716 1028 65776 1382
rect 66216 1336 66276 1594
rect 66210 1276 66216 1336
rect 66276 1276 66282 1336
rect 66216 1118 66276 1276
rect 66738 1226 66798 1684
rect 67750 1684 67764 1730
rect 67798 1730 67804 2260
rect 68766 2260 68826 2488
rect 68912 2444 68972 2708
rect 68906 2384 68912 2444
rect 68972 2384 68978 2444
rect 69276 2350 69336 2828
rect 69788 2548 69848 2918
rect 70806 2918 70818 2962
rect 70852 2962 70858 3494
rect 71820 3494 71880 3632
rect 72346 3584 72406 3634
rect 73360 3584 73420 3762
rect 73854 3634 73860 3694
rect 73920 3634 73926 3694
rect 72118 3578 72606 3584
rect 72118 3544 72130 3578
rect 72594 3544 72606 3578
rect 72118 3538 72606 3544
rect 73136 3578 73624 3584
rect 73136 3544 73148 3578
rect 73612 3544 73624 3578
rect 73136 3538 73624 3544
rect 71820 3448 71836 3494
rect 71830 2966 71836 3448
rect 70852 2918 70866 2962
rect 70082 2868 70570 2874
rect 70082 2834 70094 2868
rect 70558 2834 70570 2868
rect 70082 2828 70570 2834
rect 69782 2488 69788 2548
rect 69848 2488 69854 2548
rect 70296 2350 70356 2828
rect 70806 2776 70866 2918
rect 71822 2918 71836 2966
rect 71870 3448 71880 3494
rect 72848 3494 72894 3506
rect 73860 3494 73920 3634
rect 74154 3578 74642 3584
rect 74154 3544 74166 3578
rect 74630 3544 74642 3578
rect 74154 3538 74642 3544
rect 71870 2966 71876 3448
rect 71870 2918 71882 2966
rect 72848 2962 72854 3494
rect 71100 2868 71588 2874
rect 71100 2834 71112 2868
rect 71576 2834 71588 2868
rect 71100 2828 71588 2834
rect 70800 2716 70806 2776
rect 70866 2716 70872 2776
rect 70802 2488 70808 2548
rect 70868 2488 70874 2548
rect 69064 2344 69552 2350
rect 69064 2310 69076 2344
rect 69540 2310 69552 2344
rect 69064 2304 69552 2310
rect 70082 2344 70570 2350
rect 70082 2310 70094 2344
rect 70558 2310 70570 2344
rect 70082 2304 70570 2310
rect 68766 2216 68782 2260
rect 67798 1684 67810 1730
rect 68776 1710 68782 2216
rect 67028 1634 67516 1640
rect 67028 1600 67040 1634
rect 67504 1600 67516 1634
rect 67028 1594 67516 1600
rect 67236 1336 67296 1594
rect 67578 1488 67584 1548
rect 67644 1488 67650 1548
rect 67230 1276 67236 1336
rect 67296 1276 67302 1336
rect 67584 1296 67644 1488
rect 67750 1442 67810 1684
rect 68770 1684 68782 1710
rect 68816 2216 68826 2260
rect 69794 2260 69840 2272
rect 68816 1710 68822 2216
rect 69794 1724 69800 2260
rect 68816 1684 68830 1710
rect 68046 1634 68534 1640
rect 68046 1600 68058 1634
rect 68522 1600 68534 1634
rect 68046 1594 68534 1600
rect 67744 1382 67750 1442
rect 67810 1382 67816 1442
rect 68256 1336 68316 1594
rect 66732 1166 66738 1226
rect 66798 1166 66804 1226
rect 66010 1112 66498 1118
rect 66010 1078 66022 1112
rect 66486 1078 66498 1112
rect 66010 1072 66498 1078
rect 65716 992 65728 1028
rect 62956 402 63444 408
rect 62956 368 62968 402
rect 63432 368 63444 402
rect 62956 362 63444 368
rect 63974 402 64462 408
rect 63974 368 63986 402
rect 64450 368 64462 402
rect 63974 362 64462 368
rect 63176 196 63236 362
rect 64190 196 64250 362
rect 64184 136 64190 196
rect 64250 136 64256 196
rect 63176 130 63236 136
rect 64702 -60 64762 452
rect 65722 452 65728 992
rect 65762 992 65776 1028
rect 66738 1028 66798 1166
rect 67236 1118 67296 1276
rect 67584 1236 67810 1296
rect 68250 1276 68256 1336
rect 68316 1276 68322 1336
rect 67028 1112 67516 1118
rect 67028 1078 67040 1112
rect 67504 1078 67516 1112
rect 67028 1072 67516 1078
rect 65762 452 65768 992
rect 65722 440 65768 452
rect 66738 452 66746 1028
rect 66780 452 66798 1028
rect 67750 1028 67810 1236
rect 68256 1118 68316 1276
rect 68770 1226 68830 1684
rect 69790 1684 69800 1724
rect 69834 1724 69840 2260
rect 70808 2260 70868 2488
rect 71310 2350 71370 2828
rect 71822 2548 71882 2918
rect 72838 2918 72854 2962
rect 72888 2962 72894 3494
rect 73858 3460 73872 3494
rect 73860 3450 73872 3460
rect 72888 2918 72898 2962
rect 72118 2868 72606 2874
rect 72118 2834 72130 2868
rect 72594 2834 72606 2868
rect 72118 2828 72606 2834
rect 71816 2488 71822 2548
rect 71882 2488 71888 2548
rect 71816 2384 71822 2444
rect 71882 2384 71888 2444
rect 71100 2344 71588 2350
rect 71100 2310 71112 2344
rect 71576 2310 71588 2344
rect 71100 2304 71588 2310
rect 71318 2300 71378 2304
rect 70808 2194 70818 2260
rect 70812 1730 70818 2194
rect 69834 1684 69850 1724
rect 69064 1634 69552 1640
rect 69064 1600 69076 1634
rect 69540 1600 69552 1634
rect 69064 1594 69552 1600
rect 69282 1336 69342 1594
rect 69790 1442 69850 1684
rect 70802 1684 70818 1730
rect 70852 2194 70868 2260
rect 71822 2260 71882 2384
rect 72346 2350 72406 2828
rect 72838 2776 72898 2918
rect 73866 2918 73872 3450
rect 73906 3450 73920 3494
rect 74872 3494 74932 3762
rect 73906 2918 73912 3450
rect 74872 3440 74890 3494
rect 73866 2906 73912 2918
rect 74884 2918 74890 3440
rect 74924 3456 74936 3494
rect 74924 3440 74932 3456
rect 74924 2918 74930 3440
rect 74884 2906 74930 2918
rect 73136 2868 73624 2874
rect 73136 2834 73148 2868
rect 73612 2834 73624 2868
rect 73136 2828 73624 2834
rect 74154 2868 74642 2874
rect 74154 2834 74166 2868
rect 74630 2834 74642 2868
rect 74154 2828 74642 2834
rect 72832 2716 72838 2776
rect 72898 2716 72904 2776
rect 73358 2666 73418 2828
rect 74366 2666 74426 2828
rect 74984 2776 75044 8566
rect 75106 7652 75112 7712
rect 75172 7652 75178 7712
rect 75112 6154 75172 7652
rect 75228 7388 75288 8680
rect 75344 7430 75350 7490
rect 75410 7430 75416 7490
rect 75222 7328 75228 7388
rect 75288 7328 75294 7388
rect 75106 6094 75112 6154
rect 75172 6094 75178 6154
rect 75102 5192 75108 5252
rect 75168 5192 75174 5252
rect 75108 3928 75168 5192
rect 75228 4026 75288 7328
rect 75222 3966 75228 4026
rect 75288 3966 75294 4026
rect 75102 3868 75108 3928
rect 75168 3868 75174 3928
rect 74978 2716 74984 2776
rect 75044 2716 75050 2776
rect 73352 2606 73358 2666
rect 73418 2606 73424 2666
rect 74360 2606 74366 2666
rect 74426 2606 74432 2666
rect 75228 2550 75288 3966
rect 75350 3694 75410 7430
rect 75478 6262 75538 8784
rect 75476 6256 75538 6262
rect 75536 6196 75538 6256
rect 75476 6190 75538 6196
rect 75478 3822 75538 6190
rect 75472 3762 75478 3822
rect 75538 3762 75544 3822
rect 75344 3634 75350 3694
rect 75410 3634 75416 3694
rect 75600 2666 75660 13594
rect 75706 9784 75712 9844
rect 75772 9784 75778 9844
rect 75594 2606 75600 2666
rect 75660 2606 75666 2666
rect 72838 2488 72844 2548
rect 72904 2488 72910 2548
rect 73860 2490 75288 2550
rect 72118 2344 72606 2350
rect 72118 2310 72130 2344
rect 72594 2310 72606 2344
rect 72118 2304 72606 2310
rect 71822 2214 71836 2260
rect 70852 1730 70858 2194
rect 70852 1684 70862 1730
rect 70082 1634 70570 1640
rect 70082 1600 70094 1634
rect 70558 1600 70570 1634
rect 70082 1594 70570 1600
rect 69784 1382 69790 1442
rect 69850 1382 69856 1442
rect 70300 1336 70360 1594
rect 69276 1276 69282 1336
rect 69342 1276 69348 1336
rect 70294 1276 70300 1336
rect 70360 1276 70366 1336
rect 68764 1166 68770 1226
rect 68830 1166 68836 1226
rect 68046 1112 68534 1118
rect 68046 1078 68058 1112
rect 68522 1078 68534 1112
rect 68046 1072 68534 1078
rect 67750 992 67764 1028
rect 64992 402 65480 408
rect 64992 368 65004 402
rect 65468 368 65480 402
rect 64992 362 65480 368
rect 66010 402 66498 408
rect 66010 368 66022 402
rect 66486 368 66498 402
rect 66010 362 66498 368
rect 65206 196 65266 362
rect 66216 202 66276 362
rect 65206 130 65266 136
rect 66214 196 66276 202
rect 66274 190 66276 196
rect 66214 130 66274 136
rect 66738 -60 66798 452
rect 67758 452 67764 992
rect 67798 992 67810 1028
rect 68770 1028 68830 1166
rect 69282 1118 69342 1276
rect 70300 1118 70360 1276
rect 70802 1226 70862 1684
rect 71830 1684 71836 2214
rect 71870 2214 71882 2260
rect 72844 2260 72904 2488
rect 73136 2344 73624 2350
rect 73136 2310 73148 2344
rect 73612 2310 73624 2344
rect 73136 2304 73624 2310
rect 71870 1684 71876 2214
rect 72844 2200 72854 2260
rect 72848 1708 72854 2200
rect 71830 1672 71876 1684
rect 72842 1684 72854 1708
rect 72888 2200 72904 2260
rect 73860 2260 73920 2490
rect 74358 2350 74418 2490
rect 74154 2344 74642 2350
rect 74154 2310 74166 2344
rect 74630 2310 74642 2344
rect 74154 2304 74642 2310
rect 72888 1708 72894 2200
rect 72888 1684 72902 1708
rect 71100 1634 71588 1640
rect 71100 1600 71112 1634
rect 71576 1600 71588 1634
rect 71100 1594 71588 1600
rect 72118 1634 72606 1640
rect 72118 1600 72130 1634
rect 72594 1600 72606 1634
rect 72118 1594 72606 1600
rect 71314 1336 71374 1594
rect 71814 1382 71820 1442
rect 71880 1382 71886 1442
rect 71308 1276 71314 1336
rect 71374 1276 71380 1336
rect 70796 1166 70802 1226
rect 70862 1166 70868 1226
rect 69064 1112 69552 1118
rect 69064 1078 69076 1112
rect 69540 1078 69552 1112
rect 69064 1072 69552 1078
rect 70082 1112 70570 1118
rect 70082 1078 70094 1112
rect 70558 1078 70570 1112
rect 70082 1072 70570 1078
rect 67798 452 67804 992
rect 67758 440 67804 452
rect 68770 452 68782 1028
rect 68816 452 68830 1028
rect 69794 1028 69840 1040
rect 69794 504 69800 1028
rect 68254 408 68314 410
rect 67028 402 67516 408
rect 67028 368 67040 402
rect 67504 368 67516 402
rect 67028 362 67516 368
rect 68046 402 68534 408
rect 68046 368 68058 402
rect 68522 368 68534 402
rect 68046 362 68534 368
rect 67232 202 67292 362
rect 67230 196 67292 202
rect 67290 190 67292 196
rect 68254 196 68314 362
rect 67230 130 67290 136
rect 68254 130 68314 136
rect 68770 -60 68830 452
rect 69784 452 69800 504
rect 69834 504 69840 1028
rect 70802 1028 70862 1166
rect 71314 1118 71374 1276
rect 71100 1112 71588 1118
rect 71100 1078 71112 1112
rect 71576 1078 71588 1112
rect 71100 1072 71588 1078
rect 69834 452 69844 504
rect 69064 402 69552 408
rect 69064 368 69076 402
rect 69540 368 69552 402
rect 69064 362 69552 368
rect 69276 196 69336 362
rect 69784 304 69844 452
rect 70802 452 70818 1028
rect 70852 452 70862 1028
rect 71820 1028 71880 1382
rect 72328 1336 72388 1594
rect 72322 1276 72328 1336
rect 72388 1276 72394 1336
rect 72328 1118 72388 1276
rect 72842 1226 72902 1684
rect 73860 1684 73872 2260
rect 73906 1684 73920 2260
rect 74874 2260 74934 2490
rect 74998 2384 75004 2444
rect 75064 2384 75070 2444
rect 74874 2206 74890 2260
rect 73136 1634 73624 1640
rect 73136 1600 73148 1634
rect 73612 1600 73624 1634
rect 73136 1594 73624 1600
rect 73350 1336 73410 1594
rect 73860 1548 73920 1684
rect 74884 1684 74890 2206
rect 74924 2206 74934 2260
rect 74924 1684 74930 2206
rect 74884 1672 74930 1684
rect 74154 1634 74642 1640
rect 74154 1600 74166 1634
rect 74630 1600 74642 1634
rect 74154 1594 74642 1600
rect 73854 1488 73860 1548
rect 73920 1488 73926 1548
rect 73854 1382 73860 1442
rect 73920 1382 73926 1442
rect 73344 1276 73350 1336
rect 73410 1276 73416 1336
rect 72836 1166 72842 1226
rect 72902 1166 72908 1226
rect 72118 1112 72606 1118
rect 72118 1078 72130 1112
rect 72594 1078 72606 1112
rect 72118 1072 72606 1078
rect 71820 984 71836 1028
rect 70082 402 70570 408
rect 70082 368 70094 402
rect 70558 368 70570 402
rect 70082 362 70570 368
rect 69778 244 69784 304
rect 69844 244 69850 304
rect 70296 202 70356 362
rect 70296 196 70358 202
rect 70296 190 70298 196
rect 69276 130 69336 136
rect 70298 130 70358 136
rect 70802 -60 70862 452
rect 71830 452 71836 984
rect 71870 984 71880 1028
rect 72842 1028 72902 1166
rect 73350 1118 73410 1276
rect 73860 1226 73920 1382
rect 73860 1166 74938 1226
rect 73136 1112 73624 1118
rect 73136 1078 73148 1112
rect 73612 1078 73624 1112
rect 73136 1072 73624 1078
rect 71870 452 71876 984
rect 71830 440 71876 452
rect 72842 452 72854 1028
rect 72888 452 72902 1028
rect 73860 1028 73920 1166
rect 74376 1118 74436 1166
rect 74154 1112 74642 1118
rect 74154 1078 74166 1112
rect 74630 1078 74642 1112
rect 74154 1072 74642 1078
rect 73860 1020 73872 1028
rect 71318 408 71378 410
rect 71100 402 71588 408
rect 71100 368 71112 402
rect 71576 368 71588 402
rect 71100 362 71588 368
rect 72118 402 72606 408
rect 72118 368 72130 402
rect 72594 368 72606 402
rect 72118 362 72606 368
rect 71318 202 71378 362
rect 72332 202 72392 362
rect 71316 196 71378 202
rect 71376 190 71378 196
rect 72330 196 72392 202
rect 71316 130 71376 136
rect 72390 190 72392 196
rect 72330 130 72390 136
rect 72842 -60 72902 452
rect 73866 452 73872 1020
rect 73906 1020 73920 1028
rect 74878 1028 74938 1166
rect 73906 452 73912 1020
rect 74878 1010 74890 1028
rect 73866 440 73912 452
rect 74884 452 74890 1010
rect 74924 1010 74938 1028
rect 74924 452 74930 1010
rect 74884 440 74930 452
rect 73352 408 73412 410
rect 73136 402 73624 408
rect 73136 368 73148 402
rect 73612 368 73624 402
rect 73136 362 73624 368
rect 74154 402 74642 408
rect 74154 368 74166 402
rect 74630 368 74642 402
rect 74154 362 74642 368
rect 73352 202 73412 362
rect 75004 304 75064 2384
rect 75712 1442 75772 9784
rect 75706 1382 75712 1442
rect 75772 1382 75778 1442
rect 74998 244 75004 304
rect 75064 244 75070 304
rect 73352 196 73414 202
rect 73352 190 73354 196
rect 73354 130 73414 136
rect 76766 40 76772 14300
rect 76872 40 76878 14300
rect 43832 -106 43982 -60
rect 44028 -106 47202 -60
rect 47262 -106 53654 -60
rect 53714 -106 75756 -60
rect 75816 -106 75918 -60
rect 43832 -260 43878 -106
rect 75878 -260 75918 -106
rect 43832 -306 75918 -260
rect 40334 -746 40344 -446
rect 76156 -746 76166 -446
rect 76766 -746 76878 40
rect 39622 -752 76878 -746
rect 39622 -852 39728 -752
rect 76772 -852 76878 -752
rect 39622 -858 76878 -852
<< via1 >>
rect 11434 30286 12034 30586
rect 35066 30286 35666 30586
rect 15011 29990 31796 30204
rect 18936 28228 18996 28288
rect 20018 28228 20078 28288
rect 20976 28228 21036 28288
rect 19462 27982 19522 28042
rect 21498 27982 21558 28042
rect 17280 27050 17340 27110
rect 18444 27050 18504 27110
rect 17150 26846 17210 26906
rect 15142 24662 15202 24722
rect 18444 26846 18504 26906
rect 24040 28228 24100 28288
rect 25058 28228 25118 28288
rect 23536 27984 23596 28044
rect 20480 26946 20540 27006
rect 18930 25696 18990 25756
rect 26082 28228 26142 28288
rect 27094 28228 27154 28288
rect 25566 27984 25626 28044
rect 22516 26946 22576 27006
rect 27608 27986 27668 28046
rect 24554 27050 24614 27110
rect 24550 26846 24610 26906
rect 20986 25912 21046 25972
rect 21496 25912 21556 25972
rect 20478 25810 20542 25874
rect 19968 25696 20028 25756
rect 20980 25696 21040 25756
rect 17280 24376 17340 24436
rect 17636 21968 17696 22028
rect 17510 21358 17570 21418
rect 14626 20404 14686 20464
rect 14734 20292 14794 20352
rect 12964 19370 13024 19430
rect 15648 20404 15708 20464
rect 15518 20292 15578 20352
rect 14124 19260 14184 19320
rect 16158 19370 16218 19430
rect 12838 18282 12898 18342
rect 14640 18336 14700 18396
rect 14746 18236 14806 18296
rect 17310 19260 17370 19320
rect 15650 18336 15710 18396
rect 17502 19132 17562 19192
rect 15532 18236 15592 18296
rect 12352 17226 12412 17286
rect 12492 17050 12552 17110
rect 13286 17050 13346 17110
rect 15638 17052 15698 17112
rect 13392 16876 13452 16936
rect 17752 21358 17812 21418
rect 18438 24522 18502 24586
rect 18262 24376 18322 24436
rect 22354 25810 22418 25874
rect 28618 27986 28678 28046
rect 30152 28228 30212 28288
rect 31164 28228 31224 28288
rect 29640 27986 29700 28046
rect 26588 27050 26648 27110
rect 26586 26846 26646 26906
rect 27088 26846 27148 26906
rect 23530 25912 23590 25972
rect 21990 25704 22050 25764
rect 23014 25704 23074 25764
rect 19460 24774 19520 24834
rect 20476 24660 20540 24724
rect 24042 25704 24102 25764
rect 32182 28228 32242 28288
rect 31676 27986 31736 28046
rect 28622 26946 28682 27006
rect 28108 26846 28168 26906
rect 25568 25910 25628 25970
rect 21496 24774 21556 24834
rect 22018 24774 22078 24834
rect 22516 24774 22576 24834
rect 29134 26846 29194 26906
rect 30656 26946 30716 27006
rect 29640 26842 29700 26902
rect 30154 26842 30214 26902
rect 30658 26842 30718 26902
rect 31164 26842 31224 26902
rect 31684 26842 31744 26902
rect 26588 25812 26648 25872
rect 32696 27050 32756 27110
rect 33946 27050 34006 27110
rect 27604 25910 27664 25970
rect 28104 25910 28164 25970
rect 28618 25910 28678 25970
rect 29142 25910 29202 25970
rect 29640 25910 29700 25970
rect 30142 25910 30202 25970
rect 22990 24770 23050 24830
rect 18378 24270 18438 24330
rect 18940 24270 19000 24330
rect 19982 24270 20042 24330
rect 20982 24270 21042 24330
rect 23530 24832 23590 24834
rect 23498 24774 23590 24832
rect 23990 24774 24050 24834
rect 23498 24772 23558 24774
rect 24548 24518 24612 24582
rect 25034 24776 25094 24836
rect 24144 24270 24204 24330
rect 25566 24774 25626 24834
rect 30656 25908 30716 25968
rect 31164 25908 31224 25968
rect 31674 25908 31734 25968
rect 30146 25696 30206 25756
rect 31158 25696 31218 25756
rect 27078 24776 27138 24836
rect 26584 24376 26648 24440
rect 25154 24270 25214 24330
rect 26096 24270 26156 24330
rect 27604 24830 27664 24832
rect 27572 24772 27664 24830
rect 27572 24770 27632 24772
rect 28100 24766 28160 24826
rect 28588 24828 28648 24830
rect 28588 24770 28682 24828
rect 28622 24768 28682 24770
rect 32696 25812 32756 25872
rect 32160 25696 32220 25756
rect 29100 24766 29160 24826
rect 29640 24770 29700 24830
rect 31674 24770 31734 24830
rect 30656 24660 30720 24724
rect 33942 24522 34006 24586
rect 32690 24376 32750 24436
rect 18492 24068 18552 24128
rect 21670 24068 21730 24128
rect 19636 23132 19696 23192
rect 20140 23024 20200 23084
rect 21670 23132 21730 23192
rect 21162 23024 21222 23084
rect 22180 23024 22240 23084
rect 19632 22100 19692 22160
rect 20138 21966 20198 22026
rect 25738 24068 25798 24128
rect 23712 23132 23772 23192
rect 23204 23024 23264 23084
rect 24218 23024 24278 23084
rect 21152 21962 21212 22022
rect 22184 21970 22244 22030
rect 25738 23132 25798 23192
rect 25236 23024 25296 23084
rect 26246 23024 26306 23084
rect 23712 22100 23772 22160
rect 23182 21970 23242 22030
rect 24226 21970 24286 22030
rect 29814 24068 29874 24128
rect 27780 23132 27840 23192
rect 27268 23024 27328 23084
rect 28282 23024 28342 23084
rect 25230 21966 25290 22026
rect 26246 21966 26306 22026
rect 25030 21758 25090 21818
rect 18262 21440 18322 21500
rect 19428 21440 19488 21500
rect 17994 20394 18054 20454
rect 17752 19236 17812 19296
rect 17748 19022 17808 19082
rect 17636 17980 17696 18040
rect 12232 16726 12292 16786
rect 18130 20296 18190 20356
rect 17994 16722 18054 16782
rect 21464 21440 21524 21500
rect 21972 21436 22036 21500
rect 20446 20492 20506 20552
rect 33010 24068 33070 24128
rect 29816 23132 29876 23192
rect 29314 23024 29374 23084
rect 30324 23024 30384 23084
rect 27780 22100 27840 22160
rect 27250 21966 27310 22026
rect 28282 21970 28342 22030
rect 26766 21758 26826 21818
rect 26046 21558 26110 21622
rect 31852 23132 31912 23192
rect 31346 23024 31406 23084
rect 29298 21966 29358 22026
rect 30326 21966 30386 22026
rect 31848 22100 31908 22160
rect 31346 21966 31406 22026
rect 33804 21968 33864 22028
rect 32664 21742 32724 21802
rect 30110 21558 30174 21622
rect 31134 21558 31198 21622
rect 32146 21558 32210 21622
rect 26048 21436 26112 21500
rect 22482 20492 22542 20552
rect 22824 20494 22884 20554
rect 20446 20296 20506 20356
rect 21466 20298 21526 20358
rect 19432 20186 19492 20246
rect 21466 20186 21526 20246
rect 18414 19022 18474 19082
rect 25538 20494 25598 20554
rect 29610 21440 29670 21500
rect 31644 21440 31704 21500
rect 26556 20298 26616 20358
rect 24522 20184 24582 20244
rect 26556 20184 26616 20244
rect 20448 19132 20508 19192
rect 20448 18928 20508 18988
rect 22484 19132 22544 19192
rect 22482 19030 22542 19090
rect 22482 18928 22542 18988
rect 19430 17980 19490 18040
rect 18262 17772 18322 17832
rect 20444 17670 20504 17730
rect 24518 19236 24578 19296
rect 21466 17980 21526 18040
rect 21466 17872 21526 17932
rect 25538 19236 25598 19296
rect 25538 18930 25598 18990
rect 29612 20184 29672 20244
rect 26556 18930 26616 18990
rect 30626 20492 30686 20552
rect 31646 20184 31706 20244
rect 32662 20492 32722 20552
rect 27574 19236 27634 19296
rect 27572 18930 27632 18990
rect 22484 17988 22544 18048
rect 24286 17988 24346 18048
rect 22478 17670 22538 17730
rect 22682 17658 22742 17718
rect 19426 16722 19486 16782
rect 24520 17982 24580 18042
rect 29608 19132 29668 19192
rect 30476 19250 30536 19310
rect 30624 19140 30684 19200
rect 30476 18930 30536 18990
rect 30628 18932 30688 18992
rect 26556 17982 26616 18042
rect 26554 17872 26614 17932
rect 21462 16722 21522 16782
rect 18130 16592 18190 16652
rect 12490 16464 12550 16524
rect 13286 16464 13346 16524
rect 15638 16462 15698 16522
rect 13166 16346 13226 16406
rect 26044 17658 26104 17718
rect 31644 19030 31704 19090
rect 34240 22100 34300 22160
rect 33946 21740 34006 21800
rect 34088 21440 34148 21500
rect 33928 20298 33988 20358
rect 32664 19140 32724 19200
rect 33804 19140 33864 19200
rect 32662 18932 32722 18992
rect 27060 17658 27120 17718
rect 29610 17984 29670 18044
rect 30120 17658 30180 17718
rect 30632 17670 30692 17730
rect 31646 17984 31706 18044
rect 33928 18932 33988 18992
rect 33804 17872 33864 17932
rect 32666 17670 32726 17730
rect 29614 16722 29674 16782
rect 31650 16722 31710 16782
rect 22484 16452 22544 16512
rect 34240 20184 34300 20244
rect 34088 16452 34148 16512
rect 12720 16228 12780 16288
rect 52434 30286 53034 30586
rect 76066 30286 76666 30586
rect 56011 29990 72796 30204
rect 59936 28228 59996 28288
rect 61018 28228 61078 28288
rect 61976 28228 62036 28288
rect 60462 27982 60522 28042
rect 62498 27982 62558 28042
rect 58280 27050 58340 27110
rect 59444 27050 59504 27110
rect 58150 26846 58210 26906
rect 56142 24662 56202 24722
rect 59444 26846 59504 26906
rect 65040 28228 65100 28288
rect 66058 28228 66118 28288
rect 64536 27984 64596 28044
rect 61480 26946 61540 27006
rect 59930 25696 59990 25756
rect 67082 28228 67142 28288
rect 68094 28228 68154 28288
rect 66566 27984 66626 28044
rect 63516 26946 63576 27006
rect 68608 27986 68668 28046
rect 65554 27050 65614 27110
rect 65550 26846 65610 26906
rect 61986 25912 62046 25972
rect 62496 25912 62556 25972
rect 61478 25810 61542 25874
rect 60968 25696 61028 25756
rect 61980 25696 62040 25756
rect 58280 24376 58340 24436
rect 58636 21968 58696 22028
rect 58510 21358 58570 21418
rect 55626 20404 55686 20464
rect 55734 20292 55794 20352
rect 53964 19370 54024 19430
rect 56648 20404 56708 20464
rect 56518 20292 56578 20352
rect 55124 19260 55184 19320
rect 57158 19370 57218 19430
rect 53838 18282 53898 18342
rect 55640 18336 55700 18396
rect 55746 18236 55806 18296
rect 58310 19260 58370 19320
rect 56650 18336 56710 18396
rect 58502 19132 58562 19192
rect 56532 18236 56592 18296
rect 53352 17226 53412 17286
rect 53492 17050 53552 17110
rect 54392 16876 54452 16936
rect 58752 21358 58812 21418
rect 59438 24522 59502 24586
rect 59262 24376 59322 24436
rect 63354 25810 63418 25874
rect 69618 27986 69678 28046
rect 71152 28228 71212 28288
rect 72164 28228 72224 28288
rect 70640 27986 70700 28046
rect 67588 27050 67648 27110
rect 67586 26846 67646 26906
rect 68088 26846 68148 26906
rect 64530 25912 64590 25972
rect 62990 25704 63050 25764
rect 64014 25704 64074 25764
rect 60460 24774 60520 24834
rect 61476 24660 61540 24724
rect 65042 25704 65102 25764
rect 73182 28228 73242 28288
rect 72676 27986 72736 28046
rect 69622 26946 69682 27006
rect 69108 26846 69168 26906
rect 66568 25910 66628 25970
rect 62496 24774 62556 24834
rect 63018 24774 63078 24834
rect 63516 24774 63576 24834
rect 70134 26846 70194 26906
rect 71656 26946 71716 27006
rect 70640 26842 70700 26902
rect 71154 26842 71214 26902
rect 71658 26842 71718 26902
rect 72164 26842 72224 26902
rect 72684 26842 72744 26902
rect 67588 25812 67648 25872
rect 73696 27050 73756 27110
rect 74946 27050 75006 27110
rect 68604 25910 68664 25970
rect 69104 25910 69164 25970
rect 69618 25910 69678 25970
rect 70142 25910 70202 25970
rect 70640 25910 70700 25970
rect 71142 25910 71202 25970
rect 63990 24770 64050 24830
rect 59378 24270 59438 24330
rect 59940 24270 60000 24330
rect 60982 24270 61042 24330
rect 61982 24270 62042 24330
rect 64530 24832 64590 24834
rect 64498 24774 64590 24832
rect 64990 24774 65050 24834
rect 64498 24772 64558 24774
rect 65548 24518 65612 24582
rect 66034 24776 66094 24836
rect 65144 24270 65204 24330
rect 66566 24774 66626 24834
rect 71656 25908 71716 25968
rect 72164 25908 72224 25968
rect 72674 25908 72734 25968
rect 71146 25696 71206 25756
rect 72158 25696 72218 25756
rect 68078 24776 68138 24836
rect 67584 24376 67648 24440
rect 66154 24270 66214 24330
rect 67096 24270 67156 24330
rect 68604 24830 68664 24832
rect 68572 24772 68664 24830
rect 68572 24770 68632 24772
rect 69100 24766 69160 24826
rect 69588 24828 69648 24830
rect 69588 24770 69682 24828
rect 69622 24768 69682 24770
rect 73696 25812 73756 25872
rect 73160 25696 73220 25756
rect 70100 24766 70160 24826
rect 70640 24770 70700 24830
rect 72674 24770 72734 24830
rect 71656 24660 71720 24724
rect 74942 24522 75006 24586
rect 73690 24376 73750 24436
rect 59492 24068 59552 24128
rect 62670 24068 62730 24128
rect 60636 23132 60696 23192
rect 61140 23024 61200 23084
rect 62670 23132 62730 23192
rect 62162 23024 62222 23084
rect 63180 23024 63240 23084
rect 60632 22100 60692 22160
rect 61138 21966 61198 22026
rect 66738 24068 66798 24128
rect 64712 23132 64772 23192
rect 64204 23024 64264 23084
rect 65218 23024 65278 23084
rect 62152 21962 62212 22022
rect 63184 21970 63244 22030
rect 66738 23132 66798 23192
rect 66236 23024 66296 23084
rect 67246 23024 67306 23084
rect 64712 22100 64772 22160
rect 64182 21970 64242 22030
rect 65226 21970 65286 22030
rect 70814 24068 70874 24128
rect 68780 23132 68840 23192
rect 68268 23024 68328 23084
rect 69282 23024 69342 23084
rect 66230 21966 66290 22026
rect 67246 21966 67306 22026
rect 66030 21758 66090 21818
rect 59262 21440 59322 21500
rect 60428 21440 60488 21500
rect 58994 20394 59054 20454
rect 58752 19236 58812 19296
rect 58748 19022 58808 19082
rect 58636 17980 58696 18040
rect 53232 16726 53292 16786
rect -2680 15700 8084 15992
rect 59130 20296 59190 20356
rect 58994 16722 59054 16782
rect 62464 21440 62524 21500
rect 62972 21436 63036 21500
rect 61446 20492 61506 20552
rect 74010 24068 74070 24128
rect 70816 23132 70876 23192
rect 70314 23024 70374 23084
rect 71324 23024 71384 23084
rect 68780 22100 68840 22160
rect 68250 21966 68310 22026
rect 69282 21970 69342 22030
rect 67766 21758 67826 21818
rect 67046 21558 67110 21622
rect 72852 23132 72912 23192
rect 72346 23024 72406 23084
rect 70298 21966 70358 22026
rect 71326 21966 71386 22026
rect 72848 22100 72908 22160
rect 72346 21966 72406 22026
rect 74804 21968 74864 22028
rect 73664 21742 73724 21802
rect 71110 21558 71174 21622
rect 72134 21558 72198 21622
rect 73146 21558 73210 21622
rect 67048 21436 67112 21500
rect 63482 20492 63542 20552
rect 63824 20494 63884 20554
rect 61446 20296 61506 20356
rect 62466 20298 62526 20358
rect 60432 20186 60492 20246
rect 62466 20186 62526 20246
rect 59414 19022 59474 19082
rect 66538 20494 66598 20554
rect 70610 21440 70670 21500
rect 72644 21440 72704 21500
rect 67556 20298 67616 20358
rect 65522 20184 65582 20244
rect 67556 20184 67616 20244
rect 61448 19132 61508 19192
rect 61448 18928 61508 18988
rect 63484 19132 63544 19192
rect 63482 19030 63542 19090
rect 63482 18928 63542 18988
rect 60430 17980 60490 18040
rect 59262 17772 59322 17832
rect 61444 17670 61504 17730
rect 65518 19236 65578 19296
rect 62466 17980 62526 18040
rect 62466 17872 62526 17932
rect 66538 19236 66598 19296
rect 66538 18930 66598 18990
rect 70612 20184 70672 20244
rect 67556 18930 67616 18990
rect 71626 20492 71686 20552
rect 72646 20184 72706 20244
rect 73662 20492 73722 20552
rect 68574 19236 68634 19296
rect 68572 18930 68632 18990
rect 63484 17988 63544 18048
rect 65286 17988 65346 18048
rect 63478 17670 63538 17730
rect 63682 17658 63742 17718
rect 60426 16722 60486 16782
rect 65520 17982 65580 18042
rect 70608 19132 70668 19192
rect 71476 19250 71536 19310
rect 71624 19140 71684 19200
rect 71476 18930 71536 18990
rect 71628 18932 71688 18992
rect 67556 17982 67616 18042
rect 67554 17872 67614 17932
rect 62462 16722 62522 16782
rect 59130 16592 59190 16652
rect 54286 16464 54346 16524
rect 54166 16346 54226 16406
rect 67044 17658 67104 17718
rect 72644 19030 72704 19090
rect 75240 22100 75300 22160
rect 74946 21740 75006 21800
rect 75088 21440 75148 21500
rect 74928 20298 74988 20358
rect 73664 19140 73724 19200
rect 74804 19140 74864 19200
rect 73662 18932 73722 18992
rect 68060 17658 68120 17718
rect 70610 17984 70670 18044
rect 71120 17658 71180 17718
rect 71632 17670 71692 17730
rect 72646 17984 72706 18044
rect 74928 18932 74988 18992
rect 74804 17872 74864 17932
rect 73666 17670 73726 17730
rect 70614 16722 70674 16782
rect 72650 16722 72710 16782
rect 63484 16452 63544 16512
rect 75240 20184 75300 20244
rect 75088 16452 75148 16512
rect 53720 16228 53780 16288
rect 38320 15700 49084 15992
rect 12838 14952 12898 15012
rect 13166 14962 13226 15022
rect 12232 14816 12292 14876
rect 12352 14818 12412 14878
rect 12492 14836 12552 14896
rect 12720 14852 12780 14912
rect 12100 14688 12160 14748
rect -2276 13782 -1748 14300
rect -3342 1924 -2908 13306
rect 9388 14090 9448 14150
rect 10914 13956 10974 14016
rect 12100 7488 12160 7548
rect 7552 6562 7612 6622
rect 1442 6416 1502 6476
rect 5522 6416 5582 6476
rect 288 6288 348 6348
rect 2966 6288 3026 6348
rect 3998 6288 4058 6348
rect 1946 5326 2006 5386
rect 1446 5222 1506 5282
rect 2970 5326 3030 5386
rect 2464 5118 2524 5178
rect 288 4056 348 4116
rect 7058 6288 7118 6348
rect 4002 5326 4062 5386
rect 3482 5222 3542 5282
rect 9582 6416 9642 6476
rect 11766 6416 11826 6476
rect 8054 6288 8114 6348
rect 5002 5326 5062 5386
rect 6022 5326 6082 5386
rect 5518 5222 5578 5282
rect 4500 5118 4560 5178
rect 1938 4056 1998 4116
rect 3476 4176 3536 4236
rect 7042 5326 7102 5386
rect 6532 5118 6592 5178
rect 5008 4056 5068 4116
rect 8052 5326 8112 5386
rect 7552 5222 7612 5282
rect 9066 5326 9126 5386
rect 10084 5326 10144 5386
rect 9588 5222 9648 5282
rect 8566 5118 8626 5178
rect 6016 4056 6076 4116
rect 2464 3112 2524 3172
rect 1450 3004 1510 3064
rect 1944 2892 2004 2952
rect 3486 3004 3546 3064
rect 2968 2892 3028 2952
rect 7552 4176 7612 4236
rect 4500 3112 4560 3172
rect 4000 2892 4060 2952
rect 10610 5118 10670 5178
rect 9078 4056 9138 4116
rect 11886 5326 11946 5386
rect 11888 4670 11948 4730
rect 11766 4176 11826 4236
rect 10104 4056 10164 4116
rect 6532 3112 6592 3172
rect 5522 3004 5582 3064
rect 5000 2892 5060 2952
rect 6020 2892 6080 2952
rect 7556 3004 7616 3064
rect 7040 2892 7100 2952
rect 288 1930 348 1990
rect 2958 1930 3018 1990
rect 3990 1930 4050 1990
rect 8050 2892 8110 2952
rect 8566 3112 8626 3172
rect 10610 3112 10670 3172
rect 9592 3004 9652 3064
rect 9064 2892 9124 2952
rect 10082 2892 10142 2952
rect 7050 1930 7110 1990
rect 8046 1930 8106 1990
rect 11886 2892 11946 2952
rect 1444 1800 1504 1860
rect 5524 1800 5584 1860
rect 9584 1800 9644 1860
rect 11766 1800 11826 1860
rect 2922 434 2982 494
rect -1046 274 -986 292
rect -1046 240 -1030 274
rect -1030 240 -996 274
rect -996 240 -986 274
rect -1046 232 -986 240
rect -998 106 -986 166
rect -986 106 -952 166
rect -952 106 -938 166
rect -1046 34 -986 42
rect -1046 0 -1030 34
rect -1030 0 -996 34
rect -996 0 -986 34
rect -1046 -18 -986 0
rect 4960 434 5020 494
rect 6996 434 7056 494
rect 3940 322 4000 382
rect 9032 434 9092 494
rect 8014 322 8074 382
rect 12232 6416 12292 6476
rect 12610 14698 12670 14758
rect 12492 12006 12552 12066
rect 12492 9914 12552 9974
rect 12492 8672 12552 8732
rect 12720 13956 12780 14016
rect 13286 14954 13346 15014
rect 13166 14090 13226 14150
rect 12962 12732 13022 12792
rect 12836 11030 12896 11090
rect 12610 8570 12670 8630
rect 12492 7436 12552 7496
rect 12492 6910 12552 6970
rect 12352 6288 12412 6348
rect 12492 5326 12552 5386
rect 13174 12396 13234 12456
rect 13070 11136 13130 11196
rect 12962 10036 13022 10096
rect 13392 14818 13452 14878
rect 24204 14468 24264 14528
rect 29308 14468 29368 14528
rect 33368 14462 33428 14522
rect 14536 12732 14596 12792
rect 15550 12516 15610 12576
rect 17590 12516 17650 12576
rect 19630 12516 19690 12576
rect 21660 12516 21720 12576
rect 23700 12516 23760 12576
rect 25732 12516 25792 12576
rect 27772 12516 27832 12576
rect 29808 12516 29868 12576
rect 31842 12516 31902 12576
rect 13518 12396 13578 12456
rect 15042 12390 15102 12450
rect 13392 12274 13452 12334
rect 13286 12006 13346 12066
rect 16056 12390 16116 12450
rect 17078 12390 17138 12450
rect 18092 12390 18152 12450
rect 19118 12390 19178 12450
rect 18606 12274 18666 12334
rect 20130 12390 20190 12450
rect 21166 12390 21226 12450
rect 22172 12390 22232 12450
rect 23186 12390 23246 12450
rect 15554 11352 15614 11412
rect 15046 11242 15106 11302
rect 14536 11136 14596 11196
rect 13522 11030 13582 11090
rect 14020 11030 14080 11090
rect 14532 11030 14592 11090
rect 16068 11242 16128 11302
rect 17594 11352 17654 11412
rect 17082 11242 17142 11302
rect 16576 11136 16636 11196
rect 19626 11352 19686 11412
rect 18096 11242 18156 11302
rect 19114 11242 19174 11302
rect 18606 11136 18666 11196
rect 13392 10140 13452 10200
rect 13516 10036 13576 10096
rect 15036 10036 15096 10096
rect 15548 10036 15608 10096
rect 13286 9914 13346 9974
rect 13174 9800 13234 9860
rect 14022 9800 14082 9860
rect 15554 9802 15614 9862
rect 20140 11242 20200 11302
rect 24202 12390 24262 12450
rect 25210 12390 25270 12450
rect 26226 12390 26286 12450
rect 27250 12390 27310 12450
rect 28272 12390 28332 12450
rect 29294 12390 29354 12450
rect 28794 12274 28854 12334
rect 21658 11352 21718 11412
rect 20646 11136 20706 11196
rect 21160 11242 21220 11302
rect 20812 11030 20872 11090
rect 16570 10140 16630 10200
rect 16572 10036 16632 10096
rect 22180 11242 22240 11302
rect 23694 11352 23754 11412
rect 23182 11242 23242 11302
rect 22680 11136 22740 11196
rect 22680 11030 22740 11090
rect 24208 11242 24268 11302
rect 30312 12390 30372 12450
rect 31326 12390 31386 12450
rect 32350 12390 32410 12450
rect 32866 12274 32926 12334
rect 33998 12274 34058 12334
rect 25730 11352 25790 11412
rect 25226 11242 25286 11302
rect 24716 11136 24776 11196
rect 24718 11030 24778 11090
rect 26234 11242 26294 11302
rect 27768 11352 27828 11412
rect 27246 11242 27306 11302
rect 26752 11136 26812 11196
rect 26598 11030 26658 11090
rect 17584 10036 17644 10096
rect 17590 9802 17650 9862
rect 18604 10036 18664 10096
rect 13398 8872 13458 8932
rect 14536 8872 14596 8932
rect 13286 8672 13346 8732
rect 13180 8570 13240 8630
rect 13070 5118 13130 5178
rect 13286 7436 13346 7496
rect 13290 6910 13350 6970
rect 14534 8672 14594 8732
rect 15552 8792 15612 8852
rect 19626 10140 19686 10200
rect 29806 11352 29866 11412
rect 28278 11242 28338 11302
rect 29292 11242 29352 11302
rect 28792 11136 28852 11196
rect 25732 10140 25792 10200
rect 21662 10036 21722 10096
rect 23700 10036 23760 10096
rect 20646 9914 20706 9974
rect 22680 9914 22740 9974
rect 24710 9914 24770 9974
rect 16570 8896 16630 8956
rect 16066 8678 16126 8738
rect 17592 8792 17652 8852
rect 17070 8678 17130 8738
rect 14534 7640 14594 7700
rect 15040 7538 15100 7598
rect 18606 8896 18666 8956
rect 18082 8678 18142 8738
rect 19624 8792 19684 8852
rect 19102 8678 19162 8738
rect 19624 8680 19684 8740
rect 21658 8792 21718 8852
rect 20642 8570 20702 8630
rect 16572 7640 16632 7700
rect 16570 7436 16630 7496
rect 21660 8680 21720 8740
rect 22676 8570 22736 8630
rect 26750 10036 26810 10096
rect 30310 11242 30370 11302
rect 31842 11352 31902 11412
rect 31334 11242 31394 11302
rect 30822 11136 30882 11196
rect 30822 11032 30882 11092
rect 27768 10036 27828 10096
rect 28788 10036 28848 10096
rect 23698 8792 23758 8852
rect 23696 8680 23756 8740
rect 25732 8792 25792 8852
rect 25928 8788 25988 8848
rect 24716 8570 24776 8630
rect 25732 8680 25792 8740
rect 32354 11242 32414 11302
rect 32862 11136 32922 11196
rect 33998 11032 34058 11092
rect 30826 10140 30886 10200
rect 29804 10036 29864 10096
rect 31840 10036 31900 10096
rect 26750 8896 26810 8956
rect 25928 8570 25988 8630
rect 26222 8572 26282 8632
rect 18608 7640 18668 7700
rect 15554 7336 15614 7396
rect 17078 7430 17138 7490
rect 18100 7430 18160 7490
rect 17588 7336 17648 7396
rect 20640 7640 20700 7700
rect 20132 7538 20192 7598
rect 19114 7430 19174 7490
rect 20132 7430 20192 7490
rect 19624 7336 19684 7396
rect 15036 6412 15096 6472
rect 15946 6412 16006 6472
rect 15036 6196 15096 6256
rect 13400 6092 13460 6152
rect 13288 5326 13348 5386
rect 12838 4968 12898 5028
rect 13180 5080 13240 5140
rect 13286 4670 13346 4730
rect 16948 6412 17008 6472
rect 16074 6196 16134 6256
rect 18100 6412 18160 6472
rect 17588 6310 17648 6370
rect 17088 6196 17148 6256
rect 15034 5184 15094 5244
rect 14536 5080 14596 5140
rect 14532 4870 14592 4930
rect 16042 5184 16102 5244
rect 15552 4968 15612 5028
rect 21152 7430 21212 7490
rect 27766 8680 27826 8740
rect 27250 8572 27310 8632
rect 27768 8566 27828 8626
rect 28786 8896 28846 8956
rect 29804 8680 29864 8740
rect 30820 8788 30880 8848
rect 31324 8784 31384 8844
rect 33984 9802 34044 9862
rect 31844 8680 31904 8740
rect 29804 8566 29864 8626
rect 25222 7652 25282 7712
rect 24716 7524 24776 7584
rect 26752 7326 26812 7386
rect 19110 6412 19170 6472
rect 20116 6412 20176 6472
rect 21160 6412 21220 6472
rect 21660 6418 21720 6478
rect 20114 6196 20174 6256
rect 21154 6196 21214 6256
rect 20638 6092 20698 6152
rect 17056 5184 17116 5244
rect 18094 5184 18154 5244
rect 17590 4968 17650 5028
rect 16570 4870 16630 4930
rect 22168 6196 22228 6256
rect 23696 6418 23756 6478
rect 23176 6196 23236 6256
rect 24220 6196 24280 6256
rect 22680 6092 22740 6152
rect 31842 8566 31902 8626
rect 28264 7430 28324 7490
rect 25732 6418 25792 6478
rect 25210 6196 25270 6256
rect 26228 6196 26288 6256
rect 24718 6092 24778 6152
rect 32860 8896 32920 8956
rect 33878 8914 33938 8974
rect 34112 9784 34172 9844
rect 34478 8784 34538 8844
rect 34228 8680 34288 8740
rect 30316 7652 30376 7712
rect 30454 7656 30514 7716
rect 33984 8566 34044 8626
rect 31336 7656 31396 7716
rect 32342 7656 32402 7716
rect 29294 7430 29354 7490
rect 30454 7430 30514 7490
rect 30822 7430 30882 7490
rect 30822 7326 30882 7386
rect 32860 7652 32920 7712
rect 32860 7524 32920 7584
rect 31838 7328 31898 7388
rect 27770 6418 27830 6478
rect 27762 6310 27822 6370
rect 27262 6196 27322 6256
rect 26752 6092 26812 6152
rect 27264 6088 27324 6148
rect 28286 6088 28346 6148
rect 28786 6094 28846 6154
rect 19112 5184 19172 5244
rect 19628 5190 19688 5250
rect 21664 5190 21724 5250
rect 23696 5190 23756 5250
rect 25730 5190 25790 5250
rect 18610 4870 18670 4930
rect 13398 3848 13458 3908
rect 14538 3632 14598 3692
rect 15552 3946 15612 4006
rect 15556 3752 15616 3812
rect 16570 3848 16630 3908
rect 22680 5080 22740 5140
rect 24716 5080 24776 5140
rect 21662 4968 21722 5028
rect 20646 4870 20706 4930
rect 17588 3946 17648 4006
rect 18094 3848 18154 3908
rect 17592 3752 17652 3812
rect 19626 3946 19686 4006
rect 19116 3848 19176 3908
rect 18606 3632 18666 3692
rect 13286 2716 13346 2776
rect 13180 2590 13240 2650
rect 20138 3848 20198 3908
rect 19620 3752 19680 3812
rect 29806 6418 29866 6478
rect 29802 6310 29862 6370
rect 30294 6196 30354 6256
rect 31844 6418 31904 6478
rect 31840 6310 31900 6370
rect 31332 6196 31392 6256
rect 30820 6094 30880 6154
rect 26752 5192 26812 5252
rect 27106 5192 27166 5252
rect 26748 5080 26808 5140
rect 26258 4982 26318 5042
rect 21488 3966 21548 4026
rect 21658 3966 21718 4026
rect 21142 3848 21202 3908
rect 20640 3632 20700 3692
rect 16570 2590 16630 2650
rect 17090 2602 17150 2662
rect 15552 2488 15612 2548
rect 17588 2488 17648 2548
rect 16570 2384 16630 2444
rect 13398 1486 13458 1546
rect 13070 1382 13130 1442
rect 14534 1382 14594 1442
rect 15042 1276 15102 1336
rect 12020 322 12080 382
rect 21488 3752 21548 3812
rect 21664 3758 21724 3818
rect 27296 4982 27356 5042
rect 28272 4982 28332 5042
rect 27106 4874 27166 4934
rect 32358 6196 32418 6256
rect 32862 6094 32922 6154
rect 30824 5192 30884 5252
rect 29288 4982 29348 5042
rect 31314 4982 31374 5042
rect 28786 4870 28846 4930
rect 30822 4870 30882 4930
rect 23700 3966 23760 4026
rect 25732 3966 25792 4026
rect 27772 3966 27832 4026
rect 26750 3868 26810 3928
rect 23692 3758 23752 3818
rect 18608 2488 18668 2548
rect 19624 2488 19684 2548
rect 16568 1486 16628 1546
rect 16574 1382 16634 1442
rect 16062 1276 16122 1336
rect 15554 1166 15614 1226
rect 17086 1276 17146 1336
rect 20644 2488 20704 2548
rect 25736 3758 25796 3818
rect 27764 3758 27824 3818
rect 28790 3632 28850 3692
rect 32344 4982 32404 5042
rect 32858 4870 32918 4930
rect 29802 3758 29862 3818
rect 32856 3868 32916 3928
rect 31842 3758 31902 3818
rect 32360 3762 32420 3822
rect 33872 3762 33932 3822
rect 30820 3632 30880 3692
rect 31346 3634 31406 3694
rect 22674 2716 22734 2776
rect 24716 2716 24776 2776
rect 26752 2716 26812 2776
rect 22170 2602 22230 2662
rect 27258 2606 27318 2666
rect 21662 2488 21722 2548
rect 23692 2488 23752 2548
rect 25730 2488 25790 2548
rect 27766 2488 27826 2548
rect 21506 2384 21566 2444
rect 18604 1382 18664 1442
rect 18104 1276 18164 1336
rect 19118 1276 19178 1336
rect 17590 1166 17650 1226
rect 13398 244 13458 304
rect 14534 244 14594 304
rect 15046 136 15106 196
rect 20798 1488 20858 1548
rect 20644 1382 20704 1442
rect 20150 1276 20210 1336
rect 19628 1166 19688 1226
rect 16060 136 16120 196
rect 17082 136 17142 196
rect 21162 1276 21222 1336
rect 22676 1488 22736 1548
rect 22680 1382 22740 1442
rect 22170 1276 22230 1336
rect 21666 1166 21726 1226
rect 18604 244 18664 304
rect 18096 136 18156 196
rect 19122 136 19182 196
rect 23188 1276 23248 1336
rect 24714 1488 24774 1548
rect 24716 1382 24776 1442
rect 24214 1276 24274 1336
rect 23702 1166 23762 1226
rect 20134 136 20194 196
rect 21170 136 21230 196
rect 25216 1276 25276 1336
rect 27912 2384 27972 2444
rect 32860 3634 32920 3694
rect 28788 2488 28848 2548
rect 29806 2716 29866 2776
rect 29808 2488 29868 2548
rect 26584 1488 26644 1548
rect 26236 1276 26296 1336
rect 26750 1382 26810 1442
rect 25738 1166 25798 1226
rect 22176 136 22236 196
rect 23190 136 23250 196
rect 27256 1276 27316 1336
rect 30822 2488 30882 2548
rect 30822 2384 30882 2444
rect 31838 2716 31898 2776
rect 34112 7652 34172 7712
rect 34350 7430 34410 7490
rect 34228 7328 34288 7388
rect 34112 6094 34172 6154
rect 34108 5192 34168 5252
rect 34228 3966 34288 4026
rect 34108 3868 34168 3928
rect 33984 2716 34044 2776
rect 32358 2606 32418 2666
rect 33366 2606 33426 2666
rect 34476 6196 34536 6256
rect 34478 3762 34538 3822
rect 34350 3634 34410 3694
rect 34712 9784 34772 9844
rect 34600 2606 34660 2666
rect 31844 2488 31904 2548
rect 28790 1382 28850 1442
rect 28282 1276 28342 1336
rect 29300 1276 29360 1336
rect 27770 1166 27830 1226
rect 24206 136 24266 196
rect 25214 136 25274 196
rect 30820 1382 30880 1442
rect 30314 1276 30374 1336
rect 29802 1166 29862 1226
rect 26230 136 26290 196
rect 27254 136 27314 196
rect 31328 1276 31388 1336
rect 34004 2384 34064 2444
rect 32860 1488 32920 1548
rect 32860 1382 32920 1442
rect 32350 1276 32410 1336
rect 31842 1166 31902 1226
rect 28784 244 28844 304
rect 28276 136 28336 196
rect 29298 136 29358 196
rect 30316 136 30376 196
rect 31330 136 31390 196
rect 34712 1382 34772 1442
rect 34004 244 34064 304
rect 32354 136 32414 196
rect 53838 14952 53898 15012
rect 54166 14962 54226 15022
rect 53232 14816 53292 14876
rect 53352 14818 53412 14878
rect 53492 14836 53552 14896
rect 53720 14852 53780 14912
rect 53100 14688 53160 14748
rect 36824 13564 37424 13864
rect 37976 13564 38576 13864
rect 36928 13300 38480 13396
rect 37672 13134 37732 13194
rect 37156 12600 37216 12660
rect 38186 12600 38246 12660
rect -1198 -100 -1188 -76
rect -1188 -100 -1154 -76
rect -1154 -96 -872 -76
rect -872 -96 -836 -76
rect -836 -96 -814 -76
rect -1154 -100 -814 -96
rect -1198 -102 -814 -100
rect -1198 -136 -1116 -102
rect -1116 -136 -916 -102
rect -916 -136 -814 -102
rect -1198 -142 -814 -136
rect 2878 -260 34878 -106
rect -1266 -746 -666 -446
rect 35166 -746 35766 -446
rect 50388 14090 50448 14150
rect 51914 13956 51974 14016
rect 53100 7488 53160 7548
rect 48552 6562 48612 6622
rect 42442 6416 42502 6476
rect 46522 6416 46582 6476
rect 41288 6288 41348 6348
rect 43966 6288 44026 6348
rect 44998 6288 45058 6348
rect 42946 5326 43006 5386
rect 41288 5192 41348 5252
rect 42446 5222 42506 5282
rect 43970 5326 44030 5386
rect 43464 5118 43524 5178
rect 41288 4056 41348 4116
rect 48058 6288 48118 6348
rect 45002 5326 45062 5386
rect 44482 5222 44542 5282
rect 50582 6416 50642 6476
rect 52766 6416 52826 6476
rect 49054 6288 49114 6348
rect 46002 5326 46062 5386
rect 47022 5326 47082 5386
rect 46518 5222 46578 5282
rect 45500 5118 45560 5178
rect 42938 4056 42998 4116
rect 44476 4176 44536 4236
rect 48042 5326 48102 5386
rect 47532 5118 47592 5178
rect 46008 4056 46068 4116
rect 49052 5326 49112 5386
rect 48552 5222 48612 5282
rect 50066 5326 50126 5386
rect 51084 5326 51144 5386
rect 50588 5222 50648 5282
rect 49566 5118 49626 5178
rect 47016 4056 47076 4116
rect 43464 3112 43524 3172
rect 42450 3004 42510 3064
rect 42944 2892 43004 2952
rect 44486 3004 44546 3064
rect 43968 2892 44028 2952
rect 48552 4176 48612 4236
rect 45500 3112 45560 3172
rect 45000 2892 45060 2952
rect 51610 5118 51670 5178
rect 50078 4056 50138 4116
rect 52886 5326 52946 5386
rect 52766 4176 52826 4236
rect 51104 4056 51164 4116
rect 47532 3112 47592 3172
rect 46522 3004 46582 3064
rect 46000 2892 46060 2952
rect 47020 2892 47080 2952
rect 48556 3004 48616 3064
rect 48040 2892 48100 2952
rect 41288 1930 41348 1990
rect 43958 1930 44018 1990
rect 44990 1930 45050 1990
rect 49050 2892 49110 2952
rect 49566 3112 49626 3172
rect 51610 3112 51670 3172
rect 50592 3004 50652 3064
rect 50064 2892 50124 2952
rect 51082 2892 51142 2952
rect 48050 1930 48110 1990
rect 49046 1930 49106 1990
rect 52886 2892 52946 2952
rect 42444 1800 42504 1860
rect 46524 1800 46584 1860
rect 50584 1800 50644 1860
rect 52766 1800 52826 1860
rect 43922 434 43982 494
rect 45960 434 46020 494
rect 47996 434 48056 494
rect 44940 322 45000 382
rect 50032 434 50092 494
rect 49014 322 49074 382
rect 53232 6416 53292 6476
rect 53352 6288 53412 6348
rect 53610 14698 53670 14758
rect 53720 13956 53780 14016
rect 54286 14954 54346 15014
rect 54166 14090 54226 14150
rect 53962 12732 54022 12792
rect 53836 11030 53896 11090
rect 53610 8570 53670 8630
rect 53492 5326 53552 5386
rect 54174 12396 54234 12456
rect 54070 11136 54130 11196
rect 53962 10036 54022 10096
rect 54392 14818 54452 14878
rect 65204 14468 65264 14528
rect 70308 14468 70368 14528
rect 74368 14462 74428 14522
rect 55536 12732 55596 12792
rect 56550 12516 56610 12576
rect 58590 12516 58650 12576
rect 60630 12516 60690 12576
rect 62660 12516 62720 12576
rect 64700 12516 64760 12576
rect 66732 12516 66792 12576
rect 68772 12516 68832 12576
rect 70808 12516 70868 12576
rect 72842 12516 72902 12576
rect 54518 12396 54578 12456
rect 56042 12390 56102 12450
rect 54392 12274 54452 12334
rect 57056 12390 57116 12450
rect 58078 12390 58138 12450
rect 59092 12390 59152 12450
rect 60118 12390 60178 12450
rect 59606 12274 59666 12334
rect 61130 12390 61190 12450
rect 62166 12390 62226 12450
rect 63172 12390 63232 12450
rect 64186 12390 64246 12450
rect 56554 11352 56614 11412
rect 56046 11242 56106 11302
rect 55536 11136 55596 11196
rect 54522 11030 54582 11090
rect 55020 11030 55080 11090
rect 55532 11030 55592 11090
rect 57068 11242 57128 11302
rect 58594 11352 58654 11412
rect 58082 11242 58142 11302
rect 57576 11136 57636 11196
rect 60626 11352 60686 11412
rect 59096 11242 59156 11302
rect 60114 11242 60174 11302
rect 59606 11136 59666 11196
rect 54392 10140 54452 10200
rect 54516 10036 54576 10096
rect 56036 10036 56096 10096
rect 56548 10036 56608 10096
rect 54286 9914 54346 9974
rect 54174 9800 54234 9860
rect 55022 9800 55082 9860
rect 56554 9802 56614 9862
rect 61140 11242 61200 11302
rect 65202 12390 65262 12450
rect 66210 12390 66270 12450
rect 67226 12390 67286 12450
rect 68250 12390 68310 12450
rect 69272 12390 69332 12450
rect 70294 12390 70354 12450
rect 69794 12274 69854 12334
rect 62658 11352 62718 11412
rect 61646 11136 61706 11196
rect 62160 11242 62220 11302
rect 61812 11030 61872 11090
rect 57570 10140 57630 10200
rect 57572 10036 57632 10096
rect 63180 11242 63240 11302
rect 64694 11352 64754 11412
rect 64182 11242 64242 11302
rect 63680 11136 63740 11196
rect 63680 11030 63740 11090
rect 65208 11242 65268 11302
rect 71312 12390 71372 12450
rect 72326 12390 72386 12450
rect 73350 12390 73410 12450
rect 73866 12274 73926 12334
rect 74998 12274 75058 12334
rect 66730 11352 66790 11412
rect 66226 11242 66286 11302
rect 65716 11136 65776 11196
rect 65718 11030 65778 11090
rect 67234 11242 67294 11302
rect 68768 11352 68828 11412
rect 68246 11242 68306 11302
rect 67752 11136 67812 11196
rect 67598 11030 67658 11090
rect 58584 10036 58644 10096
rect 58590 9802 58650 9862
rect 59604 10036 59664 10096
rect 54398 8872 54458 8932
rect 55536 8872 55596 8932
rect 54286 8672 54346 8732
rect 54180 8570 54240 8630
rect 54070 5118 54130 5178
rect 54286 7436 54346 7496
rect 53838 4968 53898 5028
rect 54180 5080 54240 5140
rect 55534 8672 55594 8732
rect 56552 8792 56612 8852
rect 60626 10140 60686 10200
rect 70806 11352 70866 11412
rect 69278 11242 69338 11302
rect 70292 11242 70352 11302
rect 69792 11136 69852 11196
rect 66732 10140 66792 10200
rect 62662 10036 62722 10096
rect 64700 10036 64760 10096
rect 61646 9914 61706 9974
rect 63680 9914 63740 9974
rect 65710 9914 65770 9974
rect 57570 8896 57630 8956
rect 57066 8678 57126 8738
rect 58592 8792 58652 8852
rect 58070 8678 58130 8738
rect 55534 7640 55594 7700
rect 56040 7538 56100 7598
rect 59606 8896 59666 8956
rect 59082 8678 59142 8738
rect 60624 8792 60684 8852
rect 60102 8678 60162 8738
rect 60624 8680 60684 8740
rect 62658 8792 62718 8852
rect 61642 8570 61702 8630
rect 57572 7640 57632 7700
rect 57570 7436 57630 7496
rect 62660 8680 62720 8740
rect 63676 8570 63736 8630
rect 67750 10036 67810 10096
rect 71310 11242 71370 11302
rect 72842 11352 72902 11412
rect 72334 11242 72394 11302
rect 71822 11136 71882 11196
rect 71822 11032 71882 11092
rect 68768 10036 68828 10096
rect 69788 10036 69848 10096
rect 64698 8792 64758 8852
rect 64696 8680 64756 8740
rect 66732 8792 66792 8852
rect 66928 8788 66988 8848
rect 65716 8570 65776 8630
rect 66732 8680 66792 8740
rect 73354 11242 73414 11302
rect 73862 11136 73922 11196
rect 74998 11032 75058 11092
rect 71826 10140 71886 10200
rect 70804 10036 70864 10096
rect 72840 10036 72900 10096
rect 67750 8896 67810 8956
rect 66928 8570 66988 8630
rect 67222 8572 67282 8632
rect 59608 7640 59668 7700
rect 56554 7336 56614 7396
rect 58078 7430 58138 7490
rect 59100 7430 59160 7490
rect 58588 7336 58648 7396
rect 61640 7640 61700 7700
rect 61132 7538 61192 7598
rect 60114 7430 60174 7490
rect 61132 7430 61192 7490
rect 60624 7336 60684 7396
rect 56036 6412 56096 6472
rect 56946 6412 57006 6472
rect 56036 6196 56096 6256
rect 54400 6092 54460 6152
rect 57948 6412 58008 6472
rect 57074 6196 57134 6256
rect 59100 6412 59160 6472
rect 58588 6310 58648 6370
rect 58088 6196 58148 6256
rect 56034 5184 56094 5244
rect 55536 5080 55596 5140
rect 55532 4870 55592 4930
rect 57042 5184 57102 5244
rect 56552 4968 56612 5028
rect 62152 7430 62212 7490
rect 68766 8680 68826 8740
rect 68250 8572 68310 8632
rect 68768 8566 68828 8626
rect 69786 8896 69846 8956
rect 70804 8680 70864 8740
rect 71820 8788 71880 8848
rect 72324 8784 72384 8844
rect 74984 9802 75044 9862
rect 72844 8680 72904 8740
rect 70804 8566 70864 8626
rect 66222 7652 66282 7712
rect 65716 7524 65776 7584
rect 67752 7326 67812 7386
rect 60110 6412 60170 6472
rect 61116 6412 61176 6472
rect 62160 6412 62220 6472
rect 62660 6418 62720 6478
rect 61114 6196 61174 6256
rect 62154 6196 62214 6256
rect 61638 6092 61698 6152
rect 58056 5184 58116 5244
rect 59094 5184 59154 5244
rect 58590 4968 58650 5028
rect 57570 4870 57630 4930
rect 63168 6196 63228 6256
rect 64696 6418 64756 6478
rect 64176 6196 64236 6256
rect 65220 6196 65280 6256
rect 63680 6092 63740 6152
rect 72842 8566 72902 8626
rect 69264 7430 69324 7490
rect 66732 6418 66792 6478
rect 66210 6196 66270 6256
rect 67228 6196 67288 6256
rect 65718 6092 65778 6152
rect 73860 8896 73920 8956
rect 74878 8914 74938 8974
rect 75112 9784 75172 9844
rect 75478 8784 75538 8844
rect 75228 8680 75288 8740
rect 71316 7652 71376 7712
rect 71454 7656 71514 7716
rect 74984 8566 75044 8626
rect 72336 7656 72396 7716
rect 73342 7656 73402 7716
rect 70294 7430 70354 7490
rect 71454 7430 71514 7490
rect 71822 7430 71882 7490
rect 71822 7326 71882 7386
rect 73860 7652 73920 7712
rect 73860 7524 73920 7584
rect 72838 7328 72898 7388
rect 68770 6418 68830 6478
rect 68762 6310 68822 6370
rect 68262 6196 68322 6256
rect 67752 6092 67812 6152
rect 68264 6088 68324 6148
rect 69286 6088 69346 6148
rect 69786 6094 69846 6154
rect 60112 5184 60172 5244
rect 60628 5190 60688 5250
rect 62664 5190 62724 5250
rect 64696 5190 64756 5250
rect 66730 5190 66790 5250
rect 59610 4870 59670 4930
rect 54398 3848 54458 3908
rect 55538 3632 55598 3692
rect 56552 3946 56612 4006
rect 56556 3752 56616 3812
rect 57570 3848 57630 3908
rect 63680 5080 63740 5140
rect 65716 5080 65776 5140
rect 62662 4968 62722 5028
rect 61646 4870 61706 4930
rect 58588 3946 58648 4006
rect 59094 3848 59154 3908
rect 58592 3752 58652 3812
rect 60626 3946 60686 4006
rect 60116 3848 60176 3908
rect 59606 3632 59666 3692
rect 54286 2716 54346 2776
rect 54180 2590 54240 2650
rect 61138 3848 61198 3908
rect 60620 3752 60680 3812
rect 70806 6418 70866 6478
rect 70802 6310 70862 6370
rect 71294 6196 71354 6256
rect 72844 6418 72904 6478
rect 72840 6310 72900 6370
rect 72332 6196 72392 6256
rect 71820 6094 71880 6154
rect 67752 5192 67812 5252
rect 68106 5192 68166 5252
rect 67748 5080 67808 5140
rect 67258 4982 67318 5042
rect 62488 3966 62548 4026
rect 62658 3966 62718 4026
rect 62142 3848 62202 3908
rect 61640 3632 61700 3692
rect 57570 2590 57630 2650
rect 58090 2602 58150 2662
rect 56552 2488 56612 2548
rect 58588 2488 58648 2548
rect 57570 2384 57630 2444
rect 54398 1486 54458 1546
rect 54070 1382 54130 1442
rect 55534 1382 55594 1442
rect 56042 1276 56102 1336
rect 53020 322 53080 382
rect 62488 3752 62548 3812
rect 62664 3758 62724 3818
rect 68296 4982 68356 5042
rect 69272 4982 69332 5042
rect 68106 4874 68166 4934
rect 73358 6196 73418 6256
rect 73862 6094 73922 6154
rect 71824 5192 71884 5252
rect 70288 4982 70348 5042
rect 72314 4982 72374 5042
rect 69786 4870 69846 4930
rect 71822 4870 71882 4930
rect 64700 3966 64760 4026
rect 66732 3966 66792 4026
rect 68772 3966 68832 4026
rect 67750 3868 67810 3928
rect 64692 3758 64752 3818
rect 59608 2488 59668 2548
rect 60624 2488 60684 2548
rect 57568 1486 57628 1546
rect 57574 1382 57634 1442
rect 57062 1276 57122 1336
rect 56554 1166 56614 1226
rect 58086 1276 58146 1336
rect 61644 2488 61704 2548
rect 66736 3758 66796 3818
rect 68764 3758 68824 3818
rect 69790 3632 69850 3692
rect 73344 4982 73404 5042
rect 73858 4870 73918 4930
rect 70802 3758 70862 3818
rect 73856 3868 73916 3928
rect 72842 3758 72902 3818
rect 73360 3762 73420 3822
rect 74872 3762 74932 3822
rect 71820 3632 71880 3692
rect 72346 3634 72406 3694
rect 63674 2716 63734 2776
rect 65716 2716 65776 2776
rect 67752 2716 67812 2776
rect 63170 2602 63230 2662
rect 68258 2606 68318 2666
rect 62662 2488 62722 2548
rect 64692 2488 64752 2548
rect 66730 2488 66790 2548
rect 68766 2488 68826 2548
rect 62506 2384 62566 2444
rect 59604 1382 59664 1442
rect 59104 1276 59164 1336
rect 60118 1276 60178 1336
rect 58590 1166 58650 1226
rect 54398 244 54458 304
rect 55534 244 55594 304
rect 56046 136 56106 196
rect 61798 1488 61858 1548
rect 61644 1382 61704 1442
rect 61150 1276 61210 1336
rect 60628 1166 60688 1226
rect 57060 136 57120 196
rect 58082 136 58142 196
rect 62162 1276 62222 1336
rect 63676 1488 63736 1548
rect 63680 1382 63740 1442
rect 63170 1276 63230 1336
rect 62666 1166 62726 1226
rect 59604 244 59664 304
rect 59096 136 59156 196
rect 60122 136 60182 196
rect 64188 1276 64248 1336
rect 65714 1488 65774 1548
rect 65716 1382 65776 1442
rect 65214 1276 65274 1336
rect 64702 1166 64762 1226
rect 61134 136 61194 196
rect 62170 136 62230 196
rect 66216 1276 66276 1336
rect 68912 2384 68972 2444
rect 73860 3634 73920 3694
rect 69788 2488 69848 2548
rect 70806 2716 70866 2776
rect 70808 2488 70868 2548
rect 67584 1488 67644 1548
rect 67236 1276 67296 1336
rect 67750 1382 67810 1442
rect 66738 1166 66798 1226
rect 63176 136 63236 196
rect 64190 136 64250 196
rect 68256 1276 68316 1336
rect 71822 2488 71882 2548
rect 71822 2384 71882 2444
rect 72838 2716 72898 2776
rect 75112 7652 75172 7712
rect 75350 7430 75410 7490
rect 75228 7328 75288 7388
rect 75112 6094 75172 6154
rect 75108 5192 75168 5252
rect 75228 3966 75288 4026
rect 75108 3868 75168 3928
rect 74984 2716 75044 2776
rect 73358 2606 73418 2666
rect 74366 2606 74426 2666
rect 75476 6196 75536 6256
rect 75478 3762 75538 3822
rect 75350 3634 75410 3694
rect 75712 9784 75772 9844
rect 75600 2606 75660 2666
rect 72844 2488 72904 2548
rect 69790 1382 69850 1442
rect 69282 1276 69342 1336
rect 70300 1276 70360 1336
rect 68770 1166 68830 1226
rect 65206 136 65266 196
rect 66214 136 66274 196
rect 71820 1382 71880 1442
rect 71314 1276 71374 1336
rect 70802 1166 70862 1226
rect 67230 136 67290 196
rect 68254 136 68314 196
rect 72328 1276 72388 1336
rect 75004 2384 75064 2444
rect 73860 1488 73920 1548
rect 73860 1382 73920 1442
rect 73350 1276 73410 1336
rect 72842 1166 72902 1226
rect 69784 244 69844 304
rect 69276 136 69336 196
rect 70298 136 70358 196
rect 71316 136 71376 196
rect 72330 136 72390 196
rect 75712 1382 75772 1442
rect 75004 244 75064 304
rect 73354 136 73414 196
rect 43878 -260 75878 -106
rect 39734 -746 40334 -446
rect 76166 -746 76766 -446
<< metal2 >>
rect 11434 30586 12034 30596
rect 11434 30276 12034 30286
rect 35066 30586 35666 30596
rect 35066 30276 35666 30286
rect 52434 30586 53034 30596
rect 52434 30276 53034 30286
rect 76066 30586 76666 30596
rect 76066 30276 76666 30286
rect 14948 30204 31828 30236
rect 14948 29990 15011 30204
rect 31796 29990 31828 30204
rect 14948 29970 31828 29990
rect 55948 30204 72828 30236
rect 55948 29990 56011 30204
rect 72796 29990 72828 30204
rect 55948 29970 72828 29990
rect 14948 29968 19302 29970
rect 55948 29968 60302 29970
rect 18936 28288 18996 28294
rect 20018 28288 20078 28294
rect 20976 28288 21036 28294
rect 24040 28288 24100 28294
rect 25058 28288 25118 28294
rect 26082 28288 26142 28294
rect 27094 28288 27154 28294
rect 30152 28288 30212 28294
rect 31164 28288 31224 28294
rect 32182 28288 32242 28294
rect 18996 28228 20018 28288
rect 20078 28228 20976 28288
rect 21036 28228 24040 28288
rect 24100 28228 25058 28288
rect 25118 28228 26082 28288
rect 26142 28228 27094 28288
rect 27154 28228 30152 28288
rect 30212 28228 31164 28288
rect 31224 28228 32182 28288
rect 18936 28222 18996 28228
rect 20018 28222 20078 28228
rect 20976 28222 21036 28228
rect 24040 28222 24100 28228
rect 25058 28222 25118 28228
rect 26082 28222 26142 28228
rect 27094 28222 27154 28228
rect 30152 28222 30212 28228
rect 31164 28222 31224 28228
rect 32182 28222 32242 28228
rect 59936 28288 59996 28294
rect 61018 28288 61078 28294
rect 61976 28288 62036 28294
rect 65040 28288 65100 28294
rect 66058 28288 66118 28294
rect 67082 28288 67142 28294
rect 68094 28288 68154 28294
rect 71152 28288 71212 28294
rect 72164 28288 72224 28294
rect 73182 28288 73242 28294
rect 59996 28228 61018 28288
rect 61078 28228 61976 28288
rect 62036 28228 65040 28288
rect 65100 28228 66058 28288
rect 66118 28228 67082 28288
rect 67142 28228 68094 28288
rect 68154 28228 71152 28288
rect 71212 28228 72164 28288
rect 72224 28228 73182 28288
rect 59936 28222 59996 28228
rect 61018 28222 61078 28228
rect 61976 28222 62036 28228
rect 65040 28222 65100 28228
rect 66058 28222 66118 28228
rect 67082 28222 67142 28228
rect 68094 28222 68154 28228
rect 71152 28222 71212 28228
rect 72164 28222 72224 28228
rect 73182 28222 73242 28228
rect 19462 28042 19522 28048
rect 21498 28042 21558 28048
rect 23536 28044 23596 28050
rect 25566 28044 25626 28050
rect 27608 28046 27668 28052
rect 28618 28046 28678 28052
rect 29640 28046 29700 28052
rect 31676 28046 31736 28052
rect 19522 27982 21498 28042
rect 21558 27984 23536 28042
rect 23596 27984 25566 28044
rect 25626 27986 27608 28044
rect 27668 27986 28618 28046
rect 28678 27986 29640 28046
rect 29700 27986 31676 28046
rect 25626 27984 27806 27986
rect 21558 27982 23718 27984
rect 19462 27976 19522 27982
rect 21498 27976 21558 27982
rect 23536 27978 23596 27982
rect 25566 27978 25626 27984
rect 27608 27980 27668 27984
rect 28618 27980 28678 27986
rect 29640 27980 29700 27986
rect 31676 27980 31736 27986
rect 60462 28042 60522 28048
rect 62498 28042 62558 28048
rect 64536 28044 64596 28050
rect 66566 28044 66626 28050
rect 68608 28046 68668 28052
rect 69618 28046 69678 28052
rect 70640 28046 70700 28052
rect 72676 28046 72736 28052
rect 60522 27982 62498 28042
rect 62558 27984 64536 28042
rect 64596 27984 66566 28044
rect 66626 27986 68608 28044
rect 68668 27986 69618 28046
rect 69678 27986 70640 28046
rect 70700 27986 72676 28046
rect 66626 27984 68806 27986
rect 62558 27982 64718 27984
rect 60462 27976 60522 27982
rect 62498 27976 62558 27982
rect 64536 27978 64596 27982
rect 66566 27978 66626 27984
rect 68608 27980 68668 27984
rect 69618 27980 69678 27986
rect 70640 27980 70700 27986
rect 72676 27980 72736 27986
rect 17280 27110 17340 27116
rect 18444 27110 18504 27116
rect 24554 27110 24614 27116
rect 17340 27050 18444 27110
rect 18504 27050 24554 27110
rect 17280 27044 17340 27050
rect 18444 27044 18504 27050
rect 24554 27044 24614 27050
rect 26588 27110 26648 27116
rect 32696 27110 32756 27116
rect 33946 27110 34006 27116
rect 26648 27050 32696 27110
rect 32756 27050 33946 27110
rect 26588 27044 26648 27050
rect 32696 27044 32756 27050
rect 33946 27044 34006 27050
rect 58280 27110 58340 27116
rect 59444 27110 59504 27116
rect 65554 27110 65614 27116
rect 58340 27050 59444 27110
rect 59504 27050 65554 27110
rect 58280 27044 58340 27050
rect 59444 27044 59504 27050
rect 65554 27044 65614 27050
rect 67588 27110 67648 27116
rect 73696 27110 73756 27116
rect 74946 27110 75006 27116
rect 67648 27050 73696 27110
rect 73756 27050 74946 27110
rect 67588 27044 67648 27050
rect 73696 27044 73756 27050
rect 74946 27044 75006 27050
rect 20480 27006 20540 27012
rect 22516 27006 22576 27012
rect 28622 27006 28682 27012
rect 30656 27006 30716 27012
rect 20540 26946 22516 27006
rect 22576 26998 22994 27006
rect 23210 26998 28622 27006
rect 22576 26952 28622 26998
rect 22576 26948 25010 26952
rect 22576 26946 23984 26948
rect 24222 26946 25010 26948
rect 25226 26946 28622 26952
rect 28682 26946 30656 27006
rect 20480 26940 20540 26946
rect 22516 26940 22576 26946
rect 28622 26940 28682 26946
rect 30656 26940 30716 26946
rect 61480 27006 61540 27012
rect 63516 27006 63576 27012
rect 69622 27006 69682 27012
rect 71656 27006 71716 27012
rect 61540 26946 63516 27006
rect 63576 26998 63994 27006
rect 64210 26998 69622 27006
rect 63576 26952 69622 26998
rect 63576 26948 66010 26952
rect 63576 26946 64984 26948
rect 65222 26946 66010 26948
rect 66226 26946 69622 26952
rect 69682 26946 71656 27006
rect 61480 26940 61540 26946
rect 63516 26940 63576 26946
rect 69622 26940 69682 26946
rect 71656 26940 71716 26946
rect 17150 26906 17210 26912
rect 18444 26906 18504 26912
rect 24550 26906 24610 26912
rect 26586 26906 26646 26912
rect 17210 26846 18444 26906
rect 18504 26846 24550 26906
rect 24610 26846 26586 26906
rect 17150 26840 17210 26846
rect 18444 26840 18504 26846
rect 24550 26840 24610 26846
rect 26586 26840 26646 26846
rect 27088 26906 27148 26912
rect 28108 26906 28168 26912
rect 29134 26906 29194 26912
rect 27148 26846 28108 26906
rect 28168 26846 29134 26906
rect 27088 26840 27148 26846
rect 28108 26840 28168 26846
rect 29134 26840 29194 26846
rect 29640 26902 29700 26908
rect 30154 26902 30214 26908
rect 30658 26902 30718 26908
rect 31164 26902 31224 26908
rect 58150 26906 58210 26912
rect 59444 26906 59504 26912
rect 65550 26906 65610 26912
rect 67586 26906 67646 26912
rect 29700 26842 30154 26902
rect 30214 26842 30658 26902
rect 30718 26842 31164 26902
rect 31224 26842 31684 26902
rect 31744 26842 31750 26902
rect 58210 26846 59444 26906
rect 59504 26846 65550 26906
rect 65610 26846 67586 26906
rect 29640 26836 29700 26842
rect 30154 26836 30214 26842
rect 30658 26836 30718 26842
rect 31164 26836 31224 26842
rect 58150 26840 58210 26846
rect 59444 26840 59504 26846
rect 65550 26840 65610 26846
rect 67586 26840 67646 26846
rect 68088 26906 68148 26912
rect 69108 26906 69168 26912
rect 70134 26906 70194 26912
rect 68148 26846 69108 26906
rect 69168 26846 70134 26906
rect 68088 26840 68148 26846
rect 69108 26840 69168 26846
rect 70134 26840 70194 26846
rect 70640 26902 70700 26908
rect 71154 26902 71214 26908
rect 71658 26902 71718 26908
rect 72164 26902 72224 26908
rect 70700 26842 71154 26902
rect 71214 26842 71658 26902
rect 71718 26842 72164 26902
rect 72224 26842 72684 26902
rect 72744 26842 72750 26902
rect 70640 26836 70700 26842
rect 71154 26836 71214 26842
rect 71658 26836 71718 26842
rect 72164 26836 72224 26842
rect 21496 25972 21556 25978
rect 23530 25972 23590 25978
rect 25568 25972 25628 25976
rect 20980 25912 20986 25972
rect 21046 25912 21496 25972
rect 21556 25912 23530 25972
rect 23590 25970 25772 25972
rect 27604 25970 27664 25976
rect 28104 25970 28164 25976
rect 28618 25970 28678 25976
rect 29142 25970 29202 25976
rect 29640 25970 29700 25976
rect 30142 25970 30202 25976
rect 23590 25912 25568 25970
rect 21496 25906 21556 25912
rect 23530 25906 23590 25912
rect 25628 25910 27604 25970
rect 27664 25910 28104 25970
rect 28164 25910 28618 25970
rect 28678 25910 29142 25970
rect 29202 25910 29640 25970
rect 29700 25910 30142 25970
rect 30202 25968 30510 25970
rect 30656 25968 30716 25974
rect 31164 25968 31224 25974
rect 31674 25968 31734 25974
rect 62496 25972 62556 25978
rect 64530 25972 64590 25978
rect 66568 25972 66628 25976
rect 30202 25910 30656 25968
rect 25568 25904 25628 25910
rect 27604 25904 27664 25910
rect 28104 25904 28164 25910
rect 28618 25904 28678 25910
rect 29142 25904 29202 25910
rect 29539 25908 30054 25910
rect 29640 25904 29700 25908
rect 30142 25904 30202 25910
rect 30304 25908 30656 25910
rect 30716 25908 31164 25968
rect 31224 25908 31674 25968
rect 61980 25912 61986 25972
rect 62046 25912 62496 25972
rect 62556 25912 64530 25972
rect 64590 25970 66772 25972
rect 68604 25970 68664 25976
rect 69104 25970 69164 25976
rect 69618 25970 69678 25976
rect 70142 25970 70202 25976
rect 70640 25970 70700 25976
rect 71142 25970 71202 25976
rect 64590 25912 66568 25970
rect 30656 25902 30716 25908
rect 31164 25902 31224 25908
rect 31674 25902 31734 25908
rect 62496 25906 62556 25912
rect 64530 25906 64590 25912
rect 66628 25910 68604 25970
rect 68664 25910 69104 25970
rect 69164 25910 69618 25970
rect 69678 25910 70142 25970
rect 70202 25910 70640 25970
rect 70700 25910 71142 25970
rect 71202 25968 71510 25970
rect 71656 25968 71716 25974
rect 72164 25968 72224 25974
rect 72674 25968 72734 25974
rect 71202 25910 71656 25968
rect 66568 25904 66628 25910
rect 68604 25904 68664 25910
rect 69104 25904 69164 25910
rect 69618 25904 69678 25910
rect 70142 25904 70202 25910
rect 70539 25908 71054 25910
rect 70640 25904 70700 25908
rect 71142 25904 71202 25910
rect 71304 25908 71656 25910
rect 71716 25908 72164 25968
rect 72224 25908 72674 25968
rect 71656 25902 71716 25908
rect 72164 25902 72224 25908
rect 72674 25902 72734 25908
rect 20478 25874 20542 25880
rect 22354 25874 22418 25880
rect 20542 25810 22354 25874
rect 20478 25804 20542 25810
rect 22354 25804 22418 25810
rect 26588 25872 26648 25878
rect 32696 25872 32756 25878
rect 26648 25812 32696 25872
rect 26588 25806 26648 25812
rect 32696 25806 32756 25812
rect 61478 25874 61542 25880
rect 63354 25874 63418 25880
rect 61542 25810 63354 25874
rect 61478 25804 61542 25810
rect 63354 25804 63418 25810
rect 67588 25872 67648 25878
rect 73696 25872 73756 25878
rect 67648 25812 73696 25872
rect 67588 25806 67648 25812
rect 73696 25806 73756 25812
rect 21990 25764 22050 25770
rect 23014 25764 23074 25770
rect 24042 25764 24102 25770
rect 19968 25756 20028 25762
rect 20980 25756 21040 25762
rect 18924 25696 18930 25756
rect 18990 25696 19968 25756
rect 20028 25696 20980 25756
rect 22050 25704 23014 25764
rect 23074 25704 24042 25764
rect 62990 25764 63050 25770
rect 64014 25764 64074 25770
rect 65042 25764 65102 25770
rect 21990 25698 22050 25704
rect 23014 25698 23074 25704
rect 24042 25698 24102 25704
rect 30146 25756 30206 25762
rect 31158 25756 31218 25762
rect 32160 25756 32220 25762
rect 60968 25756 61028 25762
rect 61980 25756 62040 25762
rect 19968 25690 20028 25696
rect 20980 25690 21040 25696
rect 30206 25696 31158 25756
rect 31218 25696 32160 25756
rect 59924 25696 59930 25756
rect 59990 25696 60968 25756
rect 61028 25696 61980 25756
rect 63050 25704 64014 25764
rect 64074 25704 65042 25764
rect 62990 25698 63050 25704
rect 64014 25698 64074 25704
rect 65042 25698 65102 25704
rect 71146 25756 71206 25762
rect 72158 25756 72218 25762
rect 73160 25756 73220 25762
rect 30146 25690 30206 25696
rect 31158 25690 31218 25696
rect 32160 25690 32220 25696
rect 60968 25690 61028 25696
rect 61980 25690 62040 25696
rect 71206 25696 72158 25756
rect 72218 25696 73160 25756
rect 71146 25690 71206 25696
rect 72158 25690 72218 25696
rect 73160 25690 73220 25696
rect 19460 24834 19520 24840
rect 21496 24834 21556 24840
rect 22018 24834 22078 24840
rect 22516 24834 22576 24840
rect 23530 24834 23590 24840
rect 23990 24834 24050 24840
rect 25028 24834 25034 24836
rect 19520 24774 21496 24834
rect 21556 24774 22018 24834
rect 22078 24774 22516 24834
rect 22576 24832 23530 24834
rect 22576 24830 23498 24832
rect 22576 24774 22990 24830
rect 19460 24768 19520 24774
rect 21496 24768 21556 24774
rect 22018 24768 22078 24774
rect 22516 24768 22576 24774
rect 22984 24770 22990 24774
rect 23050 24774 23498 24830
rect 23590 24774 23990 24834
rect 24050 24776 25034 24834
rect 25094 24834 25100 24836
rect 25566 24834 25626 24840
rect 27072 24834 27078 24836
rect 25094 24776 25566 24834
rect 24050 24774 25566 24776
rect 25626 24776 27078 24834
rect 27138 24834 27144 24836
rect 27138 24832 27450 24834
rect 27604 24832 27664 24838
rect 29640 24832 29700 24836
rect 27138 24830 27604 24832
rect 27664 24830 29828 24832
rect 31674 24830 31734 24836
rect 27138 24776 27572 24830
rect 25626 24774 27572 24776
rect 23050 24770 23056 24774
rect 23492 24772 23498 24774
rect 23558 24772 23590 24774
rect 23530 24768 23590 24772
rect 23990 24768 24050 24774
rect 25566 24768 25626 24774
rect 25710 24772 27036 24774
rect 27242 24772 27572 24774
rect 27664 24826 28588 24830
rect 28648 24828 29640 24830
rect 27664 24772 28100 24826
rect 27566 24770 27572 24772
rect 27632 24770 27664 24772
rect 27604 24766 27664 24770
rect 28094 24766 28100 24772
rect 28160 24772 28588 24826
rect 28160 24766 28166 24772
rect 28582 24770 28588 24772
rect 28682 24826 29640 24828
rect 28682 24772 29100 24826
rect 28616 24768 28622 24770
rect 28682 24768 28688 24772
rect 29094 24766 29100 24772
rect 29160 24772 29640 24826
rect 29160 24766 29166 24772
rect 29700 24770 31674 24830
rect 29640 24764 29700 24770
rect 31674 24764 31734 24770
rect 60460 24834 60520 24840
rect 62496 24834 62556 24840
rect 63018 24834 63078 24840
rect 63516 24834 63576 24840
rect 64530 24834 64590 24840
rect 64990 24834 65050 24840
rect 66028 24834 66034 24836
rect 60520 24774 62496 24834
rect 62556 24774 63018 24834
rect 63078 24774 63516 24834
rect 63576 24832 64530 24834
rect 63576 24830 64498 24832
rect 63576 24774 63990 24830
rect 60460 24768 60520 24774
rect 62496 24768 62556 24774
rect 63018 24768 63078 24774
rect 63516 24768 63576 24774
rect 63984 24770 63990 24774
rect 64050 24774 64498 24830
rect 64590 24774 64990 24834
rect 65050 24776 66034 24834
rect 66094 24834 66100 24836
rect 66566 24834 66626 24840
rect 68072 24834 68078 24836
rect 66094 24776 66566 24834
rect 65050 24774 66566 24776
rect 66626 24776 68078 24834
rect 68138 24834 68144 24836
rect 68138 24832 68450 24834
rect 68604 24832 68664 24838
rect 70640 24832 70700 24836
rect 68138 24830 68604 24832
rect 68664 24830 70828 24832
rect 72674 24830 72734 24836
rect 68138 24776 68572 24830
rect 66626 24774 68572 24776
rect 64050 24770 64056 24774
rect 64492 24772 64498 24774
rect 64558 24772 64590 24774
rect 64530 24768 64590 24772
rect 64990 24768 65050 24774
rect 66566 24768 66626 24774
rect 66710 24772 68036 24774
rect 68242 24772 68572 24774
rect 68664 24826 69588 24830
rect 69648 24828 70640 24830
rect 68664 24772 69100 24826
rect 68566 24770 68572 24772
rect 68632 24770 68664 24772
rect 68604 24766 68664 24770
rect 69094 24766 69100 24772
rect 69160 24772 69588 24826
rect 69160 24766 69166 24772
rect 69582 24770 69588 24772
rect 69682 24826 70640 24828
rect 69682 24772 70100 24826
rect 69616 24768 69622 24770
rect 69682 24768 69688 24772
rect 70094 24766 70100 24772
rect 70160 24772 70640 24826
rect 70160 24766 70166 24772
rect 70700 24770 72674 24830
rect 70640 24764 70700 24770
rect 72674 24764 72734 24770
rect 15142 24724 15202 24728
rect 20476 24724 20540 24730
rect 30656 24724 30720 24730
rect 56142 24724 56202 24728
rect 61476 24724 61540 24730
rect 71656 24724 71720 24730
rect 15140 24722 20476 24724
rect 15140 24662 15142 24722
rect 15202 24662 20476 24722
rect 15140 24660 20476 24662
rect 20540 24660 30656 24724
rect 56140 24722 61476 24724
rect 56140 24662 56142 24722
rect 56202 24662 61476 24722
rect 56140 24660 61476 24662
rect 61540 24660 71656 24724
rect 15142 24656 15202 24660
rect 20476 24654 20540 24660
rect 30656 24654 30720 24660
rect 56142 24656 56202 24660
rect 61476 24654 61540 24660
rect 71656 24654 71720 24660
rect 18438 24586 18502 24592
rect 59438 24586 59502 24592
rect 18502 24582 33942 24586
rect 18502 24522 24548 24582
rect 18438 24516 18502 24522
rect 24542 24518 24548 24522
rect 24612 24522 33942 24582
rect 34006 24522 34012 24586
rect 59502 24582 74942 24586
rect 59502 24522 65548 24582
rect 24612 24518 24618 24522
rect 59438 24516 59502 24522
rect 65542 24518 65548 24522
rect 65612 24522 74942 24582
rect 75006 24522 75012 24586
rect 65612 24518 65618 24522
rect 17280 24436 17340 24442
rect 26584 24440 26648 24446
rect 17340 24376 18262 24436
rect 18322 24376 26584 24436
rect 32690 24436 32750 24442
rect 26648 24376 32690 24436
rect 17280 24370 17340 24376
rect 26584 24370 26648 24376
rect 32690 24370 32750 24376
rect 58280 24436 58340 24442
rect 67584 24440 67648 24446
rect 58340 24376 59262 24436
rect 59322 24376 67584 24436
rect 73690 24436 73750 24442
rect 67648 24376 73690 24436
rect 58280 24370 58340 24376
rect 67584 24370 67648 24376
rect 73690 24370 73750 24376
rect 18378 24330 18438 24336
rect 18940 24330 19000 24336
rect 19982 24330 20042 24336
rect 20982 24330 21042 24336
rect 24144 24330 24204 24336
rect 25154 24330 25214 24336
rect 26096 24330 26156 24336
rect 18438 24270 18940 24330
rect 19000 24270 19982 24330
rect 20042 24270 20982 24330
rect 21042 24270 24144 24330
rect 24204 24270 25154 24330
rect 25214 24270 26096 24330
rect 18378 24264 18438 24270
rect 18940 24264 19000 24270
rect 19982 24264 20042 24270
rect 20982 24264 21042 24270
rect 24144 24264 24204 24270
rect 25154 24264 25214 24270
rect 26096 24264 26156 24270
rect 59378 24330 59438 24336
rect 59940 24330 60000 24336
rect 60982 24330 61042 24336
rect 61982 24330 62042 24336
rect 65144 24330 65204 24336
rect 66154 24330 66214 24336
rect 67096 24330 67156 24336
rect 59438 24270 59940 24330
rect 60000 24270 60982 24330
rect 61042 24270 61982 24330
rect 62042 24270 65144 24330
rect 65204 24270 66154 24330
rect 66214 24270 67096 24330
rect 59378 24264 59438 24270
rect 59940 24264 60000 24270
rect 60982 24264 61042 24270
rect 61982 24264 62042 24270
rect 65144 24264 65204 24270
rect 66154 24264 66214 24270
rect 67096 24264 67156 24270
rect 18492 24128 18552 24134
rect 21670 24128 21730 24134
rect 25738 24128 25798 24134
rect 29814 24128 29874 24134
rect 33010 24128 33070 24134
rect 18552 24068 21670 24128
rect 21730 24068 25738 24128
rect 25798 24068 29814 24128
rect 29874 24068 33010 24128
rect 18492 24062 18552 24068
rect 21670 24062 21730 24068
rect 25738 24062 25798 24068
rect 29814 24062 29874 24068
rect 33010 24062 33070 24068
rect 59492 24128 59552 24134
rect 62670 24128 62730 24134
rect 66738 24128 66798 24134
rect 70814 24128 70874 24134
rect 74010 24128 74070 24134
rect 59552 24068 62670 24128
rect 62730 24068 66738 24128
rect 66798 24068 70814 24128
rect 70874 24068 74010 24128
rect 59492 24062 59552 24068
rect 62670 24062 62730 24068
rect 66738 24062 66798 24068
rect 70814 24062 70874 24068
rect 74010 24062 74070 24068
rect 19636 23192 19696 23198
rect 21670 23192 21730 23198
rect 23712 23192 23772 23198
rect 25738 23192 25798 23198
rect 27780 23192 27840 23198
rect 29816 23192 29876 23198
rect 31852 23192 31912 23198
rect 19696 23132 21670 23192
rect 21730 23132 23712 23192
rect 23772 23132 25738 23192
rect 25798 23132 27780 23192
rect 27840 23132 29816 23192
rect 29876 23132 31852 23192
rect 19636 23126 19696 23132
rect 21670 23126 21730 23132
rect 23712 23126 23772 23132
rect 25738 23126 25798 23132
rect 27780 23126 27840 23132
rect 29816 23126 29876 23132
rect 31852 23126 31912 23132
rect 60636 23192 60696 23198
rect 62670 23192 62730 23198
rect 64712 23192 64772 23198
rect 66738 23192 66798 23198
rect 68780 23192 68840 23198
rect 70816 23192 70876 23198
rect 72852 23192 72912 23198
rect 60696 23132 62670 23192
rect 62730 23132 64712 23192
rect 64772 23132 66738 23192
rect 66798 23132 68780 23192
rect 68840 23132 70816 23192
rect 70876 23132 72852 23192
rect 60636 23126 60696 23132
rect 62670 23126 62730 23132
rect 64712 23126 64772 23132
rect 66738 23126 66798 23132
rect 68780 23126 68840 23132
rect 70816 23126 70876 23132
rect 72852 23126 72912 23132
rect 20140 23084 20200 23090
rect 61140 23084 61200 23090
rect 20200 23024 21162 23084
rect 21222 23024 22180 23084
rect 22240 23024 23204 23084
rect 23264 23024 24218 23084
rect 24278 23024 25236 23084
rect 25296 23024 26246 23084
rect 26306 23024 27268 23084
rect 27328 23024 28282 23084
rect 28342 23024 29314 23084
rect 29374 23024 30324 23084
rect 30384 23024 31346 23084
rect 31406 23024 31412 23084
rect 61200 23024 62162 23084
rect 62222 23024 63180 23084
rect 63240 23024 64204 23084
rect 64264 23024 65218 23084
rect 65278 23024 66236 23084
rect 66296 23024 67246 23084
rect 67306 23024 68268 23084
rect 68328 23024 69282 23084
rect 69342 23024 70314 23084
rect 70374 23024 71324 23084
rect 71384 23024 72346 23084
rect 72406 23024 72412 23084
rect 20140 23018 20200 23024
rect 61140 23018 61200 23024
rect 19632 22160 19692 22166
rect 23712 22160 23772 22166
rect 27780 22160 27840 22166
rect 31848 22160 31908 22166
rect 34240 22160 34300 22166
rect 60632 22160 60692 22166
rect 64712 22160 64772 22166
rect 68780 22160 68840 22166
rect 72848 22160 72908 22166
rect 75240 22160 75300 22166
rect 12100 22100 19632 22160
rect 19692 22100 23712 22160
rect 23772 22100 27780 22160
rect 27840 22100 31848 22160
rect 31908 22100 34240 22160
rect -3042 15992 8228 16248
rect -3042 15700 -2680 15992
rect 8172 15700 8228 15992
rect -3042 15392 8228 15700
rect -3042 15070 9310 15392
rect 12100 14748 12160 22100
rect 19632 22094 19692 22100
rect 23712 22094 23772 22100
rect 27780 22094 27840 22100
rect 31848 22094 31908 22100
rect 34240 22094 34300 22100
rect 53100 22100 60632 22160
rect 60692 22100 64712 22160
rect 64772 22100 68780 22160
rect 68840 22100 72848 22160
rect 72908 22100 75240 22160
rect 17636 22028 17696 22034
rect 22178 22028 22184 22030
rect 17696 22026 22184 22028
rect 17696 21968 20138 22026
rect 17636 21962 17696 21968
rect 20132 21966 20138 21968
rect 20198 22022 22184 22026
rect 20198 21968 21152 22022
rect 20198 21966 20204 21968
rect 21146 21962 21152 21968
rect 21212 21970 22184 22022
rect 22244 22028 22250 22030
rect 23176 22028 23182 22030
rect 22244 21970 23182 22028
rect 23242 22028 23248 22030
rect 24220 22028 24226 22030
rect 23242 21970 24226 22028
rect 24286 22028 24292 22030
rect 28276 22028 28282 22030
rect 24286 22026 28282 22028
rect 24286 21970 25230 22026
rect 21212 21968 25230 21970
rect 21212 21962 21218 21968
rect 25224 21966 25230 21968
rect 25290 21968 26246 22026
rect 25290 21966 25296 21968
rect 26240 21966 26246 21968
rect 26306 21968 27250 22026
rect 26306 21966 26312 21968
rect 27244 21966 27250 21968
rect 27310 21970 28282 22026
rect 28342 22028 28348 22030
rect 33804 22028 33864 22034
rect 28342 22026 33804 22028
rect 28342 21970 29298 22026
rect 27310 21968 29298 21970
rect 27310 21966 27316 21968
rect 29292 21966 29298 21968
rect 29358 21968 30326 22026
rect 29358 21966 29364 21968
rect 30320 21966 30326 21968
rect 30386 21968 31346 22026
rect 30386 21966 30392 21968
rect 31340 21966 31346 21968
rect 31406 21968 33804 22026
rect 31406 21966 31412 21968
rect 33804 21962 33864 21968
rect 25030 21818 25090 21824
rect 25090 21758 26766 21818
rect 26826 21758 26832 21818
rect 32664 21804 32724 21808
rect 32662 21802 34006 21804
rect 25030 21752 25090 21758
rect 32662 21742 32664 21802
rect 32724 21800 34006 21802
rect 32724 21742 33946 21800
rect 32662 21740 33946 21742
rect 34006 21740 34012 21800
rect 32664 21736 32724 21740
rect 26046 21622 26110 21628
rect 30110 21622 30174 21628
rect 31134 21622 31198 21628
rect 32146 21622 32210 21628
rect 26110 21558 30110 21622
rect 30174 21558 31134 21622
rect 31198 21558 32146 21622
rect 26046 21552 26110 21558
rect 30110 21552 30174 21558
rect 31134 21552 31198 21558
rect 32146 21552 32210 21558
rect 18262 21500 18322 21506
rect 19428 21500 19488 21506
rect 21464 21500 21524 21506
rect 18322 21440 19428 21500
rect 19488 21440 21464 21500
rect 18262 21434 18322 21440
rect 19428 21434 19488 21440
rect 21464 21434 21524 21440
rect 21972 21500 22036 21506
rect 26048 21500 26112 21506
rect 22036 21436 26048 21500
rect 21972 21430 22036 21436
rect 26048 21430 26112 21436
rect 29610 21500 29670 21506
rect 31644 21500 31704 21506
rect 34088 21500 34148 21506
rect 29670 21440 31644 21500
rect 31704 21440 34088 21500
rect 29610 21434 29670 21440
rect 31644 21434 31704 21440
rect 34088 21434 34148 21440
rect 17510 21418 17570 21424
rect 17752 21418 17812 21424
rect 17570 21358 17752 21418
rect 17510 21352 17570 21358
rect 17752 21352 17812 21358
rect 20446 20552 20506 20558
rect 22482 20552 22542 20558
rect 20506 20492 22482 20552
rect 20446 20486 20506 20492
rect 22482 20486 22542 20492
rect 22824 20554 22884 20560
rect 25538 20554 25598 20560
rect 22884 20494 25538 20554
rect 22824 20488 22884 20494
rect 25538 20488 25598 20494
rect 30626 20552 30686 20558
rect 32662 20552 32722 20558
rect 30686 20492 32662 20552
rect 30626 20486 30686 20492
rect 14626 20464 14686 20470
rect 15648 20464 15708 20470
rect 14686 20404 15648 20464
rect 14626 20398 14686 20404
rect 15648 20398 15708 20404
rect 17994 20454 18054 20460
rect 30734 20454 30794 20492
rect 32662 20486 32722 20492
rect 18054 20394 30794 20454
rect 17994 20388 18054 20394
rect 14734 20352 14794 20358
rect 15518 20352 15578 20358
rect 14794 20292 15518 20352
rect 14734 20286 14794 20292
rect 15518 20286 15578 20292
rect 18130 20356 18190 20362
rect 20446 20356 20506 20362
rect 18190 20296 20446 20356
rect 18130 20290 18190 20296
rect 20446 20290 20506 20296
rect 21466 20358 21526 20364
rect 26556 20358 26616 20364
rect 33928 20358 33988 20364
rect 21526 20298 26556 20358
rect 26616 20298 33928 20358
rect 21466 20292 21526 20298
rect 26556 20292 26616 20298
rect 33928 20292 33988 20298
rect 19432 20246 19492 20252
rect 21466 20246 21526 20252
rect 19492 20186 21466 20246
rect 19432 20180 19492 20186
rect 21466 20180 21526 20186
rect 24522 20244 24582 20250
rect 26556 20244 26616 20250
rect 24582 20184 26556 20244
rect 24522 20178 24582 20184
rect 26556 20178 26616 20184
rect 29612 20244 29672 20250
rect 31646 20246 31706 20250
rect 31578 20244 31706 20246
rect 34240 20244 34300 20250
rect 29672 20184 31646 20244
rect 31706 20184 34240 20244
rect 29612 20178 29672 20184
rect 31578 20182 31706 20184
rect 31646 20178 31706 20182
rect 34240 20178 34300 20184
rect 12964 19430 13024 19436
rect 16158 19430 16218 19436
rect 13024 19370 16158 19430
rect 12964 19364 13024 19370
rect 16158 19364 16218 19370
rect 14124 19320 14184 19326
rect 17310 19320 17370 19326
rect 14184 19260 17310 19320
rect 30476 19310 30536 19316
rect 14124 19254 14184 19260
rect 17310 19254 17370 19260
rect 17752 19296 17812 19302
rect 24518 19296 24578 19302
rect 25538 19296 25598 19302
rect 27574 19296 27634 19302
rect 17812 19236 24518 19296
rect 24578 19236 25538 19296
rect 25598 19236 27574 19296
rect 30536 19250 34898 19310
rect 30476 19244 30536 19250
rect 17752 19230 17812 19236
rect 24518 19230 24578 19236
rect 25538 19230 25598 19236
rect 27574 19230 27634 19236
rect 30624 19200 30684 19206
rect 32664 19200 32724 19206
rect 33804 19200 33864 19206
rect 17502 19192 17562 19198
rect 22484 19192 22544 19198
rect 29608 19192 29668 19198
rect 17562 19132 20448 19192
rect 20508 19132 22484 19192
rect 22544 19132 29608 19192
rect 30684 19140 32664 19200
rect 32724 19140 33804 19200
rect 30624 19134 30684 19140
rect 32664 19134 32724 19140
rect 33804 19134 33864 19140
rect 17502 19126 17562 19132
rect 22484 19126 22544 19132
rect 29608 19126 29668 19132
rect 22482 19090 22542 19096
rect 31644 19090 31704 19096
rect 17748 19082 17808 19088
rect 18414 19082 18474 19088
rect 17808 19022 18414 19082
rect 22542 19030 31644 19090
rect 22482 19024 22542 19030
rect 31644 19024 31704 19030
rect 17748 19016 17808 19022
rect 18414 19016 18474 19022
rect 20448 18988 20508 18994
rect 22482 18988 22542 18994
rect 20508 18928 22482 18988
rect 20448 18922 20508 18928
rect 22482 18922 22542 18928
rect 25538 18990 25598 18996
rect 26556 18990 26616 18996
rect 27572 18990 27632 18996
rect 30476 18990 30536 18996
rect 25598 18930 26556 18990
rect 26616 18930 27572 18990
rect 27632 18930 30476 18990
rect 25538 18924 25598 18930
rect 26556 18924 26616 18930
rect 27572 18924 27632 18930
rect 30476 18924 30536 18930
rect 30628 18992 30688 18998
rect 32662 18992 32722 18998
rect 33928 18992 33988 18998
rect 30688 18932 32662 18992
rect 32722 18932 33928 18992
rect 33988 18932 34770 18992
rect 30628 18926 30688 18932
rect 32662 18926 32722 18932
rect 33928 18926 33988 18932
rect 14640 18396 14700 18402
rect 15650 18396 15710 18402
rect 12832 18282 12838 18342
rect 12898 18282 12904 18342
rect 14700 18336 15650 18396
rect 14640 18330 14700 18336
rect 15650 18330 15710 18336
rect 14746 18296 14806 18302
rect 15532 18296 15592 18302
rect 12346 17226 12352 17286
rect 12412 17226 12418 17286
rect 12226 16726 12232 16786
rect 12292 16726 12298 16786
rect 12232 14876 12292 16726
rect 12232 14810 12292 14816
rect 12352 14878 12412 17226
rect 12486 17050 12492 17110
rect 12552 17050 12558 17110
rect 12492 16530 12552 17050
rect 12490 16524 12552 16530
rect 12550 16464 12552 16524
rect 12490 16458 12552 16464
rect 12492 15404 12552 16458
rect 12714 16228 12720 16288
rect 12780 16228 12786 16288
rect 12492 14896 12552 15344
rect 12720 14912 12780 16228
rect 12838 15012 12898 18282
rect 14806 18236 15532 18296
rect 14746 18230 14806 18236
rect 15532 18230 15592 18236
rect 22484 18048 22544 18054
rect 24286 18048 24346 18054
rect 17636 18040 17696 18046
rect 19430 18040 19490 18046
rect 21466 18040 21526 18046
rect 17696 17980 19430 18040
rect 19490 17980 21466 18040
rect 22544 17988 24286 18048
rect 22484 17982 22544 17988
rect 24286 17982 24346 17988
rect 24520 18042 24580 18048
rect 26556 18042 26616 18048
rect 24580 17982 26556 18042
rect 17636 17974 17696 17980
rect 13286 17110 13346 17116
rect 15632 17052 15638 17112
rect 15698 17052 15704 17112
rect 13286 16524 13346 17050
rect 13386 16876 13392 16936
rect 13452 16876 13458 16936
rect 13280 16464 13286 16524
rect 13346 16464 13352 16524
rect 13160 16346 13166 16406
rect 13226 16346 13232 16406
rect 13166 15022 13226 16346
rect 13286 15430 13346 16464
rect 13269 15421 13359 15430
rect 13269 15322 13359 15331
rect 12832 14952 12838 15012
rect 12898 14952 12904 15012
rect 13286 15014 13346 15322
rect 13166 14956 13226 14962
rect 13280 14954 13286 15014
rect 13346 14954 13352 15014
rect 13392 14878 13452 16876
rect 15638 16522 15698 17052
rect 15638 16456 15698 16462
rect 12720 14846 12780 14852
rect 12492 14830 12552 14836
rect 13386 14818 13392 14878
rect 13452 14818 13458 14878
rect 12352 14812 12412 14818
rect 12610 14758 12670 14764
rect 17864 14758 17924 17980
rect 19430 17974 19490 17980
rect 21466 17974 21526 17980
rect 24520 17976 24580 17982
rect 26556 17976 26616 17982
rect 29610 18044 29670 18050
rect 31646 18044 31706 18050
rect 29670 17984 31646 18044
rect 29610 17978 29670 17984
rect 31646 17978 31706 17984
rect 21466 17932 21526 17938
rect 26554 17932 26614 17938
rect 33804 17932 33864 17938
rect 21526 17872 26554 17932
rect 26614 17872 33804 17932
rect 21466 17866 21526 17872
rect 26554 17866 26614 17872
rect 33804 17866 33864 17872
rect 18262 17832 18322 17838
rect 18322 17772 30846 17832
rect 18262 17766 18322 17772
rect 20444 17730 20504 17736
rect 22478 17730 22538 17736
rect 20504 17670 22478 17730
rect 30632 17730 30692 17736
rect 30786 17730 30846 17772
rect 32666 17730 32726 17736
rect 20444 17664 20504 17670
rect 22478 17664 22538 17670
rect 22682 17718 22742 17724
rect 22742 17658 26044 17718
rect 26104 17658 27060 17718
rect 27120 17658 30120 17718
rect 30180 17658 30186 17718
rect 30692 17670 32666 17730
rect 30632 17664 30692 17670
rect 32666 17664 32726 17670
rect 22682 17652 22742 17658
rect 17994 16782 18054 16788
rect 19426 16782 19486 16788
rect 21462 16782 21522 16788
rect 18054 16722 19426 16782
rect 19486 16722 21462 16782
rect 17994 16716 18054 16722
rect 19426 16716 19486 16722
rect 21462 16716 21522 16722
rect 29614 16782 29674 16788
rect 31650 16782 31710 16788
rect 29674 16722 31650 16782
rect 29614 16716 29674 16722
rect 18130 16652 18190 16658
rect 29744 16652 29804 16722
rect 31650 16716 31710 16722
rect 18190 16592 29804 16652
rect 18130 16586 18190 16592
rect 22484 16512 22544 16518
rect 34088 16512 34148 16518
rect 22544 16452 34088 16512
rect 22484 16446 22544 16452
rect 12670 14698 17924 14758
rect 12610 14692 12670 14698
rect 12100 14682 12160 14688
rect -3432 14300 -1262 14548
rect 24204 14528 24264 16452
rect 24204 14462 24264 14468
rect 29308 14528 29368 16452
rect 33368 14522 33428 16452
rect 34088 16446 34148 16452
rect 29308 14462 29368 14468
rect 33362 14462 33368 14522
rect 33428 14462 33434 14522
rect -3432 13782 -2276 14300
rect -1748 13782 -1262 14300
rect 9388 14150 9448 14156
rect 13166 14150 13226 14156
rect 9448 14090 13166 14150
rect 9388 14084 9448 14090
rect 13166 14084 13226 14090
rect 10914 14016 10974 14022
rect 12720 14016 12780 14022
rect 10974 13956 12720 14016
rect 10914 13950 10974 13956
rect 12720 13950 12780 13956
rect -3432 13306 -1262 13782
rect -3432 1924 -3342 13306
rect -2908 1924 -1262 13306
rect 12962 12792 13022 12798
rect 13022 12732 14536 12792
rect 14596 12732 14602 12792
rect 12962 12726 13022 12732
rect 15550 12576 15610 12582
rect 17590 12576 17650 12582
rect 19630 12576 19690 12582
rect 21660 12576 21720 12582
rect 23700 12576 23760 12582
rect 25732 12576 25792 12582
rect 27772 12576 27832 12582
rect 29808 12576 29868 12582
rect 31842 12576 31902 12582
rect 15610 12516 17590 12576
rect 17650 12516 19630 12576
rect 19690 12516 21660 12576
rect 21720 12516 23700 12576
rect 23760 12516 25732 12576
rect 25792 12516 27772 12576
rect 27832 12516 29808 12576
rect 29868 12516 31842 12576
rect 15550 12510 15610 12516
rect 17590 12510 17650 12516
rect 19630 12510 19690 12516
rect 21660 12510 21720 12516
rect 23700 12510 23760 12516
rect 25732 12510 25792 12516
rect 27772 12510 27832 12516
rect 29808 12510 29868 12516
rect 31842 12510 31902 12516
rect 13174 12456 13234 12462
rect 13518 12456 13578 12462
rect 13234 12396 13518 12456
rect 13174 12390 13234 12396
rect 13518 12390 13578 12396
rect 15042 12450 15102 12456
rect 23186 12450 23246 12456
rect 15102 12390 16056 12450
rect 16116 12390 17078 12450
rect 17138 12390 18092 12450
rect 18152 12390 19118 12450
rect 19178 12390 20130 12450
rect 20190 12390 21166 12450
rect 21226 12390 22172 12450
rect 22232 12390 23186 12450
rect 23246 12390 24202 12450
rect 24262 12390 25210 12450
rect 25270 12390 26226 12450
rect 26286 12390 27250 12450
rect 27310 12390 28272 12450
rect 28332 12390 29294 12450
rect 29354 12390 30312 12450
rect 30372 12390 31326 12450
rect 31386 12390 32350 12450
rect 32410 12390 32416 12450
rect 15042 12384 15102 12390
rect 23186 12384 23246 12390
rect 13392 12334 13452 12340
rect 18606 12334 18666 12340
rect 28794 12334 28854 12340
rect 32866 12334 32926 12340
rect 33998 12334 34058 12340
rect 13452 12274 18606 12334
rect 18666 12274 28794 12334
rect 28854 12274 32866 12334
rect 32926 12274 33998 12334
rect 13392 12268 13452 12274
rect 18606 12268 18666 12274
rect 28794 12268 28854 12274
rect 32866 12268 32926 12274
rect 33998 12268 34058 12274
rect 13286 12066 13346 12072
rect 12486 12006 12492 12066
rect 12552 12006 13286 12066
rect 13286 12000 13346 12006
rect 15554 11412 15614 11418
rect 17594 11412 17654 11418
rect 19626 11412 19686 11418
rect 21658 11412 21718 11418
rect 23694 11412 23754 11418
rect 25730 11412 25790 11418
rect 27768 11412 27828 11418
rect 29806 11412 29866 11418
rect 31842 11412 31902 11418
rect 15614 11352 17594 11412
rect 17654 11352 19626 11412
rect 19686 11352 21658 11412
rect 21718 11352 23694 11412
rect 23754 11352 25730 11412
rect 25790 11352 27768 11412
rect 27828 11352 29806 11412
rect 29866 11352 31842 11412
rect 15554 11346 15614 11352
rect 17594 11346 17654 11352
rect 19626 11346 19686 11352
rect 21658 11346 21718 11352
rect 23694 11346 23754 11352
rect 25730 11346 25790 11352
rect 27768 11346 27828 11352
rect 29806 11346 29866 11352
rect 31842 11346 31902 11352
rect 15046 11302 15106 11308
rect 16068 11302 16128 11308
rect 17082 11302 17142 11308
rect 18096 11302 18156 11308
rect 19114 11302 19174 11308
rect 20140 11302 20200 11308
rect 21160 11302 21220 11308
rect 22180 11302 22240 11308
rect 23182 11302 23242 11308
rect 24208 11302 24268 11308
rect 25226 11302 25286 11308
rect 26234 11302 26294 11308
rect 27246 11302 27306 11308
rect 28278 11302 28338 11308
rect 29292 11302 29352 11308
rect 30310 11302 30370 11308
rect 31334 11302 31394 11308
rect 32354 11302 32414 11308
rect 15106 11242 16068 11302
rect 16128 11242 17082 11302
rect 17142 11242 18096 11302
rect 18156 11242 19114 11302
rect 19174 11242 20140 11302
rect 20200 11242 21160 11302
rect 21220 11242 22180 11302
rect 22240 11242 23182 11302
rect 23242 11242 24208 11302
rect 24268 11242 25226 11302
rect 25286 11242 26234 11302
rect 26294 11242 27246 11302
rect 27306 11242 28278 11302
rect 28338 11242 29292 11302
rect 29352 11242 30310 11302
rect 30370 11242 31334 11302
rect 31394 11242 32354 11302
rect 15046 11236 15106 11242
rect 16068 11236 16128 11242
rect 17082 11236 17142 11242
rect 18096 11236 18156 11242
rect 19114 11236 19174 11242
rect 20140 11236 20200 11242
rect 21160 11236 21220 11242
rect 22180 11236 22240 11242
rect 23182 11236 23242 11242
rect 24208 11236 24268 11242
rect 25226 11236 25286 11242
rect 26234 11236 26294 11242
rect 27246 11236 27306 11242
rect 28278 11236 28338 11242
rect 29292 11236 29352 11242
rect 30310 11236 30370 11242
rect 31334 11236 31394 11242
rect 32354 11236 32414 11242
rect 13070 11196 13130 11202
rect 14536 11196 14596 11202
rect 16576 11196 16636 11202
rect 18606 11196 18666 11202
rect 20646 11196 20706 11202
rect 22680 11196 22740 11202
rect 24716 11196 24776 11202
rect 26752 11196 26812 11202
rect 28792 11196 28852 11202
rect 30822 11196 30882 11202
rect 32862 11196 32922 11202
rect 13130 11136 14536 11196
rect 14596 11136 16576 11196
rect 16636 11136 18606 11196
rect 18666 11136 20646 11196
rect 20706 11136 22680 11196
rect 22740 11136 24716 11196
rect 24776 11136 26752 11196
rect 26812 11136 28792 11196
rect 28852 11136 30822 11196
rect 30882 11136 32862 11196
rect 13070 11130 13130 11136
rect 14536 11130 14596 11136
rect 16576 11130 16636 11136
rect 18606 11130 18666 11136
rect 20646 11130 20706 11136
rect 22680 11130 22740 11136
rect 24716 11130 24776 11136
rect 26752 11130 26812 11136
rect 28792 11130 28852 11136
rect 30822 11130 30882 11136
rect 32862 11130 32922 11136
rect 13522 11090 13582 11096
rect 14020 11090 14080 11096
rect 14532 11090 14592 11096
rect 20812 11090 20872 11096
rect 22680 11090 22740 11096
rect 24718 11090 24778 11096
rect 26598 11090 26658 11096
rect 12830 11030 12836 11090
rect 12896 11030 13522 11090
rect 13582 11030 14020 11090
rect 14080 11030 14532 11090
rect 14592 11030 20812 11090
rect 20872 11030 22680 11090
rect 22740 11030 24718 11090
rect 24778 11030 26598 11090
rect 13522 11024 13582 11030
rect 14020 11024 14080 11030
rect 14532 11024 14592 11030
rect 20812 11024 20872 11030
rect 22680 11024 22740 11030
rect 24718 11024 24778 11030
rect 26598 11024 26658 11030
rect 30822 11092 30882 11098
rect 33998 11092 34058 11098
rect 30882 11032 33998 11092
rect 30822 11026 30882 11032
rect 33998 11026 34058 11032
rect 13392 10200 13452 10206
rect 16570 10200 16630 10206
rect 19626 10200 19686 10206
rect 25732 10200 25792 10206
rect 30826 10200 30886 10206
rect 13452 10140 16570 10200
rect 16630 10140 19626 10200
rect 19686 10140 25732 10200
rect 25792 10140 30826 10200
rect 13392 10134 13452 10140
rect 16570 10134 16630 10140
rect 19626 10134 19686 10140
rect 25732 10134 25792 10140
rect 30826 10134 30886 10140
rect 12962 10096 13022 10102
rect 13516 10096 13576 10102
rect 15036 10096 15096 10102
rect 13022 10036 13516 10096
rect 13576 10036 15036 10096
rect 12962 10030 13022 10036
rect 13516 10030 13576 10036
rect 15036 10030 15096 10036
rect 15548 10096 15608 10102
rect 16572 10096 16632 10102
rect 17584 10096 17644 10102
rect 18604 10096 18664 10102
rect 21662 10096 21722 10102
rect 23700 10096 23760 10102
rect 26750 10096 26810 10102
rect 27768 10096 27828 10102
rect 28788 10096 28848 10102
rect 29804 10096 29864 10102
rect 31840 10096 31900 10102
rect 15608 10036 16572 10096
rect 16632 10036 17584 10096
rect 17644 10036 18604 10096
rect 18664 10036 21662 10096
rect 21722 10036 23700 10096
rect 23760 10036 26750 10096
rect 26810 10036 27768 10096
rect 27828 10036 28788 10096
rect 28848 10036 29804 10096
rect 29864 10036 31840 10096
rect 15548 10030 15608 10036
rect 16572 10030 16632 10036
rect 17584 10030 17644 10036
rect 18604 10030 18664 10036
rect 21662 10030 21722 10036
rect 23700 10030 23760 10036
rect 26750 10030 26810 10036
rect 27768 10030 27828 10036
rect 28788 10030 28848 10036
rect 29804 10030 29864 10036
rect 31840 10030 31900 10036
rect 13286 9974 13346 9980
rect 20646 9974 20706 9980
rect 22680 9974 22740 9980
rect 24710 9974 24770 9980
rect 34710 9974 34770 18932
rect 12486 9914 12492 9974
rect 12552 9914 13286 9974
rect 13346 9914 20646 9974
rect 20706 9914 22680 9974
rect 22740 9914 24710 9974
rect 24770 9914 34708 9974
rect 34768 9914 34777 9974
rect 13286 9908 13346 9914
rect 20646 9908 20706 9914
rect 22680 9908 22740 9914
rect 24710 9908 24770 9914
rect 13174 9860 13234 9866
rect 14022 9860 14082 9866
rect 13234 9800 14022 9860
rect 13174 9794 13234 9800
rect 14022 9794 14082 9800
rect 15554 9862 15614 9868
rect 17590 9862 17650 9868
rect 33984 9862 34044 9868
rect 15614 9802 17590 9862
rect 17650 9802 33984 9862
rect 15554 9796 15614 9802
rect 17590 9796 17650 9802
rect 33984 9796 34044 9802
rect 34112 9844 34172 9850
rect 34712 9844 34772 9850
rect 34172 9784 34712 9844
rect 34112 9778 34172 9784
rect 34712 9778 34772 9784
rect 33878 8974 33938 8980
rect 34838 8974 34898 19250
rect 37958 15992 49228 16248
rect 37958 15700 38320 15992
rect 49172 15700 49228 15992
rect 37958 15392 49228 15700
rect 37958 15070 50310 15392
rect 53100 14748 53160 22100
rect 60632 22094 60692 22100
rect 64712 22094 64772 22100
rect 68780 22094 68840 22100
rect 72848 22094 72908 22100
rect 75240 22094 75300 22100
rect 58636 22028 58696 22034
rect 63178 22028 63184 22030
rect 58696 22026 63184 22028
rect 58696 21968 61138 22026
rect 58636 21962 58696 21968
rect 61132 21966 61138 21968
rect 61198 22022 63184 22026
rect 61198 21968 62152 22022
rect 61198 21966 61204 21968
rect 62146 21962 62152 21968
rect 62212 21970 63184 22022
rect 63244 22028 63250 22030
rect 64176 22028 64182 22030
rect 63244 21970 64182 22028
rect 64242 22028 64248 22030
rect 65220 22028 65226 22030
rect 64242 21970 65226 22028
rect 65286 22028 65292 22030
rect 69276 22028 69282 22030
rect 65286 22026 69282 22028
rect 65286 21970 66230 22026
rect 62212 21968 66230 21970
rect 62212 21962 62218 21968
rect 66224 21966 66230 21968
rect 66290 21968 67246 22026
rect 66290 21966 66296 21968
rect 67240 21966 67246 21968
rect 67306 21968 68250 22026
rect 67306 21966 67312 21968
rect 68244 21966 68250 21968
rect 68310 21970 69282 22026
rect 69342 22028 69348 22030
rect 74804 22028 74864 22034
rect 69342 22026 74804 22028
rect 69342 21970 70298 22026
rect 68310 21968 70298 21970
rect 68310 21966 68316 21968
rect 70292 21966 70298 21968
rect 70358 21968 71326 22026
rect 70358 21966 70364 21968
rect 71320 21966 71326 21968
rect 71386 21968 72346 22026
rect 71386 21966 71392 21968
rect 72340 21966 72346 21968
rect 72406 21968 74804 22026
rect 72406 21966 72412 21968
rect 74804 21962 74864 21968
rect 66030 21818 66090 21824
rect 66090 21758 67766 21818
rect 67826 21758 67832 21818
rect 73664 21804 73724 21808
rect 73662 21802 75006 21804
rect 66030 21752 66090 21758
rect 73662 21742 73664 21802
rect 73724 21800 75006 21802
rect 73724 21742 74946 21800
rect 73662 21740 74946 21742
rect 75006 21740 75012 21800
rect 73664 21736 73724 21740
rect 67046 21622 67110 21628
rect 71110 21622 71174 21628
rect 72134 21622 72198 21628
rect 73146 21622 73210 21628
rect 67110 21558 71110 21622
rect 71174 21558 72134 21622
rect 72198 21558 73146 21622
rect 67046 21552 67110 21558
rect 71110 21552 71174 21558
rect 72134 21552 72198 21558
rect 73146 21552 73210 21558
rect 59262 21500 59322 21506
rect 60428 21500 60488 21506
rect 62464 21500 62524 21506
rect 59322 21440 60428 21500
rect 60488 21440 62464 21500
rect 59262 21434 59322 21440
rect 60428 21434 60488 21440
rect 62464 21434 62524 21440
rect 62972 21500 63036 21506
rect 67048 21500 67112 21506
rect 63036 21436 67048 21500
rect 62972 21430 63036 21436
rect 67048 21430 67112 21436
rect 70610 21500 70670 21506
rect 72644 21500 72704 21506
rect 75088 21500 75148 21506
rect 70670 21440 72644 21500
rect 72704 21440 75088 21500
rect 70610 21434 70670 21440
rect 72644 21434 72704 21440
rect 75088 21434 75148 21440
rect 58510 21418 58570 21424
rect 58752 21418 58812 21424
rect 58570 21358 58752 21418
rect 58510 21352 58570 21358
rect 58752 21352 58812 21358
rect 61446 20552 61506 20558
rect 63482 20552 63542 20558
rect 61506 20492 63482 20552
rect 61446 20486 61506 20492
rect 63482 20486 63542 20492
rect 63824 20554 63884 20560
rect 66538 20554 66598 20560
rect 63884 20494 66538 20554
rect 63824 20488 63884 20494
rect 66538 20488 66598 20494
rect 71626 20552 71686 20558
rect 73662 20552 73722 20558
rect 71686 20492 73662 20552
rect 71626 20486 71686 20492
rect 55626 20464 55686 20470
rect 56648 20464 56708 20470
rect 55686 20404 56648 20464
rect 55626 20398 55686 20404
rect 56648 20398 56708 20404
rect 58994 20454 59054 20460
rect 71734 20454 71794 20492
rect 73662 20486 73722 20492
rect 59054 20394 71794 20454
rect 58994 20388 59054 20394
rect 55734 20352 55794 20358
rect 56518 20352 56578 20358
rect 55794 20292 56518 20352
rect 55734 20286 55794 20292
rect 56518 20286 56578 20292
rect 59130 20356 59190 20362
rect 61446 20356 61506 20362
rect 59190 20296 61446 20356
rect 59130 20290 59190 20296
rect 61446 20290 61506 20296
rect 62466 20358 62526 20364
rect 67556 20358 67616 20364
rect 74928 20358 74988 20364
rect 62526 20298 67556 20358
rect 67616 20298 74928 20358
rect 62466 20292 62526 20298
rect 67556 20292 67616 20298
rect 74928 20292 74988 20298
rect 60432 20246 60492 20252
rect 62466 20246 62526 20252
rect 60492 20186 62466 20246
rect 60432 20180 60492 20186
rect 62466 20180 62526 20186
rect 65522 20244 65582 20250
rect 67556 20244 67616 20250
rect 65582 20184 67556 20244
rect 65522 20178 65582 20184
rect 67556 20178 67616 20184
rect 70612 20244 70672 20250
rect 72646 20246 72706 20250
rect 72578 20244 72706 20246
rect 75240 20244 75300 20250
rect 70672 20184 72646 20244
rect 72706 20184 75240 20244
rect 70612 20178 70672 20184
rect 72578 20182 72706 20184
rect 72646 20178 72706 20182
rect 75240 20178 75300 20184
rect 53964 19430 54024 19436
rect 57158 19430 57218 19436
rect 54024 19370 57158 19430
rect 53964 19364 54024 19370
rect 57158 19364 57218 19370
rect 55124 19320 55184 19326
rect 58310 19320 58370 19326
rect 55184 19260 58310 19320
rect 71476 19310 71536 19316
rect 55124 19254 55184 19260
rect 58310 19254 58370 19260
rect 58752 19296 58812 19302
rect 65518 19296 65578 19302
rect 66538 19296 66598 19302
rect 68574 19296 68634 19302
rect 58812 19236 65518 19296
rect 65578 19236 66538 19296
rect 66598 19236 68574 19296
rect 71536 19250 75898 19310
rect 71476 19244 71536 19250
rect 58752 19230 58812 19236
rect 65518 19230 65578 19236
rect 66538 19230 66598 19236
rect 68574 19230 68634 19236
rect 71624 19200 71684 19206
rect 73664 19200 73724 19206
rect 74804 19200 74864 19206
rect 58502 19192 58562 19198
rect 63484 19192 63544 19198
rect 70608 19192 70668 19198
rect 58562 19132 61448 19192
rect 61508 19132 63484 19192
rect 63544 19132 70608 19192
rect 71684 19140 73664 19200
rect 73724 19140 74804 19200
rect 71624 19134 71684 19140
rect 73664 19134 73724 19140
rect 74804 19134 74864 19140
rect 58502 19126 58562 19132
rect 63484 19126 63544 19132
rect 70608 19126 70668 19132
rect 63482 19090 63542 19096
rect 72644 19090 72704 19096
rect 58748 19082 58808 19088
rect 59414 19082 59474 19088
rect 58808 19022 59414 19082
rect 63542 19030 72644 19090
rect 63482 19024 63542 19030
rect 72644 19024 72704 19030
rect 58748 19016 58808 19022
rect 59414 19016 59474 19022
rect 61448 18988 61508 18994
rect 63482 18988 63542 18994
rect 61508 18928 63482 18988
rect 61448 18922 61508 18928
rect 63482 18922 63542 18928
rect 66538 18990 66598 18996
rect 67556 18990 67616 18996
rect 68572 18990 68632 18996
rect 71476 18990 71536 18996
rect 66598 18930 67556 18990
rect 67616 18930 68572 18990
rect 68632 18930 71476 18990
rect 66538 18924 66598 18930
rect 67556 18924 67616 18930
rect 68572 18924 68632 18930
rect 71476 18924 71536 18930
rect 71628 18992 71688 18998
rect 73662 18992 73722 18998
rect 74928 18992 74988 18998
rect 71688 18932 73662 18992
rect 73722 18932 74928 18992
rect 74988 18932 75770 18992
rect 71628 18926 71688 18932
rect 73662 18926 73722 18932
rect 74928 18926 74988 18932
rect 55640 18396 55700 18402
rect 56650 18396 56710 18402
rect 53832 18282 53838 18342
rect 53898 18282 53904 18342
rect 55700 18336 56650 18396
rect 55640 18330 55700 18336
rect 56650 18330 56710 18336
rect 55746 18296 55806 18302
rect 56532 18296 56592 18302
rect 53346 17226 53352 17286
rect 53412 17226 53418 17286
rect 53226 16726 53232 16786
rect 53292 16726 53298 16786
rect 53232 14876 53292 16726
rect 53232 14810 53292 14816
rect 53352 14878 53412 17226
rect 53486 17050 53492 17110
rect 53552 17050 53558 17110
rect 53492 14896 53552 17050
rect 53714 16228 53720 16288
rect 53780 16228 53786 16288
rect 53720 14912 53780 16228
rect 53838 15012 53898 18282
rect 55806 18236 56532 18296
rect 55746 18230 55806 18236
rect 56532 18230 56592 18236
rect 63484 18048 63544 18054
rect 65286 18048 65346 18054
rect 58636 18040 58696 18046
rect 60430 18040 60490 18046
rect 62466 18040 62526 18046
rect 58696 17980 60430 18040
rect 60490 17980 62466 18040
rect 63544 17988 65286 18048
rect 63484 17982 63544 17988
rect 65286 17982 65346 17988
rect 65520 18042 65580 18048
rect 67556 18042 67616 18048
rect 65580 17982 67556 18042
rect 58636 17974 58696 17980
rect 54386 16876 54392 16936
rect 54452 16876 54458 16936
rect 54280 16464 54286 16524
rect 54346 16464 54352 16524
rect 54160 16346 54166 16406
rect 54226 16346 54232 16406
rect 54166 15022 54226 16346
rect 54286 15430 54346 16464
rect 54269 15421 54359 15430
rect 54269 15322 54359 15331
rect 53832 14952 53838 15012
rect 53898 14952 53904 15012
rect 54286 15014 54346 15322
rect 54166 14956 54226 14962
rect 54280 14954 54286 15014
rect 54346 14954 54352 15014
rect 54392 14878 54452 16876
rect 53720 14846 53780 14852
rect 53492 14830 53552 14836
rect 54386 14818 54392 14878
rect 54452 14818 54458 14878
rect 53352 14812 53412 14818
rect 53610 14758 53670 14764
rect 58864 14758 58924 17980
rect 60430 17974 60490 17980
rect 62466 17974 62526 17980
rect 65520 17976 65580 17982
rect 67556 17976 67616 17982
rect 70610 18044 70670 18050
rect 72646 18044 72706 18050
rect 70670 17984 72646 18044
rect 70610 17978 70670 17984
rect 72646 17978 72706 17984
rect 62466 17932 62526 17938
rect 67554 17932 67614 17938
rect 74804 17932 74864 17938
rect 62526 17872 67554 17932
rect 67614 17872 74804 17932
rect 62466 17866 62526 17872
rect 67554 17866 67614 17872
rect 74804 17866 74864 17872
rect 59262 17832 59322 17838
rect 59322 17772 71846 17832
rect 59262 17766 59322 17772
rect 61444 17730 61504 17736
rect 63478 17730 63538 17736
rect 61504 17670 63478 17730
rect 71632 17730 71692 17736
rect 71786 17730 71846 17772
rect 73666 17730 73726 17736
rect 61444 17664 61504 17670
rect 63478 17664 63538 17670
rect 63682 17718 63742 17724
rect 63742 17658 67044 17718
rect 67104 17658 68060 17718
rect 68120 17658 71120 17718
rect 71180 17658 71186 17718
rect 71692 17670 73666 17730
rect 71632 17664 71692 17670
rect 73666 17664 73726 17670
rect 63682 17652 63742 17658
rect 58994 16782 59054 16788
rect 60426 16782 60486 16788
rect 62462 16782 62522 16788
rect 59054 16722 60426 16782
rect 60486 16722 62462 16782
rect 58994 16716 59054 16722
rect 60426 16716 60486 16722
rect 62462 16716 62522 16722
rect 70614 16782 70674 16788
rect 72650 16782 72710 16788
rect 70674 16722 72650 16782
rect 70614 16716 70674 16722
rect 59130 16652 59190 16658
rect 70744 16652 70804 16722
rect 72650 16716 72710 16722
rect 59190 16592 70804 16652
rect 59130 16586 59190 16592
rect 63484 16512 63544 16518
rect 75088 16512 75148 16518
rect 63544 16452 75088 16512
rect 63484 16446 63544 16452
rect 53670 14698 58924 14758
rect 53610 14692 53670 14698
rect 53100 14682 53160 14688
rect 65204 14528 65264 16452
rect 65204 14462 65264 14468
rect 70308 14528 70368 16452
rect 74368 14522 74428 16452
rect 75088 16446 75148 16452
rect 70308 14462 70368 14468
rect 74362 14462 74368 14522
rect 74428 14462 74434 14522
rect 50388 14150 50448 14156
rect 54166 14150 54226 14156
rect 50448 14090 54166 14150
rect 50388 14084 50448 14090
rect 54166 14084 54226 14090
rect 51914 14016 51974 14022
rect 53720 14016 53780 14022
rect 51974 13956 53720 14016
rect 51914 13950 51974 13956
rect 53720 13950 53780 13956
rect 36824 13864 37424 13874
rect 36824 13554 37424 13564
rect 37976 13864 38576 13874
rect 37976 13554 38576 13564
rect 36890 13396 38514 13426
rect 36890 13300 36928 13396
rect 38480 13300 38514 13396
rect 36890 13272 38514 13300
rect 37672 13194 37732 13200
rect 39132 13194 39192 13203
rect 37732 13134 39132 13194
rect 37672 13128 37732 13134
rect 39132 13125 39192 13134
rect 53962 12792 54022 12798
rect 54022 12732 55536 12792
rect 55596 12732 55602 12792
rect 53962 12726 54022 12732
rect 16570 8956 16630 8962
rect 18606 8956 18666 8962
rect 26750 8956 26810 8962
rect 28786 8956 28846 8962
rect 32860 8956 32920 8962
rect 13398 8932 13458 8938
rect 14536 8932 14596 8938
rect 13458 8872 14536 8932
rect 14596 8872 15418 8932
rect 16630 8896 18606 8956
rect 18666 8896 26750 8956
rect 26810 8896 28786 8956
rect 28846 8896 32860 8956
rect 33938 8914 34898 8974
rect 37136 12660 37236 12678
rect 38186 12660 38246 12666
rect 37136 12600 37156 12660
rect 37216 12600 38186 12660
rect 33878 8908 33938 8914
rect 16570 8890 16630 8896
rect 18606 8890 18666 8896
rect 26750 8890 26810 8896
rect 28786 8890 28846 8896
rect 32860 8890 32920 8896
rect 13398 8866 13458 8872
rect 14536 8866 14596 8872
rect 13286 8732 13346 8738
rect 14534 8732 14594 8738
rect 12486 8672 12492 8732
rect 12552 8672 13286 8732
rect 13346 8672 14534 8732
rect 15358 8736 15418 8872
rect 15552 8852 15612 8858
rect 17592 8852 17652 8858
rect 19624 8852 19684 8858
rect 21658 8852 21718 8858
rect 23698 8852 23758 8858
rect 25732 8852 25792 8858
rect 15612 8792 17592 8852
rect 17652 8792 19624 8852
rect 19684 8792 21658 8852
rect 21718 8792 23698 8852
rect 23758 8792 25732 8852
rect 15552 8786 15612 8792
rect 17592 8786 17652 8792
rect 19624 8786 19684 8792
rect 21658 8786 21718 8792
rect 23698 8786 23758 8792
rect 25732 8786 25792 8792
rect 25928 8848 25988 8854
rect 30820 8848 30880 8854
rect 25988 8788 30820 8848
rect 34478 8844 34538 8850
rect 25928 8782 25988 8788
rect 30820 8782 30880 8788
rect 31318 8784 31324 8844
rect 31384 8784 34478 8844
rect 34478 8778 34538 8784
rect 16066 8738 16126 8744
rect 19624 8740 19684 8746
rect 21660 8740 21720 8746
rect 23696 8740 23756 8746
rect 25732 8740 25792 8746
rect 27766 8740 27826 8746
rect 29804 8740 29864 8746
rect 31844 8740 31904 8746
rect 34228 8740 34288 8746
rect 15358 8678 16066 8736
rect 16126 8678 17070 8738
rect 17130 8678 18082 8738
rect 18142 8678 19102 8738
rect 19162 8678 19168 8738
rect 19684 8680 21660 8740
rect 21720 8680 23696 8740
rect 23756 8680 25732 8740
rect 25792 8680 27766 8740
rect 27826 8680 29804 8740
rect 29864 8680 31844 8740
rect 31904 8680 34228 8740
rect 15358 8676 16408 8678
rect 16066 8672 16126 8676
rect 19624 8674 19684 8680
rect 21660 8674 21720 8680
rect 23696 8674 23756 8680
rect 25732 8674 25792 8680
rect 27766 8674 27826 8680
rect 29804 8674 29864 8680
rect 31844 8674 31904 8680
rect 34228 8674 34288 8680
rect 13286 8666 13346 8672
rect 14534 8666 14594 8672
rect 12610 8630 12670 8636
rect 13180 8630 13240 8636
rect 20642 8630 20702 8636
rect 22676 8630 22736 8636
rect 24716 8630 24776 8636
rect 25928 8630 25988 8636
rect 12670 8570 13180 8630
rect 13240 8570 20642 8630
rect 20702 8570 22676 8630
rect 22736 8570 24716 8630
rect 24776 8570 25928 8630
rect 12610 8564 12670 8570
rect 13180 8564 13240 8570
rect 20642 8564 20702 8570
rect 22676 8564 22736 8570
rect 24716 8564 24776 8570
rect 25928 8564 25988 8570
rect 26222 8632 26282 8638
rect 26282 8572 27250 8632
rect 27310 8572 27316 8632
rect 27768 8626 27828 8632
rect 29804 8626 29864 8632
rect 31842 8626 31902 8632
rect 33984 8626 34044 8632
rect 26222 8566 26282 8572
rect 27828 8566 29804 8626
rect 29864 8566 31842 8626
rect 31902 8566 33984 8626
rect 27768 8560 27828 8566
rect 29804 8560 29864 8566
rect 31842 8560 31902 8566
rect 33984 8560 34044 8566
rect 30316 7712 30376 7718
rect 14534 7700 14594 7706
rect 16572 7700 16632 7706
rect 18608 7700 18668 7706
rect 20640 7700 20700 7706
rect 14594 7640 16572 7700
rect 16632 7640 18608 7700
rect 18668 7640 20640 7700
rect 25216 7652 25222 7712
rect 25282 7652 30316 7712
rect 30316 7646 30376 7652
rect 30454 7716 30514 7722
rect 31336 7716 31396 7722
rect 32342 7716 32402 7722
rect 30514 7656 31336 7716
rect 31396 7656 32342 7716
rect 30454 7650 30514 7656
rect 31336 7650 31396 7656
rect 32342 7650 32402 7656
rect 32860 7712 32920 7718
rect 34112 7712 34172 7718
rect 32920 7652 34112 7712
rect 32860 7646 32920 7652
rect 34112 7646 34172 7652
rect 14534 7634 14594 7640
rect 16572 7634 16632 7640
rect 18608 7634 18668 7640
rect 20640 7634 20700 7640
rect 15040 7598 15100 7604
rect 20132 7598 20192 7604
rect 12100 7548 12160 7554
rect 15100 7538 20132 7598
rect 15040 7532 15100 7538
rect 20132 7532 20192 7538
rect 24716 7584 24776 7590
rect 32860 7584 32920 7590
rect 24776 7524 32860 7584
rect 24716 7518 24776 7524
rect 32860 7518 32920 7524
rect 13286 7496 13346 7502
rect 16570 7496 16630 7502
rect 7552 6622 7612 6628
rect 12100 6622 12160 7488
rect 12486 7436 12492 7496
rect 12552 7436 13286 7496
rect 13346 7436 16570 7496
rect 13286 7430 13346 7436
rect 16570 7430 16630 7436
rect 17078 7490 17138 7496
rect 18100 7490 18160 7496
rect 19114 7490 19174 7496
rect 20132 7490 20192 7496
rect 21152 7490 21212 7496
rect 28264 7490 28324 7496
rect 29294 7490 29354 7496
rect 30454 7490 30514 7496
rect 17138 7430 18100 7490
rect 18160 7430 19114 7490
rect 19174 7430 20132 7490
rect 20192 7430 21152 7490
rect 21212 7430 28264 7490
rect 28324 7430 29294 7490
rect 29354 7430 30454 7490
rect 17078 7424 17138 7430
rect 18100 7424 18160 7430
rect 19114 7424 19174 7430
rect 20132 7424 20192 7430
rect 21152 7424 21212 7430
rect 28264 7424 28324 7430
rect 29294 7424 29354 7430
rect 30454 7424 30514 7430
rect 30822 7490 30882 7496
rect 34350 7490 34410 7496
rect 30882 7430 34350 7490
rect 30822 7424 30882 7430
rect 34350 7424 34410 7430
rect 15554 7396 15614 7402
rect 17588 7396 17648 7402
rect 19624 7396 19684 7402
rect 15614 7336 17588 7396
rect 17648 7336 19624 7396
rect 15554 7330 15614 7336
rect 17588 7330 17648 7336
rect 19624 7330 19684 7336
rect 26752 7386 26812 7392
rect 30822 7386 30882 7392
rect 26812 7326 30822 7386
rect 26752 7320 26812 7326
rect 30822 7320 30882 7326
rect 31838 7388 31898 7394
rect 34228 7388 34288 7394
rect 31898 7328 34228 7388
rect 31838 7322 31898 7328
rect 34228 7322 34288 7328
rect 12492 6970 12552 6976
rect 12552 6910 13290 6970
rect 13350 6910 13356 6970
rect 12492 6904 12552 6910
rect 7612 6562 12160 6622
rect 7552 6556 7612 6562
rect 5522 6476 5582 6482
rect 9582 6476 9642 6482
rect 11766 6476 11826 6482
rect 12232 6476 12292 6482
rect 21660 6478 21720 6484
rect 23696 6478 23756 6484
rect 25732 6478 25792 6484
rect 27770 6478 27830 6484
rect 1436 6416 1442 6476
rect 1502 6416 5522 6476
rect 5582 6416 9582 6476
rect 9642 6416 11766 6476
rect 11826 6416 12232 6476
rect 5522 6410 5582 6416
rect 9582 6410 9642 6416
rect 11766 6410 11826 6416
rect 12232 6410 12292 6416
rect 15036 6472 15096 6478
rect 15946 6472 16006 6478
rect 16948 6472 17008 6478
rect 18100 6472 18160 6478
rect 19110 6472 19170 6478
rect 20116 6472 20176 6478
rect 21160 6472 21220 6478
rect 15096 6412 15946 6472
rect 16006 6412 16948 6472
rect 17008 6412 18100 6472
rect 18160 6412 19110 6472
rect 19170 6412 20116 6472
rect 20176 6412 21160 6472
rect 21720 6418 23696 6478
rect 23756 6418 25732 6478
rect 25792 6418 27770 6478
rect 21660 6412 21720 6418
rect 23696 6412 23756 6418
rect 25732 6412 25792 6418
rect 27770 6412 27830 6418
rect 29806 6478 29866 6484
rect 31844 6478 31904 6484
rect 29866 6418 31844 6478
rect 29806 6412 29866 6418
rect 31844 6412 31904 6418
rect 15036 6406 15096 6412
rect 15946 6406 16006 6412
rect 16948 6406 17008 6412
rect 18100 6406 18160 6412
rect 19110 6406 19170 6412
rect 20116 6406 20176 6412
rect 21160 6406 21220 6412
rect 17588 6370 17648 6376
rect 27762 6370 27822 6376
rect 29802 6370 29862 6376
rect 31840 6370 31900 6376
rect 288 6348 348 6354
rect 2966 6348 3026 6354
rect 3998 6348 4058 6354
rect 7058 6348 7118 6354
rect 8054 6348 8114 6354
rect 12352 6348 12412 6354
rect 348 6288 2966 6348
rect 3026 6288 3998 6348
rect 4058 6288 7058 6348
rect 7118 6288 8054 6348
rect 8114 6288 12352 6348
rect 17648 6310 27762 6370
rect 27822 6310 29802 6370
rect 29862 6310 31840 6370
rect 17588 6304 17648 6310
rect 27762 6304 27822 6310
rect 29802 6304 29862 6310
rect 31840 6304 31900 6310
rect 288 6282 348 6288
rect 2966 6282 3026 6288
rect 3998 6282 4058 6288
rect 7058 6282 7118 6288
rect 8054 6282 8114 6288
rect 12352 6282 12412 6288
rect 15036 6256 15096 6262
rect 17088 6256 17148 6262
rect 20114 6256 20174 6262
rect 21154 6256 21214 6262
rect 22168 6256 22228 6262
rect 23176 6256 23236 6262
rect 24220 6256 24280 6262
rect 25210 6256 25270 6262
rect 26228 6256 26288 6262
rect 27262 6256 27322 6262
rect 30294 6256 30354 6262
rect 31332 6256 31392 6262
rect 32358 6256 32418 6262
rect 15096 6196 16074 6256
rect 16134 6196 17088 6256
rect 17148 6196 20114 6256
rect 20174 6196 21154 6256
rect 21214 6196 22168 6256
rect 22228 6196 23176 6256
rect 23236 6196 24220 6256
rect 24280 6196 25210 6256
rect 25270 6196 26228 6256
rect 26288 6196 27262 6256
rect 27322 6196 30294 6256
rect 30354 6196 31332 6256
rect 31392 6196 32358 6256
rect 32418 6196 34476 6256
rect 34536 6196 34542 6256
rect 15036 6190 15096 6196
rect 17088 6190 17148 6196
rect 20114 6190 20174 6196
rect 21154 6190 21214 6196
rect 22168 6190 22228 6196
rect 23176 6190 23236 6196
rect 24220 6190 24280 6196
rect 25210 6190 25270 6196
rect 26228 6190 26288 6196
rect 27262 6190 27322 6196
rect 30294 6190 30354 6196
rect 31332 6190 31392 6196
rect 32358 6190 32418 6196
rect 20638 6152 20698 6158
rect 22680 6152 22740 6158
rect 24718 6152 24778 6158
rect 26752 6152 26812 6158
rect 28786 6154 28846 6160
rect 30820 6154 30880 6160
rect 32862 6154 32922 6160
rect 34112 6154 34172 6160
rect 13394 6092 13400 6152
rect 13460 6092 20638 6152
rect 20698 6092 22680 6152
rect 22740 6092 24718 6152
rect 24778 6092 26752 6152
rect 20638 6086 20698 6092
rect 22680 6086 22740 6092
rect 24718 6086 24778 6092
rect 26752 6086 26812 6092
rect 27264 6148 27324 6154
rect 28286 6148 28346 6154
rect 27324 6088 28286 6148
rect 28846 6094 30820 6154
rect 30880 6094 32862 6154
rect 32922 6094 34112 6154
rect 28786 6088 28846 6094
rect 30820 6088 30880 6094
rect 32862 6088 32922 6094
rect 34112 6088 34172 6094
rect 27264 6082 27324 6088
rect 28286 6082 28346 6088
rect 1946 5386 2006 5392
rect 2970 5386 3030 5392
rect 4002 5386 4062 5392
rect 5002 5386 5062 5392
rect 6022 5386 6082 5392
rect 7042 5386 7102 5392
rect 9066 5386 9126 5392
rect 11886 5386 11946 5392
rect 12492 5386 12552 5392
rect 13288 5386 13348 5392
rect 2006 5326 2970 5386
rect 3030 5326 4002 5386
rect 4062 5326 5002 5386
rect 5062 5326 6022 5386
rect 6082 5326 7042 5386
rect 7102 5326 8052 5386
rect 8112 5326 9066 5386
rect 9126 5326 10084 5386
rect 10144 5326 11886 5386
rect 11946 5326 12492 5386
rect 12552 5326 13288 5386
rect 1946 5320 2006 5326
rect 2970 5320 3030 5326
rect 4002 5320 4062 5326
rect 5002 5320 5062 5326
rect 6022 5320 6082 5326
rect 7042 5320 7102 5326
rect 9066 5320 9126 5326
rect 11886 5320 11946 5326
rect 12492 5320 12552 5326
rect 13288 5320 13348 5326
rect 1446 5282 1506 5288
rect 3482 5282 3542 5288
rect 5518 5282 5578 5288
rect 7552 5282 7612 5288
rect 9588 5282 9648 5288
rect 1506 5222 3482 5282
rect 3542 5222 5518 5282
rect 5578 5222 7552 5282
rect 7612 5222 9588 5282
rect 19628 5250 19688 5256
rect 23696 5250 23756 5256
rect 25730 5250 25790 5256
rect 1446 5216 1506 5222
rect 3482 5216 3542 5222
rect 5518 5216 5578 5222
rect 7552 5216 7612 5222
rect 9588 5216 9648 5222
rect 15034 5244 15094 5250
rect 16042 5244 16102 5250
rect 17056 5244 17116 5250
rect 18094 5244 18154 5250
rect 19112 5244 19172 5250
rect 15094 5184 16042 5244
rect 16102 5184 17056 5244
rect 17116 5184 18094 5244
rect 18154 5184 19112 5244
rect 19688 5190 21664 5250
rect 21724 5190 23696 5250
rect 23756 5190 25730 5250
rect 19628 5184 19688 5190
rect 23696 5184 23756 5190
rect 25730 5184 25790 5190
rect 26752 5252 26812 5258
rect 27106 5252 27166 5258
rect 26812 5192 27106 5252
rect 26752 5186 26812 5192
rect 27106 5186 27166 5192
rect 30824 5252 30884 5258
rect 34108 5252 34168 5258
rect 30884 5192 34108 5252
rect 34170 5192 34179 5252
rect 30824 5186 30884 5192
rect 34108 5186 34168 5192
rect 6532 5178 6592 5184
rect 13070 5178 13130 5184
rect 15034 5178 15094 5184
rect 16042 5178 16102 5184
rect 17056 5178 17116 5184
rect 18094 5178 18154 5184
rect 19112 5178 19172 5184
rect 2458 5118 2464 5178
rect 2524 5118 4500 5178
rect 4560 5118 6532 5178
rect 6592 5118 8566 5178
rect 8626 5118 10610 5178
rect 10670 5118 13070 5178
rect 6532 5112 6592 5118
rect 13070 5112 13130 5118
rect 13180 5140 13240 5146
rect 14536 5140 14596 5146
rect 22680 5140 22740 5146
rect 24716 5140 24776 5146
rect 26748 5140 26808 5146
rect 13240 5080 14536 5140
rect 14596 5080 22680 5140
rect 22740 5080 24716 5140
rect 24776 5080 26748 5140
rect 13180 5074 13240 5080
rect 14536 5074 14596 5080
rect 22680 5074 22740 5080
rect 24716 5074 24776 5080
rect 26748 5074 26808 5080
rect 26258 5042 26318 5048
rect 27296 5042 27356 5048
rect 28272 5042 28332 5048
rect 29288 5042 29348 5048
rect 31314 5042 31374 5048
rect 32344 5042 32404 5048
rect 12838 5028 12898 5034
rect 15552 5028 15612 5034
rect 17590 5028 17650 5034
rect 21662 5028 21722 5034
rect 12898 4968 15552 5028
rect 15612 4968 17590 5028
rect 17650 4968 21662 5028
rect 26318 4982 27296 5042
rect 27356 4982 28272 5042
rect 28332 4982 29288 5042
rect 29348 4982 31314 5042
rect 31374 4982 32344 5042
rect 26258 4976 26318 4982
rect 27296 4976 27356 4982
rect 28272 4976 28332 4982
rect 29288 4976 29348 4982
rect 31314 4976 31374 4982
rect 32344 4976 32404 4982
rect 12838 4962 12898 4968
rect 15552 4962 15612 4968
rect 17590 4962 17650 4968
rect 21662 4962 21722 4968
rect 14532 4930 14592 4936
rect 16570 4930 16630 4936
rect 18610 4930 18670 4936
rect 20646 4930 20706 4936
rect 26750 4930 26810 4936
rect 27100 4930 27106 4934
rect 14592 4870 16570 4930
rect 16630 4870 18610 4930
rect 18670 4870 20646 4930
rect 20706 4874 27106 4930
rect 27166 4930 27172 4934
rect 28786 4930 28846 4936
rect 30822 4930 30882 4936
rect 32858 4930 32918 4936
rect 27166 4874 28786 4930
rect 20706 4870 28786 4874
rect 28846 4870 30822 4930
rect 30882 4870 32858 4930
rect 14532 4864 14592 4870
rect 16570 4864 16630 4870
rect 18610 4864 18670 4870
rect 20646 4864 20706 4870
rect 26750 4864 26810 4870
rect 28786 4864 28846 4870
rect 30822 4864 30882 4870
rect 32858 4864 32918 4870
rect 11888 4730 11948 4736
rect 13286 4730 13346 4736
rect 11948 4670 13286 4730
rect 11888 4664 11948 4670
rect 13286 4664 13346 4670
rect 3476 4236 3536 4242
rect 7552 4236 7612 4242
rect 11766 4236 11826 4242
rect 3536 4176 7552 4236
rect 7612 4176 11766 4236
rect 3476 4170 3536 4176
rect 7552 4170 7612 4176
rect 11766 4170 11826 4176
rect 288 4116 348 4122
rect 1938 4116 1998 4122
rect 5008 4116 5068 4122
rect 6016 4116 6076 4122
rect 9078 4116 9138 4122
rect 10104 4116 10164 4122
rect 348 4056 1938 4116
rect 1998 4056 5008 4116
rect 5068 4056 6016 4116
rect 6076 4056 9078 4116
rect 9138 4056 10104 4116
rect 288 4050 348 4056
rect 1938 4050 1998 4056
rect 5008 4050 5068 4056
rect 6016 4050 6076 4056
rect 9078 4050 9138 4056
rect 10104 4050 10164 4056
rect 21658 4026 21718 4032
rect 23700 4026 23760 4032
rect 25732 4026 25792 4032
rect 27772 4026 27832 4032
rect 34228 4026 34288 4032
rect 15552 4006 15612 4012
rect 17588 4006 17648 4012
rect 19626 4006 19686 4012
rect 15612 3946 17588 4006
rect 17648 3946 19626 4006
rect 21482 3966 21488 4026
rect 21548 3966 21658 4026
rect 21718 3966 23700 4026
rect 23760 3966 25732 4026
rect 25792 3966 27772 4026
rect 27832 3966 34228 4026
rect 21658 3960 21718 3966
rect 23700 3960 23760 3966
rect 25732 3960 25792 3966
rect 27772 3960 27832 3966
rect 34228 3960 34288 3966
rect 15552 3940 15612 3946
rect 17588 3940 17648 3946
rect 19626 3940 19686 3946
rect 26750 3928 26810 3934
rect 32856 3928 32916 3934
rect 34108 3928 34168 3934
rect 13398 3908 13458 3914
rect 16570 3908 16630 3914
rect 13458 3848 16570 3908
rect 13398 3842 13458 3848
rect 16570 3842 16630 3848
rect 18094 3908 18154 3914
rect 21142 3908 21202 3914
rect 18154 3848 19116 3908
rect 19176 3848 20138 3908
rect 20198 3848 21142 3908
rect 26810 3868 32856 3928
rect 32916 3868 34108 3928
rect 26750 3862 26810 3868
rect 32856 3862 32916 3868
rect 34108 3862 34168 3868
rect 18094 3842 18154 3848
rect 21142 3842 21202 3848
rect 21664 3818 21724 3824
rect 23692 3818 23752 3824
rect 25736 3818 25796 3824
rect 27764 3818 27824 3824
rect 29802 3818 29862 3824
rect 31842 3818 31902 3824
rect 15556 3812 15616 3818
rect 17592 3812 17652 3818
rect 19620 3812 19680 3818
rect 21488 3812 21548 3818
rect 15616 3752 17592 3812
rect 17652 3752 19620 3812
rect 19680 3752 21488 3812
rect 21724 3758 23692 3818
rect 23752 3758 25736 3818
rect 25796 3758 27764 3818
rect 27824 3758 29802 3818
rect 29862 3758 31842 3818
rect 21664 3752 21724 3758
rect 23692 3752 23752 3758
rect 25736 3752 25796 3758
rect 27764 3752 27824 3758
rect 29802 3752 29862 3758
rect 31842 3752 31902 3758
rect 32360 3822 32420 3828
rect 33872 3822 33932 3828
rect 34478 3822 34538 3828
rect 32420 3762 33872 3822
rect 33932 3762 34478 3822
rect 32360 3756 32420 3762
rect 33872 3756 33932 3762
rect 34478 3756 34538 3762
rect 15556 3746 15616 3752
rect 17592 3746 17652 3752
rect 19620 3746 19680 3752
rect 21488 3746 21548 3752
rect 14538 3692 14598 3698
rect 18606 3692 18666 3698
rect 20640 3692 20700 3698
rect 28790 3692 28850 3698
rect 30820 3692 30880 3698
rect 32860 3694 32920 3700
rect 34350 3694 34410 3700
rect 14598 3632 18606 3692
rect 18666 3632 20640 3692
rect 20700 3632 28790 3692
rect 28850 3632 30820 3692
rect 31340 3634 31346 3694
rect 31406 3634 32860 3694
rect 32920 3634 34350 3694
rect 14538 3626 14598 3632
rect 18606 3626 18666 3632
rect 20640 3626 20700 3632
rect 28790 3626 28850 3632
rect 30820 3626 30880 3632
rect 32860 3628 32920 3634
rect 34350 3628 34410 3634
rect 10610 3172 10670 3178
rect 2458 3112 2464 3172
rect 2524 3112 4500 3172
rect 4560 3112 6532 3172
rect 6592 3112 8566 3172
rect 8626 3112 10610 3172
rect 10610 3106 10670 3112
rect 1450 3064 1510 3070
rect 3486 3064 3546 3070
rect 5522 3064 5582 3070
rect 7556 3064 7616 3070
rect 9592 3064 9652 3070
rect 1510 3004 3486 3064
rect 3546 3004 5522 3064
rect 5582 3004 7556 3064
rect 7616 3004 9592 3064
rect 1450 2998 1510 3004
rect 3486 2998 3546 3004
rect 5522 2998 5582 3004
rect 7556 2998 7616 3004
rect 9592 2998 9652 3004
rect 1944 2952 2004 2958
rect 2968 2952 3028 2958
rect 4000 2952 4060 2958
rect 5000 2952 5060 2958
rect 6020 2952 6080 2958
rect 7040 2952 7100 2958
rect 9064 2952 9124 2958
rect 11886 2952 11946 2958
rect 2004 2892 2968 2952
rect 3028 2892 4000 2952
rect 4060 2892 5000 2952
rect 5060 2892 6020 2952
rect 6080 2892 7040 2952
rect 7100 2892 8050 2952
rect 8110 2892 9064 2952
rect 9124 2892 10082 2952
rect 10142 2892 11886 2952
rect 1944 2886 2004 2892
rect 2968 2886 3028 2892
rect 4000 2886 4060 2892
rect 5000 2886 5060 2892
rect 6020 2886 6080 2892
rect 7040 2886 7100 2892
rect 9064 2886 9124 2892
rect 11886 2776 11946 2892
rect 13286 2776 13346 2782
rect 22674 2776 22734 2782
rect 24716 2776 24776 2782
rect 26752 2776 26812 2782
rect 11886 2716 13286 2776
rect 13346 2716 22674 2776
rect 22734 2716 24716 2776
rect 24776 2716 26752 2776
rect 13286 2710 13346 2716
rect 22674 2710 22734 2716
rect 24716 2710 24776 2716
rect 26752 2710 26812 2716
rect 29806 2776 29866 2782
rect 31838 2776 31898 2782
rect 33984 2776 34044 2782
rect 29866 2716 31838 2776
rect 31898 2716 33984 2776
rect 29806 2710 29866 2716
rect 31838 2710 31898 2716
rect 33984 2710 34044 2716
rect 17090 2662 17150 2668
rect 22170 2662 22230 2668
rect 13180 2650 13240 2656
rect 16570 2650 16630 2656
rect 13240 2590 16570 2650
rect 17150 2602 22170 2662
rect 17090 2596 17150 2602
rect 22170 2596 22230 2602
rect 27258 2666 27318 2672
rect 32358 2666 32418 2672
rect 27318 2606 32358 2666
rect 27258 2600 27318 2606
rect 32358 2600 32418 2606
rect 33366 2666 33426 2672
rect 34600 2666 34660 2672
rect 33426 2606 34600 2666
rect 33366 2600 33426 2606
rect 34600 2600 34660 2606
rect 13180 2584 13240 2590
rect 16570 2584 16630 2590
rect 15552 2548 15612 2554
rect 17588 2548 17648 2554
rect 18608 2548 18668 2554
rect 19624 2548 19684 2554
rect 20644 2548 20704 2554
rect 21662 2548 21722 2554
rect 23692 2548 23752 2554
rect 25730 2548 25790 2554
rect 27766 2548 27826 2554
rect 28788 2548 28848 2554
rect 29808 2548 29868 2554
rect 30822 2548 30882 2554
rect 31844 2548 31904 2554
rect 15612 2488 17588 2548
rect 17648 2488 18608 2548
rect 18668 2488 19624 2548
rect 19684 2488 20644 2548
rect 20704 2488 21662 2548
rect 21722 2488 23692 2548
rect 23752 2488 25730 2548
rect 25790 2488 27766 2548
rect 27826 2488 28788 2548
rect 28848 2488 29808 2548
rect 29868 2488 30822 2548
rect 30882 2488 31844 2548
rect 15552 2482 15612 2488
rect 17588 2482 17648 2488
rect 18608 2482 18668 2488
rect 19624 2482 19684 2488
rect 20644 2482 20704 2488
rect 21662 2482 21722 2488
rect 23692 2482 23752 2488
rect 25730 2482 25790 2488
rect 27766 2482 27826 2488
rect 28788 2482 28848 2488
rect 29808 2482 29868 2488
rect 30822 2482 30882 2488
rect 31844 2482 31904 2488
rect 16570 2444 16630 2450
rect 21506 2444 21566 2450
rect 27912 2444 27972 2450
rect 30822 2444 30882 2450
rect 34004 2444 34064 2450
rect 16630 2384 21506 2444
rect 21566 2384 27912 2444
rect 27972 2384 30822 2444
rect 30882 2384 34004 2444
rect 16570 2378 16630 2384
rect 21506 2378 21566 2384
rect 27912 2378 27972 2384
rect 30822 2378 30882 2384
rect 34004 2378 34064 2384
rect -3432 1842 -1262 1924
rect 264 1913 273 2003
rect 363 1990 372 2003
rect 2958 1990 3018 1996
rect 3990 1990 4050 1996
rect 7050 1990 7110 1996
rect 8046 1990 8106 1996
rect 363 1930 2958 1990
rect 3018 1930 3990 1990
rect 4050 1930 7050 1990
rect 7110 1930 8046 1990
rect 363 1913 372 1930
rect 2958 1924 3018 1930
rect 3990 1924 4050 1930
rect 7050 1924 7110 1930
rect 8046 1924 8106 1930
rect 5524 1860 5584 1866
rect 9584 1860 9644 1866
rect 11766 1860 11826 1866
rect 1438 1800 1444 1860
rect 1504 1800 5524 1860
rect 5584 1800 9584 1860
rect 9644 1800 11766 1860
rect 5524 1794 5584 1800
rect 9584 1794 9644 1800
rect 11766 1794 11826 1800
rect 13398 1546 13458 1552
rect 16568 1546 16628 1552
rect 13458 1486 16568 1546
rect 13398 1480 13458 1486
rect 16568 1480 16628 1486
rect 20798 1548 20858 1554
rect 22676 1548 22736 1554
rect 24714 1548 24774 1554
rect 26584 1548 26644 1554
rect 32860 1548 32920 1554
rect 20858 1488 22676 1548
rect 22736 1488 24714 1548
rect 24774 1488 26584 1548
rect 26644 1488 32860 1548
rect 20798 1482 20858 1488
rect 22676 1482 22736 1488
rect 24714 1482 24774 1488
rect 26584 1482 26644 1488
rect 32860 1482 32920 1488
rect 13070 1442 13130 1448
rect 14534 1442 14594 1448
rect 16574 1442 16634 1448
rect 18604 1442 18664 1448
rect 20644 1442 20704 1448
rect 22680 1442 22740 1448
rect 24716 1442 24776 1448
rect 26750 1442 26810 1448
rect 28790 1442 28850 1448
rect 30820 1442 30880 1448
rect 32860 1442 32920 1448
rect 34712 1442 34772 1448
rect 13130 1382 14534 1442
rect 14594 1382 16574 1442
rect 16634 1382 18604 1442
rect 18664 1382 20644 1442
rect 20704 1382 22680 1442
rect 22740 1382 24716 1442
rect 24776 1382 26750 1442
rect 26810 1382 28790 1442
rect 28850 1382 30820 1442
rect 30880 1382 32860 1442
rect 32920 1382 34712 1442
rect 13070 1376 13130 1382
rect 14534 1376 14594 1382
rect 16574 1376 16634 1382
rect 18604 1376 18664 1382
rect 20644 1376 20704 1382
rect 22680 1376 22740 1382
rect 24716 1376 24776 1382
rect 26750 1376 26810 1382
rect 28790 1376 28850 1382
rect 30820 1376 30880 1382
rect 32860 1376 32920 1382
rect 34712 1376 34772 1382
rect 15042 1336 15102 1342
rect 16062 1336 16122 1342
rect 17086 1336 17146 1342
rect 18104 1336 18164 1342
rect 19118 1336 19178 1342
rect 20150 1336 20210 1342
rect 21162 1336 21222 1342
rect 22170 1336 22230 1342
rect 23188 1336 23248 1342
rect 24214 1336 24274 1342
rect 25216 1336 25276 1342
rect 26236 1336 26296 1342
rect 27256 1336 27316 1342
rect 28282 1336 28342 1342
rect 29300 1336 29360 1342
rect 30314 1336 30374 1342
rect 31328 1336 31388 1342
rect 32350 1336 32410 1342
rect 15102 1276 16062 1336
rect 16122 1276 17086 1336
rect 17146 1276 18104 1336
rect 18164 1276 19118 1336
rect 19178 1276 20150 1336
rect 20210 1276 21162 1336
rect 21222 1276 22170 1336
rect 22230 1276 23188 1336
rect 23248 1276 24214 1336
rect 24274 1276 25216 1336
rect 25276 1276 26236 1336
rect 26296 1276 27256 1336
rect 27316 1276 28282 1336
rect 28342 1276 29300 1336
rect 29360 1276 30314 1336
rect 30374 1276 31328 1336
rect 31388 1276 32350 1336
rect 15042 1270 15102 1276
rect 16062 1270 16122 1276
rect 17086 1270 17146 1276
rect 18104 1270 18164 1276
rect 19118 1270 19178 1276
rect 20150 1270 20210 1276
rect 21162 1270 21222 1276
rect 22170 1270 22230 1276
rect 23188 1270 23248 1276
rect 24214 1270 24274 1276
rect 25216 1270 25276 1276
rect 26236 1270 26296 1276
rect 27256 1270 27316 1276
rect 28282 1270 28342 1276
rect 29300 1270 29360 1276
rect 30314 1270 30374 1276
rect 31328 1270 31388 1276
rect 32350 1270 32410 1276
rect 15554 1226 15614 1232
rect 17590 1226 17650 1232
rect 19628 1226 19688 1232
rect 21666 1226 21726 1232
rect 23702 1226 23762 1232
rect 25738 1226 25798 1232
rect 27770 1226 27830 1232
rect 29802 1226 29862 1232
rect 31842 1226 31902 1232
rect 15614 1166 17590 1226
rect 17650 1166 19628 1226
rect 19688 1166 21666 1226
rect 21726 1166 23702 1226
rect 23762 1166 25738 1226
rect 25798 1166 27770 1226
rect 27830 1166 29802 1226
rect 29862 1166 31842 1226
rect 15554 1160 15614 1166
rect 17590 1160 17650 1166
rect 19628 1160 19688 1166
rect 21666 1160 21726 1166
rect 23702 1160 23762 1166
rect 25738 1160 25798 1166
rect 27770 1160 27830 1166
rect 29802 1160 29862 1166
rect 31842 1160 31902 1166
rect 2922 494 2982 500
rect 4960 494 5020 500
rect 6996 494 7056 500
rect 9032 494 9092 500
rect 2982 434 4960 494
rect 5020 434 6996 494
rect 7056 434 9032 494
rect 2922 428 2982 434
rect 4960 428 5020 434
rect 6996 428 7056 434
rect 9032 428 9092 434
rect 3940 382 4000 388
rect 8014 382 8074 388
rect 12020 382 12080 388
rect 4000 322 8014 382
rect 8074 322 12020 382
rect 3940 316 4000 322
rect 8014 316 8074 322
rect 12020 316 12080 322
rect 13398 304 13458 310
rect 14534 304 14594 310
rect 18604 304 18664 310
rect 28784 304 28844 310
rect 34004 304 34064 310
rect -1046 292 -986 298
rect -986 232 -694 292
rect 13458 244 14534 304
rect 14594 244 18604 304
rect 18664 244 28784 304
rect 28844 244 34004 304
rect 37136 254 37236 12600
rect 38186 12594 38246 12600
rect 56550 12576 56610 12582
rect 58590 12576 58650 12582
rect 60630 12576 60690 12582
rect 62660 12576 62720 12582
rect 64700 12576 64760 12582
rect 66732 12576 66792 12582
rect 68772 12576 68832 12582
rect 70808 12576 70868 12582
rect 72842 12576 72902 12582
rect 56610 12516 58590 12576
rect 58650 12516 60630 12576
rect 60690 12516 62660 12576
rect 62720 12516 64700 12576
rect 64760 12516 66732 12576
rect 66792 12516 68772 12576
rect 68832 12516 70808 12576
rect 70868 12516 72842 12576
rect 56550 12510 56610 12516
rect 58590 12510 58650 12516
rect 60630 12510 60690 12516
rect 62660 12510 62720 12516
rect 64700 12510 64760 12516
rect 66732 12510 66792 12516
rect 68772 12510 68832 12516
rect 70808 12510 70868 12516
rect 72842 12510 72902 12516
rect 54174 12456 54234 12462
rect 54518 12456 54578 12462
rect 54234 12396 54518 12456
rect 54174 12390 54234 12396
rect 54518 12390 54578 12396
rect 56042 12450 56102 12456
rect 64186 12450 64246 12456
rect 56102 12390 57056 12450
rect 57116 12390 58078 12450
rect 58138 12390 59092 12450
rect 59152 12390 60118 12450
rect 60178 12390 61130 12450
rect 61190 12390 62166 12450
rect 62226 12390 63172 12450
rect 63232 12390 64186 12450
rect 64246 12390 65202 12450
rect 65262 12390 66210 12450
rect 66270 12390 67226 12450
rect 67286 12390 68250 12450
rect 68310 12390 69272 12450
rect 69332 12390 70294 12450
rect 70354 12390 71312 12450
rect 71372 12390 72326 12450
rect 72386 12390 73350 12450
rect 73410 12390 73416 12450
rect 56042 12384 56102 12390
rect 64186 12384 64246 12390
rect 54392 12334 54452 12340
rect 59606 12334 59666 12340
rect 69794 12334 69854 12340
rect 73866 12334 73926 12340
rect 74998 12334 75058 12340
rect 54452 12274 59606 12334
rect 59666 12274 69794 12334
rect 69854 12274 73866 12334
rect 73926 12274 74998 12334
rect 54392 12268 54452 12274
rect 59606 12268 59666 12274
rect 69794 12268 69854 12274
rect 73866 12268 73926 12274
rect 74998 12268 75058 12274
rect 56554 11412 56614 11418
rect 58594 11412 58654 11418
rect 60626 11412 60686 11418
rect 62658 11412 62718 11418
rect 64694 11412 64754 11418
rect 66730 11412 66790 11418
rect 68768 11412 68828 11418
rect 70806 11412 70866 11418
rect 72842 11412 72902 11418
rect 56614 11352 58594 11412
rect 58654 11352 60626 11412
rect 60686 11352 62658 11412
rect 62718 11352 64694 11412
rect 64754 11352 66730 11412
rect 66790 11352 68768 11412
rect 68828 11352 70806 11412
rect 70866 11352 72842 11412
rect 56554 11346 56614 11352
rect 58594 11346 58654 11352
rect 60626 11346 60686 11352
rect 62658 11346 62718 11352
rect 64694 11346 64754 11352
rect 66730 11346 66790 11352
rect 68768 11346 68828 11352
rect 70806 11346 70866 11352
rect 72842 11346 72902 11352
rect 56046 11302 56106 11308
rect 57068 11302 57128 11308
rect 58082 11302 58142 11308
rect 59096 11302 59156 11308
rect 60114 11302 60174 11308
rect 61140 11302 61200 11308
rect 62160 11302 62220 11308
rect 63180 11302 63240 11308
rect 64182 11302 64242 11308
rect 65208 11302 65268 11308
rect 66226 11302 66286 11308
rect 67234 11302 67294 11308
rect 68246 11302 68306 11308
rect 69278 11302 69338 11308
rect 70292 11302 70352 11308
rect 71310 11302 71370 11308
rect 72334 11302 72394 11308
rect 73354 11302 73414 11308
rect 56106 11242 57068 11302
rect 57128 11242 58082 11302
rect 58142 11242 59096 11302
rect 59156 11242 60114 11302
rect 60174 11242 61140 11302
rect 61200 11242 62160 11302
rect 62220 11242 63180 11302
rect 63240 11242 64182 11302
rect 64242 11242 65208 11302
rect 65268 11242 66226 11302
rect 66286 11242 67234 11302
rect 67294 11242 68246 11302
rect 68306 11242 69278 11302
rect 69338 11242 70292 11302
rect 70352 11242 71310 11302
rect 71370 11242 72334 11302
rect 72394 11242 73354 11302
rect 56046 11236 56106 11242
rect 57068 11236 57128 11242
rect 58082 11236 58142 11242
rect 59096 11236 59156 11242
rect 60114 11236 60174 11242
rect 61140 11236 61200 11242
rect 62160 11236 62220 11242
rect 63180 11236 63240 11242
rect 64182 11236 64242 11242
rect 65208 11236 65268 11242
rect 66226 11236 66286 11242
rect 67234 11236 67294 11242
rect 68246 11236 68306 11242
rect 69278 11236 69338 11242
rect 70292 11236 70352 11242
rect 71310 11236 71370 11242
rect 72334 11236 72394 11242
rect 73354 11236 73414 11242
rect 54070 11196 54130 11202
rect 55536 11196 55596 11202
rect 57576 11196 57636 11202
rect 59606 11196 59666 11202
rect 61646 11196 61706 11202
rect 63680 11196 63740 11202
rect 65716 11196 65776 11202
rect 67752 11196 67812 11202
rect 69792 11196 69852 11202
rect 71822 11196 71882 11202
rect 73862 11196 73922 11202
rect 54130 11136 55536 11196
rect 55596 11136 57576 11196
rect 57636 11136 59606 11196
rect 59666 11136 61646 11196
rect 61706 11136 63680 11196
rect 63740 11136 65716 11196
rect 65776 11136 67752 11196
rect 67812 11136 69792 11196
rect 69852 11136 71822 11196
rect 71882 11136 73862 11196
rect 54070 11130 54130 11136
rect 55536 11130 55596 11136
rect 57576 11130 57636 11136
rect 59606 11130 59666 11136
rect 61646 11130 61706 11136
rect 63680 11130 63740 11136
rect 65716 11130 65776 11136
rect 67752 11130 67812 11136
rect 69792 11130 69852 11136
rect 71822 11130 71882 11136
rect 73862 11130 73922 11136
rect 54522 11090 54582 11096
rect 55020 11090 55080 11096
rect 55532 11090 55592 11096
rect 61812 11090 61872 11096
rect 63680 11090 63740 11096
rect 65718 11090 65778 11096
rect 67598 11090 67658 11096
rect 53830 11030 53836 11090
rect 53896 11030 54522 11090
rect 54582 11030 55020 11090
rect 55080 11030 55532 11090
rect 55592 11030 61812 11090
rect 61872 11030 63680 11090
rect 63740 11030 65718 11090
rect 65778 11030 67598 11090
rect 54522 11024 54582 11030
rect 55020 11024 55080 11030
rect 55532 11024 55592 11030
rect 61812 11024 61872 11030
rect 63680 11024 63740 11030
rect 65718 11024 65778 11030
rect 67598 11024 67658 11030
rect 71822 11092 71882 11098
rect 74998 11092 75058 11098
rect 71882 11032 74998 11092
rect 71822 11026 71882 11032
rect 74998 11026 75058 11032
rect 54392 10200 54452 10206
rect 57570 10200 57630 10206
rect 60626 10200 60686 10206
rect 66732 10200 66792 10206
rect 71826 10200 71886 10206
rect 54452 10140 57570 10200
rect 57630 10140 60626 10200
rect 60686 10140 66732 10200
rect 66792 10140 71826 10200
rect 54392 10134 54452 10140
rect 57570 10134 57630 10140
rect 60626 10134 60686 10140
rect 66732 10134 66792 10140
rect 71826 10134 71886 10140
rect 53962 10096 54022 10102
rect 54516 10096 54576 10102
rect 56036 10096 56096 10102
rect 54022 10036 54516 10096
rect 54576 10036 56036 10096
rect 53962 10030 54022 10036
rect 54516 10030 54576 10036
rect 56036 10030 56096 10036
rect 56548 10096 56608 10102
rect 57572 10096 57632 10102
rect 58584 10096 58644 10102
rect 59604 10096 59664 10102
rect 62662 10096 62722 10102
rect 64700 10096 64760 10102
rect 67750 10096 67810 10102
rect 68768 10096 68828 10102
rect 69788 10096 69848 10102
rect 70804 10096 70864 10102
rect 72840 10096 72900 10102
rect 56608 10036 57572 10096
rect 57632 10036 58584 10096
rect 58644 10036 59604 10096
rect 59664 10036 62662 10096
rect 62722 10036 64700 10096
rect 64760 10036 67750 10096
rect 67810 10036 68768 10096
rect 68828 10036 69788 10096
rect 69848 10036 70804 10096
rect 70864 10036 72840 10096
rect 56548 10030 56608 10036
rect 57572 10030 57632 10036
rect 58584 10030 58644 10036
rect 59604 10030 59664 10036
rect 62662 10030 62722 10036
rect 64700 10030 64760 10036
rect 67750 10030 67810 10036
rect 68768 10030 68828 10036
rect 69788 10030 69848 10036
rect 70804 10030 70864 10036
rect 72840 10030 72900 10036
rect 54286 9974 54346 9980
rect 61646 9974 61706 9980
rect 63680 9974 63740 9980
rect 65710 9974 65770 9980
rect 75710 9974 75770 18932
rect 54346 9914 61646 9974
rect 61706 9914 63680 9974
rect 63740 9914 65710 9974
rect 65770 9914 75770 9974
rect 54286 9908 54346 9914
rect 61646 9908 61706 9914
rect 63680 9908 63740 9914
rect 65710 9908 65770 9914
rect 54174 9860 54234 9866
rect 55022 9860 55082 9866
rect 54234 9800 55022 9860
rect 54174 9794 54234 9800
rect 55022 9794 55082 9800
rect 56554 9862 56614 9868
rect 58590 9862 58650 9868
rect 74984 9862 75044 9868
rect 56614 9802 58590 9862
rect 58650 9802 74984 9862
rect 56554 9796 56614 9802
rect 58590 9796 58650 9802
rect 74984 9796 75044 9802
rect 75112 9844 75172 9850
rect 75712 9844 75772 9850
rect 75172 9784 75712 9844
rect 75112 9778 75172 9784
rect 75712 9778 75772 9784
rect 74878 8974 74938 8980
rect 75838 8974 75898 19250
rect 57570 8956 57630 8962
rect 59606 8956 59666 8962
rect 67750 8956 67810 8962
rect 69786 8956 69846 8962
rect 73860 8956 73920 8962
rect 54398 8932 54458 8938
rect 55536 8932 55596 8938
rect 54458 8872 55536 8932
rect 55596 8872 56418 8932
rect 57630 8896 59606 8956
rect 59666 8896 67750 8956
rect 67810 8896 69786 8956
rect 69846 8896 73860 8956
rect 74938 8914 75898 8974
rect 74878 8908 74938 8914
rect 57570 8890 57630 8896
rect 59606 8890 59666 8896
rect 67750 8890 67810 8896
rect 69786 8890 69846 8896
rect 73860 8890 73920 8896
rect 54398 8866 54458 8872
rect 55536 8866 55596 8872
rect 54286 8732 54346 8738
rect 55534 8732 55594 8738
rect 54346 8672 55534 8732
rect 56358 8736 56418 8872
rect 56552 8852 56612 8858
rect 58592 8852 58652 8858
rect 60624 8852 60684 8858
rect 62658 8852 62718 8858
rect 64698 8852 64758 8858
rect 66732 8852 66792 8858
rect 56612 8792 58592 8852
rect 58652 8792 60624 8852
rect 60684 8792 62658 8852
rect 62718 8792 64698 8852
rect 64758 8792 66732 8852
rect 56552 8786 56612 8792
rect 58592 8786 58652 8792
rect 60624 8786 60684 8792
rect 62658 8786 62718 8792
rect 64698 8786 64758 8792
rect 66732 8786 66792 8792
rect 66928 8848 66988 8854
rect 71820 8848 71880 8854
rect 66988 8788 71820 8848
rect 75478 8844 75538 8850
rect 66928 8782 66988 8788
rect 71820 8782 71880 8788
rect 72318 8784 72324 8844
rect 72384 8784 75478 8844
rect 75478 8778 75538 8784
rect 57066 8738 57126 8744
rect 60624 8740 60684 8746
rect 62660 8740 62720 8746
rect 64696 8740 64756 8746
rect 66732 8740 66792 8746
rect 68766 8740 68826 8746
rect 70804 8740 70864 8746
rect 72844 8740 72904 8746
rect 75228 8740 75288 8746
rect 56358 8678 57066 8736
rect 57126 8678 58070 8738
rect 58130 8678 59082 8738
rect 59142 8678 60102 8738
rect 60162 8678 60168 8738
rect 60684 8680 62660 8740
rect 62720 8680 64696 8740
rect 64756 8680 66732 8740
rect 66792 8680 68766 8740
rect 68826 8680 70804 8740
rect 70864 8680 72844 8740
rect 72904 8680 75228 8740
rect 56358 8676 57408 8678
rect 57066 8672 57126 8676
rect 60624 8674 60684 8680
rect 62660 8674 62720 8680
rect 64696 8674 64756 8680
rect 66732 8674 66792 8680
rect 68766 8674 68826 8680
rect 70804 8674 70864 8680
rect 72844 8674 72904 8680
rect 75228 8674 75288 8680
rect 54286 8666 54346 8672
rect 55534 8666 55594 8672
rect 53610 8630 53670 8636
rect 54180 8630 54240 8636
rect 61642 8630 61702 8636
rect 63676 8630 63736 8636
rect 65716 8630 65776 8636
rect 66928 8630 66988 8636
rect 53670 8570 54180 8630
rect 54240 8570 61642 8630
rect 61702 8570 63676 8630
rect 63736 8570 65716 8630
rect 65776 8570 66928 8630
rect 53610 8564 53670 8570
rect 54180 8564 54240 8570
rect 61642 8564 61702 8570
rect 63676 8564 63736 8570
rect 65716 8564 65776 8570
rect 66928 8564 66988 8570
rect 67222 8632 67282 8638
rect 67282 8572 68250 8632
rect 68310 8572 68316 8632
rect 68768 8626 68828 8632
rect 70804 8626 70864 8632
rect 72842 8626 72902 8632
rect 74984 8626 75044 8632
rect 67222 8566 67282 8572
rect 68828 8566 70804 8626
rect 70864 8566 72842 8626
rect 72902 8566 74984 8626
rect 68768 8560 68828 8566
rect 70804 8560 70864 8566
rect 72842 8560 72902 8566
rect 74984 8560 75044 8566
rect 71316 7712 71376 7718
rect 55534 7700 55594 7706
rect 57572 7700 57632 7706
rect 59608 7700 59668 7706
rect 61640 7700 61700 7706
rect 55594 7640 57572 7700
rect 57632 7640 59608 7700
rect 59668 7640 61640 7700
rect 66216 7652 66222 7712
rect 66282 7652 71316 7712
rect 71316 7646 71376 7652
rect 71454 7716 71514 7722
rect 72336 7716 72396 7722
rect 73342 7716 73402 7722
rect 71514 7656 72336 7716
rect 72396 7656 73342 7716
rect 71454 7650 71514 7656
rect 72336 7650 72396 7656
rect 73342 7650 73402 7656
rect 73860 7712 73920 7718
rect 75112 7712 75172 7718
rect 73920 7652 75112 7712
rect 73860 7646 73920 7652
rect 75112 7646 75172 7652
rect 55534 7634 55594 7640
rect 57572 7634 57632 7640
rect 59608 7634 59668 7640
rect 61640 7634 61700 7640
rect 56040 7598 56100 7604
rect 61132 7598 61192 7604
rect 53100 7548 53160 7554
rect 56100 7538 61132 7598
rect 56040 7532 56100 7538
rect 61132 7532 61192 7538
rect 65716 7584 65776 7590
rect 73860 7584 73920 7590
rect 65776 7524 73860 7584
rect 65716 7518 65776 7524
rect 73860 7518 73920 7524
rect 48552 6622 48612 6628
rect 53100 6622 53160 7488
rect 54286 7496 54346 7502
rect 57570 7496 57630 7502
rect 54346 7436 57570 7496
rect 54286 7430 54346 7436
rect 57570 7430 57630 7436
rect 58078 7490 58138 7496
rect 59100 7490 59160 7496
rect 60114 7490 60174 7496
rect 61132 7490 61192 7496
rect 62152 7490 62212 7496
rect 69264 7490 69324 7496
rect 70294 7490 70354 7496
rect 71454 7490 71514 7496
rect 58138 7430 59100 7490
rect 59160 7430 60114 7490
rect 60174 7430 61132 7490
rect 61192 7430 62152 7490
rect 62212 7430 69264 7490
rect 69324 7430 70294 7490
rect 70354 7430 71454 7490
rect 58078 7424 58138 7430
rect 59100 7424 59160 7430
rect 60114 7424 60174 7430
rect 61132 7424 61192 7430
rect 62152 7424 62212 7430
rect 69264 7424 69324 7430
rect 70294 7424 70354 7430
rect 71454 7424 71514 7430
rect 71822 7490 71882 7496
rect 75350 7490 75410 7496
rect 71882 7430 75350 7490
rect 71822 7424 71882 7430
rect 75350 7424 75410 7430
rect 56554 7396 56614 7402
rect 58588 7396 58648 7402
rect 60624 7396 60684 7402
rect 56614 7336 58588 7396
rect 58648 7336 60624 7396
rect 56554 7330 56614 7336
rect 58588 7330 58648 7336
rect 60624 7330 60684 7336
rect 67752 7386 67812 7392
rect 71822 7386 71882 7392
rect 67812 7326 71822 7386
rect 67752 7320 67812 7326
rect 71822 7320 71882 7326
rect 72838 7388 72898 7394
rect 75228 7388 75288 7394
rect 72898 7328 75228 7388
rect 72838 7322 72898 7328
rect 75228 7322 75288 7328
rect 48612 6562 53160 6622
rect 48552 6556 48612 6562
rect 46522 6476 46582 6482
rect 50582 6476 50642 6482
rect 52766 6476 52826 6482
rect 53232 6476 53292 6482
rect 62660 6478 62720 6484
rect 64696 6478 64756 6484
rect 66732 6478 66792 6484
rect 68770 6478 68830 6484
rect 42436 6416 42442 6476
rect 42502 6416 46522 6476
rect 46582 6416 50582 6476
rect 50642 6416 52766 6476
rect 52826 6416 53232 6476
rect 46522 6410 46582 6416
rect 50582 6410 50642 6416
rect 52766 6410 52826 6416
rect 53232 6410 53292 6416
rect 56036 6472 56096 6478
rect 56946 6472 57006 6478
rect 57948 6472 58008 6478
rect 59100 6472 59160 6478
rect 60110 6472 60170 6478
rect 61116 6472 61176 6478
rect 62160 6472 62220 6478
rect 56096 6412 56946 6472
rect 57006 6412 57948 6472
rect 58008 6412 59100 6472
rect 59160 6412 60110 6472
rect 60170 6412 61116 6472
rect 61176 6412 62160 6472
rect 62720 6418 64696 6478
rect 64756 6418 66732 6478
rect 66792 6418 68770 6478
rect 62660 6412 62720 6418
rect 64696 6412 64756 6418
rect 66732 6412 66792 6418
rect 68770 6412 68830 6418
rect 70806 6478 70866 6484
rect 72844 6478 72904 6484
rect 70866 6418 72844 6478
rect 70806 6412 70866 6418
rect 72844 6412 72904 6418
rect 56036 6406 56096 6412
rect 56946 6406 57006 6412
rect 57948 6406 58008 6412
rect 59100 6406 59160 6412
rect 60110 6406 60170 6412
rect 61116 6406 61176 6412
rect 62160 6406 62220 6412
rect 58588 6370 58648 6376
rect 68762 6370 68822 6376
rect 70802 6370 70862 6376
rect 72840 6370 72900 6376
rect 41288 6348 41348 6354
rect 43966 6348 44026 6354
rect 44998 6348 45058 6354
rect 48058 6348 48118 6354
rect 49054 6348 49114 6354
rect 53352 6348 53412 6354
rect 41279 6288 41288 6348
rect 41348 6288 43966 6348
rect 44026 6288 44998 6348
rect 45058 6288 48058 6348
rect 48118 6288 49054 6348
rect 49114 6288 53352 6348
rect 58648 6310 68762 6370
rect 68822 6310 70802 6370
rect 70862 6310 72840 6370
rect 58588 6304 58648 6310
rect 68762 6304 68822 6310
rect 70802 6304 70862 6310
rect 72840 6304 72900 6310
rect 41288 6282 41348 6288
rect 43966 6282 44026 6288
rect 44998 6282 45058 6288
rect 48058 6282 48118 6288
rect 49054 6282 49114 6288
rect 53352 6282 53412 6288
rect 56036 6256 56096 6262
rect 58088 6256 58148 6262
rect 61114 6256 61174 6262
rect 62154 6256 62214 6262
rect 63168 6256 63228 6262
rect 64176 6256 64236 6262
rect 65220 6256 65280 6262
rect 66210 6256 66270 6262
rect 67228 6256 67288 6262
rect 68262 6256 68322 6262
rect 71294 6256 71354 6262
rect 72332 6256 72392 6262
rect 73358 6256 73418 6262
rect 56096 6196 57074 6256
rect 57134 6196 58088 6256
rect 58148 6196 61114 6256
rect 61174 6196 62154 6256
rect 62214 6196 63168 6256
rect 63228 6196 64176 6256
rect 64236 6196 65220 6256
rect 65280 6196 66210 6256
rect 66270 6196 67228 6256
rect 67288 6196 68262 6256
rect 68322 6196 71294 6256
rect 71354 6196 72332 6256
rect 72392 6196 73358 6256
rect 73418 6196 75476 6256
rect 75536 6196 75542 6256
rect 56036 6190 56096 6196
rect 58088 6190 58148 6196
rect 61114 6190 61174 6196
rect 62154 6190 62214 6196
rect 63168 6190 63228 6196
rect 64176 6190 64236 6196
rect 65220 6190 65280 6196
rect 66210 6190 66270 6196
rect 67228 6190 67288 6196
rect 68262 6190 68322 6196
rect 71294 6190 71354 6196
rect 72332 6190 72392 6196
rect 73358 6190 73418 6196
rect 61638 6152 61698 6158
rect 63680 6152 63740 6158
rect 65718 6152 65778 6158
rect 67752 6152 67812 6158
rect 69786 6154 69846 6160
rect 71820 6154 71880 6160
rect 73862 6154 73922 6160
rect 75112 6154 75172 6160
rect 54394 6092 54400 6152
rect 54460 6092 61638 6152
rect 61698 6092 63680 6152
rect 63740 6092 65718 6152
rect 65778 6092 67752 6152
rect 61638 6086 61698 6092
rect 63680 6086 63740 6092
rect 65718 6086 65778 6092
rect 67752 6086 67812 6092
rect 68264 6148 68324 6154
rect 69286 6148 69346 6154
rect 68324 6088 69286 6148
rect 69846 6094 71820 6154
rect 71880 6094 73862 6154
rect 73922 6094 75112 6154
rect 69786 6088 69846 6094
rect 71820 6088 71880 6094
rect 73862 6088 73922 6094
rect 75112 6088 75172 6094
rect 68264 6082 68324 6088
rect 69286 6082 69346 6088
rect 42946 5386 43006 5392
rect 43970 5386 44030 5392
rect 45002 5386 45062 5392
rect 46002 5386 46062 5392
rect 47022 5386 47082 5392
rect 48042 5386 48102 5392
rect 50066 5386 50126 5392
rect 52886 5386 52946 5392
rect 53492 5386 53552 5392
rect 43006 5326 43970 5386
rect 44030 5326 45002 5386
rect 45062 5326 46002 5386
rect 46062 5326 47022 5386
rect 47082 5326 48042 5386
rect 48102 5326 49052 5386
rect 49112 5326 50066 5386
rect 50126 5326 51084 5386
rect 51144 5326 52886 5386
rect 52946 5326 53492 5386
rect 42946 5320 43006 5326
rect 43970 5320 44030 5326
rect 45002 5320 45062 5326
rect 46002 5320 46062 5326
rect 47022 5320 47082 5326
rect 48042 5320 48102 5326
rect 50066 5320 50126 5326
rect 52886 5320 52946 5326
rect 53492 5320 53552 5326
rect 42446 5282 42506 5288
rect 44482 5282 44542 5288
rect 46518 5282 46578 5288
rect 48552 5282 48612 5288
rect 50588 5282 50648 5288
rect 41288 5252 41348 5261
rect 41282 5192 41288 5252
rect 41348 5192 41354 5252
rect 42506 5222 44482 5282
rect 44542 5222 46518 5282
rect 46578 5222 48552 5282
rect 48612 5222 50588 5282
rect 60628 5250 60688 5256
rect 64696 5250 64756 5256
rect 66730 5250 66790 5256
rect 42446 5216 42506 5222
rect 44482 5216 44542 5222
rect 46518 5216 46578 5222
rect 48552 5216 48612 5222
rect 50588 5216 50648 5222
rect 56034 5244 56094 5250
rect 57042 5244 57102 5250
rect 58056 5244 58116 5250
rect 59094 5244 59154 5250
rect 60112 5244 60172 5250
rect 41288 5183 41348 5192
rect 56094 5184 57042 5244
rect 57102 5184 58056 5244
rect 58116 5184 59094 5244
rect 59154 5184 60112 5244
rect 60688 5190 62664 5250
rect 62724 5190 64696 5250
rect 64756 5190 66730 5250
rect 60628 5184 60688 5190
rect 64696 5184 64756 5190
rect 66730 5184 66790 5190
rect 67752 5252 67812 5258
rect 68106 5252 68166 5258
rect 67812 5192 68106 5252
rect 67752 5186 67812 5192
rect 68106 5186 68166 5192
rect 71824 5252 71884 5258
rect 75108 5252 75168 5258
rect 71884 5192 75108 5252
rect 71824 5186 71884 5192
rect 75108 5186 75168 5192
rect 47532 5178 47592 5184
rect 54070 5178 54130 5184
rect 56034 5178 56094 5184
rect 57042 5178 57102 5184
rect 58056 5178 58116 5184
rect 59094 5178 59154 5184
rect 60112 5178 60172 5184
rect 43458 5118 43464 5178
rect 43524 5118 45500 5178
rect 45560 5118 47532 5178
rect 47592 5118 49566 5178
rect 49626 5118 51610 5178
rect 51670 5118 54070 5178
rect 47532 5112 47592 5118
rect 54070 5112 54130 5118
rect 54180 5140 54240 5146
rect 55536 5140 55596 5146
rect 63680 5140 63740 5146
rect 65716 5140 65776 5146
rect 67748 5140 67808 5146
rect 54240 5080 55536 5140
rect 55596 5080 63680 5140
rect 63740 5080 65716 5140
rect 65776 5080 67748 5140
rect 54180 5074 54240 5080
rect 55536 5074 55596 5080
rect 63680 5074 63740 5080
rect 65716 5074 65776 5080
rect 67748 5074 67808 5080
rect 67258 5042 67318 5048
rect 68296 5042 68356 5048
rect 69272 5042 69332 5048
rect 70288 5042 70348 5048
rect 72314 5042 72374 5048
rect 73344 5042 73404 5048
rect 53838 5028 53898 5034
rect 56552 5028 56612 5034
rect 58590 5028 58650 5034
rect 62662 5028 62722 5034
rect 53898 4968 56552 5028
rect 56612 4968 58590 5028
rect 58650 4968 62662 5028
rect 67318 4982 68296 5042
rect 68356 4982 69272 5042
rect 69332 4982 70288 5042
rect 70348 4982 72314 5042
rect 72374 4982 73344 5042
rect 67258 4976 67318 4982
rect 68296 4976 68356 4982
rect 69272 4976 69332 4982
rect 70288 4976 70348 4982
rect 72314 4976 72374 4982
rect 73344 4976 73404 4982
rect 53838 4962 53898 4968
rect 56552 4962 56612 4968
rect 58590 4962 58650 4968
rect 62662 4962 62722 4968
rect 55532 4930 55592 4936
rect 57570 4930 57630 4936
rect 59610 4930 59670 4936
rect 61646 4930 61706 4936
rect 67750 4930 67810 4936
rect 68100 4930 68106 4934
rect 55592 4870 57570 4930
rect 57630 4870 59610 4930
rect 59670 4870 61646 4930
rect 61706 4874 68106 4930
rect 68166 4930 68172 4934
rect 69786 4930 69846 4936
rect 71822 4930 71882 4936
rect 73858 4930 73918 4936
rect 68166 4874 69786 4930
rect 61706 4870 69786 4874
rect 69846 4870 71822 4930
rect 71882 4870 73858 4930
rect 55532 4864 55592 4870
rect 57570 4864 57630 4870
rect 59610 4864 59670 4870
rect 61646 4864 61706 4870
rect 67750 4864 67810 4870
rect 69786 4864 69846 4870
rect 71822 4864 71882 4870
rect 73858 4864 73918 4870
rect 44476 4236 44536 4242
rect 48552 4236 48612 4242
rect 52766 4236 52826 4242
rect 44536 4176 48552 4236
rect 48612 4176 52766 4236
rect 44476 4170 44536 4176
rect 48552 4170 48612 4176
rect 52766 4170 52826 4176
rect 41288 4116 41348 4122
rect 42938 4116 42998 4122
rect 46008 4116 46068 4122
rect 47016 4116 47076 4122
rect 50078 4116 50138 4122
rect 51104 4116 51164 4122
rect 41348 4056 42938 4116
rect 42998 4056 46008 4116
rect 46068 4056 47016 4116
rect 47076 4056 50078 4116
rect 50138 4056 51104 4116
rect 41288 4050 41348 4056
rect 42938 4050 42998 4056
rect 46008 4050 46068 4056
rect 47016 4050 47076 4056
rect 50078 4050 50138 4056
rect 51104 4050 51164 4056
rect 62658 4026 62718 4032
rect 64700 4026 64760 4032
rect 66732 4026 66792 4032
rect 68772 4026 68832 4032
rect 75228 4026 75288 4032
rect 56552 4006 56612 4012
rect 58588 4006 58648 4012
rect 60626 4006 60686 4012
rect 56612 3946 58588 4006
rect 58648 3946 60626 4006
rect 62482 3966 62488 4026
rect 62548 3966 62658 4026
rect 62718 3966 64700 4026
rect 64760 3966 66732 4026
rect 66792 3966 68772 4026
rect 68832 3966 75228 4026
rect 62658 3960 62718 3966
rect 64700 3960 64760 3966
rect 66732 3960 66792 3966
rect 68772 3960 68832 3966
rect 75228 3960 75288 3966
rect 56552 3940 56612 3946
rect 58588 3940 58648 3946
rect 60626 3940 60686 3946
rect 67750 3928 67810 3934
rect 73856 3928 73916 3934
rect 75108 3928 75168 3934
rect 54398 3908 54458 3914
rect 57570 3908 57630 3914
rect 54458 3848 57570 3908
rect 54398 3842 54458 3848
rect 57570 3842 57630 3848
rect 59094 3908 59154 3914
rect 62142 3908 62202 3914
rect 59154 3848 60116 3908
rect 60176 3848 61138 3908
rect 61198 3848 62142 3908
rect 67810 3868 73856 3928
rect 73916 3868 75108 3928
rect 67750 3862 67810 3868
rect 73856 3862 73916 3868
rect 75108 3862 75168 3868
rect 59094 3842 59154 3848
rect 62142 3842 62202 3848
rect 62664 3818 62724 3824
rect 64692 3818 64752 3824
rect 66736 3818 66796 3824
rect 68764 3818 68824 3824
rect 70802 3818 70862 3824
rect 72842 3818 72902 3824
rect 56556 3812 56616 3818
rect 58592 3812 58652 3818
rect 60620 3812 60680 3818
rect 62488 3812 62548 3818
rect 56616 3752 58592 3812
rect 58652 3752 60620 3812
rect 60680 3752 62488 3812
rect 62724 3758 64692 3818
rect 64752 3758 66736 3818
rect 66796 3758 68764 3818
rect 68824 3758 70802 3818
rect 70862 3758 72842 3818
rect 62664 3752 62724 3758
rect 64692 3752 64752 3758
rect 66736 3752 66796 3758
rect 68764 3752 68824 3758
rect 70802 3752 70862 3758
rect 72842 3752 72902 3758
rect 73360 3822 73420 3828
rect 74872 3822 74932 3828
rect 75478 3822 75538 3828
rect 73420 3762 74872 3822
rect 74932 3762 75478 3822
rect 73360 3756 73420 3762
rect 74872 3756 74932 3762
rect 75478 3756 75538 3762
rect 56556 3746 56616 3752
rect 58592 3746 58652 3752
rect 60620 3746 60680 3752
rect 62488 3746 62548 3752
rect 55538 3692 55598 3698
rect 59606 3692 59666 3698
rect 61640 3692 61700 3698
rect 69790 3692 69850 3698
rect 71820 3692 71880 3698
rect 73860 3694 73920 3700
rect 75350 3694 75410 3700
rect 55598 3632 59606 3692
rect 59666 3632 61640 3692
rect 61700 3632 69790 3692
rect 69850 3632 71820 3692
rect 72340 3634 72346 3694
rect 72406 3634 73860 3694
rect 73920 3634 75350 3694
rect 55538 3626 55598 3632
rect 59606 3626 59666 3632
rect 61640 3626 61700 3632
rect 69790 3626 69850 3632
rect 71820 3626 71880 3632
rect 73860 3628 73920 3634
rect 75350 3628 75410 3634
rect 51610 3172 51670 3178
rect 43458 3112 43464 3172
rect 43524 3112 45500 3172
rect 45560 3112 47532 3172
rect 47592 3112 49566 3172
rect 49626 3112 51610 3172
rect 51610 3106 51670 3112
rect 42450 3064 42510 3070
rect 44486 3064 44546 3070
rect 46522 3064 46582 3070
rect 48556 3064 48616 3070
rect 50592 3064 50652 3070
rect 42510 3004 44486 3064
rect 44546 3004 46522 3064
rect 46582 3004 48556 3064
rect 48616 3004 50592 3064
rect 42450 2998 42510 3004
rect 44486 2998 44546 3004
rect 46522 2998 46582 3004
rect 48556 2998 48616 3004
rect 50592 2998 50652 3004
rect 42944 2952 43004 2958
rect 43968 2952 44028 2958
rect 45000 2952 45060 2958
rect 46000 2952 46060 2958
rect 47020 2952 47080 2958
rect 48040 2952 48100 2958
rect 50064 2952 50124 2958
rect 52886 2952 52946 2958
rect 43004 2892 43968 2952
rect 44028 2892 45000 2952
rect 45060 2892 46000 2952
rect 46060 2892 47020 2952
rect 47080 2892 48040 2952
rect 48100 2892 49050 2952
rect 49110 2892 50064 2952
rect 50124 2892 51082 2952
rect 51142 2892 52886 2952
rect 52946 2892 53274 2952
rect 42944 2886 43004 2892
rect 43968 2886 44028 2892
rect 45000 2886 45060 2892
rect 46000 2886 46060 2892
rect 47020 2886 47080 2892
rect 48040 2886 48100 2892
rect 50064 2886 50124 2892
rect 52886 2886 52946 2892
rect 54286 2776 54346 2782
rect 63674 2776 63734 2782
rect 65716 2776 65776 2782
rect 67752 2776 67812 2782
rect 54346 2716 63674 2776
rect 63734 2716 65716 2776
rect 65776 2716 67752 2776
rect 54286 2710 54346 2716
rect 63674 2710 63734 2716
rect 65716 2710 65776 2716
rect 67752 2710 67812 2716
rect 70806 2776 70866 2782
rect 72838 2776 72898 2782
rect 74984 2776 75044 2782
rect 70866 2716 72838 2776
rect 72898 2716 74984 2776
rect 70806 2710 70866 2716
rect 72838 2710 72898 2716
rect 74984 2710 75044 2716
rect 58090 2662 58150 2668
rect 63170 2662 63230 2668
rect 54180 2650 54240 2656
rect 57570 2650 57630 2656
rect 54240 2590 57570 2650
rect 58150 2602 63170 2662
rect 58090 2596 58150 2602
rect 63170 2596 63230 2602
rect 68258 2666 68318 2672
rect 73358 2666 73418 2672
rect 68318 2606 73358 2666
rect 68258 2600 68318 2606
rect 73358 2600 73418 2606
rect 74366 2666 74426 2672
rect 75600 2666 75660 2672
rect 74426 2606 75600 2666
rect 74366 2600 74426 2606
rect 75600 2600 75660 2606
rect 54180 2584 54240 2590
rect 57570 2584 57630 2590
rect 56552 2548 56612 2554
rect 58588 2548 58648 2554
rect 59608 2548 59668 2554
rect 60624 2548 60684 2554
rect 61644 2548 61704 2554
rect 62662 2548 62722 2554
rect 64692 2548 64752 2554
rect 66730 2548 66790 2554
rect 68766 2548 68826 2554
rect 69788 2548 69848 2554
rect 70808 2548 70868 2554
rect 71822 2548 71882 2554
rect 72844 2548 72904 2554
rect 56612 2488 58588 2548
rect 58648 2488 59608 2548
rect 59668 2488 60624 2548
rect 60684 2488 61644 2548
rect 61704 2488 62662 2548
rect 62722 2488 64692 2548
rect 64752 2488 66730 2548
rect 66790 2488 68766 2548
rect 68826 2488 69788 2548
rect 69848 2488 70808 2548
rect 70868 2488 71822 2548
rect 71882 2488 72844 2548
rect 56552 2482 56612 2488
rect 58588 2482 58648 2488
rect 59608 2482 59668 2488
rect 60624 2482 60684 2488
rect 61644 2482 61704 2488
rect 62662 2482 62722 2488
rect 64692 2482 64752 2488
rect 66730 2482 66790 2488
rect 68766 2482 68826 2488
rect 69788 2482 69848 2488
rect 70808 2482 70868 2488
rect 71822 2482 71882 2488
rect 72844 2482 72904 2488
rect 57570 2444 57630 2450
rect 62506 2444 62566 2450
rect 68912 2444 68972 2450
rect 71822 2444 71882 2450
rect 75004 2444 75064 2450
rect 57630 2384 62506 2444
rect 62566 2384 68912 2444
rect 68972 2384 71822 2444
rect 71882 2384 75004 2444
rect 57570 2378 57630 2384
rect 62506 2378 62566 2384
rect 68912 2378 68972 2384
rect 71822 2378 71882 2384
rect 75004 2378 75064 2384
rect 41288 1990 41348 1996
rect 43958 1990 44018 1996
rect 44990 1990 45050 1996
rect 48050 1990 48110 1996
rect 49046 1990 49106 1996
rect 41348 1930 43958 1990
rect 44018 1930 44990 1990
rect 45050 1930 48050 1990
rect 48110 1930 49046 1990
rect 41288 1924 41348 1930
rect 43958 1924 44018 1930
rect 44990 1924 45050 1930
rect 48050 1924 48110 1930
rect 49046 1924 49106 1930
rect 46524 1860 46584 1866
rect 50584 1860 50644 1866
rect 52766 1860 52826 1866
rect 42438 1800 42444 1860
rect 42504 1800 46524 1860
rect 46584 1800 50584 1860
rect 50644 1800 52766 1860
rect 46524 1794 46584 1800
rect 50584 1794 50644 1800
rect 52766 1794 52826 1800
rect 54398 1546 54458 1552
rect 57568 1546 57628 1552
rect 54458 1486 57568 1546
rect 54398 1480 54458 1486
rect 57568 1480 57628 1486
rect 61798 1548 61858 1554
rect 63676 1548 63736 1554
rect 65714 1548 65774 1554
rect 67584 1548 67644 1554
rect 73860 1548 73920 1554
rect 61858 1488 63676 1548
rect 63736 1488 65714 1548
rect 65774 1488 67584 1548
rect 67644 1488 73860 1548
rect 61798 1482 61858 1488
rect 63676 1482 63736 1488
rect 65714 1482 65774 1488
rect 67584 1482 67644 1488
rect 73860 1482 73920 1488
rect 54070 1442 54130 1448
rect 55534 1442 55594 1448
rect 57574 1442 57634 1448
rect 59604 1442 59664 1448
rect 61644 1442 61704 1448
rect 63680 1442 63740 1448
rect 65716 1442 65776 1448
rect 67750 1442 67810 1448
rect 69790 1442 69850 1448
rect 71820 1442 71880 1448
rect 73860 1442 73920 1448
rect 75712 1442 75772 1448
rect 54130 1382 55534 1442
rect 55594 1382 57574 1442
rect 57634 1382 59604 1442
rect 59664 1382 61644 1442
rect 61704 1382 63680 1442
rect 63740 1382 65716 1442
rect 65776 1382 67750 1442
rect 67810 1382 69790 1442
rect 69850 1382 71820 1442
rect 71880 1382 73860 1442
rect 73920 1382 75712 1442
rect 54070 1376 54130 1382
rect 55534 1376 55594 1382
rect 57574 1376 57634 1382
rect 59604 1376 59664 1382
rect 61644 1376 61704 1382
rect 63680 1376 63740 1382
rect 65716 1376 65776 1382
rect 67750 1376 67810 1382
rect 69790 1376 69850 1382
rect 71820 1376 71880 1382
rect 73860 1376 73920 1382
rect 75712 1376 75772 1382
rect 56042 1336 56102 1342
rect 57062 1336 57122 1342
rect 58086 1336 58146 1342
rect 59104 1336 59164 1342
rect 60118 1336 60178 1342
rect 61150 1336 61210 1342
rect 62162 1336 62222 1342
rect 63170 1336 63230 1342
rect 64188 1336 64248 1342
rect 65214 1336 65274 1342
rect 66216 1336 66276 1342
rect 67236 1336 67296 1342
rect 68256 1336 68316 1342
rect 69282 1336 69342 1342
rect 70300 1336 70360 1342
rect 71314 1336 71374 1342
rect 72328 1336 72388 1342
rect 73350 1336 73410 1342
rect 56102 1276 57062 1336
rect 57122 1276 58086 1336
rect 58146 1276 59104 1336
rect 59164 1276 60118 1336
rect 60178 1276 61150 1336
rect 61210 1276 62162 1336
rect 62222 1276 63170 1336
rect 63230 1276 64188 1336
rect 64248 1276 65214 1336
rect 65274 1276 66216 1336
rect 66276 1276 67236 1336
rect 67296 1276 68256 1336
rect 68316 1276 69282 1336
rect 69342 1276 70300 1336
rect 70360 1276 71314 1336
rect 71374 1276 72328 1336
rect 72388 1276 73350 1336
rect 56042 1270 56102 1276
rect 57062 1270 57122 1276
rect 58086 1270 58146 1276
rect 59104 1270 59164 1276
rect 60118 1270 60178 1276
rect 61150 1270 61210 1276
rect 62162 1270 62222 1276
rect 63170 1270 63230 1276
rect 64188 1270 64248 1276
rect 65214 1270 65274 1276
rect 66216 1270 66276 1276
rect 67236 1270 67296 1276
rect 68256 1270 68316 1276
rect 69282 1270 69342 1276
rect 70300 1270 70360 1276
rect 71314 1270 71374 1276
rect 72328 1270 72388 1276
rect 73350 1270 73410 1276
rect 56554 1226 56614 1232
rect 58590 1226 58650 1232
rect 60628 1226 60688 1232
rect 62666 1226 62726 1232
rect 64702 1226 64762 1232
rect 66738 1226 66798 1232
rect 68770 1226 68830 1232
rect 70802 1226 70862 1232
rect 72842 1226 72902 1232
rect 56614 1166 58590 1226
rect 58650 1166 60628 1226
rect 60688 1166 62666 1226
rect 62726 1166 64702 1226
rect 64762 1166 66738 1226
rect 66798 1166 68770 1226
rect 68830 1166 70802 1226
rect 70862 1166 72842 1226
rect 56554 1160 56614 1166
rect 58590 1160 58650 1166
rect 60628 1160 60688 1166
rect 62666 1160 62726 1166
rect 64702 1160 64762 1166
rect 66738 1160 66798 1166
rect 68770 1160 68830 1166
rect 70802 1160 70862 1166
rect 72842 1160 72902 1166
rect 43922 494 43982 500
rect 45960 494 46020 500
rect 47996 494 48056 500
rect 50032 494 50092 500
rect 43982 434 45960 494
rect 46020 434 47996 494
rect 48056 434 50032 494
rect 43922 428 43982 434
rect 45960 428 46020 434
rect 47996 428 48056 434
rect 50032 428 50092 434
rect 44940 382 45000 388
rect 49014 382 49074 388
rect 53020 382 53080 388
rect 45000 322 49014 382
rect 49074 322 53020 382
rect 44940 316 45000 322
rect 49014 316 49074 322
rect 53020 316 53080 322
rect 54398 304 54458 310
rect 55534 304 55594 310
rect 59604 304 59664 310
rect 69784 304 69844 310
rect 75004 304 75064 310
rect 13398 238 13458 244
rect 14534 238 14594 244
rect 18604 238 18664 244
rect 28784 238 28844 244
rect 34004 238 34064 244
rect -1046 226 -986 232
rect -1012 168 -922 180
rect -1012 104 -1000 168
rect -934 104 -922 168
rect -1012 94 -922 104
rect -1046 42 -986 48
rect -834 42 -774 232
rect 15046 196 15106 202
rect 23190 196 23250 202
rect 15106 136 16060 196
rect 16120 136 17082 196
rect 17142 136 18096 196
rect 18156 136 19122 196
rect 19182 136 20134 196
rect 20194 136 21170 196
rect 21230 136 22176 196
rect 22236 136 23190 196
rect 23250 136 24206 196
rect 24266 136 25214 196
rect 25274 136 26230 196
rect 26290 136 27254 196
rect 27314 136 28276 196
rect 28336 136 29298 196
rect 29358 136 30316 196
rect 30376 136 31330 196
rect 31390 136 32354 196
rect 32414 136 32420 196
rect 37127 154 37136 254
rect 37236 154 37245 254
rect 54458 244 55534 304
rect 55594 244 59604 304
rect 59664 244 69784 304
rect 69844 244 75004 304
rect 54398 238 54458 244
rect 55534 238 55594 244
rect 59604 238 59664 244
rect 69784 238 69844 244
rect 75004 238 75064 244
rect 56046 196 56106 202
rect 64190 196 64250 202
rect 56106 136 57060 196
rect 57120 136 58082 196
rect 58142 136 59096 196
rect 59156 136 60122 196
rect 60182 136 61134 196
rect 61194 136 62170 196
rect 62230 136 63176 196
rect 63236 136 64190 196
rect 64250 136 65206 196
rect 65266 136 66214 196
rect 66274 136 67230 196
rect 67290 136 68254 196
rect 68314 136 69276 196
rect 69336 136 70298 196
rect 70358 136 71316 196
rect 71376 136 72330 196
rect 72390 136 73354 196
rect 73414 136 73420 196
rect 15046 130 15106 136
rect 23190 130 23250 136
rect 56046 130 56106 136
rect 64190 130 64250 136
rect -986 -18 -774 42
rect -1046 -24 -986 -18
rect -1212 -76 -806 -64
rect -1212 -142 -1198 -76
rect -814 -142 -806 -76
rect -1212 -154 -806 -142
rect 2832 -106 34918 -60
rect 2832 -260 2878 -106
rect 34878 -260 34918 -106
rect 2832 -306 34918 -260
rect 43832 -106 75918 -60
rect 43832 -260 43878 -106
rect 75878 -260 75918 -106
rect 43832 -306 75918 -260
rect -1266 -446 -666 -436
rect -1266 -756 -666 -746
rect 35166 -446 35766 -436
rect 35166 -756 35766 -746
rect 39734 -446 40334 -436
rect 39734 -756 40334 -746
rect 76166 -446 76766 -436
rect 76166 -756 76766 -746
<< via2 >>
rect 11434 30286 12034 30586
rect 35066 30286 35666 30586
rect 52434 30286 53034 30586
rect 76066 30286 76666 30586
rect 15011 29990 31796 30204
rect 56011 29990 72796 30204
rect -2680 15700 8084 15992
rect 8084 15700 8172 15992
rect 12492 15344 12552 15404
rect 13269 15331 13359 15421
rect -2276 13782 -1748 14300
rect -3342 1924 -2908 13306
rect 34708 9914 34768 9974
rect 38320 15700 49084 15992
rect 49084 15700 49172 15992
rect 54269 15331 54359 15421
rect 36824 13564 37424 13864
rect 37976 13564 38576 13864
rect 36928 13300 38480 13396
rect 39132 13134 39192 13194
rect 34110 5192 34168 5252
rect 34168 5192 34170 5252
rect 273 1990 363 2003
rect 273 1930 288 1990
rect 288 1930 348 1990
rect 348 1930 363 1990
rect 273 1913 363 1930
rect 41288 6288 41348 6348
rect 41288 5192 41348 5252
rect -1000 166 -934 168
rect -1000 106 -998 166
rect -998 106 -938 166
rect -938 106 -934 166
rect -1000 104 -934 106
rect 37136 154 37236 254
rect -1198 -142 -814 -76
rect 2878 -260 34878 -106
rect 43878 -260 75878 -106
rect -1266 -746 -666 -446
rect 35166 -746 35766 -446
rect 39734 -746 40334 -446
rect 76166 -746 76766 -446
<< metal3 >>
rect 11424 30586 12044 30591
rect 11424 30286 11434 30586
rect 12034 30286 12044 30586
rect 11424 30281 12044 30286
rect 35056 30586 35676 30591
rect 35056 30286 35066 30586
rect 35666 30286 35676 30586
rect 35056 30281 35676 30286
rect 52424 30586 53044 30591
rect 52424 30286 52434 30586
rect 53034 30286 53044 30586
rect 52424 30281 53044 30286
rect 76056 30586 76676 30591
rect 76056 30286 76066 30586
rect 76666 30286 76676 30586
rect 76056 30281 76676 30286
rect 14948 30204 31828 30236
rect 14948 29990 15011 30204
rect 31796 29990 31828 30204
rect 14948 29970 31828 29990
rect 55948 30204 72828 30236
rect 55948 29990 56011 30204
rect 72796 29990 72828 30204
rect 55948 29970 72828 29990
rect 14948 29968 19302 29970
rect 55948 29968 60302 29970
rect -4218 29310 10822 29456
rect -4218 29300 9976 29310
rect -4218 28610 -4066 29300
rect -3370 28612 9976 29300
rect 10666 28612 10822 29310
rect -3370 28610 10822 28612
rect -4218 28280 10822 28610
rect -4218 15618 -3036 28280
rect -2748 17080 9158 28020
rect 9522 17080 10822 28280
rect -2748 15992 10822 17080
rect 8172 15700 10822 15992
rect 8084 15618 10822 15700
rect -4218 15392 10822 15618
rect 36782 29310 51822 29456
rect 36782 29300 50976 29310
rect 36782 28610 36934 29300
rect 37630 28612 50976 29300
rect 51666 28612 51822 29310
rect 37630 28610 51822 28612
rect 36782 28280 51822 28610
rect 36782 15618 37964 28280
rect 38252 17080 50158 28020
rect 50522 17080 51822 28280
rect 38252 15992 51822 17080
rect 49172 15700 51822 15992
rect 49084 15618 51822 15700
rect 13265 15426 13363 15431
rect 12430 15424 12624 15426
rect 13264 15425 13364 15426
rect 12430 15409 12636 15424
rect -4218 15292 9324 15392
rect 12430 15345 12487 15409
rect 12557 15345 12636 15409
rect 12430 15344 12492 15345
rect 12552 15344 12636 15345
rect 12430 15328 12636 15344
rect 12430 15324 12624 15328
rect 13264 15327 13265 15425
rect 13363 15327 13364 15425
rect 13264 15326 13364 15327
rect 36782 15392 51822 15618
rect 54265 15426 54363 15431
rect 54264 15425 54364 15426
rect 13265 15321 13363 15326
rect -4218 14610 -4064 15292
rect -3730 14610 9324 15292
rect -4218 14544 9324 14610
rect -16568 14454 9324 14544
rect 36782 15292 50324 15392
rect 54264 15327 54265 15425
rect 54363 15327 54364 15425
rect 54264 15326 54364 15327
rect 54265 15321 54363 15326
rect 36782 14610 36936 15292
rect 37270 14610 50324 15292
rect 36782 14454 50324 14610
rect -16568 14398 -1528 14454
rect -16568 14388 -2374 14398
rect -16568 13698 -16416 14388
rect -15720 13700 -2374 14388
rect -1684 13700 -1528 14398
rect 52113 14346 52211 14351
rect 39110 14345 52212 14346
rect 39110 14247 52113 14345
rect 52211 14247 52212 14345
rect 39110 14246 52212 14247
rect -15720 13698 -1528 13700
rect -16568 13368 -1528 13698
rect 36814 13864 37434 13869
rect 36814 13564 36824 13864
rect 37424 13564 37434 13864
rect 36814 13559 37434 13564
rect 37966 13864 38586 13869
rect 37966 13564 37976 13864
rect 38576 13564 38586 13864
rect 37966 13559 38586 13564
rect -16568 706 -15386 13368
rect -15066 1844 -3376 12976
rect -2828 1844 -1528 13368
rect 36890 13396 38514 13426
rect 36890 13300 36928 13396
rect 38480 13300 38514 13396
rect 36890 13272 38514 13300
rect 39110 13194 39210 14246
rect 52113 14241 52211 14246
rect 39110 13134 39132 13194
rect 39192 13134 39210 13194
rect 39110 13114 39210 13134
rect 34688 9974 41370 9992
rect 34688 9914 34708 9974
rect 34768 9914 41370 9974
rect 34688 9892 41370 9914
rect 41270 6348 41370 9892
rect 41270 6288 41288 6348
rect 41348 6288 41370 6348
rect 41270 6270 41370 6288
rect 34086 5252 41380 5270
rect 34086 5192 34110 5252
rect 34170 5192 41288 5252
rect 41348 5192 41380 5252
rect 34086 5170 41380 5192
rect -15066 1070 -1528 1844
rect -4132 706 -1528 1070
rect -16568 360 -1528 706
rect 268 2003 368 2008
rect 268 1913 273 2003
rect 363 1913 368 2003
rect 268 634 368 1913
rect -1016 514 -916 520
rect 268 513 370 634
rect 263 415 269 513
rect 367 415 373 513
rect 268 414 370 415
rect -16568 -458 -2656 360
rect -1016 168 -916 414
rect -1016 104 -1000 168
rect -934 104 -916 168
rect 270 254 370 414
rect 37131 254 37241 259
rect 270 154 37136 254
rect 37236 154 37241 254
rect 37131 149 37241 154
rect -1016 94 -916 104
rect -1212 -76 -806 -64
rect -1212 -142 -1198 -76
rect -814 -142 -806 -76
rect -1212 -154 -806 -142
rect 2832 -106 34918 -60
rect 2832 -260 2878 -106
rect 34878 -260 34918 -106
rect 2832 -306 34918 -260
rect 43832 -106 75918 -60
rect 43832 -260 43878 -106
rect 75878 -260 75918 -106
rect 43832 -306 75918 -260
rect -1276 -446 -656 -441
rect -1276 -746 -1266 -446
rect -666 -746 -656 -446
rect -1276 -751 -656 -746
rect 35156 -446 35776 -441
rect 35156 -746 35166 -446
rect 35766 -746 35776 -446
rect 35156 -751 35776 -746
rect 39724 -446 40344 -441
rect 39724 -746 39734 -446
rect 40334 -746 40344 -446
rect 39724 -751 40344 -746
rect 76156 -446 76776 -441
rect 76156 -746 76166 -446
rect 76766 -746 76776 -446
rect 76156 -751 76776 -746
<< via3 >>
rect 11434 30286 12034 30586
rect 35066 30286 35666 30586
rect 52434 30286 53034 30586
rect 76066 30286 76666 30586
rect 15011 29990 31796 30204
rect 56011 29990 72796 30204
rect -4066 28610 -3370 29300
rect 9976 28612 10666 29310
rect -3036 28020 9522 28280
rect -3036 15992 -2748 28020
rect 9158 17080 9522 28020
rect -3036 15700 -2680 15992
rect -2680 15700 8084 15992
rect -3036 15618 8084 15700
rect 36934 28610 37630 29300
rect 50976 28612 51666 29310
rect 37964 28020 50522 28280
rect 37964 15992 38252 28020
rect 50158 17080 50522 28020
rect 37964 15700 38320 15992
rect 38320 15700 49084 15992
rect 37964 15618 49084 15700
rect 12487 15404 12557 15409
rect 12487 15345 12492 15404
rect 12492 15345 12552 15404
rect 12552 15345 12557 15404
rect 13265 15421 13363 15425
rect 13265 15331 13269 15421
rect 13269 15331 13359 15421
rect 13359 15331 13363 15421
rect 13265 15327 13363 15331
rect -4064 14610 -3730 15292
rect 54265 15421 54363 15425
rect 54265 15331 54269 15421
rect 54269 15331 54359 15421
rect 54359 15331 54363 15421
rect 54265 15327 54363 15331
rect 36936 14610 37270 15292
rect -16416 13698 -15720 14388
rect -2374 14300 -1684 14398
rect -2374 13782 -2276 14300
rect -2276 13782 -1748 14300
rect -1748 13782 -1684 14300
rect -2374 13700 -1684 13782
rect 52113 14247 52211 14345
rect 36824 13564 37424 13864
rect 37976 13564 38576 13864
rect -15386 13306 -2828 13368
rect -15386 12976 -3342 13306
rect -15386 1070 -15066 12976
rect -3376 1924 -3342 12976
rect -3342 1924 -2908 13306
rect -2908 1924 -2828 13306
rect -3376 1844 -2828 1924
rect 36928 13300 38480 13396
rect -15386 706 -4132 1070
rect -1016 414 -916 514
rect 269 415 367 513
rect -1198 -142 -814 -76
rect 2878 -260 34878 -106
rect 43878 -260 75878 -106
rect -1266 -746 -666 -446
rect 35166 -746 35766 -446
rect 39734 -746 40334 -446
rect 76166 -746 76766 -446
<< mimcap >>
rect -3032 29306 3168 29356
rect -3032 29006 2818 29306
rect 3118 29006 3168 29306
rect -3032 28956 3168 29006
rect 3368 29306 9568 29356
rect 3368 29006 9218 29306
rect 9518 29006 9568 29306
rect 3368 28956 9568 29006
rect 37968 29306 44168 29356
rect 37968 29006 43818 29306
rect 44118 29006 44168 29306
rect 37968 28956 44168 29006
rect 44368 29306 50568 29356
rect 44368 29006 50218 29306
rect 50518 29006 50568 29306
rect 44368 28956 50568 29006
rect -4118 28224 -3318 28274
rect -4118 22524 -3668 28224
rect -3368 22524 -3318 28224
rect 9926 28224 10726 28274
rect -2178 27306 3022 27356
rect -2178 22606 2672 27306
rect 2972 22606 3022 27306
rect -2178 22556 3022 22606
rect 3422 27306 8622 27356
rect 3422 22606 8272 27306
rect 8572 22606 8622 27306
rect 3422 22556 8622 22606
rect -4118 22474 -3318 22524
rect 9926 22524 10376 28224
rect 10676 22524 10726 28224
rect 9926 22474 10726 22524
rect 36882 28224 37682 28274
rect 36882 22524 37332 28224
rect 37632 22524 37682 28224
rect 50926 28224 51726 28274
rect 38822 27306 44022 27356
rect 38822 22606 43672 27306
rect 43972 22606 44022 27306
rect 38822 22556 44022 22606
rect 44422 27306 49622 27356
rect 44422 22606 49272 27306
rect 49572 22606 49622 27306
rect 44422 22556 49622 22606
rect 36882 22474 37682 22524
rect 50926 22524 51376 28224
rect 51676 22524 51726 28224
rect 50926 22474 51726 22524
rect -4118 21732 -3318 21782
rect -4118 16032 -3668 21732
rect -3368 16032 -3318 21732
rect -2178 21706 3022 21756
rect -2178 17006 2672 21706
rect 2972 17006 3022 21706
rect -2178 16956 3022 17006
rect 3422 21706 8622 21756
rect 3422 17006 8272 21706
rect 8572 17006 8622 21706
rect 3422 16956 8622 17006
rect 9926 21732 10726 21782
rect -4118 15982 -3318 16032
rect 9926 16032 10376 21732
rect 10676 16032 10726 21732
rect 9926 15982 10726 16032
rect 36882 21732 37682 21782
rect 36882 16032 37332 21732
rect 37632 16032 37682 21732
rect 38822 21706 44022 21756
rect 38822 17006 43672 21706
rect 43972 17006 44022 21706
rect 38822 16956 44022 17006
rect 44422 21706 49622 21756
rect 44422 17006 49272 21706
rect 49572 17006 49622 21706
rect 44422 16956 49622 17006
rect 50926 21732 51726 21782
rect 36882 15982 37682 16032
rect 50926 16032 51376 21732
rect 51676 16032 51726 21732
rect 50926 15982 51726 16032
rect -3532 15306 2668 15356
rect -3532 15006 2318 15306
rect 2618 15006 2668 15306
rect -3532 14956 2668 15006
rect 2868 15306 9068 15356
rect 2868 15006 8718 15306
rect 9018 15006 9068 15306
rect 2868 14956 9068 15006
rect 37468 15306 43668 15356
rect 37468 15006 43318 15306
rect 43618 15006 43668 15306
rect 37468 14956 43668 15006
rect 43868 15306 50068 15356
rect 43868 15006 49718 15306
rect 50018 15006 50068 15306
rect 43868 14956 50068 15006
rect -15382 14294 -9182 14344
rect -15382 13994 -9532 14294
rect -9232 13994 -9182 14294
rect -15382 13944 -9182 13994
rect -8982 14294 -2782 14344
rect -8982 13994 -3132 14294
rect -2832 13994 -2782 14294
rect -8982 13944 -2782 13994
rect -16468 13312 -15668 13362
rect -16468 7612 -16018 13312
rect -15718 7612 -15668 13312
rect -2424 13312 -1624 13362
rect -14528 12394 -9328 12444
rect -14528 7694 -9678 12394
rect -9378 7694 -9328 12394
rect -14528 7644 -9328 7694
rect -8928 12394 -3728 12444
rect -8928 7694 -4078 12394
rect -3778 7694 -3728 12394
rect -8928 7644 -3728 7694
rect -16468 7562 -15668 7612
rect -2424 7612 -1974 13312
rect -1674 7612 -1624 13312
rect -2424 7562 -1624 7612
rect -16468 6820 -15668 6870
rect -16468 1120 -16018 6820
rect -15718 1120 -15668 6820
rect -14528 6794 -9328 6844
rect -14528 2094 -9678 6794
rect -9378 2094 -9328 6794
rect -14528 2044 -9328 2094
rect -8928 6794 -3728 6844
rect -8928 2094 -4078 6794
rect -3778 2094 -3728 6794
rect -8928 2044 -3728 2094
rect -2424 6820 -1624 6870
rect -16468 1070 -15668 1120
rect -2424 1120 -1974 6820
rect -1674 1120 -1624 6820
rect -2424 1070 -1624 1120
rect -15882 394 -9682 444
rect -15882 94 -10032 394
rect -9732 94 -9682 394
rect -15882 44 -9682 94
rect -9482 394 -3282 444
rect -9482 94 -3632 394
rect -3332 94 -3282 394
rect -9482 44 -3282 94
<< mimcapcontact >>
rect 2818 29006 3118 29306
rect 9218 29006 9518 29306
rect 43818 29006 44118 29306
rect 50218 29006 50518 29306
rect -3668 22524 -3368 28224
rect 2672 22606 2972 27306
rect 8272 22606 8572 27306
rect 10376 22524 10676 28224
rect 37332 22524 37632 28224
rect 43672 22606 43972 27306
rect 49272 22606 49572 27306
rect 51376 22524 51676 28224
rect -3668 16032 -3368 21732
rect 2672 17006 2972 21706
rect 8272 17006 8572 21706
rect 10376 16032 10676 21732
rect 37332 16032 37632 21732
rect 43672 17006 43972 21706
rect 49272 17006 49572 21706
rect 51376 16032 51676 21732
rect 2318 15006 2618 15306
rect 8718 15006 9018 15306
rect 43318 15006 43618 15306
rect 49718 15006 50018 15306
rect -9532 13994 -9232 14294
rect -3132 13994 -2832 14294
rect -16018 7612 -15718 13312
rect -9678 7694 -9378 12394
rect -4078 7694 -3778 12394
rect -1974 7612 -1674 13312
rect -16018 1120 -15718 6820
rect -9678 2094 -9378 6794
rect -4078 2094 -3778 6794
rect -1974 1120 -1674 6820
rect -10032 94 -9732 394
rect -3632 94 -3332 394
<< metal4 >>
rect -4218 30586 35232 30770
rect 36032 30586 76950 30770
rect -4218 30286 11434 30586
rect 12034 30286 35066 30586
rect 36032 30286 52434 30586
rect 53034 30286 76066 30586
rect 76666 30286 76950 30586
rect -4218 30204 35232 30286
rect -4218 29990 15011 30204
rect 31796 29990 35232 30204
rect -4218 29970 35232 29990
rect 36032 30204 76950 30286
rect 36032 29990 56011 30204
rect 72796 29990 76950 30204
rect 36032 29970 76950 29990
rect -4218 29310 10822 29456
rect -4218 29306 9976 29310
rect -4218 29300 2818 29306
rect -4218 28610 -4066 29300
rect -3370 29006 2818 29300
rect 3118 29006 9218 29306
rect 9518 29006 9976 29306
rect -3370 28612 9976 29006
rect 10666 28612 10822 29310
rect -3370 28610 10822 28612
rect -4218 28280 10822 28610
rect -4218 28224 -3036 28280
rect -4218 22524 -3668 28224
rect -3368 22524 -3036 28224
rect 9522 28224 10822 28280
rect -4218 21732 -3036 22524
rect -4218 16032 -3668 21732
rect -3368 16032 -3036 21732
rect -4218 15618 -3036 16032
rect -2278 27306 8722 27456
rect -2278 22606 2672 27306
rect 2972 22606 8272 27306
rect 8572 22606 8722 27306
rect -2278 21706 8722 22606
rect -2278 17006 2672 21706
rect 2972 17006 8272 21706
rect 8572 17006 8722 21706
rect -2278 16554 8722 17006
rect 9522 22524 10376 28224
rect 10676 22524 10822 28224
rect 9522 21732 10822 22524
rect 9522 16934 10376 21732
rect -2278 16457 9623 16554
rect -2278 16456 8722 16457
rect -2548 15992 8228 16074
rect 8116 15618 8228 15992
rect -4218 15532 8228 15618
rect -4216 15392 8228 15532
rect -4216 15306 9228 15392
rect -4216 15292 2318 15306
rect -4216 14610 -4064 15292
rect -3730 15006 2318 15292
rect 2618 15006 8718 15306
rect 9018 15006 9228 15306
rect -3730 14610 9228 15006
rect 9526 14970 9623 16457
rect 9892 16032 10376 16934
rect 10676 16032 10822 21732
rect 9892 15522 10822 16032
rect 36782 29310 51822 29456
rect 36782 29306 50976 29310
rect 36782 29300 43818 29306
rect 36782 28610 36934 29300
rect 37630 29006 43818 29300
rect 44118 29006 50218 29306
rect 50518 29006 50976 29306
rect 37630 28612 50976 29006
rect 51666 28612 51822 29310
rect 37630 28610 51822 28612
rect 36782 28280 51822 28610
rect 36782 28224 37964 28280
rect 36782 22524 37332 28224
rect 37632 22524 37964 28224
rect 50522 28224 51822 28280
rect 36782 21732 37964 22524
rect 36782 16032 37332 21732
rect 37632 16032 37964 21732
rect 36782 15618 37964 16032
rect 38722 27306 49722 27456
rect 38722 22606 43672 27306
rect 43972 22606 49272 27306
rect 49572 22606 49722 27306
rect 38722 21706 49722 22606
rect 38722 17006 43672 21706
rect 43972 17006 49272 21706
rect 49572 17006 49722 21706
rect 38722 16554 49722 17006
rect 50522 22524 51376 28224
rect 51676 22524 51822 28224
rect 50522 21732 51822 22524
rect 50522 16934 51376 21732
rect 38722 16457 50623 16554
rect 38722 16456 49722 16457
rect 38452 15992 49228 16074
rect 49116 15618 49228 15992
rect 36782 15532 49228 15618
rect 11176 15425 13364 15426
rect 11176 15409 13265 15425
rect 11176 15345 12487 15409
rect 12557 15345 13265 15409
rect 11176 15327 13265 15345
rect 13363 15327 13364 15425
rect 11176 15326 13364 15327
rect 36784 15392 49228 15532
rect 11176 14970 11276 15326
rect 9526 14870 11276 14970
rect 36784 15306 50228 15392
rect 36784 15292 43318 15306
rect -4216 14544 9228 14610
rect -16568 14454 9228 14544
rect 36784 14610 36936 15292
rect 37270 15006 43318 15292
rect 43618 15006 49718 15306
rect 50018 15006 50228 15306
rect 37270 14610 50228 15006
rect 50526 14970 50623 16457
rect 50892 16032 51376 16934
rect 51676 16032 51822 21732
rect 50892 15522 51822 16032
rect 52112 15425 54364 15426
rect 52112 15327 54265 15425
rect 54363 15327 54364 15425
rect 52112 15326 54364 15327
rect 52112 14970 52276 15326
rect 50526 14870 52276 14970
rect 36784 14454 50228 14610
rect -16568 14398 -1528 14454
rect -16568 14388 -2374 14398
rect -16568 13698 -16416 14388
rect -15720 14294 -2374 14388
rect -15720 13994 -9532 14294
rect -9232 13994 -3132 14294
rect -2832 13994 -2374 14294
rect -15720 13700 -2374 13994
rect -1684 13700 -1528 14398
rect 52112 14345 52212 14870
rect 52112 14247 52113 14345
rect 52211 14247 52212 14345
rect 52112 14246 52212 14247
rect 35516 14048 36670 14050
rect -15720 13698 -1528 13700
rect -16568 13368 -1528 13698
rect -16568 13312 -15386 13368
rect -16568 7612 -16018 13312
rect -15718 7612 -15386 13312
rect -2828 13312 -1528 13368
rect -16568 6820 -15386 7612
rect -16568 1120 -16018 6820
rect -15718 1120 -15386 6820
rect -16568 706 -15386 1120
rect -15066 12934 -3376 12976
rect -15066 1084 -15016 12934
rect -14628 12394 -3628 12544
rect -14628 7694 -9678 12394
rect -9378 7694 -4078 12394
rect -3778 7694 -3628 12394
rect -14628 6794 -3628 7694
rect -14628 2094 -9678 6794
rect -9378 2094 -4078 6794
rect -3778 2094 -3628 6794
rect -14628 1544 -3628 2094
rect -3388 1844 -3376 12934
rect -2828 7612 -1974 13312
rect -1674 7612 -1528 13312
rect 35232 14028 38760 14048
rect 35232 13276 35256 14028
rect 36008 13864 38760 14028
rect 36008 13564 36824 13864
rect 37424 13564 37976 13864
rect 38576 13564 38760 13864
rect 36008 13396 38760 13564
rect 36008 13300 36928 13396
rect 38480 13300 38760 13396
rect 36008 13276 38760 13300
rect 35232 13248 38760 13276
rect -2828 6820 -1528 7612
rect -2828 1844 -1974 6820
rect -3388 1760 -1974 1844
rect -3754 1496 -3628 1544
rect -3754 1396 -2814 1496
rect -15066 1070 -3244 1084
rect -4132 706 -3244 1070
rect -16568 620 -3244 706
rect -16566 394 -3244 620
rect -16566 94 -10032 394
rect -9732 94 -3632 394
rect -3332 94 -3244 394
rect -2914 340 -2814 1396
rect -2458 1120 -1974 1760
rect -1674 1120 -1528 6820
rect -2458 1002 -1528 1120
rect -2458 610 -1952 1002
rect -1017 514 -915 515
rect -1400 414 -1016 514
rect -916 513 368 514
rect -916 415 269 513
rect 367 415 368 513
rect -916 414 368 415
rect -1400 340 -1300 414
rect -1017 413 -915 414
rect -2914 240 -1300 340
rect -16566 38 -3244 94
rect -16566 -358 -16436 38
rect -16034 -30 -3244 38
rect -16034 -76 76950 -30
rect -16034 -142 -1198 -76
rect -814 -106 76950 -76
rect -814 -142 2878 -106
rect -16034 -260 2878 -142
rect 34878 -260 43878 -106
rect 75878 -260 76950 -106
rect -16034 -358 76950 -260
rect -16566 -446 76950 -358
rect -16566 -746 -1266 -446
rect -666 -746 35166 -446
rect 35766 -746 39734 -446
rect 40334 -746 76166 -446
rect 76766 -746 76950 -446
rect -16566 -830 76950 -746
<< via4 >>
rect 35232 30586 36032 30770
rect 35232 30286 35666 30586
rect 35666 30286 36032 30586
rect 35232 29970 36032 30286
rect -4066 28610 -3370 29300
rect 9976 28612 10666 29310
rect -3036 28020 9522 28280
rect -3036 15992 -2748 28020
rect -2748 27816 9158 28020
rect -2748 15992 -2548 27816
rect 9066 17080 9158 27816
rect 9158 17080 9522 28020
rect 9066 16934 9522 17080
rect -3036 15618 8084 15992
rect 8084 15618 8116 15992
rect -4064 14610 -3730 15292
rect 36934 28610 37630 29300
rect 50976 28612 51666 29310
rect 37964 28020 50522 28280
rect 37964 15992 38252 28020
rect 38252 27816 50158 28020
rect 38252 15992 38452 27816
rect 50066 17080 50158 27816
rect 50158 17080 50522 28020
rect 50066 16934 50522 17080
rect 37964 15618 49084 15992
rect 49084 15618 49116 15992
rect 36936 14610 37270 15292
rect -16416 13698 -15720 14388
rect -2374 13700 -1684 14398
rect -15386 12976 -2828 13368
rect -15386 1070 -15066 12976
rect -3376 1844 -2828 12976
rect 35256 13276 36008 14028
rect -15386 706 -4134 1070
rect -16436 -358 -16034 38
<< mimcap2 >>
rect -3032 28906 2768 29356
rect -3032 28606 -2982 28906
rect 2718 28606 2768 28906
rect -3032 28556 2768 28606
rect 3368 28906 9168 29356
rect 3368 28606 3418 28906
rect 9118 28606 9168 28906
rect 3368 28556 9168 28606
rect 37968 28906 43768 29356
rect 37968 28606 38018 28906
rect 43718 28606 43768 28906
rect 37968 28556 43768 28606
rect 44368 28906 50168 29356
rect 44368 28606 44418 28906
rect 50118 28606 50168 28906
rect 44368 28556 50168 28606
rect -4118 22424 -3718 28274
rect -4118 22124 -4068 22424
rect -3768 22124 -3718 22424
rect -2178 22506 2622 27356
rect -2178 22206 -2128 22506
rect 2572 22206 2622 22506
rect -2178 22156 2622 22206
rect 3422 22506 8222 27356
rect 3422 22206 3472 22506
rect 8172 22206 8222 22506
rect 3422 22156 8222 22206
rect 9926 22424 10326 28274
rect -4118 22074 -3718 22124
rect 9926 22124 9976 22424
rect 10276 22124 10326 22424
rect 9926 22074 10326 22124
rect 36882 22424 37282 28274
rect 36882 22124 36932 22424
rect 37232 22124 37282 22424
rect 38822 22506 43622 27356
rect 38822 22206 38872 22506
rect 43572 22206 43622 22506
rect 38822 22156 43622 22206
rect 44422 22506 49222 27356
rect 44422 22206 44472 22506
rect 49172 22206 49222 22506
rect 44422 22156 49222 22206
rect 50926 22424 51326 28274
rect 36882 22074 37282 22124
rect 50926 22124 50976 22424
rect 51276 22124 51326 22424
rect 50926 22074 51326 22124
rect -4118 15932 -3718 21782
rect -2178 16906 2622 21756
rect -2178 16606 -2128 16906
rect 2572 16606 2622 16906
rect -2178 16556 2622 16606
rect 3422 16906 8222 21756
rect 3422 16606 3472 16906
rect 8172 16606 8222 16906
rect 3422 16556 8222 16606
rect -4118 15632 -4068 15932
rect -3768 15632 -3718 15932
rect -4118 15582 -3718 15632
rect 9926 15932 10326 21782
rect 9926 15646 9976 15932
rect 10276 15646 10326 15932
rect 9926 15582 10326 15646
rect 36882 15932 37282 21782
rect 38822 16906 43622 21756
rect 38822 16606 38872 16906
rect 43572 16606 43622 16906
rect 38822 16556 43622 16606
rect 44422 16906 49222 21756
rect 44422 16606 44472 16906
rect 49172 16606 49222 16906
rect 44422 16556 49222 16606
rect 36882 15632 36932 15932
rect 37232 15632 37282 15932
rect 36882 15582 37282 15632
rect 50926 15932 51326 21782
rect 50926 15646 50976 15932
rect 51276 15646 51326 15932
rect 50926 15582 51326 15646
rect -3532 14906 2268 15356
rect -3532 14606 -3482 14906
rect 2218 14606 2268 14906
rect -3532 14556 2268 14606
rect 2868 14906 8668 15356
rect 2868 14606 2918 14906
rect 8618 14606 8668 14906
rect 2868 14556 8668 14606
rect 37468 14906 43268 15356
rect 37468 14606 37518 14906
rect 43218 14606 43268 14906
rect 37468 14556 43268 14606
rect 43868 14906 49668 15356
rect 43868 14606 43918 14906
rect 49618 14606 49668 14906
rect 43868 14556 49668 14606
rect -15382 13894 -9582 14344
rect -15382 13594 -15332 13894
rect -9632 13594 -9582 13894
rect -15382 13544 -9582 13594
rect -8982 13894 -3182 14344
rect -8982 13594 -8932 13894
rect -3232 13594 -3182 13894
rect -8982 13544 -3182 13594
rect -16468 7512 -16068 13362
rect -16468 7212 -16418 7512
rect -16118 7212 -16068 7512
rect -14528 7594 -9728 12444
rect -14528 7294 -14478 7594
rect -9778 7294 -9728 7594
rect -14528 7244 -9728 7294
rect -8928 7594 -4128 12444
rect -8928 7294 -8878 7594
rect -4178 7294 -4128 7594
rect -8928 7244 -4128 7294
rect -2424 7512 -2024 13362
rect -16468 7162 -16068 7212
rect -2424 7212 -2374 7512
rect -2074 7212 -2024 7512
rect -2424 7162 -2024 7212
rect -16468 1020 -16068 6870
rect -14528 1994 -9728 6844
rect -14528 1694 -14478 1994
rect -9778 1694 -9728 1994
rect -14528 1644 -9728 1694
rect -8928 1994 -4128 6844
rect -8928 1694 -8878 1994
rect -4178 1694 -4128 1994
rect -8928 1644 -4128 1694
rect -16468 720 -16418 1020
rect -16118 720 -16068 1020
rect -16468 670 -16068 720
rect -2424 1020 -2024 6870
rect -2424 720 -2374 1020
rect -2074 720 -2024 1020
rect -2424 670 -2024 720
rect -15882 -6 -10082 444
rect -15882 -306 -15832 -6
rect -10132 -306 -10082 -6
rect -15882 -356 -10082 -306
rect -9482 -6 -3682 444
rect -9482 -306 -9432 -6
rect -3732 -306 -3682 -6
rect -9482 -356 -3682 -306
<< mimcap2contact >>
rect -2982 28606 2718 28906
rect 3418 28606 9118 28906
rect 38018 28606 43718 28906
rect 44418 28606 50118 28906
rect -4068 22124 -3768 22424
rect -2128 22206 2572 22506
rect 3472 22206 8172 22506
rect 9976 22124 10276 22424
rect 36932 22124 37232 22424
rect 38872 22206 43572 22506
rect 44472 22206 49172 22506
rect 50976 22124 51276 22424
rect -2128 16606 2572 16906
rect 3472 16606 8172 16906
rect -4068 15632 -3768 15932
rect 9976 15646 10276 15932
rect 38872 16606 43572 16906
rect 44472 16606 49172 16906
rect 36932 15632 37232 15932
rect 50976 15646 51276 15932
rect -3482 14606 2218 14906
rect 2918 14606 8618 14906
rect 37518 14606 43218 14906
rect 43918 14606 49618 14906
rect -15332 13594 -9632 13894
rect -8932 13594 -3232 13894
rect -16418 7212 -16118 7512
rect -14478 7294 -9778 7594
rect -8878 7294 -4178 7594
rect -2374 7212 -2074 7512
rect -14478 1694 -9778 1994
rect -8878 1694 -4178 1994
rect -16418 720 -16118 1020
rect -2374 720 -2074 1020
rect -15832 -306 -10132 -6
rect -9432 -306 -3732 -6
<< metal5 >>
rect 35208 30770 36056 30794
rect 35208 29970 35232 30770
rect 36032 29970 36056 30770
rect 35208 29946 36056 29970
rect -4218 29310 10822 29456
rect -4218 29300 9976 29310
rect -4218 28610 -4066 29300
rect -3370 28906 9976 29300
rect -3370 28610 -2982 28906
rect -4218 28606 -2982 28610
rect 2718 28606 3418 28906
rect 9118 28612 9976 28906
rect 10666 28612 10822 29310
rect 9118 28606 10822 28612
rect -4218 28280 10822 28606
rect -4218 22424 -3036 28280
rect -4218 22124 -4068 22424
rect -3768 22124 -3036 22424
rect -4218 15932 -3036 22124
rect -2548 22506 9066 27816
rect -2548 22206 -2128 22506
rect 2572 22206 3472 22506
rect 8172 22206 9066 22506
rect -2548 16934 9066 22206
rect 9522 22424 10822 28280
rect 9522 22124 9976 22424
rect 10276 22124 10822 22424
rect 9522 16934 10822 22124
rect -2548 16906 10822 16934
rect -2548 16606 -2128 16906
rect 2572 16606 3472 16906
rect 8172 16852 10822 16906
rect 8172 16606 8224 16852
rect -2548 15992 8224 16606
rect -4218 15632 -4068 15932
rect -3768 15632 -3036 15932
rect -4218 15618 -3036 15632
rect 8116 15618 8224 15992
rect -4218 15388 8224 15618
rect 9878 15932 10822 16852
rect 9878 15646 9976 15932
rect 10276 15646 10822 15932
rect 9878 15606 10822 15646
rect -4218 15292 9122 15388
rect -4218 14610 -4064 15292
rect -3730 14906 9122 15292
rect -3730 14610 -3482 14906
rect -4218 14606 -3482 14610
rect 2218 14606 2918 14906
rect 8618 14606 9122 14906
rect -4218 14544 9122 14606
rect -16568 14454 9122 14544
rect -16568 14398 -1528 14454
rect -16568 14388 -2374 14398
rect -16568 13698 -16416 14388
rect -15720 13894 -2374 14388
rect -15720 13698 -15332 13894
rect -16568 13594 -15332 13698
rect -9632 13594 -8932 13894
rect -3232 13700 -2374 13894
rect -1684 13700 -1528 14398
rect -3232 13594 -1528 13700
rect -16568 13368 -1528 13594
rect -16568 7512 -15386 13368
rect -16568 7212 -16418 7512
rect -16118 7212 -15386 7512
rect -16568 1020 -15386 7212
rect -15066 7594 -3376 12976
rect -15066 7294 -14478 7594
rect -9778 7294 -8878 7594
rect -4178 7294 -3376 7594
rect -15066 1994 -3376 7294
rect -15066 1694 -14478 1994
rect -9778 1694 -8878 1994
rect -4178 1844 -3376 1994
rect -2828 7512 -1528 13368
rect 35232 14028 36032 29946
rect 36782 29310 51822 29456
rect 36782 29300 50976 29310
rect 36782 28610 36934 29300
rect 37630 28906 50976 29300
rect 37630 28610 38018 28906
rect 36782 28606 38018 28610
rect 43718 28606 44418 28906
rect 50118 28612 50976 28906
rect 51666 28612 51822 29310
rect 50118 28606 51822 28612
rect 36782 28280 51822 28606
rect 36782 22424 37964 28280
rect 36782 22124 36932 22424
rect 37232 22124 37964 22424
rect 36782 15932 37964 22124
rect 38452 22506 50066 27816
rect 38452 22206 38872 22506
rect 43572 22206 44472 22506
rect 49172 22206 50066 22506
rect 38452 16934 50066 22206
rect 50522 22424 51822 28280
rect 50522 22124 50976 22424
rect 51276 22124 51822 22424
rect 50522 16934 51822 22124
rect 38452 16906 51822 16934
rect 38452 16606 38872 16906
rect 43572 16606 44472 16906
rect 49172 16852 51822 16906
rect 49172 16606 49224 16852
rect 38452 15992 49224 16606
rect 36782 15632 36932 15932
rect 37232 15632 37964 15932
rect 36782 15618 37964 15632
rect 49116 15618 49224 15992
rect 36782 15388 49224 15618
rect 50878 15932 51822 16852
rect 50878 15646 50976 15932
rect 51276 15646 51822 15932
rect 50878 15606 51822 15646
rect 36782 15292 50122 15388
rect 36782 14610 36936 15292
rect 37270 14906 50122 15292
rect 37270 14610 37518 14906
rect 36782 14606 37518 14610
rect 43218 14606 43918 14906
rect 49618 14606 50122 14906
rect 36782 14454 50122 14606
rect 35232 13276 35256 14028
rect 36008 13276 36032 14028
rect 35232 13252 36032 13276
rect -2828 7212 -2374 7512
rect -2074 7212 -1528 7512
rect -2828 1844 -1528 7212
rect -4178 1694 -1528 1844
rect -15066 1070 -1528 1694
rect -16568 720 -16418 1020
rect -16118 720 -15386 1020
rect -16568 706 -15386 720
rect -4134 1020 -1528 1070
rect -4134 720 -2374 1020
rect -2074 720 -1528 1020
rect -4134 706 -1528 720
rect -16568 360 -1528 706
rect -16568 38 -2656 360
rect -16568 -358 -16436 38
rect -16034 -6 -2656 38
rect -16034 -306 -15832 -6
rect -10132 -306 -9432 -6
rect -3732 -306 -2656 -6
rect -16034 -358 -2656 -306
rect -16568 -458 -2656 -358
<< labels >>
flabel metal2 38146 12624 38158 12636 1 FreeSans 480 0 0 0 vpeakh
port 6 n
flabel metal1 37310 12672 37326 12682 1 FreeSans 480 0 0 0 verr
flabel metal4 37536 14028 37548 14038 1 FreeSans 480 0 0 0 VDD
port 4 n power bidirectional
flabel metal2 -742 256 -736 264 1 FreeSans 480 0 0 0 rst
port 7 n
flabel metal2 53200 2918 53216 2930 1 FreeSans 480 0 0 0 vin
port 1 n
flabel metal2 12516 15272 12528 15284 1 FreeSans 480 0 0 0 vpeak_out
port 3 n
flabel metal4 36274 -344 36322 -292 1 FreeSans 480 0 0 0 VSS
port 5 n ground bidirectional
flabel metal1 8324 1414 8342 1424 1 FreeSans 480 0 0 0 ibiasn2
port 8 n
flabel metal1 47952 1414 47972 1428 1 FreeSans 480 0 0 0 ibiasn1
port 2 n
flabel metal4 -1544 284 -1530 294 1 FreeSans 480 0 0 0 vpeak
flabel metal1 2872 14018 2872 14018 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal1 4744 7344 4744 7344 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal1 34130 7052 34154 7082 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal1 34506 7900 34506 7900 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias3
flabel metal1 34250 8106 34250 8106 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 34386 3874 34386 3874 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias4
flabel metal1 13088 8268 13116 8298 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal1 13406 11610 13438 11650 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 14272 14472 14362 14502 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal1 13194 8008 13232 8044 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 33888 9740 33924 9770 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal1 304 4830 332 4874 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 11904 4834 11936 4872 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal1 5748 1404 5844 1440 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/ibiasn
flabel metal1 10898 4130 10946 4154 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal4 30 -374 56 -352 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal2 4386 6436 4434 6452 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal1 1462 4202 1494 4230 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal4 -754 30280 -728 30374 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal4 11544 15368 11564 15388 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 33558 17998 33564 18016 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 18448 24820 18480 24852 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
flabel metal1 13882 21362 13954 21392 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 16606 21370 16648 21392 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 15160 21332 15186 21370 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 14648 17324 14678 17350 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 15656 17320 15686 17354 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal2 31122 21980 31184 22008 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 27160 24184 27212 24210 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 21396 23142 21464 23172 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 21620 22110 21672 22144 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 19274 28254 19274 28254 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 20252 27992 20282 28020 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal1 17296 26980 17330 27002 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 18684 26856 18742 26892 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal2 20710 24676 20788 24710 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 28460 20510 28496 20538 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 22816 16462 22870 16496 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal2 23240 21450 23322 21482 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal2 27790 18940 27852 18970 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal2 27382 19252 27446 19284 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal1 18274 21290 18314 21324 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 33344 19152 33406 19184 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal2 31458 19042 31508 19078 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 31510 17994 31602 18026 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 18568 20322 18568 20322 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 18438 16736 18494 16770 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
flabel metal1 43872 14018 43872 14018 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias1
flabel metal1 45744 7344 45744 7344 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias2
flabel metal1 75130 7052 75154 7082 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/VSS
flabel metal1 75506 7900 75506 7900 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias3
flabel metal1 75250 8106 75250 8106 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascnm
flabel metal1 75386 3874 75386 3874 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias4
flabel metal1 54088 8268 54116 8298 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vtail_cascn
flabel metal1 54406 11610 54438 11650 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascnp
flabel metal1 55272 14472 55362 14502 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M8d
flabel metal1 54194 8008 54232 8044 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vmirror
flabel metal1 74888 9740 74924 9770 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M16d
flabel metal1 41304 4830 41332 4874 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vip
flabel metal1 52904 4834 52936 4872 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vim
flabel metal1 46748 1404 46844 1440 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/ibiasn
flabel metal1 51898 4130 51946 4154 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vtail_cascn
flabel metal4 41030 -374 41056 -352 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_1/VSS
flabel metal2 45386 6436 45434 6452 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascpp
flabel metal1 42462 4202 42494 4230 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascpm
flabel metal4 40246 30280 40272 30374 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_1/VDD
flabel metal4 52544 15368 52564 15388 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vo
flabel metal1 74558 17998 74564 18016 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vo
flabel metal1 59448 24820 59480 24852 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M9d
flabel metal1 54882 21362 54954 21392 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascnm
flabel metal1 57606 21370 57648 21392 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascnp
flabel metal1 56160 21332 56186 21370 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vtail_cascp
flabel metal1 55648 17324 55678 17350 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vip
flabel metal1 56656 17320 56686 17354 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vim
flabel metal2 72122 21980 72184 22008 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vmirror
flabel metal1 68160 24184 68212 24210 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/VDD
flabel metal2 62396 23142 62464 23172 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascpp
flabel metal2 62620 22110 62672 22144 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascpm
flabel metal2 60274 28254 60274 28254 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias1
flabel metal2 61252 27992 61282 28020 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/VDD
flabel metal1 58296 26980 58330 27002 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M7d
flabel metal2 59684 26856 59742 26892 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M13d
flabel metal2 61710 24676 61788 24710 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vtail_cascp
flabel metal1 69460 20510 69496 20538 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/VDD
flabel metal2 63816 16462 63870 16496 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M8d
flabel metal2 64240 21450 64322 21482 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias2
flabel metal2 68790 18940 68852 18970 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M16d
flabel metal2 68382 19252 68446 19284 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M13d
flabel metal1 59274 21290 59314 21324 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M7d
flabel metal2 74344 19152 74406 19184 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vmirror
flabel metal2 72458 19042 72508 19078 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascpm
flabel metal2 72510 17994 72602 18026 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vcascpp
flabel metal2 59568 20322 59568 20322 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/vbias1
flabel metal2 59438 16736 59494 16770 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_1/M9d
<< end >>
