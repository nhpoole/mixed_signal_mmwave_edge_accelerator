magic
tech sky130A
magscale 1 2
timestamp 1622264460
<< error_p >>
rect -13822 13650 -13762 15250
rect -13742 13650 -13682 15250
rect -12103 13650 -12043 15250
rect -12023 13650 -11963 15250
rect -10384 13650 -10324 15250
rect -10304 13650 -10244 15250
rect -8665 13650 -8605 15250
rect -8585 13650 -8525 15250
rect -6946 13650 -6886 15250
rect -6866 13650 -6806 15250
rect -5227 13650 -5167 15250
rect -5147 13650 -5087 15250
rect -3508 13650 -3448 15250
rect -3428 13650 -3368 15250
rect -1789 13650 -1729 15250
rect -1709 13650 -1649 15250
rect -70 13650 -10 15250
rect 10 13650 70 15250
rect 1649 13650 1709 15250
rect 1729 13650 1789 15250
rect 3368 13650 3428 15250
rect 3448 13650 3508 15250
rect 5087 13650 5147 15250
rect 5167 13650 5227 15250
rect 6806 13650 6866 15250
rect 6886 13650 6946 15250
rect 8525 13650 8585 15250
rect 8605 13650 8665 15250
rect 10244 13650 10304 15250
rect 10324 13650 10384 15250
rect 11963 13650 12023 15250
rect 12043 13650 12103 15250
rect 13682 13650 13742 15250
rect 13762 13650 13822 15250
rect -13822 11950 -13762 13550
rect -13742 11950 -13682 13550
rect -12103 11950 -12043 13550
rect -12023 11950 -11963 13550
rect -10384 11950 -10324 13550
rect -10304 11950 -10244 13550
rect -8665 11950 -8605 13550
rect -8585 11950 -8525 13550
rect -6946 11950 -6886 13550
rect -6866 11950 -6806 13550
rect -5227 11950 -5167 13550
rect -5147 11950 -5087 13550
rect -3508 11950 -3448 13550
rect -3428 11950 -3368 13550
rect -1789 11950 -1729 13550
rect -1709 11950 -1649 13550
rect -70 11950 -10 13550
rect 10 11950 70 13550
rect 1649 11950 1709 13550
rect 1729 11950 1789 13550
rect 3368 11950 3428 13550
rect 3448 11950 3508 13550
rect 5087 11950 5147 13550
rect 5167 11950 5227 13550
rect 6806 11950 6866 13550
rect 6886 11950 6946 13550
rect 8525 11950 8585 13550
rect 8605 11950 8665 13550
rect 10244 11950 10304 13550
rect 10324 11950 10384 13550
rect 11963 11950 12023 13550
rect 12043 11950 12103 13550
rect 13682 11950 13742 13550
rect 13762 11950 13822 13550
rect -13822 10250 -13762 11850
rect -13742 10250 -13682 11850
rect -12103 10250 -12043 11850
rect -12023 10250 -11963 11850
rect -10384 10250 -10324 11850
rect -10304 10250 -10244 11850
rect -8665 10250 -8605 11850
rect -8585 10250 -8525 11850
rect -6946 10250 -6886 11850
rect -6866 10250 -6806 11850
rect -5227 10250 -5167 11850
rect -5147 10250 -5087 11850
rect -3508 10250 -3448 11850
rect -3428 10250 -3368 11850
rect -1789 10250 -1729 11850
rect -1709 10250 -1649 11850
rect -70 10250 -10 11850
rect 10 10250 70 11850
rect 1649 10250 1709 11850
rect 1729 10250 1789 11850
rect 3368 10250 3428 11850
rect 3448 10250 3508 11850
rect 5087 10250 5147 11850
rect 5167 10250 5227 11850
rect 6806 10250 6866 11850
rect 6886 10250 6946 11850
rect 8525 10250 8585 11850
rect 8605 10250 8665 11850
rect 10244 10250 10304 11850
rect 10324 10250 10384 11850
rect 11963 10250 12023 11850
rect 12043 10250 12103 11850
rect 13682 10250 13742 11850
rect 13762 10250 13822 11850
rect -13822 8550 -13762 10150
rect -13742 8550 -13682 10150
rect -12103 8550 -12043 10150
rect -12023 8550 -11963 10150
rect -10384 8550 -10324 10150
rect -10304 8550 -10244 10150
rect -8665 8550 -8605 10150
rect -8585 8550 -8525 10150
rect -6946 8550 -6886 10150
rect -6866 8550 -6806 10150
rect -5227 8550 -5167 10150
rect -5147 8550 -5087 10150
rect -3508 8550 -3448 10150
rect -3428 8550 -3368 10150
rect -1789 8550 -1729 10150
rect -1709 8550 -1649 10150
rect -70 8550 -10 10150
rect 10 8550 70 10150
rect 1649 8550 1709 10150
rect 1729 8550 1789 10150
rect 3368 8550 3428 10150
rect 3448 8550 3508 10150
rect 5087 8550 5147 10150
rect 5167 8550 5227 10150
rect 6806 8550 6866 10150
rect 6886 8550 6946 10150
rect 8525 8550 8585 10150
rect 8605 8550 8665 10150
rect 10244 8550 10304 10150
rect 10324 8550 10384 10150
rect 11963 8550 12023 10150
rect 12043 8550 12103 10150
rect 13682 8550 13742 10150
rect 13762 8550 13822 10150
rect -13822 6850 -13762 8450
rect -13742 6850 -13682 8450
rect -12103 6850 -12043 8450
rect -12023 6850 -11963 8450
rect -10384 6850 -10324 8450
rect -10304 6850 -10244 8450
rect -8665 6850 -8605 8450
rect -8585 6850 -8525 8450
rect -6946 6850 -6886 8450
rect -6866 6850 -6806 8450
rect -5227 6850 -5167 8450
rect -5147 6850 -5087 8450
rect -3508 6850 -3448 8450
rect -3428 6850 -3368 8450
rect -1789 6850 -1729 8450
rect -1709 6850 -1649 8450
rect -70 6850 -10 8450
rect 10 6850 70 8450
rect 1649 6850 1709 8450
rect 1729 6850 1789 8450
rect 3368 6850 3428 8450
rect 3448 6850 3508 8450
rect 5087 6850 5147 8450
rect 5167 6850 5227 8450
rect 6806 6850 6866 8450
rect 6886 6850 6946 8450
rect 8525 6850 8585 8450
rect 8605 6850 8665 8450
rect 10244 6850 10304 8450
rect 10324 6850 10384 8450
rect 11963 6850 12023 8450
rect 12043 6850 12103 8450
rect 13682 6850 13742 8450
rect 13762 6850 13822 8450
rect -13822 5150 -13762 6750
rect -13742 5150 -13682 6750
rect -12103 5150 -12043 6750
rect -12023 5150 -11963 6750
rect -10384 5150 -10324 6750
rect -10304 5150 -10244 6750
rect -8665 5150 -8605 6750
rect -8585 5150 -8525 6750
rect -6946 5150 -6886 6750
rect -6866 5150 -6806 6750
rect -5227 5150 -5167 6750
rect -5147 5150 -5087 6750
rect -3508 5150 -3448 6750
rect -3428 5150 -3368 6750
rect -1789 5150 -1729 6750
rect -1709 5150 -1649 6750
rect -70 5150 -10 6750
rect 10 5150 70 6750
rect 1649 5150 1709 6750
rect 1729 5150 1789 6750
rect 3368 5150 3428 6750
rect 3448 5150 3508 6750
rect 5087 5150 5147 6750
rect 5167 5150 5227 6750
rect 6806 5150 6866 6750
rect 6886 5150 6946 6750
rect 8525 5150 8585 6750
rect 8605 5150 8665 6750
rect 10244 5150 10304 6750
rect 10324 5150 10384 6750
rect 11963 5150 12023 6750
rect 12043 5150 12103 6750
rect 13682 5150 13742 6750
rect 13762 5150 13822 6750
rect -13822 3450 -13762 5050
rect -13742 3450 -13682 5050
rect -12103 3450 -12043 5050
rect -12023 3450 -11963 5050
rect -10384 3450 -10324 5050
rect -10304 3450 -10244 5050
rect -8665 3450 -8605 5050
rect -8585 3450 -8525 5050
rect -6946 3450 -6886 5050
rect -6866 3450 -6806 5050
rect -5227 3450 -5167 5050
rect -5147 3450 -5087 5050
rect -3508 3450 -3448 5050
rect -3428 3450 -3368 5050
rect -1789 3450 -1729 5050
rect -1709 3450 -1649 5050
rect -70 3450 -10 5050
rect 10 3450 70 5050
rect 1649 3450 1709 5050
rect 1729 3450 1789 5050
rect 3368 3450 3428 5050
rect 3448 3450 3508 5050
rect 5087 3450 5147 5050
rect 5167 3450 5227 5050
rect 6806 3450 6866 5050
rect 6886 3450 6946 5050
rect 8525 3450 8585 5050
rect 8605 3450 8665 5050
rect 10244 3450 10304 5050
rect 10324 3450 10384 5050
rect 11963 3450 12023 5050
rect 12043 3450 12103 5050
rect 13682 3450 13742 5050
rect 13762 3450 13822 5050
rect -13822 1750 -13762 3350
rect -13742 1750 -13682 3350
rect -12103 1750 -12043 3350
rect -12023 1750 -11963 3350
rect -10384 1750 -10324 3350
rect -10304 1750 -10244 3350
rect -8665 1750 -8605 3350
rect -8585 1750 -8525 3350
rect -6946 1750 -6886 3350
rect -6866 1750 -6806 3350
rect -5227 1750 -5167 3350
rect -5147 1750 -5087 3350
rect -3508 1750 -3448 3350
rect -3428 1750 -3368 3350
rect -1789 1750 -1729 3350
rect -1709 1750 -1649 3350
rect -70 1750 -10 3350
rect 10 1750 70 3350
rect 1649 1750 1709 3350
rect 1729 1750 1789 3350
rect 3368 1750 3428 3350
rect 3448 1750 3508 3350
rect 5087 1750 5147 3350
rect 5167 1750 5227 3350
rect 6806 1750 6866 3350
rect 6886 1750 6946 3350
rect 8525 1750 8585 3350
rect 8605 1750 8665 3350
rect 10244 1750 10304 3350
rect 10324 1750 10384 3350
rect 11963 1750 12023 3350
rect 12043 1750 12103 3350
rect 13682 1750 13742 3350
rect 13762 1750 13822 3350
rect -13822 50 -13762 1650
rect -13742 50 -13682 1650
rect -12103 50 -12043 1650
rect -12023 50 -11963 1650
rect -10384 50 -10324 1650
rect -10304 50 -10244 1650
rect -8665 50 -8605 1650
rect -8585 50 -8525 1650
rect -6946 50 -6886 1650
rect -6866 50 -6806 1650
rect -5227 50 -5167 1650
rect -5147 50 -5087 1650
rect -3508 50 -3448 1650
rect -3428 50 -3368 1650
rect -1789 50 -1729 1650
rect -1709 50 -1649 1650
rect -70 50 -10 1650
rect 10 50 70 1650
rect 1649 50 1709 1650
rect 1729 50 1789 1650
rect 3368 50 3428 1650
rect 3448 50 3508 1650
rect 5087 50 5147 1650
rect 5167 50 5227 1650
rect 6806 50 6866 1650
rect 6886 50 6946 1650
rect 8525 50 8585 1650
rect 8605 50 8665 1650
rect 10244 50 10304 1650
rect 10324 50 10384 1650
rect 11963 50 12023 1650
rect 12043 50 12103 1650
rect 13682 50 13742 1650
rect 13762 50 13822 1650
rect -13822 -1650 -13762 -50
rect -13742 -1650 -13682 -50
rect -12103 -1650 -12043 -50
rect -12023 -1650 -11963 -50
rect -10384 -1650 -10324 -50
rect -10304 -1650 -10244 -50
rect -8665 -1650 -8605 -50
rect -8585 -1650 -8525 -50
rect -6946 -1650 -6886 -50
rect -6866 -1650 -6806 -50
rect -5227 -1650 -5167 -50
rect -5147 -1650 -5087 -50
rect -3508 -1650 -3448 -50
rect -3428 -1650 -3368 -50
rect -1789 -1650 -1729 -50
rect -1709 -1650 -1649 -50
rect -70 -1650 -10 -50
rect 10 -1650 70 -50
rect 1649 -1650 1709 -50
rect 1729 -1650 1789 -50
rect 3368 -1650 3428 -50
rect 3448 -1650 3508 -50
rect 5087 -1650 5147 -50
rect 5167 -1650 5227 -50
rect 6806 -1650 6866 -50
rect 6886 -1650 6946 -50
rect 8525 -1650 8585 -50
rect 8605 -1650 8665 -50
rect 10244 -1650 10304 -50
rect 10324 -1650 10384 -50
rect 11963 -1650 12023 -50
rect 12043 -1650 12103 -50
rect 13682 -1650 13742 -50
rect 13762 -1650 13822 -50
rect -13822 -3350 -13762 -1750
rect -13742 -3350 -13682 -1750
rect -12103 -3350 -12043 -1750
rect -12023 -3350 -11963 -1750
rect -10384 -3350 -10324 -1750
rect -10304 -3350 -10244 -1750
rect -8665 -3350 -8605 -1750
rect -8585 -3350 -8525 -1750
rect -6946 -3350 -6886 -1750
rect -6866 -3350 -6806 -1750
rect -5227 -3350 -5167 -1750
rect -5147 -3350 -5087 -1750
rect -3508 -3350 -3448 -1750
rect -3428 -3350 -3368 -1750
rect -1789 -3350 -1729 -1750
rect -1709 -3350 -1649 -1750
rect -70 -3350 -10 -1750
rect 10 -3350 70 -1750
rect 1649 -3350 1709 -1750
rect 1729 -3350 1789 -1750
rect 3368 -3350 3428 -1750
rect 3448 -3350 3508 -1750
rect 5087 -3350 5147 -1750
rect 5167 -3350 5227 -1750
rect 6806 -3350 6866 -1750
rect 6886 -3350 6946 -1750
rect 8525 -3350 8585 -1750
rect 8605 -3350 8665 -1750
rect 10244 -3350 10304 -1750
rect 10324 -3350 10384 -1750
rect 11963 -3350 12023 -1750
rect 12043 -3350 12103 -1750
rect 13682 -3350 13742 -1750
rect 13762 -3350 13822 -1750
rect -13822 -5050 -13762 -3450
rect -13742 -5050 -13682 -3450
rect -12103 -5050 -12043 -3450
rect -12023 -5050 -11963 -3450
rect -10384 -5050 -10324 -3450
rect -10304 -5050 -10244 -3450
rect -8665 -5050 -8605 -3450
rect -8585 -5050 -8525 -3450
rect -6946 -5050 -6886 -3450
rect -6866 -5050 -6806 -3450
rect -5227 -5050 -5167 -3450
rect -5147 -5050 -5087 -3450
rect -3508 -5050 -3448 -3450
rect -3428 -5050 -3368 -3450
rect -1789 -5050 -1729 -3450
rect -1709 -5050 -1649 -3450
rect -70 -5050 -10 -3450
rect 10 -5050 70 -3450
rect 1649 -5050 1709 -3450
rect 1729 -5050 1789 -3450
rect 3368 -5050 3428 -3450
rect 3448 -5050 3508 -3450
rect 5087 -5050 5147 -3450
rect 5167 -5050 5227 -3450
rect 6806 -5050 6866 -3450
rect 6886 -5050 6946 -3450
rect 8525 -5050 8585 -3450
rect 8605 -5050 8665 -3450
rect 10244 -5050 10304 -3450
rect 10324 -5050 10384 -3450
rect 11963 -5050 12023 -3450
rect 12043 -5050 12103 -3450
rect 13682 -5050 13742 -3450
rect 13762 -5050 13822 -3450
rect -13822 -6750 -13762 -5150
rect -13742 -6750 -13682 -5150
rect -12103 -6750 -12043 -5150
rect -12023 -6750 -11963 -5150
rect -10384 -6750 -10324 -5150
rect -10304 -6750 -10244 -5150
rect -8665 -6750 -8605 -5150
rect -8585 -6750 -8525 -5150
rect -6946 -6750 -6886 -5150
rect -6866 -6750 -6806 -5150
rect -5227 -6750 -5167 -5150
rect -5147 -6750 -5087 -5150
rect -3508 -6750 -3448 -5150
rect -3428 -6750 -3368 -5150
rect -1789 -6750 -1729 -5150
rect -1709 -6750 -1649 -5150
rect -70 -6750 -10 -5150
rect 10 -6750 70 -5150
rect 1649 -6750 1709 -5150
rect 1729 -6750 1789 -5150
rect 3368 -6750 3428 -5150
rect 3448 -6750 3508 -5150
rect 5087 -6750 5147 -5150
rect 5167 -6750 5227 -5150
rect 6806 -6750 6866 -5150
rect 6886 -6750 6946 -5150
rect 8525 -6750 8585 -5150
rect 8605 -6750 8665 -5150
rect 10244 -6750 10304 -5150
rect 10324 -6750 10384 -5150
rect 11963 -6750 12023 -5150
rect 12043 -6750 12103 -5150
rect 13682 -6750 13742 -5150
rect 13762 -6750 13822 -5150
rect -13822 -8450 -13762 -6850
rect -13742 -8450 -13682 -6850
rect -12103 -8450 -12043 -6850
rect -12023 -8450 -11963 -6850
rect -10384 -8450 -10324 -6850
rect -10304 -8450 -10244 -6850
rect -8665 -8450 -8605 -6850
rect -8585 -8450 -8525 -6850
rect -6946 -8450 -6886 -6850
rect -6866 -8450 -6806 -6850
rect -5227 -8450 -5167 -6850
rect -5147 -8450 -5087 -6850
rect -3508 -8450 -3448 -6850
rect -3428 -8450 -3368 -6850
rect -1789 -8450 -1729 -6850
rect -1709 -8450 -1649 -6850
rect -70 -8450 -10 -6850
rect 10 -8450 70 -6850
rect 1649 -8450 1709 -6850
rect 1729 -8450 1789 -6850
rect 3368 -8450 3428 -6850
rect 3448 -8450 3508 -6850
rect 5087 -8450 5147 -6850
rect 5167 -8450 5227 -6850
rect 6806 -8450 6866 -6850
rect 6886 -8450 6946 -6850
rect 8525 -8450 8585 -6850
rect 8605 -8450 8665 -6850
rect 10244 -8450 10304 -6850
rect 10324 -8450 10384 -6850
rect 11963 -8450 12023 -6850
rect 12043 -8450 12103 -6850
rect 13682 -8450 13742 -6850
rect 13762 -8450 13822 -6850
rect -13822 -10150 -13762 -8550
rect -13742 -10150 -13682 -8550
rect -12103 -10150 -12043 -8550
rect -12023 -10150 -11963 -8550
rect -10384 -10150 -10324 -8550
rect -10304 -10150 -10244 -8550
rect -8665 -10150 -8605 -8550
rect -8585 -10150 -8525 -8550
rect -6946 -10150 -6886 -8550
rect -6866 -10150 -6806 -8550
rect -5227 -10150 -5167 -8550
rect -5147 -10150 -5087 -8550
rect -3508 -10150 -3448 -8550
rect -3428 -10150 -3368 -8550
rect -1789 -10150 -1729 -8550
rect -1709 -10150 -1649 -8550
rect -70 -10150 -10 -8550
rect 10 -10150 70 -8550
rect 1649 -10150 1709 -8550
rect 1729 -10150 1789 -8550
rect 3368 -10150 3428 -8550
rect 3448 -10150 3508 -8550
rect 5087 -10150 5147 -8550
rect 5167 -10150 5227 -8550
rect 6806 -10150 6866 -8550
rect 6886 -10150 6946 -8550
rect 8525 -10150 8585 -8550
rect 8605 -10150 8665 -8550
rect 10244 -10150 10304 -8550
rect 10324 -10150 10384 -8550
rect 11963 -10150 12023 -8550
rect 12043 -10150 12103 -8550
rect 13682 -10150 13742 -8550
rect 13762 -10150 13822 -8550
rect -13822 -11850 -13762 -10250
rect -13742 -11850 -13682 -10250
rect -12103 -11850 -12043 -10250
rect -12023 -11850 -11963 -10250
rect -10384 -11850 -10324 -10250
rect -10304 -11850 -10244 -10250
rect -8665 -11850 -8605 -10250
rect -8585 -11850 -8525 -10250
rect -6946 -11850 -6886 -10250
rect -6866 -11850 -6806 -10250
rect -5227 -11850 -5167 -10250
rect -5147 -11850 -5087 -10250
rect -3508 -11850 -3448 -10250
rect -3428 -11850 -3368 -10250
rect -1789 -11850 -1729 -10250
rect -1709 -11850 -1649 -10250
rect -70 -11850 -10 -10250
rect 10 -11850 70 -10250
rect 1649 -11850 1709 -10250
rect 1729 -11850 1789 -10250
rect 3368 -11850 3428 -10250
rect 3448 -11850 3508 -10250
rect 5087 -11850 5147 -10250
rect 5167 -11850 5227 -10250
rect 6806 -11850 6866 -10250
rect 6886 -11850 6946 -10250
rect 8525 -11850 8585 -10250
rect 8605 -11850 8665 -10250
rect 10244 -11850 10304 -10250
rect 10324 -11850 10384 -10250
rect 11963 -11850 12023 -10250
rect 12043 -11850 12103 -10250
rect 13682 -11850 13742 -10250
rect 13762 -11850 13822 -10250
rect -13822 -13550 -13762 -11950
rect -13742 -13550 -13682 -11950
rect -12103 -13550 -12043 -11950
rect -12023 -13550 -11963 -11950
rect -10384 -13550 -10324 -11950
rect -10304 -13550 -10244 -11950
rect -8665 -13550 -8605 -11950
rect -8585 -13550 -8525 -11950
rect -6946 -13550 -6886 -11950
rect -6866 -13550 -6806 -11950
rect -5227 -13550 -5167 -11950
rect -5147 -13550 -5087 -11950
rect -3508 -13550 -3448 -11950
rect -3428 -13550 -3368 -11950
rect -1789 -13550 -1729 -11950
rect -1709 -13550 -1649 -11950
rect -70 -13550 -10 -11950
rect 10 -13550 70 -11950
rect 1649 -13550 1709 -11950
rect 1729 -13550 1789 -11950
rect 3368 -13550 3428 -11950
rect 3448 -13550 3508 -11950
rect 5087 -13550 5147 -11950
rect 5167 -13550 5227 -11950
rect 6806 -13550 6866 -11950
rect 6886 -13550 6946 -11950
rect 8525 -13550 8585 -11950
rect 8605 -13550 8665 -11950
rect 10244 -13550 10304 -11950
rect 10324 -13550 10384 -11950
rect 11963 -13550 12023 -11950
rect 12043 -13550 12103 -11950
rect 13682 -13550 13742 -11950
rect 13762 -13550 13822 -11950
rect -13822 -15250 -13762 -13650
rect -13742 -15250 -13682 -13650
rect -12103 -15250 -12043 -13650
rect -12023 -15250 -11963 -13650
rect -10384 -15250 -10324 -13650
rect -10304 -15250 -10244 -13650
rect -8665 -15250 -8605 -13650
rect -8585 -15250 -8525 -13650
rect -6946 -15250 -6886 -13650
rect -6866 -15250 -6806 -13650
rect -5227 -15250 -5167 -13650
rect -5147 -15250 -5087 -13650
rect -3508 -15250 -3448 -13650
rect -3428 -15250 -3368 -13650
rect -1789 -15250 -1729 -13650
rect -1709 -15250 -1649 -13650
rect -70 -15250 -10 -13650
rect 10 -15250 70 -13650
rect 1649 -15250 1709 -13650
rect 1729 -15250 1789 -13650
rect 3368 -15250 3428 -13650
rect 3448 -15250 3508 -13650
rect 5087 -15250 5147 -13650
rect 5167 -15250 5227 -13650
rect 6806 -15250 6866 -13650
rect 6886 -15250 6946 -13650
rect 8525 -15250 8585 -13650
rect 8605 -15250 8665 -13650
rect 10244 -15250 10304 -13650
rect 10324 -15250 10384 -13650
rect 11963 -15250 12023 -13650
rect 12043 -15250 12103 -13650
rect 13682 -15250 13742 -13650
rect 13762 -15250 13822 -13650
<< metal3 >>
rect -15461 15222 -13762 15250
rect -15461 13678 -13846 15222
rect -13782 13678 -13762 15222
rect -15461 13650 -13762 13678
rect -13742 15222 -12043 15250
rect -13742 13678 -12127 15222
rect -12063 13678 -12043 15222
rect -13742 13650 -12043 13678
rect -12023 15222 -10324 15250
rect -12023 13678 -10408 15222
rect -10344 13678 -10324 15222
rect -12023 13650 -10324 13678
rect -10304 15222 -8605 15250
rect -10304 13678 -8689 15222
rect -8625 13678 -8605 15222
rect -10304 13650 -8605 13678
rect -8585 15222 -6886 15250
rect -8585 13678 -6970 15222
rect -6906 13678 -6886 15222
rect -8585 13650 -6886 13678
rect -6866 15222 -5167 15250
rect -6866 13678 -5251 15222
rect -5187 13678 -5167 15222
rect -6866 13650 -5167 13678
rect -5147 15222 -3448 15250
rect -5147 13678 -3532 15222
rect -3468 13678 -3448 15222
rect -5147 13650 -3448 13678
rect -3428 15222 -1729 15250
rect -3428 13678 -1813 15222
rect -1749 13678 -1729 15222
rect -3428 13650 -1729 13678
rect -1709 15222 -10 15250
rect -1709 13678 -94 15222
rect -30 13678 -10 15222
rect -1709 13650 -10 13678
rect 10 15222 1709 15250
rect 10 13678 1625 15222
rect 1689 13678 1709 15222
rect 10 13650 1709 13678
rect 1729 15222 3428 15250
rect 1729 13678 3344 15222
rect 3408 13678 3428 15222
rect 1729 13650 3428 13678
rect 3448 15222 5147 15250
rect 3448 13678 5063 15222
rect 5127 13678 5147 15222
rect 3448 13650 5147 13678
rect 5167 15222 6866 15250
rect 5167 13678 6782 15222
rect 6846 13678 6866 15222
rect 5167 13650 6866 13678
rect 6886 15222 8585 15250
rect 6886 13678 8501 15222
rect 8565 13678 8585 15222
rect 6886 13650 8585 13678
rect 8605 15222 10304 15250
rect 8605 13678 10220 15222
rect 10284 13678 10304 15222
rect 8605 13650 10304 13678
rect 10324 15222 12023 15250
rect 10324 13678 11939 15222
rect 12003 13678 12023 15222
rect 10324 13650 12023 13678
rect 12043 15222 13742 15250
rect 12043 13678 13658 15222
rect 13722 13678 13742 15222
rect 12043 13650 13742 13678
rect 13762 15222 15461 15250
rect 13762 13678 15377 15222
rect 15441 13678 15461 15222
rect 13762 13650 15461 13678
rect -15461 13522 -13762 13550
rect -15461 11978 -13846 13522
rect -13782 11978 -13762 13522
rect -15461 11950 -13762 11978
rect -13742 13522 -12043 13550
rect -13742 11978 -12127 13522
rect -12063 11978 -12043 13522
rect -13742 11950 -12043 11978
rect -12023 13522 -10324 13550
rect -12023 11978 -10408 13522
rect -10344 11978 -10324 13522
rect -12023 11950 -10324 11978
rect -10304 13522 -8605 13550
rect -10304 11978 -8689 13522
rect -8625 11978 -8605 13522
rect -10304 11950 -8605 11978
rect -8585 13522 -6886 13550
rect -8585 11978 -6970 13522
rect -6906 11978 -6886 13522
rect -8585 11950 -6886 11978
rect -6866 13522 -5167 13550
rect -6866 11978 -5251 13522
rect -5187 11978 -5167 13522
rect -6866 11950 -5167 11978
rect -5147 13522 -3448 13550
rect -5147 11978 -3532 13522
rect -3468 11978 -3448 13522
rect -5147 11950 -3448 11978
rect -3428 13522 -1729 13550
rect -3428 11978 -1813 13522
rect -1749 11978 -1729 13522
rect -3428 11950 -1729 11978
rect -1709 13522 -10 13550
rect -1709 11978 -94 13522
rect -30 11978 -10 13522
rect -1709 11950 -10 11978
rect 10 13522 1709 13550
rect 10 11978 1625 13522
rect 1689 11978 1709 13522
rect 10 11950 1709 11978
rect 1729 13522 3428 13550
rect 1729 11978 3344 13522
rect 3408 11978 3428 13522
rect 1729 11950 3428 11978
rect 3448 13522 5147 13550
rect 3448 11978 5063 13522
rect 5127 11978 5147 13522
rect 3448 11950 5147 11978
rect 5167 13522 6866 13550
rect 5167 11978 6782 13522
rect 6846 11978 6866 13522
rect 5167 11950 6866 11978
rect 6886 13522 8585 13550
rect 6886 11978 8501 13522
rect 8565 11978 8585 13522
rect 6886 11950 8585 11978
rect 8605 13522 10304 13550
rect 8605 11978 10220 13522
rect 10284 11978 10304 13522
rect 8605 11950 10304 11978
rect 10324 13522 12023 13550
rect 10324 11978 11939 13522
rect 12003 11978 12023 13522
rect 10324 11950 12023 11978
rect 12043 13522 13742 13550
rect 12043 11978 13658 13522
rect 13722 11978 13742 13522
rect 12043 11950 13742 11978
rect 13762 13522 15461 13550
rect 13762 11978 15377 13522
rect 15441 11978 15461 13522
rect 13762 11950 15461 11978
rect -15461 11822 -13762 11850
rect -15461 10278 -13846 11822
rect -13782 10278 -13762 11822
rect -15461 10250 -13762 10278
rect -13742 11822 -12043 11850
rect -13742 10278 -12127 11822
rect -12063 10278 -12043 11822
rect -13742 10250 -12043 10278
rect -12023 11822 -10324 11850
rect -12023 10278 -10408 11822
rect -10344 10278 -10324 11822
rect -12023 10250 -10324 10278
rect -10304 11822 -8605 11850
rect -10304 10278 -8689 11822
rect -8625 10278 -8605 11822
rect -10304 10250 -8605 10278
rect -8585 11822 -6886 11850
rect -8585 10278 -6970 11822
rect -6906 10278 -6886 11822
rect -8585 10250 -6886 10278
rect -6866 11822 -5167 11850
rect -6866 10278 -5251 11822
rect -5187 10278 -5167 11822
rect -6866 10250 -5167 10278
rect -5147 11822 -3448 11850
rect -5147 10278 -3532 11822
rect -3468 10278 -3448 11822
rect -5147 10250 -3448 10278
rect -3428 11822 -1729 11850
rect -3428 10278 -1813 11822
rect -1749 10278 -1729 11822
rect -3428 10250 -1729 10278
rect -1709 11822 -10 11850
rect -1709 10278 -94 11822
rect -30 10278 -10 11822
rect -1709 10250 -10 10278
rect 10 11822 1709 11850
rect 10 10278 1625 11822
rect 1689 10278 1709 11822
rect 10 10250 1709 10278
rect 1729 11822 3428 11850
rect 1729 10278 3344 11822
rect 3408 10278 3428 11822
rect 1729 10250 3428 10278
rect 3448 11822 5147 11850
rect 3448 10278 5063 11822
rect 5127 10278 5147 11822
rect 3448 10250 5147 10278
rect 5167 11822 6866 11850
rect 5167 10278 6782 11822
rect 6846 10278 6866 11822
rect 5167 10250 6866 10278
rect 6886 11822 8585 11850
rect 6886 10278 8501 11822
rect 8565 10278 8585 11822
rect 6886 10250 8585 10278
rect 8605 11822 10304 11850
rect 8605 10278 10220 11822
rect 10284 10278 10304 11822
rect 8605 10250 10304 10278
rect 10324 11822 12023 11850
rect 10324 10278 11939 11822
rect 12003 10278 12023 11822
rect 10324 10250 12023 10278
rect 12043 11822 13742 11850
rect 12043 10278 13658 11822
rect 13722 10278 13742 11822
rect 12043 10250 13742 10278
rect 13762 11822 15461 11850
rect 13762 10278 15377 11822
rect 15441 10278 15461 11822
rect 13762 10250 15461 10278
rect -15461 10122 -13762 10150
rect -15461 8578 -13846 10122
rect -13782 8578 -13762 10122
rect -15461 8550 -13762 8578
rect -13742 10122 -12043 10150
rect -13742 8578 -12127 10122
rect -12063 8578 -12043 10122
rect -13742 8550 -12043 8578
rect -12023 10122 -10324 10150
rect -12023 8578 -10408 10122
rect -10344 8578 -10324 10122
rect -12023 8550 -10324 8578
rect -10304 10122 -8605 10150
rect -10304 8578 -8689 10122
rect -8625 8578 -8605 10122
rect -10304 8550 -8605 8578
rect -8585 10122 -6886 10150
rect -8585 8578 -6970 10122
rect -6906 8578 -6886 10122
rect -8585 8550 -6886 8578
rect -6866 10122 -5167 10150
rect -6866 8578 -5251 10122
rect -5187 8578 -5167 10122
rect -6866 8550 -5167 8578
rect -5147 10122 -3448 10150
rect -5147 8578 -3532 10122
rect -3468 8578 -3448 10122
rect -5147 8550 -3448 8578
rect -3428 10122 -1729 10150
rect -3428 8578 -1813 10122
rect -1749 8578 -1729 10122
rect -3428 8550 -1729 8578
rect -1709 10122 -10 10150
rect -1709 8578 -94 10122
rect -30 8578 -10 10122
rect -1709 8550 -10 8578
rect 10 10122 1709 10150
rect 10 8578 1625 10122
rect 1689 8578 1709 10122
rect 10 8550 1709 8578
rect 1729 10122 3428 10150
rect 1729 8578 3344 10122
rect 3408 8578 3428 10122
rect 1729 8550 3428 8578
rect 3448 10122 5147 10150
rect 3448 8578 5063 10122
rect 5127 8578 5147 10122
rect 3448 8550 5147 8578
rect 5167 10122 6866 10150
rect 5167 8578 6782 10122
rect 6846 8578 6866 10122
rect 5167 8550 6866 8578
rect 6886 10122 8585 10150
rect 6886 8578 8501 10122
rect 8565 8578 8585 10122
rect 6886 8550 8585 8578
rect 8605 10122 10304 10150
rect 8605 8578 10220 10122
rect 10284 8578 10304 10122
rect 8605 8550 10304 8578
rect 10324 10122 12023 10150
rect 10324 8578 11939 10122
rect 12003 8578 12023 10122
rect 10324 8550 12023 8578
rect 12043 10122 13742 10150
rect 12043 8578 13658 10122
rect 13722 8578 13742 10122
rect 12043 8550 13742 8578
rect 13762 10122 15461 10150
rect 13762 8578 15377 10122
rect 15441 8578 15461 10122
rect 13762 8550 15461 8578
rect -15461 8422 -13762 8450
rect -15461 6878 -13846 8422
rect -13782 6878 -13762 8422
rect -15461 6850 -13762 6878
rect -13742 8422 -12043 8450
rect -13742 6878 -12127 8422
rect -12063 6878 -12043 8422
rect -13742 6850 -12043 6878
rect -12023 8422 -10324 8450
rect -12023 6878 -10408 8422
rect -10344 6878 -10324 8422
rect -12023 6850 -10324 6878
rect -10304 8422 -8605 8450
rect -10304 6878 -8689 8422
rect -8625 6878 -8605 8422
rect -10304 6850 -8605 6878
rect -8585 8422 -6886 8450
rect -8585 6878 -6970 8422
rect -6906 6878 -6886 8422
rect -8585 6850 -6886 6878
rect -6866 8422 -5167 8450
rect -6866 6878 -5251 8422
rect -5187 6878 -5167 8422
rect -6866 6850 -5167 6878
rect -5147 8422 -3448 8450
rect -5147 6878 -3532 8422
rect -3468 6878 -3448 8422
rect -5147 6850 -3448 6878
rect -3428 8422 -1729 8450
rect -3428 6878 -1813 8422
rect -1749 6878 -1729 8422
rect -3428 6850 -1729 6878
rect -1709 8422 -10 8450
rect -1709 6878 -94 8422
rect -30 6878 -10 8422
rect -1709 6850 -10 6878
rect 10 8422 1709 8450
rect 10 6878 1625 8422
rect 1689 6878 1709 8422
rect 10 6850 1709 6878
rect 1729 8422 3428 8450
rect 1729 6878 3344 8422
rect 3408 6878 3428 8422
rect 1729 6850 3428 6878
rect 3448 8422 5147 8450
rect 3448 6878 5063 8422
rect 5127 6878 5147 8422
rect 3448 6850 5147 6878
rect 5167 8422 6866 8450
rect 5167 6878 6782 8422
rect 6846 6878 6866 8422
rect 5167 6850 6866 6878
rect 6886 8422 8585 8450
rect 6886 6878 8501 8422
rect 8565 6878 8585 8422
rect 6886 6850 8585 6878
rect 8605 8422 10304 8450
rect 8605 6878 10220 8422
rect 10284 6878 10304 8422
rect 8605 6850 10304 6878
rect 10324 8422 12023 8450
rect 10324 6878 11939 8422
rect 12003 6878 12023 8422
rect 10324 6850 12023 6878
rect 12043 8422 13742 8450
rect 12043 6878 13658 8422
rect 13722 6878 13742 8422
rect 12043 6850 13742 6878
rect 13762 8422 15461 8450
rect 13762 6878 15377 8422
rect 15441 6878 15461 8422
rect 13762 6850 15461 6878
rect -15461 6722 -13762 6750
rect -15461 5178 -13846 6722
rect -13782 5178 -13762 6722
rect -15461 5150 -13762 5178
rect -13742 6722 -12043 6750
rect -13742 5178 -12127 6722
rect -12063 5178 -12043 6722
rect -13742 5150 -12043 5178
rect -12023 6722 -10324 6750
rect -12023 5178 -10408 6722
rect -10344 5178 -10324 6722
rect -12023 5150 -10324 5178
rect -10304 6722 -8605 6750
rect -10304 5178 -8689 6722
rect -8625 5178 -8605 6722
rect -10304 5150 -8605 5178
rect -8585 6722 -6886 6750
rect -8585 5178 -6970 6722
rect -6906 5178 -6886 6722
rect -8585 5150 -6886 5178
rect -6866 6722 -5167 6750
rect -6866 5178 -5251 6722
rect -5187 5178 -5167 6722
rect -6866 5150 -5167 5178
rect -5147 6722 -3448 6750
rect -5147 5178 -3532 6722
rect -3468 5178 -3448 6722
rect -5147 5150 -3448 5178
rect -3428 6722 -1729 6750
rect -3428 5178 -1813 6722
rect -1749 5178 -1729 6722
rect -3428 5150 -1729 5178
rect -1709 6722 -10 6750
rect -1709 5178 -94 6722
rect -30 5178 -10 6722
rect -1709 5150 -10 5178
rect 10 6722 1709 6750
rect 10 5178 1625 6722
rect 1689 5178 1709 6722
rect 10 5150 1709 5178
rect 1729 6722 3428 6750
rect 1729 5178 3344 6722
rect 3408 5178 3428 6722
rect 1729 5150 3428 5178
rect 3448 6722 5147 6750
rect 3448 5178 5063 6722
rect 5127 5178 5147 6722
rect 3448 5150 5147 5178
rect 5167 6722 6866 6750
rect 5167 5178 6782 6722
rect 6846 5178 6866 6722
rect 5167 5150 6866 5178
rect 6886 6722 8585 6750
rect 6886 5178 8501 6722
rect 8565 5178 8585 6722
rect 6886 5150 8585 5178
rect 8605 6722 10304 6750
rect 8605 5178 10220 6722
rect 10284 5178 10304 6722
rect 8605 5150 10304 5178
rect 10324 6722 12023 6750
rect 10324 5178 11939 6722
rect 12003 5178 12023 6722
rect 10324 5150 12023 5178
rect 12043 6722 13742 6750
rect 12043 5178 13658 6722
rect 13722 5178 13742 6722
rect 12043 5150 13742 5178
rect 13762 6722 15461 6750
rect 13762 5178 15377 6722
rect 15441 5178 15461 6722
rect 13762 5150 15461 5178
rect -15461 5022 -13762 5050
rect -15461 3478 -13846 5022
rect -13782 3478 -13762 5022
rect -15461 3450 -13762 3478
rect -13742 5022 -12043 5050
rect -13742 3478 -12127 5022
rect -12063 3478 -12043 5022
rect -13742 3450 -12043 3478
rect -12023 5022 -10324 5050
rect -12023 3478 -10408 5022
rect -10344 3478 -10324 5022
rect -12023 3450 -10324 3478
rect -10304 5022 -8605 5050
rect -10304 3478 -8689 5022
rect -8625 3478 -8605 5022
rect -10304 3450 -8605 3478
rect -8585 5022 -6886 5050
rect -8585 3478 -6970 5022
rect -6906 3478 -6886 5022
rect -8585 3450 -6886 3478
rect -6866 5022 -5167 5050
rect -6866 3478 -5251 5022
rect -5187 3478 -5167 5022
rect -6866 3450 -5167 3478
rect -5147 5022 -3448 5050
rect -5147 3478 -3532 5022
rect -3468 3478 -3448 5022
rect -5147 3450 -3448 3478
rect -3428 5022 -1729 5050
rect -3428 3478 -1813 5022
rect -1749 3478 -1729 5022
rect -3428 3450 -1729 3478
rect -1709 5022 -10 5050
rect -1709 3478 -94 5022
rect -30 3478 -10 5022
rect -1709 3450 -10 3478
rect 10 5022 1709 5050
rect 10 3478 1625 5022
rect 1689 3478 1709 5022
rect 10 3450 1709 3478
rect 1729 5022 3428 5050
rect 1729 3478 3344 5022
rect 3408 3478 3428 5022
rect 1729 3450 3428 3478
rect 3448 5022 5147 5050
rect 3448 3478 5063 5022
rect 5127 3478 5147 5022
rect 3448 3450 5147 3478
rect 5167 5022 6866 5050
rect 5167 3478 6782 5022
rect 6846 3478 6866 5022
rect 5167 3450 6866 3478
rect 6886 5022 8585 5050
rect 6886 3478 8501 5022
rect 8565 3478 8585 5022
rect 6886 3450 8585 3478
rect 8605 5022 10304 5050
rect 8605 3478 10220 5022
rect 10284 3478 10304 5022
rect 8605 3450 10304 3478
rect 10324 5022 12023 5050
rect 10324 3478 11939 5022
rect 12003 3478 12023 5022
rect 10324 3450 12023 3478
rect 12043 5022 13742 5050
rect 12043 3478 13658 5022
rect 13722 3478 13742 5022
rect 12043 3450 13742 3478
rect 13762 5022 15461 5050
rect 13762 3478 15377 5022
rect 15441 3478 15461 5022
rect 13762 3450 15461 3478
rect -15461 3322 -13762 3350
rect -15461 1778 -13846 3322
rect -13782 1778 -13762 3322
rect -15461 1750 -13762 1778
rect -13742 3322 -12043 3350
rect -13742 1778 -12127 3322
rect -12063 1778 -12043 3322
rect -13742 1750 -12043 1778
rect -12023 3322 -10324 3350
rect -12023 1778 -10408 3322
rect -10344 1778 -10324 3322
rect -12023 1750 -10324 1778
rect -10304 3322 -8605 3350
rect -10304 1778 -8689 3322
rect -8625 1778 -8605 3322
rect -10304 1750 -8605 1778
rect -8585 3322 -6886 3350
rect -8585 1778 -6970 3322
rect -6906 1778 -6886 3322
rect -8585 1750 -6886 1778
rect -6866 3322 -5167 3350
rect -6866 1778 -5251 3322
rect -5187 1778 -5167 3322
rect -6866 1750 -5167 1778
rect -5147 3322 -3448 3350
rect -5147 1778 -3532 3322
rect -3468 1778 -3448 3322
rect -5147 1750 -3448 1778
rect -3428 3322 -1729 3350
rect -3428 1778 -1813 3322
rect -1749 1778 -1729 3322
rect -3428 1750 -1729 1778
rect -1709 3322 -10 3350
rect -1709 1778 -94 3322
rect -30 1778 -10 3322
rect -1709 1750 -10 1778
rect 10 3322 1709 3350
rect 10 1778 1625 3322
rect 1689 1778 1709 3322
rect 10 1750 1709 1778
rect 1729 3322 3428 3350
rect 1729 1778 3344 3322
rect 3408 1778 3428 3322
rect 1729 1750 3428 1778
rect 3448 3322 5147 3350
rect 3448 1778 5063 3322
rect 5127 1778 5147 3322
rect 3448 1750 5147 1778
rect 5167 3322 6866 3350
rect 5167 1778 6782 3322
rect 6846 1778 6866 3322
rect 5167 1750 6866 1778
rect 6886 3322 8585 3350
rect 6886 1778 8501 3322
rect 8565 1778 8585 3322
rect 6886 1750 8585 1778
rect 8605 3322 10304 3350
rect 8605 1778 10220 3322
rect 10284 1778 10304 3322
rect 8605 1750 10304 1778
rect 10324 3322 12023 3350
rect 10324 1778 11939 3322
rect 12003 1778 12023 3322
rect 10324 1750 12023 1778
rect 12043 3322 13742 3350
rect 12043 1778 13658 3322
rect 13722 1778 13742 3322
rect 12043 1750 13742 1778
rect 13762 3322 15461 3350
rect 13762 1778 15377 3322
rect 15441 1778 15461 3322
rect 13762 1750 15461 1778
rect -15461 1622 -13762 1650
rect -15461 78 -13846 1622
rect -13782 78 -13762 1622
rect -15461 50 -13762 78
rect -13742 1622 -12043 1650
rect -13742 78 -12127 1622
rect -12063 78 -12043 1622
rect -13742 50 -12043 78
rect -12023 1622 -10324 1650
rect -12023 78 -10408 1622
rect -10344 78 -10324 1622
rect -12023 50 -10324 78
rect -10304 1622 -8605 1650
rect -10304 78 -8689 1622
rect -8625 78 -8605 1622
rect -10304 50 -8605 78
rect -8585 1622 -6886 1650
rect -8585 78 -6970 1622
rect -6906 78 -6886 1622
rect -8585 50 -6886 78
rect -6866 1622 -5167 1650
rect -6866 78 -5251 1622
rect -5187 78 -5167 1622
rect -6866 50 -5167 78
rect -5147 1622 -3448 1650
rect -5147 78 -3532 1622
rect -3468 78 -3448 1622
rect -5147 50 -3448 78
rect -3428 1622 -1729 1650
rect -3428 78 -1813 1622
rect -1749 78 -1729 1622
rect -3428 50 -1729 78
rect -1709 1622 -10 1650
rect -1709 78 -94 1622
rect -30 78 -10 1622
rect -1709 50 -10 78
rect 10 1622 1709 1650
rect 10 78 1625 1622
rect 1689 78 1709 1622
rect 10 50 1709 78
rect 1729 1622 3428 1650
rect 1729 78 3344 1622
rect 3408 78 3428 1622
rect 1729 50 3428 78
rect 3448 1622 5147 1650
rect 3448 78 5063 1622
rect 5127 78 5147 1622
rect 3448 50 5147 78
rect 5167 1622 6866 1650
rect 5167 78 6782 1622
rect 6846 78 6866 1622
rect 5167 50 6866 78
rect 6886 1622 8585 1650
rect 6886 78 8501 1622
rect 8565 78 8585 1622
rect 6886 50 8585 78
rect 8605 1622 10304 1650
rect 8605 78 10220 1622
rect 10284 78 10304 1622
rect 8605 50 10304 78
rect 10324 1622 12023 1650
rect 10324 78 11939 1622
rect 12003 78 12023 1622
rect 10324 50 12023 78
rect 12043 1622 13742 1650
rect 12043 78 13658 1622
rect 13722 78 13742 1622
rect 12043 50 13742 78
rect 13762 1622 15461 1650
rect 13762 78 15377 1622
rect 15441 78 15461 1622
rect 13762 50 15461 78
rect -15461 -78 -13762 -50
rect -15461 -1622 -13846 -78
rect -13782 -1622 -13762 -78
rect -15461 -1650 -13762 -1622
rect -13742 -78 -12043 -50
rect -13742 -1622 -12127 -78
rect -12063 -1622 -12043 -78
rect -13742 -1650 -12043 -1622
rect -12023 -78 -10324 -50
rect -12023 -1622 -10408 -78
rect -10344 -1622 -10324 -78
rect -12023 -1650 -10324 -1622
rect -10304 -78 -8605 -50
rect -10304 -1622 -8689 -78
rect -8625 -1622 -8605 -78
rect -10304 -1650 -8605 -1622
rect -8585 -78 -6886 -50
rect -8585 -1622 -6970 -78
rect -6906 -1622 -6886 -78
rect -8585 -1650 -6886 -1622
rect -6866 -78 -5167 -50
rect -6866 -1622 -5251 -78
rect -5187 -1622 -5167 -78
rect -6866 -1650 -5167 -1622
rect -5147 -78 -3448 -50
rect -5147 -1622 -3532 -78
rect -3468 -1622 -3448 -78
rect -5147 -1650 -3448 -1622
rect -3428 -78 -1729 -50
rect -3428 -1622 -1813 -78
rect -1749 -1622 -1729 -78
rect -3428 -1650 -1729 -1622
rect -1709 -78 -10 -50
rect -1709 -1622 -94 -78
rect -30 -1622 -10 -78
rect -1709 -1650 -10 -1622
rect 10 -78 1709 -50
rect 10 -1622 1625 -78
rect 1689 -1622 1709 -78
rect 10 -1650 1709 -1622
rect 1729 -78 3428 -50
rect 1729 -1622 3344 -78
rect 3408 -1622 3428 -78
rect 1729 -1650 3428 -1622
rect 3448 -78 5147 -50
rect 3448 -1622 5063 -78
rect 5127 -1622 5147 -78
rect 3448 -1650 5147 -1622
rect 5167 -78 6866 -50
rect 5167 -1622 6782 -78
rect 6846 -1622 6866 -78
rect 5167 -1650 6866 -1622
rect 6886 -78 8585 -50
rect 6886 -1622 8501 -78
rect 8565 -1622 8585 -78
rect 6886 -1650 8585 -1622
rect 8605 -78 10304 -50
rect 8605 -1622 10220 -78
rect 10284 -1622 10304 -78
rect 8605 -1650 10304 -1622
rect 10324 -78 12023 -50
rect 10324 -1622 11939 -78
rect 12003 -1622 12023 -78
rect 10324 -1650 12023 -1622
rect 12043 -78 13742 -50
rect 12043 -1622 13658 -78
rect 13722 -1622 13742 -78
rect 12043 -1650 13742 -1622
rect 13762 -78 15461 -50
rect 13762 -1622 15377 -78
rect 15441 -1622 15461 -78
rect 13762 -1650 15461 -1622
rect -15461 -1778 -13762 -1750
rect -15461 -3322 -13846 -1778
rect -13782 -3322 -13762 -1778
rect -15461 -3350 -13762 -3322
rect -13742 -1778 -12043 -1750
rect -13742 -3322 -12127 -1778
rect -12063 -3322 -12043 -1778
rect -13742 -3350 -12043 -3322
rect -12023 -1778 -10324 -1750
rect -12023 -3322 -10408 -1778
rect -10344 -3322 -10324 -1778
rect -12023 -3350 -10324 -3322
rect -10304 -1778 -8605 -1750
rect -10304 -3322 -8689 -1778
rect -8625 -3322 -8605 -1778
rect -10304 -3350 -8605 -3322
rect -8585 -1778 -6886 -1750
rect -8585 -3322 -6970 -1778
rect -6906 -3322 -6886 -1778
rect -8585 -3350 -6886 -3322
rect -6866 -1778 -5167 -1750
rect -6866 -3322 -5251 -1778
rect -5187 -3322 -5167 -1778
rect -6866 -3350 -5167 -3322
rect -5147 -1778 -3448 -1750
rect -5147 -3322 -3532 -1778
rect -3468 -3322 -3448 -1778
rect -5147 -3350 -3448 -3322
rect -3428 -1778 -1729 -1750
rect -3428 -3322 -1813 -1778
rect -1749 -3322 -1729 -1778
rect -3428 -3350 -1729 -3322
rect -1709 -1778 -10 -1750
rect -1709 -3322 -94 -1778
rect -30 -3322 -10 -1778
rect -1709 -3350 -10 -3322
rect 10 -1778 1709 -1750
rect 10 -3322 1625 -1778
rect 1689 -3322 1709 -1778
rect 10 -3350 1709 -3322
rect 1729 -1778 3428 -1750
rect 1729 -3322 3344 -1778
rect 3408 -3322 3428 -1778
rect 1729 -3350 3428 -3322
rect 3448 -1778 5147 -1750
rect 3448 -3322 5063 -1778
rect 5127 -3322 5147 -1778
rect 3448 -3350 5147 -3322
rect 5167 -1778 6866 -1750
rect 5167 -3322 6782 -1778
rect 6846 -3322 6866 -1778
rect 5167 -3350 6866 -3322
rect 6886 -1778 8585 -1750
rect 6886 -3322 8501 -1778
rect 8565 -3322 8585 -1778
rect 6886 -3350 8585 -3322
rect 8605 -1778 10304 -1750
rect 8605 -3322 10220 -1778
rect 10284 -3322 10304 -1778
rect 8605 -3350 10304 -3322
rect 10324 -1778 12023 -1750
rect 10324 -3322 11939 -1778
rect 12003 -3322 12023 -1778
rect 10324 -3350 12023 -3322
rect 12043 -1778 13742 -1750
rect 12043 -3322 13658 -1778
rect 13722 -3322 13742 -1778
rect 12043 -3350 13742 -3322
rect 13762 -1778 15461 -1750
rect 13762 -3322 15377 -1778
rect 15441 -3322 15461 -1778
rect 13762 -3350 15461 -3322
rect -15461 -3478 -13762 -3450
rect -15461 -5022 -13846 -3478
rect -13782 -5022 -13762 -3478
rect -15461 -5050 -13762 -5022
rect -13742 -3478 -12043 -3450
rect -13742 -5022 -12127 -3478
rect -12063 -5022 -12043 -3478
rect -13742 -5050 -12043 -5022
rect -12023 -3478 -10324 -3450
rect -12023 -5022 -10408 -3478
rect -10344 -5022 -10324 -3478
rect -12023 -5050 -10324 -5022
rect -10304 -3478 -8605 -3450
rect -10304 -5022 -8689 -3478
rect -8625 -5022 -8605 -3478
rect -10304 -5050 -8605 -5022
rect -8585 -3478 -6886 -3450
rect -8585 -5022 -6970 -3478
rect -6906 -5022 -6886 -3478
rect -8585 -5050 -6886 -5022
rect -6866 -3478 -5167 -3450
rect -6866 -5022 -5251 -3478
rect -5187 -5022 -5167 -3478
rect -6866 -5050 -5167 -5022
rect -5147 -3478 -3448 -3450
rect -5147 -5022 -3532 -3478
rect -3468 -5022 -3448 -3478
rect -5147 -5050 -3448 -5022
rect -3428 -3478 -1729 -3450
rect -3428 -5022 -1813 -3478
rect -1749 -5022 -1729 -3478
rect -3428 -5050 -1729 -5022
rect -1709 -3478 -10 -3450
rect -1709 -5022 -94 -3478
rect -30 -5022 -10 -3478
rect -1709 -5050 -10 -5022
rect 10 -3478 1709 -3450
rect 10 -5022 1625 -3478
rect 1689 -5022 1709 -3478
rect 10 -5050 1709 -5022
rect 1729 -3478 3428 -3450
rect 1729 -5022 3344 -3478
rect 3408 -5022 3428 -3478
rect 1729 -5050 3428 -5022
rect 3448 -3478 5147 -3450
rect 3448 -5022 5063 -3478
rect 5127 -5022 5147 -3478
rect 3448 -5050 5147 -5022
rect 5167 -3478 6866 -3450
rect 5167 -5022 6782 -3478
rect 6846 -5022 6866 -3478
rect 5167 -5050 6866 -5022
rect 6886 -3478 8585 -3450
rect 6886 -5022 8501 -3478
rect 8565 -5022 8585 -3478
rect 6886 -5050 8585 -5022
rect 8605 -3478 10304 -3450
rect 8605 -5022 10220 -3478
rect 10284 -5022 10304 -3478
rect 8605 -5050 10304 -5022
rect 10324 -3478 12023 -3450
rect 10324 -5022 11939 -3478
rect 12003 -5022 12023 -3478
rect 10324 -5050 12023 -5022
rect 12043 -3478 13742 -3450
rect 12043 -5022 13658 -3478
rect 13722 -5022 13742 -3478
rect 12043 -5050 13742 -5022
rect 13762 -3478 15461 -3450
rect 13762 -5022 15377 -3478
rect 15441 -5022 15461 -3478
rect 13762 -5050 15461 -5022
rect -15461 -5178 -13762 -5150
rect -15461 -6722 -13846 -5178
rect -13782 -6722 -13762 -5178
rect -15461 -6750 -13762 -6722
rect -13742 -5178 -12043 -5150
rect -13742 -6722 -12127 -5178
rect -12063 -6722 -12043 -5178
rect -13742 -6750 -12043 -6722
rect -12023 -5178 -10324 -5150
rect -12023 -6722 -10408 -5178
rect -10344 -6722 -10324 -5178
rect -12023 -6750 -10324 -6722
rect -10304 -5178 -8605 -5150
rect -10304 -6722 -8689 -5178
rect -8625 -6722 -8605 -5178
rect -10304 -6750 -8605 -6722
rect -8585 -5178 -6886 -5150
rect -8585 -6722 -6970 -5178
rect -6906 -6722 -6886 -5178
rect -8585 -6750 -6886 -6722
rect -6866 -5178 -5167 -5150
rect -6866 -6722 -5251 -5178
rect -5187 -6722 -5167 -5178
rect -6866 -6750 -5167 -6722
rect -5147 -5178 -3448 -5150
rect -5147 -6722 -3532 -5178
rect -3468 -6722 -3448 -5178
rect -5147 -6750 -3448 -6722
rect -3428 -5178 -1729 -5150
rect -3428 -6722 -1813 -5178
rect -1749 -6722 -1729 -5178
rect -3428 -6750 -1729 -6722
rect -1709 -5178 -10 -5150
rect -1709 -6722 -94 -5178
rect -30 -6722 -10 -5178
rect -1709 -6750 -10 -6722
rect 10 -5178 1709 -5150
rect 10 -6722 1625 -5178
rect 1689 -6722 1709 -5178
rect 10 -6750 1709 -6722
rect 1729 -5178 3428 -5150
rect 1729 -6722 3344 -5178
rect 3408 -6722 3428 -5178
rect 1729 -6750 3428 -6722
rect 3448 -5178 5147 -5150
rect 3448 -6722 5063 -5178
rect 5127 -6722 5147 -5178
rect 3448 -6750 5147 -6722
rect 5167 -5178 6866 -5150
rect 5167 -6722 6782 -5178
rect 6846 -6722 6866 -5178
rect 5167 -6750 6866 -6722
rect 6886 -5178 8585 -5150
rect 6886 -6722 8501 -5178
rect 8565 -6722 8585 -5178
rect 6886 -6750 8585 -6722
rect 8605 -5178 10304 -5150
rect 8605 -6722 10220 -5178
rect 10284 -6722 10304 -5178
rect 8605 -6750 10304 -6722
rect 10324 -5178 12023 -5150
rect 10324 -6722 11939 -5178
rect 12003 -6722 12023 -5178
rect 10324 -6750 12023 -6722
rect 12043 -5178 13742 -5150
rect 12043 -6722 13658 -5178
rect 13722 -6722 13742 -5178
rect 12043 -6750 13742 -6722
rect 13762 -5178 15461 -5150
rect 13762 -6722 15377 -5178
rect 15441 -6722 15461 -5178
rect 13762 -6750 15461 -6722
rect -15461 -6878 -13762 -6850
rect -15461 -8422 -13846 -6878
rect -13782 -8422 -13762 -6878
rect -15461 -8450 -13762 -8422
rect -13742 -6878 -12043 -6850
rect -13742 -8422 -12127 -6878
rect -12063 -8422 -12043 -6878
rect -13742 -8450 -12043 -8422
rect -12023 -6878 -10324 -6850
rect -12023 -8422 -10408 -6878
rect -10344 -8422 -10324 -6878
rect -12023 -8450 -10324 -8422
rect -10304 -6878 -8605 -6850
rect -10304 -8422 -8689 -6878
rect -8625 -8422 -8605 -6878
rect -10304 -8450 -8605 -8422
rect -8585 -6878 -6886 -6850
rect -8585 -8422 -6970 -6878
rect -6906 -8422 -6886 -6878
rect -8585 -8450 -6886 -8422
rect -6866 -6878 -5167 -6850
rect -6866 -8422 -5251 -6878
rect -5187 -8422 -5167 -6878
rect -6866 -8450 -5167 -8422
rect -5147 -6878 -3448 -6850
rect -5147 -8422 -3532 -6878
rect -3468 -8422 -3448 -6878
rect -5147 -8450 -3448 -8422
rect -3428 -6878 -1729 -6850
rect -3428 -8422 -1813 -6878
rect -1749 -8422 -1729 -6878
rect -3428 -8450 -1729 -8422
rect -1709 -6878 -10 -6850
rect -1709 -8422 -94 -6878
rect -30 -8422 -10 -6878
rect -1709 -8450 -10 -8422
rect 10 -6878 1709 -6850
rect 10 -8422 1625 -6878
rect 1689 -8422 1709 -6878
rect 10 -8450 1709 -8422
rect 1729 -6878 3428 -6850
rect 1729 -8422 3344 -6878
rect 3408 -8422 3428 -6878
rect 1729 -8450 3428 -8422
rect 3448 -6878 5147 -6850
rect 3448 -8422 5063 -6878
rect 5127 -8422 5147 -6878
rect 3448 -8450 5147 -8422
rect 5167 -6878 6866 -6850
rect 5167 -8422 6782 -6878
rect 6846 -8422 6866 -6878
rect 5167 -8450 6866 -8422
rect 6886 -6878 8585 -6850
rect 6886 -8422 8501 -6878
rect 8565 -8422 8585 -6878
rect 6886 -8450 8585 -8422
rect 8605 -6878 10304 -6850
rect 8605 -8422 10220 -6878
rect 10284 -8422 10304 -6878
rect 8605 -8450 10304 -8422
rect 10324 -6878 12023 -6850
rect 10324 -8422 11939 -6878
rect 12003 -8422 12023 -6878
rect 10324 -8450 12023 -8422
rect 12043 -6878 13742 -6850
rect 12043 -8422 13658 -6878
rect 13722 -8422 13742 -6878
rect 12043 -8450 13742 -8422
rect 13762 -6878 15461 -6850
rect 13762 -8422 15377 -6878
rect 15441 -8422 15461 -6878
rect 13762 -8450 15461 -8422
rect -15461 -8578 -13762 -8550
rect -15461 -10122 -13846 -8578
rect -13782 -10122 -13762 -8578
rect -15461 -10150 -13762 -10122
rect -13742 -8578 -12043 -8550
rect -13742 -10122 -12127 -8578
rect -12063 -10122 -12043 -8578
rect -13742 -10150 -12043 -10122
rect -12023 -8578 -10324 -8550
rect -12023 -10122 -10408 -8578
rect -10344 -10122 -10324 -8578
rect -12023 -10150 -10324 -10122
rect -10304 -8578 -8605 -8550
rect -10304 -10122 -8689 -8578
rect -8625 -10122 -8605 -8578
rect -10304 -10150 -8605 -10122
rect -8585 -8578 -6886 -8550
rect -8585 -10122 -6970 -8578
rect -6906 -10122 -6886 -8578
rect -8585 -10150 -6886 -10122
rect -6866 -8578 -5167 -8550
rect -6866 -10122 -5251 -8578
rect -5187 -10122 -5167 -8578
rect -6866 -10150 -5167 -10122
rect -5147 -8578 -3448 -8550
rect -5147 -10122 -3532 -8578
rect -3468 -10122 -3448 -8578
rect -5147 -10150 -3448 -10122
rect -3428 -8578 -1729 -8550
rect -3428 -10122 -1813 -8578
rect -1749 -10122 -1729 -8578
rect -3428 -10150 -1729 -10122
rect -1709 -8578 -10 -8550
rect -1709 -10122 -94 -8578
rect -30 -10122 -10 -8578
rect -1709 -10150 -10 -10122
rect 10 -8578 1709 -8550
rect 10 -10122 1625 -8578
rect 1689 -10122 1709 -8578
rect 10 -10150 1709 -10122
rect 1729 -8578 3428 -8550
rect 1729 -10122 3344 -8578
rect 3408 -10122 3428 -8578
rect 1729 -10150 3428 -10122
rect 3448 -8578 5147 -8550
rect 3448 -10122 5063 -8578
rect 5127 -10122 5147 -8578
rect 3448 -10150 5147 -10122
rect 5167 -8578 6866 -8550
rect 5167 -10122 6782 -8578
rect 6846 -10122 6866 -8578
rect 5167 -10150 6866 -10122
rect 6886 -8578 8585 -8550
rect 6886 -10122 8501 -8578
rect 8565 -10122 8585 -8578
rect 6886 -10150 8585 -10122
rect 8605 -8578 10304 -8550
rect 8605 -10122 10220 -8578
rect 10284 -10122 10304 -8578
rect 8605 -10150 10304 -10122
rect 10324 -8578 12023 -8550
rect 10324 -10122 11939 -8578
rect 12003 -10122 12023 -8578
rect 10324 -10150 12023 -10122
rect 12043 -8578 13742 -8550
rect 12043 -10122 13658 -8578
rect 13722 -10122 13742 -8578
rect 12043 -10150 13742 -10122
rect 13762 -8578 15461 -8550
rect 13762 -10122 15377 -8578
rect 15441 -10122 15461 -8578
rect 13762 -10150 15461 -10122
rect -15461 -10278 -13762 -10250
rect -15461 -11822 -13846 -10278
rect -13782 -11822 -13762 -10278
rect -15461 -11850 -13762 -11822
rect -13742 -10278 -12043 -10250
rect -13742 -11822 -12127 -10278
rect -12063 -11822 -12043 -10278
rect -13742 -11850 -12043 -11822
rect -12023 -10278 -10324 -10250
rect -12023 -11822 -10408 -10278
rect -10344 -11822 -10324 -10278
rect -12023 -11850 -10324 -11822
rect -10304 -10278 -8605 -10250
rect -10304 -11822 -8689 -10278
rect -8625 -11822 -8605 -10278
rect -10304 -11850 -8605 -11822
rect -8585 -10278 -6886 -10250
rect -8585 -11822 -6970 -10278
rect -6906 -11822 -6886 -10278
rect -8585 -11850 -6886 -11822
rect -6866 -10278 -5167 -10250
rect -6866 -11822 -5251 -10278
rect -5187 -11822 -5167 -10278
rect -6866 -11850 -5167 -11822
rect -5147 -10278 -3448 -10250
rect -5147 -11822 -3532 -10278
rect -3468 -11822 -3448 -10278
rect -5147 -11850 -3448 -11822
rect -3428 -10278 -1729 -10250
rect -3428 -11822 -1813 -10278
rect -1749 -11822 -1729 -10278
rect -3428 -11850 -1729 -11822
rect -1709 -10278 -10 -10250
rect -1709 -11822 -94 -10278
rect -30 -11822 -10 -10278
rect -1709 -11850 -10 -11822
rect 10 -10278 1709 -10250
rect 10 -11822 1625 -10278
rect 1689 -11822 1709 -10278
rect 10 -11850 1709 -11822
rect 1729 -10278 3428 -10250
rect 1729 -11822 3344 -10278
rect 3408 -11822 3428 -10278
rect 1729 -11850 3428 -11822
rect 3448 -10278 5147 -10250
rect 3448 -11822 5063 -10278
rect 5127 -11822 5147 -10278
rect 3448 -11850 5147 -11822
rect 5167 -10278 6866 -10250
rect 5167 -11822 6782 -10278
rect 6846 -11822 6866 -10278
rect 5167 -11850 6866 -11822
rect 6886 -10278 8585 -10250
rect 6886 -11822 8501 -10278
rect 8565 -11822 8585 -10278
rect 6886 -11850 8585 -11822
rect 8605 -10278 10304 -10250
rect 8605 -11822 10220 -10278
rect 10284 -11822 10304 -10278
rect 8605 -11850 10304 -11822
rect 10324 -10278 12023 -10250
rect 10324 -11822 11939 -10278
rect 12003 -11822 12023 -10278
rect 10324 -11850 12023 -11822
rect 12043 -10278 13742 -10250
rect 12043 -11822 13658 -10278
rect 13722 -11822 13742 -10278
rect 12043 -11850 13742 -11822
rect 13762 -10278 15461 -10250
rect 13762 -11822 15377 -10278
rect 15441 -11822 15461 -10278
rect 13762 -11850 15461 -11822
rect -15461 -11978 -13762 -11950
rect -15461 -13522 -13846 -11978
rect -13782 -13522 -13762 -11978
rect -15461 -13550 -13762 -13522
rect -13742 -11978 -12043 -11950
rect -13742 -13522 -12127 -11978
rect -12063 -13522 -12043 -11978
rect -13742 -13550 -12043 -13522
rect -12023 -11978 -10324 -11950
rect -12023 -13522 -10408 -11978
rect -10344 -13522 -10324 -11978
rect -12023 -13550 -10324 -13522
rect -10304 -11978 -8605 -11950
rect -10304 -13522 -8689 -11978
rect -8625 -13522 -8605 -11978
rect -10304 -13550 -8605 -13522
rect -8585 -11978 -6886 -11950
rect -8585 -13522 -6970 -11978
rect -6906 -13522 -6886 -11978
rect -8585 -13550 -6886 -13522
rect -6866 -11978 -5167 -11950
rect -6866 -13522 -5251 -11978
rect -5187 -13522 -5167 -11978
rect -6866 -13550 -5167 -13522
rect -5147 -11978 -3448 -11950
rect -5147 -13522 -3532 -11978
rect -3468 -13522 -3448 -11978
rect -5147 -13550 -3448 -13522
rect -3428 -11978 -1729 -11950
rect -3428 -13522 -1813 -11978
rect -1749 -13522 -1729 -11978
rect -3428 -13550 -1729 -13522
rect -1709 -11978 -10 -11950
rect -1709 -13522 -94 -11978
rect -30 -13522 -10 -11978
rect -1709 -13550 -10 -13522
rect 10 -11978 1709 -11950
rect 10 -13522 1625 -11978
rect 1689 -13522 1709 -11978
rect 10 -13550 1709 -13522
rect 1729 -11978 3428 -11950
rect 1729 -13522 3344 -11978
rect 3408 -13522 3428 -11978
rect 1729 -13550 3428 -13522
rect 3448 -11978 5147 -11950
rect 3448 -13522 5063 -11978
rect 5127 -13522 5147 -11978
rect 3448 -13550 5147 -13522
rect 5167 -11978 6866 -11950
rect 5167 -13522 6782 -11978
rect 6846 -13522 6866 -11978
rect 5167 -13550 6866 -13522
rect 6886 -11978 8585 -11950
rect 6886 -13522 8501 -11978
rect 8565 -13522 8585 -11978
rect 6886 -13550 8585 -13522
rect 8605 -11978 10304 -11950
rect 8605 -13522 10220 -11978
rect 10284 -13522 10304 -11978
rect 8605 -13550 10304 -13522
rect 10324 -11978 12023 -11950
rect 10324 -13522 11939 -11978
rect 12003 -13522 12023 -11978
rect 10324 -13550 12023 -13522
rect 12043 -11978 13742 -11950
rect 12043 -13522 13658 -11978
rect 13722 -13522 13742 -11978
rect 12043 -13550 13742 -13522
rect 13762 -11978 15461 -11950
rect 13762 -13522 15377 -11978
rect 15441 -13522 15461 -11978
rect 13762 -13550 15461 -13522
rect -15461 -13678 -13762 -13650
rect -15461 -15222 -13846 -13678
rect -13782 -15222 -13762 -13678
rect -15461 -15250 -13762 -15222
rect -13742 -13678 -12043 -13650
rect -13742 -15222 -12127 -13678
rect -12063 -15222 -12043 -13678
rect -13742 -15250 -12043 -15222
rect -12023 -13678 -10324 -13650
rect -12023 -15222 -10408 -13678
rect -10344 -15222 -10324 -13678
rect -12023 -15250 -10324 -15222
rect -10304 -13678 -8605 -13650
rect -10304 -15222 -8689 -13678
rect -8625 -15222 -8605 -13678
rect -10304 -15250 -8605 -15222
rect -8585 -13678 -6886 -13650
rect -8585 -15222 -6970 -13678
rect -6906 -15222 -6886 -13678
rect -8585 -15250 -6886 -15222
rect -6866 -13678 -5167 -13650
rect -6866 -15222 -5251 -13678
rect -5187 -15222 -5167 -13678
rect -6866 -15250 -5167 -15222
rect -5147 -13678 -3448 -13650
rect -5147 -15222 -3532 -13678
rect -3468 -15222 -3448 -13678
rect -5147 -15250 -3448 -15222
rect -3428 -13678 -1729 -13650
rect -3428 -15222 -1813 -13678
rect -1749 -15222 -1729 -13678
rect -3428 -15250 -1729 -15222
rect -1709 -13678 -10 -13650
rect -1709 -15222 -94 -13678
rect -30 -15222 -10 -13678
rect -1709 -15250 -10 -15222
rect 10 -13678 1709 -13650
rect 10 -15222 1625 -13678
rect 1689 -15222 1709 -13678
rect 10 -15250 1709 -15222
rect 1729 -13678 3428 -13650
rect 1729 -15222 3344 -13678
rect 3408 -15222 3428 -13678
rect 1729 -15250 3428 -15222
rect 3448 -13678 5147 -13650
rect 3448 -15222 5063 -13678
rect 5127 -15222 5147 -13678
rect 3448 -15250 5147 -15222
rect 5167 -13678 6866 -13650
rect 5167 -15222 6782 -13678
rect 6846 -15222 6866 -13678
rect 5167 -15250 6866 -15222
rect 6886 -13678 8585 -13650
rect 6886 -15222 8501 -13678
rect 8565 -15222 8585 -13678
rect 6886 -15250 8585 -15222
rect 8605 -13678 10304 -13650
rect 8605 -15222 10220 -13678
rect 10284 -15222 10304 -13678
rect 8605 -15250 10304 -15222
rect 10324 -13678 12023 -13650
rect 10324 -15222 11939 -13678
rect 12003 -15222 12023 -13678
rect 10324 -15250 12023 -15222
rect 12043 -13678 13742 -13650
rect 12043 -15222 13658 -13678
rect 13722 -15222 13742 -13678
rect 12043 -15250 13742 -15222
rect 13762 -13678 15461 -13650
rect 13762 -15222 15377 -13678
rect 15441 -15222 15461 -13678
rect 13762 -15250 15461 -15222
<< via3 >>
rect -13846 13678 -13782 15222
rect -12127 13678 -12063 15222
rect -10408 13678 -10344 15222
rect -8689 13678 -8625 15222
rect -6970 13678 -6906 15222
rect -5251 13678 -5187 15222
rect -3532 13678 -3468 15222
rect -1813 13678 -1749 15222
rect -94 13678 -30 15222
rect 1625 13678 1689 15222
rect 3344 13678 3408 15222
rect 5063 13678 5127 15222
rect 6782 13678 6846 15222
rect 8501 13678 8565 15222
rect 10220 13678 10284 15222
rect 11939 13678 12003 15222
rect 13658 13678 13722 15222
rect 15377 13678 15441 15222
rect -13846 11978 -13782 13522
rect -12127 11978 -12063 13522
rect -10408 11978 -10344 13522
rect -8689 11978 -8625 13522
rect -6970 11978 -6906 13522
rect -5251 11978 -5187 13522
rect -3532 11978 -3468 13522
rect -1813 11978 -1749 13522
rect -94 11978 -30 13522
rect 1625 11978 1689 13522
rect 3344 11978 3408 13522
rect 5063 11978 5127 13522
rect 6782 11978 6846 13522
rect 8501 11978 8565 13522
rect 10220 11978 10284 13522
rect 11939 11978 12003 13522
rect 13658 11978 13722 13522
rect 15377 11978 15441 13522
rect -13846 10278 -13782 11822
rect -12127 10278 -12063 11822
rect -10408 10278 -10344 11822
rect -8689 10278 -8625 11822
rect -6970 10278 -6906 11822
rect -5251 10278 -5187 11822
rect -3532 10278 -3468 11822
rect -1813 10278 -1749 11822
rect -94 10278 -30 11822
rect 1625 10278 1689 11822
rect 3344 10278 3408 11822
rect 5063 10278 5127 11822
rect 6782 10278 6846 11822
rect 8501 10278 8565 11822
rect 10220 10278 10284 11822
rect 11939 10278 12003 11822
rect 13658 10278 13722 11822
rect 15377 10278 15441 11822
rect -13846 8578 -13782 10122
rect -12127 8578 -12063 10122
rect -10408 8578 -10344 10122
rect -8689 8578 -8625 10122
rect -6970 8578 -6906 10122
rect -5251 8578 -5187 10122
rect -3532 8578 -3468 10122
rect -1813 8578 -1749 10122
rect -94 8578 -30 10122
rect 1625 8578 1689 10122
rect 3344 8578 3408 10122
rect 5063 8578 5127 10122
rect 6782 8578 6846 10122
rect 8501 8578 8565 10122
rect 10220 8578 10284 10122
rect 11939 8578 12003 10122
rect 13658 8578 13722 10122
rect 15377 8578 15441 10122
rect -13846 6878 -13782 8422
rect -12127 6878 -12063 8422
rect -10408 6878 -10344 8422
rect -8689 6878 -8625 8422
rect -6970 6878 -6906 8422
rect -5251 6878 -5187 8422
rect -3532 6878 -3468 8422
rect -1813 6878 -1749 8422
rect -94 6878 -30 8422
rect 1625 6878 1689 8422
rect 3344 6878 3408 8422
rect 5063 6878 5127 8422
rect 6782 6878 6846 8422
rect 8501 6878 8565 8422
rect 10220 6878 10284 8422
rect 11939 6878 12003 8422
rect 13658 6878 13722 8422
rect 15377 6878 15441 8422
rect -13846 5178 -13782 6722
rect -12127 5178 -12063 6722
rect -10408 5178 -10344 6722
rect -8689 5178 -8625 6722
rect -6970 5178 -6906 6722
rect -5251 5178 -5187 6722
rect -3532 5178 -3468 6722
rect -1813 5178 -1749 6722
rect -94 5178 -30 6722
rect 1625 5178 1689 6722
rect 3344 5178 3408 6722
rect 5063 5178 5127 6722
rect 6782 5178 6846 6722
rect 8501 5178 8565 6722
rect 10220 5178 10284 6722
rect 11939 5178 12003 6722
rect 13658 5178 13722 6722
rect 15377 5178 15441 6722
rect -13846 3478 -13782 5022
rect -12127 3478 -12063 5022
rect -10408 3478 -10344 5022
rect -8689 3478 -8625 5022
rect -6970 3478 -6906 5022
rect -5251 3478 -5187 5022
rect -3532 3478 -3468 5022
rect -1813 3478 -1749 5022
rect -94 3478 -30 5022
rect 1625 3478 1689 5022
rect 3344 3478 3408 5022
rect 5063 3478 5127 5022
rect 6782 3478 6846 5022
rect 8501 3478 8565 5022
rect 10220 3478 10284 5022
rect 11939 3478 12003 5022
rect 13658 3478 13722 5022
rect 15377 3478 15441 5022
rect -13846 1778 -13782 3322
rect -12127 1778 -12063 3322
rect -10408 1778 -10344 3322
rect -8689 1778 -8625 3322
rect -6970 1778 -6906 3322
rect -5251 1778 -5187 3322
rect -3532 1778 -3468 3322
rect -1813 1778 -1749 3322
rect -94 1778 -30 3322
rect 1625 1778 1689 3322
rect 3344 1778 3408 3322
rect 5063 1778 5127 3322
rect 6782 1778 6846 3322
rect 8501 1778 8565 3322
rect 10220 1778 10284 3322
rect 11939 1778 12003 3322
rect 13658 1778 13722 3322
rect 15377 1778 15441 3322
rect -13846 78 -13782 1622
rect -12127 78 -12063 1622
rect -10408 78 -10344 1622
rect -8689 78 -8625 1622
rect -6970 78 -6906 1622
rect -5251 78 -5187 1622
rect -3532 78 -3468 1622
rect -1813 78 -1749 1622
rect -94 78 -30 1622
rect 1625 78 1689 1622
rect 3344 78 3408 1622
rect 5063 78 5127 1622
rect 6782 78 6846 1622
rect 8501 78 8565 1622
rect 10220 78 10284 1622
rect 11939 78 12003 1622
rect 13658 78 13722 1622
rect 15377 78 15441 1622
rect -13846 -1622 -13782 -78
rect -12127 -1622 -12063 -78
rect -10408 -1622 -10344 -78
rect -8689 -1622 -8625 -78
rect -6970 -1622 -6906 -78
rect -5251 -1622 -5187 -78
rect -3532 -1622 -3468 -78
rect -1813 -1622 -1749 -78
rect -94 -1622 -30 -78
rect 1625 -1622 1689 -78
rect 3344 -1622 3408 -78
rect 5063 -1622 5127 -78
rect 6782 -1622 6846 -78
rect 8501 -1622 8565 -78
rect 10220 -1622 10284 -78
rect 11939 -1622 12003 -78
rect 13658 -1622 13722 -78
rect 15377 -1622 15441 -78
rect -13846 -3322 -13782 -1778
rect -12127 -3322 -12063 -1778
rect -10408 -3322 -10344 -1778
rect -8689 -3322 -8625 -1778
rect -6970 -3322 -6906 -1778
rect -5251 -3322 -5187 -1778
rect -3532 -3322 -3468 -1778
rect -1813 -3322 -1749 -1778
rect -94 -3322 -30 -1778
rect 1625 -3322 1689 -1778
rect 3344 -3322 3408 -1778
rect 5063 -3322 5127 -1778
rect 6782 -3322 6846 -1778
rect 8501 -3322 8565 -1778
rect 10220 -3322 10284 -1778
rect 11939 -3322 12003 -1778
rect 13658 -3322 13722 -1778
rect 15377 -3322 15441 -1778
rect -13846 -5022 -13782 -3478
rect -12127 -5022 -12063 -3478
rect -10408 -5022 -10344 -3478
rect -8689 -5022 -8625 -3478
rect -6970 -5022 -6906 -3478
rect -5251 -5022 -5187 -3478
rect -3532 -5022 -3468 -3478
rect -1813 -5022 -1749 -3478
rect -94 -5022 -30 -3478
rect 1625 -5022 1689 -3478
rect 3344 -5022 3408 -3478
rect 5063 -5022 5127 -3478
rect 6782 -5022 6846 -3478
rect 8501 -5022 8565 -3478
rect 10220 -5022 10284 -3478
rect 11939 -5022 12003 -3478
rect 13658 -5022 13722 -3478
rect 15377 -5022 15441 -3478
rect -13846 -6722 -13782 -5178
rect -12127 -6722 -12063 -5178
rect -10408 -6722 -10344 -5178
rect -8689 -6722 -8625 -5178
rect -6970 -6722 -6906 -5178
rect -5251 -6722 -5187 -5178
rect -3532 -6722 -3468 -5178
rect -1813 -6722 -1749 -5178
rect -94 -6722 -30 -5178
rect 1625 -6722 1689 -5178
rect 3344 -6722 3408 -5178
rect 5063 -6722 5127 -5178
rect 6782 -6722 6846 -5178
rect 8501 -6722 8565 -5178
rect 10220 -6722 10284 -5178
rect 11939 -6722 12003 -5178
rect 13658 -6722 13722 -5178
rect 15377 -6722 15441 -5178
rect -13846 -8422 -13782 -6878
rect -12127 -8422 -12063 -6878
rect -10408 -8422 -10344 -6878
rect -8689 -8422 -8625 -6878
rect -6970 -8422 -6906 -6878
rect -5251 -8422 -5187 -6878
rect -3532 -8422 -3468 -6878
rect -1813 -8422 -1749 -6878
rect -94 -8422 -30 -6878
rect 1625 -8422 1689 -6878
rect 3344 -8422 3408 -6878
rect 5063 -8422 5127 -6878
rect 6782 -8422 6846 -6878
rect 8501 -8422 8565 -6878
rect 10220 -8422 10284 -6878
rect 11939 -8422 12003 -6878
rect 13658 -8422 13722 -6878
rect 15377 -8422 15441 -6878
rect -13846 -10122 -13782 -8578
rect -12127 -10122 -12063 -8578
rect -10408 -10122 -10344 -8578
rect -8689 -10122 -8625 -8578
rect -6970 -10122 -6906 -8578
rect -5251 -10122 -5187 -8578
rect -3532 -10122 -3468 -8578
rect -1813 -10122 -1749 -8578
rect -94 -10122 -30 -8578
rect 1625 -10122 1689 -8578
rect 3344 -10122 3408 -8578
rect 5063 -10122 5127 -8578
rect 6782 -10122 6846 -8578
rect 8501 -10122 8565 -8578
rect 10220 -10122 10284 -8578
rect 11939 -10122 12003 -8578
rect 13658 -10122 13722 -8578
rect 15377 -10122 15441 -8578
rect -13846 -11822 -13782 -10278
rect -12127 -11822 -12063 -10278
rect -10408 -11822 -10344 -10278
rect -8689 -11822 -8625 -10278
rect -6970 -11822 -6906 -10278
rect -5251 -11822 -5187 -10278
rect -3532 -11822 -3468 -10278
rect -1813 -11822 -1749 -10278
rect -94 -11822 -30 -10278
rect 1625 -11822 1689 -10278
rect 3344 -11822 3408 -10278
rect 5063 -11822 5127 -10278
rect 6782 -11822 6846 -10278
rect 8501 -11822 8565 -10278
rect 10220 -11822 10284 -10278
rect 11939 -11822 12003 -10278
rect 13658 -11822 13722 -10278
rect 15377 -11822 15441 -10278
rect -13846 -13522 -13782 -11978
rect -12127 -13522 -12063 -11978
rect -10408 -13522 -10344 -11978
rect -8689 -13522 -8625 -11978
rect -6970 -13522 -6906 -11978
rect -5251 -13522 -5187 -11978
rect -3532 -13522 -3468 -11978
rect -1813 -13522 -1749 -11978
rect -94 -13522 -30 -11978
rect 1625 -13522 1689 -11978
rect 3344 -13522 3408 -11978
rect 5063 -13522 5127 -11978
rect 6782 -13522 6846 -11978
rect 8501 -13522 8565 -11978
rect 10220 -13522 10284 -11978
rect 11939 -13522 12003 -11978
rect 13658 -13522 13722 -11978
rect 15377 -13522 15441 -11978
rect -13846 -15222 -13782 -13678
rect -12127 -15222 -12063 -13678
rect -10408 -15222 -10344 -13678
rect -8689 -15222 -8625 -13678
rect -6970 -15222 -6906 -13678
rect -5251 -15222 -5187 -13678
rect -3532 -15222 -3468 -13678
rect -1813 -15222 -1749 -13678
rect -94 -15222 -30 -13678
rect 1625 -15222 1689 -13678
rect 3344 -15222 3408 -13678
rect 5063 -15222 5127 -13678
rect 6782 -15222 6846 -13678
rect 8501 -15222 8565 -13678
rect 10220 -15222 10284 -13678
rect 11939 -15222 12003 -13678
rect 13658 -15222 13722 -13678
rect 15377 -15222 15441 -13678
<< mimcap >>
rect -15361 15110 -13961 15150
rect -15361 13790 -15321 15110
rect -14001 13790 -13961 15110
rect -15361 13750 -13961 13790
rect -13642 15110 -12242 15150
rect -13642 13790 -13602 15110
rect -12282 13790 -12242 15110
rect -13642 13750 -12242 13790
rect -11923 15110 -10523 15150
rect -11923 13790 -11883 15110
rect -10563 13790 -10523 15110
rect -11923 13750 -10523 13790
rect -10204 15110 -8804 15150
rect -10204 13790 -10164 15110
rect -8844 13790 -8804 15110
rect -10204 13750 -8804 13790
rect -8485 15110 -7085 15150
rect -8485 13790 -8445 15110
rect -7125 13790 -7085 15110
rect -8485 13750 -7085 13790
rect -6766 15110 -5366 15150
rect -6766 13790 -6726 15110
rect -5406 13790 -5366 15110
rect -6766 13750 -5366 13790
rect -5047 15110 -3647 15150
rect -5047 13790 -5007 15110
rect -3687 13790 -3647 15110
rect -5047 13750 -3647 13790
rect -3328 15110 -1928 15150
rect -3328 13790 -3288 15110
rect -1968 13790 -1928 15110
rect -3328 13750 -1928 13790
rect -1609 15110 -209 15150
rect -1609 13790 -1569 15110
rect -249 13790 -209 15110
rect -1609 13750 -209 13790
rect 110 15110 1510 15150
rect 110 13790 150 15110
rect 1470 13790 1510 15110
rect 110 13750 1510 13790
rect 1829 15110 3229 15150
rect 1829 13790 1869 15110
rect 3189 13790 3229 15110
rect 1829 13750 3229 13790
rect 3548 15110 4948 15150
rect 3548 13790 3588 15110
rect 4908 13790 4948 15110
rect 3548 13750 4948 13790
rect 5267 15110 6667 15150
rect 5267 13790 5307 15110
rect 6627 13790 6667 15110
rect 5267 13750 6667 13790
rect 6986 15110 8386 15150
rect 6986 13790 7026 15110
rect 8346 13790 8386 15110
rect 6986 13750 8386 13790
rect 8705 15110 10105 15150
rect 8705 13790 8745 15110
rect 10065 13790 10105 15110
rect 8705 13750 10105 13790
rect 10424 15110 11824 15150
rect 10424 13790 10464 15110
rect 11784 13790 11824 15110
rect 10424 13750 11824 13790
rect 12143 15110 13543 15150
rect 12143 13790 12183 15110
rect 13503 13790 13543 15110
rect 12143 13750 13543 13790
rect 13862 15110 15262 15150
rect 13862 13790 13902 15110
rect 15222 13790 15262 15110
rect 13862 13750 15262 13790
rect -15361 13410 -13961 13450
rect -15361 12090 -15321 13410
rect -14001 12090 -13961 13410
rect -15361 12050 -13961 12090
rect -13642 13410 -12242 13450
rect -13642 12090 -13602 13410
rect -12282 12090 -12242 13410
rect -13642 12050 -12242 12090
rect -11923 13410 -10523 13450
rect -11923 12090 -11883 13410
rect -10563 12090 -10523 13410
rect -11923 12050 -10523 12090
rect -10204 13410 -8804 13450
rect -10204 12090 -10164 13410
rect -8844 12090 -8804 13410
rect -10204 12050 -8804 12090
rect -8485 13410 -7085 13450
rect -8485 12090 -8445 13410
rect -7125 12090 -7085 13410
rect -8485 12050 -7085 12090
rect -6766 13410 -5366 13450
rect -6766 12090 -6726 13410
rect -5406 12090 -5366 13410
rect -6766 12050 -5366 12090
rect -5047 13410 -3647 13450
rect -5047 12090 -5007 13410
rect -3687 12090 -3647 13410
rect -5047 12050 -3647 12090
rect -3328 13410 -1928 13450
rect -3328 12090 -3288 13410
rect -1968 12090 -1928 13410
rect -3328 12050 -1928 12090
rect -1609 13410 -209 13450
rect -1609 12090 -1569 13410
rect -249 12090 -209 13410
rect -1609 12050 -209 12090
rect 110 13410 1510 13450
rect 110 12090 150 13410
rect 1470 12090 1510 13410
rect 110 12050 1510 12090
rect 1829 13410 3229 13450
rect 1829 12090 1869 13410
rect 3189 12090 3229 13410
rect 1829 12050 3229 12090
rect 3548 13410 4948 13450
rect 3548 12090 3588 13410
rect 4908 12090 4948 13410
rect 3548 12050 4948 12090
rect 5267 13410 6667 13450
rect 5267 12090 5307 13410
rect 6627 12090 6667 13410
rect 5267 12050 6667 12090
rect 6986 13410 8386 13450
rect 6986 12090 7026 13410
rect 8346 12090 8386 13410
rect 6986 12050 8386 12090
rect 8705 13410 10105 13450
rect 8705 12090 8745 13410
rect 10065 12090 10105 13410
rect 8705 12050 10105 12090
rect 10424 13410 11824 13450
rect 10424 12090 10464 13410
rect 11784 12090 11824 13410
rect 10424 12050 11824 12090
rect 12143 13410 13543 13450
rect 12143 12090 12183 13410
rect 13503 12090 13543 13410
rect 12143 12050 13543 12090
rect 13862 13410 15262 13450
rect 13862 12090 13902 13410
rect 15222 12090 15262 13410
rect 13862 12050 15262 12090
rect -15361 11710 -13961 11750
rect -15361 10390 -15321 11710
rect -14001 10390 -13961 11710
rect -15361 10350 -13961 10390
rect -13642 11710 -12242 11750
rect -13642 10390 -13602 11710
rect -12282 10390 -12242 11710
rect -13642 10350 -12242 10390
rect -11923 11710 -10523 11750
rect -11923 10390 -11883 11710
rect -10563 10390 -10523 11710
rect -11923 10350 -10523 10390
rect -10204 11710 -8804 11750
rect -10204 10390 -10164 11710
rect -8844 10390 -8804 11710
rect -10204 10350 -8804 10390
rect -8485 11710 -7085 11750
rect -8485 10390 -8445 11710
rect -7125 10390 -7085 11710
rect -8485 10350 -7085 10390
rect -6766 11710 -5366 11750
rect -6766 10390 -6726 11710
rect -5406 10390 -5366 11710
rect -6766 10350 -5366 10390
rect -5047 11710 -3647 11750
rect -5047 10390 -5007 11710
rect -3687 10390 -3647 11710
rect -5047 10350 -3647 10390
rect -3328 11710 -1928 11750
rect -3328 10390 -3288 11710
rect -1968 10390 -1928 11710
rect -3328 10350 -1928 10390
rect -1609 11710 -209 11750
rect -1609 10390 -1569 11710
rect -249 10390 -209 11710
rect -1609 10350 -209 10390
rect 110 11710 1510 11750
rect 110 10390 150 11710
rect 1470 10390 1510 11710
rect 110 10350 1510 10390
rect 1829 11710 3229 11750
rect 1829 10390 1869 11710
rect 3189 10390 3229 11710
rect 1829 10350 3229 10390
rect 3548 11710 4948 11750
rect 3548 10390 3588 11710
rect 4908 10390 4948 11710
rect 3548 10350 4948 10390
rect 5267 11710 6667 11750
rect 5267 10390 5307 11710
rect 6627 10390 6667 11710
rect 5267 10350 6667 10390
rect 6986 11710 8386 11750
rect 6986 10390 7026 11710
rect 8346 10390 8386 11710
rect 6986 10350 8386 10390
rect 8705 11710 10105 11750
rect 8705 10390 8745 11710
rect 10065 10390 10105 11710
rect 8705 10350 10105 10390
rect 10424 11710 11824 11750
rect 10424 10390 10464 11710
rect 11784 10390 11824 11710
rect 10424 10350 11824 10390
rect 12143 11710 13543 11750
rect 12143 10390 12183 11710
rect 13503 10390 13543 11710
rect 12143 10350 13543 10390
rect 13862 11710 15262 11750
rect 13862 10390 13902 11710
rect 15222 10390 15262 11710
rect 13862 10350 15262 10390
rect -15361 10010 -13961 10050
rect -15361 8690 -15321 10010
rect -14001 8690 -13961 10010
rect -15361 8650 -13961 8690
rect -13642 10010 -12242 10050
rect -13642 8690 -13602 10010
rect -12282 8690 -12242 10010
rect -13642 8650 -12242 8690
rect -11923 10010 -10523 10050
rect -11923 8690 -11883 10010
rect -10563 8690 -10523 10010
rect -11923 8650 -10523 8690
rect -10204 10010 -8804 10050
rect -10204 8690 -10164 10010
rect -8844 8690 -8804 10010
rect -10204 8650 -8804 8690
rect -8485 10010 -7085 10050
rect -8485 8690 -8445 10010
rect -7125 8690 -7085 10010
rect -8485 8650 -7085 8690
rect -6766 10010 -5366 10050
rect -6766 8690 -6726 10010
rect -5406 8690 -5366 10010
rect -6766 8650 -5366 8690
rect -5047 10010 -3647 10050
rect -5047 8690 -5007 10010
rect -3687 8690 -3647 10010
rect -5047 8650 -3647 8690
rect -3328 10010 -1928 10050
rect -3328 8690 -3288 10010
rect -1968 8690 -1928 10010
rect -3328 8650 -1928 8690
rect -1609 10010 -209 10050
rect -1609 8690 -1569 10010
rect -249 8690 -209 10010
rect -1609 8650 -209 8690
rect 110 10010 1510 10050
rect 110 8690 150 10010
rect 1470 8690 1510 10010
rect 110 8650 1510 8690
rect 1829 10010 3229 10050
rect 1829 8690 1869 10010
rect 3189 8690 3229 10010
rect 1829 8650 3229 8690
rect 3548 10010 4948 10050
rect 3548 8690 3588 10010
rect 4908 8690 4948 10010
rect 3548 8650 4948 8690
rect 5267 10010 6667 10050
rect 5267 8690 5307 10010
rect 6627 8690 6667 10010
rect 5267 8650 6667 8690
rect 6986 10010 8386 10050
rect 6986 8690 7026 10010
rect 8346 8690 8386 10010
rect 6986 8650 8386 8690
rect 8705 10010 10105 10050
rect 8705 8690 8745 10010
rect 10065 8690 10105 10010
rect 8705 8650 10105 8690
rect 10424 10010 11824 10050
rect 10424 8690 10464 10010
rect 11784 8690 11824 10010
rect 10424 8650 11824 8690
rect 12143 10010 13543 10050
rect 12143 8690 12183 10010
rect 13503 8690 13543 10010
rect 12143 8650 13543 8690
rect 13862 10010 15262 10050
rect 13862 8690 13902 10010
rect 15222 8690 15262 10010
rect 13862 8650 15262 8690
rect -15361 8310 -13961 8350
rect -15361 6990 -15321 8310
rect -14001 6990 -13961 8310
rect -15361 6950 -13961 6990
rect -13642 8310 -12242 8350
rect -13642 6990 -13602 8310
rect -12282 6990 -12242 8310
rect -13642 6950 -12242 6990
rect -11923 8310 -10523 8350
rect -11923 6990 -11883 8310
rect -10563 6990 -10523 8310
rect -11923 6950 -10523 6990
rect -10204 8310 -8804 8350
rect -10204 6990 -10164 8310
rect -8844 6990 -8804 8310
rect -10204 6950 -8804 6990
rect -8485 8310 -7085 8350
rect -8485 6990 -8445 8310
rect -7125 6990 -7085 8310
rect -8485 6950 -7085 6990
rect -6766 8310 -5366 8350
rect -6766 6990 -6726 8310
rect -5406 6990 -5366 8310
rect -6766 6950 -5366 6990
rect -5047 8310 -3647 8350
rect -5047 6990 -5007 8310
rect -3687 6990 -3647 8310
rect -5047 6950 -3647 6990
rect -3328 8310 -1928 8350
rect -3328 6990 -3288 8310
rect -1968 6990 -1928 8310
rect -3328 6950 -1928 6990
rect -1609 8310 -209 8350
rect -1609 6990 -1569 8310
rect -249 6990 -209 8310
rect -1609 6950 -209 6990
rect 110 8310 1510 8350
rect 110 6990 150 8310
rect 1470 6990 1510 8310
rect 110 6950 1510 6990
rect 1829 8310 3229 8350
rect 1829 6990 1869 8310
rect 3189 6990 3229 8310
rect 1829 6950 3229 6990
rect 3548 8310 4948 8350
rect 3548 6990 3588 8310
rect 4908 6990 4948 8310
rect 3548 6950 4948 6990
rect 5267 8310 6667 8350
rect 5267 6990 5307 8310
rect 6627 6990 6667 8310
rect 5267 6950 6667 6990
rect 6986 8310 8386 8350
rect 6986 6990 7026 8310
rect 8346 6990 8386 8310
rect 6986 6950 8386 6990
rect 8705 8310 10105 8350
rect 8705 6990 8745 8310
rect 10065 6990 10105 8310
rect 8705 6950 10105 6990
rect 10424 8310 11824 8350
rect 10424 6990 10464 8310
rect 11784 6990 11824 8310
rect 10424 6950 11824 6990
rect 12143 8310 13543 8350
rect 12143 6990 12183 8310
rect 13503 6990 13543 8310
rect 12143 6950 13543 6990
rect 13862 8310 15262 8350
rect 13862 6990 13902 8310
rect 15222 6990 15262 8310
rect 13862 6950 15262 6990
rect -15361 6610 -13961 6650
rect -15361 5290 -15321 6610
rect -14001 5290 -13961 6610
rect -15361 5250 -13961 5290
rect -13642 6610 -12242 6650
rect -13642 5290 -13602 6610
rect -12282 5290 -12242 6610
rect -13642 5250 -12242 5290
rect -11923 6610 -10523 6650
rect -11923 5290 -11883 6610
rect -10563 5290 -10523 6610
rect -11923 5250 -10523 5290
rect -10204 6610 -8804 6650
rect -10204 5290 -10164 6610
rect -8844 5290 -8804 6610
rect -10204 5250 -8804 5290
rect -8485 6610 -7085 6650
rect -8485 5290 -8445 6610
rect -7125 5290 -7085 6610
rect -8485 5250 -7085 5290
rect -6766 6610 -5366 6650
rect -6766 5290 -6726 6610
rect -5406 5290 -5366 6610
rect -6766 5250 -5366 5290
rect -5047 6610 -3647 6650
rect -5047 5290 -5007 6610
rect -3687 5290 -3647 6610
rect -5047 5250 -3647 5290
rect -3328 6610 -1928 6650
rect -3328 5290 -3288 6610
rect -1968 5290 -1928 6610
rect -3328 5250 -1928 5290
rect -1609 6610 -209 6650
rect -1609 5290 -1569 6610
rect -249 5290 -209 6610
rect -1609 5250 -209 5290
rect 110 6610 1510 6650
rect 110 5290 150 6610
rect 1470 5290 1510 6610
rect 110 5250 1510 5290
rect 1829 6610 3229 6650
rect 1829 5290 1869 6610
rect 3189 5290 3229 6610
rect 1829 5250 3229 5290
rect 3548 6610 4948 6650
rect 3548 5290 3588 6610
rect 4908 5290 4948 6610
rect 3548 5250 4948 5290
rect 5267 6610 6667 6650
rect 5267 5290 5307 6610
rect 6627 5290 6667 6610
rect 5267 5250 6667 5290
rect 6986 6610 8386 6650
rect 6986 5290 7026 6610
rect 8346 5290 8386 6610
rect 6986 5250 8386 5290
rect 8705 6610 10105 6650
rect 8705 5290 8745 6610
rect 10065 5290 10105 6610
rect 8705 5250 10105 5290
rect 10424 6610 11824 6650
rect 10424 5290 10464 6610
rect 11784 5290 11824 6610
rect 10424 5250 11824 5290
rect 12143 6610 13543 6650
rect 12143 5290 12183 6610
rect 13503 5290 13543 6610
rect 12143 5250 13543 5290
rect 13862 6610 15262 6650
rect 13862 5290 13902 6610
rect 15222 5290 15262 6610
rect 13862 5250 15262 5290
rect -15361 4910 -13961 4950
rect -15361 3590 -15321 4910
rect -14001 3590 -13961 4910
rect -15361 3550 -13961 3590
rect -13642 4910 -12242 4950
rect -13642 3590 -13602 4910
rect -12282 3590 -12242 4910
rect -13642 3550 -12242 3590
rect -11923 4910 -10523 4950
rect -11923 3590 -11883 4910
rect -10563 3590 -10523 4910
rect -11923 3550 -10523 3590
rect -10204 4910 -8804 4950
rect -10204 3590 -10164 4910
rect -8844 3590 -8804 4910
rect -10204 3550 -8804 3590
rect -8485 4910 -7085 4950
rect -8485 3590 -8445 4910
rect -7125 3590 -7085 4910
rect -8485 3550 -7085 3590
rect -6766 4910 -5366 4950
rect -6766 3590 -6726 4910
rect -5406 3590 -5366 4910
rect -6766 3550 -5366 3590
rect -5047 4910 -3647 4950
rect -5047 3590 -5007 4910
rect -3687 3590 -3647 4910
rect -5047 3550 -3647 3590
rect -3328 4910 -1928 4950
rect -3328 3590 -3288 4910
rect -1968 3590 -1928 4910
rect -3328 3550 -1928 3590
rect -1609 4910 -209 4950
rect -1609 3590 -1569 4910
rect -249 3590 -209 4910
rect -1609 3550 -209 3590
rect 110 4910 1510 4950
rect 110 3590 150 4910
rect 1470 3590 1510 4910
rect 110 3550 1510 3590
rect 1829 4910 3229 4950
rect 1829 3590 1869 4910
rect 3189 3590 3229 4910
rect 1829 3550 3229 3590
rect 3548 4910 4948 4950
rect 3548 3590 3588 4910
rect 4908 3590 4948 4910
rect 3548 3550 4948 3590
rect 5267 4910 6667 4950
rect 5267 3590 5307 4910
rect 6627 3590 6667 4910
rect 5267 3550 6667 3590
rect 6986 4910 8386 4950
rect 6986 3590 7026 4910
rect 8346 3590 8386 4910
rect 6986 3550 8386 3590
rect 8705 4910 10105 4950
rect 8705 3590 8745 4910
rect 10065 3590 10105 4910
rect 8705 3550 10105 3590
rect 10424 4910 11824 4950
rect 10424 3590 10464 4910
rect 11784 3590 11824 4910
rect 10424 3550 11824 3590
rect 12143 4910 13543 4950
rect 12143 3590 12183 4910
rect 13503 3590 13543 4910
rect 12143 3550 13543 3590
rect 13862 4910 15262 4950
rect 13862 3590 13902 4910
rect 15222 3590 15262 4910
rect 13862 3550 15262 3590
rect -15361 3210 -13961 3250
rect -15361 1890 -15321 3210
rect -14001 1890 -13961 3210
rect -15361 1850 -13961 1890
rect -13642 3210 -12242 3250
rect -13642 1890 -13602 3210
rect -12282 1890 -12242 3210
rect -13642 1850 -12242 1890
rect -11923 3210 -10523 3250
rect -11923 1890 -11883 3210
rect -10563 1890 -10523 3210
rect -11923 1850 -10523 1890
rect -10204 3210 -8804 3250
rect -10204 1890 -10164 3210
rect -8844 1890 -8804 3210
rect -10204 1850 -8804 1890
rect -8485 3210 -7085 3250
rect -8485 1890 -8445 3210
rect -7125 1890 -7085 3210
rect -8485 1850 -7085 1890
rect -6766 3210 -5366 3250
rect -6766 1890 -6726 3210
rect -5406 1890 -5366 3210
rect -6766 1850 -5366 1890
rect -5047 3210 -3647 3250
rect -5047 1890 -5007 3210
rect -3687 1890 -3647 3210
rect -5047 1850 -3647 1890
rect -3328 3210 -1928 3250
rect -3328 1890 -3288 3210
rect -1968 1890 -1928 3210
rect -3328 1850 -1928 1890
rect -1609 3210 -209 3250
rect -1609 1890 -1569 3210
rect -249 1890 -209 3210
rect -1609 1850 -209 1890
rect 110 3210 1510 3250
rect 110 1890 150 3210
rect 1470 1890 1510 3210
rect 110 1850 1510 1890
rect 1829 3210 3229 3250
rect 1829 1890 1869 3210
rect 3189 1890 3229 3210
rect 1829 1850 3229 1890
rect 3548 3210 4948 3250
rect 3548 1890 3588 3210
rect 4908 1890 4948 3210
rect 3548 1850 4948 1890
rect 5267 3210 6667 3250
rect 5267 1890 5307 3210
rect 6627 1890 6667 3210
rect 5267 1850 6667 1890
rect 6986 3210 8386 3250
rect 6986 1890 7026 3210
rect 8346 1890 8386 3210
rect 6986 1850 8386 1890
rect 8705 3210 10105 3250
rect 8705 1890 8745 3210
rect 10065 1890 10105 3210
rect 8705 1850 10105 1890
rect 10424 3210 11824 3250
rect 10424 1890 10464 3210
rect 11784 1890 11824 3210
rect 10424 1850 11824 1890
rect 12143 3210 13543 3250
rect 12143 1890 12183 3210
rect 13503 1890 13543 3210
rect 12143 1850 13543 1890
rect 13862 3210 15262 3250
rect 13862 1890 13902 3210
rect 15222 1890 15262 3210
rect 13862 1850 15262 1890
rect -15361 1510 -13961 1550
rect -15361 190 -15321 1510
rect -14001 190 -13961 1510
rect -15361 150 -13961 190
rect -13642 1510 -12242 1550
rect -13642 190 -13602 1510
rect -12282 190 -12242 1510
rect -13642 150 -12242 190
rect -11923 1510 -10523 1550
rect -11923 190 -11883 1510
rect -10563 190 -10523 1510
rect -11923 150 -10523 190
rect -10204 1510 -8804 1550
rect -10204 190 -10164 1510
rect -8844 190 -8804 1510
rect -10204 150 -8804 190
rect -8485 1510 -7085 1550
rect -8485 190 -8445 1510
rect -7125 190 -7085 1510
rect -8485 150 -7085 190
rect -6766 1510 -5366 1550
rect -6766 190 -6726 1510
rect -5406 190 -5366 1510
rect -6766 150 -5366 190
rect -5047 1510 -3647 1550
rect -5047 190 -5007 1510
rect -3687 190 -3647 1510
rect -5047 150 -3647 190
rect -3328 1510 -1928 1550
rect -3328 190 -3288 1510
rect -1968 190 -1928 1510
rect -3328 150 -1928 190
rect -1609 1510 -209 1550
rect -1609 190 -1569 1510
rect -249 190 -209 1510
rect -1609 150 -209 190
rect 110 1510 1510 1550
rect 110 190 150 1510
rect 1470 190 1510 1510
rect 110 150 1510 190
rect 1829 1510 3229 1550
rect 1829 190 1869 1510
rect 3189 190 3229 1510
rect 1829 150 3229 190
rect 3548 1510 4948 1550
rect 3548 190 3588 1510
rect 4908 190 4948 1510
rect 3548 150 4948 190
rect 5267 1510 6667 1550
rect 5267 190 5307 1510
rect 6627 190 6667 1510
rect 5267 150 6667 190
rect 6986 1510 8386 1550
rect 6986 190 7026 1510
rect 8346 190 8386 1510
rect 6986 150 8386 190
rect 8705 1510 10105 1550
rect 8705 190 8745 1510
rect 10065 190 10105 1510
rect 8705 150 10105 190
rect 10424 1510 11824 1550
rect 10424 190 10464 1510
rect 11784 190 11824 1510
rect 10424 150 11824 190
rect 12143 1510 13543 1550
rect 12143 190 12183 1510
rect 13503 190 13543 1510
rect 12143 150 13543 190
rect 13862 1510 15262 1550
rect 13862 190 13902 1510
rect 15222 190 15262 1510
rect 13862 150 15262 190
rect -15361 -190 -13961 -150
rect -15361 -1510 -15321 -190
rect -14001 -1510 -13961 -190
rect -15361 -1550 -13961 -1510
rect -13642 -190 -12242 -150
rect -13642 -1510 -13602 -190
rect -12282 -1510 -12242 -190
rect -13642 -1550 -12242 -1510
rect -11923 -190 -10523 -150
rect -11923 -1510 -11883 -190
rect -10563 -1510 -10523 -190
rect -11923 -1550 -10523 -1510
rect -10204 -190 -8804 -150
rect -10204 -1510 -10164 -190
rect -8844 -1510 -8804 -190
rect -10204 -1550 -8804 -1510
rect -8485 -190 -7085 -150
rect -8485 -1510 -8445 -190
rect -7125 -1510 -7085 -190
rect -8485 -1550 -7085 -1510
rect -6766 -190 -5366 -150
rect -6766 -1510 -6726 -190
rect -5406 -1510 -5366 -190
rect -6766 -1550 -5366 -1510
rect -5047 -190 -3647 -150
rect -5047 -1510 -5007 -190
rect -3687 -1510 -3647 -190
rect -5047 -1550 -3647 -1510
rect -3328 -190 -1928 -150
rect -3328 -1510 -3288 -190
rect -1968 -1510 -1928 -190
rect -3328 -1550 -1928 -1510
rect -1609 -190 -209 -150
rect -1609 -1510 -1569 -190
rect -249 -1510 -209 -190
rect -1609 -1550 -209 -1510
rect 110 -190 1510 -150
rect 110 -1510 150 -190
rect 1470 -1510 1510 -190
rect 110 -1550 1510 -1510
rect 1829 -190 3229 -150
rect 1829 -1510 1869 -190
rect 3189 -1510 3229 -190
rect 1829 -1550 3229 -1510
rect 3548 -190 4948 -150
rect 3548 -1510 3588 -190
rect 4908 -1510 4948 -190
rect 3548 -1550 4948 -1510
rect 5267 -190 6667 -150
rect 5267 -1510 5307 -190
rect 6627 -1510 6667 -190
rect 5267 -1550 6667 -1510
rect 6986 -190 8386 -150
rect 6986 -1510 7026 -190
rect 8346 -1510 8386 -190
rect 6986 -1550 8386 -1510
rect 8705 -190 10105 -150
rect 8705 -1510 8745 -190
rect 10065 -1510 10105 -190
rect 8705 -1550 10105 -1510
rect 10424 -190 11824 -150
rect 10424 -1510 10464 -190
rect 11784 -1510 11824 -190
rect 10424 -1550 11824 -1510
rect 12143 -190 13543 -150
rect 12143 -1510 12183 -190
rect 13503 -1510 13543 -190
rect 12143 -1550 13543 -1510
rect 13862 -190 15262 -150
rect 13862 -1510 13902 -190
rect 15222 -1510 15262 -190
rect 13862 -1550 15262 -1510
rect -15361 -1890 -13961 -1850
rect -15361 -3210 -15321 -1890
rect -14001 -3210 -13961 -1890
rect -15361 -3250 -13961 -3210
rect -13642 -1890 -12242 -1850
rect -13642 -3210 -13602 -1890
rect -12282 -3210 -12242 -1890
rect -13642 -3250 -12242 -3210
rect -11923 -1890 -10523 -1850
rect -11923 -3210 -11883 -1890
rect -10563 -3210 -10523 -1890
rect -11923 -3250 -10523 -3210
rect -10204 -1890 -8804 -1850
rect -10204 -3210 -10164 -1890
rect -8844 -3210 -8804 -1890
rect -10204 -3250 -8804 -3210
rect -8485 -1890 -7085 -1850
rect -8485 -3210 -8445 -1890
rect -7125 -3210 -7085 -1890
rect -8485 -3250 -7085 -3210
rect -6766 -1890 -5366 -1850
rect -6766 -3210 -6726 -1890
rect -5406 -3210 -5366 -1890
rect -6766 -3250 -5366 -3210
rect -5047 -1890 -3647 -1850
rect -5047 -3210 -5007 -1890
rect -3687 -3210 -3647 -1890
rect -5047 -3250 -3647 -3210
rect -3328 -1890 -1928 -1850
rect -3328 -3210 -3288 -1890
rect -1968 -3210 -1928 -1890
rect -3328 -3250 -1928 -3210
rect -1609 -1890 -209 -1850
rect -1609 -3210 -1569 -1890
rect -249 -3210 -209 -1890
rect -1609 -3250 -209 -3210
rect 110 -1890 1510 -1850
rect 110 -3210 150 -1890
rect 1470 -3210 1510 -1890
rect 110 -3250 1510 -3210
rect 1829 -1890 3229 -1850
rect 1829 -3210 1869 -1890
rect 3189 -3210 3229 -1890
rect 1829 -3250 3229 -3210
rect 3548 -1890 4948 -1850
rect 3548 -3210 3588 -1890
rect 4908 -3210 4948 -1890
rect 3548 -3250 4948 -3210
rect 5267 -1890 6667 -1850
rect 5267 -3210 5307 -1890
rect 6627 -3210 6667 -1890
rect 5267 -3250 6667 -3210
rect 6986 -1890 8386 -1850
rect 6986 -3210 7026 -1890
rect 8346 -3210 8386 -1890
rect 6986 -3250 8386 -3210
rect 8705 -1890 10105 -1850
rect 8705 -3210 8745 -1890
rect 10065 -3210 10105 -1890
rect 8705 -3250 10105 -3210
rect 10424 -1890 11824 -1850
rect 10424 -3210 10464 -1890
rect 11784 -3210 11824 -1890
rect 10424 -3250 11824 -3210
rect 12143 -1890 13543 -1850
rect 12143 -3210 12183 -1890
rect 13503 -3210 13543 -1890
rect 12143 -3250 13543 -3210
rect 13862 -1890 15262 -1850
rect 13862 -3210 13902 -1890
rect 15222 -3210 15262 -1890
rect 13862 -3250 15262 -3210
rect -15361 -3590 -13961 -3550
rect -15361 -4910 -15321 -3590
rect -14001 -4910 -13961 -3590
rect -15361 -4950 -13961 -4910
rect -13642 -3590 -12242 -3550
rect -13642 -4910 -13602 -3590
rect -12282 -4910 -12242 -3590
rect -13642 -4950 -12242 -4910
rect -11923 -3590 -10523 -3550
rect -11923 -4910 -11883 -3590
rect -10563 -4910 -10523 -3590
rect -11923 -4950 -10523 -4910
rect -10204 -3590 -8804 -3550
rect -10204 -4910 -10164 -3590
rect -8844 -4910 -8804 -3590
rect -10204 -4950 -8804 -4910
rect -8485 -3590 -7085 -3550
rect -8485 -4910 -8445 -3590
rect -7125 -4910 -7085 -3590
rect -8485 -4950 -7085 -4910
rect -6766 -3590 -5366 -3550
rect -6766 -4910 -6726 -3590
rect -5406 -4910 -5366 -3590
rect -6766 -4950 -5366 -4910
rect -5047 -3590 -3647 -3550
rect -5047 -4910 -5007 -3590
rect -3687 -4910 -3647 -3590
rect -5047 -4950 -3647 -4910
rect -3328 -3590 -1928 -3550
rect -3328 -4910 -3288 -3590
rect -1968 -4910 -1928 -3590
rect -3328 -4950 -1928 -4910
rect -1609 -3590 -209 -3550
rect -1609 -4910 -1569 -3590
rect -249 -4910 -209 -3590
rect -1609 -4950 -209 -4910
rect 110 -3590 1510 -3550
rect 110 -4910 150 -3590
rect 1470 -4910 1510 -3590
rect 110 -4950 1510 -4910
rect 1829 -3590 3229 -3550
rect 1829 -4910 1869 -3590
rect 3189 -4910 3229 -3590
rect 1829 -4950 3229 -4910
rect 3548 -3590 4948 -3550
rect 3548 -4910 3588 -3590
rect 4908 -4910 4948 -3590
rect 3548 -4950 4948 -4910
rect 5267 -3590 6667 -3550
rect 5267 -4910 5307 -3590
rect 6627 -4910 6667 -3590
rect 5267 -4950 6667 -4910
rect 6986 -3590 8386 -3550
rect 6986 -4910 7026 -3590
rect 8346 -4910 8386 -3590
rect 6986 -4950 8386 -4910
rect 8705 -3590 10105 -3550
rect 8705 -4910 8745 -3590
rect 10065 -4910 10105 -3590
rect 8705 -4950 10105 -4910
rect 10424 -3590 11824 -3550
rect 10424 -4910 10464 -3590
rect 11784 -4910 11824 -3590
rect 10424 -4950 11824 -4910
rect 12143 -3590 13543 -3550
rect 12143 -4910 12183 -3590
rect 13503 -4910 13543 -3590
rect 12143 -4950 13543 -4910
rect 13862 -3590 15262 -3550
rect 13862 -4910 13902 -3590
rect 15222 -4910 15262 -3590
rect 13862 -4950 15262 -4910
rect -15361 -5290 -13961 -5250
rect -15361 -6610 -15321 -5290
rect -14001 -6610 -13961 -5290
rect -15361 -6650 -13961 -6610
rect -13642 -5290 -12242 -5250
rect -13642 -6610 -13602 -5290
rect -12282 -6610 -12242 -5290
rect -13642 -6650 -12242 -6610
rect -11923 -5290 -10523 -5250
rect -11923 -6610 -11883 -5290
rect -10563 -6610 -10523 -5290
rect -11923 -6650 -10523 -6610
rect -10204 -5290 -8804 -5250
rect -10204 -6610 -10164 -5290
rect -8844 -6610 -8804 -5290
rect -10204 -6650 -8804 -6610
rect -8485 -5290 -7085 -5250
rect -8485 -6610 -8445 -5290
rect -7125 -6610 -7085 -5290
rect -8485 -6650 -7085 -6610
rect -6766 -5290 -5366 -5250
rect -6766 -6610 -6726 -5290
rect -5406 -6610 -5366 -5290
rect -6766 -6650 -5366 -6610
rect -5047 -5290 -3647 -5250
rect -5047 -6610 -5007 -5290
rect -3687 -6610 -3647 -5290
rect -5047 -6650 -3647 -6610
rect -3328 -5290 -1928 -5250
rect -3328 -6610 -3288 -5290
rect -1968 -6610 -1928 -5290
rect -3328 -6650 -1928 -6610
rect -1609 -5290 -209 -5250
rect -1609 -6610 -1569 -5290
rect -249 -6610 -209 -5290
rect -1609 -6650 -209 -6610
rect 110 -5290 1510 -5250
rect 110 -6610 150 -5290
rect 1470 -6610 1510 -5290
rect 110 -6650 1510 -6610
rect 1829 -5290 3229 -5250
rect 1829 -6610 1869 -5290
rect 3189 -6610 3229 -5290
rect 1829 -6650 3229 -6610
rect 3548 -5290 4948 -5250
rect 3548 -6610 3588 -5290
rect 4908 -6610 4948 -5290
rect 3548 -6650 4948 -6610
rect 5267 -5290 6667 -5250
rect 5267 -6610 5307 -5290
rect 6627 -6610 6667 -5290
rect 5267 -6650 6667 -6610
rect 6986 -5290 8386 -5250
rect 6986 -6610 7026 -5290
rect 8346 -6610 8386 -5290
rect 6986 -6650 8386 -6610
rect 8705 -5290 10105 -5250
rect 8705 -6610 8745 -5290
rect 10065 -6610 10105 -5290
rect 8705 -6650 10105 -6610
rect 10424 -5290 11824 -5250
rect 10424 -6610 10464 -5290
rect 11784 -6610 11824 -5290
rect 10424 -6650 11824 -6610
rect 12143 -5290 13543 -5250
rect 12143 -6610 12183 -5290
rect 13503 -6610 13543 -5290
rect 12143 -6650 13543 -6610
rect 13862 -5290 15262 -5250
rect 13862 -6610 13902 -5290
rect 15222 -6610 15262 -5290
rect 13862 -6650 15262 -6610
rect -15361 -6990 -13961 -6950
rect -15361 -8310 -15321 -6990
rect -14001 -8310 -13961 -6990
rect -15361 -8350 -13961 -8310
rect -13642 -6990 -12242 -6950
rect -13642 -8310 -13602 -6990
rect -12282 -8310 -12242 -6990
rect -13642 -8350 -12242 -8310
rect -11923 -6990 -10523 -6950
rect -11923 -8310 -11883 -6990
rect -10563 -8310 -10523 -6990
rect -11923 -8350 -10523 -8310
rect -10204 -6990 -8804 -6950
rect -10204 -8310 -10164 -6990
rect -8844 -8310 -8804 -6990
rect -10204 -8350 -8804 -8310
rect -8485 -6990 -7085 -6950
rect -8485 -8310 -8445 -6990
rect -7125 -8310 -7085 -6990
rect -8485 -8350 -7085 -8310
rect -6766 -6990 -5366 -6950
rect -6766 -8310 -6726 -6990
rect -5406 -8310 -5366 -6990
rect -6766 -8350 -5366 -8310
rect -5047 -6990 -3647 -6950
rect -5047 -8310 -5007 -6990
rect -3687 -8310 -3647 -6990
rect -5047 -8350 -3647 -8310
rect -3328 -6990 -1928 -6950
rect -3328 -8310 -3288 -6990
rect -1968 -8310 -1928 -6990
rect -3328 -8350 -1928 -8310
rect -1609 -6990 -209 -6950
rect -1609 -8310 -1569 -6990
rect -249 -8310 -209 -6990
rect -1609 -8350 -209 -8310
rect 110 -6990 1510 -6950
rect 110 -8310 150 -6990
rect 1470 -8310 1510 -6990
rect 110 -8350 1510 -8310
rect 1829 -6990 3229 -6950
rect 1829 -8310 1869 -6990
rect 3189 -8310 3229 -6990
rect 1829 -8350 3229 -8310
rect 3548 -6990 4948 -6950
rect 3548 -8310 3588 -6990
rect 4908 -8310 4948 -6990
rect 3548 -8350 4948 -8310
rect 5267 -6990 6667 -6950
rect 5267 -8310 5307 -6990
rect 6627 -8310 6667 -6990
rect 5267 -8350 6667 -8310
rect 6986 -6990 8386 -6950
rect 6986 -8310 7026 -6990
rect 8346 -8310 8386 -6990
rect 6986 -8350 8386 -8310
rect 8705 -6990 10105 -6950
rect 8705 -8310 8745 -6990
rect 10065 -8310 10105 -6990
rect 8705 -8350 10105 -8310
rect 10424 -6990 11824 -6950
rect 10424 -8310 10464 -6990
rect 11784 -8310 11824 -6990
rect 10424 -8350 11824 -8310
rect 12143 -6990 13543 -6950
rect 12143 -8310 12183 -6990
rect 13503 -8310 13543 -6990
rect 12143 -8350 13543 -8310
rect 13862 -6990 15262 -6950
rect 13862 -8310 13902 -6990
rect 15222 -8310 15262 -6990
rect 13862 -8350 15262 -8310
rect -15361 -8690 -13961 -8650
rect -15361 -10010 -15321 -8690
rect -14001 -10010 -13961 -8690
rect -15361 -10050 -13961 -10010
rect -13642 -8690 -12242 -8650
rect -13642 -10010 -13602 -8690
rect -12282 -10010 -12242 -8690
rect -13642 -10050 -12242 -10010
rect -11923 -8690 -10523 -8650
rect -11923 -10010 -11883 -8690
rect -10563 -10010 -10523 -8690
rect -11923 -10050 -10523 -10010
rect -10204 -8690 -8804 -8650
rect -10204 -10010 -10164 -8690
rect -8844 -10010 -8804 -8690
rect -10204 -10050 -8804 -10010
rect -8485 -8690 -7085 -8650
rect -8485 -10010 -8445 -8690
rect -7125 -10010 -7085 -8690
rect -8485 -10050 -7085 -10010
rect -6766 -8690 -5366 -8650
rect -6766 -10010 -6726 -8690
rect -5406 -10010 -5366 -8690
rect -6766 -10050 -5366 -10010
rect -5047 -8690 -3647 -8650
rect -5047 -10010 -5007 -8690
rect -3687 -10010 -3647 -8690
rect -5047 -10050 -3647 -10010
rect -3328 -8690 -1928 -8650
rect -3328 -10010 -3288 -8690
rect -1968 -10010 -1928 -8690
rect -3328 -10050 -1928 -10010
rect -1609 -8690 -209 -8650
rect -1609 -10010 -1569 -8690
rect -249 -10010 -209 -8690
rect -1609 -10050 -209 -10010
rect 110 -8690 1510 -8650
rect 110 -10010 150 -8690
rect 1470 -10010 1510 -8690
rect 110 -10050 1510 -10010
rect 1829 -8690 3229 -8650
rect 1829 -10010 1869 -8690
rect 3189 -10010 3229 -8690
rect 1829 -10050 3229 -10010
rect 3548 -8690 4948 -8650
rect 3548 -10010 3588 -8690
rect 4908 -10010 4948 -8690
rect 3548 -10050 4948 -10010
rect 5267 -8690 6667 -8650
rect 5267 -10010 5307 -8690
rect 6627 -10010 6667 -8690
rect 5267 -10050 6667 -10010
rect 6986 -8690 8386 -8650
rect 6986 -10010 7026 -8690
rect 8346 -10010 8386 -8690
rect 6986 -10050 8386 -10010
rect 8705 -8690 10105 -8650
rect 8705 -10010 8745 -8690
rect 10065 -10010 10105 -8690
rect 8705 -10050 10105 -10010
rect 10424 -8690 11824 -8650
rect 10424 -10010 10464 -8690
rect 11784 -10010 11824 -8690
rect 10424 -10050 11824 -10010
rect 12143 -8690 13543 -8650
rect 12143 -10010 12183 -8690
rect 13503 -10010 13543 -8690
rect 12143 -10050 13543 -10010
rect 13862 -8690 15262 -8650
rect 13862 -10010 13902 -8690
rect 15222 -10010 15262 -8690
rect 13862 -10050 15262 -10010
rect -15361 -10390 -13961 -10350
rect -15361 -11710 -15321 -10390
rect -14001 -11710 -13961 -10390
rect -15361 -11750 -13961 -11710
rect -13642 -10390 -12242 -10350
rect -13642 -11710 -13602 -10390
rect -12282 -11710 -12242 -10390
rect -13642 -11750 -12242 -11710
rect -11923 -10390 -10523 -10350
rect -11923 -11710 -11883 -10390
rect -10563 -11710 -10523 -10390
rect -11923 -11750 -10523 -11710
rect -10204 -10390 -8804 -10350
rect -10204 -11710 -10164 -10390
rect -8844 -11710 -8804 -10390
rect -10204 -11750 -8804 -11710
rect -8485 -10390 -7085 -10350
rect -8485 -11710 -8445 -10390
rect -7125 -11710 -7085 -10390
rect -8485 -11750 -7085 -11710
rect -6766 -10390 -5366 -10350
rect -6766 -11710 -6726 -10390
rect -5406 -11710 -5366 -10390
rect -6766 -11750 -5366 -11710
rect -5047 -10390 -3647 -10350
rect -5047 -11710 -5007 -10390
rect -3687 -11710 -3647 -10390
rect -5047 -11750 -3647 -11710
rect -3328 -10390 -1928 -10350
rect -3328 -11710 -3288 -10390
rect -1968 -11710 -1928 -10390
rect -3328 -11750 -1928 -11710
rect -1609 -10390 -209 -10350
rect -1609 -11710 -1569 -10390
rect -249 -11710 -209 -10390
rect -1609 -11750 -209 -11710
rect 110 -10390 1510 -10350
rect 110 -11710 150 -10390
rect 1470 -11710 1510 -10390
rect 110 -11750 1510 -11710
rect 1829 -10390 3229 -10350
rect 1829 -11710 1869 -10390
rect 3189 -11710 3229 -10390
rect 1829 -11750 3229 -11710
rect 3548 -10390 4948 -10350
rect 3548 -11710 3588 -10390
rect 4908 -11710 4948 -10390
rect 3548 -11750 4948 -11710
rect 5267 -10390 6667 -10350
rect 5267 -11710 5307 -10390
rect 6627 -11710 6667 -10390
rect 5267 -11750 6667 -11710
rect 6986 -10390 8386 -10350
rect 6986 -11710 7026 -10390
rect 8346 -11710 8386 -10390
rect 6986 -11750 8386 -11710
rect 8705 -10390 10105 -10350
rect 8705 -11710 8745 -10390
rect 10065 -11710 10105 -10390
rect 8705 -11750 10105 -11710
rect 10424 -10390 11824 -10350
rect 10424 -11710 10464 -10390
rect 11784 -11710 11824 -10390
rect 10424 -11750 11824 -11710
rect 12143 -10390 13543 -10350
rect 12143 -11710 12183 -10390
rect 13503 -11710 13543 -10390
rect 12143 -11750 13543 -11710
rect 13862 -10390 15262 -10350
rect 13862 -11710 13902 -10390
rect 15222 -11710 15262 -10390
rect 13862 -11750 15262 -11710
rect -15361 -12090 -13961 -12050
rect -15361 -13410 -15321 -12090
rect -14001 -13410 -13961 -12090
rect -15361 -13450 -13961 -13410
rect -13642 -12090 -12242 -12050
rect -13642 -13410 -13602 -12090
rect -12282 -13410 -12242 -12090
rect -13642 -13450 -12242 -13410
rect -11923 -12090 -10523 -12050
rect -11923 -13410 -11883 -12090
rect -10563 -13410 -10523 -12090
rect -11923 -13450 -10523 -13410
rect -10204 -12090 -8804 -12050
rect -10204 -13410 -10164 -12090
rect -8844 -13410 -8804 -12090
rect -10204 -13450 -8804 -13410
rect -8485 -12090 -7085 -12050
rect -8485 -13410 -8445 -12090
rect -7125 -13410 -7085 -12090
rect -8485 -13450 -7085 -13410
rect -6766 -12090 -5366 -12050
rect -6766 -13410 -6726 -12090
rect -5406 -13410 -5366 -12090
rect -6766 -13450 -5366 -13410
rect -5047 -12090 -3647 -12050
rect -5047 -13410 -5007 -12090
rect -3687 -13410 -3647 -12090
rect -5047 -13450 -3647 -13410
rect -3328 -12090 -1928 -12050
rect -3328 -13410 -3288 -12090
rect -1968 -13410 -1928 -12090
rect -3328 -13450 -1928 -13410
rect -1609 -12090 -209 -12050
rect -1609 -13410 -1569 -12090
rect -249 -13410 -209 -12090
rect -1609 -13450 -209 -13410
rect 110 -12090 1510 -12050
rect 110 -13410 150 -12090
rect 1470 -13410 1510 -12090
rect 110 -13450 1510 -13410
rect 1829 -12090 3229 -12050
rect 1829 -13410 1869 -12090
rect 3189 -13410 3229 -12090
rect 1829 -13450 3229 -13410
rect 3548 -12090 4948 -12050
rect 3548 -13410 3588 -12090
rect 4908 -13410 4948 -12090
rect 3548 -13450 4948 -13410
rect 5267 -12090 6667 -12050
rect 5267 -13410 5307 -12090
rect 6627 -13410 6667 -12090
rect 5267 -13450 6667 -13410
rect 6986 -12090 8386 -12050
rect 6986 -13410 7026 -12090
rect 8346 -13410 8386 -12090
rect 6986 -13450 8386 -13410
rect 8705 -12090 10105 -12050
rect 8705 -13410 8745 -12090
rect 10065 -13410 10105 -12090
rect 8705 -13450 10105 -13410
rect 10424 -12090 11824 -12050
rect 10424 -13410 10464 -12090
rect 11784 -13410 11824 -12090
rect 10424 -13450 11824 -13410
rect 12143 -12090 13543 -12050
rect 12143 -13410 12183 -12090
rect 13503 -13410 13543 -12090
rect 12143 -13450 13543 -13410
rect 13862 -12090 15262 -12050
rect 13862 -13410 13902 -12090
rect 15222 -13410 15262 -12090
rect 13862 -13450 15262 -13410
rect -15361 -13790 -13961 -13750
rect -15361 -15110 -15321 -13790
rect -14001 -15110 -13961 -13790
rect -15361 -15150 -13961 -15110
rect -13642 -13790 -12242 -13750
rect -13642 -15110 -13602 -13790
rect -12282 -15110 -12242 -13790
rect -13642 -15150 -12242 -15110
rect -11923 -13790 -10523 -13750
rect -11923 -15110 -11883 -13790
rect -10563 -15110 -10523 -13790
rect -11923 -15150 -10523 -15110
rect -10204 -13790 -8804 -13750
rect -10204 -15110 -10164 -13790
rect -8844 -15110 -8804 -13790
rect -10204 -15150 -8804 -15110
rect -8485 -13790 -7085 -13750
rect -8485 -15110 -8445 -13790
rect -7125 -15110 -7085 -13790
rect -8485 -15150 -7085 -15110
rect -6766 -13790 -5366 -13750
rect -6766 -15110 -6726 -13790
rect -5406 -15110 -5366 -13790
rect -6766 -15150 -5366 -15110
rect -5047 -13790 -3647 -13750
rect -5047 -15110 -5007 -13790
rect -3687 -15110 -3647 -13790
rect -5047 -15150 -3647 -15110
rect -3328 -13790 -1928 -13750
rect -3328 -15110 -3288 -13790
rect -1968 -15110 -1928 -13790
rect -3328 -15150 -1928 -15110
rect -1609 -13790 -209 -13750
rect -1609 -15110 -1569 -13790
rect -249 -15110 -209 -13790
rect -1609 -15150 -209 -15110
rect 110 -13790 1510 -13750
rect 110 -15110 150 -13790
rect 1470 -15110 1510 -13790
rect 110 -15150 1510 -15110
rect 1829 -13790 3229 -13750
rect 1829 -15110 1869 -13790
rect 3189 -15110 3229 -13790
rect 1829 -15150 3229 -15110
rect 3548 -13790 4948 -13750
rect 3548 -15110 3588 -13790
rect 4908 -15110 4948 -13790
rect 3548 -15150 4948 -15110
rect 5267 -13790 6667 -13750
rect 5267 -15110 5307 -13790
rect 6627 -15110 6667 -13790
rect 5267 -15150 6667 -15110
rect 6986 -13790 8386 -13750
rect 6986 -15110 7026 -13790
rect 8346 -15110 8386 -13790
rect 6986 -15150 8386 -15110
rect 8705 -13790 10105 -13750
rect 8705 -15110 8745 -13790
rect 10065 -15110 10105 -13790
rect 8705 -15150 10105 -15110
rect 10424 -13790 11824 -13750
rect 10424 -15110 10464 -13790
rect 11784 -15110 11824 -13790
rect 10424 -15150 11824 -15110
rect 12143 -13790 13543 -13750
rect 12143 -15110 12183 -13790
rect 13503 -15110 13543 -13790
rect 12143 -15150 13543 -15110
rect 13862 -13790 15262 -13750
rect 13862 -15110 13902 -13790
rect 15222 -15110 15262 -13790
rect 13862 -15150 15262 -15110
<< mimcapcontact >>
rect -15321 13790 -14001 15110
rect -13602 13790 -12282 15110
rect -11883 13790 -10563 15110
rect -10164 13790 -8844 15110
rect -8445 13790 -7125 15110
rect -6726 13790 -5406 15110
rect -5007 13790 -3687 15110
rect -3288 13790 -1968 15110
rect -1569 13790 -249 15110
rect 150 13790 1470 15110
rect 1869 13790 3189 15110
rect 3588 13790 4908 15110
rect 5307 13790 6627 15110
rect 7026 13790 8346 15110
rect 8745 13790 10065 15110
rect 10464 13790 11784 15110
rect 12183 13790 13503 15110
rect 13902 13790 15222 15110
rect -15321 12090 -14001 13410
rect -13602 12090 -12282 13410
rect -11883 12090 -10563 13410
rect -10164 12090 -8844 13410
rect -8445 12090 -7125 13410
rect -6726 12090 -5406 13410
rect -5007 12090 -3687 13410
rect -3288 12090 -1968 13410
rect -1569 12090 -249 13410
rect 150 12090 1470 13410
rect 1869 12090 3189 13410
rect 3588 12090 4908 13410
rect 5307 12090 6627 13410
rect 7026 12090 8346 13410
rect 8745 12090 10065 13410
rect 10464 12090 11784 13410
rect 12183 12090 13503 13410
rect 13902 12090 15222 13410
rect -15321 10390 -14001 11710
rect -13602 10390 -12282 11710
rect -11883 10390 -10563 11710
rect -10164 10390 -8844 11710
rect -8445 10390 -7125 11710
rect -6726 10390 -5406 11710
rect -5007 10390 -3687 11710
rect -3288 10390 -1968 11710
rect -1569 10390 -249 11710
rect 150 10390 1470 11710
rect 1869 10390 3189 11710
rect 3588 10390 4908 11710
rect 5307 10390 6627 11710
rect 7026 10390 8346 11710
rect 8745 10390 10065 11710
rect 10464 10390 11784 11710
rect 12183 10390 13503 11710
rect 13902 10390 15222 11710
rect -15321 8690 -14001 10010
rect -13602 8690 -12282 10010
rect -11883 8690 -10563 10010
rect -10164 8690 -8844 10010
rect -8445 8690 -7125 10010
rect -6726 8690 -5406 10010
rect -5007 8690 -3687 10010
rect -3288 8690 -1968 10010
rect -1569 8690 -249 10010
rect 150 8690 1470 10010
rect 1869 8690 3189 10010
rect 3588 8690 4908 10010
rect 5307 8690 6627 10010
rect 7026 8690 8346 10010
rect 8745 8690 10065 10010
rect 10464 8690 11784 10010
rect 12183 8690 13503 10010
rect 13902 8690 15222 10010
rect -15321 6990 -14001 8310
rect -13602 6990 -12282 8310
rect -11883 6990 -10563 8310
rect -10164 6990 -8844 8310
rect -8445 6990 -7125 8310
rect -6726 6990 -5406 8310
rect -5007 6990 -3687 8310
rect -3288 6990 -1968 8310
rect -1569 6990 -249 8310
rect 150 6990 1470 8310
rect 1869 6990 3189 8310
rect 3588 6990 4908 8310
rect 5307 6990 6627 8310
rect 7026 6990 8346 8310
rect 8745 6990 10065 8310
rect 10464 6990 11784 8310
rect 12183 6990 13503 8310
rect 13902 6990 15222 8310
rect -15321 5290 -14001 6610
rect -13602 5290 -12282 6610
rect -11883 5290 -10563 6610
rect -10164 5290 -8844 6610
rect -8445 5290 -7125 6610
rect -6726 5290 -5406 6610
rect -5007 5290 -3687 6610
rect -3288 5290 -1968 6610
rect -1569 5290 -249 6610
rect 150 5290 1470 6610
rect 1869 5290 3189 6610
rect 3588 5290 4908 6610
rect 5307 5290 6627 6610
rect 7026 5290 8346 6610
rect 8745 5290 10065 6610
rect 10464 5290 11784 6610
rect 12183 5290 13503 6610
rect 13902 5290 15222 6610
rect -15321 3590 -14001 4910
rect -13602 3590 -12282 4910
rect -11883 3590 -10563 4910
rect -10164 3590 -8844 4910
rect -8445 3590 -7125 4910
rect -6726 3590 -5406 4910
rect -5007 3590 -3687 4910
rect -3288 3590 -1968 4910
rect -1569 3590 -249 4910
rect 150 3590 1470 4910
rect 1869 3590 3189 4910
rect 3588 3590 4908 4910
rect 5307 3590 6627 4910
rect 7026 3590 8346 4910
rect 8745 3590 10065 4910
rect 10464 3590 11784 4910
rect 12183 3590 13503 4910
rect 13902 3590 15222 4910
rect -15321 1890 -14001 3210
rect -13602 1890 -12282 3210
rect -11883 1890 -10563 3210
rect -10164 1890 -8844 3210
rect -8445 1890 -7125 3210
rect -6726 1890 -5406 3210
rect -5007 1890 -3687 3210
rect -3288 1890 -1968 3210
rect -1569 1890 -249 3210
rect 150 1890 1470 3210
rect 1869 1890 3189 3210
rect 3588 1890 4908 3210
rect 5307 1890 6627 3210
rect 7026 1890 8346 3210
rect 8745 1890 10065 3210
rect 10464 1890 11784 3210
rect 12183 1890 13503 3210
rect 13902 1890 15222 3210
rect -15321 190 -14001 1510
rect -13602 190 -12282 1510
rect -11883 190 -10563 1510
rect -10164 190 -8844 1510
rect -8445 190 -7125 1510
rect -6726 190 -5406 1510
rect -5007 190 -3687 1510
rect -3288 190 -1968 1510
rect -1569 190 -249 1510
rect 150 190 1470 1510
rect 1869 190 3189 1510
rect 3588 190 4908 1510
rect 5307 190 6627 1510
rect 7026 190 8346 1510
rect 8745 190 10065 1510
rect 10464 190 11784 1510
rect 12183 190 13503 1510
rect 13902 190 15222 1510
rect -15321 -1510 -14001 -190
rect -13602 -1510 -12282 -190
rect -11883 -1510 -10563 -190
rect -10164 -1510 -8844 -190
rect -8445 -1510 -7125 -190
rect -6726 -1510 -5406 -190
rect -5007 -1510 -3687 -190
rect -3288 -1510 -1968 -190
rect -1569 -1510 -249 -190
rect 150 -1510 1470 -190
rect 1869 -1510 3189 -190
rect 3588 -1510 4908 -190
rect 5307 -1510 6627 -190
rect 7026 -1510 8346 -190
rect 8745 -1510 10065 -190
rect 10464 -1510 11784 -190
rect 12183 -1510 13503 -190
rect 13902 -1510 15222 -190
rect -15321 -3210 -14001 -1890
rect -13602 -3210 -12282 -1890
rect -11883 -3210 -10563 -1890
rect -10164 -3210 -8844 -1890
rect -8445 -3210 -7125 -1890
rect -6726 -3210 -5406 -1890
rect -5007 -3210 -3687 -1890
rect -3288 -3210 -1968 -1890
rect -1569 -3210 -249 -1890
rect 150 -3210 1470 -1890
rect 1869 -3210 3189 -1890
rect 3588 -3210 4908 -1890
rect 5307 -3210 6627 -1890
rect 7026 -3210 8346 -1890
rect 8745 -3210 10065 -1890
rect 10464 -3210 11784 -1890
rect 12183 -3210 13503 -1890
rect 13902 -3210 15222 -1890
rect -15321 -4910 -14001 -3590
rect -13602 -4910 -12282 -3590
rect -11883 -4910 -10563 -3590
rect -10164 -4910 -8844 -3590
rect -8445 -4910 -7125 -3590
rect -6726 -4910 -5406 -3590
rect -5007 -4910 -3687 -3590
rect -3288 -4910 -1968 -3590
rect -1569 -4910 -249 -3590
rect 150 -4910 1470 -3590
rect 1869 -4910 3189 -3590
rect 3588 -4910 4908 -3590
rect 5307 -4910 6627 -3590
rect 7026 -4910 8346 -3590
rect 8745 -4910 10065 -3590
rect 10464 -4910 11784 -3590
rect 12183 -4910 13503 -3590
rect 13902 -4910 15222 -3590
rect -15321 -6610 -14001 -5290
rect -13602 -6610 -12282 -5290
rect -11883 -6610 -10563 -5290
rect -10164 -6610 -8844 -5290
rect -8445 -6610 -7125 -5290
rect -6726 -6610 -5406 -5290
rect -5007 -6610 -3687 -5290
rect -3288 -6610 -1968 -5290
rect -1569 -6610 -249 -5290
rect 150 -6610 1470 -5290
rect 1869 -6610 3189 -5290
rect 3588 -6610 4908 -5290
rect 5307 -6610 6627 -5290
rect 7026 -6610 8346 -5290
rect 8745 -6610 10065 -5290
rect 10464 -6610 11784 -5290
rect 12183 -6610 13503 -5290
rect 13902 -6610 15222 -5290
rect -15321 -8310 -14001 -6990
rect -13602 -8310 -12282 -6990
rect -11883 -8310 -10563 -6990
rect -10164 -8310 -8844 -6990
rect -8445 -8310 -7125 -6990
rect -6726 -8310 -5406 -6990
rect -5007 -8310 -3687 -6990
rect -3288 -8310 -1968 -6990
rect -1569 -8310 -249 -6990
rect 150 -8310 1470 -6990
rect 1869 -8310 3189 -6990
rect 3588 -8310 4908 -6990
rect 5307 -8310 6627 -6990
rect 7026 -8310 8346 -6990
rect 8745 -8310 10065 -6990
rect 10464 -8310 11784 -6990
rect 12183 -8310 13503 -6990
rect 13902 -8310 15222 -6990
rect -15321 -10010 -14001 -8690
rect -13602 -10010 -12282 -8690
rect -11883 -10010 -10563 -8690
rect -10164 -10010 -8844 -8690
rect -8445 -10010 -7125 -8690
rect -6726 -10010 -5406 -8690
rect -5007 -10010 -3687 -8690
rect -3288 -10010 -1968 -8690
rect -1569 -10010 -249 -8690
rect 150 -10010 1470 -8690
rect 1869 -10010 3189 -8690
rect 3588 -10010 4908 -8690
rect 5307 -10010 6627 -8690
rect 7026 -10010 8346 -8690
rect 8745 -10010 10065 -8690
rect 10464 -10010 11784 -8690
rect 12183 -10010 13503 -8690
rect 13902 -10010 15222 -8690
rect -15321 -11710 -14001 -10390
rect -13602 -11710 -12282 -10390
rect -11883 -11710 -10563 -10390
rect -10164 -11710 -8844 -10390
rect -8445 -11710 -7125 -10390
rect -6726 -11710 -5406 -10390
rect -5007 -11710 -3687 -10390
rect -3288 -11710 -1968 -10390
rect -1569 -11710 -249 -10390
rect 150 -11710 1470 -10390
rect 1869 -11710 3189 -10390
rect 3588 -11710 4908 -10390
rect 5307 -11710 6627 -10390
rect 7026 -11710 8346 -10390
rect 8745 -11710 10065 -10390
rect 10464 -11710 11784 -10390
rect 12183 -11710 13503 -10390
rect 13902 -11710 15222 -10390
rect -15321 -13410 -14001 -12090
rect -13602 -13410 -12282 -12090
rect -11883 -13410 -10563 -12090
rect -10164 -13410 -8844 -12090
rect -8445 -13410 -7125 -12090
rect -6726 -13410 -5406 -12090
rect -5007 -13410 -3687 -12090
rect -3288 -13410 -1968 -12090
rect -1569 -13410 -249 -12090
rect 150 -13410 1470 -12090
rect 1869 -13410 3189 -12090
rect 3588 -13410 4908 -12090
rect 5307 -13410 6627 -12090
rect 7026 -13410 8346 -12090
rect 8745 -13410 10065 -12090
rect 10464 -13410 11784 -12090
rect 12183 -13410 13503 -12090
rect 13902 -13410 15222 -12090
rect -15321 -15110 -14001 -13790
rect -13602 -15110 -12282 -13790
rect -11883 -15110 -10563 -13790
rect -10164 -15110 -8844 -13790
rect -8445 -15110 -7125 -13790
rect -6726 -15110 -5406 -13790
rect -5007 -15110 -3687 -13790
rect -3288 -15110 -1968 -13790
rect -1569 -15110 -249 -13790
rect 150 -15110 1470 -13790
rect 1869 -15110 3189 -13790
rect 3588 -15110 4908 -13790
rect 5307 -15110 6627 -13790
rect 7026 -15110 8346 -13790
rect 8745 -15110 10065 -13790
rect 10464 -15110 11784 -13790
rect 12183 -15110 13503 -13790
rect 13902 -15110 15222 -13790
<< metal4 >>
rect -13862 15222 -13766 15238
rect -15322 15110 -14000 15111
rect -15322 13790 -15321 15110
rect -14001 13790 -14000 15110
rect -15322 13789 -14000 13790
rect -13862 13678 -13846 15222
rect -13782 13678 -13766 15222
rect -12143 15222 -12047 15238
rect -13603 15110 -12281 15111
rect -13603 13790 -13602 15110
rect -12282 13790 -12281 15110
rect -13603 13789 -12281 13790
rect -13862 13662 -13766 13678
rect -12143 13678 -12127 15222
rect -12063 13678 -12047 15222
rect -10424 15222 -10328 15238
rect -11884 15110 -10562 15111
rect -11884 13790 -11883 15110
rect -10563 13790 -10562 15110
rect -11884 13789 -10562 13790
rect -12143 13662 -12047 13678
rect -10424 13678 -10408 15222
rect -10344 13678 -10328 15222
rect -8705 15222 -8609 15238
rect -10165 15110 -8843 15111
rect -10165 13790 -10164 15110
rect -8844 13790 -8843 15110
rect -10165 13789 -8843 13790
rect -10424 13662 -10328 13678
rect -8705 13678 -8689 15222
rect -8625 13678 -8609 15222
rect -6986 15222 -6890 15238
rect -8446 15110 -7124 15111
rect -8446 13790 -8445 15110
rect -7125 13790 -7124 15110
rect -8446 13789 -7124 13790
rect -8705 13662 -8609 13678
rect -6986 13678 -6970 15222
rect -6906 13678 -6890 15222
rect -5267 15222 -5171 15238
rect -6727 15110 -5405 15111
rect -6727 13790 -6726 15110
rect -5406 13790 -5405 15110
rect -6727 13789 -5405 13790
rect -6986 13662 -6890 13678
rect -5267 13678 -5251 15222
rect -5187 13678 -5171 15222
rect -3548 15222 -3452 15238
rect -5008 15110 -3686 15111
rect -5008 13790 -5007 15110
rect -3687 13790 -3686 15110
rect -5008 13789 -3686 13790
rect -5267 13662 -5171 13678
rect -3548 13678 -3532 15222
rect -3468 13678 -3452 15222
rect -1829 15222 -1733 15238
rect -3289 15110 -1967 15111
rect -3289 13790 -3288 15110
rect -1968 13790 -1967 15110
rect -3289 13789 -1967 13790
rect -3548 13662 -3452 13678
rect -1829 13678 -1813 15222
rect -1749 13678 -1733 15222
rect -110 15222 -14 15238
rect -1570 15110 -248 15111
rect -1570 13790 -1569 15110
rect -249 13790 -248 15110
rect -1570 13789 -248 13790
rect -1829 13662 -1733 13678
rect -110 13678 -94 15222
rect -30 13678 -14 15222
rect 1609 15222 1705 15238
rect 149 15110 1471 15111
rect 149 13790 150 15110
rect 1470 13790 1471 15110
rect 149 13789 1471 13790
rect -110 13662 -14 13678
rect 1609 13678 1625 15222
rect 1689 13678 1705 15222
rect 3328 15222 3424 15238
rect 1868 15110 3190 15111
rect 1868 13790 1869 15110
rect 3189 13790 3190 15110
rect 1868 13789 3190 13790
rect 1609 13662 1705 13678
rect 3328 13678 3344 15222
rect 3408 13678 3424 15222
rect 5047 15222 5143 15238
rect 3587 15110 4909 15111
rect 3587 13790 3588 15110
rect 4908 13790 4909 15110
rect 3587 13789 4909 13790
rect 3328 13662 3424 13678
rect 5047 13678 5063 15222
rect 5127 13678 5143 15222
rect 6766 15222 6862 15238
rect 5306 15110 6628 15111
rect 5306 13790 5307 15110
rect 6627 13790 6628 15110
rect 5306 13789 6628 13790
rect 5047 13662 5143 13678
rect 6766 13678 6782 15222
rect 6846 13678 6862 15222
rect 8485 15222 8581 15238
rect 7025 15110 8347 15111
rect 7025 13790 7026 15110
rect 8346 13790 8347 15110
rect 7025 13789 8347 13790
rect 6766 13662 6862 13678
rect 8485 13678 8501 15222
rect 8565 13678 8581 15222
rect 10204 15222 10300 15238
rect 8744 15110 10066 15111
rect 8744 13790 8745 15110
rect 10065 13790 10066 15110
rect 8744 13789 10066 13790
rect 8485 13662 8581 13678
rect 10204 13678 10220 15222
rect 10284 13678 10300 15222
rect 11923 15222 12019 15238
rect 10463 15110 11785 15111
rect 10463 13790 10464 15110
rect 11784 13790 11785 15110
rect 10463 13789 11785 13790
rect 10204 13662 10300 13678
rect 11923 13678 11939 15222
rect 12003 13678 12019 15222
rect 13642 15222 13738 15238
rect 12182 15110 13504 15111
rect 12182 13790 12183 15110
rect 13503 13790 13504 15110
rect 12182 13789 13504 13790
rect 11923 13662 12019 13678
rect 13642 13678 13658 15222
rect 13722 13678 13738 15222
rect 15361 15222 15457 15238
rect 13901 15110 15223 15111
rect 13901 13790 13902 15110
rect 15222 13790 15223 15110
rect 13901 13789 15223 13790
rect 13642 13662 13738 13678
rect 15361 13678 15377 15222
rect 15441 13678 15457 15222
rect 15361 13662 15457 13678
rect -13862 13522 -13766 13538
rect -15322 13410 -14000 13411
rect -15322 12090 -15321 13410
rect -14001 12090 -14000 13410
rect -15322 12089 -14000 12090
rect -13862 11978 -13846 13522
rect -13782 11978 -13766 13522
rect -12143 13522 -12047 13538
rect -13603 13410 -12281 13411
rect -13603 12090 -13602 13410
rect -12282 12090 -12281 13410
rect -13603 12089 -12281 12090
rect -13862 11962 -13766 11978
rect -12143 11978 -12127 13522
rect -12063 11978 -12047 13522
rect -10424 13522 -10328 13538
rect -11884 13410 -10562 13411
rect -11884 12090 -11883 13410
rect -10563 12090 -10562 13410
rect -11884 12089 -10562 12090
rect -12143 11962 -12047 11978
rect -10424 11978 -10408 13522
rect -10344 11978 -10328 13522
rect -8705 13522 -8609 13538
rect -10165 13410 -8843 13411
rect -10165 12090 -10164 13410
rect -8844 12090 -8843 13410
rect -10165 12089 -8843 12090
rect -10424 11962 -10328 11978
rect -8705 11978 -8689 13522
rect -8625 11978 -8609 13522
rect -6986 13522 -6890 13538
rect -8446 13410 -7124 13411
rect -8446 12090 -8445 13410
rect -7125 12090 -7124 13410
rect -8446 12089 -7124 12090
rect -8705 11962 -8609 11978
rect -6986 11978 -6970 13522
rect -6906 11978 -6890 13522
rect -5267 13522 -5171 13538
rect -6727 13410 -5405 13411
rect -6727 12090 -6726 13410
rect -5406 12090 -5405 13410
rect -6727 12089 -5405 12090
rect -6986 11962 -6890 11978
rect -5267 11978 -5251 13522
rect -5187 11978 -5171 13522
rect -3548 13522 -3452 13538
rect -5008 13410 -3686 13411
rect -5008 12090 -5007 13410
rect -3687 12090 -3686 13410
rect -5008 12089 -3686 12090
rect -5267 11962 -5171 11978
rect -3548 11978 -3532 13522
rect -3468 11978 -3452 13522
rect -1829 13522 -1733 13538
rect -3289 13410 -1967 13411
rect -3289 12090 -3288 13410
rect -1968 12090 -1967 13410
rect -3289 12089 -1967 12090
rect -3548 11962 -3452 11978
rect -1829 11978 -1813 13522
rect -1749 11978 -1733 13522
rect -110 13522 -14 13538
rect -1570 13410 -248 13411
rect -1570 12090 -1569 13410
rect -249 12090 -248 13410
rect -1570 12089 -248 12090
rect -1829 11962 -1733 11978
rect -110 11978 -94 13522
rect -30 11978 -14 13522
rect 1609 13522 1705 13538
rect 149 13410 1471 13411
rect 149 12090 150 13410
rect 1470 12090 1471 13410
rect 149 12089 1471 12090
rect -110 11962 -14 11978
rect 1609 11978 1625 13522
rect 1689 11978 1705 13522
rect 3328 13522 3424 13538
rect 1868 13410 3190 13411
rect 1868 12090 1869 13410
rect 3189 12090 3190 13410
rect 1868 12089 3190 12090
rect 1609 11962 1705 11978
rect 3328 11978 3344 13522
rect 3408 11978 3424 13522
rect 5047 13522 5143 13538
rect 3587 13410 4909 13411
rect 3587 12090 3588 13410
rect 4908 12090 4909 13410
rect 3587 12089 4909 12090
rect 3328 11962 3424 11978
rect 5047 11978 5063 13522
rect 5127 11978 5143 13522
rect 6766 13522 6862 13538
rect 5306 13410 6628 13411
rect 5306 12090 5307 13410
rect 6627 12090 6628 13410
rect 5306 12089 6628 12090
rect 5047 11962 5143 11978
rect 6766 11978 6782 13522
rect 6846 11978 6862 13522
rect 8485 13522 8581 13538
rect 7025 13410 8347 13411
rect 7025 12090 7026 13410
rect 8346 12090 8347 13410
rect 7025 12089 8347 12090
rect 6766 11962 6862 11978
rect 8485 11978 8501 13522
rect 8565 11978 8581 13522
rect 10204 13522 10300 13538
rect 8744 13410 10066 13411
rect 8744 12090 8745 13410
rect 10065 12090 10066 13410
rect 8744 12089 10066 12090
rect 8485 11962 8581 11978
rect 10204 11978 10220 13522
rect 10284 11978 10300 13522
rect 11923 13522 12019 13538
rect 10463 13410 11785 13411
rect 10463 12090 10464 13410
rect 11784 12090 11785 13410
rect 10463 12089 11785 12090
rect 10204 11962 10300 11978
rect 11923 11978 11939 13522
rect 12003 11978 12019 13522
rect 13642 13522 13738 13538
rect 12182 13410 13504 13411
rect 12182 12090 12183 13410
rect 13503 12090 13504 13410
rect 12182 12089 13504 12090
rect 11923 11962 12019 11978
rect 13642 11978 13658 13522
rect 13722 11978 13738 13522
rect 15361 13522 15457 13538
rect 13901 13410 15223 13411
rect 13901 12090 13902 13410
rect 15222 12090 15223 13410
rect 13901 12089 15223 12090
rect 13642 11962 13738 11978
rect 15361 11978 15377 13522
rect 15441 11978 15457 13522
rect 15361 11962 15457 11978
rect -13862 11822 -13766 11838
rect -15322 11710 -14000 11711
rect -15322 10390 -15321 11710
rect -14001 10390 -14000 11710
rect -15322 10389 -14000 10390
rect -13862 10278 -13846 11822
rect -13782 10278 -13766 11822
rect -12143 11822 -12047 11838
rect -13603 11710 -12281 11711
rect -13603 10390 -13602 11710
rect -12282 10390 -12281 11710
rect -13603 10389 -12281 10390
rect -13862 10262 -13766 10278
rect -12143 10278 -12127 11822
rect -12063 10278 -12047 11822
rect -10424 11822 -10328 11838
rect -11884 11710 -10562 11711
rect -11884 10390 -11883 11710
rect -10563 10390 -10562 11710
rect -11884 10389 -10562 10390
rect -12143 10262 -12047 10278
rect -10424 10278 -10408 11822
rect -10344 10278 -10328 11822
rect -8705 11822 -8609 11838
rect -10165 11710 -8843 11711
rect -10165 10390 -10164 11710
rect -8844 10390 -8843 11710
rect -10165 10389 -8843 10390
rect -10424 10262 -10328 10278
rect -8705 10278 -8689 11822
rect -8625 10278 -8609 11822
rect -6986 11822 -6890 11838
rect -8446 11710 -7124 11711
rect -8446 10390 -8445 11710
rect -7125 10390 -7124 11710
rect -8446 10389 -7124 10390
rect -8705 10262 -8609 10278
rect -6986 10278 -6970 11822
rect -6906 10278 -6890 11822
rect -5267 11822 -5171 11838
rect -6727 11710 -5405 11711
rect -6727 10390 -6726 11710
rect -5406 10390 -5405 11710
rect -6727 10389 -5405 10390
rect -6986 10262 -6890 10278
rect -5267 10278 -5251 11822
rect -5187 10278 -5171 11822
rect -3548 11822 -3452 11838
rect -5008 11710 -3686 11711
rect -5008 10390 -5007 11710
rect -3687 10390 -3686 11710
rect -5008 10389 -3686 10390
rect -5267 10262 -5171 10278
rect -3548 10278 -3532 11822
rect -3468 10278 -3452 11822
rect -1829 11822 -1733 11838
rect -3289 11710 -1967 11711
rect -3289 10390 -3288 11710
rect -1968 10390 -1967 11710
rect -3289 10389 -1967 10390
rect -3548 10262 -3452 10278
rect -1829 10278 -1813 11822
rect -1749 10278 -1733 11822
rect -110 11822 -14 11838
rect -1570 11710 -248 11711
rect -1570 10390 -1569 11710
rect -249 10390 -248 11710
rect -1570 10389 -248 10390
rect -1829 10262 -1733 10278
rect -110 10278 -94 11822
rect -30 10278 -14 11822
rect 1609 11822 1705 11838
rect 149 11710 1471 11711
rect 149 10390 150 11710
rect 1470 10390 1471 11710
rect 149 10389 1471 10390
rect -110 10262 -14 10278
rect 1609 10278 1625 11822
rect 1689 10278 1705 11822
rect 3328 11822 3424 11838
rect 1868 11710 3190 11711
rect 1868 10390 1869 11710
rect 3189 10390 3190 11710
rect 1868 10389 3190 10390
rect 1609 10262 1705 10278
rect 3328 10278 3344 11822
rect 3408 10278 3424 11822
rect 5047 11822 5143 11838
rect 3587 11710 4909 11711
rect 3587 10390 3588 11710
rect 4908 10390 4909 11710
rect 3587 10389 4909 10390
rect 3328 10262 3424 10278
rect 5047 10278 5063 11822
rect 5127 10278 5143 11822
rect 6766 11822 6862 11838
rect 5306 11710 6628 11711
rect 5306 10390 5307 11710
rect 6627 10390 6628 11710
rect 5306 10389 6628 10390
rect 5047 10262 5143 10278
rect 6766 10278 6782 11822
rect 6846 10278 6862 11822
rect 8485 11822 8581 11838
rect 7025 11710 8347 11711
rect 7025 10390 7026 11710
rect 8346 10390 8347 11710
rect 7025 10389 8347 10390
rect 6766 10262 6862 10278
rect 8485 10278 8501 11822
rect 8565 10278 8581 11822
rect 10204 11822 10300 11838
rect 8744 11710 10066 11711
rect 8744 10390 8745 11710
rect 10065 10390 10066 11710
rect 8744 10389 10066 10390
rect 8485 10262 8581 10278
rect 10204 10278 10220 11822
rect 10284 10278 10300 11822
rect 11923 11822 12019 11838
rect 10463 11710 11785 11711
rect 10463 10390 10464 11710
rect 11784 10390 11785 11710
rect 10463 10389 11785 10390
rect 10204 10262 10300 10278
rect 11923 10278 11939 11822
rect 12003 10278 12019 11822
rect 13642 11822 13738 11838
rect 12182 11710 13504 11711
rect 12182 10390 12183 11710
rect 13503 10390 13504 11710
rect 12182 10389 13504 10390
rect 11923 10262 12019 10278
rect 13642 10278 13658 11822
rect 13722 10278 13738 11822
rect 15361 11822 15457 11838
rect 13901 11710 15223 11711
rect 13901 10390 13902 11710
rect 15222 10390 15223 11710
rect 13901 10389 15223 10390
rect 13642 10262 13738 10278
rect 15361 10278 15377 11822
rect 15441 10278 15457 11822
rect 15361 10262 15457 10278
rect -13862 10122 -13766 10138
rect -15322 10010 -14000 10011
rect -15322 8690 -15321 10010
rect -14001 8690 -14000 10010
rect -15322 8689 -14000 8690
rect -13862 8578 -13846 10122
rect -13782 8578 -13766 10122
rect -12143 10122 -12047 10138
rect -13603 10010 -12281 10011
rect -13603 8690 -13602 10010
rect -12282 8690 -12281 10010
rect -13603 8689 -12281 8690
rect -13862 8562 -13766 8578
rect -12143 8578 -12127 10122
rect -12063 8578 -12047 10122
rect -10424 10122 -10328 10138
rect -11884 10010 -10562 10011
rect -11884 8690 -11883 10010
rect -10563 8690 -10562 10010
rect -11884 8689 -10562 8690
rect -12143 8562 -12047 8578
rect -10424 8578 -10408 10122
rect -10344 8578 -10328 10122
rect -8705 10122 -8609 10138
rect -10165 10010 -8843 10011
rect -10165 8690 -10164 10010
rect -8844 8690 -8843 10010
rect -10165 8689 -8843 8690
rect -10424 8562 -10328 8578
rect -8705 8578 -8689 10122
rect -8625 8578 -8609 10122
rect -6986 10122 -6890 10138
rect -8446 10010 -7124 10011
rect -8446 8690 -8445 10010
rect -7125 8690 -7124 10010
rect -8446 8689 -7124 8690
rect -8705 8562 -8609 8578
rect -6986 8578 -6970 10122
rect -6906 8578 -6890 10122
rect -5267 10122 -5171 10138
rect -6727 10010 -5405 10011
rect -6727 8690 -6726 10010
rect -5406 8690 -5405 10010
rect -6727 8689 -5405 8690
rect -6986 8562 -6890 8578
rect -5267 8578 -5251 10122
rect -5187 8578 -5171 10122
rect -3548 10122 -3452 10138
rect -5008 10010 -3686 10011
rect -5008 8690 -5007 10010
rect -3687 8690 -3686 10010
rect -5008 8689 -3686 8690
rect -5267 8562 -5171 8578
rect -3548 8578 -3532 10122
rect -3468 8578 -3452 10122
rect -1829 10122 -1733 10138
rect -3289 10010 -1967 10011
rect -3289 8690 -3288 10010
rect -1968 8690 -1967 10010
rect -3289 8689 -1967 8690
rect -3548 8562 -3452 8578
rect -1829 8578 -1813 10122
rect -1749 8578 -1733 10122
rect -110 10122 -14 10138
rect -1570 10010 -248 10011
rect -1570 8690 -1569 10010
rect -249 8690 -248 10010
rect -1570 8689 -248 8690
rect -1829 8562 -1733 8578
rect -110 8578 -94 10122
rect -30 8578 -14 10122
rect 1609 10122 1705 10138
rect 149 10010 1471 10011
rect 149 8690 150 10010
rect 1470 8690 1471 10010
rect 149 8689 1471 8690
rect -110 8562 -14 8578
rect 1609 8578 1625 10122
rect 1689 8578 1705 10122
rect 3328 10122 3424 10138
rect 1868 10010 3190 10011
rect 1868 8690 1869 10010
rect 3189 8690 3190 10010
rect 1868 8689 3190 8690
rect 1609 8562 1705 8578
rect 3328 8578 3344 10122
rect 3408 8578 3424 10122
rect 5047 10122 5143 10138
rect 3587 10010 4909 10011
rect 3587 8690 3588 10010
rect 4908 8690 4909 10010
rect 3587 8689 4909 8690
rect 3328 8562 3424 8578
rect 5047 8578 5063 10122
rect 5127 8578 5143 10122
rect 6766 10122 6862 10138
rect 5306 10010 6628 10011
rect 5306 8690 5307 10010
rect 6627 8690 6628 10010
rect 5306 8689 6628 8690
rect 5047 8562 5143 8578
rect 6766 8578 6782 10122
rect 6846 8578 6862 10122
rect 8485 10122 8581 10138
rect 7025 10010 8347 10011
rect 7025 8690 7026 10010
rect 8346 8690 8347 10010
rect 7025 8689 8347 8690
rect 6766 8562 6862 8578
rect 8485 8578 8501 10122
rect 8565 8578 8581 10122
rect 10204 10122 10300 10138
rect 8744 10010 10066 10011
rect 8744 8690 8745 10010
rect 10065 8690 10066 10010
rect 8744 8689 10066 8690
rect 8485 8562 8581 8578
rect 10204 8578 10220 10122
rect 10284 8578 10300 10122
rect 11923 10122 12019 10138
rect 10463 10010 11785 10011
rect 10463 8690 10464 10010
rect 11784 8690 11785 10010
rect 10463 8689 11785 8690
rect 10204 8562 10300 8578
rect 11923 8578 11939 10122
rect 12003 8578 12019 10122
rect 13642 10122 13738 10138
rect 12182 10010 13504 10011
rect 12182 8690 12183 10010
rect 13503 8690 13504 10010
rect 12182 8689 13504 8690
rect 11923 8562 12019 8578
rect 13642 8578 13658 10122
rect 13722 8578 13738 10122
rect 15361 10122 15457 10138
rect 13901 10010 15223 10011
rect 13901 8690 13902 10010
rect 15222 8690 15223 10010
rect 13901 8689 15223 8690
rect 13642 8562 13738 8578
rect 15361 8578 15377 10122
rect 15441 8578 15457 10122
rect 15361 8562 15457 8578
rect -13862 8422 -13766 8438
rect -15322 8310 -14000 8311
rect -15322 6990 -15321 8310
rect -14001 6990 -14000 8310
rect -15322 6989 -14000 6990
rect -13862 6878 -13846 8422
rect -13782 6878 -13766 8422
rect -12143 8422 -12047 8438
rect -13603 8310 -12281 8311
rect -13603 6990 -13602 8310
rect -12282 6990 -12281 8310
rect -13603 6989 -12281 6990
rect -13862 6862 -13766 6878
rect -12143 6878 -12127 8422
rect -12063 6878 -12047 8422
rect -10424 8422 -10328 8438
rect -11884 8310 -10562 8311
rect -11884 6990 -11883 8310
rect -10563 6990 -10562 8310
rect -11884 6989 -10562 6990
rect -12143 6862 -12047 6878
rect -10424 6878 -10408 8422
rect -10344 6878 -10328 8422
rect -8705 8422 -8609 8438
rect -10165 8310 -8843 8311
rect -10165 6990 -10164 8310
rect -8844 6990 -8843 8310
rect -10165 6989 -8843 6990
rect -10424 6862 -10328 6878
rect -8705 6878 -8689 8422
rect -8625 6878 -8609 8422
rect -6986 8422 -6890 8438
rect -8446 8310 -7124 8311
rect -8446 6990 -8445 8310
rect -7125 6990 -7124 8310
rect -8446 6989 -7124 6990
rect -8705 6862 -8609 6878
rect -6986 6878 -6970 8422
rect -6906 6878 -6890 8422
rect -5267 8422 -5171 8438
rect -6727 8310 -5405 8311
rect -6727 6990 -6726 8310
rect -5406 6990 -5405 8310
rect -6727 6989 -5405 6990
rect -6986 6862 -6890 6878
rect -5267 6878 -5251 8422
rect -5187 6878 -5171 8422
rect -3548 8422 -3452 8438
rect -5008 8310 -3686 8311
rect -5008 6990 -5007 8310
rect -3687 6990 -3686 8310
rect -5008 6989 -3686 6990
rect -5267 6862 -5171 6878
rect -3548 6878 -3532 8422
rect -3468 6878 -3452 8422
rect -1829 8422 -1733 8438
rect -3289 8310 -1967 8311
rect -3289 6990 -3288 8310
rect -1968 6990 -1967 8310
rect -3289 6989 -1967 6990
rect -3548 6862 -3452 6878
rect -1829 6878 -1813 8422
rect -1749 6878 -1733 8422
rect -110 8422 -14 8438
rect -1570 8310 -248 8311
rect -1570 6990 -1569 8310
rect -249 6990 -248 8310
rect -1570 6989 -248 6990
rect -1829 6862 -1733 6878
rect -110 6878 -94 8422
rect -30 6878 -14 8422
rect 1609 8422 1705 8438
rect 149 8310 1471 8311
rect 149 6990 150 8310
rect 1470 6990 1471 8310
rect 149 6989 1471 6990
rect -110 6862 -14 6878
rect 1609 6878 1625 8422
rect 1689 6878 1705 8422
rect 3328 8422 3424 8438
rect 1868 8310 3190 8311
rect 1868 6990 1869 8310
rect 3189 6990 3190 8310
rect 1868 6989 3190 6990
rect 1609 6862 1705 6878
rect 3328 6878 3344 8422
rect 3408 6878 3424 8422
rect 5047 8422 5143 8438
rect 3587 8310 4909 8311
rect 3587 6990 3588 8310
rect 4908 6990 4909 8310
rect 3587 6989 4909 6990
rect 3328 6862 3424 6878
rect 5047 6878 5063 8422
rect 5127 6878 5143 8422
rect 6766 8422 6862 8438
rect 5306 8310 6628 8311
rect 5306 6990 5307 8310
rect 6627 6990 6628 8310
rect 5306 6989 6628 6990
rect 5047 6862 5143 6878
rect 6766 6878 6782 8422
rect 6846 6878 6862 8422
rect 8485 8422 8581 8438
rect 7025 8310 8347 8311
rect 7025 6990 7026 8310
rect 8346 6990 8347 8310
rect 7025 6989 8347 6990
rect 6766 6862 6862 6878
rect 8485 6878 8501 8422
rect 8565 6878 8581 8422
rect 10204 8422 10300 8438
rect 8744 8310 10066 8311
rect 8744 6990 8745 8310
rect 10065 6990 10066 8310
rect 8744 6989 10066 6990
rect 8485 6862 8581 6878
rect 10204 6878 10220 8422
rect 10284 6878 10300 8422
rect 11923 8422 12019 8438
rect 10463 8310 11785 8311
rect 10463 6990 10464 8310
rect 11784 6990 11785 8310
rect 10463 6989 11785 6990
rect 10204 6862 10300 6878
rect 11923 6878 11939 8422
rect 12003 6878 12019 8422
rect 13642 8422 13738 8438
rect 12182 8310 13504 8311
rect 12182 6990 12183 8310
rect 13503 6990 13504 8310
rect 12182 6989 13504 6990
rect 11923 6862 12019 6878
rect 13642 6878 13658 8422
rect 13722 6878 13738 8422
rect 15361 8422 15457 8438
rect 13901 8310 15223 8311
rect 13901 6990 13902 8310
rect 15222 6990 15223 8310
rect 13901 6989 15223 6990
rect 13642 6862 13738 6878
rect 15361 6878 15377 8422
rect 15441 6878 15457 8422
rect 15361 6862 15457 6878
rect -13862 6722 -13766 6738
rect -15322 6610 -14000 6611
rect -15322 5290 -15321 6610
rect -14001 5290 -14000 6610
rect -15322 5289 -14000 5290
rect -13862 5178 -13846 6722
rect -13782 5178 -13766 6722
rect -12143 6722 -12047 6738
rect -13603 6610 -12281 6611
rect -13603 5290 -13602 6610
rect -12282 5290 -12281 6610
rect -13603 5289 -12281 5290
rect -13862 5162 -13766 5178
rect -12143 5178 -12127 6722
rect -12063 5178 -12047 6722
rect -10424 6722 -10328 6738
rect -11884 6610 -10562 6611
rect -11884 5290 -11883 6610
rect -10563 5290 -10562 6610
rect -11884 5289 -10562 5290
rect -12143 5162 -12047 5178
rect -10424 5178 -10408 6722
rect -10344 5178 -10328 6722
rect -8705 6722 -8609 6738
rect -10165 6610 -8843 6611
rect -10165 5290 -10164 6610
rect -8844 5290 -8843 6610
rect -10165 5289 -8843 5290
rect -10424 5162 -10328 5178
rect -8705 5178 -8689 6722
rect -8625 5178 -8609 6722
rect -6986 6722 -6890 6738
rect -8446 6610 -7124 6611
rect -8446 5290 -8445 6610
rect -7125 5290 -7124 6610
rect -8446 5289 -7124 5290
rect -8705 5162 -8609 5178
rect -6986 5178 -6970 6722
rect -6906 5178 -6890 6722
rect -5267 6722 -5171 6738
rect -6727 6610 -5405 6611
rect -6727 5290 -6726 6610
rect -5406 5290 -5405 6610
rect -6727 5289 -5405 5290
rect -6986 5162 -6890 5178
rect -5267 5178 -5251 6722
rect -5187 5178 -5171 6722
rect -3548 6722 -3452 6738
rect -5008 6610 -3686 6611
rect -5008 5290 -5007 6610
rect -3687 5290 -3686 6610
rect -5008 5289 -3686 5290
rect -5267 5162 -5171 5178
rect -3548 5178 -3532 6722
rect -3468 5178 -3452 6722
rect -1829 6722 -1733 6738
rect -3289 6610 -1967 6611
rect -3289 5290 -3288 6610
rect -1968 5290 -1967 6610
rect -3289 5289 -1967 5290
rect -3548 5162 -3452 5178
rect -1829 5178 -1813 6722
rect -1749 5178 -1733 6722
rect -110 6722 -14 6738
rect -1570 6610 -248 6611
rect -1570 5290 -1569 6610
rect -249 5290 -248 6610
rect -1570 5289 -248 5290
rect -1829 5162 -1733 5178
rect -110 5178 -94 6722
rect -30 5178 -14 6722
rect 1609 6722 1705 6738
rect 149 6610 1471 6611
rect 149 5290 150 6610
rect 1470 5290 1471 6610
rect 149 5289 1471 5290
rect -110 5162 -14 5178
rect 1609 5178 1625 6722
rect 1689 5178 1705 6722
rect 3328 6722 3424 6738
rect 1868 6610 3190 6611
rect 1868 5290 1869 6610
rect 3189 5290 3190 6610
rect 1868 5289 3190 5290
rect 1609 5162 1705 5178
rect 3328 5178 3344 6722
rect 3408 5178 3424 6722
rect 5047 6722 5143 6738
rect 3587 6610 4909 6611
rect 3587 5290 3588 6610
rect 4908 5290 4909 6610
rect 3587 5289 4909 5290
rect 3328 5162 3424 5178
rect 5047 5178 5063 6722
rect 5127 5178 5143 6722
rect 6766 6722 6862 6738
rect 5306 6610 6628 6611
rect 5306 5290 5307 6610
rect 6627 5290 6628 6610
rect 5306 5289 6628 5290
rect 5047 5162 5143 5178
rect 6766 5178 6782 6722
rect 6846 5178 6862 6722
rect 8485 6722 8581 6738
rect 7025 6610 8347 6611
rect 7025 5290 7026 6610
rect 8346 5290 8347 6610
rect 7025 5289 8347 5290
rect 6766 5162 6862 5178
rect 8485 5178 8501 6722
rect 8565 5178 8581 6722
rect 10204 6722 10300 6738
rect 8744 6610 10066 6611
rect 8744 5290 8745 6610
rect 10065 5290 10066 6610
rect 8744 5289 10066 5290
rect 8485 5162 8581 5178
rect 10204 5178 10220 6722
rect 10284 5178 10300 6722
rect 11923 6722 12019 6738
rect 10463 6610 11785 6611
rect 10463 5290 10464 6610
rect 11784 5290 11785 6610
rect 10463 5289 11785 5290
rect 10204 5162 10300 5178
rect 11923 5178 11939 6722
rect 12003 5178 12019 6722
rect 13642 6722 13738 6738
rect 12182 6610 13504 6611
rect 12182 5290 12183 6610
rect 13503 5290 13504 6610
rect 12182 5289 13504 5290
rect 11923 5162 12019 5178
rect 13642 5178 13658 6722
rect 13722 5178 13738 6722
rect 15361 6722 15457 6738
rect 13901 6610 15223 6611
rect 13901 5290 13902 6610
rect 15222 5290 15223 6610
rect 13901 5289 15223 5290
rect 13642 5162 13738 5178
rect 15361 5178 15377 6722
rect 15441 5178 15457 6722
rect 15361 5162 15457 5178
rect -13862 5022 -13766 5038
rect -15322 4910 -14000 4911
rect -15322 3590 -15321 4910
rect -14001 3590 -14000 4910
rect -15322 3589 -14000 3590
rect -13862 3478 -13846 5022
rect -13782 3478 -13766 5022
rect -12143 5022 -12047 5038
rect -13603 4910 -12281 4911
rect -13603 3590 -13602 4910
rect -12282 3590 -12281 4910
rect -13603 3589 -12281 3590
rect -13862 3462 -13766 3478
rect -12143 3478 -12127 5022
rect -12063 3478 -12047 5022
rect -10424 5022 -10328 5038
rect -11884 4910 -10562 4911
rect -11884 3590 -11883 4910
rect -10563 3590 -10562 4910
rect -11884 3589 -10562 3590
rect -12143 3462 -12047 3478
rect -10424 3478 -10408 5022
rect -10344 3478 -10328 5022
rect -8705 5022 -8609 5038
rect -10165 4910 -8843 4911
rect -10165 3590 -10164 4910
rect -8844 3590 -8843 4910
rect -10165 3589 -8843 3590
rect -10424 3462 -10328 3478
rect -8705 3478 -8689 5022
rect -8625 3478 -8609 5022
rect -6986 5022 -6890 5038
rect -8446 4910 -7124 4911
rect -8446 3590 -8445 4910
rect -7125 3590 -7124 4910
rect -8446 3589 -7124 3590
rect -8705 3462 -8609 3478
rect -6986 3478 -6970 5022
rect -6906 3478 -6890 5022
rect -5267 5022 -5171 5038
rect -6727 4910 -5405 4911
rect -6727 3590 -6726 4910
rect -5406 3590 -5405 4910
rect -6727 3589 -5405 3590
rect -6986 3462 -6890 3478
rect -5267 3478 -5251 5022
rect -5187 3478 -5171 5022
rect -3548 5022 -3452 5038
rect -5008 4910 -3686 4911
rect -5008 3590 -5007 4910
rect -3687 3590 -3686 4910
rect -5008 3589 -3686 3590
rect -5267 3462 -5171 3478
rect -3548 3478 -3532 5022
rect -3468 3478 -3452 5022
rect -1829 5022 -1733 5038
rect -3289 4910 -1967 4911
rect -3289 3590 -3288 4910
rect -1968 3590 -1967 4910
rect -3289 3589 -1967 3590
rect -3548 3462 -3452 3478
rect -1829 3478 -1813 5022
rect -1749 3478 -1733 5022
rect -110 5022 -14 5038
rect -1570 4910 -248 4911
rect -1570 3590 -1569 4910
rect -249 3590 -248 4910
rect -1570 3589 -248 3590
rect -1829 3462 -1733 3478
rect -110 3478 -94 5022
rect -30 3478 -14 5022
rect 1609 5022 1705 5038
rect 149 4910 1471 4911
rect 149 3590 150 4910
rect 1470 3590 1471 4910
rect 149 3589 1471 3590
rect -110 3462 -14 3478
rect 1609 3478 1625 5022
rect 1689 3478 1705 5022
rect 3328 5022 3424 5038
rect 1868 4910 3190 4911
rect 1868 3590 1869 4910
rect 3189 3590 3190 4910
rect 1868 3589 3190 3590
rect 1609 3462 1705 3478
rect 3328 3478 3344 5022
rect 3408 3478 3424 5022
rect 5047 5022 5143 5038
rect 3587 4910 4909 4911
rect 3587 3590 3588 4910
rect 4908 3590 4909 4910
rect 3587 3589 4909 3590
rect 3328 3462 3424 3478
rect 5047 3478 5063 5022
rect 5127 3478 5143 5022
rect 6766 5022 6862 5038
rect 5306 4910 6628 4911
rect 5306 3590 5307 4910
rect 6627 3590 6628 4910
rect 5306 3589 6628 3590
rect 5047 3462 5143 3478
rect 6766 3478 6782 5022
rect 6846 3478 6862 5022
rect 8485 5022 8581 5038
rect 7025 4910 8347 4911
rect 7025 3590 7026 4910
rect 8346 3590 8347 4910
rect 7025 3589 8347 3590
rect 6766 3462 6862 3478
rect 8485 3478 8501 5022
rect 8565 3478 8581 5022
rect 10204 5022 10300 5038
rect 8744 4910 10066 4911
rect 8744 3590 8745 4910
rect 10065 3590 10066 4910
rect 8744 3589 10066 3590
rect 8485 3462 8581 3478
rect 10204 3478 10220 5022
rect 10284 3478 10300 5022
rect 11923 5022 12019 5038
rect 10463 4910 11785 4911
rect 10463 3590 10464 4910
rect 11784 3590 11785 4910
rect 10463 3589 11785 3590
rect 10204 3462 10300 3478
rect 11923 3478 11939 5022
rect 12003 3478 12019 5022
rect 13642 5022 13738 5038
rect 12182 4910 13504 4911
rect 12182 3590 12183 4910
rect 13503 3590 13504 4910
rect 12182 3589 13504 3590
rect 11923 3462 12019 3478
rect 13642 3478 13658 5022
rect 13722 3478 13738 5022
rect 15361 5022 15457 5038
rect 13901 4910 15223 4911
rect 13901 3590 13902 4910
rect 15222 3590 15223 4910
rect 13901 3589 15223 3590
rect 13642 3462 13738 3478
rect 15361 3478 15377 5022
rect 15441 3478 15457 5022
rect 15361 3462 15457 3478
rect -13862 3322 -13766 3338
rect -15322 3210 -14000 3211
rect -15322 1890 -15321 3210
rect -14001 1890 -14000 3210
rect -15322 1889 -14000 1890
rect -13862 1778 -13846 3322
rect -13782 1778 -13766 3322
rect -12143 3322 -12047 3338
rect -13603 3210 -12281 3211
rect -13603 1890 -13602 3210
rect -12282 1890 -12281 3210
rect -13603 1889 -12281 1890
rect -13862 1762 -13766 1778
rect -12143 1778 -12127 3322
rect -12063 1778 -12047 3322
rect -10424 3322 -10328 3338
rect -11884 3210 -10562 3211
rect -11884 1890 -11883 3210
rect -10563 1890 -10562 3210
rect -11884 1889 -10562 1890
rect -12143 1762 -12047 1778
rect -10424 1778 -10408 3322
rect -10344 1778 -10328 3322
rect -8705 3322 -8609 3338
rect -10165 3210 -8843 3211
rect -10165 1890 -10164 3210
rect -8844 1890 -8843 3210
rect -10165 1889 -8843 1890
rect -10424 1762 -10328 1778
rect -8705 1778 -8689 3322
rect -8625 1778 -8609 3322
rect -6986 3322 -6890 3338
rect -8446 3210 -7124 3211
rect -8446 1890 -8445 3210
rect -7125 1890 -7124 3210
rect -8446 1889 -7124 1890
rect -8705 1762 -8609 1778
rect -6986 1778 -6970 3322
rect -6906 1778 -6890 3322
rect -5267 3322 -5171 3338
rect -6727 3210 -5405 3211
rect -6727 1890 -6726 3210
rect -5406 1890 -5405 3210
rect -6727 1889 -5405 1890
rect -6986 1762 -6890 1778
rect -5267 1778 -5251 3322
rect -5187 1778 -5171 3322
rect -3548 3322 -3452 3338
rect -5008 3210 -3686 3211
rect -5008 1890 -5007 3210
rect -3687 1890 -3686 3210
rect -5008 1889 -3686 1890
rect -5267 1762 -5171 1778
rect -3548 1778 -3532 3322
rect -3468 1778 -3452 3322
rect -1829 3322 -1733 3338
rect -3289 3210 -1967 3211
rect -3289 1890 -3288 3210
rect -1968 1890 -1967 3210
rect -3289 1889 -1967 1890
rect -3548 1762 -3452 1778
rect -1829 1778 -1813 3322
rect -1749 1778 -1733 3322
rect -110 3322 -14 3338
rect -1570 3210 -248 3211
rect -1570 1890 -1569 3210
rect -249 1890 -248 3210
rect -1570 1889 -248 1890
rect -1829 1762 -1733 1778
rect -110 1778 -94 3322
rect -30 1778 -14 3322
rect 1609 3322 1705 3338
rect 149 3210 1471 3211
rect 149 1890 150 3210
rect 1470 1890 1471 3210
rect 149 1889 1471 1890
rect -110 1762 -14 1778
rect 1609 1778 1625 3322
rect 1689 1778 1705 3322
rect 3328 3322 3424 3338
rect 1868 3210 3190 3211
rect 1868 1890 1869 3210
rect 3189 1890 3190 3210
rect 1868 1889 3190 1890
rect 1609 1762 1705 1778
rect 3328 1778 3344 3322
rect 3408 1778 3424 3322
rect 5047 3322 5143 3338
rect 3587 3210 4909 3211
rect 3587 1890 3588 3210
rect 4908 1890 4909 3210
rect 3587 1889 4909 1890
rect 3328 1762 3424 1778
rect 5047 1778 5063 3322
rect 5127 1778 5143 3322
rect 6766 3322 6862 3338
rect 5306 3210 6628 3211
rect 5306 1890 5307 3210
rect 6627 1890 6628 3210
rect 5306 1889 6628 1890
rect 5047 1762 5143 1778
rect 6766 1778 6782 3322
rect 6846 1778 6862 3322
rect 8485 3322 8581 3338
rect 7025 3210 8347 3211
rect 7025 1890 7026 3210
rect 8346 1890 8347 3210
rect 7025 1889 8347 1890
rect 6766 1762 6862 1778
rect 8485 1778 8501 3322
rect 8565 1778 8581 3322
rect 10204 3322 10300 3338
rect 8744 3210 10066 3211
rect 8744 1890 8745 3210
rect 10065 1890 10066 3210
rect 8744 1889 10066 1890
rect 8485 1762 8581 1778
rect 10204 1778 10220 3322
rect 10284 1778 10300 3322
rect 11923 3322 12019 3338
rect 10463 3210 11785 3211
rect 10463 1890 10464 3210
rect 11784 1890 11785 3210
rect 10463 1889 11785 1890
rect 10204 1762 10300 1778
rect 11923 1778 11939 3322
rect 12003 1778 12019 3322
rect 13642 3322 13738 3338
rect 12182 3210 13504 3211
rect 12182 1890 12183 3210
rect 13503 1890 13504 3210
rect 12182 1889 13504 1890
rect 11923 1762 12019 1778
rect 13642 1778 13658 3322
rect 13722 1778 13738 3322
rect 15361 3322 15457 3338
rect 13901 3210 15223 3211
rect 13901 1890 13902 3210
rect 15222 1890 15223 3210
rect 13901 1889 15223 1890
rect 13642 1762 13738 1778
rect 15361 1778 15377 3322
rect 15441 1778 15457 3322
rect 15361 1762 15457 1778
rect -13862 1622 -13766 1638
rect -15322 1510 -14000 1511
rect -15322 190 -15321 1510
rect -14001 190 -14000 1510
rect -15322 189 -14000 190
rect -13862 78 -13846 1622
rect -13782 78 -13766 1622
rect -12143 1622 -12047 1638
rect -13603 1510 -12281 1511
rect -13603 190 -13602 1510
rect -12282 190 -12281 1510
rect -13603 189 -12281 190
rect -13862 62 -13766 78
rect -12143 78 -12127 1622
rect -12063 78 -12047 1622
rect -10424 1622 -10328 1638
rect -11884 1510 -10562 1511
rect -11884 190 -11883 1510
rect -10563 190 -10562 1510
rect -11884 189 -10562 190
rect -12143 62 -12047 78
rect -10424 78 -10408 1622
rect -10344 78 -10328 1622
rect -8705 1622 -8609 1638
rect -10165 1510 -8843 1511
rect -10165 190 -10164 1510
rect -8844 190 -8843 1510
rect -10165 189 -8843 190
rect -10424 62 -10328 78
rect -8705 78 -8689 1622
rect -8625 78 -8609 1622
rect -6986 1622 -6890 1638
rect -8446 1510 -7124 1511
rect -8446 190 -8445 1510
rect -7125 190 -7124 1510
rect -8446 189 -7124 190
rect -8705 62 -8609 78
rect -6986 78 -6970 1622
rect -6906 78 -6890 1622
rect -5267 1622 -5171 1638
rect -6727 1510 -5405 1511
rect -6727 190 -6726 1510
rect -5406 190 -5405 1510
rect -6727 189 -5405 190
rect -6986 62 -6890 78
rect -5267 78 -5251 1622
rect -5187 78 -5171 1622
rect -3548 1622 -3452 1638
rect -5008 1510 -3686 1511
rect -5008 190 -5007 1510
rect -3687 190 -3686 1510
rect -5008 189 -3686 190
rect -5267 62 -5171 78
rect -3548 78 -3532 1622
rect -3468 78 -3452 1622
rect -1829 1622 -1733 1638
rect -3289 1510 -1967 1511
rect -3289 190 -3288 1510
rect -1968 190 -1967 1510
rect -3289 189 -1967 190
rect -3548 62 -3452 78
rect -1829 78 -1813 1622
rect -1749 78 -1733 1622
rect -110 1622 -14 1638
rect -1570 1510 -248 1511
rect -1570 190 -1569 1510
rect -249 190 -248 1510
rect -1570 189 -248 190
rect -1829 62 -1733 78
rect -110 78 -94 1622
rect -30 78 -14 1622
rect 1609 1622 1705 1638
rect 149 1510 1471 1511
rect 149 190 150 1510
rect 1470 190 1471 1510
rect 149 189 1471 190
rect -110 62 -14 78
rect 1609 78 1625 1622
rect 1689 78 1705 1622
rect 3328 1622 3424 1638
rect 1868 1510 3190 1511
rect 1868 190 1869 1510
rect 3189 190 3190 1510
rect 1868 189 3190 190
rect 1609 62 1705 78
rect 3328 78 3344 1622
rect 3408 78 3424 1622
rect 5047 1622 5143 1638
rect 3587 1510 4909 1511
rect 3587 190 3588 1510
rect 4908 190 4909 1510
rect 3587 189 4909 190
rect 3328 62 3424 78
rect 5047 78 5063 1622
rect 5127 78 5143 1622
rect 6766 1622 6862 1638
rect 5306 1510 6628 1511
rect 5306 190 5307 1510
rect 6627 190 6628 1510
rect 5306 189 6628 190
rect 5047 62 5143 78
rect 6766 78 6782 1622
rect 6846 78 6862 1622
rect 8485 1622 8581 1638
rect 7025 1510 8347 1511
rect 7025 190 7026 1510
rect 8346 190 8347 1510
rect 7025 189 8347 190
rect 6766 62 6862 78
rect 8485 78 8501 1622
rect 8565 78 8581 1622
rect 10204 1622 10300 1638
rect 8744 1510 10066 1511
rect 8744 190 8745 1510
rect 10065 190 10066 1510
rect 8744 189 10066 190
rect 8485 62 8581 78
rect 10204 78 10220 1622
rect 10284 78 10300 1622
rect 11923 1622 12019 1638
rect 10463 1510 11785 1511
rect 10463 190 10464 1510
rect 11784 190 11785 1510
rect 10463 189 11785 190
rect 10204 62 10300 78
rect 11923 78 11939 1622
rect 12003 78 12019 1622
rect 13642 1622 13738 1638
rect 12182 1510 13504 1511
rect 12182 190 12183 1510
rect 13503 190 13504 1510
rect 12182 189 13504 190
rect 11923 62 12019 78
rect 13642 78 13658 1622
rect 13722 78 13738 1622
rect 15361 1622 15457 1638
rect 13901 1510 15223 1511
rect 13901 190 13902 1510
rect 15222 190 15223 1510
rect 13901 189 15223 190
rect 13642 62 13738 78
rect 15361 78 15377 1622
rect 15441 78 15457 1622
rect 15361 62 15457 78
rect -13862 -78 -13766 -62
rect -15322 -190 -14000 -189
rect -15322 -1510 -15321 -190
rect -14001 -1510 -14000 -190
rect -15322 -1511 -14000 -1510
rect -13862 -1622 -13846 -78
rect -13782 -1622 -13766 -78
rect -12143 -78 -12047 -62
rect -13603 -190 -12281 -189
rect -13603 -1510 -13602 -190
rect -12282 -1510 -12281 -190
rect -13603 -1511 -12281 -1510
rect -13862 -1638 -13766 -1622
rect -12143 -1622 -12127 -78
rect -12063 -1622 -12047 -78
rect -10424 -78 -10328 -62
rect -11884 -190 -10562 -189
rect -11884 -1510 -11883 -190
rect -10563 -1510 -10562 -190
rect -11884 -1511 -10562 -1510
rect -12143 -1638 -12047 -1622
rect -10424 -1622 -10408 -78
rect -10344 -1622 -10328 -78
rect -8705 -78 -8609 -62
rect -10165 -190 -8843 -189
rect -10165 -1510 -10164 -190
rect -8844 -1510 -8843 -190
rect -10165 -1511 -8843 -1510
rect -10424 -1638 -10328 -1622
rect -8705 -1622 -8689 -78
rect -8625 -1622 -8609 -78
rect -6986 -78 -6890 -62
rect -8446 -190 -7124 -189
rect -8446 -1510 -8445 -190
rect -7125 -1510 -7124 -190
rect -8446 -1511 -7124 -1510
rect -8705 -1638 -8609 -1622
rect -6986 -1622 -6970 -78
rect -6906 -1622 -6890 -78
rect -5267 -78 -5171 -62
rect -6727 -190 -5405 -189
rect -6727 -1510 -6726 -190
rect -5406 -1510 -5405 -190
rect -6727 -1511 -5405 -1510
rect -6986 -1638 -6890 -1622
rect -5267 -1622 -5251 -78
rect -5187 -1622 -5171 -78
rect -3548 -78 -3452 -62
rect -5008 -190 -3686 -189
rect -5008 -1510 -5007 -190
rect -3687 -1510 -3686 -190
rect -5008 -1511 -3686 -1510
rect -5267 -1638 -5171 -1622
rect -3548 -1622 -3532 -78
rect -3468 -1622 -3452 -78
rect -1829 -78 -1733 -62
rect -3289 -190 -1967 -189
rect -3289 -1510 -3288 -190
rect -1968 -1510 -1967 -190
rect -3289 -1511 -1967 -1510
rect -3548 -1638 -3452 -1622
rect -1829 -1622 -1813 -78
rect -1749 -1622 -1733 -78
rect -110 -78 -14 -62
rect -1570 -190 -248 -189
rect -1570 -1510 -1569 -190
rect -249 -1510 -248 -190
rect -1570 -1511 -248 -1510
rect -1829 -1638 -1733 -1622
rect -110 -1622 -94 -78
rect -30 -1622 -14 -78
rect 1609 -78 1705 -62
rect 149 -190 1471 -189
rect 149 -1510 150 -190
rect 1470 -1510 1471 -190
rect 149 -1511 1471 -1510
rect -110 -1638 -14 -1622
rect 1609 -1622 1625 -78
rect 1689 -1622 1705 -78
rect 3328 -78 3424 -62
rect 1868 -190 3190 -189
rect 1868 -1510 1869 -190
rect 3189 -1510 3190 -190
rect 1868 -1511 3190 -1510
rect 1609 -1638 1705 -1622
rect 3328 -1622 3344 -78
rect 3408 -1622 3424 -78
rect 5047 -78 5143 -62
rect 3587 -190 4909 -189
rect 3587 -1510 3588 -190
rect 4908 -1510 4909 -190
rect 3587 -1511 4909 -1510
rect 3328 -1638 3424 -1622
rect 5047 -1622 5063 -78
rect 5127 -1622 5143 -78
rect 6766 -78 6862 -62
rect 5306 -190 6628 -189
rect 5306 -1510 5307 -190
rect 6627 -1510 6628 -190
rect 5306 -1511 6628 -1510
rect 5047 -1638 5143 -1622
rect 6766 -1622 6782 -78
rect 6846 -1622 6862 -78
rect 8485 -78 8581 -62
rect 7025 -190 8347 -189
rect 7025 -1510 7026 -190
rect 8346 -1510 8347 -190
rect 7025 -1511 8347 -1510
rect 6766 -1638 6862 -1622
rect 8485 -1622 8501 -78
rect 8565 -1622 8581 -78
rect 10204 -78 10300 -62
rect 8744 -190 10066 -189
rect 8744 -1510 8745 -190
rect 10065 -1510 10066 -190
rect 8744 -1511 10066 -1510
rect 8485 -1638 8581 -1622
rect 10204 -1622 10220 -78
rect 10284 -1622 10300 -78
rect 11923 -78 12019 -62
rect 10463 -190 11785 -189
rect 10463 -1510 10464 -190
rect 11784 -1510 11785 -190
rect 10463 -1511 11785 -1510
rect 10204 -1638 10300 -1622
rect 11923 -1622 11939 -78
rect 12003 -1622 12019 -78
rect 13642 -78 13738 -62
rect 12182 -190 13504 -189
rect 12182 -1510 12183 -190
rect 13503 -1510 13504 -190
rect 12182 -1511 13504 -1510
rect 11923 -1638 12019 -1622
rect 13642 -1622 13658 -78
rect 13722 -1622 13738 -78
rect 15361 -78 15457 -62
rect 13901 -190 15223 -189
rect 13901 -1510 13902 -190
rect 15222 -1510 15223 -190
rect 13901 -1511 15223 -1510
rect 13642 -1638 13738 -1622
rect 15361 -1622 15377 -78
rect 15441 -1622 15457 -78
rect 15361 -1638 15457 -1622
rect -13862 -1778 -13766 -1762
rect -15322 -1890 -14000 -1889
rect -15322 -3210 -15321 -1890
rect -14001 -3210 -14000 -1890
rect -15322 -3211 -14000 -3210
rect -13862 -3322 -13846 -1778
rect -13782 -3322 -13766 -1778
rect -12143 -1778 -12047 -1762
rect -13603 -1890 -12281 -1889
rect -13603 -3210 -13602 -1890
rect -12282 -3210 -12281 -1890
rect -13603 -3211 -12281 -3210
rect -13862 -3338 -13766 -3322
rect -12143 -3322 -12127 -1778
rect -12063 -3322 -12047 -1778
rect -10424 -1778 -10328 -1762
rect -11884 -1890 -10562 -1889
rect -11884 -3210 -11883 -1890
rect -10563 -3210 -10562 -1890
rect -11884 -3211 -10562 -3210
rect -12143 -3338 -12047 -3322
rect -10424 -3322 -10408 -1778
rect -10344 -3322 -10328 -1778
rect -8705 -1778 -8609 -1762
rect -10165 -1890 -8843 -1889
rect -10165 -3210 -10164 -1890
rect -8844 -3210 -8843 -1890
rect -10165 -3211 -8843 -3210
rect -10424 -3338 -10328 -3322
rect -8705 -3322 -8689 -1778
rect -8625 -3322 -8609 -1778
rect -6986 -1778 -6890 -1762
rect -8446 -1890 -7124 -1889
rect -8446 -3210 -8445 -1890
rect -7125 -3210 -7124 -1890
rect -8446 -3211 -7124 -3210
rect -8705 -3338 -8609 -3322
rect -6986 -3322 -6970 -1778
rect -6906 -3322 -6890 -1778
rect -5267 -1778 -5171 -1762
rect -6727 -1890 -5405 -1889
rect -6727 -3210 -6726 -1890
rect -5406 -3210 -5405 -1890
rect -6727 -3211 -5405 -3210
rect -6986 -3338 -6890 -3322
rect -5267 -3322 -5251 -1778
rect -5187 -3322 -5171 -1778
rect -3548 -1778 -3452 -1762
rect -5008 -1890 -3686 -1889
rect -5008 -3210 -5007 -1890
rect -3687 -3210 -3686 -1890
rect -5008 -3211 -3686 -3210
rect -5267 -3338 -5171 -3322
rect -3548 -3322 -3532 -1778
rect -3468 -3322 -3452 -1778
rect -1829 -1778 -1733 -1762
rect -3289 -1890 -1967 -1889
rect -3289 -3210 -3288 -1890
rect -1968 -3210 -1967 -1890
rect -3289 -3211 -1967 -3210
rect -3548 -3338 -3452 -3322
rect -1829 -3322 -1813 -1778
rect -1749 -3322 -1733 -1778
rect -110 -1778 -14 -1762
rect -1570 -1890 -248 -1889
rect -1570 -3210 -1569 -1890
rect -249 -3210 -248 -1890
rect -1570 -3211 -248 -3210
rect -1829 -3338 -1733 -3322
rect -110 -3322 -94 -1778
rect -30 -3322 -14 -1778
rect 1609 -1778 1705 -1762
rect 149 -1890 1471 -1889
rect 149 -3210 150 -1890
rect 1470 -3210 1471 -1890
rect 149 -3211 1471 -3210
rect -110 -3338 -14 -3322
rect 1609 -3322 1625 -1778
rect 1689 -3322 1705 -1778
rect 3328 -1778 3424 -1762
rect 1868 -1890 3190 -1889
rect 1868 -3210 1869 -1890
rect 3189 -3210 3190 -1890
rect 1868 -3211 3190 -3210
rect 1609 -3338 1705 -3322
rect 3328 -3322 3344 -1778
rect 3408 -3322 3424 -1778
rect 5047 -1778 5143 -1762
rect 3587 -1890 4909 -1889
rect 3587 -3210 3588 -1890
rect 4908 -3210 4909 -1890
rect 3587 -3211 4909 -3210
rect 3328 -3338 3424 -3322
rect 5047 -3322 5063 -1778
rect 5127 -3322 5143 -1778
rect 6766 -1778 6862 -1762
rect 5306 -1890 6628 -1889
rect 5306 -3210 5307 -1890
rect 6627 -3210 6628 -1890
rect 5306 -3211 6628 -3210
rect 5047 -3338 5143 -3322
rect 6766 -3322 6782 -1778
rect 6846 -3322 6862 -1778
rect 8485 -1778 8581 -1762
rect 7025 -1890 8347 -1889
rect 7025 -3210 7026 -1890
rect 8346 -3210 8347 -1890
rect 7025 -3211 8347 -3210
rect 6766 -3338 6862 -3322
rect 8485 -3322 8501 -1778
rect 8565 -3322 8581 -1778
rect 10204 -1778 10300 -1762
rect 8744 -1890 10066 -1889
rect 8744 -3210 8745 -1890
rect 10065 -3210 10066 -1890
rect 8744 -3211 10066 -3210
rect 8485 -3338 8581 -3322
rect 10204 -3322 10220 -1778
rect 10284 -3322 10300 -1778
rect 11923 -1778 12019 -1762
rect 10463 -1890 11785 -1889
rect 10463 -3210 10464 -1890
rect 11784 -3210 11785 -1890
rect 10463 -3211 11785 -3210
rect 10204 -3338 10300 -3322
rect 11923 -3322 11939 -1778
rect 12003 -3322 12019 -1778
rect 13642 -1778 13738 -1762
rect 12182 -1890 13504 -1889
rect 12182 -3210 12183 -1890
rect 13503 -3210 13504 -1890
rect 12182 -3211 13504 -3210
rect 11923 -3338 12019 -3322
rect 13642 -3322 13658 -1778
rect 13722 -3322 13738 -1778
rect 15361 -1778 15457 -1762
rect 13901 -1890 15223 -1889
rect 13901 -3210 13902 -1890
rect 15222 -3210 15223 -1890
rect 13901 -3211 15223 -3210
rect 13642 -3338 13738 -3322
rect 15361 -3322 15377 -1778
rect 15441 -3322 15457 -1778
rect 15361 -3338 15457 -3322
rect -13862 -3478 -13766 -3462
rect -15322 -3590 -14000 -3589
rect -15322 -4910 -15321 -3590
rect -14001 -4910 -14000 -3590
rect -15322 -4911 -14000 -4910
rect -13862 -5022 -13846 -3478
rect -13782 -5022 -13766 -3478
rect -12143 -3478 -12047 -3462
rect -13603 -3590 -12281 -3589
rect -13603 -4910 -13602 -3590
rect -12282 -4910 -12281 -3590
rect -13603 -4911 -12281 -4910
rect -13862 -5038 -13766 -5022
rect -12143 -5022 -12127 -3478
rect -12063 -5022 -12047 -3478
rect -10424 -3478 -10328 -3462
rect -11884 -3590 -10562 -3589
rect -11884 -4910 -11883 -3590
rect -10563 -4910 -10562 -3590
rect -11884 -4911 -10562 -4910
rect -12143 -5038 -12047 -5022
rect -10424 -5022 -10408 -3478
rect -10344 -5022 -10328 -3478
rect -8705 -3478 -8609 -3462
rect -10165 -3590 -8843 -3589
rect -10165 -4910 -10164 -3590
rect -8844 -4910 -8843 -3590
rect -10165 -4911 -8843 -4910
rect -10424 -5038 -10328 -5022
rect -8705 -5022 -8689 -3478
rect -8625 -5022 -8609 -3478
rect -6986 -3478 -6890 -3462
rect -8446 -3590 -7124 -3589
rect -8446 -4910 -8445 -3590
rect -7125 -4910 -7124 -3590
rect -8446 -4911 -7124 -4910
rect -8705 -5038 -8609 -5022
rect -6986 -5022 -6970 -3478
rect -6906 -5022 -6890 -3478
rect -5267 -3478 -5171 -3462
rect -6727 -3590 -5405 -3589
rect -6727 -4910 -6726 -3590
rect -5406 -4910 -5405 -3590
rect -6727 -4911 -5405 -4910
rect -6986 -5038 -6890 -5022
rect -5267 -5022 -5251 -3478
rect -5187 -5022 -5171 -3478
rect -3548 -3478 -3452 -3462
rect -5008 -3590 -3686 -3589
rect -5008 -4910 -5007 -3590
rect -3687 -4910 -3686 -3590
rect -5008 -4911 -3686 -4910
rect -5267 -5038 -5171 -5022
rect -3548 -5022 -3532 -3478
rect -3468 -5022 -3452 -3478
rect -1829 -3478 -1733 -3462
rect -3289 -3590 -1967 -3589
rect -3289 -4910 -3288 -3590
rect -1968 -4910 -1967 -3590
rect -3289 -4911 -1967 -4910
rect -3548 -5038 -3452 -5022
rect -1829 -5022 -1813 -3478
rect -1749 -5022 -1733 -3478
rect -110 -3478 -14 -3462
rect -1570 -3590 -248 -3589
rect -1570 -4910 -1569 -3590
rect -249 -4910 -248 -3590
rect -1570 -4911 -248 -4910
rect -1829 -5038 -1733 -5022
rect -110 -5022 -94 -3478
rect -30 -5022 -14 -3478
rect 1609 -3478 1705 -3462
rect 149 -3590 1471 -3589
rect 149 -4910 150 -3590
rect 1470 -4910 1471 -3590
rect 149 -4911 1471 -4910
rect -110 -5038 -14 -5022
rect 1609 -5022 1625 -3478
rect 1689 -5022 1705 -3478
rect 3328 -3478 3424 -3462
rect 1868 -3590 3190 -3589
rect 1868 -4910 1869 -3590
rect 3189 -4910 3190 -3590
rect 1868 -4911 3190 -4910
rect 1609 -5038 1705 -5022
rect 3328 -5022 3344 -3478
rect 3408 -5022 3424 -3478
rect 5047 -3478 5143 -3462
rect 3587 -3590 4909 -3589
rect 3587 -4910 3588 -3590
rect 4908 -4910 4909 -3590
rect 3587 -4911 4909 -4910
rect 3328 -5038 3424 -5022
rect 5047 -5022 5063 -3478
rect 5127 -5022 5143 -3478
rect 6766 -3478 6862 -3462
rect 5306 -3590 6628 -3589
rect 5306 -4910 5307 -3590
rect 6627 -4910 6628 -3590
rect 5306 -4911 6628 -4910
rect 5047 -5038 5143 -5022
rect 6766 -5022 6782 -3478
rect 6846 -5022 6862 -3478
rect 8485 -3478 8581 -3462
rect 7025 -3590 8347 -3589
rect 7025 -4910 7026 -3590
rect 8346 -4910 8347 -3590
rect 7025 -4911 8347 -4910
rect 6766 -5038 6862 -5022
rect 8485 -5022 8501 -3478
rect 8565 -5022 8581 -3478
rect 10204 -3478 10300 -3462
rect 8744 -3590 10066 -3589
rect 8744 -4910 8745 -3590
rect 10065 -4910 10066 -3590
rect 8744 -4911 10066 -4910
rect 8485 -5038 8581 -5022
rect 10204 -5022 10220 -3478
rect 10284 -5022 10300 -3478
rect 11923 -3478 12019 -3462
rect 10463 -3590 11785 -3589
rect 10463 -4910 10464 -3590
rect 11784 -4910 11785 -3590
rect 10463 -4911 11785 -4910
rect 10204 -5038 10300 -5022
rect 11923 -5022 11939 -3478
rect 12003 -5022 12019 -3478
rect 13642 -3478 13738 -3462
rect 12182 -3590 13504 -3589
rect 12182 -4910 12183 -3590
rect 13503 -4910 13504 -3590
rect 12182 -4911 13504 -4910
rect 11923 -5038 12019 -5022
rect 13642 -5022 13658 -3478
rect 13722 -5022 13738 -3478
rect 15361 -3478 15457 -3462
rect 13901 -3590 15223 -3589
rect 13901 -4910 13902 -3590
rect 15222 -4910 15223 -3590
rect 13901 -4911 15223 -4910
rect 13642 -5038 13738 -5022
rect 15361 -5022 15377 -3478
rect 15441 -5022 15457 -3478
rect 15361 -5038 15457 -5022
rect -13862 -5178 -13766 -5162
rect -15322 -5290 -14000 -5289
rect -15322 -6610 -15321 -5290
rect -14001 -6610 -14000 -5290
rect -15322 -6611 -14000 -6610
rect -13862 -6722 -13846 -5178
rect -13782 -6722 -13766 -5178
rect -12143 -5178 -12047 -5162
rect -13603 -5290 -12281 -5289
rect -13603 -6610 -13602 -5290
rect -12282 -6610 -12281 -5290
rect -13603 -6611 -12281 -6610
rect -13862 -6738 -13766 -6722
rect -12143 -6722 -12127 -5178
rect -12063 -6722 -12047 -5178
rect -10424 -5178 -10328 -5162
rect -11884 -5290 -10562 -5289
rect -11884 -6610 -11883 -5290
rect -10563 -6610 -10562 -5290
rect -11884 -6611 -10562 -6610
rect -12143 -6738 -12047 -6722
rect -10424 -6722 -10408 -5178
rect -10344 -6722 -10328 -5178
rect -8705 -5178 -8609 -5162
rect -10165 -5290 -8843 -5289
rect -10165 -6610 -10164 -5290
rect -8844 -6610 -8843 -5290
rect -10165 -6611 -8843 -6610
rect -10424 -6738 -10328 -6722
rect -8705 -6722 -8689 -5178
rect -8625 -6722 -8609 -5178
rect -6986 -5178 -6890 -5162
rect -8446 -5290 -7124 -5289
rect -8446 -6610 -8445 -5290
rect -7125 -6610 -7124 -5290
rect -8446 -6611 -7124 -6610
rect -8705 -6738 -8609 -6722
rect -6986 -6722 -6970 -5178
rect -6906 -6722 -6890 -5178
rect -5267 -5178 -5171 -5162
rect -6727 -5290 -5405 -5289
rect -6727 -6610 -6726 -5290
rect -5406 -6610 -5405 -5290
rect -6727 -6611 -5405 -6610
rect -6986 -6738 -6890 -6722
rect -5267 -6722 -5251 -5178
rect -5187 -6722 -5171 -5178
rect -3548 -5178 -3452 -5162
rect -5008 -5290 -3686 -5289
rect -5008 -6610 -5007 -5290
rect -3687 -6610 -3686 -5290
rect -5008 -6611 -3686 -6610
rect -5267 -6738 -5171 -6722
rect -3548 -6722 -3532 -5178
rect -3468 -6722 -3452 -5178
rect -1829 -5178 -1733 -5162
rect -3289 -5290 -1967 -5289
rect -3289 -6610 -3288 -5290
rect -1968 -6610 -1967 -5290
rect -3289 -6611 -1967 -6610
rect -3548 -6738 -3452 -6722
rect -1829 -6722 -1813 -5178
rect -1749 -6722 -1733 -5178
rect -110 -5178 -14 -5162
rect -1570 -5290 -248 -5289
rect -1570 -6610 -1569 -5290
rect -249 -6610 -248 -5290
rect -1570 -6611 -248 -6610
rect -1829 -6738 -1733 -6722
rect -110 -6722 -94 -5178
rect -30 -6722 -14 -5178
rect 1609 -5178 1705 -5162
rect 149 -5290 1471 -5289
rect 149 -6610 150 -5290
rect 1470 -6610 1471 -5290
rect 149 -6611 1471 -6610
rect -110 -6738 -14 -6722
rect 1609 -6722 1625 -5178
rect 1689 -6722 1705 -5178
rect 3328 -5178 3424 -5162
rect 1868 -5290 3190 -5289
rect 1868 -6610 1869 -5290
rect 3189 -6610 3190 -5290
rect 1868 -6611 3190 -6610
rect 1609 -6738 1705 -6722
rect 3328 -6722 3344 -5178
rect 3408 -6722 3424 -5178
rect 5047 -5178 5143 -5162
rect 3587 -5290 4909 -5289
rect 3587 -6610 3588 -5290
rect 4908 -6610 4909 -5290
rect 3587 -6611 4909 -6610
rect 3328 -6738 3424 -6722
rect 5047 -6722 5063 -5178
rect 5127 -6722 5143 -5178
rect 6766 -5178 6862 -5162
rect 5306 -5290 6628 -5289
rect 5306 -6610 5307 -5290
rect 6627 -6610 6628 -5290
rect 5306 -6611 6628 -6610
rect 5047 -6738 5143 -6722
rect 6766 -6722 6782 -5178
rect 6846 -6722 6862 -5178
rect 8485 -5178 8581 -5162
rect 7025 -5290 8347 -5289
rect 7025 -6610 7026 -5290
rect 8346 -6610 8347 -5290
rect 7025 -6611 8347 -6610
rect 6766 -6738 6862 -6722
rect 8485 -6722 8501 -5178
rect 8565 -6722 8581 -5178
rect 10204 -5178 10300 -5162
rect 8744 -5290 10066 -5289
rect 8744 -6610 8745 -5290
rect 10065 -6610 10066 -5290
rect 8744 -6611 10066 -6610
rect 8485 -6738 8581 -6722
rect 10204 -6722 10220 -5178
rect 10284 -6722 10300 -5178
rect 11923 -5178 12019 -5162
rect 10463 -5290 11785 -5289
rect 10463 -6610 10464 -5290
rect 11784 -6610 11785 -5290
rect 10463 -6611 11785 -6610
rect 10204 -6738 10300 -6722
rect 11923 -6722 11939 -5178
rect 12003 -6722 12019 -5178
rect 13642 -5178 13738 -5162
rect 12182 -5290 13504 -5289
rect 12182 -6610 12183 -5290
rect 13503 -6610 13504 -5290
rect 12182 -6611 13504 -6610
rect 11923 -6738 12019 -6722
rect 13642 -6722 13658 -5178
rect 13722 -6722 13738 -5178
rect 15361 -5178 15457 -5162
rect 13901 -5290 15223 -5289
rect 13901 -6610 13902 -5290
rect 15222 -6610 15223 -5290
rect 13901 -6611 15223 -6610
rect 13642 -6738 13738 -6722
rect 15361 -6722 15377 -5178
rect 15441 -6722 15457 -5178
rect 15361 -6738 15457 -6722
rect -13862 -6878 -13766 -6862
rect -15322 -6990 -14000 -6989
rect -15322 -8310 -15321 -6990
rect -14001 -8310 -14000 -6990
rect -15322 -8311 -14000 -8310
rect -13862 -8422 -13846 -6878
rect -13782 -8422 -13766 -6878
rect -12143 -6878 -12047 -6862
rect -13603 -6990 -12281 -6989
rect -13603 -8310 -13602 -6990
rect -12282 -8310 -12281 -6990
rect -13603 -8311 -12281 -8310
rect -13862 -8438 -13766 -8422
rect -12143 -8422 -12127 -6878
rect -12063 -8422 -12047 -6878
rect -10424 -6878 -10328 -6862
rect -11884 -6990 -10562 -6989
rect -11884 -8310 -11883 -6990
rect -10563 -8310 -10562 -6990
rect -11884 -8311 -10562 -8310
rect -12143 -8438 -12047 -8422
rect -10424 -8422 -10408 -6878
rect -10344 -8422 -10328 -6878
rect -8705 -6878 -8609 -6862
rect -10165 -6990 -8843 -6989
rect -10165 -8310 -10164 -6990
rect -8844 -8310 -8843 -6990
rect -10165 -8311 -8843 -8310
rect -10424 -8438 -10328 -8422
rect -8705 -8422 -8689 -6878
rect -8625 -8422 -8609 -6878
rect -6986 -6878 -6890 -6862
rect -8446 -6990 -7124 -6989
rect -8446 -8310 -8445 -6990
rect -7125 -8310 -7124 -6990
rect -8446 -8311 -7124 -8310
rect -8705 -8438 -8609 -8422
rect -6986 -8422 -6970 -6878
rect -6906 -8422 -6890 -6878
rect -5267 -6878 -5171 -6862
rect -6727 -6990 -5405 -6989
rect -6727 -8310 -6726 -6990
rect -5406 -8310 -5405 -6990
rect -6727 -8311 -5405 -8310
rect -6986 -8438 -6890 -8422
rect -5267 -8422 -5251 -6878
rect -5187 -8422 -5171 -6878
rect -3548 -6878 -3452 -6862
rect -5008 -6990 -3686 -6989
rect -5008 -8310 -5007 -6990
rect -3687 -8310 -3686 -6990
rect -5008 -8311 -3686 -8310
rect -5267 -8438 -5171 -8422
rect -3548 -8422 -3532 -6878
rect -3468 -8422 -3452 -6878
rect -1829 -6878 -1733 -6862
rect -3289 -6990 -1967 -6989
rect -3289 -8310 -3288 -6990
rect -1968 -8310 -1967 -6990
rect -3289 -8311 -1967 -8310
rect -3548 -8438 -3452 -8422
rect -1829 -8422 -1813 -6878
rect -1749 -8422 -1733 -6878
rect -110 -6878 -14 -6862
rect -1570 -6990 -248 -6989
rect -1570 -8310 -1569 -6990
rect -249 -8310 -248 -6990
rect -1570 -8311 -248 -8310
rect -1829 -8438 -1733 -8422
rect -110 -8422 -94 -6878
rect -30 -8422 -14 -6878
rect 1609 -6878 1705 -6862
rect 149 -6990 1471 -6989
rect 149 -8310 150 -6990
rect 1470 -8310 1471 -6990
rect 149 -8311 1471 -8310
rect -110 -8438 -14 -8422
rect 1609 -8422 1625 -6878
rect 1689 -8422 1705 -6878
rect 3328 -6878 3424 -6862
rect 1868 -6990 3190 -6989
rect 1868 -8310 1869 -6990
rect 3189 -8310 3190 -6990
rect 1868 -8311 3190 -8310
rect 1609 -8438 1705 -8422
rect 3328 -8422 3344 -6878
rect 3408 -8422 3424 -6878
rect 5047 -6878 5143 -6862
rect 3587 -6990 4909 -6989
rect 3587 -8310 3588 -6990
rect 4908 -8310 4909 -6990
rect 3587 -8311 4909 -8310
rect 3328 -8438 3424 -8422
rect 5047 -8422 5063 -6878
rect 5127 -8422 5143 -6878
rect 6766 -6878 6862 -6862
rect 5306 -6990 6628 -6989
rect 5306 -8310 5307 -6990
rect 6627 -8310 6628 -6990
rect 5306 -8311 6628 -8310
rect 5047 -8438 5143 -8422
rect 6766 -8422 6782 -6878
rect 6846 -8422 6862 -6878
rect 8485 -6878 8581 -6862
rect 7025 -6990 8347 -6989
rect 7025 -8310 7026 -6990
rect 8346 -8310 8347 -6990
rect 7025 -8311 8347 -8310
rect 6766 -8438 6862 -8422
rect 8485 -8422 8501 -6878
rect 8565 -8422 8581 -6878
rect 10204 -6878 10300 -6862
rect 8744 -6990 10066 -6989
rect 8744 -8310 8745 -6990
rect 10065 -8310 10066 -6990
rect 8744 -8311 10066 -8310
rect 8485 -8438 8581 -8422
rect 10204 -8422 10220 -6878
rect 10284 -8422 10300 -6878
rect 11923 -6878 12019 -6862
rect 10463 -6990 11785 -6989
rect 10463 -8310 10464 -6990
rect 11784 -8310 11785 -6990
rect 10463 -8311 11785 -8310
rect 10204 -8438 10300 -8422
rect 11923 -8422 11939 -6878
rect 12003 -8422 12019 -6878
rect 13642 -6878 13738 -6862
rect 12182 -6990 13504 -6989
rect 12182 -8310 12183 -6990
rect 13503 -8310 13504 -6990
rect 12182 -8311 13504 -8310
rect 11923 -8438 12019 -8422
rect 13642 -8422 13658 -6878
rect 13722 -8422 13738 -6878
rect 15361 -6878 15457 -6862
rect 13901 -6990 15223 -6989
rect 13901 -8310 13902 -6990
rect 15222 -8310 15223 -6990
rect 13901 -8311 15223 -8310
rect 13642 -8438 13738 -8422
rect 15361 -8422 15377 -6878
rect 15441 -8422 15457 -6878
rect 15361 -8438 15457 -8422
rect -13862 -8578 -13766 -8562
rect -15322 -8690 -14000 -8689
rect -15322 -10010 -15321 -8690
rect -14001 -10010 -14000 -8690
rect -15322 -10011 -14000 -10010
rect -13862 -10122 -13846 -8578
rect -13782 -10122 -13766 -8578
rect -12143 -8578 -12047 -8562
rect -13603 -8690 -12281 -8689
rect -13603 -10010 -13602 -8690
rect -12282 -10010 -12281 -8690
rect -13603 -10011 -12281 -10010
rect -13862 -10138 -13766 -10122
rect -12143 -10122 -12127 -8578
rect -12063 -10122 -12047 -8578
rect -10424 -8578 -10328 -8562
rect -11884 -8690 -10562 -8689
rect -11884 -10010 -11883 -8690
rect -10563 -10010 -10562 -8690
rect -11884 -10011 -10562 -10010
rect -12143 -10138 -12047 -10122
rect -10424 -10122 -10408 -8578
rect -10344 -10122 -10328 -8578
rect -8705 -8578 -8609 -8562
rect -10165 -8690 -8843 -8689
rect -10165 -10010 -10164 -8690
rect -8844 -10010 -8843 -8690
rect -10165 -10011 -8843 -10010
rect -10424 -10138 -10328 -10122
rect -8705 -10122 -8689 -8578
rect -8625 -10122 -8609 -8578
rect -6986 -8578 -6890 -8562
rect -8446 -8690 -7124 -8689
rect -8446 -10010 -8445 -8690
rect -7125 -10010 -7124 -8690
rect -8446 -10011 -7124 -10010
rect -8705 -10138 -8609 -10122
rect -6986 -10122 -6970 -8578
rect -6906 -10122 -6890 -8578
rect -5267 -8578 -5171 -8562
rect -6727 -8690 -5405 -8689
rect -6727 -10010 -6726 -8690
rect -5406 -10010 -5405 -8690
rect -6727 -10011 -5405 -10010
rect -6986 -10138 -6890 -10122
rect -5267 -10122 -5251 -8578
rect -5187 -10122 -5171 -8578
rect -3548 -8578 -3452 -8562
rect -5008 -8690 -3686 -8689
rect -5008 -10010 -5007 -8690
rect -3687 -10010 -3686 -8690
rect -5008 -10011 -3686 -10010
rect -5267 -10138 -5171 -10122
rect -3548 -10122 -3532 -8578
rect -3468 -10122 -3452 -8578
rect -1829 -8578 -1733 -8562
rect -3289 -8690 -1967 -8689
rect -3289 -10010 -3288 -8690
rect -1968 -10010 -1967 -8690
rect -3289 -10011 -1967 -10010
rect -3548 -10138 -3452 -10122
rect -1829 -10122 -1813 -8578
rect -1749 -10122 -1733 -8578
rect -110 -8578 -14 -8562
rect -1570 -8690 -248 -8689
rect -1570 -10010 -1569 -8690
rect -249 -10010 -248 -8690
rect -1570 -10011 -248 -10010
rect -1829 -10138 -1733 -10122
rect -110 -10122 -94 -8578
rect -30 -10122 -14 -8578
rect 1609 -8578 1705 -8562
rect 149 -8690 1471 -8689
rect 149 -10010 150 -8690
rect 1470 -10010 1471 -8690
rect 149 -10011 1471 -10010
rect -110 -10138 -14 -10122
rect 1609 -10122 1625 -8578
rect 1689 -10122 1705 -8578
rect 3328 -8578 3424 -8562
rect 1868 -8690 3190 -8689
rect 1868 -10010 1869 -8690
rect 3189 -10010 3190 -8690
rect 1868 -10011 3190 -10010
rect 1609 -10138 1705 -10122
rect 3328 -10122 3344 -8578
rect 3408 -10122 3424 -8578
rect 5047 -8578 5143 -8562
rect 3587 -8690 4909 -8689
rect 3587 -10010 3588 -8690
rect 4908 -10010 4909 -8690
rect 3587 -10011 4909 -10010
rect 3328 -10138 3424 -10122
rect 5047 -10122 5063 -8578
rect 5127 -10122 5143 -8578
rect 6766 -8578 6862 -8562
rect 5306 -8690 6628 -8689
rect 5306 -10010 5307 -8690
rect 6627 -10010 6628 -8690
rect 5306 -10011 6628 -10010
rect 5047 -10138 5143 -10122
rect 6766 -10122 6782 -8578
rect 6846 -10122 6862 -8578
rect 8485 -8578 8581 -8562
rect 7025 -8690 8347 -8689
rect 7025 -10010 7026 -8690
rect 8346 -10010 8347 -8690
rect 7025 -10011 8347 -10010
rect 6766 -10138 6862 -10122
rect 8485 -10122 8501 -8578
rect 8565 -10122 8581 -8578
rect 10204 -8578 10300 -8562
rect 8744 -8690 10066 -8689
rect 8744 -10010 8745 -8690
rect 10065 -10010 10066 -8690
rect 8744 -10011 10066 -10010
rect 8485 -10138 8581 -10122
rect 10204 -10122 10220 -8578
rect 10284 -10122 10300 -8578
rect 11923 -8578 12019 -8562
rect 10463 -8690 11785 -8689
rect 10463 -10010 10464 -8690
rect 11784 -10010 11785 -8690
rect 10463 -10011 11785 -10010
rect 10204 -10138 10300 -10122
rect 11923 -10122 11939 -8578
rect 12003 -10122 12019 -8578
rect 13642 -8578 13738 -8562
rect 12182 -8690 13504 -8689
rect 12182 -10010 12183 -8690
rect 13503 -10010 13504 -8690
rect 12182 -10011 13504 -10010
rect 11923 -10138 12019 -10122
rect 13642 -10122 13658 -8578
rect 13722 -10122 13738 -8578
rect 15361 -8578 15457 -8562
rect 13901 -8690 15223 -8689
rect 13901 -10010 13902 -8690
rect 15222 -10010 15223 -8690
rect 13901 -10011 15223 -10010
rect 13642 -10138 13738 -10122
rect 15361 -10122 15377 -8578
rect 15441 -10122 15457 -8578
rect 15361 -10138 15457 -10122
rect -13862 -10278 -13766 -10262
rect -15322 -10390 -14000 -10389
rect -15322 -11710 -15321 -10390
rect -14001 -11710 -14000 -10390
rect -15322 -11711 -14000 -11710
rect -13862 -11822 -13846 -10278
rect -13782 -11822 -13766 -10278
rect -12143 -10278 -12047 -10262
rect -13603 -10390 -12281 -10389
rect -13603 -11710 -13602 -10390
rect -12282 -11710 -12281 -10390
rect -13603 -11711 -12281 -11710
rect -13862 -11838 -13766 -11822
rect -12143 -11822 -12127 -10278
rect -12063 -11822 -12047 -10278
rect -10424 -10278 -10328 -10262
rect -11884 -10390 -10562 -10389
rect -11884 -11710 -11883 -10390
rect -10563 -11710 -10562 -10390
rect -11884 -11711 -10562 -11710
rect -12143 -11838 -12047 -11822
rect -10424 -11822 -10408 -10278
rect -10344 -11822 -10328 -10278
rect -8705 -10278 -8609 -10262
rect -10165 -10390 -8843 -10389
rect -10165 -11710 -10164 -10390
rect -8844 -11710 -8843 -10390
rect -10165 -11711 -8843 -11710
rect -10424 -11838 -10328 -11822
rect -8705 -11822 -8689 -10278
rect -8625 -11822 -8609 -10278
rect -6986 -10278 -6890 -10262
rect -8446 -10390 -7124 -10389
rect -8446 -11710 -8445 -10390
rect -7125 -11710 -7124 -10390
rect -8446 -11711 -7124 -11710
rect -8705 -11838 -8609 -11822
rect -6986 -11822 -6970 -10278
rect -6906 -11822 -6890 -10278
rect -5267 -10278 -5171 -10262
rect -6727 -10390 -5405 -10389
rect -6727 -11710 -6726 -10390
rect -5406 -11710 -5405 -10390
rect -6727 -11711 -5405 -11710
rect -6986 -11838 -6890 -11822
rect -5267 -11822 -5251 -10278
rect -5187 -11822 -5171 -10278
rect -3548 -10278 -3452 -10262
rect -5008 -10390 -3686 -10389
rect -5008 -11710 -5007 -10390
rect -3687 -11710 -3686 -10390
rect -5008 -11711 -3686 -11710
rect -5267 -11838 -5171 -11822
rect -3548 -11822 -3532 -10278
rect -3468 -11822 -3452 -10278
rect -1829 -10278 -1733 -10262
rect -3289 -10390 -1967 -10389
rect -3289 -11710 -3288 -10390
rect -1968 -11710 -1967 -10390
rect -3289 -11711 -1967 -11710
rect -3548 -11838 -3452 -11822
rect -1829 -11822 -1813 -10278
rect -1749 -11822 -1733 -10278
rect -110 -10278 -14 -10262
rect -1570 -10390 -248 -10389
rect -1570 -11710 -1569 -10390
rect -249 -11710 -248 -10390
rect -1570 -11711 -248 -11710
rect -1829 -11838 -1733 -11822
rect -110 -11822 -94 -10278
rect -30 -11822 -14 -10278
rect 1609 -10278 1705 -10262
rect 149 -10390 1471 -10389
rect 149 -11710 150 -10390
rect 1470 -11710 1471 -10390
rect 149 -11711 1471 -11710
rect -110 -11838 -14 -11822
rect 1609 -11822 1625 -10278
rect 1689 -11822 1705 -10278
rect 3328 -10278 3424 -10262
rect 1868 -10390 3190 -10389
rect 1868 -11710 1869 -10390
rect 3189 -11710 3190 -10390
rect 1868 -11711 3190 -11710
rect 1609 -11838 1705 -11822
rect 3328 -11822 3344 -10278
rect 3408 -11822 3424 -10278
rect 5047 -10278 5143 -10262
rect 3587 -10390 4909 -10389
rect 3587 -11710 3588 -10390
rect 4908 -11710 4909 -10390
rect 3587 -11711 4909 -11710
rect 3328 -11838 3424 -11822
rect 5047 -11822 5063 -10278
rect 5127 -11822 5143 -10278
rect 6766 -10278 6862 -10262
rect 5306 -10390 6628 -10389
rect 5306 -11710 5307 -10390
rect 6627 -11710 6628 -10390
rect 5306 -11711 6628 -11710
rect 5047 -11838 5143 -11822
rect 6766 -11822 6782 -10278
rect 6846 -11822 6862 -10278
rect 8485 -10278 8581 -10262
rect 7025 -10390 8347 -10389
rect 7025 -11710 7026 -10390
rect 8346 -11710 8347 -10390
rect 7025 -11711 8347 -11710
rect 6766 -11838 6862 -11822
rect 8485 -11822 8501 -10278
rect 8565 -11822 8581 -10278
rect 10204 -10278 10300 -10262
rect 8744 -10390 10066 -10389
rect 8744 -11710 8745 -10390
rect 10065 -11710 10066 -10390
rect 8744 -11711 10066 -11710
rect 8485 -11838 8581 -11822
rect 10204 -11822 10220 -10278
rect 10284 -11822 10300 -10278
rect 11923 -10278 12019 -10262
rect 10463 -10390 11785 -10389
rect 10463 -11710 10464 -10390
rect 11784 -11710 11785 -10390
rect 10463 -11711 11785 -11710
rect 10204 -11838 10300 -11822
rect 11923 -11822 11939 -10278
rect 12003 -11822 12019 -10278
rect 13642 -10278 13738 -10262
rect 12182 -10390 13504 -10389
rect 12182 -11710 12183 -10390
rect 13503 -11710 13504 -10390
rect 12182 -11711 13504 -11710
rect 11923 -11838 12019 -11822
rect 13642 -11822 13658 -10278
rect 13722 -11822 13738 -10278
rect 15361 -10278 15457 -10262
rect 13901 -10390 15223 -10389
rect 13901 -11710 13902 -10390
rect 15222 -11710 15223 -10390
rect 13901 -11711 15223 -11710
rect 13642 -11838 13738 -11822
rect 15361 -11822 15377 -10278
rect 15441 -11822 15457 -10278
rect 15361 -11838 15457 -11822
rect -13862 -11978 -13766 -11962
rect -15322 -12090 -14000 -12089
rect -15322 -13410 -15321 -12090
rect -14001 -13410 -14000 -12090
rect -15322 -13411 -14000 -13410
rect -13862 -13522 -13846 -11978
rect -13782 -13522 -13766 -11978
rect -12143 -11978 -12047 -11962
rect -13603 -12090 -12281 -12089
rect -13603 -13410 -13602 -12090
rect -12282 -13410 -12281 -12090
rect -13603 -13411 -12281 -13410
rect -13862 -13538 -13766 -13522
rect -12143 -13522 -12127 -11978
rect -12063 -13522 -12047 -11978
rect -10424 -11978 -10328 -11962
rect -11884 -12090 -10562 -12089
rect -11884 -13410 -11883 -12090
rect -10563 -13410 -10562 -12090
rect -11884 -13411 -10562 -13410
rect -12143 -13538 -12047 -13522
rect -10424 -13522 -10408 -11978
rect -10344 -13522 -10328 -11978
rect -8705 -11978 -8609 -11962
rect -10165 -12090 -8843 -12089
rect -10165 -13410 -10164 -12090
rect -8844 -13410 -8843 -12090
rect -10165 -13411 -8843 -13410
rect -10424 -13538 -10328 -13522
rect -8705 -13522 -8689 -11978
rect -8625 -13522 -8609 -11978
rect -6986 -11978 -6890 -11962
rect -8446 -12090 -7124 -12089
rect -8446 -13410 -8445 -12090
rect -7125 -13410 -7124 -12090
rect -8446 -13411 -7124 -13410
rect -8705 -13538 -8609 -13522
rect -6986 -13522 -6970 -11978
rect -6906 -13522 -6890 -11978
rect -5267 -11978 -5171 -11962
rect -6727 -12090 -5405 -12089
rect -6727 -13410 -6726 -12090
rect -5406 -13410 -5405 -12090
rect -6727 -13411 -5405 -13410
rect -6986 -13538 -6890 -13522
rect -5267 -13522 -5251 -11978
rect -5187 -13522 -5171 -11978
rect -3548 -11978 -3452 -11962
rect -5008 -12090 -3686 -12089
rect -5008 -13410 -5007 -12090
rect -3687 -13410 -3686 -12090
rect -5008 -13411 -3686 -13410
rect -5267 -13538 -5171 -13522
rect -3548 -13522 -3532 -11978
rect -3468 -13522 -3452 -11978
rect -1829 -11978 -1733 -11962
rect -3289 -12090 -1967 -12089
rect -3289 -13410 -3288 -12090
rect -1968 -13410 -1967 -12090
rect -3289 -13411 -1967 -13410
rect -3548 -13538 -3452 -13522
rect -1829 -13522 -1813 -11978
rect -1749 -13522 -1733 -11978
rect -110 -11978 -14 -11962
rect -1570 -12090 -248 -12089
rect -1570 -13410 -1569 -12090
rect -249 -13410 -248 -12090
rect -1570 -13411 -248 -13410
rect -1829 -13538 -1733 -13522
rect -110 -13522 -94 -11978
rect -30 -13522 -14 -11978
rect 1609 -11978 1705 -11962
rect 149 -12090 1471 -12089
rect 149 -13410 150 -12090
rect 1470 -13410 1471 -12090
rect 149 -13411 1471 -13410
rect -110 -13538 -14 -13522
rect 1609 -13522 1625 -11978
rect 1689 -13522 1705 -11978
rect 3328 -11978 3424 -11962
rect 1868 -12090 3190 -12089
rect 1868 -13410 1869 -12090
rect 3189 -13410 3190 -12090
rect 1868 -13411 3190 -13410
rect 1609 -13538 1705 -13522
rect 3328 -13522 3344 -11978
rect 3408 -13522 3424 -11978
rect 5047 -11978 5143 -11962
rect 3587 -12090 4909 -12089
rect 3587 -13410 3588 -12090
rect 4908 -13410 4909 -12090
rect 3587 -13411 4909 -13410
rect 3328 -13538 3424 -13522
rect 5047 -13522 5063 -11978
rect 5127 -13522 5143 -11978
rect 6766 -11978 6862 -11962
rect 5306 -12090 6628 -12089
rect 5306 -13410 5307 -12090
rect 6627 -13410 6628 -12090
rect 5306 -13411 6628 -13410
rect 5047 -13538 5143 -13522
rect 6766 -13522 6782 -11978
rect 6846 -13522 6862 -11978
rect 8485 -11978 8581 -11962
rect 7025 -12090 8347 -12089
rect 7025 -13410 7026 -12090
rect 8346 -13410 8347 -12090
rect 7025 -13411 8347 -13410
rect 6766 -13538 6862 -13522
rect 8485 -13522 8501 -11978
rect 8565 -13522 8581 -11978
rect 10204 -11978 10300 -11962
rect 8744 -12090 10066 -12089
rect 8744 -13410 8745 -12090
rect 10065 -13410 10066 -12090
rect 8744 -13411 10066 -13410
rect 8485 -13538 8581 -13522
rect 10204 -13522 10220 -11978
rect 10284 -13522 10300 -11978
rect 11923 -11978 12019 -11962
rect 10463 -12090 11785 -12089
rect 10463 -13410 10464 -12090
rect 11784 -13410 11785 -12090
rect 10463 -13411 11785 -13410
rect 10204 -13538 10300 -13522
rect 11923 -13522 11939 -11978
rect 12003 -13522 12019 -11978
rect 13642 -11978 13738 -11962
rect 12182 -12090 13504 -12089
rect 12182 -13410 12183 -12090
rect 13503 -13410 13504 -12090
rect 12182 -13411 13504 -13410
rect 11923 -13538 12019 -13522
rect 13642 -13522 13658 -11978
rect 13722 -13522 13738 -11978
rect 15361 -11978 15457 -11962
rect 13901 -12090 15223 -12089
rect 13901 -13410 13902 -12090
rect 15222 -13410 15223 -12090
rect 13901 -13411 15223 -13410
rect 13642 -13538 13738 -13522
rect 15361 -13522 15377 -11978
rect 15441 -13522 15457 -11978
rect 15361 -13538 15457 -13522
rect -13862 -13678 -13766 -13662
rect -15322 -13790 -14000 -13789
rect -15322 -15110 -15321 -13790
rect -14001 -15110 -14000 -13790
rect -15322 -15111 -14000 -15110
rect -13862 -15222 -13846 -13678
rect -13782 -15222 -13766 -13678
rect -12143 -13678 -12047 -13662
rect -13603 -13790 -12281 -13789
rect -13603 -15110 -13602 -13790
rect -12282 -15110 -12281 -13790
rect -13603 -15111 -12281 -15110
rect -13862 -15238 -13766 -15222
rect -12143 -15222 -12127 -13678
rect -12063 -15222 -12047 -13678
rect -10424 -13678 -10328 -13662
rect -11884 -13790 -10562 -13789
rect -11884 -15110 -11883 -13790
rect -10563 -15110 -10562 -13790
rect -11884 -15111 -10562 -15110
rect -12143 -15238 -12047 -15222
rect -10424 -15222 -10408 -13678
rect -10344 -15222 -10328 -13678
rect -8705 -13678 -8609 -13662
rect -10165 -13790 -8843 -13789
rect -10165 -15110 -10164 -13790
rect -8844 -15110 -8843 -13790
rect -10165 -15111 -8843 -15110
rect -10424 -15238 -10328 -15222
rect -8705 -15222 -8689 -13678
rect -8625 -15222 -8609 -13678
rect -6986 -13678 -6890 -13662
rect -8446 -13790 -7124 -13789
rect -8446 -15110 -8445 -13790
rect -7125 -15110 -7124 -13790
rect -8446 -15111 -7124 -15110
rect -8705 -15238 -8609 -15222
rect -6986 -15222 -6970 -13678
rect -6906 -15222 -6890 -13678
rect -5267 -13678 -5171 -13662
rect -6727 -13790 -5405 -13789
rect -6727 -15110 -6726 -13790
rect -5406 -15110 -5405 -13790
rect -6727 -15111 -5405 -15110
rect -6986 -15238 -6890 -15222
rect -5267 -15222 -5251 -13678
rect -5187 -15222 -5171 -13678
rect -3548 -13678 -3452 -13662
rect -5008 -13790 -3686 -13789
rect -5008 -15110 -5007 -13790
rect -3687 -15110 -3686 -13790
rect -5008 -15111 -3686 -15110
rect -5267 -15238 -5171 -15222
rect -3548 -15222 -3532 -13678
rect -3468 -15222 -3452 -13678
rect -1829 -13678 -1733 -13662
rect -3289 -13790 -1967 -13789
rect -3289 -15110 -3288 -13790
rect -1968 -15110 -1967 -13790
rect -3289 -15111 -1967 -15110
rect -3548 -15238 -3452 -15222
rect -1829 -15222 -1813 -13678
rect -1749 -15222 -1733 -13678
rect -110 -13678 -14 -13662
rect -1570 -13790 -248 -13789
rect -1570 -15110 -1569 -13790
rect -249 -15110 -248 -13790
rect -1570 -15111 -248 -15110
rect -1829 -15238 -1733 -15222
rect -110 -15222 -94 -13678
rect -30 -15222 -14 -13678
rect 1609 -13678 1705 -13662
rect 149 -13790 1471 -13789
rect 149 -15110 150 -13790
rect 1470 -15110 1471 -13790
rect 149 -15111 1471 -15110
rect -110 -15238 -14 -15222
rect 1609 -15222 1625 -13678
rect 1689 -15222 1705 -13678
rect 3328 -13678 3424 -13662
rect 1868 -13790 3190 -13789
rect 1868 -15110 1869 -13790
rect 3189 -15110 3190 -13790
rect 1868 -15111 3190 -15110
rect 1609 -15238 1705 -15222
rect 3328 -15222 3344 -13678
rect 3408 -15222 3424 -13678
rect 5047 -13678 5143 -13662
rect 3587 -13790 4909 -13789
rect 3587 -15110 3588 -13790
rect 4908 -15110 4909 -13790
rect 3587 -15111 4909 -15110
rect 3328 -15238 3424 -15222
rect 5047 -15222 5063 -13678
rect 5127 -15222 5143 -13678
rect 6766 -13678 6862 -13662
rect 5306 -13790 6628 -13789
rect 5306 -15110 5307 -13790
rect 6627 -15110 6628 -13790
rect 5306 -15111 6628 -15110
rect 5047 -15238 5143 -15222
rect 6766 -15222 6782 -13678
rect 6846 -15222 6862 -13678
rect 8485 -13678 8581 -13662
rect 7025 -13790 8347 -13789
rect 7025 -15110 7026 -13790
rect 8346 -15110 8347 -13790
rect 7025 -15111 8347 -15110
rect 6766 -15238 6862 -15222
rect 8485 -15222 8501 -13678
rect 8565 -15222 8581 -13678
rect 10204 -13678 10300 -13662
rect 8744 -13790 10066 -13789
rect 8744 -15110 8745 -13790
rect 10065 -15110 10066 -13790
rect 8744 -15111 10066 -15110
rect 8485 -15238 8581 -15222
rect 10204 -15222 10220 -13678
rect 10284 -15222 10300 -13678
rect 11923 -13678 12019 -13662
rect 10463 -13790 11785 -13789
rect 10463 -15110 10464 -13790
rect 11784 -15110 11785 -13790
rect 10463 -15111 11785 -15110
rect 10204 -15238 10300 -15222
rect 11923 -15222 11939 -13678
rect 12003 -15222 12019 -13678
rect 13642 -13678 13738 -13662
rect 12182 -13790 13504 -13789
rect 12182 -15110 12183 -13790
rect 13503 -15110 13504 -13790
rect 12182 -15111 13504 -15110
rect 11923 -15238 12019 -15222
rect 13642 -15222 13658 -13678
rect 13722 -15222 13738 -13678
rect 15361 -13678 15457 -13662
rect 13901 -13790 15223 -13789
rect 13901 -15110 13902 -13790
rect 15222 -15110 15223 -13790
rect 13901 -15111 15223 -15110
rect 13642 -15238 13738 -15222
rect 15361 -15222 15377 -13678
rect 15441 -15222 15457 -13678
rect 15361 -15238 15457 -15222
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 13762 13650 15362 15250
string parameters w 7.00 l 7.00 val 103.32 carea 2.00 cperi 0.19 nx 18 ny 18 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
