magic
tech sky130A
timestamp 1622084130
<< viali >>
rect 232 -28 256 -5
rect 282 -29 306 -5
<< metal1 >>
rect 130 112 201 160
rect 152 -5 262 -2
rect 152 -28 232 -5
rect 256 -28 262 -5
rect 152 -32 262 -28
rect 276 -5 359 -2
rect 276 -29 282 -5
rect 306 -29 359 -5
rect 276 -32 359 -29
rect 91 -160 203 -112
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1620951057
transform 1 0 325 0 1 -136
box -19 -24 65 296
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1620951057
transform 1 0 197 0 1 -136
box -19 -24 157 296
<< labels >>
flabel metal1 143 135 145 136 1 FreeSans 240 0 0 0 VDD
flabel metal1 139 -137 142 -135 1 FreeSans 240 0 0 0 VSS
flabel metal1 166 -19 169 -16 1 FreeSans 240 0 0 0 A
flabel metal1 336 -17 338 -15 1 FreeSans 240 0 0 0 Y
<< end >>
