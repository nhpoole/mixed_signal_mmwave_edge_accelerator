magic
tech sky130A
magscale 1 2
timestamp 1622230511
<< viali >>
rect 73 497 107 531
rect 1519 414 1561 456
rect -202 290 -154 338
rect 1835 283 1869 317
<< metal1 >>
rect 1698 570 2104 668
rect 61 531 119 537
rect 61 530 73 531
rect -366 498 73 530
rect 61 497 73 498
rect 107 497 119 531
rect 61 491 119 497
rect 1507 456 1980 462
rect 1507 414 1519 456
rect 1561 414 1980 456
rect 1507 408 1980 414
rect -342 338 -142 344
rect -342 290 -202 338
rect -154 290 -142 338
rect 1186 314 1192 378
rect 1256 314 1262 378
rect 1823 322 1881 323
rect 1823 317 2062 322
rect -342 284 -142 290
rect 1823 283 1835 317
rect 1869 283 2062 317
rect 1823 278 2062 283
rect 1823 277 1881 278
rect 1858 22 2116 118
<< via1 >>
rect 1192 314 1256 378
<< metal2 >>
rect 1192 378 1256 384
rect 1256 314 1460 378
rect 1192 308 1256 314
rect 1396 -118 1460 314
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_0
timestamp 1620951057
transform 1 0 -224 0 1 72
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1620951057
transform 1 0 -316 0 1 72
box -38 -48 130 592
<< labels >>
flabel metal1 -300 312 -294 320 1 FreeSans 480 0 0 0 CLK
flabel metal1 -320 512 -312 516 1 FreeSans 480 0 0 0 D
flabel metal2 1414 -50 1424 -42 1 FreeSans 480 0 0 0 RN
flabel metal1 1948 434 1956 440 1 FreeSans 480 0 0 0 Q
flabel metal1 2002 298 2010 304 1 FreeSans 480 0 0 0 QB
flabel metal1 2052 604 2060 610 1 FreeSans 480 0 0 0 VDD
flabel metal1 2048 68 2066 76 1 FreeSans 480 0 0 0 VSS
<< end >>
