magic
tech sky130A
magscale 1 2
timestamp 1620882364
<< locali >>
rect 668 780 800 798
rect 668 694 718 780
rect 780 694 800 780
rect 668 682 800 694
<< viali >>
rect 718 694 780 780
rect -98 215 -50 263
rect 246 215 294 263
<< metal1 >>
rect 864 922 1234 958
rect -234 886 1234 922
rect -234 874 934 886
rect -234 263 -186 874
rect 668 780 800 798
rect 668 760 718 780
rect 98 712 718 760
rect 98 534 146 712
rect 668 694 718 712
rect 780 760 800 780
rect 780 712 878 760
rect 940 754 988 806
rect 1062 754 1068 756
rect 780 694 800 712
rect 668 682 800 694
rect 940 706 1068 754
rect 940 672 988 706
rect 1062 704 1068 706
rect 1120 704 1126 756
rect 868 578 940 604
rect 1162 578 1234 886
rect 868 506 1234 578
rect 620 352 626 404
rect 678 352 684 404
rect -104 263 -44 275
rect -234 215 -98 263
rect -50 215 -44 263
rect -104 203 -44 215
rect 240 263 300 275
rect 240 215 246 263
rect 294 215 418 263
rect 240 203 300 215
rect 628 162 676 352
rect 870 306 942 506
rect 870 234 1232 306
rect 628 114 878 162
rect 1062 158 1068 160
rect 940 110 1068 158
rect 1062 108 1068 110
rect 1120 108 1126 160
rect 1160 42 1232 234
rect -76 -48 -70 4
rect -18 -48 -12 4
rect 880 -30 1232 42
<< via1 >>
rect 1068 704 1120 756
rect 626 352 678 404
rect 1068 108 1120 160
rect -70 -48 -18 4
<< metal2 >>
rect 1068 756 1120 762
rect 1120 706 1330 754
rect 1068 698 1120 704
rect 626 404 678 410
rect 1282 402 1330 706
rect 678 354 1330 402
rect 626 346 678 352
rect 1068 160 1120 166
rect 1120 110 1370 158
rect 1068 102 1120 108
rect -70 4 -18 10
rect -70 -54 -18 -48
rect -68 -180 -20 -54
rect 1322 -180 1370 110
rect -68 -228 1370 -180
use sky130_fd_pr__pfet_01v8_hvt_UU5H43  sky130_fd_pr__pfet_01v8_hvt_UU5H43_0
timestamp 1620878641
transform 1 0 907 0 1 739
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_82JX4H  sky130_fd_pr__nfet_01v8_82JX4H_0
timestamp 1620878641
transform 1 0 909 0 1 135
box -211 -275 211 275
use inv1  inv1_0
timestamp 1608267076
transform 1 0 0 0 1 0
box -101 -48 314 592
<< labels >>
flabel metal1 -214 658 -214 658 1 FreeSans 480 0 0 0 in
port 1 n
flabel metal2 1312 536 1312 536 1 FreeSans 480 0 0 0 out
port 3 n
flabel metal1 326 734 326 734 1 FreeSans 480 0 0 0 VDD
port 4 n
flabel metal2 512 -206 512 -206 1 FreeSans 480 0 0 0 VSS
port 5 n
flabel metal1 392 236 392 236 1 FreeSans 480 0 0 0 out2
port 6 n
<< end >>
