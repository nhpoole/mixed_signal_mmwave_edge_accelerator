magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -194 -500 194 500
<< nwell >>
rect -194 -500 194 500
<< pmoshvt >>
rect -100 -400 100 400
<< pdiff >>
rect -158 388 -100 400
rect -158 -388 -146 388
rect -112 -388 -100 388
rect -158 -400 -100 -388
rect 100 388 158 400
rect 100 -388 112 388
rect 146 -388 158 388
rect 100 -400 158 -388
<< pdiffc >>
rect -146 -388 -112 388
rect 112 -388 146 388
<< poly >>
rect -66 481 66 497
rect -66 464 -50 481
rect -100 447 -50 464
rect 50 464 66 481
rect 50 447 100 464
rect -100 400 100 447
rect -100 -447 100 -400
rect -100 -464 -50 -447
rect -66 -481 -50 -464
rect 50 -464 100 -447
rect 50 -481 66 -464
rect -66 -497 66 -481
<< polycont >>
rect -50 447 50 481
rect -50 -481 50 -447
<< locali >>
rect -66 447 -50 481
rect 50 447 66 481
rect -146 388 -112 404
rect -146 -404 -112 -388
rect 112 388 146 404
rect 112 -404 146 -388
rect -66 -481 -50 -447
rect 50 -481 66 -447
<< viali >>
rect -42 447 42 481
rect -146 -388 -112 388
rect 112 -388 146 388
rect -42 -481 42 -447
<< metal1 >>
rect -54 481 54 487
rect -54 447 -42 481
rect 42 447 54 481
rect -54 441 54 447
rect -152 388 -106 400
rect -152 -388 -146 388
rect -112 -388 -106 388
rect -152 -400 -106 -388
rect 106 388 152 400
rect 106 -388 112 388
rect 146 -388 152 388
rect 106 -400 152 -388
rect -54 -447 54 -441
rect -54 -481 -42 -447
rect 42 -481 54 -447
rect -54 -487 54 -481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string parameters w 4 l 1 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
