magic
tech sky130A
magscale 1 2
timestamp 1620412613
<< nwell >>
rect -8209 -400 8209 400
<< pmoslvt >>
rect -8115 -300 -7155 300
rect -7097 -300 -6137 300
rect -6079 -300 -5119 300
rect -5061 -300 -4101 300
rect -4043 -300 -3083 300
rect -3025 -300 -2065 300
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
rect 2065 -300 3025 300
rect 3083 -300 4043 300
rect 4101 -300 5061 300
rect 5119 -300 6079 300
rect 6137 -300 7097 300
rect 7155 -300 8115 300
<< pdiff >>
rect -8173 288 -8115 300
rect -8173 -288 -8161 288
rect -8127 -288 -8115 288
rect -8173 -300 -8115 -288
rect -7155 288 -7097 300
rect -7155 -288 -7143 288
rect -7109 -288 -7097 288
rect -7155 -300 -7097 -288
rect -6137 288 -6079 300
rect -6137 -288 -6125 288
rect -6091 -288 -6079 288
rect -6137 -300 -6079 -288
rect -5119 288 -5061 300
rect -5119 -288 -5107 288
rect -5073 -288 -5061 288
rect -5119 -300 -5061 -288
rect -4101 288 -4043 300
rect -4101 -288 -4089 288
rect -4055 -288 -4043 288
rect -4101 -300 -4043 -288
rect -3083 288 -3025 300
rect -3083 -288 -3071 288
rect -3037 -288 -3025 288
rect -3083 -300 -3025 -288
rect -2065 288 -2007 300
rect -2065 -288 -2053 288
rect -2019 -288 -2007 288
rect -2065 -300 -2007 -288
rect -1047 288 -989 300
rect -1047 -288 -1035 288
rect -1001 -288 -989 288
rect -1047 -300 -989 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 989 288 1047 300
rect 989 -288 1001 288
rect 1035 -288 1047 288
rect 989 -300 1047 -288
rect 2007 288 2065 300
rect 2007 -288 2019 288
rect 2053 -288 2065 288
rect 2007 -300 2065 -288
rect 3025 288 3083 300
rect 3025 -288 3037 288
rect 3071 -288 3083 288
rect 3025 -300 3083 -288
rect 4043 288 4101 300
rect 4043 -288 4055 288
rect 4089 -288 4101 288
rect 4043 -300 4101 -288
rect 5061 288 5119 300
rect 5061 -288 5073 288
rect 5107 -288 5119 288
rect 5061 -300 5119 -288
rect 6079 288 6137 300
rect 6079 -288 6091 288
rect 6125 -288 6137 288
rect 6079 -300 6137 -288
rect 7097 288 7155 300
rect 7097 -288 7109 288
rect 7143 -288 7155 288
rect 7097 -300 7155 -288
rect 8115 288 8173 300
rect 8115 -288 8127 288
rect 8161 -288 8173 288
rect 8115 -300 8173 -288
<< pdiffc >>
rect -8161 -288 -8127 288
rect -7143 -288 -7109 288
rect -6125 -288 -6091 288
rect -5107 -288 -5073 288
rect -4089 -288 -4055 288
rect -3071 -288 -3037 288
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect 3037 -288 3071 288
rect 4055 -288 4089 288
rect 5073 -288 5107 288
rect 6091 -288 6125 288
rect 7109 -288 7143 288
rect 8127 -288 8161 288
<< poly >>
rect -7929 381 -7341 397
rect -7929 364 -7913 381
rect -8115 347 -7913 364
rect -7357 364 -7341 381
rect -6911 381 -6323 397
rect -6911 364 -6895 381
rect -7357 347 -7155 364
rect -8115 300 -7155 347
rect -7097 347 -6895 364
rect -6339 364 -6323 381
rect -5893 381 -5305 397
rect -5893 364 -5877 381
rect -6339 347 -6137 364
rect -7097 300 -6137 347
rect -6079 347 -5877 364
rect -5321 364 -5305 381
rect -4875 381 -4287 397
rect -4875 364 -4859 381
rect -5321 347 -5119 364
rect -6079 300 -5119 347
rect -5061 347 -4859 364
rect -4303 364 -4287 381
rect -3857 381 -3269 397
rect -3857 364 -3841 381
rect -4303 347 -4101 364
rect -5061 300 -4101 347
rect -4043 347 -3841 364
rect -3285 364 -3269 381
rect -2839 381 -2251 397
rect -2839 364 -2823 381
rect -3285 347 -3083 364
rect -4043 300 -3083 347
rect -3025 347 -2823 364
rect -2267 364 -2251 381
rect -1821 381 -1233 397
rect -1821 364 -1805 381
rect -2267 347 -2065 364
rect -3025 300 -2065 347
rect -2007 347 -1805 364
rect -1249 364 -1233 381
rect -803 381 -215 397
rect -803 364 -787 381
rect -1249 347 -1047 364
rect -2007 300 -1047 347
rect -989 347 -787 364
rect -231 364 -215 381
rect 215 381 803 397
rect 215 364 231 381
rect -231 347 -29 364
rect -989 300 -29 347
rect 29 347 231 364
rect 787 364 803 381
rect 1233 381 1821 397
rect 1233 364 1249 381
rect 787 347 989 364
rect 29 300 989 347
rect 1047 347 1249 364
rect 1805 364 1821 381
rect 2251 381 2839 397
rect 2251 364 2267 381
rect 1805 347 2007 364
rect 1047 300 2007 347
rect 2065 347 2267 364
rect 2823 364 2839 381
rect 3269 381 3857 397
rect 3269 364 3285 381
rect 2823 347 3025 364
rect 2065 300 3025 347
rect 3083 347 3285 364
rect 3841 364 3857 381
rect 4287 381 4875 397
rect 4287 364 4303 381
rect 3841 347 4043 364
rect 3083 300 4043 347
rect 4101 347 4303 364
rect 4859 364 4875 381
rect 5305 381 5893 397
rect 5305 364 5321 381
rect 4859 347 5061 364
rect 4101 300 5061 347
rect 5119 347 5321 364
rect 5877 364 5893 381
rect 6323 381 6911 397
rect 6323 364 6339 381
rect 5877 347 6079 364
rect 5119 300 6079 347
rect 6137 347 6339 364
rect 6895 364 6911 381
rect 7341 381 7929 397
rect 7341 364 7357 381
rect 6895 347 7097 364
rect 6137 300 7097 347
rect 7155 347 7357 364
rect 7913 364 7929 381
rect 7913 347 8115 364
rect 7155 300 8115 347
rect -8115 -347 -7155 -300
rect -8115 -364 -7913 -347
rect -7929 -381 -7913 -364
rect -7357 -364 -7155 -347
rect -7097 -347 -6137 -300
rect -7097 -364 -6895 -347
rect -7357 -381 -7341 -364
rect -7929 -397 -7341 -381
rect -6911 -381 -6895 -364
rect -6339 -364 -6137 -347
rect -6079 -347 -5119 -300
rect -6079 -364 -5877 -347
rect -6339 -381 -6323 -364
rect -6911 -397 -6323 -381
rect -5893 -381 -5877 -364
rect -5321 -364 -5119 -347
rect -5061 -347 -4101 -300
rect -5061 -364 -4859 -347
rect -5321 -381 -5305 -364
rect -5893 -397 -5305 -381
rect -4875 -381 -4859 -364
rect -4303 -364 -4101 -347
rect -4043 -347 -3083 -300
rect -4043 -364 -3841 -347
rect -4303 -381 -4287 -364
rect -4875 -397 -4287 -381
rect -3857 -381 -3841 -364
rect -3285 -364 -3083 -347
rect -3025 -347 -2065 -300
rect -3025 -364 -2823 -347
rect -3285 -381 -3269 -364
rect -3857 -397 -3269 -381
rect -2839 -381 -2823 -364
rect -2267 -364 -2065 -347
rect -2007 -347 -1047 -300
rect -2007 -364 -1805 -347
rect -2267 -381 -2251 -364
rect -2839 -397 -2251 -381
rect -1821 -381 -1805 -364
rect -1249 -364 -1047 -347
rect -989 -347 -29 -300
rect -989 -364 -787 -347
rect -1249 -381 -1233 -364
rect -1821 -397 -1233 -381
rect -803 -381 -787 -364
rect -231 -364 -29 -347
rect 29 -347 989 -300
rect 29 -364 231 -347
rect -231 -381 -215 -364
rect -803 -397 -215 -381
rect 215 -381 231 -364
rect 787 -364 989 -347
rect 1047 -347 2007 -300
rect 1047 -364 1249 -347
rect 787 -381 803 -364
rect 215 -397 803 -381
rect 1233 -381 1249 -364
rect 1805 -364 2007 -347
rect 2065 -347 3025 -300
rect 2065 -364 2267 -347
rect 1805 -381 1821 -364
rect 1233 -397 1821 -381
rect 2251 -381 2267 -364
rect 2823 -364 3025 -347
rect 3083 -347 4043 -300
rect 3083 -364 3285 -347
rect 2823 -381 2839 -364
rect 2251 -397 2839 -381
rect 3269 -381 3285 -364
rect 3841 -364 4043 -347
rect 4101 -347 5061 -300
rect 4101 -364 4303 -347
rect 3841 -381 3857 -364
rect 3269 -397 3857 -381
rect 4287 -381 4303 -364
rect 4859 -364 5061 -347
rect 5119 -347 6079 -300
rect 5119 -364 5321 -347
rect 4859 -381 4875 -364
rect 4287 -397 4875 -381
rect 5305 -381 5321 -364
rect 5877 -364 6079 -347
rect 6137 -347 7097 -300
rect 6137 -364 6339 -347
rect 5877 -381 5893 -364
rect 5305 -397 5893 -381
rect 6323 -381 6339 -364
rect 6895 -364 7097 -347
rect 7155 -347 8115 -300
rect 7155 -364 7357 -347
rect 6895 -381 6911 -364
rect 6323 -397 6911 -381
rect 7341 -381 7357 -364
rect 7913 -364 8115 -347
rect 7913 -381 7929 -364
rect 7341 -397 7929 -381
<< polycont >>
rect -7913 347 -7357 381
rect -6895 347 -6339 381
rect -5877 347 -5321 381
rect -4859 347 -4303 381
rect -3841 347 -3285 381
rect -2823 347 -2267 381
rect -1805 347 -1249 381
rect -787 347 -231 381
rect 231 347 787 381
rect 1249 347 1805 381
rect 2267 347 2823 381
rect 3285 347 3841 381
rect 4303 347 4859 381
rect 5321 347 5877 381
rect 6339 347 6895 381
rect 7357 347 7913 381
rect -7913 -381 -7357 -347
rect -6895 -381 -6339 -347
rect -5877 -381 -5321 -347
rect -4859 -381 -4303 -347
rect -3841 -381 -3285 -347
rect -2823 -381 -2267 -347
rect -1805 -381 -1249 -347
rect -787 -381 -231 -347
rect 231 -381 787 -347
rect 1249 -381 1805 -347
rect 2267 -381 2823 -347
rect 3285 -381 3841 -347
rect 4303 -381 4859 -347
rect 5321 -381 5877 -347
rect 6339 -381 6895 -347
rect 7357 -381 7913 -347
<< locali >>
rect -7929 347 -7913 381
rect -7357 347 -7341 381
rect -6911 347 -6895 381
rect -6339 347 -6323 381
rect -5893 347 -5877 381
rect -5321 347 -5305 381
rect -4875 347 -4859 381
rect -4303 347 -4287 381
rect -3857 347 -3841 381
rect -3285 347 -3269 381
rect -2839 347 -2823 381
rect -2267 347 -2251 381
rect -1821 347 -1805 381
rect -1249 347 -1233 381
rect -803 347 -787 381
rect -231 347 -215 381
rect 215 347 231 381
rect 787 347 803 381
rect 1233 347 1249 381
rect 1805 347 1821 381
rect 2251 347 2267 381
rect 2823 347 2839 381
rect 3269 347 3285 381
rect 3841 347 3857 381
rect 4287 347 4303 381
rect 4859 347 4875 381
rect 5305 347 5321 381
rect 5877 347 5893 381
rect 6323 347 6339 381
rect 6895 347 6911 381
rect 7341 347 7357 381
rect 7913 347 7929 381
rect -8161 288 -8127 304
rect -8161 -304 -8127 -288
rect -7143 288 -7109 304
rect -7143 -304 -7109 -288
rect -6125 288 -6091 304
rect -6125 -304 -6091 -288
rect -5107 288 -5073 304
rect -5107 -304 -5073 -288
rect -4089 288 -4055 304
rect -4089 -304 -4055 -288
rect -3071 288 -3037 304
rect -3071 -304 -3037 -288
rect -2053 288 -2019 304
rect -2053 -304 -2019 -288
rect -1035 288 -1001 304
rect -1035 -304 -1001 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 1001 288 1035 304
rect 1001 -304 1035 -288
rect 2019 288 2053 304
rect 2019 -304 2053 -288
rect 3037 288 3071 304
rect 3037 -304 3071 -288
rect 4055 288 4089 304
rect 4055 -304 4089 -288
rect 5073 288 5107 304
rect 5073 -304 5107 -288
rect 6091 288 6125 304
rect 6091 -304 6125 -288
rect 7109 288 7143 304
rect 7109 -304 7143 -288
rect 8127 288 8161 304
rect 8127 -304 8161 -288
rect -7929 -381 -7913 -347
rect -7357 -381 -7341 -347
rect -6911 -381 -6895 -347
rect -6339 -381 -6323 -347
rect -5893 -381 -5877 -347
rect -5321 -381 -5305 -347
rect -4875 -381 -4859 -347
rect -4303 -381 -4287 -347
rect -3857 -381 -3841 -347
rect -3285 -381 -3269 -347
rect -2839 -381 -2823 -347
rect -2267 -381 -2251 -347
rect -1821 -381 -1805 -347
rect -1249 -381 -1233 -347
rect -803 -381 -787 -347
rect -231 -381 -215 -347
rect 215 -381 231 -347
rect 787 -381 803 -347
rect 1233 -381 1249 -347
rect 1805 -381 1821 -347
rect 2251 -381 2267 -347
rect 2823 -381 2839 -347
rect 3269 -381 3285 -347
rect 3841 -381 3857 -347
rect 4287 -381 4303 -347
rect 4859 -381 4875 -347
rect 5305 -381 5321 -347
rect 5877 -381 5893 -347
rect 6323 -381 6339 -347
rect 6895 -381 6911 -347
rect 7341 -381 7357 -347
rect 7913 -381 7929 -347
<< viali >>
rect -7867 347 -7403 381
rect -6849 347 -6385 381
rect -5831 347 -5367 381
rect -4813 347 -4349 381
rect -3795 347 -3331 381
rect -2777 347 -2313 381
rect -1759 347 -1295 381
rect -741 347 -277 381
rect 277 347 741 381
rect 1295 347 1759 381
rect 2313 347 2777 381
rect 3331 347 3795 381
rect 4349 347 4813 381
rect 5367 347 5831 381
rect 6385 347 6849 381
rect 7403 347 7867 381
rect -8161 -288 -8127 288
rect -7143 -288 -7109 288
rect -6125 -288 -6091 288
rect -5107 -288 -5073 288
rect -4089 -288 -4055 288
rect -3071 -288 -3037 288
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect 3037 -288 3071 288
rect 4055 -288 4089 288
rect 5073 -288 5107 288
rect 6091 -288 6125 288
rect 7109 -288 7143 288
rect 8127 -288 8161 288
rect -7867 -381 -7403 -347
rect -6849 -381 -6385 -347
rect -5831 -381 -5367 -347
rect -4813 -381 -4349 -347
rect -3795 -381 -3331 -347
rect -2777 -381 -2313 -347
rect -1759 -381 -1295 -347
rect -741 -381 -277 -347
rect 277 -381 741 -347
rect 1295 -381 1759 -347
rect 2313 -381 2777 -347
rect 3331 -381 3795 -347
rect 4349 -381 4813 -347
rect 5367 -381 5831 -347
rect 6385 -381 6849 -347
rect 7403 -381 7867 -347
<< metal1 >>
rect -7879 381 -7391 387
rect -7879 347 -7867 381
rect -7403 347 -7391 381
rect -7879 341 -7391 347
rect -6861 381 -6373 387
rect -6861 347 -6849 381
rect -6385 347 -6373 381
rect -6861 341 -6373 347
rect -5843 381 -5355 387
rect -5843 347 -5831 381
rect -5367 347 -5355 381
rect -5843 341 -5355 347
rect -4825 381 -4337 387
rect -4825 347 -4813 381
rect -4349 347 -4337 381
rect -4825 341 -4337 347
rect -3807 381 -3319 387
rect -3807 347 -3795 381
rect -3331 347 -3319 381
rect -3807 341 -3319 347
rect -2789 381 -2301 387
rect -2789 347 -2777 381
rect -2313 347 -2301 381
rect -2789 341 -2301 347
rect -1771 381 -1283 387
rect -1771 347 -1759 381
rect -1295 347 -1283 381
rect -1771 341 -1283 347
rect -753 381 -265 387
rect -753 347 -741 381
rect -277 347 -265 381
rect -753 341 -265 347
rect 265 381 753 387
rect 265 347 277 381
rect 741 347 753 381
rect 265 341 753 347
rect 1283 381 1771 387
rect 1283 347 1295 381
rect 1759 347 1771 381
rect 1283 341 1771 347
rect 2301 381 2789 387
rect 2301 347 2313 381
rect 2777 347 2789 381
rect 2301 341 2789 347
rect 3319 381 3807 387
rect 3319 347 3331 381
rect 3795 347 3807 381
rect 3319 341 3807 347
rect 4337 381 4825 387
rect 4337 347 4349 381
rect 4813 347 4825 381
rect 4337 341 4825 347
rect 5355 381 5843 387
rect 5355 347 5367 381
rect 5831 347 5843 381
rect 5355 341 5843 347
rect 6373 381 6861 387
rect 6373 347 6385 381
rect 6849 347 6861 381
rect 6373 341 6861 347
rect 7391 381 7879 387
rect 7391 347 7403 381
rect 7867 347 7879 381
rect 7391 341 7879 347
rect -8167 288 -8121 300
rect -8167 -288 -8161 288
rect -8127 -288 -8121 288
rect -8167 -300 -8121 -288
rect -7149 288 -7103 300
rect -7149 -288 -7143 288
rect -7109 -288 -7103 288
rect -7149 -300 -7103 -288
rect -6131 288 -6085 300
rect -6131 -288 -6125 288
rect -6091 -288 -6085 288
rect -6131 -300 -6085 -288
rect -5113 288 -5067 300
rect -5113 -288 -5107 288
rect -5073 -288 -5067 288
rect -5113 -300 -5067 -288
rect -4095 288 -4049 300
rect -4095 -288 -4089 288
rect -4055 -288 -4049 288
rect -4095 -300 -4049 -288
rect -3077 288 -3031 300
rect -3077 -288 -3071 288
rect -3037 -288 -3031 288
rect -3077 -300 -3031 -288
rect -2059 288 -2013 300
rect -2059 -288 -2053 288
rect -2019 -288 -2013 288
rect -2059 -300 -2013 -288
rect -1041 288 -995 300
rect -1041 -288 -1035 288
rect -1001 -288 -995 288
rect -1041 -300 -995 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 995 288 1041 300
rect 995 -288 1001 288
rect 1035 -288 1041 288
rect 995 -300 1041 -288
rect 2013 288 2059 300
rect 2013 -288 2019 288
rect 2053 -288 2059 288
rect 2013 -300 2059 -288
rect 3031 288 3077 300
rect 3031 -288 3037 288
rect 3071 -288 3077 288
rect 3031 -300 3077 -288
rect 4049 288 4095 300
rect 4049 -288 4055 288
rect 4089 -288 4095 288
rect 4049 -300 4095 -288
rect 5067 288 5113 300
rect 5067 -288 5073 288
rect 5107 -288 5113 288
rect 5067 -300 5113 -288
rect 6085 288 6131 300
rect 6085 -288 6091 288
rect 6125 -288 6131 288
rect 6085 -300 6131 -288
rect 7103 288 7149 300
rect 7103 -288 7109 288
rect 7143 -288 7149 288
rect 7103 -300 7149 -288
rect 8121 288 8167 300
rect 8121 -288 8127 288
rect 8161 -288 8167 288
rect 8121 -300 8167 -288
rect -7879 -347 -7391 -341
rect -7879 -381 -7867 -347
rect -7403 -381 -7391 -347
rect -7879 -387 -7391 -381
rect -6861 -347 -6373 -341
rect -6861 -381 -6849 -347
rect -6385 -381 -6373 -347
rect -6861 -387 -6373 -381
rect -5843 -347 -5355 -341
rect -5843 -381 -5831 -347
rect -5367 -381 -5355 -347
rect -5843 -387 -5355 -381
rect -4825 -347 -4337 -341
rect -4825 -381 -4813 -347
rect -4349 -381 -4337 -347
rect -4825 -387 -4337 -381
rect -3807 -347 -3319 -341
rect -3807 -381 -3795 -347
rect -3331 -381 -3319 -347
rect -3807 -387 -3319 -381
rect -2789 -347 -2301 -341
rect -2789 -381 -2777 -347
rect -2313 -381 -2301 -347
rect -2789 -387 -2301 -381
rect -1771 -347 -1283 -341
rect -1771 -381 -1759 -347
rect -1295 -381 -1283 -347
rect -1771 -387 -1283 -381
rect -753 -347 -265 -341
rect -753 -381 -741 -347
rect -277 -381 -265 -347
rect -753 -387 -265 -381
rect 265 -347 753 -341
rect 265 -381 277 -347
rect 741 -381 753 -347
rect 265 -387 753 -381
rect 1283 -347 1771 -341
rect 1283 -381 1295 -347
rect 1759 -381 1771 -347
rect 1283 -387 1771 -381
rect 2301 -347 2789 -341
rect 2301 -381 2313 -347
rect 2777 -381 2789 -347
rect 2301 -387 2789 -381
rect 3319 -347 3807 -341
rect 3319 -381 3331 -347
rect 3795 -381 3807 -347
rect 3319 -387 3807 -381
rect 4337 -347 4825 -341
rect 4337 -381 4349 -347
rect 4813 -381 4825 -347
rect 4337 -387 4825 -381
rect 5355 -347 5843 -341
rect 5355 -381 5367 -347
rect 5831 -381 5843 -347
rect 5355 -387 5843 -381
rect 6373 -347 6861 -341
rect 6373 -381 6385 -347
rect 6849 -381 6861 -347
rect 6373 -387 6861 -381
rect 7391 -347 7879 -341
rect 7391 -381 7403 -347
rect 7867 -381 7879 -347
rect 7391 -387 7879 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 3 l 4.8 m 1 nf 16 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
