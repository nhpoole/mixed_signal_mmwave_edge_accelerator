magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -3361 -1660 3361 1660
<< nwell >>
rect -2101 -400 2101 400
<< pmoslvt >>
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
<< pdiff >>
rect -2065 255 -2007 300
rect -2065 221 -2053 255
rect -2019 221 -2007 255
rect -2065 187 -2007 221
rect -2065 153 -2053 187
rect -2019 153 -2007 187
rect -2065 119 -2007 153
rect -2065 85 -2053 119
rect -2019 85 -2007 119
rect -2065 51 -2007 85
rect -2065 17 -2053 51
rect -2019 17 -2007 51
rect -2065 -17 -2007 17
rect -2065 -51 -2053 -17
rect -2019 -51 -2007 -17
rect -2065 -85 -2007 -51
rect -2065 -119 -2053 -85
rect -2019 -119 -2007 -85
rect -2065 -153 -2007 -119
rect -2065 -187 -2053 -153
rect -2019 -187 -2007 -153
rect -2065 -221 -2007 -187
rect -2065 -255 -2053 -221
rect -2019 -255 -2007 -221
rect -2065 -300 -2007 -255
rect -1047 255 -989 300
rect -1047 221 -1035 255
rect -1001 221 -989 255
rect -1047 187 -989 221
rect -1047 153 -1035 187
rect -1001 153 -989 187
rect -1047 119 -989 153
rect -1047 85 -1035 119
rect -1001 85 -989 119
rect -1047 51 -989 85
rect -1047 17 -1035 51
rect -1001 17 -989 51
rect -1047 -17 -989 17
rect -1047 -51 -1035 -17
rect -1001 -51 -989 -17
rect -1047 -85 -989 -51
rect -1047 -119 -1035 -85
rect -1001 -119 -989 -85
rect -1047 -153 -989 -119
rect -1047 -187 -1035 -153
rect -1001 -187 -989 -153
rect -1047 -221 -989 -187
rect -1047 -255 -1035 -221
rect -1001 -255 -989 -221
rect -1047 -300 -989 -255
rect -29 255 29 300
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -300 29 -255
rect 989 255 1047 300
rect 989 221 1001 255
rect 1035 221 1047 255
rect 989 187 1047 221
rect 989 153 1001 187
rect 1035 153 1047 187
rect 989 119 1047 153
rect 989 85 1001 119
rect 1035 85 1047 119
rect 989 51 1047 85
rect 989 17 1001 51
rect 1035 17 1047 51
rect 989 -17 1047 17
rect 989 -51 1001 -17
rect 1035 -51 1047 -17
rect 989 -85 1047 -51
rect 989 -119 1001 -85
rect 1035 -119 1047 -85
rect 989 -153 1047 -119
rect 989 -187 1001 -153
rect 1035 -187 1047 -153
rect 989 -221 1047 -187
rect 989 -255 1001 -221
rect 1035 -255 1047 -221
rect 989 -300 1047 -255
rect 2007 255 2065 300
rect 2007 221 2019 255
rect 2053 221 2065 255
rect 2007 187 2065 221
rect 2007 153 2019 187
rect 2053 153 2065 187
rect 2007 119 2065 153
rect 2007 85 2019 119
rect 2053 85 2065 119
rect 2007 51 2065 85
rect 2007 17 2019 51
rect 2053 17 2065 51
rect 2007 -17 2065 17
rect 2007 -51 2019 -17
rect 2053 -51 2065 -17
rect 2007 -85 2065 -51
rect 2007 -119 2019 -85
rect 2053 -119 2065 -85
rect 2007 -153 2065 -119
rect 2007 -187 2019 -153
rect 2053 -187 2065 -153
rect 2007 -221 2065 -187
rect 2007 -255 2019 -221
rect 2053 -255 2065 -221
rect 2007 -300 2065 -255
<< pdiffc >>
rect -2053 221 -2019 255
rect -2053 153 -2019 187
rect -2053 85 -2019 119
rect -2053 17 -2019 51
rect -2053 -51 -2019 -17
rect -2053 -119 -2019 -85
rect -2053 -187 -2019 -153
rect -2053 -255 -2019 -221
rect -1035 221 -1001 255
rect -1035 153 -1001 187
rect -1035 85 -1001 119
rect -1035 17 -1001 51
rect -1035 -51 -1001 -17
rect -1035 -119 -1001 -85
rect -1035 -187 -1001 -153
rect -1035 -255 -1001 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 1001 221 1035 255
rect 1001 153 1035 187
rect 1001 85 1035 119
rect 1001 17 1035 51
rect 1001 -51 1035 -17
rect 1001 -119 1035 -85
rect 1001 -187 1035 -153
rect 1001 -255 1035 -221
rect 2019 221 2053 255
rect 2019 153 2053 187
rect 2019 85 2053 119
rect 2019 17 2053 51
rect 2019 -51 2053 -17
rect 2019 -119 2053 -85
rect 2019 -187 2053 -153
rect 2019 -255 2053 -221
<< poly >>
rect -1821 381 -1233 397
rect -1821 364 -1782 381
rect -2007 347 -1782 364
rect -1748 347 -1714 381
rect -1680 347 -1646 381
rect -1612 347 -1578 381
rect -1544 347 -1510 381
rect -1476 347 -1442 381
rect -1408 347 -1374 381
rect -1340 347 -1306 381
rect -1272 364 -1233 381
rect -803 381 -215 397
rect -803 364 -764 381
rect -1272 347 -1047 364
rect -2007 300 -1047 347
rect -989 347 -764 364
rect -730 347 -696 381
rect -662 347 -628 381
rect -594 347 -560 381
rect -526 347 -492 381
rect -458 347 -424 381
rect -390 347 -356 381
rect -322 347 -288 381
rect -254 364 -215 381
rect 215 381 803 397
rect 215 364 254 381
rect -254 347 -29 364
rect -989 300 -29 347
rect 29 347 254 364
rect 288 347 322 381
rect 356 347 390 381
rect 424 347 458 381
rect 492 347 526 381
rect 560 347 594 381
rect 628 347 662 381
rect 696 347 730 381
rect 764 364 803 381
rect 1233 381 1821 397
rect 1233 364 1272 381
rect 764 347 989 364
rect 29 300 989 347
rect 1047 347 1272 364
rect 1306 347 1340 381
rect 1374 347 1408 381
rect 1442 347 1476 381
rect 1510 347 1544 381
rect 1578 347 1612 381
rect 1646 347 1680 381
rect 1714 347 1748 381
rect 1782 364 1821 381
rect 1782 347 2007 364
rect 1047 300 2007 347
rect -2007 -347 -1047 -300
rect -2007 -364 -1782 -347
rect -1821 -381 -1782 -364
rect -1748 -381 -1714 -347
rect -1680 -381 -1646 -347
rect -1612 -381 -1578 -347
rect -1544 -381 -1510 -347
rect -1476 -381 -1442 -347
rect -1408 -381 -1374 -347
rect -1340 -381 -1306 -347
rect -1272 -364 -1047 -347
rect -989 -347 -29 -300
rect -989 -364 -764 -347
rect -1272 -381 -1233 -364
rect -1821 -397 -1233 -381
rect -803 -381 -764 -364
rect -730 -381 -696 -347
rect -662 -381 -628 -347
rect -594 -381 -560 -347
rect -526 -381 -492 -347
rect -458 -381 -424 -347
rect -390 -381 -356 -347
rect -322 -381 -288 -347
rect -254 -364 -29 -347
rect 29 -347 989 -300
rect 29 -364 254 -347
rect -254 -381 -215 -364
rect -803 -397 -215 -381
rect 215 -381 254 -364
rect 288 -381 322 -347
rect 356 -381 390 -347
rect 424 -381 458 -347
rect 492 -381 526 -347
rect 560 -381 594 -347
rect 628 -381 662 -347
rect 696 -381 730 -347
rect 764 -364 989 -347
rect 1047 -347 2007 -300
rect 1047 -364 1272 -347
rect 764 -381 803 -364
rect 215 -397 803 -381
rect 1233 -381 1272 -364
rect 1306 -381 1340 -347
rect 1374 -381 1408 -347
rect 1442 -381 1476 -347
rect 1510 -381 1544 -347
rect 1578 -381 1612 -347
rect 1646 -381 1680 -347
rect 1714 -381 1748 -347
rect 1782 -364 2007 -347
rect 1782 -381 1821 -364
rect 1233 -397 1821 -381
<< polycont >>
rect -1782 347 -1748 381
rect -1714 347 -1680 381
rect -1646 347 -1612 381
rect -1578 347 -1544 381
rect -1510 347 -1476 381
rect -1442 347 -1408 381
rect -1374 347 -1340 381
rect -1306 347 -1272 381
rect -764 347 -730 381
rect -696 347 -662 381
rect -628 347 -594 381
rect -560 347 -526 381
rect -492 347 -458 381
rect -424 347 -390 381
rect -356 347 -322 381
rect -288 347 -254 381
rect 254 347 288 381
rect 322 347 356 381
rect 390 347 424 381
rect 458 347 492 381
rect 526 347 560 381
rect 594 347 628 381
rect 662 347 696 381
rect 730 347 764 381
rect 1272 347 1306 381
rect 1340 347 1374 381
rect 1408 347 1442 381
rect 1476 347 1510 381
rect 1544 347 1578 381
rect 1612 347 1646 381
rect 1680 347 1714 381
rect 1748 347 1782 381
rect -1782 -381 -1748 -347
rect -1714 -381 -1680 -347
rect -1646 -381 -1612 -347
rect -1578 -381 -1544 -347
rect -1510 -381 -1476 -347
rect -1442 -381 -1408 -347
rect -1374 -381 -1340 -347
rect -1306 -381 -1272 -347
rect -764 -381 -730 -347
rect -696 -381 -662 -347
rect -628 -381 -594 -347
rect -560 -381 -526 -347
rect -492 -381 -458 -347
rect -424 -381 -390 -347
rect -356 -381 -322 -347
rect -288 -381 -254 -347
rect 254 -381 288 -347
rect 322 -381 356 -347
rect 390 -381 424 -347
rect 458 -381 492 -347
rect 526 -381 560 -347
rect 594 -381 628 -347
rect 662 -381 696 -347
rect 730 -381 764 -347
rect 1272 -381 1306 -347
rect 1340 -381 1374 -347
rect 1408 -381 1442 -347
rect 1476 -381 1510 -347
rect 1544 -381 1578 -347
rect 1612 -381 1646 -347
rect 1680 -381 1714 -347
rect 1748 -381 1782 -347
<< locali >>
rect -1821 347 -1782 381
rect -1748 347 -1724 381
rect -1680 347 -1652 381
rect -1612 347 -1580 381
rect -1544 347 -1510 381
rect -1474 347 -1442 381
rect -1402 347 -1374 381
rect -1330 347 -1306 381
rect -1272 347 -1233 381
rect -803 347 -764 381
rect -730 347 -706 381
rect -662 347 -634 381
rect -594 347 -562 381
rect -526 347 -492 381
rect -456 347 -424 381
rect -384 347 -356 381
rect -312 347 -288 381
rect -254 347 -215 381
rect 215 347 254 381
rect 288 347 312 381
rect 356 347 384 381
rect 424 347 456 381
rect 492 347 526 381
rect 562 347 594 381
rect 634 347 662 381
rect 706 347 730 381
rect 764 347 803 381
rect 1233 347 1272 381
rect 1306 347 1330 381
rect 1374 347 1402 381
rect 1442 347 1474 381
rect 1510 347 1544 381
rect 1580 347 1612 381
rect 1652 347 1680 381
rect 1724 347 1748 381
rect 1782 347 1821 381
rect -2053 269 -2019 304
rect -2053 197 -2019 221
rect -2053 125 -2019 153
rect -2053 53 -2019 85
rect -2053 -17 -2019 17
rect -2053 -85 -2019 -53
rect -2053 -153 -2019 -125
rect -2053 -221 -2019 -197
rect -2053 -304 -2019 -269
rect -1035 269 -1001 304
rect -1035 197 -1001 221
rect -1035 125 -1001 153
rect -1035 53 -1001 85
rect -1035 -17 -1001 17
rect -1035 -85 -1001 -53
rect -1035 -153 -1001 -125
rect -1035 -221 -1001 -197
rect -1035 -304 -1001 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 1001 269 1035 304
rect 1001 197 1035 221
rect 1001 125 1035 153
rect 1001 53 1035 85
rect 1001 -17 1035 17
rect 1001 -85 1035 -53
rect 1001 -153 1035 -125
rect 1001 -221 1035 -197
rect 1001 -304 1035 -269
rect 2019 269 2053 304
rect 2019 197 2053 221
rect 2019 125 2053 153
rect 2019 53 2053 85
rect 2019 -17 2053 17
rect 2019 -85 2053 -53
rect 2019 -153 2053 -125
rect 2019 -221 2053 -197
rect 2019 -304 2053 -269
rect -1821 -381 -1782 -347
rect -1748 -381 -1724 -347
rect -1680 -381 -1652 -347
rect -1612 -381 -1580 -347
rect -1544 -381 -1510 -347
rect -1474 -381 -1442 -347
rect -1402 -381 -1374 -347
rect -1330 -381 -1306 -347
rect -1272 -381 -1233 -347
rect -803 -381 -764 -347
rect -730 -381 -706 -347
rect -662 -381 -634 -347
rect -594 -381 -562 -347
rect -526 -381 -492 -347
rect -456 -381 -424 -347
rect -384 -381 -356 -347
rect -312 -381 -288 -347
rect -254 -381 -215 -347
rect 215 -381 254 -347
rect 288 -381 312 -347
rect 356 -381 384 -347
rect 424 -381 456 -347
rect 492 -381 526 -347
rect 562 -381 594 -347
rect 634 -381 662 -347
rect 706 -381 730 -347
rect 764 -381 803 -347
rect 1233 -381 1272 -347
rect 1306 -381 1330 -347
rect 1374 -381 1402 -347
rect 1442 -381 1474 -347
rect 1510 -381 1544 -347
rect 1580 -381 1612 -347
rect 1652 -381 1680 -347
rect 1724 -381 1748 -347
rect 1782 -381 1821 -347
<< viali >>
rect -1724 347 -1714 381
rect -1714 347 -1690 381
rect -1652 347 -1646 381
rect -1646 347 -1618 381
rect -1580 347 -1578 381
rect -1578 347 -1546 381
rect -1508 347 -1476 381
rect -1476 347 -1474 381
rect -1436 347 -1408 381
rect -1408 347 -1402 381
rect -1364 347 -1340 381
rect -1340 347 -1330 381
rect -706 347 -696 381
rect -696 347 -672 381
rect -634 347 -628 381
rect -628 347 -600 381
rect -562 347 -560 381
rect -560 347 -528 381
rect -490 347 -458 381
rect -458 347 -456 381
rect -418 347 -390 381
rect -390 347 -384 381
rect -346 347 -322 381
rect -322 347 -312 381
rect 312 347 322 381
rect 322 347 346 381
rect 384 347 390 381
rect 390 347 418 381
rect 456 347 458 381
rect 458 347 490 381
rect 528 347 560 381
rect 560 347 562 381
rect 600 347 628 381
rect 628 347 634 381
rect 672 347 696 381
rect 696 347 706 381
rect 1330 347 1340 381
rect 1340 347 1364 381
rect 1402 347 1408 381
rect 1408 347 1436 381
rect 1474 347 1476 381
rect 1476 347 1508 381
rect 1546 347 1578 381
rect 1578 347 1580 381
rect 1618 347 1646 381
rect 1646 347 1652 381
rect 1690 347 1714 381
rect 1714 347 1724 381
rect -2053 255 -2019 269
rect -2053 235 -2019 255
rect -2053 187 -2019 197
rect -2053 163 -2019 187
rect -2053 119 -2019 125
rect -2053 91 -2019 119
rect -2053 51 -2019 53
rect -2053 19 -2019 51
rect -2053 -51 -2019 -19
rect -2053 -53 -2019 -51
rect -2053 -119 -2019 -91
rect -2053 -125 -2019 -119
rect -2053 -187 -2019 -163
rect -2053 -197 -2019 -187
rect -2053 -255 -2019 -235
rect -2053 -269 -2019 -255
rect -1035 255 -1001 269
rect -1035 235 -1001 255
rect -1035 187 -1001 197
rect -1035 163 -1001 187
rect -1035 119 -1001 125
rect -1035 91 -1001 119
rect -1035 51 -1001 53
rect -1035 19 -1001 51
rect -1035 -51 -1001 -19
rect -1035 -53 -1001 -51
rect -1035 -119 -1001 -91
rect -1035 -125 -1001 -119
rect -1035 -187 -1001 -163
rect -1035 -197 -1001 -187
rect -1035 -255 -1001 -235
rect -1035 -269 -1001 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 1001 255 1035 269
rect 1001 235 1035 255
rect 1001 187 1035 197
rect 1001 163 1035 187
rect 1001 119 1035 125
rect 1001 91 1035 119
rect 1001 51 1035 53
rect 1001 19 1035 51
rect 1001 -51 1035 -19
rect 1001 -53 1035 -51
rect 1001 -119 1035 -91
rect 1001 -125 1035 -119
rect 1001 -187 1035 -163
rect 1001 -197 1035 -187
rect 1001 -255 1035 -235
rect 1001 -269 1035 -255
rect 2019 255 2053 269
rect 2019 235 2053 255
rect 2019 187 2053 197
rect 2019 163 2053 187
rect 2019 119 2053 125
rect 2019 91 2053 119
rect 2019 51 2053 53
rect 2019 19 2053 51
rect 2019 -51 2053 -19
rect 2019 -53 2053 -51
rect 2019 -119 2053 -91
rect 2019 -125 2053 -119
rect 2019 -187 2053 -163
rect 2019 -197 2053 -187
rect 2019 -255 2053 -235
rect 2019 -269 2053 -255
rect -1724 -381 -1714 -347
rect -1714 -381 -1690 -347
rect -1652 -381 -1646 -347
rect -1646 -381 -1618 -347
rect -1580 -381 -1578 -347
rect -1578 -381 -1546 -347
rect -1508 -381 -1476 -347
rect -1476 -381 -1474 -347
rect -1436 -381 -1408 -347
rect -1408 -381 -1402 -347
rect -1364 -381 -1340 -347
rect -1340 -381 -1330 -347
rect -706 -381 -696 -347
rect -696 -381 -672 -347
rect -634 -381 -628 -347
rect -628 -381 -600 -347
rect -562 -381 -560 -347
rect -560 -381 -528 -347
rect -490 -381 -458 -347
rect -458 -381 -456 -347
rect -418 -381 -390 -347
rect -390 -381 -384 -347
rect -346 -381 -322 -347
rect -322 -381 -312 -347
rect 312 -381 322 -347
rect 322 -381 346 -347
rect 384 -381 390 -347
rect 390 -381 418 -347
rect 456 -381 458 -347
rect 458 -381 490 -347
rect 528 -381 560 -347
rect 560 -381 562 -347
rect 600 -381 628 -347
rect 628 -381 634 -347
rect 672 -381 696 -347
rect 696 -381 706 -347
rect 1330 -381 1340 -347
rect 1340 -381 1364 -347
rect 1402 -381 1408 -347
rect 1408 -381 1436 -347
rect 1474 -381 1476 -347
rect 1476 -381 1508 -347
rect 1546 -381 1578 -347
rect 1578 -381 1580 -347
rect 1618 -381 1646 -347
rect 1646 -381 1652 -347
rect 1690 -381 1714 -347
rect 1714 -381 1724 -347
<< metal1 >>
rect -1771 381 -1283 387
rect -1771 347 -1724 381
rect -1690 347 -1652 381
rect -1618 347 -1580 381
rect -1546 347 -1508 381
rect -1474 347 -1436 381
rect -1402 347 -1364 381
rect -1330 347 -1283 381
rect -1771 341 -1283 347
rect -753 381 -265 387
rect -753 347 -706 381
rect -672 347 -634 381
rect -600 347 -562 381
rect -528 347 -490 381
rect -456 347 -418 381
rect -384 347 -346 381
rect -312 347 -265 381
rect -753 341 -265 347
rect 265 381 753 387
rect 265 347 312 381
rect 346 347 384 381
rect 418 347 456 381
rect 490 347 528 381
rect 562 347 600 381
rect 634 347 672 381
rect 706 347 753 381
rect 265 341 753 347
rect 1283 381 1771 387
rect 1283 347 1330 381
rect 1364 347 1402 381
rect 1436 347 1474 381
rect 1508 347 1546 381
rect 1580 347 1618 381
rect 1652 347 1690 381
rect 1724 347 1771 381
rect 1283 341 1771 347
rect -2059 269 -2013 300
rect -2059 235 -2053 269
rect -2019 235 -2013 269
rect -2059 197 -2013 235
rect -2059 163 -2053 197
rect -2019 163 -2013 197
rect -2059 125 -2013 163
rect -2059 91 -2053 125
rect -2019 91 -2013 125
rect -2059 53 -2013 91
rect -2059 19 -2053 53
rect -2019 19 -2013 53
rect -2059 -19 -2013 19
rect -2059 -53 -2053 -19
rect -2019 -53 -2013 -19
rect -2059 -91 -2013 -53
rect -2059 -125 -2053 -91
rect -2019 -125 -2013 -91
rect -2059 -163 -2013 -125
rect -2059 -197 -2053 -163
rect -2019 -197 -2013 -163
rect -2059 -235 -2013 -197
rect -2059 -269 -2053 -235
rect -2019 -269 -2013 -235
rect -2059 -300 -2013 -269
rect -1041 269 -995 300
rect -1041 235 -1035 269
rect -1001 235 -995 269
rect -1041 197 -995 235
rect -1041 163 -1035 197
rect -1001 163 -995 197
rect -1041 125 -995 163
rect -1041 91 -1035 125
rect -1001 91 -995 125
rect -1041 53 -995 91
rect -1041 19 -1035 53
rect -1001 19 -995 53
rect -1041 -19 -995 19
rect -1041 -53 -1035 -19
rect -1001 -53 -995 -19
rect -1041 -91 -995 -53
rect -1041 -125 -1035 -91
rect -1001 -125 -995 -91
rect -1041 -163 -995 -125
rect -1041 -197 -1035 -163
rect -1001 -197 -995 -163
rect -1041 -235 -995 -197
rect -1041 -269 -1035 -235
rect -1001 -269 -995 -235
rect -1041 -300 -995 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 995 269 1041 300
rect 995 235 1001 269
rect 1035 235 1041 269
rect 995 197 1041 235
rect 995 163 1001 197
rect 1035 163 1041 197
rect 995 125 1041 163
rect 995 91 1001 125
rect 1035 91 1041 125
rect 995 53 1041 91
rect 995 19 1001 53
rect 1035 19 1041 53
rect 995 -19 1041 19
rect 995 -53 1001 -19
rect 1035 -53 1041 -19
rect 995 -91 1041 -53
rect 995 -125 1001 -91
rect 1035 -125 1041 -91
rect 995 -163 1041 -125
rect 995 -197 1001 -163
rect 1035 -197 1041 -163
rect 995 -235 1041 -197
rect 995 -269 1001 -235
rect 1035 -269 1041 -235
rect 995 -300 1041 -269
rect 2013 269 2059 300
rect 2013 235 2019 269
rect 2053 235 2059 269
rect 2013 197 2059 235
rect 2013 163 2019 197
rect 2053 163 2059 197
rect 2013 125 2059 163
rect 2013 91 2019 125
rect 2053 91 2059 125
rect 2013 53 2059 91
rect 2013 19 2019 53
rect 2053 19 2059 53
rect 2013 -19 2059 19
rect 2013 -53 2019 -19
rect 2053 -53 2059 -19
rect 2013 -91 2059 -53
rect 2013 -125 2019 -91
rect 2053 -125 2059 -91
rect 2013 -163 2059 -125
rect 2013 -197 2019 -163
rect 2053 -197 2059 -163
rect 2013 -235 2059 -197
rect 2013 -269 2019 -235
rect 2053 -269 2059 -235
rect 2013 -300 2059 -269
rect -1771 -347 -1283 -341
rect -1771 -381 -1724 -347
rect -1690 -381 -1652 -347
rect -1618 -381 -1580 -347
rect -1546 -381 -1508 -347
rect -1474 -381 -1436 -347
rect -1402 -381 -1364 -347
rect -1330 -381 -1283 -347
rect -1771 -387 -1283 -381
rect -753 -347 -265 -341
rect -753 -381 -706 -347
rect -672 -381 -634 -347
rect -600 -381 -562 -347
rect -528 -381 -490 -347
rect -456 -381 -418 -347
rect -384 -381 -346 -347
rect -312 -381 -265 -347
rect -753 -387 -265 -381
rect 265 -347 753 -341
rect 265 -381 312 -347
rect 346 -381 384 -347
rect 418 -381 456 -347
rect 490 -381 528 -347
rect 562 -381 600 -347
rect 634 -381 672 -347
rect 706 -381 753 -347
rect 265 -387 753 -381
rect 1283 -347 1771 -341
rect 1283 -381 1330 -347
rect 1364 -381 1402 -347
rect 1436 -381 1474 -347
rect 1508 -381 1546 -347
rect 1580 -381 1618 -347
rect 1652 -381 1690 -347
rect 1724 -381 1771 -347
rect 1283 -387 1771 -381
<< end >>
