* Stimulus file.

.param vdd=1.8 vctrl=1 Wpbias=16 Wnbias=1 Wpint=6 Wnint=0.5 Wpinv=6 Wninv=0.5 Lpmos=64 Lnmos=64 Mpmos=1 Mnmos=1

vdd VDD GND 'vdd'
*vip vip GND pwl(0 'vincm' 10n 'vincm' 11n 'vincm+5m' 50n 'vincm+5m' 51n 'vincm-5m' 90n 'vincm-5m' 91n 'vincm+5m' 130n 'vincm+5m')
*vim vim GND pwl(0 'vincm' 10n 'vincm' 11n 'vincm-5m' 50n 'vincm-5m' 51n 'vincm+5m' 90n 'vincm+5m' 91n 'vincm-5m' 130n 'vincm-5m')
*vip vip GND dc 'vincm+vsig' ac 0.5 0
*vim vim GND dc 'vincm-vsig' ac 0.5 180
vctrl vctrl GND 'vctrl'
*vintest vin_test GND pulse(0 'vdd' 0.1u 0.1u 0.1u 10u 20u)

*.measure tran cs1_rise_delay
*+   TRIG v(vin)  VAL='vdd/2' FALL=1
*+   TARG v(vcs0) VAL='vdd/2' RISE=1
*.measure tran cs1_fall_delay
*+   TRIG v(vin)  VAL='vdd/2' RISE=1
*+   TARG v(vcs0) VAL='vdd/2' FALL=1
*.measure tran vout1_rise_delay
*+   TRIG v(vcs1)  VAL='vdd/2' FALL=1
*+   TARG v(vout1) VAL='vdd/2' RISE=1
*.measure tran vout1_fall_delay
*+   TRIG v(vcs1)  VAL='vdd/2' RISE=1
*+   TARG v(vout1) VAL='vdd/2' FALL=1

.ic v(vin)=0
*.options savecurrents
.save vin x7.qint1 x7.qbint1 x7.q1 x7.qb1 x7.qint2 x7.qbint2
+   x8.qint1 x8.qbint1 x8.q1 x8.qb1 x8.qint2 x8.qbint2
+   x9.qint1 x9.qbint1 x9.q1 x9.qb1 x9.qint2 x9.qbint2

.tran 0.01u 10m

.control
let ctrl = 1.2
while ctrl < 1.3
    set ctrl = $&ctrl
    alter vctrl dc ctrl
    save vin vin2 vin_buf vdff1 vdff2 vdff3 vdff4 vdff5 vdff6 vdff7 vout
    +   x7.qint1 x7.qbint1 x7.q1 x7.qb1 x7.qint2 x7.qbint2
    +   x8.qint1 x8.qbint1 x8.q1 x8.qb1 x8.qint2 x8.qbint2
    +   x9.qint1 x9.qbint1 x9.q1 x9.qb1 x9.qint2 x9.qbint2
    run
    write cs_ring_osc_div_tran_{$ctrl}.raw vin vin2 vin_buf vdff1 vdff2 vdff3 vdff4 vdff5 vdff6 vdff7 vout
    +   x7.qint1 x7.qbint1 x7.q1 x7.qb1 x7.qint2 x7.qbint2
    +   x8.qint1 x8.qbint1 x8.q1 x8.qb1 x8.qint2 x8.qbint2
    +   x9.qint1 x9.qbint1 x9.q1 x9.qb1 x9.qint2 x9.qbint2
    let ctrl = ctrl + 0.1
end
quit
.endc
