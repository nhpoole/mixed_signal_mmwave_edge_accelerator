magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1296 -1277 3068 2731
<< nwell >>
rect -36 679 1808 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 1772 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1566 1130 1600 1397
rect 1670 1322 1704 1397
rect 64 674 98 740
rect 814 724 848 1096
rect 814 690 865 724
rect 814 318 848 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1566 17 1600 218
rect 1670 17 1704 92
rect 0 -17 1772 17
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m14_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m14_w2_000_sli_dli_da_p_0
timestamp 1626486988
transform 1 0 54 0 1 963
box -59 -56 1613 454
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m14_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m14_w2_000_sli_dli_da_p_0
timestamp 1626486988
transform 1 0 54 0 1 51
box -26 -26 1580 456
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1626486988
transform 1 0 48 0 1 674
box 0 0 66 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1626486988
transform 1 0 1662 0 1 51
box -26 -26 76 108
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1626486988
transform 1 0 1662 0 1 1281
box -59 -43 109 125
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 848 707 848 707 4 Z
rlabel locali s 886 0 886 0 4 gnd
rlabel locali s 886 1414 886 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1772 1414
<< end >>
