magic
tech sky130A
magscale 1 2
timestamp 1625985445
<< nwell >>
rect -11247 15506 -9306 16346
rect -7803 15507 -7200 15828
<< viali >>
rect -7288 15458 -7240 15506
rect -7184 15462 -7136 15510
<< metal1 >>
rect -4458 30288 -4398 30294
rect -4458 16436 -4398 30228
rect -11018 16376 -9518 16436
rect -8284 16376 -7916 16436
rect -7856 16376 -7850 16436
rect -4464 16376 -4458 16436
rect -4398 16376 -4392 16436
rect -7540 15742 -7332 15838
rect -7490 15506 -7228 15512
rect -7490 15458 -7288 15506
rect -7240 15458 -7228 15506
rect -7490 15452 -7228 15458
rect -7196 15510 -7030 15516
rect -7196 15462 -7184 15510
rect -7136 15462 -7030 15510
rect -7196 15456 -7030 15462
rect -7528 15198 -7326 15294
rect -9694 14740 -9688 14760
rect -11068 14680 -9566 14740
rect -8452 14680 -1320 14740
rect 664 1564 1066 1624
<< via1 >>
rect -4458 30228 -4398 30288
rect -7916 16376 -7856 16436
rect -4458 16376 -4398 16436
<< metal2 >>
rect -4458 30288 -4398 30297
rect -4464 30228 -4458 30288
rect -4398 30228 -4392 30288
rect -4458 30219 -4398 30228
rect -7916 16436 -7856 16442
rect -4458 16436 -4398 16442
rect -7856 16376 -4458 16436
rect -7916 16370 -7856 16376
rect -4458 16370 -4398 16376
rect -13297 15502 -13288 15562
rect -13228 15502 -11530 15562
rect -9675 15502 -9666 15562
rect -9606 15502 -8926 15562
rect -12495 15353 -12486 15413
rect -12426 15353 -11732 15413
rect -9859 15353 -9850 15413
rect -9790 15353 -9164 15413
rect -10082 14806 -7716 14866
rect -13105 14576 -13015 14580
rect -9874 14576 -9774 14585
rect -13110 14571 -9874 14576
rect -13110 14481 -13105 14571
rect -13015 14481 -9874 14571
rect -13110 14476 -9874 14481
rect -9774 14476 -9766 14576
rect -13105 14472 -13015 14476
rect -9874 14467 -9774 14476
rect -13499 14354 -13409 14358
rect -9686 14354 -9586 14363
rect -13504 14349 -9686 14354
rect -13504 14259 -13499 14349
rect -13409 14259 -9686 14349
rect -13504 14254 -9686 14259
rect -13499 14250 -13409 14254
rect -9686 14245 -9586 14254
rect -11022 11009 -10932 11014
rect -11026 10929 -11017 11009
rect -10937 10929 -10928 11009
rect -6664 11001 -6578 11006
rect -11022 10869 -10932 10929
rect -6668 10925 -6659 11001
rect -6583 10925 -6574 11001
rect -6664 10871 -6578 10925
rect -11022 10779 -8595 10869
rect -6664 10785 -4371 10871
rect -8685 10703 -8595 10779
rect -8685 10604 -8595 10613
rect -4457 10689 -4371 10785
rect -4457 10594 -4371 10603
rect -1851 6458 -1842 6518
rect -1782 6458 480 6518
rect -1566 5556 -1506 5565
rect -1506 5496 2058 5556
rect -1566 5487 -1506 5496
rect -10744 3789 -10642 3794
rect -6568 3791 -6474 3796
rect -10748 3697 -10739 3789
rect -10647 3697 -10638 3789
rect -6572 3707 -6563 3791
rect -6479 3707 -6470 3791
rect -10744 3649 -10642 3697
rect -10744 3547 -8631 3649
rect -8733 3485 -8631 3547
rect -6568 3639 -6474 3707
rect -6568 3545 -4455 3639
rect -8733 3374 -8631 3383
rect -4549 3473 -4455 3545
rect -4549 3370 -4455 3379
<< via2 >>
rect -4458 30228 -4398 30288
rect -13288 15502 -13228 15562
rect -9666 15502 -9606 15562
rect -12486 15353 -12426 15413
rect -9850 15353 -9790 15413
rect -13105 14481 -13015 14571
rect -9874 14476 -9774 14576
rect -13499 14259 -13409 14349
rect -9686 14254 -9586 14354
rect -11017 10929 -10937 11009
rect -6659 10925 -6583 11001
rect -8685 10613 -8595 10703
rect -4457 10603 -4371 10689
rect -1842 6458 -1782 6518
rect -1566 5496 -1506 5556
rect -10739 3697 -10647 3789
rect -6563 3707 -6479 3791
rect -8733 3383 -8631 3485
rect -4549 3379 -4455 3473
<< metal3 >>
rect -4486 30293 -4350 30322
rect -4486 30229 -4463 30293
rect -4393 30229 -4350 30293
rect -4486 30228 -4458 30229
rect -4398 30228 -4350 30229
rect -4486 30192 -4350 30228
rect -13310 15562 -13210 15584
rect -13310 15502 -13288 15562
rect -13228 15502 -13210 15562
rect -13504 14349 -13404 14354
rect -13504 14259 -13499 14349
rect -13409 14259 -13404 14349
rect -13504 3497 -13404 14259
rect -13310 5903 -13210 15502
rect -9686 15562 -9586 15580
rect -9686 15502 -9666 15562
rect -9606 15502 -9586 15562
rect -12510 15413 -12410 15434
rect -12510 15353 -12486 15413
rect -12426 15353 -12410 15413
rect -12510 14688 -12410 15353
rect -12510 14582 -12410 14588
rect -9874 15413 -9774 15436
rect -9874 15353 -9850 15413
rect -9790 15353 -9774 15413
rect -9874 14581 -9774 15353
rect -9879 14576 -9769 14581
rect -13110 14571 -13010 14576
rect -13110 14481 -13105 14571
rect -13015 14481 -13010 14571
rect -13110 10725 -13010 14481
rect -9879 14476 -9874 14576
rect -9774 14476 -9769 14576
rect -9879 14471 -9769 14476
rect -9686 14359 -9586 15502
rect 10952 14470 11052 14476
rect -1600 14370 10952 14470
rect -9691 14354 -9581 14359
rect -9691 14254 -9686 14354
rect -9586 14254 -9581 14354
rect -9691 14249 -9581 14254
rect -11124 14114 -10954 14120
rect -12012 14010 -11124 14012
rect -12572 13944 -11124 14010
rect -8772 14118 -8612 14124
rect -10954 13958 -8772 14012
rect -6398 14122 -6256 14128
rect -8612 13980 -6398 14012
rect -4024 14106 -3862 14112
rect -6256 13980 -4024 14012
rect -8612 13958 -4024 13980
rect -10954 13944 -4024 13958
rect -3862 14010 -2864 14012
rect -3862 13944 -2610 14010
rect -12572 13408 -2610 13944
rect -12572 11918 -11971 13408
rect -10026 13056 -7214 13156
rect -10026 12694 -9896 13056
rect -7314 12716 -7214 13056
rect -10026 12562 -9926 12694
rect -12700 11820 -12694 11918
rect -12596 11820 -11971 11918
rect -13115 10627 -13109 10725
rect -13011 10627 -13005 10725
rect -13110 10626 -13010 10627
rect -12572 9826 -11971 11820
rect -3213 11908 -2610 13408
rect -1858 12903 -1758 12904
rect -1863 12805 -1857 12903
rect -1759 12805 -1753 12903
rect -3213 11786 -2562 11908
rect -2440 11786 -2434 11908
rect -11022 11009 -10932 11046
rect -9332 11021 -9232 11294
rect -5192 11029 -5092 11278
rect -11022 10929 -11017 11009
rect -10937 10929 -10932 11009
rect -11022 10924 -10932 10929
rect -9337 10923 -9331 11021
rect -9233 10923 -9227 11021
rect -6664 11001 -6578 11028
rect -6664 10925 -6659 11001
rect -6583 10925 -6578 11001
rect -5197 10931 -5191 11029
rect -5093 10931 -5087 11029
rect -5192 10930 -5092 10931
rect -9332 10922 -9232 10923
rect -6664 10920 -6578 10925
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10881 -7570 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -7570 10881
rect -8102 10782 -7570 10783
rect -3901 10880 -3803 10885
rect -3400 10880 -3300 10886
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -3902 10879 -3400 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3400 10879
rect -3902 10780 -3400 10781
rect -3901 10775 -3803 10780
rect -3400 10774 -3300 10780
rect -10156 10725 -10056 10726
rect -5956 10725 -5856 10726
rect -10161 10627 -10155 10725
rect -10057 10627 -10051 10725
rect -8690 10703 -8590 10708
rect -10156 10588 -10056 10627
rect -8690 10613 -8685 10703
rect -8595 10613 -8590 10703
rect -5961 10627 -5955 10725
rect -5857 10627 -5851 10725
rect -4462 10689 -4366 10694
rect -8690 10608 -8590 10613
rect -10156 10476 -10002 10588
rect -12678 9708 -12672 9826
rect -12554 9708 -11971 9826
rect -13100 8615 -13000 8616
rect -13105 8517 -13099 8615
rect -13001 8517 -12995 8615
rect -13315 5805 -13309 5903
rect -13211 5805 -13205 5903
rect -13310 5804 -13210 5805
rect -13509 3399 -13503 3497
rect -13405 3399 -13399 3497
rect -13504 3398 -13404 3399
rect -13100 1627 -13000 8517
rect -12572 8256 -11971 9708
rect -10102 8616 -10002 10476
rect -8685 10421 -8595 10608
rect -5956 10476 -5856 10627
rect -4462 10603 -4457 10689
rect -4371 10603 -4366 10689
rect -4462 10598 -4366 10603
rect -4457 10357 -4371 10598
rect -3213 9850 -2610 11786
rect -3213 9742 -2534 9850
rect -2426 9742 -2420 9850
rect -7192 8616 -7092 9154
rect -10510 8516 -10504 8616
rect -10404 8516 -7092 8616
rect -3213 8256 -2610 9742
rect -12572 7654 -2610 8256
rect -12572 7652 -2956 7654
rect -11068 7570 -10886 7652
rect -11068 7402 -11061 7570
rect -10893 7402 -10886 7570
rect -8768 7570 -8586 7652
rect -8768 7402 -8761 7570
rect -8593 7402 -8586 7570
rect -6468 7570 -6286 7652
rect -6468 7402 -6461 7570
rect -6293 7402 -6286 7570
rect -4048 7570 -3866 7652
rect -4048 7402 -4041 7570
rect -3873 7402 -3866 7570
rect -11062 7401 -10892 7402
rect -8762 7401 -8592 7402
rect -6462 7401 -6292 7402
rect -4042 7401 -3872 7402
rect -11062 6884 -10892 6890
rect -11950 6778 -11062 6782
rect -12509 6714 -11062 6778
rect -8762 6884 -8592 6890
rect -10892 6714 -8762 6782
rect -6462 6884 -6292 6890
rect -8592 6714 -6462 6782
rect -4042 6884 -3872 6890
rect -6292 6714 -4042 6782
rect -3872 6778 -2802 6782
rect -3872 6714 -2548 6778
rect -12509 6178 -2548 6714
rect -12509 4688 -11909 6178
rect -11530 5804 -11524 5904
rect -11424 5804 -7198 5904
rect -10006 5428 -9906 5804
rect -7298 5478 -7198 5804
rect -12638 4590 -12632 4688
rect -12534 4590 -11909 4688
rect -12509 2596 -11909 4590
rect -3151 4678 -2548 6178
rect -1858 6518 -1758 12805
rect -1600 8863 -1500 14370
rect 10952 14364 11052 14370
rect -1605 8765 -1599 8863
rect -1501 8765 -1495 8863
rect -1600 8764 -1500 8765
rect -1858 6458 -1842 6518
rect -1782 6458 -1758 6518
rect -1858 5665 -1758 6458
rect -1863 5567 -1857 5665
rect -1759 5567 -1753 5665
rect -1858 5566 -1758 5567
rect -1586 5556 -1486 5594
rect -1586 5496 -1566 5556
rect -1506 5496 -1486 5556
rect -3151 4556 -2500 4678
rect -2378 4556 -2372 4678
rect -10744 3789 -10642 3844
rect -9304 3797 -9204 4022
rect -10744 3697 -10739 3789
rect -10647 3697 -10642 3789
rect -9309 3699 -9303 3797
rect -9205 3699 -9199 3797
rect -6568 3791 -6474 3830
rect -5084 3801 -4984 4060
rect -6568 3707 -6563 3791
rect -6479 3707 -6474 3791
rect -6568 3702 -6474 3707
rect -5089 3703 -5083 3801
rect -4985 3703 -4979 3801
rect -5084 3702 -4984 3703
rect -9304 3698 -9204 3699
rect -10744 3692 -10642 3697
rect -8085 3644 -7987 3649
rect -7554 3644 -7454 3650
rect -3845 3644 -3747 3649
rect -3344 3644 -3244 3650
rect -8086 3643 -7554 3644
rect -8086 3545 -8085 3643
rect -7987 3545 -7554 3643
rect -8086 3544 -7554 3545
rect -3846 3643 -3344 3644
rect -3846 3545 -3845 3643
rect -3747 3545 -3344 3643
rect -3846 3544 -3344 3545
rect -8085 3539 -7987 3544
rect -7554 3538 -7454 3544
rect -3845 3539 -3747 3544
rect -3344 3538 -3244 3544
rect -5940 3501 -5840 3502
rect -10180 3497 -10080 3498
rect -10185 3399 -10179 3497
rect -10081 3399 -10075 3497
rect -8738 3485 -8626 3490
rect -10180 3350 -10080 3399
rect -8738 3383 -8733 3485
rect -8631 3383 -8626 3485
rect -8738 3378 -8626 3383
rect -10180 3238 -10026 3350
rect -12616 2478 -12610 2596
rect -12492 2478 -11909 2596
rect -13103 1529 -13097 1627
rect -12999 1529 -12993 1627
rect -13100 1528 -13000 1529
rect -12509 1028 -11909 2478
rect -10126 1378 -10026 3238
rect -8733 3109 -8631 3378
rect -7176 3254 -7174 3446
rect -5945 3403 -5939 3501
rect -5841 3403 -5835 3501
rect -4554 3473 -4450 3478
rect -5940 3238 -5840 3403
rect -4554 3379 -4549 3473
rect -4455 3379 -4450 3473
rect -4554 3374 -4450 3379
rect -4549 3065 -4455 3374
rect -3151 2620 -2548 4556
rect -3151 2512 -2472 2620
rect -2364 2512 -2358 2620
rect -7176 1378 -7076 1916
rect -10126 1278 -7076 1378
rect -3151 1028 -2548 2512
rect -1586 1625 -1486 5496
rect -1591 1527 -1585 1625
rect -1487 1527 -1481 1625
rect -1586 1526 -1486 1527
rect -12509 484 -2548 1028
rect -12509 422 -11094 484
rect -10918 422 -8682 484
rect -11094 302 -10918 308
rect -8506 422 -6362 484
rect -8682 302 -8506 308
rect -6186 422 -3962 484
rect -6362 302 -6186 308
rect -3786 424 -2548 484
rect -3786 422 -3061 424
rect -3962 302 -3786 308
<< via3 >>
rect -4463 30288 -4393 30293
rect -4463 30229 -4458 30288
rect -4458 30229 -4398 30288
rect -4398 30229 -4393 30288
rect -12510 14588 -12410 14688
rect 10952 14370 11052 14470
rect -11124 13944 -10954 14114
rect -8772 13958 -8612 14118
rect -6398 13980 -6256 14122
rect -4024 13944 -3862 14106
rect -12694 11820 -12596 11918
rect -13109 10627 -13011 10725
rect -1857 12805 -1759 12903
rect -2562 11786 -2440 11908
rect -9331 10923 -9233 11021
rect -5191 10931 -5093 11029
rect -8101 10783 -8003 10881
rect -7570 10782 -7470 10882
rect -3901 10781 -3803 10879
rect -3400 10780 -3300 10880
rect -10155 10627 -10057 10725
rect -5955 10627 -5857 10725
rect -12672 9708 -12554 9826
rect -13099 8517 -13001 8615
rect -13309 5805 -13211 5903
rect -13503 3399 -13405 3497
rect -2534 9742 -2426 9850
rect -10504 8516 -10404 8616
rect -11061 7402 -10893 7570
rect -8761 7402 -8593 7570
rect -6461 7402 -6293 7570
rect -4041 7402 -3873 7570
rect -11062 6714 -10892 6884
rect -8762 6714 -8592 6884
rect -6462 6714 -6292 6884
rect -4042 6714 -3872 6884
rect -11524 5804 -11424 5904
rect -12632 4590 -12534 4688
rect -1599 8765 -1501 8863
rect -1857 5567 -1759 5665
rect -2500 4556 -2378 4678
rect -9303 3699 -9205 3797
rect -5083 3703 -4985 3801
rect -8085 3545 -7987 3643
rect -7554 3544 -7454 3644
rect -3845 3545 -3747 3643
rect -3344 3544 -3244 3644
rect -10179 3399 -10081 3497
rect -12610 2478 -12492 2596
rect -13097 1529 -12999 1627
rect -5939 3403 -5841 3501
rect -2472 2512 -2364 2620
rect -1585 1527 -1487 1625
rect -11094 308 -10918 484
rect -8682 308 -8506 484
rect -6362 308 -6186 484
rect -3962 308 -3786 484
<< metal4 >>
rect -4928 30293 -3252 30940
rect -4928 30229 -4463 30293
rect -4393 30229 -3252 30293
rect -4928 30140 -3252 30229
rect -12511 14688 -12409 14689
rect -12511 14588 -12510 14688
rect -12410 14588 -12409 14688
rect -12511 14587 -12409 14588
rect -12510 13220 -12410 14587
rect 10952 14471 11052 15140
rect 10951 14470 11053 14471
rect 10951 14370 10952 14470
rect 11052 14370 11053 14470
rect 10951 14369 11053 14370
rect -6399 14122 -6255 14123
rect -8773 14118 -8611 14119
rect -11125 14114 -10953 14115
rect -11125 13944 -11124 14114
rect -10954 13944 -10953 14114
rect -8773 13958 -8772 14118
rect -8612 13958 -8611 14118
rect -6399 13980 -6398 14122
rect -6256 13980 -6255 14122
rect -6399 13979 -6255 13980
rect -4025 14106 -3861 14107
rect -8773 13957 -8611 13958
rect -11125 13943 -10953 13944
rect -11124 13605 -10954 13943
rect -8772 13654 -8612 13957
rect -6398 13705 -6256 13979
rect -4025 13944 -4024 14106
rect -3862 13944 -3861 14106
rect -4025 13943 -3861 13944
rect -4024 13667 -3862 13943
rect -12510 13120 -10034 13220
rect -10134 12904 -10034 13120
rect -10134 12903 -1758 12904
rect -10134 12805 -1857 12903
rect -1759 12805 -1758 12903
rect -10134 12804 -1758 12805
rect -10134 12450 -10034 12804
rect -12695 11918 -12595 11919
rect -12695 11820 -12694 11918
rect -12596 11820 -12243 11918
rect -12695 11819 -12595 11820
rect -8246 11784 -7706 11884
rect -9332 11021 -9232 11022
rect -9332 10923 -9331 11021
rect -9233 10923 -9232 11021
rect -9332 10726 -9232 10923
rect -13110 10725 -9232 10726
rect -13110 10627 -13109 10725
rect -13011 10627 -10155 10725
rect -10057 10627 -9232 10725
rect -13110 10626 -9232 10627
rect -8102 10881 -8002 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -8002 10881
rect -8102 10382 -8002 10783
rect -12673 9826 -12553 9827
rect -12673 9708 -12672 9826
rect -12554 9708 -12205 9826
rect -12673 9707 -12553 9708
rect -10152 8864 -10052 9244
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12450 -5834 12804
rect -4046 11784 -3506 11884
rect -5192 11029 -5092 11030
rect -5192 10931 -5191 11029
rect -5093 10931 -5092 11029
rect -7571 10882 -7469 10883
rect -7571 10782 -7570 10882
rect -7470 10782 -7469 10882
rect -7571 10781 -7469 10782
rect -5192 10726 -5092 10931
rect -5956 10725 -5092 10726
rect -5956 10627 -5955 10725
rect -5857 10627 -5092 10725
rect -5956 10626 -5092 10627
rect -3902 10879 -3802 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3802 10879
rect -3902 10382 -3802 10781
rect -5952 8864 -5852 9244
rect -3606 8864 -3506 11784
rect -3400 10881 -3300 12804
rect -2563 11908 -2439 11909
rect -2879 11786 -2562 11908
rect -2440 11786 -2439 11908
rect -2563 11785 -2439 11786
rect -3401 10880 -3299 10881
rect -3401 10780 -3400 10880
rect -3300 10780 -3299 10880
rect -3401 10779 -3299 10780
rect -2535 9850 -2425 9851
rect -2922 9742 -2534 9850
rect -2426 9742 -2425 9850
rect -2535 9741 -2425 9742
rect -10152 8863 -1500 8864
rect -10152 8765 -1599 8863
rect -1501 8765 -1500 8863
rect -10152 8764 -1500 8765
rect -10505 8616 -10403 8617
rect -13100 8615 -10504 8616
rect -13100 8517 -13099 8615
rect -13001 8517 -10504 8615
rect -13100 8516 -10504 8517
rect -10404 8516 -10403 8616
rect -10505 8515 -10403 8516
rect -11062 7570 -10892 7927
rect -11062 7402 -11061 7570
rect -10893 7402 -10892 7570
rect -11062 6885 -10892 7402
rect -8762 7570 -8592 7927
rect -8762 7402 -8761 7570
rect -8593 7402 -8592 7570
rect -8762 6885 -8592 7402
rect -6462 7570 -6292 7927
rect -6462 7402 -6461 7570
rect -6293 7402 -6292 7570
rect -6462 6885 -6292 7402
rect -4042 7570 -3872 7927
rect -4042 7402 -4041 7570
rect -3873 7402 -3872 7570
rect -4042 6885 -3872 7402
rect -11063 6884 -10891 6885
rect -11063 6714 -11062 6884
rect -10892 6714 -10891 6884
rect -11063 6713 -10891 6714
rect -8763 6884 -8591 6885
rect -8763 6714 -8762 6884
rect -8592 6714 -8591 6884
rect -8763 6713 -8591 6714
rect -6463 6884 -6291 6885
rect -6463 6714 -6462 6884
rect -6292 6714 -6291 6884
rect -6463 6713 -6291 6714
rect -4043 6884 -3871 6885
rect -4043 6714 -4042 6884
rect -3872 6714 -3871 6884
rect -4043 6713 -3871 6714
rect -11062 6375 -10892 6713
rect -8762 6375 -8592 6713
rect -6462 6375 -6292 6713
rect -4042 6375 -3872 6713
rect -11525 5904 -11423 5905
rect -13310 5903 -11524 5904
rect -13310 5805 -13309 5903
rect -13211 5805 -11524 5903
rect -13310 5804 -11524 5805
rect -11424 5804 -11423 5904
rect -11525 5803 -11423 5804
rect -10158 5665 -1758 5666
rect -10158 5567 -1857 5665
rect -1759 5567 -1758 5665
rect -10158 5566 -1758 5567
rect -10158 5212 -10058 5566
rect -12633 4688 -12533 4689
rect -12633 4590 -12632 4688
rect -12534 4590 -12181 4688
rect -12633 4589 -12533 4590
rect -8230 4546 -7690 4646
rect -9304 3797 -9204 3798
rect -9304 3699 -9303 3797
rect -9205 3699 -9204 3797
rect -9304 3498 -9204 3699
rect -13504 3497 -9204 3498
rect -13504 3399 -13503 3497
rect -13405 3399 -10179 3497
rect -10081 3399 -9204 3497
rect -13504 3398 -9204 3399
rect -8086 3643 -7986 3644
rect -8086 3545 -8085 3643
rect -7987 3545 -7986 3643
rect -8086 3144 -7986 3545
rect -12611 2596 -12491 2597
rect -12611 2478 -12610 2596
rect -12492 2478 -12143 2596
rect -12611 2477 -12491 2478
rect -10176 1628 -10076 2006
rect -13098 1627 -9512 1628
rect -13098 1529 -13097 1627
rect -12999 1626 -9512 1627
rect -7790 1626 -7690 4546
rect -7554 3645 -7454 5566
rect -5918 5212 -5818 5566
rect -3990 4546 -3450 4646
rect -5084 3801 -4984 3802
rect -5084 3703 -5083 3801
rect -4985 3703 -4984 3801
rect -7555 3644 -7453 3645
rect -7555 3544 -7554 3644
rect -7454 3544 -7453 3644
rect -7555 3543 -7453 3544
rect -5084 3502 -4984 3703
rect -5940 3501 -4984 3502
rect -5940 3403 -5939 3501
rect -5841 3403 -4984 3501
rect -5940 3402 -4984 3403
rect -3846 3643 -3746 3644
rect -3846 3545 -3845 3643
rect -3747 3545 -3746 3643
rect -3846 3144 -3746 3545
rect -5936 1626 -5836 2006
rect -3550 1626 -3450 4546
rect -3344 3645 -3244 5566
rect -2501 4678 -2377 4679
rect -2817 4556 -2500 4678
rect -2378 4556 -2377 4678
rect -2501 4555 -2377 4556
rect -3345 3644 -3243 3645
rect -3345 3544 -3344 3644
rect -3244 3544 -3243 3644
rect -3345 3543 -3243 3544
rect -2473 2620 -2363 2621
rect -2860 2512 -2472 2620
rect -2364 2512 -2363 2620
rect -2473 2511 -2363 2512
rect -12999 1625 -1486 1626
rect -12999 1529 -1585 1625
rect -13098 1528 -1585 1529
rect -10176 1527 -1585 1528
rect -1487 1527 -1486 1625
rect -10176 1526 -1486 1527
rect -11094 485 -10918 750
rect -8682 485 -8506 750
rect -6362 485 -6186 750
rect -3962 485 -3786 750
rect -11095 484 -10917 485
rect -11095 308 -11094 484
rect -10918 308 -10917 484
rect -11095 307 -10917 308
rect -8683 484 -8505 485
rect -8683 308 -8682 484
rect -8506 308 -8505 484
rect -8683 307 -8505 308
rect -6363 484 -6185 485
rect -6363 308 -6362 484
rect -6186 308 -6185 484
rect -6363 307 -6185 308
rect -3963 484 -3785 485
rect -3963 308 -3962 484
rect -3786 308 -3785 484
rect -3963 307 -3785 308
rect -11094 140 -10918 307
rect -8682 140 -8506 307
rect -6362 140 -6186 307
rect -3962 140 -3786 307
rect -13514 -660 -1808 140
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_4
timestamp 1624477805
transform 1 0 -12158 0 1 2542
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_7
timestamp 1624477805
transform 1 0 -8632 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_4
timestamp 1624477805
transform -1 0 -11077 0 1 724
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_0
timestamp 1624477805
transform 1 0 -8594 0 1 724
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_6
timestamp 1624477805
transform 1 0 -10672 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_9
timestamp 1624477805
transform 1 0 -6432 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_7
timestamp 1624477805
transform 1 0 -3823 0 1 726
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_3
timestamp 1624477805
transform -1 0 -6306 0 1 726
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_8
timestamp 1624477805
transform 1 0 -4392 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_7
timestamp 1624477805
transform -1 0 -2902 0 1 2544
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_5
timestamp 1624477805
transform 1 0 -12158 0 1 4646
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_0
timestamp 1624477805
transform -1 0 -11139 0 1 7954
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_4
timestamp 1624477805
transform 1 0 -8632 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_5
timestamp 1624477805
transform -1 0 -11077 0 1 6480
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_1
timestamp 1624477805
transform 1 0 -8594 0 1 6480
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_5
timestamp 1624477805
transform 1 0 -10672 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_4
timestamp 1624477805
transform 1 0 -8656 0 1 7954
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_10
timestamp 1624477805
transform 1 0 -6432 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_2
timestamp 1624477805
transform -1 0 -6306 0 1 6482
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_6
timestamp 1624477805
transform 1 0 -3823 0 1 6482
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_11
timestamp 1624477805
transform 1 0 -4392 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_5
timestamp 1624477805
transform -1 0 -6368 0 1 7956
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_1
timestamp 1624477805
transform 1 0 -3885 0 1 7956
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_6
timestamp 1624477805
transform -1 0 -2902 0 1 4648
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_2
timestamp 1624477805
transform 1 0 -12220 0 1 9772
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_3
timestamp 1624477805
transform 1 0 -12220 0 1 11876
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_0
timestamp 1624477805
transform 1 0 -10734 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_1
timestamp 1624477805
transform 1 0 -8694 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_12
timestamp 1624477805
transform 1 0 -10734 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_14
timestamp 1624477805
transform 1 0 -8694 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_2
timestamp 1624477805
transform 1 0 -6494 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_3
timestamp 1624477805
transform 1 0 -4454 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_13
timestamp 1624477805
transform 1 0 -6494 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_15
timestamp 1624477805
transform 1 0 -4454 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_0
timestamp 1624477805
transform -1 0 -2964 0 1 9774
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_1
timestamp 1624477805
transform -1 0 -2964 0 1 11878
box -350 -900 244 900
use txgate  txgate_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/txgate
timestamp 1625985445
transform 1 0 -86501 0 1 -42680
box 74185 57360 76542 59116
use txgate  txgate_1
timestamp 1625985445
transform 1 0 -83901 0 1 -42680
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_2
timestamp 1624477805
transform -1 0 -11139 0 1 13710
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_6
timestamp 1624477805
transform 1 0 -8656 0 1 13710
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_3
timestamp 1624477805
transform 1 0 -3885 0 1 13712
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_7
timestamp 1624477805
transform -1 0 -6368 0 1 13712
box -950 -300 818 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 -7070 0 1 15246
box -38 -48 314 592
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624477805
transform 1 0 10912 0 1 26540
box -15168 -27258 25000 4400
<< labels >>
flabel metal4 -5616 -342 -5562 -296 1 FreeSans 480 0 0 0 VSS
flabel metal4 -9816 8794 -9798 8822 1 FreeSans 480 0 0 0 vse
flabel metal4 -9746 12834 -9732 12846 1 FreeSans 480 0 0 0 vip
flabel metal1 704 1582 716 1600 1 FreeSans 480 0 0 0 ibiasn
flabel metal4 -4738 30526 -4712 30558 1 FreeSans 480 0 0 0 VDD
flabel metal1 -7056 15480 -7054 15484 1 FreeSans 480 0 0 0 rst_n
flabel metal1 -7332 15474 -7328 15480 1 FreeSans 480 0 0 0 rst
flabel metal3 -9542 5852 -9520 5872 1 FreeSans 480 0 0 0 vdiffp
flabel metal4 -9702 5600 -9680 5618 1 FreeSans 480 0 0 0 vip
flabel metal4 -9786 1568 -9770 1582 1 FreeSans 480 0 0 0 vim
flabel metal3 -9812 1318 -9800 1332 1 FreeSans 480 0 0 0 vdiffm
flabel metal3 -9752 13102 -9732 13118 1 FreeSans 480 0 0 0 vocm
flabel metal3 -9862 8562 -9854 8578 1 FreeSans 480 0 0 0 vim
<< end >>
