magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2812 -7339 24942 6535
<< nwell >>
rect 9590 3318 13304 5174
rect 9590 -5978 13120 -4122
<< metal1 >>
rect 4664 -2764 4724 -2754
rect 4664 -2816 4668 -2764
rect 4720 -2816 4724 -2764
rect 4664 -3466 4724 -2816
rect 5690 -2766 5762 -2762
rect 5690 -2818 5700 -2766
rect 5752 -2818 5762 -2766
rect 5690 -2822 5762 -2818
rect 6602 -2822 6792 -2762
rect 5052 -3716 5112 -3398
rect 5308 -3716 5368 -3402
rect 5696 -3410 5756 -2822
rect 6080 -3716 6140 -3400
rect 6342 -3716 6402 -3404
rect 6732 -3414 6792 -2822
rect 16854 -3712 16914 -3430
rect 16848 -3716 16920 -3712
rect 5046 -3720 5118 -3716
rect 5046 -3772 5056 -3720
rect 5108 -3772 5118 -3720
rect 5046 -3776 5118 -3772
rect 5302 -3720 5374 -3716
rect 5302 -3772 5312 -3720
rect 5364 -3772 5374 -3720
rect 5302 -3776 5374 -3772
rect 6074 -3720 6146 -3716
rect 6074 -3772 6084 -3720
rect 6136 -3772 6146 -3720
rect 6074 -3776 6146 -3772
rect 6336 -3720 6408 -3716
rect 6336 -3772 6346 -3720
rect 6398 -3772 6408 -3720
rect 16848 -3768 16858 -3716
rect 16910 -3768 16920 -3716
rect 16848 -3772 16920 -3768
rect 6336 -3776 6408 -3772
<< via1 >>
rect 4668 -2816 4720 -2764
rect 5700 -2818 5752 -2766
rect 5056 -3772 5108 -3720
rect 5312 -3772 5364 -3720
rect 6084 -3772 6136 -3720
rect 6346 -3772 6398 -3720
rect 16858 -3768 16910 -3716
<< metal2 >>
rect 16973 3262 17051 3264
rect 16973 3206 16984 3262
rect 17040 3206 17051 3262
rect 16973 3204 17051 3206
rect 16982 3128 17042 3204
rect 4659 2986 4737 2988
rect 4659 2930 4670 2986
rect 4726 2930 4737 2986
rect 4659 2928 4737 2930
rect 11488 2871 11588 2876
rect 11484 2854 11592 2871
rect 11484 2798 11510 2854
rect 11566 2798 11592 2854
rect 11484 2781 11592 2798
rect 16459 2854 17164 2856
rect 16459 2798 16470 2854
rect 16526 2798 17164 2854
rect 16459 2796 17164 2798
rect 4998 2686 5184 2746
rect 9642 2740 9702 2749
rect 9578 2738 9702 2740
rect 9578 2682 9644 2738
rect 9700 2682 9702 2738
rect 9578 2680 9702 2682
rect 9642 2671 9702 2680
rect 1489 2008 1796 2010
rect 1489 1952 1500 2008
rect 1556 1952 1796 2008
rect 4732 1956 5170 2016
rect 1489 1950 1796 1952
rect 6792 1050 6954 1110
rect 6772 -1914 6930 -1854
rect 4268 -2764 4928 -2760
rect 4268 -2816 4668 -2764
rect 4720 -2816 4928 -2764
rect 4268 -2820 4928 -2816
rect 5696 -2766 5756 -2756
rect 5696 -2818 5700 -2766
rect 5752 -2818 5756 -2766
rect 4268 -2916 4328 -2820
rect 5696 -2828 5756 -2818
rect 4259 -2918 4337 -2916
rect 4259 -2974 4270 -2918
rect 4326 -2974 4337 -2918
rect 4259 -2976 4337 -2974
rect 11488 -3464 11588 2781
rect 17734 2744 18213 2746
rect 17734 2688 18146 2744
rect 18202 2688 18213 2744
rect 17734 2686 18213 2688
rect 18156 1956 18980 2016
rect 11691 1894 11809 1916
rect 11691 1838 11722 1894
rect 11778 1838 11809 1894
rect 11691 1816 11809 1838
rect 11700 -2625 11800 1816
rect 18920 1684 18980 1956
rect 18911 1682 18989 1684
rect 18911 1626 18922 1682
rect 18978 1626 18989 1682
rect 18911 1624 18989 1626
rect 18536 1050 18740 1110
rect 18578 -1914 18742 -1854
rect 16979 -2404 17057 -2402
rect 16979 -2460 16990 -2404
rect 17046 -2460 17057 -2404
rect 16979 -2462 17057 -2460
rect 16988 -2522 17048 -2462
rect 16898 -2582 17048 -2522
rect 11696 -2642 11804 -2625
rect 11696 -2698 11722 -2642
rect 11778 -2698 11804 -2642
rect 11696 -2715 11804 -2698
rect 11700 -2720 11800 -2715
rect 16070 -2820 16720 -2760
rect 9286 -3486 9707 -3484
rect 5045 -3492 5304 -3490
rect 5045 -3548 5056 -3492
rect 5112 -3548 5304 -3492
rect 9286 -3542 9640 -3486
rect 9696 -3542 9707 -3486
rect 9286 -3544 9707 -3542
rect 11479 -3486 11597 -3464
rect 16070 -3480 16130 -2820
rect 11479 -3542 11510 -3486
rect 11566 -3542 11597 -3486
rect 16061 -3482 16139 -3480
rect 16061 -3538 16072 -3482
rect 16128 -3538 16139 -3482
rect 16061 -3540 16139 -3538
rect 21084 -3486 21509 -3484
rect 5045 -3550 5304 -3548
rect 11479 -3564 11597 -3542
rect 21084 -3542 21442 -3486
rect 21498 -3542 21509 -3486
rect 21084 -3544 21509 -3542
rect 5052 -3716 5112 -3710
rect 5308 -3716 5368 -3710
rect 6080 -3716 6140 -3710
rect 6342 -3716 6402 -3710
rect 16854 -3712 16914 -3706
rect 16845 -3714 16923 -3712
rect 5052 -3720 5492 -3716
rect 5052 -3772 5056 -3720
rect 5108 -3772 5312 -3720
rect 5364 -3772 5492 -3720
rect 5052 -3776 5492 -3772
rect 5980 -3718 6411 -3716
rect 5980 -3720 6344 -3718
rect 5980 -3772 6084 -3720
rect 6136 -3772 6344 -3720
rect 5980 -3774 6344 -3772
rect 6400 -3774 6411 -3718
rect 16845 -3770 16856 -3714
rect 16912 -3770 16923 -3714
rect 16845 -3772 16923 -3770
rect 5980 -3776 6411 -3774
rect 5052 -3782 5112 -3776
rect 5308 -3782 5368 -3776
rect 6080 -3782 6140 -3776
rect 6342 -3782 6402 -3776
rect 16854 -3778 16914 -3772
<< via2 >>
rect 16984 3206 17040 3262
rect 4670 2930 4726 2986
rect 11510 2798 11566 2854
rect 16470 2798 16526 2854
rect 9644 2682 9700 2738
rect 1500 1952 1556 2008
rect 4270 -2974 4326 -2918
rect 18146 2688 18202 2744
rect 11722 1838 11778 1894
rect 18922 1626 18978 1682
rect 16990 -2460 17046 -2404
rect 11722 -2698 11778 -2642
rect 5056 -3548 5112 -3492
rect 9640 -3542 9696 -3486
rect 11510 -3542 11566 -3486
rect 16072 -3538 16128 -3482
rect 21442 -3542 21498 -3486
rect 6344 -3720 6400 -3718
rect 6344 -3772 6346 -3720
rect 6346 -3772 6398 -3720
rect 6398 -3772 6400 -3720
rect 6344 -3774 6400 -3772
rect 16856 -3716 16912 -3714
rect 16856 -3768 16858 -3716
rect 16858 -3768 16910 -3716
rect 16910 -3768 16912 -3716
rect 16856 -3770 16912 -3768
<< metal3 >>
rect 9620 3262 17070 3284
rect 9620 3206 16984 3262
rect 17040 3206 17070 3262
rect 9620 3184 17070 3206
rect -592 2986 4752 3008
rect -592 2930 4670 2986
rect 4726 2930 4752 2986
rect -592 2908 4752 2930
rect -592 -3466 -492 2908
rect 9620 2738 9720 3184
rect 11488 2854 16550 2876
rect 11488 2798 11510 2854
rect 11566 2798 16470 2854
rect 16526 2798 16550 2854
rect 11488 2776 16550 2798
rect 9620 2682 9644 2738
rect 9700 2682 9720 2738
rect 9620 2660 9720 2682
rect 18128 2744 23682 2764
rect 18128 2688 18146 2744
rect 18202 2688 23682 2744
rect 18128 2664 23682 2688
rect -330 2008 1580 2030
rect -330 1952 1500 2008
rect 1556 1952 1580 2008
rect -330 1930 1580 1952
rect -330 -2450 -230 1930
rect 11695 1916 11805 1921
rect 7896 1894 16354 1916
rect 7896 1838 11722 1894
rect 11778 1838 16354 1894
rect 7896 1816 16354 1838
rect 11695 1811 11805 1816
rect 18890 1682 23412 1706
rect 18890 1626 18922 1682
rect 18978 1626 23412 1682
rect 18890 1606 23412 1626
rect 23312 -2384 23412 1606
rect 16958 -2404 23412 -2384
rect -330 -2550 3908 -2450
rect 16958 -2460 16990 -2404
rect 17046 -2460 23412 -2404
rect 16958 -2484 23412 -2460
rect 3808 -2896 3908 -2550
rect 7972 -2642 16034 -2620
rect 7972 -2698 11722 -2642
rect 11778 -2698 16034 -2642
rect 7972 -2720 16034 -2698
rect 3808 -2918 4358 -2896
rect 3808 -2974 4270 -2918
rect 4326 -2974 4358 -2918
rect 3808 -2996 4358 -2974
rect 11483 -3464 11593 -3459
rect -592 -3492 5138 -3466
rect -592 -3548 5056 -3492
rect 5112 -3548 5138 -3492
rect -592 -3566 5138 -3548
rect 9614 -3482 16158 -3464
rect 23582 -3466 23682 2664
rect 9614 -3486 16072 -3482
rect 9614 -3542 9640 -3486
rect 9696 -3542 11510 -3486
rect 11566 -3538 16072 -3486
rect 16128 -3538 16158 -3482
rect 11566 -3542 16158 -3538
rect 9614 -3564 16158 -3542
rect 21422 -3486 23682 -3466
rect 21422 -3542 21442 -3486
rect 21498 -3542 23682 -3486
rect 11483 -3569 11593 -3564
rect 21422 -3566 23682 -3542
rect 6324 -3714 16934 -3696
rect 6324 -3718 16856 -3714
rect 6324 -3774 6344 -3718
rect 6400 -3770 16856 -3718
rect 16912 -3770 16934 -3714
rect 6400 -3774 16934 -3770
rect 6324 -3796 16934 -3774
<< metal4 >>
rect -1528 5094 1572 5216
rect -1528 4538 -1406 5094
rect -850 4538 1572 5094
rect -1528 4416 1572 4538
rect 9840 4416 12720 5216
rect 11292 -180 12036 434
rect -12 -624 23288 -180
rect 11292 -1242 12036 -624
rect -1528 -5344 1572 -5220
rect -1528 -5900 -1406 -5344
rect -850 -5900 1572 -5344
rect -1528 -6020 1572 -5900
rect 9904 -6020 12650 -5220
<< via4 >>
rect -1406 4538 -850 5094
rect -1406 -5900 -850 -5344
<< metal5 >>
rect -1552 5094 -704 5240
rect -1552 4538 -1406 5094
rect -850 4538 -704 5094
rect -1552 4392 -704 4538
rect -1528 -5344 -728 4392
rect -1528 -5900 -1406 -5344
rect -850 -5900 -728 -5344
rect -1528 -6022 -728 -5900
use gm_c_stage  gm_c_stage_3
timestamp 1626486988
transform 1 0 12188 0 1 2736
box -400 -3100 11100 2480
use gm_c_stage  gm_c_stage_2
timestamp 1626486988
transform 1 0 12188 0 -1 -3540
box -400 -3100 11100 2480
use gm_c_stage  gm_c_stage_1
timestamp 1626486988
transform 1 0 388 0 -1 -3540
box -400 -3100 11100 2480
use gm_c_stage  gm_c_stage_0
timestamp 1626486988
transform 1 0 388 0 1 2736
box -400 -3100 11100 2480
<< labels >>
flabel metal2 s 4746 1978 4762 1992 1 FreeSans 600 0 0 0 vip
flabel metal2 s 5012 2710 5020 2724 1 FreeSans 600 0 0 0 vim
flabel metal3 s 11604 1874 11614 1882 1 FreeSans 600 0 0 0 vocm
flabel metal4 s 11516 5188 11546 5206 1 FreeSans 600 0 0 0 VDD
flabel metal4 s 11416 -406 11440 -390 1 FreeSans 600 0 0 0 VSS
flabel metal3 s 23620 1100 23640 1116 1 FreeSans 600 0 0 0 vfiltm
flabel metal3 s 23360 1060 23382 1076 1 FreeSans 600 0 0 0 vfiltp
flabel metal3 s -562 1138 -542 1158 1 FreeSans 600 0 0 0 vintp
flabel metal3 s -290 1124 -268 1144 1 FreeSans 600 0 0 0 vintm
flabel metal2 s 6858 1072 6874 1080 1 FreeSans 600 0 0 0 ibiasn1
flabel metal2 s 6844 -1890 6870 -1878 1 FreeSans 600 0 0 0 ibiasn2
flabel metal2 s 18656 -1896 18670 -1880 1 FreeSans 600 0 0 0 ibiasn3
flabel metal2 s 18640 1074 18656 1084 1 FreeSans 600 0 0 0 ibiasn4
<< end >>
