magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2110 -2060 2109 2060
<< metal3 >>
rect -850 627 849 800
rect -850 563 765 627
rect 829 563 849 627
rect -850 547 849 563
rect -850 483 765 547
rect 829 483 849 547
rect -850 467 849 483
rect -850 403 765 467
rect 829 403 849 467
rect -850 387 849 403
rect -850 323 765 387
rect 829 323 849 387
rect -850 307 849 323
rect -850 243 765 307
rect 829 243 849 307
rect -850 227 849 243
rect -850 163 765 227
rect 829 163 849 227
rect -850 147 849 163
rect -850 83 765 147
rect 829 83 849 147
rect -850 67 849 83
rect -850 3 765 67
rect 829 3 849 67
rect -850 -13 849 3
rect -850 -77 765 -13
rect 829 -77 849 -13
rect -850 -93 849 -77
rect -850 -157 765 -93
rect 829 -157 849 -93
rect -850 -173 849 -157
rect -850 -237 765 -173
rect 829 -237 849 -173
rect -850 -253 849 -237
rect -850 -317 765 -253
rect 829 -317 849 -253
rect -850 -333 849 -317
rect -850 -397 765 -333
rect 829 -397 849 -333
rect -850 -413 849 -397
rect -850 -477 765 -413
rect 829 -477 849 -413
rect -850 -493 849 -477
rect -850 -557 765 -493
rect 829 -557 849 -493
rect -850 -573 849 -557
rect -850 -637 765 -573
rect 829 -637 849 -573
rect -850 -800 849 -637
<< via3 >>
rect 765 563 829 627
rect 765 483 829 547
rect 765 403 829 467
rect 765 323 829 387
rect 765 243 829 307
rect 765 163 829 227
rect 765 83 829 147
rect 765 3 829 67
rect 765 -77 829 -13
rect 765 -157 829 -93
rect 765 -237 829 -173
rect 765 -317 829 -253
rect 765 -397 829 -333
rect 765 -477 829 -413
rect 765 -557 829 -493
rect 765 -637 829 -573
<< mimcap >>
rect -750 632 650 700
rect -750 -632 -682 632
rect 582 -632 650 632
rect -750 -700 650 -632
<< mimcapcontact >>
rect -682 -632 582 632
<< metal4 >>
rect -711 632 611 661
rect -711 -632 -682 632
rect 582 -632 611 632
rect -711 -661 611 -632
rect 749 627 845 662
rect 749 563 765 627
rect 829 563 845 627
rect 749 547 845 563
rect 749 483 765 547
rect 829 483 845 547
rect 749 467 845 483
rect 749 403 765 467
rect 829 403 845 467
rect 749 387 845 403
rect 749 323 765 387
rect 829 323 845 387
rect 749 307 845 323
rect 749 243 765 307
rect 829 243 845 307
rect 749 227 845 243
rect 749 163 765 227
rect 829 163 845 227
rect 749 147 845 163
rect 749 83 765 147
rect 829 83 845 147
rect 749 67 845 83
rect 749 3 765 67
rect 829 3 845 67
rect 749 -13 845 3
rect 749 -77 765 -13
rect 829 -77 845 -13
rect 749 -93 845 -77
rect 749 -157 765 -93
rect 829 -157 845 -93
rect 749 -173 845 -157
rect 749 -237 765 -173
rect 829 -237 845 -173
rect 749 -253 845 -237
rect 749 -317 765 -253
rect 829 -317 845 -253
rect 749 -333 845 -317
rect 749 -397 765 -333
rect 829 -397 845 -333
rect 749 -413 845 -397
rect 749 -477 765 -413
rect 829 -477 845 -413
rect 749 -493 845 -477
rect 749 -557 765 -493
rect 829 -557 845 -493
rect 749 -573 845 -557
rect 749 -637 765 -573
rect 829 -637 845 -573
rect 749 -662 845 -637
<< properties >>
string FIXED_BBOX -850 -800 750 800
<< end >>
