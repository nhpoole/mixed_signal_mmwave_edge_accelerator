magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1155 -300 1155 300
<< nwell >>
rect -1155 -300 1155 300
<< pmos >>
rect -1061 -200 -901 200
rect -843 -200 -683 200
rect -625 -200 -465 200
rect -407 -200 -247 200
rect -189 -200 -29 200
rect 29 -200 189 200
rect 247 -200 407 200
rect 465 -200 625 200
rect 683 -200 843 200
rect 901 -200 1061 200
<< pdiff >>
rect -1119 188 -1061 200
rect -1119 -188 -1107 188
rect -1073 -188 -1061 188
rect -1119 -200 -1061 -188
rect -901 188 -843 200
rect -901 -188 -889 188
rect -855 -188 -843 188
rect -901 -200 -843 -188
rect -683 188 -625 200
rect -683 -188 -671 188
rect -637 -188 -625 188
rect -683 -200 -625 -188
rect -465 188 -407 200
rect -465 -188 -453 188
rect -419 -188 -407 188
rect -465 -200 -407 -188
rect -247 188 -189 200
rect -247 -188 -235 188
rect -201 -188 -189 188
rect -247 -200 -189 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 189 188 247 200
rect 189 -188 201 188
rect 235 -188 247 188
rect 189 -200 247 -188
rect 407 188 465 200
rect 407 -188 419 188
rect 453 -188 465 188
rect 407 -200 465 -188
rect 625 188 683 200
rect 625 -188 637 188
rect 671 -188 683 188
rect 625 -200 683 -188
rect 843 188 901 200
rect 843 -188 855 188
rect 889 -188 901 188
rect 843 -200 901 -188
rect 1061 188 1119 200
rect 1061 -188 1073 188
rect 1107 -188 1119 188
rect 1061 -200 1119 -188
<< pdiffc >>
rect -1107 -188 -1073 188
rect -889 -188 -855 188
rect -671 -188 -637 188
rect -453 -188 -419 188
rect -235 -188 -201 188
rect -17 -188 17 188
rect 201 -188 235 188
rect 419 -188 453 188
rect 637 -188 671 188
rect 855 -188 889 188
rect 1073 -188 1107 188
<< poly >>
rect -1035 281 -927 297
rect -1035 264 -1019 281
rect -1061 247 -1019 264
rect -943 264 -927 281
rect -817 281 -709 297
rect -817 264 -801 281
rect -943 247 -901 264
rect -1061 200 -901 247
rect -843 247 -801 264
rect -725 264 -709 281
rect -599 281 -491 297
rect -599 264 -583 281
rect -725 247 -683 264
rect -843 200 -683 247
rect -625 247 -583 264
rect -507 264 -491 281
rect -381 281 -273 297
rect -381 264 -365 281
rect -507 247 -465 264
rect -625 200 -465 247
rect -407 247 -365 264
rect -289 264 -273 281
rect -163 281 -55 297
rect -163 264 -147 281
rect -289 247 -247 264
rect -407 200 -247 247
rect -189 247 -147 264
rect -71 264 -55 281
rect 55 281 163 297
rect 55 264 71 281
rect -71 247 -29 264
rect -189 200 -29 247
rect 29 247 71 264
rect 147 264 163 281
rect 273 281 381 297
rect 273 264 289 281
rect 147 247 189 264
rect 29 200 189 247
rect 247 247 289 264
rect 365 264 381 281
rect 491 281 599 297
rect 491 264 507 281
rect 365 247 407 264
rect 247 200 407 247
rect 465 247 507 264
rect 583 264 599 281
rect 709 281 817 297
rect 709 264 725 281
rect 583 247 625 264
rect 465 200 625 247
rect 683 247 725 264
rect 801 264 817 281
rect 927 281 1035 297
rect 927 264 943 281
rect 801 247 843 264
rect 683 200 843 247
rect 901 247 943 264
rect 1019 264 1035 281
rect 1019 247 1061 264
rect 901 200 1061 247
rect -1061 -247 -901 -200
rect -1061 -264 -1019 -247
rect -1035 -281 -1019 -264
rect -943 -264 -901 -247
rect -843 -247 -683 -200
rect -843 -264 -801 -247
rect -943 -281 -927 -264
rect -1035 -297 -927 -281
rect -817 -281 -801 -264
rect -725 -264 -683 -247
rect -625 -247 -465 -200
rect -625 -264 -583 -247
rect -725 -281 -709 -264
rect -817 -297 -709 -281
rect -599 -281 -583 -264
rect -507 -264 -465 -247
rect -407 -247 -247 -200
rect -407 -264 -365 -247
rect -507 -281 -491 -264
rect -599 -297 -491 -281
rect -381 -281 -365 -264
rect -289 -264 -247 -247
rect -189 -247 -29 -200
rect -189 -264 -147 -247
rect -289 -281 -273 -264
rect -381 -297 -273 -281
rect -163 -281 -147 -264
rect -71 -264 -29 -247
rect 29 -247 189 -200
rect 29 -264 71 -247
rect -71 -281 -55 -264
rect -163 -297 -55 -281
rect 55 -281 71 -264
rect 147 -264 189 -247
rect 247 -247 407 -200
rect 247 -264 289 -247
rect 147 -281 163 -264
rect 55 -297 163 -281
rect 273 -281 289 -264
rect 365 -264 407 -247
rect 465 -247 625 -200
rect 465 -264 507 -247
rect 365 -281 381 -264
rect 273 -297 381 -281
rect 491 -281 507 -264
rect 583 -264 625 -247
rect 683 -247 843 -200
rect 683 -264 725 -247
rect 583 -281 599 -264
rect 491 -297 599 -281
rect 709 -281 725 -264
rect 801 -264 843 -247
rect 901 -247 1061 -200
rect 901 -264 943 -247
rect 801 -281 817 -264
rect 709 -297 817 -281
rect 927 -281 943 -264
rect 1019 -264 1061 -247
rect 1019 -281 1035 -264
rect 927 -297 1035 -281
<< polycont >>
rect -1019 247 -943 281
rect -801 247 -725 281
rect -583 247 -507 281
rect -365 247 -289 281
rect -147 247 -71 281
rect 71 247 147 281
rect 289 247 365 281
rect 507 247 583 281
rect 725 247 801 281
rect 943 247 1019 281
rect -1019 -281 -943 -247
rect -801 -281 -725 -247
rect -583 -281 -507 -247
rect -365 -281 -289 -247
rect -147 -281 -71 -247
rect 71 -281 147 -247
rect 289 -281 365 -247
rect 507 -281 583 -247
rect 725 -281 801 -247
rect 943 -281 1019 -247
<< locali >>
rect -1035 247 -1019 281
rect -943 247 -927 281
rect -817 247 -801 281
rect -725 247 -709 281
rect -599 247 -583 281
rect -507 247 -491 281
rect -381 247 -365 281
rect -289 247 -273 281
rect -163 247 -147 281
rect -71 247 -55 281
rect 55 247 71 281
rect 147 247 163 281
rect 273 247 289 281
rect 365 247 381 281
rect 491 247 507 281
rect 583 247 599 281
rect 709 247 725 281
rect 801 247 817 281
rect 927 247 943 281
rect 1019 247 1035 281
rect -1107 188 -1073 204
rect -1107 -204 -1073 -188
rect -889 188 -855 204
rect -889 -204 -855 -188
rect -671 188 -637 204
rect -671 -204 -637 -188
rect -453 188 -419 204
rect -453 -204 -419 -188
rect -235 188 -201 204
rect -235 -204 -201 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 201 188 235 204
rect 201 -204 235 -188
rect 419 188 453 204
rect 419 -204 453 -188
rect 637 188 671 204
rect 637 -204 671 -188
rect 855 188 889 204
rect 855 -204 889 -188
rect 1073 188 1107 204
rect 1073 -204 1107 -188
rect -1035 -281 -1019 -247
rect -943 -281 -927 -247
rect -817 -281 -801 -247
rect -725 -281 -709 -247
rect -599 -281 -583 -247
rect -507 -281 -491 -247
rect -381 -281 -365 -247
rect -289 -281 -273 -247
rect -163 -281 -147 -247
rect -71 -281 -55 -247
rect 55 -281 71 -247
rect 147 -281 163 -247
rect 273 -281 289 -247
rect 365 -281 381 -247
rect 491 -281 507 -247
rect 583 -281 599 -247
rect 709 -281 725 -247
rect 801 -281 817 -247
rect 927 -281 943 -247
rect 1019 -281 1035 -247
<< viali >>
rect -1013 247 -949 281
rect -795 247 -731 281
rect -577 247 -513 281
rect -359 247 -295 281
rect -141 247 -77 281
rect 77 247 141 281
rect 295 247 359 281
rect 513 247 577 281
rect 731 247 795 281
rect 949 247 1013 281
rect -1107 -188 -1073 188
rect -889 -188 -855 188
rect -671 -188 -637 188
rect -453 -188 -419 188
rect -235 -188 -201 188
rect -17 -188 17 188
rect 201 -188 235 188
rect 419 -188 453 188
rect 637 -188 671 188
rect 855 -188 889 188
rect 1073 -188 1107 188
rect -1013 -281 -949 -247
rect -795 -281 -731 -247
rect -577 -281 -513 -247
rect -359 -281 -295 -247
rect -141 -281 -77 -247
rect 77 -281 141 -247
rect 295 -281 359 -247
rect 513 -281 577 -247
rect 731 -281 795 -247
rect 949 -281 1013 -247
<< metal1 >>
rect -1025 281 -937 287
rect -1025 247 -1013 281
rect -949 247 -937 281
rect -1025 241 -937 247
rect -807 281 -719 287
rect -807 247 -795 281
rect -731 247 -719 281
rect -807 241 -719 247
rect -589 281 -501 287
rect -589 247 -577 281
rect -513 247 -501 281
rect -589 241 -501 247
rect -371 281 -283 287
rect -371 247 -359 281
rect -295 247 -283 281
rect -371 241 -283 247
rect -153 281 -65 287
rect -153 247 -141 281
rect -77 247 -65 281
rect -153 241 -65 247
rect 65 281 153 287
rect 65 247 77 281
rect 141 247 153 281
rect 65 241 153 247
rect 283 281 371 287
rect 283 247 295 281
rect 359 247 371 281
rect 283 241 371 247
rect 501 281 589 287
rect 501 247 513 281
rect 577 247 589 281
rect 501 241 589 247
rect 719 281 807 287
rect 719 247 731 281
rect 795 247 807 281
rect 719 241 807 247
rect 937 281 1025 287
rect 937 247 949 281
rect 1013 247 1025 281
rect 937 241 1025 247
rect -1113 188 -1067 200
rect -1113 -188 -1107 188
rect -1073 -188 -1067 188
rect -1113 -200 -1067 -188
rect -895 188 -849 200
rect -895 -188 -889 188
rect -855 -188 -849 188
rect -895 -200 -849 -188
rect -677 188 -631 200
rect -677 -188 -671 188
rect -637 -188 -631 188
rect -677 -200 -631 -188
rect -459 188 -413 200
rect -459 -188 -453 188
rect -419 -188 -413 188
rect -459 -200 -413 -188
rect -241 188 -195 200
rect -241 -188 -235 188
rect -201 -188 -195 188
rect -241 -200 -195 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 195 188 241 200
rect 195 -188 201 188
rect 235 -188 241 188
rect 195 -200 241 -188
rect 413 188 459 200
rect 413 -188 419 188
rect 453 -188 459 188
rect 413 -200 459 -188
rect 631 188 677 200
rect 631 -188 637 188
rect 671 -188 677 188
rect 631 -200 677 -188
rect 849 188 895 200
rect 849 -188 855 188
rect 889 -188 895 188
rect 849 -200 895 -188
rect 1067 188 1113 200
rect 1067 -188 1073 188
rect 1107 -188 1113 188
rect 1067 -200 1113 -188
rect -1025 -247 -937 -241
rect -1025 -281 -1013 -247
rect -949 -281 -937 -247
rect -1025 -287 -937 -281
rect -807 -247 -719 -241
rect -807 -281 -795 -247
rect -731 -281 -719 -247
rect -807 -287 -719 -281
rect -589 -247 -501 -241
rect -589 -281 -577 -247
rect -513 -281 -501 -247
rect -589 -287 -501 -281
rect -371 -247 -283 -241
rect -371 -281 -359 -247
rect -295 -281 -283 -247
rect -371 -287 -283 -281
rect -153 -247 -65 -241
rect -153 -281 -141 -247
rect -77 -281 -65 -247
rect -153 -287 -65 -281
rect 65 -247 153 -241
rect 65 -281 77 -247
rect 141 -281 153 -247
rect 65 -287 153 -281
rect 283 -247 371 -241
rect 283 -281 295 -247
rect 359 -281 371 -247
rect 283 -287 371 -281
rect 501 -247 589 -241
rect 501 -281 513 -247
rect 577 -281 589 -247
rect 501 -287 589 -281
rect 719 -247 807 -241
rect 719 -281 731 -247
rect 795 -281 807 -247
rect 719 -287 807 -281
rect 937 -247 1025 -241
rect 937 -281 949 -247
rect 1013 -281 1025 -247
rect 937 -287 1025 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 2 l 0.8 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
