magic
tech sky130A
magscale 1 2
timestamp 1620511006
<< nwell >>
rect -7700 -400 7700 400
<< pmos >>
rect -7606 -300 -6646 300
rect -6588 -300 -5628 300
rect -5570 -300 -4610 300
rect -4552 -300 -3592 300
rect -3534 -300 -2574 300
rect -2516 -300 -1556 300
rect -1498 -300 -538 300
rect -480 -300 480 300
rect 538 -300 1498 300
rect 1556 -300 2516 300
rect 2574 -300 3534 300
rect 3592 -300 4552 300
rect 4610 -300 5570 300
rect 5628 -300 6588 300
rect 6646 -300 7606 300
<< pdiff >>
rect -7664 288 -7606 300
rect -7664 -288 -7652 288
rect -7618 -288 -7606 288
rect -7664 -300 -7606 -288
rect -6646 288 -6588 300
rect -6646 -288 -6634 288
rect -6600 -288 -6588 288
rect -6646 -300 -6588 -288
rect -5628 288 -5570 300
rect -5628 -288 -5616 288
rect -5582 -288 -5570 288
rect -5628 -300 -5570 -288
rect -4610 288 -4552 300
rect -4610 -288 -4598 288
rect -4564 -288 -4552 288
rect -4610 -300 -4552 -288
rect -3592 288 -3534 300
rect -3592 -288 -3580 288
rect -3546 -288 -3534 288
rect -3592 -300 -3534 -288
rect -2574 288 -2516 300
rect -2574 -288 -2562 288
rect -2528 -288 -2516 288
rect -2574 -300 -2516 -288
rect -1556 288 -1498 300
rect -1556 -288 -1544 288
rect -1510 -288 -1498 288
rect -1556 -300 -1498 -288
rect -538 288 -480 300
rect -538 -288 -526 288
rect -492 -288 -480 288
rect -538 -300 -480 -288
rect 480 288 538 300
rect 480 -288 492 288
rect 526 -288 538 288
rect 480 -300 538 -288
rect 1498 288 1556 300
rect 1498 -288 1510 288
rect 1544 -288 1556 288
rect 1498 -300 1556 -288
rect 2516 288 2574 300
rect 2516 -288 2528 288
rect 2562 -288 2574 288
rect 2516 -300 2574 -288
rect 3534 288 3592 300
rect 3534 -288 3546 288
rect 3580 -288 3592 288
rect 3534 -300 3592 -288
rect 4552 288 4610 300
rect 4552 -288 4564 288
rect 4598 -288 4610 288
rect 4552 -300 4610 -288
rect 5570 288 5628 300
rect 5570 -288 5582 288
rect 5616 -288 5628 288
rect 5570 -300 5628 -288
rect 6588 288 6646 300
rect 6588 -288 6600 288
rect 6634 -288 6646 288
rect 6588 -300 6646 -288
rect 7606 288 7664 300
rect 7606 -288 7618 288
rect 7652 -288 7664 288
rect 7606 -300 7664 -288
<< pdiffc >>
rect -7652 -288 -7618 288
rect -6634 -288 -6600 288
rect -5616 -288 -5582 288
rect -4598 -288 -4564 288
rect -3580 -288 -3546 288
rect -2562 -288 -2528 288
rect -1544 -288 -1510 288
rect -526 -288 -492 288
rect 492 -288 526 288
rect 1510 -288 1544 288
rect 2528 -288 2562 288
rect 3546 -288 3580 288
rect 4564 -288 4598 288
rect 5582 -288 5616 288
rect 6600 -288 6634 288
rect 7618 -288 7652 288
<< poly >>
rect -7420 381 -6832 397
rect -7420 364 -7404 381
rect -7606 347 -7404 364
rect -6848 364 -6832 381
rect -6402 381 -5814 397
rect -6402 364 -6386 381
rect -6848 347 -6646 364
rect -7606 300 -6646 347
rect -6588 347 -6386 364
rect -5830 364 -5814 381
rect -5384 381 -4796 397
rect -5384 364 -5368 381
rect -5830 347 -5628 364
rect -6588 300 -5628 347
rect -5570 347 -5368 364
rect -4812 364 -4796 381
rect -4366 381 -3778 397
rect -4366 364 -4350 381
rect -4812 347 -4610 364
rect -5570 300 -4610 347
rect -4552 347 -4350 364
rect -3794 364 -3778 381
rect -3348 381 -2760 397
rect -3348 364 -3332 381
rect -3794 347 -3592 364
rect -4552 300 -3592 347
rect -3534 347 -3332 364
rect -2776 364 -2760 381
rect -2330 381 -1742 397
rect -2330 364 -2314 381
rect -2776 347 -2574 364
rect -3534 300 -2574 347
rect -2516 347 -2314 364
rect -1758 364 -1742 381
rect -1312 381 -724 397
rect -1312 364 -1296 381
rect -1758 347 -1556 364
rect -2516 300 -1556 347
rect -1498 347 -1296 364
rect -740 364 -724 381
rect -294 381 294 397
rect -294 364 -278 381
rect -740 347 -538 364
rect -1498 300 -538 347
rect -480 347 -278 364
rect 278 364 294 381
rect 724 381 1312 397
rect 724 364 740 381
rect 278 347 480 364
rect -480 300 480 347
rect 538 347 740 364
rect 1296 364 1312 381
rect 1742 381 2330 397
rect 1742 364 1758 381
rect 1296 347 1498 364
rect 538 300 1498 347
rect 1556 347 1758 364
rect 2314 364 2330 381
rect 2760 381 3348 397
rect 2760 364 2776 381
rect 2314 347 2516 364
rect 1556 300 2516 347
rect 2574 347 2776 364
rect 3332 364 3348 381
rect 3778 381 4366 397
rect 3778 364 3794 381
rect 3332 347 3534 364
rect 2574 300 3534 347
rect 3592 347 3794 364
rect 4350 364 4366 381
rect 4796 381 5384 397
rect 4796 364 4812 381
rect 4350 347 4552 364
rect 3592 300 4552 347
rect 4610 347 4812 364
rect 5368 364 5384 381
rect 5814 381 6402 397
rect 5814 364 5830 381
rect 5368 347 5570 364
rect 4610 300 5570 347
rect 5628 347 5830 364
rect 6386 364 6402 381
rect 6832 381 7420 397
rect 6832 364 6848 381
rect 6386 347 6588 364
rect 5628 300 6588 347
rect 6646 347 6848 364
rect 7404 364 7420 381
rect 7404 347 7606 364
rect 6646 300 7606 347
rect -7606 -347 -6646 -300
rect -7606 -364 -7404 -347
rect -7420 -381 -7404 -364
rect -6848 -364 -6646 -347
rect -6588 -347 -5628 -300
rect -6588 -364 -6386 -347
rect -6848 -381 -6832 -364
rect -7420 -397 -6832 -381
rect -6402 -381 -6386 -364
rect -5830 -364 -5628 -347
rect -5570 -347 -4610 -300
rect -5570 -364 -5368 -347
rect -5830 -381 -5814 -364
rect -6402 -397 -5814 -381
rect -5384 -381 -5368 -364
rect -4812 -364 -4610 -347
rect -4552 -347 -3592 -300
rect -4552 -364 -4350 -347
rect -4812 -381 -4796 -364
rect -5384 -397 -4796 -381
rect -4366 -381 -4350 -364
rect -3794 -364 -3592 -347
rect -3534 -347 -2574 -300
rect -3534 -364 -3332 -347
rect -3794 -381 -3778 -364
rect -4366 -397 -3778 -381
rect -3348 -381 -3332 -364
rect -2776 -364 -2574 -347
rect -2516 -347 -1556 -300
rect -2516 -364 -2314 -347
rect -2776 -381 -2760 -364
rect -3348 -397 -2760 -381
rect -2330 -381 -2314 -364
rect -1758 -364 -1556 -347
rect -1498 -347 -538 -300
rect -1498 -364 -1296 -347
rect -1758 -381 -1742 -364
rect -2330 -397 -1742 -381
rect -1312 -381 -1296 -364
rect -740 -364 -538 -347
rect -480 -347 480 -300
rect -480 -364 -278 -347
rect -740 -381 -724 -364
rect -1312 -397 -724 -381
rect -294 -381 -278 -364
rect 278 -364 480 -347
rect 538 -347 1498 -300
rect 538 -364 740 -347
rect 278 -381 294 -364
rect -294 -397 294 -381
rect 724 -381 740 -364
rect 1296 -364 1498 -347
rect 1556 -347 2516 -300
rect 1556 -364 1758 -347
rect 1296 -381 1312 -364
rect 724 -397 1312 -381
rect 1742 -381 1758 -364
rect 2314 -364 2516 -347
rect 2574 -347 3534 -300
rect 2574 -364 2776 -347
rect 2314 -381 2330 -364
rect 1742 -397 2330 -381
rect 2760 -381 2776 -364
rect 3332 -364 3534 -347
rect 3592 -347 4552 -300
rect 3592 -364 3794 -347
rect 3332 -381 3348 -364
rect 2760 -397 3348 -381
rect 3778 -381 3794 -364
rect 4350 -364 4552 -347
rect 4610 -347 5570 -300
rect 4610 -364 4812 -347
rect 4350 -381 4366 -364
rect 3778 -397 4366 -381
rect 4796 -381 4812 -364
rect 5368 -364 5570 -347
rect 5628 -347 6588 -300
rect 5628 -364 5830 -347
rect 5368 -381 5384 -364
rect 4796 -397 5384 -381
rect 5814 -381 5830 -364
rect 6386 -364 6588 -347
rect 6646 -347 7606 -300
rect 6646 -364 6848 -347
rect 6386 -381 6402 -364
rect 5814 -397 6402 -381
rect 6832 -381 6848 -364
rect 7404 -364 7606 -347
rect 7404 -381 7420 -364
rect 6832 -397 7420 -381
<< polycont >>
rect -7404 347 -6848 381
rect -6386 347 -5830 381
rect -5368 347 -4812 381
rect -4350 347 -3794 381
rect -3332 347 -2776 381
rect -2314 347 -1758 381
rect -1296 347 -740 381
rect -278 347 278 381
rect 740 347 1296 381
rect 1758 347 2314 381
rect 2776 347 3332 381
rect 3794 347 4350 381
rect 4812 347 5368 381
rect 5830 347 6386 381
rect 6848 347 7404 381
rect -7404 -381 -6848 -347
rect -6386 -381 -5830 -347
rect -5368 -381 -4812 -347
rect -4350 -381 -3794 -347
rect -3332 -381 -2776 -347
rect -2314 -381 -1758 -347
rect -1296 -381 -740 -347
rect -278 -381 278 -347
rect 740 -381 1296 -347
rect 1758 -381 2314 -347
rect 2776 -381 3332 -347
rect 3794 -381 4350 -347
rect 4812 -381 5368 -347
rect 5830 -381 6386 -347
rect 6848 -381 7404 -347
<< locali >>
rect -7420 347 -7404 381
rect -6848 347 -6832 381
rect -6402 347 -6386 381
rect -5830 347 -5814 381
rect -5384 347 -5368 381
rect -4812 347 -4796 381
rect -4366 347 -4350 381
rect -3794 347 -3778 381
rect -3348 347 -3332 381
rect -2776 347 -2760 381
rect -2330 347 -2314 381
rect -1758 347 -1742 381
rect -1312 347 -1296 381
rect -740 347 -724 381
rect -294 347 -278 381
rect 278 347 294 381
rect 724 347 740 381
rect 1296 347 1312 381
rect 1742 347 1758 381
rect 2314 347 2330 381
rect 2760 347 2776 381
rect 3332 347 3348 381
rect 3778 347 3794 381
rect 4350 347 4366 381
rect 4796 347 4812 381
rect 5368 347 5384 381
rect 5814 347 5830 381
rect 6386 347 6402 381
rect 6832 347 6848 381
rect 7404 347 7420 381
rect -7652 288 -7618 304
rect -7652 -304 -7618 -288
rect -6634 288 -6600 304
rect -6634 -304 -6600 -288
rect -5616 288 -5582 304
rect -5616 -304 -5582 -288
rect -4598 288 -4564 304
rect -4598 -304 -4564 -288
rect -3580 288 -3546 304
rect -3580 -304 -3546 -288
rect -2562 288 -2528 304
rect -2562 -304 -2528 -288
rect -1544 288 -1510 304
rect -1544 -304 -1510 -288
rect -526 288 -492 304
rect -526 -304 -492 -288
rect 492 288 526 304
rect 492 -304 526 -288
rect 1510 288 1544 304
rect 1510 -304 1544 -288
rect 2528 288 2562 304
rect 2528 -304 2562 -288
rect 3546 288 3580 304
rect 3546 -304 3580 -288
rect 4564 288 4598 304
rect 4564 -304 4598 -288
rect 5582 288 5616 304
rect 5582 -304 5616 -288
rect 6600 288 6634 304
rect 6600 -304 6634 -288
rect 7618 288 7652 304
rect 7618 -304 7652 -288
rect -7420 -381 -7404 -347
rect -6848 -381 -6832 -347
rect -6402 -381 -6386 -347
rect -5830 -381 -5814 -347
rect -5384 -381 -5368 -347
rect -4812 -381 -4796 -347
rect -4366 -381 -4350 -347
rect -3794 -381 -3778 -347
rect -3348 -381 -3332 -347
rect -2776 -381 -2760 -347
rect -2330 -381 -2314 -347
rect -1758 -381 -1742 -347
rect -1312 -381 -1296 -347
rect -740 -381 -724 -347
rect -294 -381 -278 -347
rect 278 -381 294 -347
rect 724 -381 740 -347
rect 1296 -381 1312 -347
rect 1742 -381 1758 -347
rect 2314 -381 2330 -347
rect 2760 -381 2776 -347
rect 3332 -381 3348 -347
rect 3778 -381 3794 -347
rect 4350 -381 4366 -347
rect 4796 -381 4812 -347
rect 5368 -381 5384 -347
rect 5814 -381 5830 -347
rect 6386 -381 6402 -347
rect 6832 -381 6848 -347
rect 7404 -381 7420 -347
<< viali >>
rect -7358 347 -6894 381
rect -6340 347 -5876 381
rect -5322 347 -4858 381
rect -4304 347 -3840 381
rect -3286 347 -2822 381
rect -2268 347 -1804 381
rect -1250 347 -786 381
rect -232 347 232 381
rect 786 347 1250 381
rect 1804 347 2268 381
rect 2822 347 3286 381
rect 3840 347 4304 381
rect 4858 347 5322 381
rect 5876 347 6340 381
rect 6894 347 7358 381
rect -7652 -288 -7618 288
rect -6634 -288 -6600 288
rect -5616 -288 -5582 288
rect -4598 -288 -4564 288
rect -3580 -288 -3546 288
rect -2562 -288 -2528 288
rect -1544 -288 -1510 288
rect -526 -288 -492 288
rect 492 -288 526 288
rect 1510 -288 1544 288
rect 2528 -288 2562 288
rect 3546 -288 3580 288
rect 4564 -288 4598 288
rect 5582 -288 5616 288
rect 6600 -288 6634 288
rect 7618 -288 7652 288
rect -7358 -381 -6894 -347
rect -6340 -381 -5876 -347
rect -5322 -381 -4858 -347
rect -4304 -381 -3840 -347
rect -3286 -381 -2822 -347
rect -2268 -381 -1804 -347
rect -1250 -381 -786 -347
rect -232 -381 232 -347
rect 786 -381 1250 -347
rect 1804 -381 2268 -347
rect 2822 -381 3286 -347
rect 3840 -381 4304 -347
rect 4858 -381 5322 -347
rect 5876 -381 6340 -347
rect 6894 -381 7358 -347
<< metal1 >>
rect -7370 381 -6882 387
rect -7370 347 -7358 381
rect -6894 347 -6882 381
rect -7370 341 -6882 347
rect -6352 381 -5864 387
rect -6352 347 -6340 381
rect -5876 347 -5864 381
rect -6352 341 -5864 347
rect -5334 381 -4846 387
rect -5334 347 -5322 381
rect -4858 347 -4846 381
rect -5334 341 -4846 347
rect -4316 381 -3828 387
rect -4316 347 -4304 381
rect -3840 347 -3828 381
rect -4316 341 -3828 347
rect -3298 381 -2810 387
rect -3298 347 -3286 381
rect -2822 347 -2810 381
rect -3298 341 -2810 347
rect -2280 381 -1792 387
rect -2280 347 -2268 381
rect -1804 347 -1792 381
rect -2280 341 -1792 347
rect -1262 381 -774 387
rect -1262 347 -1250 381
rect -786 347 -774 381
rect -1262 341 -774 347
rect -244 381 244 387
rect -244 347 -232 381
rect 232 347 244 381
rect -244 341 244 347
rect 774 381 1262 387
rect 774 347 786 381
rect 1250 347 1262 381
rect 774 341 1262 347
rect 1792 381 2280 387
rect 1792 347 1804 381
rect 2268 347 2280 381
rect 1792 341 2280 347
rect 2810 381 3298 387
rect 2810 347 2822 381
rect 3286 347 3298 381
rect 2810 341 3298 347
rect 3828 381 4316 387
rect 3828 347 3840 381
rect 4304 347 4316 381
rect 3828 341 4316 347
rect 4846 381 5334 387
rect 4846 347 4858 381
rect 5322 347 5334 381
rect 4846 341 5334 347
rect 5864 381 6352 387
rect 5864 347 5876 381
rect 6340 347 6352 381
rect 5864 341 6352 347
rect 6882 381 7370 387
rect 6882 347 6894 381
rect 7358 347 7370 381
rect 6882 341 7370 347
rect -7658 288 -7612 300
rect -7658 -288 -7652 288
rect -7618 -288 -7612 288
rect -7658 -300 -7612 -288
rect -6640 288 -6594 300
rect -6640 -288 -6634 288
rect -6600 -288 -6594 288
rect -6640 -300 -6594 -288
rect -5622 288 -5576 300
rect -5622 -288 -5616 288
rect -5582 -288 -5576 288
rect -5622 -300 -5576 -288
rect -4604 288 -4558 300
rect -4604 -288 -4598 288
rect -4564 -288 -4558 288
rect -4604 -300 -4558 -288
rect -3586 288 -3540 300
rect -3586 -288 -3580 288
rect -3546 -288 -3540 288
rect -3586 -300 -3540 -288
rect -2568 288 -2522 300
rect -2568 -288 -2562 288
rect -2528 -288 -2522 288
rect -2568 -300 -2522 -288
rect -1550 288 -1504 300
rect -1550 -288 -1544 288
rect -1510 -288 -1504 288
rect -1550 -300 -1504 -288
rect -532 288 -486 300
rect -532 -288 -526 288
rect -492 -288 -486 288
rect -532 -300 -486 -288
rect 486 288 532 300
rect 486 -288 492 288
rect 526 -288 532 288
rect 486 -300 532 -288
rect 1504 288 1550 300
rect 1504 -288 1510 288
rect 1544 -288 1550 288
rect 1504 -300 1550 -288
rect 2522 288 2568 300
rect 2522 -288 2528 288
rect 2562 -288 2568 288
rect 2522 -300 2568 -288
rect 3540 288 3586 300
rect 3540 -288 3546 288
rect 3580 -288 3586 288
rect 3540 -300 3586 -288
rect 4558 288 4604 300
rect 4558 -288 4564 288
rect 4598 -288 4604 288
rect 4558 -300 4604 -288
rect 5576 288 5622 300
rect 5576 -288 5582 288
rect 5616 -288 5622 288
rect 5576 -300 5622 -288
rect 6594 288 6640 300
rect 6594 -288 6600 288
rect 6634 -288 6640 288
rect 6594 -300 6640 -288
rect 7612 288 7658 300
rect 7612 -288 7618 288
rect 7652 -288 7658 288
rect 7612 -300 7658 -288
rect -7370 -347 -6882 -341
rect -7370 -381 -7358 -347
rect -6894 -381 -6882 -347
rect -7370 -387 -6882 -381
rect -6352 -347 -5864 -341
rect -6352 -381 -6340 -347
rect -5876 -381 -5864 -347
rect -6352 -387 -5864 -381
rect -5334 -347 -4846 -341
rect -5334 -381 -5322 -347
rect -4858 -381 -4846 -347
rect -5334 -387 -4846 -381
rect -4316 -347 -3828 -341
rect -4316 -381 -4304 -347
rect -3840 -381 -3828 -347
rect -4316 -387 -3828 -381
rect -3298 -347 -2810 -341
rect -3298 -381 -3286 -347
rect -2822 -381 -2810 -347
rect -3298 -387 -2810 -381
rect -2280 -347 -1792 -341
rect -2280 -381 -2268 -347
rect -1804 -381 -1792 -347
rect -2280 -387 -1792 -381
rect -1262 -347 -774 -341
rect -1262 -381 -1250 -347
rect -786 -381 -774 -347
rect -1262 -387 -774 -381
rect -244 -347 244 -341
rect -244 -381 -232 -347
rect 232 -381 244 -347
rect -244 -387 244 -381
rect 774 -347 1262 -341
rect 774 -381 786 -347
rect 1250 -381 1262 -347
rect 774 -387 1262 -381
rect 1792 -347 2280 -341
rect 1792 -381 1804 -347
rect 2268 -381 2280 -347
rect 1792 -387 2280 -381
rect 2810 -347 3298 -341
rect 2810 -381 2822 -347
rect 3286 -381 3298 -347
rect 2810 -387 3298 -381
rect 3828 -347 4316 -341
rect 3828 -381 3840 -347
rect 4304 -381 4316 -347
rect 3828 -387 4316 -381
rect 4846 -347 5334 -341
rect 4846 -381 4858 -347
rect 5322 -381 5334 -347
rect 4846 -387 5334 -381
rect 5864 -347 6352 -341
rect 5864 -381 5876 -347
rect 6340 -381 6352 -347
rect 5864 -387 6352 -381
rect 6882 -347 7370 -341
rect 6882 -381 6894 -347
rect 7358 -381 7370 -347
rect 6882 -387 7370 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 3 l 4.8 m 1 nf 15 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
