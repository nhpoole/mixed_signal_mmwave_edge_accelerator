magic
tech sky130A
timestamp 1624477805
<< pwell >>
rect 35 63 93 120
<< psubdiff >>
rect 44 100 85 112
rect 44 83 56 100
rect 73 83 85 100
rect 44 71 85 83
<< psubdiffcont >>
rect 56 83 73 100
<< locali >>
rect 44 100 85 112
rect 44 83 56 100
rect 73 83 85 100
rect 44 71 85 83
<< end >>
