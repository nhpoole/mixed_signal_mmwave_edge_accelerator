magic
tech sky130A
magscale 1 2
timestamp 1621481787
<< error_p >>
rect -1279 1000 777 1028
rect -1279 -1000 -1251 1000
rect -1235 960 733 984
rect -1211 936 733 960
rect -1211 -936 -1187 936
rect 685 -936 733 936
rect -1211 -960 733 -936
rect 709 -984 733 -960
rect 749 -1000 777 1000
rect -1279 -1028 777 -1000
<< mimcap2 >>
rect -1251 960 749 1000
rect -1251 -960 -1211 960
rect 709 -960 749 960
rect -1251 -1000 749 -960
<< mimcap2contact >>
rect -1211 -960 709 960
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -1351 -1100 849 1100
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
