magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1335 -1309 13342 19691
<< locali >>
rect 9082 11295 11998 11329
rect 3678 9881 11998 9915
rect 3678 8467 11998 8501
rect 3842 7350 3876 7832
rect 3657 7316 3876 7350
rect 6424 7053 11998 7087
rect 5992 5639 11998 5673
rect 4704 4225 11998 4259
rect 4704 2811 11998 2845
rect 3639 2541 3824 2575
rect 3639 2176 3673 2541
rect 3506 2142 3673 2176
rect 5072 1397 11998 1431
<< metal1 >>
rect 11966 11286 12030 11338
rect 2736 10629 3391 10657
rect 7586 10579 7650 10631
rect 11966 9872 12030 9924
rect 2652 9139 3391 9167
rect 3474 9127 3538 9179
rect 11966 8458 12030 8510
rect 2820 8200 3439 8228
rect 2652 7952 3539 7980
rect 8054 7751 8118 7803
rect 11966 7044 12030 7096
rect 5036 6337 5100 6389
rect 2736 6160 3672 6188
rect 2568 6036 3539 6064
rect 2904 5912 3406 5940
rect 11966 5630 12030 5682
rect 2652 5372 3406 5400
rect 2736 5248 3539 5276
rect 2988 5124 3672 5152
rect 4820 4923 4884 4975
rect 1553 4308 2652 4336
rect 11966 4216 12030 4268
rect 383 4148 3072 4176
rect 4178 3493 4242 3545
rect 3156 3332 3539 3360
rect 3072 3084 3439 3112
rect 11966 2802 12030 2854
rect 3875 2284 3939 2336
rect 3072 2145 3391 2173
rect 4546 2111 4610 2163
rect 11966 1388 12030 1440
rect 3359 643 3423 695
rect 9530 681 9594 733
rect 11966 -26 12030 26
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4322 1567 6401
rect 369 2828 397 4162
rect 137 2238 203 2290
rect 137 538 203 590
rect 2554 0 2582 11352
rect 2638 0 2666 11352
rect 2722 0 2750 11352
rect 2806 0 2834 11352
rect 2890 0 2918 11352
rect 2974 0 3002 11352
rect 3058 0 3086 11352
rect 3142 0 3170 11352
rect 11970 11288 12026 11336
rect 7618 10591 12082 10619
rect 11970 9874 12026 9922
rect 3492 8587 3520 9153
rect 11970 8460 12026 8508
rect 8086 7763 12082 7791
rect 11970 7046 12026 7094
rect 5068 6349 12082 6377
rect 11970 5632 12026 5680
rect 4852 4935 12082 4963
rect 11970 4218 12026 4266
rect 4182 3495 4238 3543
rect 11970 2804 12026 2852
rect 3879 2286 3935 2334
rect 4564 1571 4592 2137
rect 11970 1390 12026 1438
rect 9562 707 12082 721
rect 9548 693 12082 707
rect 3377 655 3405 683
rect 9548 141 9576 693
rect 11970 -24 12026 24
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 11949 11263 12047 11361
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 11949 9849 12047 9947
rect 2568 8557 3506 8617
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 11949 8435 12047 8533
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 11949 7021 12047 7119
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 11949 5607 12047 5705
rect 11949 4193 12047 4291
rect 2820 3489 4210 3549
rect -49 2779 49 2877
rect 11949 2779 12047 2877
rect 2378 2295 2988 2355
rect 3156 2280 3907 2340
rect 1872 1913 2904 1973
rect 2736 1541 4578 1601
rect -49 1365 49 1463
rect 11949 1365 12047 1463
rect 1872 855 3156 915
rect 3072 111 9562 171
rect -49 -49 49 49
rect 11949 -49 12047 49
use sky130_sram_2kbyte_1rw1r_32x512_8_dff_buf_array  sky130_sram_2kbyte_1rw1r_32x512_8_dff_buf_array_0
timestamp 1626486988
transform 1 0 0 0 1 0
box -49 -49 2590 2877
use sky130_sram_2kbyte_1rw1r_32x512_8_pand3  sky130_sram_2kbyte_1rw1r_32x512_8_pand3_0
timestamp 1626486988
transform 1 0 3310 0 1 5656
box -36 -17 3150 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1_1
timestamp 1626486988
transform 1 0 3678 0 -1 2828
box -36 -17 1430 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1_0
timestamp 1626486988
transform 1 0 3310 0 1 2828
box -36 -17 1430 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_delay_chain  sky130_sram_2kbyte_1rw1r_32x512_8_delay_chain_0
timestamp 1626486988
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
use sky130_sram_2kbyte_1rw1r_32x512_8_pand3_0  sky130_sram_2kbyte_1rw1r_32x512_8_pand3_0_0
timestamp 1626486988
transform 1 0 3310 0 -1 5656
box -36 -17 2718 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_2  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_2_0
timestamp 1626486988
transform 1 0 3310 0 1 0
box -36 -17 8724 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pnand2_1  sky130_sram_2kbyte_1rw1r_32x512_8_pnand2_1_0
timestamp 1626486988
transform 1 0 3310 0 -1 8484
box -36 -17 504 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_1  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_1_1
timestamp 1626486988
transform 1 0 3310 0 1 8484
box -36 -17 404 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_1  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_1_0
timestamp 1626486988
transform 1 0 3310 0 -1 2828
box -36 -17 404 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3_1
timestamp 1626486988
transform 1 0 3310 0 -1 11312
box -36 -17 5808 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3_0
timestamp 1626486988
transform 1 0 3778 0 -1 8484
box -36 -17 5808 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 11966 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626486988
transform 1 0 11969 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_0
timestamp 1626486988
transform 1 0 9529 0 1 104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 8054 0 1 7745
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626486988
transform 1 0 9530 0 1 675
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626486988
transform 1 0 9533 0 1 674
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626486988
transform 1 0 11965 0 1 8447
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626486988
transform 1 0 11966 0 1 8452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626486988
transform 1 0 11969 0 1 8451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626486988
transform 1 0 9530 0 1 675
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626486988
transform 1 0 9533 0 1 674
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1626486988
transform 1 0 8057 0 1 7744
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626486988
transform 1 0 11965 0 1 8447
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626486988
transform 1 0 11966 0 1 8452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1626486988
transform 1 0 11969 0 1 8451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626486988
transform 1 0 11965 0 1 7033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626486988
transform 1 0 11966 0 1 7038
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1626486988
transform 1 0 11969 0 1 7037
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626486988
transform 1 0 11965 0 1 5619
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626486988
transform 1 0 11966 0 1 5624
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1626486988
transform 1 0 11969 0 1 5623
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626486988
transform 1 0 11965 0 1 7033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626486988
transform 1 0 11966 0 1 7038
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1626486988
transform 1 0 11969 0 1 7037
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626486988
transform 1 0 11965 0 1 5619
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626486988
transform 1 0 11966 0 1 5624
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1626486988
transform 1 0 11969 0 1 5623
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626486988
transform 1 0 11965 0 1 4205
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626486988
transform 1 0 11966 0 1 4210
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1626486988
transform 1 0 11969 0 1 4209
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626486988
transform 1 0 11965 0 1 2791
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626486988
transform 1 0 11966 0 1 2796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1626486988
transform 1 0 11969 0 1 2795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626486988
transform 1 0 11965 0 1 4205
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626486988
transform 1 0 11966 0 1 4210
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1626486988
transform 1 0 11969 0 1 4209
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626486988
transform 1 0 11965 0 1 2791
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626486988
transform 1 0 11966 0 1 2796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1626486988
transform 1 0 11969 0 1 2795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626486988
transform 1 0 11965 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1626486988
transform 1 0 11966 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1626486988
transform 1 0 11969 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626486988
transform 1 0 11965 0 1 -37
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1626486988
transform 1 0 11966 0 1 -32
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1626486988
transform 1 0 11969 0 1 -33
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626486988
transform 1 0 11965 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1626486988
transform 1 0 3040 0 1 4130
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1626486988
transform 1 0 351 0 1 4130
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626486988
transform 1 0 2345 0 1 2288
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_1
timestamp 1626486988
transform 1 0 2955 0 1 2288
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626486988
transform 1 0 1839 0 1 1906
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_2
timestamp 1626486988
transform 1 0 2871 0 1 1906
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626486988
transform 1 0 1839 0 1 848
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_3
timestamp 1626486988
transform 1 0 3123 0 1 848
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1626486988
transform 1 0 4178 0 1 3487
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1626486988
transform 1 0 4181 0 1 3486
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626486988
transform 1 0 4177 0 1 3482
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1626486988
transform 1 0 4178 0 1 3487
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1626486988
transform 1 0 4181 0 1 3486
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_4
timestamp 1626486988
transform 1 0 2787 0 1 3482
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1626486988
transform 1 0 3510 0 1 3313
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1626486988
transform 1 0 3124 0 1 3314
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1626486988
transform 1 0 3410 0 1 3065
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1626486988
transform 1 0 3040 0 1 3066
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1626486988
transform 1 0 4546 0 1 2105
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_20
timestamp 1626486988
transform 1 0 4549 0 1 2104
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_5
timestamp 1626486988
transform 1 0 2703 0 1 1534
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_6
timestamp 1626486988
transform 1 0 4545 0 1 1534
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1626486988
transform 1 0 3874 0 1 2273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1626486988
transform 1 0 3875 0 1 2278
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_21
timestamp 1626486988
transform 1 0 3878 0 1 2277
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1626486988
transform 1 0 3874 0 1 2273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1626486988
transform 1 0 3875 0 1 2278
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_22
timestamp 1626486988
transform 1 0 3878 0 1 2277
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_7
timestamp 1626486988
transform 1 0 3123 0 1 2273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_23
timestamp 1626486988
transform 1 0 3362 0 1 2126
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1626486988
transform 1 0 3040 0 1 2127
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_8
timestamp 1626486988
transform 1 0 3039 0 1 104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1626486988
transform 1 0 3359 0 1 637
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_24
timestamp 1626486988
transform 1 0 3362 0 1 636
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_25
timestamp 1626486988
transform 1 0 3510 0 1 7933
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1626486988
transform 1 0 2620 0 1 7934
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_26
timestamp 1626486988
transform 1 0 3410 0 1 8181
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1626486988
transform 1 0 2788 0 1 8182
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1626486988
transform 1 0 2620 0 1 4290
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1626486988
transform 1 0 1521 0 1 4290
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1626486988
transform 1 0 4820 0 1 4917
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_27
timestamp 1626486988
transform 1 0 4823 0 1 4916
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_28
timestamp 1626486988
transform 1 0 3643 0 1 5105
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1626486988
transform 1 0 2956 0 1 5106
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_29
timestamp 1626486988
transform 1 0 3510 0 1 5229
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1626486988
transform 1 0 2704 0 1 5230
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_30
timestamp 1626486988
transform 1 0 3377 0 1 5353
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1626486988
transform 1 0 2620 0 1 5354
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1626486988
transform 1 0 5036 0 1 6331
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_31
timestamp 1626486988
transform 1 0 5039 0 1 6330
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_32
timestamp 1626486988
transform 1 0 3643 0 1 6141
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_36
timestamp 1626486988
transform 1 0 2704 0 1 6142
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_33
timestamp 1626486988
transform 1 0 3510 0 1 6017
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_37
timestamp 1626486988
transform 1 0 2536 0 1 6018
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_34
timestamp 1626486988
transform 1 0 3377 0 1 5893
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_38
timestamp 1626486988
transform 1 0 2872 0 1 5894
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_35
timestamp 1626486988
transform 1 0 3362 0 1 9120
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_39
timestamp 1626486988
transform 1 0 2620 0 1 9121
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_40
timestamp 1626486988
transform 1 0 3474 0 1 9121
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_36
timestamp 1626486988
transform 1 0 3477 0 1 9120
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_9
timestamp 1626486988
transform 1 0 2535 0 1 8550
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_10
timestamp 1626486988
transform 1 0 3473 0 1 8550
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_41
timestamp 1626486988
transform 1 0 2704 0 1 10611
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_37
timestamp 1626486988
transform 1 0 3362 0 1 10610
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1626486988
transform 1 0 11965 0 1 11275
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_42
timestamp 1626486988
transform 1 0 11966 0 1 11280
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_38
timestamp 1626486988
transform 1 0 11969 0 1 11279
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1626486988
transform 1 0 11965 0 1 9861
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_43
timestamp 1626486988
transform 1 0 11966 0 1 9866
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_39
timestamp 1626486988
transform 1 0 11969 0 1 9865
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1626486988
transform 1 0 11965 0 1 9861
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_44
timestamp 1626486988
transform 1 0 11966 0 1 9866
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_40
timestamp 1626486988
transform 1 0 11969 0 1 9865
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_45
timestamp 1626486988
transform 1 0 7586 0 1 10573
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_41
timestamp 1626486988
transform 1 0 7589 0 1 10572
box 0 0 58 66
<< labels >>
rlabel metal3 s 1343 11263 1441 11361 4 vdd
rlabel metal3 s 11949 4193 12047 4291 4 vdd
rlabel metal3 s 607 8435 705 8533 4 vdd
rlabel metal3 s 607 11263 705 11361 4 vdd
rlabel metal3 s 1343 5607 1441 5705 4 vdd
rlabel metal3 s 607 5607 705 5705 4 vdd
rlabel metal3 s 1343 16919 1441 17017 4 vdd
rlabel metal3 s 1343 14091 1441 14189 4 vdd
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s 607 14091 705 14189 4 vdd
rlabel metal3 s 11949 1365 12047 1463 4 vdd
rlabel metal3 s 11949 9849 12047 9947 4 vdd
rlabel metal3 s 11949 7021 12047 7119 4 vdd
rlabel metal3 s 607 16919 705 17017 4 vdd
rlabel metal3 s 1343 8435 1441 8533 4 vdd
rlabel metal3 s 11949 2779 12047 2877 4 gnd
rlabel metal3 s 11949 5607 12047 5705 4 gnd
rlabel metal3 s 1343 7021 1441 7119 4 gnd
rlabel metal3 s 607 15505 705 15603 4 gnd
rlabel metal3 s 1343 9849 1441 9947 4 gnd
rlabel metal3 s -49 2779 49 2877 4 gnd
rlabel metal3 s 1343 12677 1441 12775 4 gnd
rlabel metal3 s 1343 18333 1441 18431 4 gnd
rlabel metal3 s 11949 8435 12047 8533 4 gnd
rlabel metal3 s 11949 11263 12047 11361 4 gnd
rlabel metal3 s 607 9849 705 9947 4 gnd
rlabel metal3 s 607 18333 705 18431 4 gnd
rlabel metal3 s 607 7021 705 7119 4 gnd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal3 s 1343 15505 1441 15603 4 gnd
rlabel metal3 s 11949 -49 12047 49 4 gnd
rlabel metal3 s 607 12677 705 12775 4 gnd
rlabel metal2 s 137 538 203 590 4 csb
rlabel metal2 s 137 2238 203 2290 4 web
rlabel metal2 s 7618 10591 12082 10619 4 wl_en
rlabel metal2 s 5068 6349 12082 6377 4 w_en
rlabel metal2 s 4852 4935 12082 4963 4 s_en
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
rlabel metal2 s 8086 7763 12082 7791 4 p_en_bar
rlabel metal2 s 3377 655 3405 683 4 clk
rlabel metal2 s 9562 693 12082 721 4 clk_buf
<< properties >>
string FIXED_BBOX 0 0 12082 18542
<< end >>
