../../30-open-magic-gds2spice-nobbox/outputs/design_extracted.spice