

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO deconv_kernel_estimator_top_level 
  PIN clk 
    ANTENNAPARTIALMETALAREA 6.3938 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.808 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 8.9508 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.208 LAYER met3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met3 ; 
    ANTENNAMAXAREACAR 16.6087 LAYER met3 ;
    ANTENNAMAXSIDEAREACAR 86.8212 LAYER met3 ;
    ANTENNAMAXCUTCAR 0.158681 LAYER via3 ;
  END clk
  PIN rst_n 
    ANTENNAPARTIALMETALAREA 73.5824 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 367.633 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.3518 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4 ; 
    ANTENNAMAXAREACAR 37.3026 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 189.04 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4 ;
  END rst_n
  PIN load_en 
    ANTENNAPARTIALMETALAREA 69.7464 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 348.453 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 37.8747 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 202.464 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4 ; 
    ANTENNAMAXAREACAR 58.3144 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 302.811 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END load_en
  PIN debug_en 
    ANTENNAPARTIALMETALAREA 47.3156 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 236.299 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ; 
    ANTENNAMAXAREACAR 18.8909 LAYER met3 ;
    ANTENNAMAXSIDEAREACAR 97.8239 LAYER met3 ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3 ;
  END debug_en
  PIN serial_in 
    ANTENNAPARTIALMETALAREA 72.3112 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 361.277 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.315 LAYER met4 ; 
    ANTENNAMAXAREACAR 27.3717 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 142.159 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.417143 LAYER via4 ;
  END serial_in
  PIN sram_select[1] 
    ANTENNAPARTIALMETALAREA 151.739 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 758.415 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4 ; 
    ANTENNAMAXAREACAR 39.2394 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 202.122 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4 ;
  END sram_select[1]
  PIN sram_select[0] 
    ANTENNAPARTIALMETALAREA 94.3528 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 471.485 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.3518 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4 ; 
    ANTENNAMAXAREACAR 55.8402 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 288.254 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4 ;
  END sram_select[0]
  PIN frequency_adc_done 
    ANTENNAPARTIALMETALAREA 132.259 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 661.014 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.5588 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4 ; 
    ANTENNAMAXAREACAR 41.7831 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 216.089 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4 ;
  END frequency_adc_done
  PIN amplitude_adc_done 
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 32.071 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 171.512 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNADIFFAREA 2.6082 LAYER met5 ; 
    ANTENNAPARTIALMETALAREA 684.832 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 1031.09 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7672 LAYER met5 ; 
    ANTENNAMAXAREACAR 257.092 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 402.468 LAYER met5 ;
  END amplitude_adc_done
  PIN sig_frequency[7] 
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 32.254 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 172.488 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.5558 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.976 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNADIFFAREA 2.6082 LAYER met5 ; 
    ANTENNAPARTIALMETALAREA 682.624 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 1027.78 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7672 LAYER met5 ; 
    ANTENNAMAXAREACAR 253.162 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 384.625 LAYER met5 ;
  END sig_frequency[7]
  PIN sig_frequency[6] 
    ANTENNAPARTIALMETALAREA 1.4026 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.734 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 143.665 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 766.68 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4 ; 
    ANTENNAMAXAREACAR 31.1539 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 157.504 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via4 ;
  END sig_frequency[6]
  PIN sig_frequency[5] 
    ANTENNAPARTIALMETALAREA 19.177 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 95.606 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 7.873 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 10.7808 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.968 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4 ; 
    ANTENNAMAXAREACAR 62.6131 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 327.776 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via4 ;
  END sig_frequency[5]
  PIN sig_frequency[4] 
    ANTENNAPARTIALMETALAREA 36.747 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 183.456 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4 ; 
    ANTENNAMAXAREACAR 43.9033 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 225.135 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4 ;
  END sig_frequency[4]
  PIN sig_frequency[3] 
    ANTENNAPARTIALMETALAREA 60.4773 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 301.872 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 72.94 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 389.48 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 12.9288 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 69.424 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4 ; 
    ANTENNAMAXAREACAR 70.4721 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 367.642 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.450101 LAYER via4 ;
  END sig_frequency[3]
  PIN sig_frequency[2] 
    ANTENNAPARTIALMETALAREA 0.5746 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.765 LAYER met2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ; 
    ANTENNAMAXAREACAR 43.3657 LAYER met2 ;
    ANTENNAMAXSIDEAREACAR 212.211 LAYER met2 ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2 ;
  END sig_frequency[2]
  PIN sig_frequency[1] 
    ANTENNAPARTIALMETALAREA 1.0521 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0995 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNADIFFAREA 0.8694 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0284 LAYER met4 ; 
    ANTENNAMAXAREACAR 98.2655 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 474.81 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.166152 LAYER via4 ;
  END sig_frequency[1]
  PIN sig_frequency[0] 
    ANTENNAPARTIALMETALAREA 117 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 584.721 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ; 
    ANTENNAMAXAREACAR 67.2619 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 346.528 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4 ;
  END sig_frequency[0]
  PIN sig_amplitude[7] 
    ANTENNAPARTIALMETALAREA 12.7036 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.056 LAYER met2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2 ; 
    ANTENNAMAXAREACAR 65.0117 LAYER met2 ;
    ANTENNAMAXSIDEAREACAR 318.707 LAYER met2 ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2 ;
  END sig_amplitude[7]
  PIN sig_amplitude[6] 
    ANTENNAPARTIALMETALAREA 149.769 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 748.682 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4 ; 
    ANTENNAMAXAREACAR 55.7883 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 285.249 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4 ;
  END sig_amplitude[6]
  PIN sig_amplitude[5] 
    ANTENNAPARTIALMETALAREA 2.2882 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.333 LAYER met2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2 ; 
    ANTENNAMAXAREACAR 41.7883 LAYER met2 ;
    ANTENNAMAXSIDEAREACAR 204.077 LAYER met2 ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2 ;
  END sig_amplitude[5]
  PIN sig_amplitude[4] 
    ANTENNAPARTIALMETALAREA 102.02 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 509.82 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4 ; 
    ANTENNAMAXAREACAR 38.2798 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 197.324 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4 ;
  END sig_amplitude[4]
  PIN sig_amplitude[3] 
    ANTENNAPARTIALMETALAREA 6.3903 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7905 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 26.626 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 142.472 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.5558 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.976 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNADIFFAREA 2.6082 LAYER met5 ; 
    ANTENNAPARTIALMETALAREA 702.496 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 1057.58 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8212 LAYER met5 ; 
    ANTENNAMAXAREACAR 256.51 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 393.526 LAYER met5 ;
  END sig_amplitude[3]
  PIN sig_amplitude[2] 
    ANTENNAPARTIALMETALAREA 61.8679 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 309.06 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4 ; 
    ANTENNAMAXAREACAR 36.1521 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 186.399 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4 ;
  END sig_amplitude[2]
  PIN sig_amplitude[1] 
    ANTENNAPARTIALMETALAREA 16.2263 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 80.7345 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 154.774 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 825.928 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 25.0648 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 130.024 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 38.24 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 65.04 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met5 ; 
    ANTENNAMAXAREACAR 267.897 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 700.784 LAYER met5 ;
  END sig_amplitude[1]
  PIN sig_amplitude[0] 
    ANTENNAPARTIALMETALAREA 15.796 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 78.701 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 26.812 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 143.464 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNADIFFAREA 2.6082 LAYER met5 ; 
    ANTENNAPARTIALMETALAREA 711.232 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 1070.69 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7672 LAYER met5 ; 
    ANTENNAMAXAREACAR 264.447 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 405.11 LAYER met5 ;
  END sig_amplitude[0]
  PIN adc_bypass_en 
    ANTENNAPARTIALMETALAREA 45.5446 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 227.444 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNADIFFAREA 0.4347 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6477 LAYER met4 ; 
    ANTENNAMAXAREACAR 61.0385 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 292.772 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.293933 LAYER via4 ;
  END adc_bypass_en
  PIN serial_out 
    ANTENNADIFFAREA 0.4455 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 91.4218 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 456.883 LAYER met2 ;
  END serial_out
  PIN serial_out_valid 
    ANTENNAPARTIALMETALAREA 10.8619 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.1485 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 31.933 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 170.776 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.6408 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNADIFFAREA 0.429 LAYER met5 ; 
    ANTENNAPARTIALMETALAREA 671.584 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 1011.22 LAYER met5 ;
  END serial_out_valid
  PIN freq_eval_done 
    ANTENNADIFFAREA 0.7952 LAYER met2 ; 
    ANTENNAPARTIALMETALAREA 146.33 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 731.423 LAYER met2 ;
  END freq_eval_done
END deconv_kernel_estimator_top_level

END LIBRARY
