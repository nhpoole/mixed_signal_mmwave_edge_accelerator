* Stimulus file.

.include ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota/se_fold_casc_wide_swing_ota_pex.spice
.include se_fold_casc_wide_swing_ota_lvs.spice

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice

.param vincm=1.4 vsig=0 vdd=1.8

x0 vip vim vo ibiasn VDD VSS se_fold_casc_wide_swing_ota_flat
*x1 vip vim vo ibiasn VDD VSS se_fold_casc_wide_swing_ota_lvs
vdd VDD VSS 'vdd'
vss VSS 0 0
vip vip VSS dc 'vincm+vsig' ac 1 0
vim vim VSS dc 'vincm-vsig'
ibias VDD ibiasn 10u

.options savecurrents
.save all
+ @m.xm5.msky130_fd_pr__nfet_01v8[id]
+ @m.xm5.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm7.msky130_fd_pr__nfet_01v8[id]
+ @m.xm7.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm10.msky130_fd_pr__nfet_01v8[id]
+ @m.xm10.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__pfet_01v8[id]
+ @m.xm12.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__pfet_01v8[cgd]
+ @m.xm15.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm15.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm15.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm27.msky130_fd_pr__nfet_01v8[id]
+ @m.xm27.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm31.msky130_fd_pr__pfet_01v8[id]
+ @m.xm31.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm31.msky130_fd_pr__pfet_01v8[cgd]
+ @m.xm32.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm32.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm32.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm33.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm33.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm34.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm34.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm35.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm35.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm36.msky130_fd_pr__pfet_01v8[id]
+ @m.xm36.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm37.msky130_fd_pr__pfet_01v8[id]
+ @m.xm37.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm38.msky130_fd_pr__pfet_01v8[id]
+ @m.xm38.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm39.msky130_fd_pr__pfet_01v8[id]
+ @m.xm39.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm40.msky130_fd_pr__pfet_01v8[id]
+ @m.xm40.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm41.msky130_fd_pr__nfet_01v8[id]
+ @m.xm41.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm42.msky130_fd_pr__nfet_01v8[id]
+ @m.xm42.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm43.msky130_fd_pr__nfet_01v8[id]
+ @m.xm43.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm44.msky130_fd_pr__nfet_01v8[id]
+ @m.xm44.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm45.msky130_fd_pr__nfet_01v8[id]
+ @m.xm45.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm51.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm51.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm51.msky130_fd_pr__nfet_01v8_lvt[cgd]
+ @m.xm53.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm53.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm53.msky130_fd_pr__nfet_01v8_lvt[cgd]

+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm1.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm2.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm6.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm8.msky130_fd_pr__pfet_01v8[id]
+ @m.xm8.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm8.msky130_fd_pr__pfet_01v8[cgd]
+ @m.xm9.msky130_fd_pr__pfet_01v8[id]
+ @m.xm9.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm9.msky130_fd_pr__pfet_01v8[cgd]
+ @m.xm11.msky130_fd_pr__nfet_01v8[id]
+ @m.xm11.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm11.msky130_fd_pr__nfet_01v8[cgd]
+ @m.xm13.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm13.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm14.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm14.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm16.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm16.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm17.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm17.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm18.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm18.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm19.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm19.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm20.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm20.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm21.msky130_fd_pr__nfet_01v8[id]
+ @m.xm21.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm22.msky130_fd_pr__nfet_01v8[id]
+ @m.xm22.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm23.msky130_fd_pr__pfet_01v8[id]
+ @m.xm23.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm24.msky130_fd_pr__pfet_01v8[id]
+ @m.xm24.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm25.msky130_fd_pr__pfet_01v8[id]
+ @m.xm25.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm26.msky130_fd_pr__nfet_01v8[id]
+ @m.xm26.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm28.msky130_fd_pr__nfet_01v8[id]
+ @m.xm28.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm28.msky130_fd_pr__nfet_01v8[cgd]
+ @m.xm29.msky130_fd_pr__nfet_01v8[id]
+ @m.xm29.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm30.msky130_fd_pr__pfet_01v8[id]
+ @m.xm30.msky130_fd_pr__pfet_01v8[vth]

*.op
*.print all
*write se_fold_casc_wide_swing_ota_lvs_op.raw

* Control Block 1
*.control
*    op
*    print all
*    ac dec 100 0.1 1g
*    *noise v(vo) vip dec 100 1 10meg
*    run
*    write se_fold_casc_wide_swing_ota_lvs_ac.raw
*    *setplot noise1
*    *write se_fold_casc_wide_swing_ota_lvs_noise1.raw v(onoise_spectrum) v(inoise_spectrum)
*    *setplot noise2
*    *write se_fold_casc_wide_swing_ota_lvs_noise2.raw v(onoise_total) v(inoise_total)
*    quit
*.endc

* Control Block 2
.ac dec 100 0.1 1g
.control
    let incm = 0.4
    while incm < 1.5
        set incm = $&incm
        alter @vip[dc]=$incm
        alter @vim[dc]=$incm
        run
        write se_fold_casc_wide_swing_ota_lvs_ac_{$incm}.raw
        let incm = incm + 0.1
    end
    quit
.endc

* Control Block 3
*.ac dec 100 0.1 1g
*.control
*    let temperature = -40
*    while temperature < 130
*        set temp = $&temperature
*        run
*        write se_fold_casc_wide_swing_ota_lvs_temp_{$temp}.raw
*        let temperature = temperature + 10
*    end
*    quit
*.endc

* Control Block 4
*.ac dec 100 0.1 1g
*.control
*    let supply = 1.62
*    while supply < 2
*        alterparam vdd = {$&supply}
*        reset
*        run
*        write se_fold_casc_wide_swing_ota_lvs_vdd_{$&supply}.raw
*        let supply = supply + 0.04
*    end
*    quit
*.endc