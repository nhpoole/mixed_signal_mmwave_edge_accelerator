magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -6360 436 10710 11660
<< nwell >>
rect -5058 4282 5458 10358
<< pwell >>
rect -5048 4116 5448 4268
rect -5048 1904 -4896 4116
rect 5296 1904 5448 4116
rect -5048 1752 5448 1904
<< psubdiff >>
rect -5022 4209 5422 4242
rect -5022 4175 -4849 4209
rect -4815 4175 -4781 4209
rect -4747 4175 -4713 4209
rect -4679 4175 -4645 4209
rect -4611 4175 -4577 4209
rect -4543 4175 -4509 4209
rect -4475 4175 -4441 4209
rect -4407 4175 -4373 4209
rect -4339 4175 -4305 4209
rect -4271 4175 -4237 4209
rect -4203 4175 -4169 4209
rect -4135 4175 -4101 4209
rect -4067 4175 -4033 4209
rect -3999 4175 -3965 4209
rect -3931 4175 -3897 4209
rect -3863 4175 -3829 4209
rect -3795 4175 -3761 4209
rect -3727 4175 -3693 4209
rect -3659 4175 -3625 4209
rect -3591 4175 -3557 4209
rect -3523 4175 -3489 4209
rect -3455 4175 -3421 4209
rect -3387 4175 -3353 4209
rect -3319 4175 -3285 4209
rect -3251 4175 -3217 4209
rect -3183 4175 -3149 4209
rect -3115 4175 -3081 4209
rect -3047 4175 -3013 4209
rect -2979 4175 -2945 4209
rect -2911 4175 -2877 4209
rect -2843 4175 -2809 4209
rect -2775 4175 -2741 4209
rect -2707 4175 -2673 4209
rect -2639 4175 -2605 4209
rect -2571 4175 -2537 4209
rect -2503 4175 -2469 4209
rect -2435 4175 -2401 4209
rect -2367 4175 -2333 4209
rect -2299 4175 -2265 4209
rect -2231 4175 -2197 4209
rect -2163 4175 -2129 4209
rect -2095 4175 -2061 4209
rect -2027 4175 -1993 4209
rect -1959 4175 -1925 4209
rect -1891 4175 -1857 4209
rect -1823 4175 -1789 4209
rect -1755 4175 -1721 4209
rect -1687 4175 -1653 4209
rect -1619 4175 -1585 4209
rect -1551 4175 -1517 4209
rect -1483 4175 -1449 4209
rect -1415 4175 -1381 4209
rect -1347 4175 -1313 4209
rect -1279 4175 -1245 4209
rect -1211 4175 -1177 4209
rect -1143 4175 -1109 4209
rect -1075 4175 -1041 4209
rect -1007 4175 -973 4209
rect -939 4175 -905 4209
rect -871 4175 -837 4209
rect -803 4175 -769 4209
rect -735 4175 -701 4209
rect -667 4175 -633 4209
rect -599 4175 -565 4209
rect -531 4175 -497 4209
rect -463 4175 -429 4209
rect -395 4175 -361 4209
rect -327 4175 -293 4209
rect -259 4175 -225 4209
rect -191 4175 -157 4209
rect -123 4175 -89 4209
rect -55 4175 -21 4209
rect 13 4175 47 4209
rect 81 4175 115 4209
rect 149 4175 183 4209
rect 217 4175 251 4209
rect 285 4175 319 4209
rect 353 4175 387 4209
rect 421 4175 455 4209
rect 489 4175 523 4209
rect 557 4175 591 4209
rect 625 4175 659 4209
rect 693 4175 727 4209
rect 761 4175 795 4209
rect 829 4175 863 4209
rect 897 4175 931 4209
rect 965 4175 999 4209
rect 1033 4175 1067 4209
rect 1101 4175 1135 4209
rect 1169 4175 1203 4209
rect 1237 4175 1271 4209
rect 1305 4175 1339 4209
rect 1373 4175 1407 4209
rect 1441 4175 1475 4209
rect 1509 4175 1543 4209
rect 1577 4175 1611 4209
rect 1645 4175 1679 4209
rect 1713 4175 1747 4209
rect 1781 4175 1815 4209
rect 1849 4175 1883 4209
rect 1917 4175 1951 4209
rect 1985 4175 2019 4209
rect 2053 4175 2087 4209
rect 2121 4175 2155 4209
rect 2189 4175 2223 4209
rect 2257 4175 2291 4209
rect 2325 4175 2359 4209
rect 2393 4175 2427 4209
rect 2461 4175 2495 4209
rect 2529 4175 2563 4209
rect 2597 4175 2631 4209
rect 2665 4175 2699 4209
rect 2733 4175 2767 4209
rect 2801 4175 2835 4209
rect 2869 4175 2903 4209
rect 2937 4175 2971 4209
rect 3005 4175 3039 4209
rect 3073 4175 3107 4209
rect 3141 4175 3175 4209
rect 3209 4175 3243 4209
rect 3277 4175 3311 4209
rect 3345 4175 3379 4209
rect 3413 4175 3447 4209
rect 3481 4175 3515 4209
rect 3549 4175 3583 4209
rect 3617 4175 3651 4209
rect 3685 4175 3719 4209
rect 3753 4175 3787 4209
rect 3821 4175 3855 4209
rect 3889 4175 3923 4209
rect 3957 4175 3991 4209
rect 4025 4175 4059 4209
rect 4093 4175 4127 4209
rect 4161 4175 4195 4209
rect 4229 4175 4263 4209
rect 4297 4175 4331 4209
rect 4365 4175 4399 4209
rect 4433 4175 4467 4209
rect 4501 4175 4535 4209
rect 4569 4175 4603 4209
rect 4637 4175 4671 4209
rect 4705 4175 4739 4209
rect 4773 4175 4807 4209
rect 4841 4175 4875 4209
rect 4909 4175 4943 4209
rect 4977 4175 5011 4209
rect 5045 4175 5079 4209
rect 5113 4175 5147 4209
rect 5181 4175 5215 4209
rect 5249 4175 5422 4209
rect -5022 4142 5422 4175
rect -5022 4047 -4922 4142
rect -5022 4013 -4989 4047
rect -4955 4013 -4922 4047
rect -5022 3979 -4922 4013
rect -5022 3945 -4989 3979
rect -4955 3945 -4922 3979
rect -5022 3911 -4922 3945
rect -5022 3877 -4989 3911
rect -4955 3877 -4922 3911
rect -5022 3843 -4922 3877
rect -5022 3809 -4989 3843
rect -4955 3809 -4922 3843
rect -5022 3775 -4922 3809
rect -5022 3741 -4989 3775
rect -4955 3741 -4922 3775
rect -5022 3707 -4922 3741
rect -5022 3673 -4989 3707
rect -4955 3673 -4922 3707
rect -5022 3639 -4922 3673
rect -5022 3605 -4989 3639
rect -4955 3605 -4922 3639
rect -5022 3571 -4922 3605
rect -5022 3537 -4989 3571
rect -4955 3537 -4922 3571
rect -5022 3503 -4922 3537
rect -5022 3469 -4989 3503
rect -4955 3469 -4922 3503
rect -5022 3435 -4922 3469
rect -5022 3401 -4989 3435
rect -4955 3401 -4922 3435
rect -5022 3367 -4922 3401
rect -5022 3333 -4989 3367
rect -4955 3333 -4922 3367
rect -5022 3299 -4922 3333
rect -5022 3265 -4989 3299
rect -4955 3265 -4922 3299
rect -5022 3231 -4922 3265
rect -5022 3197 -4989 3231
rect -4955 3197 -4922 3231
rect -5022 3163 -4922 3197
rect -5022 3129 -4989 3163
rect -4955 3129 -4922 3163
rect -5022 3095 -4922 3129
rect -5022 3061 -4989 3095
rect -4955 3061 -4922 3095
rect -5022 3027 -4922 3061
rect -5022 2993 -4989 3027
rect -4955 2993 -4922 3027
rect -5022 2959 -4922 2993
rect -5022 2925 -4989 2959
rect -4955 2925 -4922 2959
rect -5022 2891 -4922 2925
rect -5022 2857 -4989 2891
rect -4955 2857 -4922 2891
rect -5022 2823 -4922 2857
rect -5022 2789 -4989 2823
rect -4955 2789 -4922 2823
rect -5022 2755 -4922 2789
rect -5022 2721 -4989 2755
rect -4955 2721 -4922 2755
rect -5022 2687 -4922 2721
rect -5022 2653 -4989 2687
rect -4955 2653 -4922 2687
rect -5022 2619 -4922 2653
rect -5022 2585 -4989 2619
rect -4955 2585 -4922 2619
rect -5022 2551 -4922 2585
rect -5022 2517 -4989 2551
rect -4955 2517 -4922 2551
rect -5022 2483 -4922 2517
rect -5022 2449 -4989 2483
rect -4955 2449 -4922 2483
rect -5022 2415 -4922 2449
rect -5022 2381 -4989 2415
rect -4955 2381 -4922 2415
rect -5022 2347 -4922 2381
rect -5022 2313 -4989 2347
rect -4955 2313 -4922 2347
rect -5022 2279 -4922 2313
rect -5022 2245 -4989 2279
rect -4955 2245 -4922 2279
rect -5022 2211 -4922 2245
rect -5022 2177 -4989 2211
rect -4955 2177 -4922 2211
rect -5022 2143 -4922 2177
rect -5022 2109 -4989 2143
rect -4955 2109 -4922 2143
rect -5022 2075 -4922 2109
rect -5022 2041 -4989 2075
rect -4955 2041 -4922 2075
rect -5022 2007 -4922 2041
rect -5022 1973 -4989 2007
rect -4955 1973 -4922 2007
rect -5022 1878 -4922 1973
rect 5322 4047 5422 4142
rect 5322 4013 5355 4047
rect 5389 4013 5422 4047
rect 5322 3979 5422 4013
rect 5322 3945 5355 3979
rect 5389 3945 5422 3979
rect 5322 3911 5422 3945
rect 5322 3877 5355 3911
rect 5389 3877 5422 3911
rect 5322 3843 5422 3877
rect 5322 3809 5355 3843
rect 5389 3809 5422 3843
rect 5322 3775 5422 3809
rect 5322 3741 5355 3775
rect 5389 3741 5422 3775
rect 5322 3707 5422 3741
rect 5322 3673 5355 3707
rect 5389 3673 5422 3707
rect 5322 3639 5422 3673
rect 5322 3605 5355 3639
rect 5389 3605 5422 3639
rect 5322 3571 5422 3605
rect 5322 3537 5355 3571
rect 5389 3537 5422 3571
rect 5322 3503 5422 3537
rect 5322 3469 5355 3503
rect 5389 3469 5422 3503
rect 5322 3435 5422 3469
rect 5322 3401 5355 3435
rect 5389 3401 5422 3435
rect 5322 3367 5422 3401
rect 5322 3333 5355 3367
rect 5389 3333 5422 3367
rect 5322 3299 5422 3333
rect 5322 3265 5355 3299
rect 5389 3265 5422 3299
rect 5322 3231 5422 3265
rect 5322 3197 5355 3231
rect 5389 3197 5422 3231
rect 5322 3163 5422 3197
rect 5322 3129 5355 3163
rect 5389 3129 5422 3163
rect 5322 3095 5422 3129
rect 5322 3061 5355 3095
rect 5389 3061 5422 3095
rect 5322 3027 5422 3061
rect 5322 2993 5355 3027
rect 5389 2993 5422 3027
rect 5322 2959 5422 2993
rect 5322 2925 5355 2959
rect 5389 2925 5422 2959
rect 5322 2891 5422 2925
rect 5322 2857 5355 2891
rect 5389 2857 5422 2891
rect 5322 2823 5422 2857
rect 5322 2789 5355 2823
rect 5389 2789 5422 2823
rect 5322 2755 5422 2789
rect 5322 2721 5355 2755
rect 5389 2721 5422 2755
rect 5322 2687 5422 2721
rect 5322 2653 5355 2687
rect 5389 2653 5422 2687
rect 5322 2619 5422 2653
rect 5322 2585 5355 2619
rect 5389 2585 5422 2619
rect 5322 2551 5422 2585
rect 5322 2517 5355 2551
rect 5389 2517 5422 2551
rect 5322 2483 5422 2517
rect 5322 2449 5355 2483
rect 5389 2449 5422 2483
rect 5322 2415 5422 2449
rect 5322 2381 5355 2415
rect 5389 2381 5422 2415
rect 5322 2347 5422 2381
rect 5322 2313 5355 2347
rect 5389 2313 5422 2347
rect 5322 2279 5422 2313
rect 5322 2245 5355 2279
rect 5389 2245 5422 2279
rect 5322 2211 5422 2245
rect 5322 2177 5355 2211
rect 5389 2177 5422 2211
rect 5322 2143 5422 2177
rect 5322 2109 5355 2143
rect 5389 2109 5422 2143
rect 5322 2075 5422 2109
rect 5322 2041 5355 2075
rect 5389 2041 5422 2075
rect 5322 2007 5422 2041
rect 5322 1973 5355 2007
rect 5389 1973 5422 2007
rect 5322 1878 5422 1973
rect -5022 1845 5422 1878
rect -5022 1811 -4849 1845
rect -4815 1811 -4781 1845
rect -4747 1811 -4713 1845
rect -4679 1811 -4645 1845
rect -4611 1811 -4577 1845
rect -4543 1811 -4509 1845
rect -4475 1811 -4441 1845
rect -4407 1811 -4373 1845
rect -4339 1811 -4305 1845
rect -4271 1811 -4237 1845
rect -4203 1811 -4169 1845
rect -4135 1811 -4101 1845
rect -4067 1811 -4033 1845
rect -3999 1811 -3965 1845
rect -3931 1811 -3897 1845
rect -3863 1811 -3829 1845
rect -3795 1811 -3761 1845
rect -3727 1811 -3693 1845
rect -3659 1811 -3625 1845
rect -3591 1811 -3557 1845
rect -3523 1811 -3489 1845
rect -3455 1811 -3421 1845
rect -3387 1811 -3353 1845
rect -3319 1811 -3285 1845
rect -3251 1811 -3217 1845
rect -3183 1811 -3149 1845
rect -3115 1811 -3081 1845
rect -3047 1811 -3013 1845
rect -2979 1811 -2945 1845
rect -2911 1811 -2877 1845
rect -2843 1811 -2809 1845
rect -2775 1811 -2741 1845
rect -2707 1811 -2673 1845
rect -2639 1811 -2605 1845
rect -2571 1811 -2537 1845
rect -2503 1811 -2469 1845
rect -2435 1811 -2401 1845
rect -2367 1811 -2333 1845
rect -2299 1811 -2265 1845
rect -2231 1811 -2197 1845
rect -2163 1811 -2129 1845
rect -2095 1811 -2061 1845
rect -2027 1811 -1993 1845
rect -1959 1811 -1925 1845
rect -1891 1811 -1857 1845
rect -1823 1811 -1789 1845
rect -1755 1811 -1721 1845
rect -1687 1811 -1653 1845
rect -1619 1811 -1585 1845
rect -1551 1811 -1517 1845
rect -1483 1811 -1449 1845
rect -1415 1811 -1381 1845
rect -1347 1811 -1313 1845
rect -1279 1811 -1245 1845
rect -1211 1811 -1177 1845
rect -1143 1811 -1109 1845
rect -1075 1811 -1041 1845
rect -1007 1811 -973 1845
rect -939 1811 -905 1845
rect -871 1811 -837 1845
rect -803 1811 -769 1845
rect -735 1811 -701 1845
rect -667 1811 -633 1845
rect -599 1811 -565 1845
rect -531 1811 -497 1845
rect -463 1811 -429 1845
rect -395 1811 -361 1845
rect -327 1811 -293 1845
rect -259 1811 -225 1845
rect -191 1811 -157 1845
rect -123 1811 -89 1845
rect -55 1811 -21 1845
rect 13 1811 47 1845
rect 81 1811 115 1845
rect 149 1811 183 1845
rect 217 1811 251 1845
rect 285 1811 319 1845
rect 353 1811 387 1845
rect 421 1811 455 1845
rect 489 1811 523 1845
rect 557 1811 591 1845
rect 625 1811 659 1845
rect 693 1811 727 1845
rect 761 1811 795 1845
rect 829 1811 863 1845
rect 897 1811 931 1845
rect 965 1811 999 1845
rect 1033 1811 1067 1845
rect 1101 1811 1135 1845
rect 1169 1811 1203 1845
rect 1237 1811 1271 1845
rect 1305 1811 1339 1845
rect 1373 1811 1407 1845
rect 1441 1811 1475 1845
rect 1509 1811 1543 1845
rect 1577 1811 1611 1845
rect 1645 1811 1679 1845
rect 1713 1811 1747 1845
rect 1781 1811 1815 1845
rect 1849 1811 1883 1845
rect 1917 1811 1951 1845
rect 1985 1811 2019 1845
rect 2053 1811 2087 1845
rect 2121 1811 2155 1845
rect 2189 1811 2223 1845
rect 2257 1811 2291 1845
rect 2325 1811 2359 1845
rect 2393 1811 2427 1845
rect 2461 1811 2495 1845
rect 2529 1811 2563 1845
rect 2597 1811 2631 1845
rect 2665 1811 2699 1845
rect 2733 1811 2767 1845
rect 2801 1811 2835 1845
rect 2869 1811 2903 1845
rect 2937 1811 2971 1845
rect 3005 1811 3039 1845
rect 3073 1811 3107 1845
rect 3141 1811 3175 1845
rect 3209 1811 3243 1845
rect 3277 1811 3311 1845
rect 3345 1811 3379 1845
rect 3413 1811 3447 1845
rect 3481 1811 3515 1845
rect 3549 1811 3583 1845
rect 3617 1811 3651 1845
rect 3685 1811 3719 1845
rect 3753 1811 3787 1845
rect 3821 1811 3855 1845
rect 3889 1811 3923 1845
rect 3957 1811 3991 1845
rect 4025 1811 4059 1845
rect 4093 1811 4127 1845
rect 4161 1811 4195 1845
rect 4229 1811 4263 1845
rect 4297 1811 4331 1845
rect 4365 1811 4399 1845
rect 4433 1811 4467 1845
rect 4501 1811 4535 1845
rect 4569 1811 4603 1845
rect 4637 1811 4671 1845
rect 4705 1811 4739 1845
rect 4773 1811 4807 1845
rect 4841 1811 4875 1845
rect 4909 1811 4943 1845
rect 4977 1811 5011 1845
rect 5045 1811 5079 1845
rect 5113 1811 5147 1845
rect 5181 1811 5215 1845
rect 5249 1811 5422 1845
rect -5022 1778 5422 1811
<< nsubdiff >>
rect -5022 10289 5422 10322
rect -5022 10255 -4849 10289
rect -4815 10255 -4781 10289
rect -4747 10255 -4713 10289
rect -4679 10255 -4645 10289
rect -4611 10255 -4577 10289
rect -4543 10255 -4509 10289
rect -4475 10255 -4441 10289
rect -4407 10255 -4373 10289
rect -4339 10255 -4305 10289
rect -4271 10255 -4237 10289
rect -4203 10255 -4169 10289
rect -4135 10255 -4101 10289
rect -4067 10255 -4033 10289
rect -3999 10255 -3965 10289
rect -3931 10255 -3897 10289
rect -3863 10255 -3829 10289
rect -3795 10255 -3761 10289
rect -3727 10255 -3693 10289
rect -3659 10255 -3625 10289
rect -3591 10255 -3557 10289
rect -3523 10255 -3489 10289
rect -3455 10255 -3421 10289
rect -3387 10255 -3353 10289
rect -3319 10255 -3285 10289
rect -3251 10255 -3217 10289
rect -3183 10255 -3149 10289
rect -3115 10255 -3081 10289
rect -3047 10255 -3013 10289
rect -2979 10255 -2945 10289
rect -2911 10255 -2877 10289
rect -2843 10255 -2809 10289
rect -2775 10255 -2741 10289
rect -2707 10255 -2673 10289
rect -2639 10255 -2605 10289
rect -2571 10255 -2537 10289
rect -2503 10255 -2469 10289
rect -2435 10255 -2401 10289
rect -2367 10255 -2333 10289
rect -2299 10255 -2265 10289
rect -2231 10255 -2197 10289
rect -2163 10255 -2129 10289
rect -2095 10255 -2061 10289
rect -2027 10255 -1993 10289
rect -1959 10255 -1925 10289
rect -1891 10255 -1857 10289
rect -1823 10255 -1789 10289
rect -1755 10255 -1721 10289
rect -1687 10255 -1653 10289
rect -1619 10255 -1585 10289
rect -1551 10255 -1517 10289
rect -1483 10255 -1449 10289
rect -1415 10255 -1381 10289
rect -1347 10255 -1313 10289
rect -1279 10255 -1245 10289
rect -1211 10255 -1177 10289
rect -1143 10255 -1109 10289
rect -1075 10255 -1041 10289
rect -1007 10255 -973 10289
rect -939 10255 -905 10289
rect -871 10255 -837 10289
rect -803 10255 -769 10289
rect -735 10255 -701 10289
rect -667 10255 -633 10289
rect -599 10255 -565 10289
rect -531 10255 -497 10289
rect -463 10255 -429 10289
rect -395 10255 -361 10289
rect -327 10255 -293 10289
rect -259 10255 -225 10289
rect -191 10255 -157 10289
rect -123 10255 -89 10289
rect -55 10255 -21 10289
rect 13 10255 47 10289
rect 81 10255 115 10289
rect 149 10255 183 10289
rect 217 10255 251 10289
rect 285 10255 319 10289
rect 353 10255 387 10289
rect 421 10255 455 10289
rect 489 10255 523 10289
rect 557 10255 591 10289
rect 625 10255 659 10289
rect 693 10255 727 10289
rect 761 10255 795 10289
rect 829 10255 863 10289
rect 897 10255 931 10289
rect 965 10255 999 10289
rect 1033 10255 1067 10289
rect 1101 10255 1135 10289
rect 1169 10255 1203 10289
rect 1237 10255 1271 10289
rect 1305 10255 1339 10289
rect 1373 10255 1407 10289
rect 1441 10255 1475 10289
rect 1509 10255 1543 10289
rect 1577 10255 1611 10289
rect 1645 10255 1679 10289
rect 1713 10255 1747 10289
rect 1781 10255 1815 10289
rect 1849 10255 1883 10289
rect 1917 10255 1951 10289
rect 1985 10255 2019 10289
rect 2053 10255 2087 10289
rect 2121 10255 2155 10289
rect 2189 10255 2223 10289
rect 2257 10255 2291 10289
rect 2325 10255 2359 10289
rect 2393 10255 2427 10289
rect 2461 10255 2495 10289
rect 2529 10255 2563 10289
rect 2597 10255 2631 10289
rect 2665 10255 2699 10289
rect 2733 10255 2767 10289
rect 2801 10255 2835 10289
rect 2869 10255 2903 10289
rect 2937 10255 2971 10289
rect 3005 10255 3039 10289
rect 3073 10255 3107 10289
rect 3141 10255 3175 10289
rect 3209 10255 3243 10289
rect 3277 10255 3311 10289
rect 3345 10255 3379 10289
rect 3413 10255 3447 10289
rect 3481 10255 3515 10289
rect 3549 10255 3583 10289
rect 3617 10255 3651 10289
rect 3685 10255 3719 10289
rect 3753 10255 3787 10289
rect 3821 10255 3855 10289
rect 3889 10255 3923 10289
rect 3957 10255 3991 10289
rect 4025 10255 4059 10289
rect 4093 10255 4127 10289
rect 4161 10255 4195 10289
rect 4229 10255 4263 10289
rect 4297 10255 4331 10289
rect 4365 10255 4399 10289
rect 4433 10255 4467 10289
rect 4501 10255 4535 10289
rect 4569 10255 4603 10289
rect 4637 10255 4671 10289
rect 4705 10255 4739 10289
rect 4773 10255 4807 10289
rect 4841 10255 4875 10289
rect 4909 10255 4943 10289
rect 4977 10255 5011 10289
rect 5045 10255 5079 10289
rect 5113 10255 5147 10289
rect 5181 10255 5215 10289
rect 5249 10255 5422 10289
rect -5022 10222 5422 10255
rect -5022 10137 -4922 10222
rect -5022 10103 -4989 10137
rect -4955 10103 -4922 10137
rect -5022 10069 -4922 10103
rect -5022 10035 -4989 10069
rect -4955 10035 -4922 10069
rect -5022 10001 -4922 10035
rect -5022 9967 -4989 10001
rect -4955 9967 -4922 10001
rect -5022 9933 -4922 9967
rect -5022 9899 -4989 9933
rect -4955 9899 -4922 9933
rect -5022 9865 -4922 9899
rect -5022 9831 -4989 9865
rect -4955 9831 -4922 9865
rect -5022 9797 -4922 9831
rect -5022 9763 -4989 9797
rect -4955 9763 -4922 9797
rect -5022 9729 -4922 9763
rect -5022 9695 -4989 9729
rect -4955 9695 -4922 9729
rect -5022 9661 -4922 9695
rect -5022 9627 -4989 9661
rect -4955 9627 -4922 9661
rect -5022 9593 -4922 9627
rect -5022 9559 -4989 9593
rect -4955 9559 -4922 9593
rect -5022 9525 -4922 9559
rect -5022 9491 -4989 9525
rect -4955 9491 -4922 9525
rect -5022 9457 -4922 9491
rect -5022 9423 -4989 9457
rect -4955 9423 -4922 9457
rect -5022 9389 -4922 9423
rect -5022 9355 -4989 9389
rect -4955 9355 -4922 9389
rect -5022 9321 -4922 9355
rect -5022 9287 -4989 9321
rect -4955 9287 -4922 9321
rect -5022 9253 -4922 9287
rect -5022 9219 -4989 9253
rect -4955 9219 -4922 9253
rect -5022 9185 -4922 9219
rect -5022 9151 -4989 9185
rect -4955 9151 -4922 9185
rect -5022 9117 -4922 9151
rect -5022 9083 -4989 9117
rect -4955 9083 -4922 9117
rect -5022 9049 -4922 9083
rect -5022 9015 -4989 9049
rect -4955 9015 -4922 9049
rect -5022 8981 -4922 9015
rect -5022 8947 -4989 8981
rect -4955 8947 -4922 8981
rect -5022 8913 -4922 8947
rect -5022 8879 -4989 8913
rect -4955 8879 -4922 8913
rect -5022 8845 -4922 8879
rect -5022 8811 -4989 8845
rect -4955 8811 -4922 8845
rect -5022 8777 -4922 8811
rect -5022 8743 -4989 8777
rect -4955 8743 -4922 8777
rect -5022 8709 -4922 8743
rect -5022 8675 -4989 8709
rect -4955 8675 -4922 8709
rect -5022 8641 -4922 8675
rect -5022 8607 -4989 8641
rect -4955 8607 -4922 8641
rect -5022 8573 -4922 8607
rect -5022 8539 -4989 8573
rect -4955 8539 -4922 8573
rect -5022 8505 -4922 8539
rect -5022 8471 -4989 8505
rect -4955 8471 -4922 8505
rect -5022 8437 -4922 8471
rect -5022 8403 -4989 8437
rect -4955 8403 -4922 8437
rect -5022 8369 -4922 8403
rect -5022 8335 -4989 8369
rect -4955 8335 -4922 8369
rect -5022 8301 -4922 8335
rect -5022 8267 -4989 8301
rect -4955 8267 -4922 8301
rect -5022 8233 -4922 8267
rect -5022 8199 -4989 8233
rect -4955 8199 -4922 8233
rect -5022 8165 -4922 8199
rect -5022 8131 -4989 8165
rect -4955 8131 -4922 8165
rect -5022 8097 -4922 8131
rect -5022 8063 -4989 8097
rect -4955 8063 -4922 8097
rect -5022 8029 -4922 8063
rect -5022 7995 -4989 8029
rect -4955 7995 -4922 8029
rect -5022 7961 -4922 7995
rect -5022 7927 -4989 7961
rect -4955 7927 -4922 7961
rect -5022 7893 -4922 7927
rect -5022 7859 -4989 7893
rect -4955 7859 -4922 7893
rect -5022 7825 -4922 7859
rect -5022 7791 -4989 7825
rect -4955 7791 -4922 7825
rect -5022 7757 -4922 7791
rect -5022 7723 -4989 7757
rect -4955 7723 -4922 7757
rect -5022 7689 -4922 7723
rect -5022 7655 -4989 7689
rect -4955 7655 -4922 7689
rect -5022 7621 -4922 7655
rect -5022 7587 -4989 7621
rect -4955 7587 -4922 7621
rect -5022 7553 -4922 7587
rect -5022 7519 -4989 7553
rect -4955 7519 -4922 7553
rect -5022 7485 -4922 7519
rect -5022 7451 -4989 7485
rect -4955 7451 -4922 7485
rect -5022 7417 -4922 7451
rect -5022 7383 -4989 7417
rect -4955 7383 -4922 7417
rect -5022 7349 -4922 7383
rect -5022 7315 -4989 7349
rect -4955 7315 -4922 7349
rect -5022 7281 -4922 7315
rect -5022 7247 -4989 7281
rect -4955 7247 -4922 7281
rect -5022 7213 -4922 7247
rect -5022 7179 -4989 7213
rect -4955 7179 -4922 7213
rect -5022 7145 -4922 7179
rect -5022 7111 -4989 7145
rect -4955 7111 -4922 7145
rect -5022 7077 -4922 7111
rect -5022 7043 -4989 7077
rect -4955 7043 -4922 7077
rect -5022 7009 -4922 7043
rect -5022 6975 -4989 7009
rect -4955 6975 -4922 7009
rect -5022 6941 -4922 6975
rect -5022 6907 -4989 6941
rect -4955 6907 -4922 6941
rect -5022 6873 -4922 6907
rect -5022 6839 -4989 6873
rect -4955 6839 -4922 6873
rect -5022 6805 -4922 6839
rect -5022 6771 -4989 6805
rect -4955 6771 -4922 6805
rect -5022 6737 -4922 6771
rect -5022 6703 -4989 6737
rect -4955 6703 -4922 6737
rect -5022 6669 -4922 6703
rect -5022 6635 -4989 6669
rect -4955 6635 -4922 6669
rect -5022 6601 -4922 6635
rect -5022 6567 -4989 6601
rect -4955 6567 -4922 6601
rect -5022 6533 -4922 6567
rect -5022 6499 -4989 6533
rect -4955 6499 -4922 6533
rect -5022 6465 -4922 6499
rect -5022 6431 -4989 6465
rect -4955 6431 -4922 6465
rect -5022 6397 -4922 6431
rect -5022 6363 -4989 6397
rect -4955 6363 -4922 6397
rect -5022 6329 -4922 6363
rect -5022 6295 -4989 6329
rect -4955 6295 -4922 6329
rect -5022 6261 -4922 6295
rect -5022 6227 -4989 6261
rect -4955 6227 -4922 6261
rect -5022 6193 -4922 6227
rect -5022 6159 -4989 6193
rect -4955 6159 -4922 6193
rect -5022 6125 -4922 6159
rect -5022 6091 -4989 6125
rect -4955 6091 -4922 6125
rect -5022 6057 -4922 6091
rect -5022 6023 -4989 6057
rect -4955 6023 -4922 6057
rect -5022 5989 -4922 6023
rect -5022 5955 -4989 5989
rect -4955 5955 -4922 5989
rect -5022 5921 -4922 5955
rect -5022 5887 -4989 5921
rect -4955 5887 -4922 5921
rect -5022 5853 -4922 5887
rect -5022 5819 -4989 5853
rect -4955 5819 -4922 5853
rect -5022 5785 -4922 5819
rect -5022 5751 -4989 5785
rect -4955 5751 -4922 5785
rect -5022 5717 -4922 5751
rect -5022 5683 -4989 5717
rect -4955 5683 -4922 5717
rect -5022 5649 -4922 5683
rect -5022 5615 -4989 5649
rect -4955 5615 -4922 5649
rect -5022 5581 -4922 5615
rect -5022 5547 -4989 5581
rect -4955 5547 -4922 5581
rect -5022 5513 -4922 5547
rect -5022 5479 -4989 5513
rect -4955 5479 -4922 5513
rect -5022 5445 -4922 5479
rect -5022 5411 -4989 5445
rect -4955 5411 -4922 5445
rect -5022 5377 -4922 5411
rect -5022 5343 -4989 5377
rect -4955 5343 -4922 5377
rect -5022 5309 -4922 5343
rect -5022 5275 -4989 5309
rect -4955 5275 -4922 5309
rect -5022 5241 -4922 5275
rect -5022 5207 -4989 5241
rect -4955 5207 -4922 5241
rect -5022 5173 -4922 5207
rect -5022 5139 -4989 5173
rect -4955 5139 -4922 5173
rect -5022 5105 -4922 5139
rect -5022 5071 -4989 5105
rect -4955 5071 -4922 5105
rect -5022 5037 -4922 5071
rect -5022 5003 -4989 5037
rect -4955 5003 -4922 5037
rect -5022 4969 -4922 5003
rect -5022 4935 -4989 4969
rect -4955 4935 -4922 4969
rect -5022 4901 -4922 4935
rect -5022 4867 -4989 4901
rect -4955 4867 -4922 4901
rect -5022 4833 -4922 4867
rect -5022 4799 -4989 4833
rect -4955 4799 -4922 4833
rect -5022 4765 -4922 4799
rect -5022 4731 -4989 4765
rect -4955 4731 -4922 4765
rect -5022 4697 -4922 4731
rect -5022 4663 -4989 4697
rect -4955 4663 -4922 4697
rect -5022 4578 -4922 4663
rect 5322 10137 5422 10222
rect 5322 10103 5355 10137
rect 5389 10103 5422 10137
rect 5322 10069 5422 10103
rect 5322 10035 5355 10069
rect 5389 10035 5422 10069
rect 5322 10001 5422 10035
rect 5322 9967 5355 10001
rect 5389 9967 5422 10001
rect 5322 9933 5422 9967
rect 5322 9899 5355 9933
rect 5389 9899 5422 9933
rect 5322 9865 5422 9899
rect 5322 9831 5355 9865
rect 5389 9831 5422 9865
rect 5322 9797 5422 9831
rect 5322 9763 5355 9797
rect 5389 9763 5422 9797
rect 5322 9729 5422 9763
rect 5322 9695 5355 9729
rect 5389 9695 5422 9729
rect 5322 9661 5422 9695
rect 5322 9627 5355 9661
rect 5389 9627 5422 9661
rect 5322 9593 5422 9627
rect 5322 9559 5355 9593
rect 5389 9559 5422 9593
rect 5322 9525 5422 9559
rect 5322 9491 5355 9525
rect 5389 9491 5422 9525
rect 5322 9457 5422 9491
rect 5322 9423 5355 9457
rect 5389 9423 5422 9457
rect 5322 9389 5422 9423
rect 5322 9355 5355 9389
rect 5389 9355 5422 9389
rect 5322 9321 5422 9355
rect 5322 9287 5355 9321
rect 5389 9287 5422 9321
rect 5322 9253 5422 9287
rect 5322 9219 5355 9253
rect 5389 9219 5422 9253
rect 5322 9185 5422 9219
rect 5322 9151 5355 9185
rect 5389 9151 5422 9185
rect 5322 9117 5422 9151
rect 5322 9083 5355 9117
rect 5389 9083 5422 9117
rect 5322 9049 5422 9083
rect 5322 9015 5355 9049
rect 5389 9015 5422 9049
rect 5322 8981 5422 9015
rect 5322 8947 5355 8981
rect 5389 8947 5422 8981
rect 5322 8913 5422 8947
rect 5322 8879 5355 8913
rect 5389 8879 5422 8913
rect 5322 8845 5422 8879
rect 5322 8811 5355 8845
rect 5389 8811 5422 8845
rect 5322 8777 5422 8811
rect 5322 8743 5355 8777
rect 5389 8743 5422 8777
rect 5322 8709 5422 8743
rect 5322 8675 5355 8709
rect 5389 8675 5422 8709
rect 5322 8641 5422 8675
rect 5322 8607 5355 8641
rect 5389 8607 5422 8641
rect 5322 8573 5422 8607
rect 5322 8539 5355 8573
rect 5389 8539 5422 8573
rect 5322 8505 5422 8539
rect 5322 8471 5355 8505
rect 5389 8471 5422 8505
rect 5322 8437 5422 8471
rect 5322 8403 5355 8437
rect 5389 8403 5422 8437
rect 5322 8369 5422 8403
rect 5322 8335 5355 8369
rect 5389 8335 5422 8369
rect 5322 8301 5422 8335
rect 5322 8267 5355 8301
rect 5389 8267 5422 8301
rect 5322 8233 5422 8267
rect 5322 8199 5355 8233
rect 5389 8199 5422 8233
rect 5322 8165 5422 8199
rect 5322 8131 5355 8165
rect 5389 8131 5422 8165
rect 5322 8097 5422 8131
rect 5322 8063 5355 8097
rect 5389 8063 5422 8097
rect 5322 8029 5422 8063
rect 5322 7995 5355 8029
rect 5389 7995 5422 8029
rect 5322 7961 5422 7995
rect 5322 7927 5355 7961
rect 5389 7927 5422 7961
rect 5322 7893 5422 7927
rect 5322 7859 5355 7893
rect 5389 7859 5422 7893
rect 5322 7825 5422 7859
rect 5322 7791 5355 7825
rect 5389 7791 5422 7825
rect 5322 7757 5422 7791
rect 5322 7723 5355 7757
rect 5389 7723 5422 7757
rect 5322 7689 5422 7723
rect 5322 7655 5355 7689
rect 5389 7655 5422 7689
rect 5322 7621 5422 7655
rect 5322 7587 5355 7621
rect 5389 7587 5422 7621
rect 5322 7553 5422 7587
rect 5322 7519 5355 7553
rect 5389 7519 5422 7553
rect 5322 7485 5422 7519
rect 5322 7451 5355 7485
rect 5389 7451 5422 7485
rect 5322 7417 5422 7451
rect 5322 7383 5355 7417
rect 5389 7383 5422 7417
rect 5322 7349 5422 7383
rect 5322 7315 5355 7349
rect 5389 7315 5422 7349
rect 5322 7281 5422 7315
rect 5322 7247 5355 7281
rect 5389 7247 5422 7281
rect 5322 7213 5422 7247
rect 5322 7179 5355 7213
rect 5389 7179 5422 7213
rect 5322 7145 5422 7179
rect 5322 7111 5355 7145
rect 5389 7111 5422 7145
rect 5322 7077 5422 7111
rect 5322 7043 5355 7077
rect 5389 7043 5422 7077
rect 5322 7009 5422 7043
rect 5322 6975 5355 7009
rect 5389 6975 5422 7009
rect 5322 6941 5422 6975
rect 5322 6907 5355 6941
rect 5389 6907 5422 6941
rect 5322 6873 5422 6907
rect 5322 6839 5355 6873
rect 5389 6839 5422 6873
rect 5322 6805 5422 6839
rect 5322 6771 5355 6805
rect 5389 6771 5422 6805
rect 5322 6737 5422 6771
rect 5322 6703 5355 6737
rect 5389 6703 5422 6737
rect 5322 6669 5422 6703
rect 5322 6635 5355 6669
rect 5389 6635 5422 6669
rect 5322 6601 5422 6635
rect 5322 6567 5355 6601
rect 5389 6567 5422 6601
rect 5322 6533 5422 6567
rect 5322 6499 5355 6533
rect 5389 6499 5422 6533
rect 5322 6465 5422 6499
rect 5322 6431 5355 6465
rect 5389 6431 5422 6465
rect 5322 6397 5422 6431
rect 5322 6363 5355 6397
rect 5389 6363 5422 6397
rect 5322 6329 5422 6363
rect 5322 6295 5355 6329
rect 5389 6295 5422 6329
rect 5322 6261 5422 6295
rect 5322 6227 5355 6261
rect 5389 6227 5422 6261
rect 5322 6193 5422 6227
rect 5322 6159 5355 6193
rect 5389 6159 5422 6193
rect 5322 6125 5422 6159
rect 5322 6091 5355 6125
rect 5389 6091 5422 6125
rect 5322 6057 5422 6091
rect 5322 6023 5355 6057
rect 5389 6023 5422 6057
rect 5322 5989 5422 6023
rect 5322 5955 5355 5989
rect 5389 5955 5422 5989
rect 5322 5921 5422 5955
rect 5322 5887 5355 5921
rect 5389 5887 5422 5921
rect 5322 5853 5422 5887
rect 5322 5819 5355 5853
rect 5389 5819 5422 5853
rect 5322 5785 5422 5819
rect 5322 5751 5355 5785
rect 5389 5751 5422 5785
rect 5322 5717 5422 5751
rect 5322 5683 5355 5717
rect 5389 5683 5422 5717
rect 5322 5649 5422 5683
rect 5322 5615 5355 5649
rect 5389 5615 5422 5649
rect 5322 5581 5422 5615
rect 5322 5547 5355 5581
rect 5389 5547 5422 5581
rect 5322 5513 5422 5547
rect 5322 5479 5355 5513
rect 5389 5479 5422 5513
rect 5322 5445 5422 5479
rect 5322 5411 5355 5445
rect 5389 5411 5422 5445
rect 5322 5377 5422 5411
rect 5322 5343 5355 5377
rect 5389 5343 5422 5377
rect 5322 5309 5422 5343
rect 5322 5275 5355 5309
rect 5389 5275 5422 5309
rect 5322 5241 5422 5275
rect 5322 5207 5355 5241
rect 5389 5207 5422 5241
rect 5322 5173 5422 5207
rect 5322 5139 5355 5173
rect 5389 5139 5422 5173
rect 5322 5105 5422 5139
rect 5322 5071 5355 5105
rect 5389 5071 5422 5105
rect 5322 5037 5422 5071
rect 5322 5003 5355 5037
rect 5389 5003 5422 5037
rect 5322 4969 5422 5003
rect 5322 4935 5355 4969
rect 5389 4935 5422 4969
rect 5322 4901 5422 4935
rect 5322 4867 5355 4901
rect 5389 4867 5422 4901
rect 5322 4833 5422 4867
rect 5322 4799 5355 4833
rect 5389 4799 5422 4833
rect 5322 4765 5422 4799
rect 5322 4731 5355 4765
rect 5389 4731 5422 4765
rect 5322 4697 5422 4731
rect 5322 4663 5355 4697
rect 5389 4663 5422 4697
rect 5322 4578 5422 4663
rect -5022 4545 5422 4578
rect -5022 4511 -4849 4545
rect -4815 4511 -4781 4545
rect -4747 4511 -4713 4545
rect -4679 4511 -4645 4545
rect -4611 4511 -4577 4545
rect -4543 4511 -4509 4545
rect -4475 4511 -4441 4545
rect -4407 4511 -4373 4545
rect -4339 4511 -4305 4545
rect -4271 4511 -4237 4545
rect -4203 4511 -4169 4545
rect -4135 4511 -4101 4545
rect -4067 4511 -4033 4545
rect -3999 4511 -3965 4545
rect -3931 4511 -3897 4545
rect -3863 4511 -3829 4545
rect -3795 4511 -3761 4545
rect -3727 4511 -3693 4545
rect -3659 4511 -3625 4545
rect -3591 4511 -3557 4545
rect -3523 4511 -3489 4545
rect -3455 4511 -3421 4545
rect -3387 4511 -3353 4545
rect -3319 4511 -3285 4545
rect -3251 4511 -3217 4545
rect -3183 4511 -3149 4545
rect -3115 4511 -3081 4545
rect -3047 4511 -3013 4545
rect -2979 4511 -2945 4545
rect -2911 4511 -2877 4545
rect -2843 4511 -2809 4545
rect -2775 4511 -2741 4545
rect -2707 4511 -2673 4545
rect -2639 4511 -2605 4545
rect -2571 4511 -2537 4545
rect -2503 4511 -2469 4545
rect -2435 4511 -2401 4545
rect -2367 4511 -2333 4545
rect -2299 4511 -2265 4545
rect -2231 4511 -2197 4545
rect -2163 4511 -2129 4545
rect -2095 4511 -2061 4545
rect -2027 4511 -1993 4545
rect -1959 4511 -1925 4545
rect -1891 4511 -1857 4545
rect -1823 4511 -1789 4545
rect -1755 4511 -1721 4545
rect -1687 4511 -1653 4545
rect -1619 4511 -1585 4545
rect -1551 4511 -1517 4545
rect -1483 4511 -1449 4545
rect -1415 4511 -1381 4545
rect -1347 4511 -1313 4545
rect -1279 4511 -1245 4545
rect -1211 4511 -1177 4545
rect -1143 4511 -1109 4545
rect -1075 4511 -1041 4545
rect -1007 4511 -973 4545
rect -939 4511 -905 4545
rect -871 4511 -837 4545
rect -803 4511 -769 4545
rect -735 4511 -701 4545
rect -667 4511 -633 4545
rect -599 4511 -565 4545
rect -531 4511 -497 4545
rect -463 4511 -429 4545
rect -395 4511 -361 4545
rect -327 4511 -293 4545
rect -259 4511 -225 4545
rect -191 4511 -157 4545
rect -123 4511 -89 4545
rect -55 4511 -21 4545
rect 13 4511 47 4545
rect 81 4511 115 4545
rect 149 4511 183 4545
rect 217 4511 251 4545
rect 285 4511 319 4545
rect 353 4511 387 4545
rect 421 4511 455 4545
rect 489 4511 523 4545
rect 557 4511 591 4545
rect 625 4511 659 4545
rect 693 4511 727 4545
rect 761 4511 795 4545
rect 829 4511 863 4545
rect 897 4511 931 4545
rect 965 4511 999 4545
rect 1033 4511 1067 4545
rect 1101 4511 1135 4545
rect 1169 4511 1203 4545
rect 1237 4511 1271 4545
rect 1305 4511 1339 4545
rect 1373 4511 1407 4545
rect 1441 4511 1475 4545
rect 1509 4511 1543 4545
rect 1577 4511 1611 4545
rect 1645 4511 1679 4545
rect 1713 4511 1747 4545
rect 1781 4511 1815 4545
rect 1849 4511 1883 4545
rect 1917 4511 1951 4545
rect 1985 4511 2019 4545
rect 2053 4511 2087 4545
rect 2121 4511 2155 4545
rect 2189 4511 2223 4545
rect 2257 4511 2291 4545
rect 2325 4511 2359 4545
rect 2393 4511 2427 4545
rect 2461 4511 2495 4545
rect 2529 4511 2563 4545
rect 2597 4511 2631 4545
rect 2665 4511 2699 4545
rect 2733 4511 2767 4545
rect 2801 4511 2835 4545
rect 2869 4511 2903 4545
rect 2937 4511 2971 4545
rect 3005 4511 3039 4545
rect 3073 4511 3107 4545
rect 3141 4511 3175 4545
rect 3209 4511 3243 4545
rect 3277 4511 3311 4545
rect 3345 4511 3379 4545
rect 3413 4511 3447 4545
rect 3481 4511 3515 4545
rect 3549 4511 3583 4545
rect 3617 4511 3651 4545
rect 3685 4511 3719 4545
rect 3753 4511 3787 4545
rect 3821 4511 3855 4545
rect 3889 4511 3923 4545
rect 3957 4511 3991 4545
rect 4025 4511 4059 4545
rect 4093 4511 4127 4545
rect 4161 4511 4195 4545
rect 4229 4511 4263 4545
rect 4297 4511 4331 4545
rect 4365 4511 4399 4545
rect 4433 4511 4467 4545
rect 4501 4511 4535 4545
rect 4569 4511 4603 4545
rect 4637 4511 4671 4545
rect 4705 4511 4739 4545
rect 4773 4511 4807 4545
rect 4841 4511 4875 4545
rect 4909 4511 4943 4545
rect 4977 4511 5011 4545
rect 5045 4511 5079 4545
rect 5113 4511 5147 4545
rect 5181 4511 5215 4545
rect 5249 4511 5422 4545
rect -5022 4478 5422 4511
<< psubdiffcont >>
rect -4849 4175 -4815 4209
rect -4781 4175 -4747 4209
rect -4713 4175 -4679 4209
rect -4645 4175 -4611 4209
rect -4577 4175 -4543 4209
rect -4509 4175 -4475 4209
rect -4441 4175 -4407 4209
rect -4373 4175 -4339 4209
rect -4305 4175 -4271 4209
rect -4237 4175 -4203 4209
rect -4169 4175 -4135 4209
rect -4101 4175 -4067 4209
rect -4033 4175 -3999 4209
rect -3965 4175 -3931 4209
rect -3897 4175 -3863 4209
rect -3829 4175 -3795 4209
rect -3761 4175 -3727 4209
rect -3693 4175 -3659 4209
rect -3625 4175 -3591 4209
rect -3557 4175 -3523 4209
rect -3489 4175 -3455 4209
rect -3421 4175 -3387 4209
rect -3353 4175 -3319 4209
rect -3285 4175 -3251 4209
rect -3217 4175 -3183 4209
rect -3149 4175 -3115 4209
rect -3081 4175 -3047 4209
rect -3013 4175 -2979 4209
rect -2945 4175 -2911 4209
rect -2877 4175 -2843 4209
rect -2809 4175 -2775 4209
rect -2741 4175 -2707 4209
rect -2673 4175 -2639 4209
rect -2605 4175 -2571 4209
rect -2537 4175 -2503 4209
rect -2469 4175 -2435 4209
rect -2401 4175 -2367 4209
rect -2333 4175 -2299 4209
rect -2265 4175 -2231 4209
rect -2197 4175 -2163 4209
rect -2129 4175 -2095 4209
rect -2061 4175 -2027 4209
rect -1993 4175 -1959 4209
rect -1925 4175 -1891 4209
rect -1857 4175 -1823 4209
rect -1789 4175 -1755 4209
rect -1721 4175 -1687 4209
rect -1653 4175 -1619 4209
rect -1585 4175 -1551 4209
rect -1517 4175 -1483 4209
rect -1449 4175 -1415 4209
rect -1381 4175 -1347 4209
rect -1313 4175 -1279 4209
rect -1245 4175 -1211 4209
rect -1177 4175 -1143 4209
rect -1109 4175 -1075 4209
rect -1041 4175 -1007 4209
rect -973 4175 -939 4209
rect -905 4175 -871 4209
rect -837 4175 -803 4209
rect -769 4175 -735 4209
rect -701 4175 -667 4209
rect -633 4175 -599 4209
rect -565 4175 -531 4209
rect -497 4175 -463 4209
rect -429 4175 -395 4209
rect -361 4175 -327 4209
rect -293 4175 -259 4209
rect -225 4175 -191 4209
rect -157 4175 -123 4209
rect -89 4175 -55 4209
rect -21 4175 13 4209
rect 47 4175 81 4209
rect 115 4175 149 4209
rect 183 4175 217 4209
rect 251 4175 285 4209
rect 319 4175 353 4209
rect 387 4175 421 4209
rect 455 4175 489 4209
rect 523 4175 557 4209
rect 591 4175 625 4209
rect 659 4175 693 4209
rect 727 4175 761 4209
rect 795 4175 829 4209
rect 863 4175 897 4209
rect 931 4175 965 4209
rect 999 4175 1033 4209
rect 1067 4175 1101 4209
rect 1135 4175 1169 4209
rect 1203 4175 1237 4209
rect 1271 4175 1305 4209
rect 1339 4175 1373 4209
rect 1407 4175 1441 4209
rect 1475 4175 1509 4209
rect 1543 4175 1577 4209
rect 1611 4175 1645 4209
rect 1679 4175 1713 4209
rect 1747 4175 1781 4209
rect 1815 4175 1849 4209
rect 1883 4175 1917 4209
rect 1951 4175 1985 4209
rect 2019 4175 2053 4209
rect 2087 4175 2121 4209
rect 2155 4175 2189 4209
rect 2223 4175 2257 4209
rect 2291 4175 2325 4209
rect 2359 4175 2393 4209
rect 2427 4175 2461 4209
rect 2495 4175 2529 4209
rect 2563 4175 2597 4209
rect 2631 4175 2665 4209
rect 2699 4175 2733 4209
rect 2767 4175 2801 4209
rect 2835 4175 2869 4209
rect 2903 4175 2937 4209
rect 2971 4175 3005 4209
rect 3039 4175 3073 4209
rect 3107 4175 3141 4209
rect 3175 4175 3209 4209
rect 3243 4175 3277 4209
rect 3311 4175 3345 4209
rect 3379 4175 3413 4209
rect 3447 4175 3481 4209
rect 3515 4175 3549 4209
rect 3583 4175 3617 4209
rect 3651 4175 3685 4209
rect 3719 4175 3753 4209
rect 3787 4175 3821 4209
rect 3855 4175 3889 4209
rect 3923 4175 3957 4209
rect 3991 4175 4025 4209
rect 4059 4175 4093 4209
rect 4127 4175 4161 4209
rect 4195 4175 4229 4209
rect 4263 4175 4297 4209
rect 4331 4175 4365 4209
rect 4399 4175 4433 4209
rect 4467 4175 4501 4209
rect 4535 4175 4569 4209
rect 4603 4175 4637 4209
rect 4671 4175 4705 4209
rect 4739 4175 4773 4209
rect 4807 4175 4841 4209
rect 4875 4175 4909 4209
rect 4943 4175 4977 4209
rect 5011 4175 5045 4209
rect 5079 4175 5113 4209
rect 5147 4175 5181 4209
rect 5215 4175 5249 4209
rect -4989 4013 -4955 4047
rect -4989 3945 -4955 3979
rect -4989 3877 -4955 3911
rect -4989 3809 -4955 3843
rect -4989 3741 -4955 3775
rect -4989 3673 -4955 3707
rect -4989 3605 -4955 3639
rect -4989 3537 -4955 3571
rect -4989 3469 -4955 3503
rect -4989 3401 -4955 3435
rect -4989 3333 -4955 3367
rect -4989 3265 -4955 3299
rect -4989 3197 -4955 3231
rect -4989 3129 -4955 3163
rect -4989 3061 -4955 3095
rect -4989 2993 -4955 3027
rect -4989 2925 -4955 2959
rect -4989 2857 -4955 2891
rect -4989 2789 -4955 2823
rect -4989 2721 -4955 2755
rect -4989 2653 -4955 2687
rect -4989 2585 -4955 2619
rect -4989 2517 -4955 2551
rect -4989 2449 -4955 2483
rect -4989 2381 -4955 2415
rect -4989 2313 -4955 2347
rect -4989 2245 -4955 2279
rect -4989 2177 -4955 2211
rect -4989 2109 -4955 2143
rect -4989 2041 -4955 2075
rect -4989 1973 -4955 2007
rect 5355 4013 5389 4047
rect 5355 3945 5389 3979
rect 5355 3877 5389 3911
rect 5355 3809 5389 3843
rect 5355 3741 5389 3775
rect 5355 3673 5389 3707
rect 5355 3605 5389 3639
rect 5355 3537 5389 3571
rect 5355 3469 5389 3503
rect 5355 3401 5389 3435
rect 5355 3333 5389 3367
rect 5355 3265 5389 3299
rect 5355 3197 5389 3231
rect 5355 3129 5389 3163
rect 5355 3061 5389 3095
rect 5355 2993 5389 3027
rect 5355 2925 5389 2959
rect 5355 2857 5389 2891
rect 5355 2789 5389 2823
rect 5355 2721 5389 2755
rect 5355 2653 5389 2687
rect 5355 2585 5389 2619
rect 5355 2517 5389 2551
rect 5355 2449 5389 2483
rect 5355 2381 5389 2415
rect 5355 2313 5389 2347
rect 5355 2245 5389 2279
rect 5355 2177 5389 2211
rect 5355 2109 5389 2143
rect 5355 2041 5389 2075
rect 5355 1973 5389 2007
rect -4849 1811 -4815 1845
rect -4781 1811 -4747 1845
rect -4713 1811 -4679 1845
rect -4645 1811 -4611 1845
rect -4577 1811 -4543 1845
rect -4509 1811 -4475 1845
rect -4441 1811 -4407 1845
rect -4373 1811 -4339 1845
rect -4305 1811 -4271 1845
rect -4237 1811 -4203 1845
rect -4169 1811 -4135 1845
rect -4101 1811 -4067 1845
rect -4033 1811 -3999 1845
rect -3965 1811 -3931 1845
rect -3897 1811 -3863 1845
rect -3829 1811 -3795 1845
rect -3761 1811 -3727 1845
rect -3693 1811 -3659 1845
rect -3625 1811 -3591 1845
rect -3557 1811 -3523 1845
rect -3489 1811 -3455 1845
rect -3421 1811 -3387 1845
rect -3353 1811 -3319 1845
rect -3285 1811 -3251 1845
rect -3217 1811 -3183 1845
rect -3149 1811 -3115 1845
rect -3081 1811 -3047 1845
rect -3013 1811 -2979 1845
rect -2945 1811 -2911 1845
rect -2877 1811 -2843 1845
rect -2809 1811 -2775 1845
rect -2741 1811 -2707 1845
rect -2673 1811 -2639 1845
rect -2605 1811 -2571 1845
rect -2537 1811 -2503 1845
rect -2469 1811 -2435 1845
rect -2401 1811 -2367 1845
rect -2333 1811 -2299 1845
rect -2265 1811 -2231 1845
rect -2197 1811 -2163 1845
rect -2129 1811 -2095 1845
rect -2061 1811 -2027 1845
rect -1993 1811 -1959 1845
rect -1925 1811 -1891 1845
rect -1857 1811 -1823 1845
rect -1789 1811 -1755 1845
rect -1721 1811 -1687 1845
rect -1653 1811 -1619 1845
rect -1585 1811 -1551 1845
rect -1517 1811 -1483 1845
rect -1449 1811 -1415 1845
rect -1381 1811 -1347 1845
rect -1313 1811 -1279 1845
rect -1245 1811 -1211 1845
rect -1177 1811 -1143 1845
rect -1109 1811 -1075 1845
rect -1041 1811 -1007 1845
rect -973 1811 -939 1845
rect -905 1811 -871 1845
rect -837 1811 -803 1845
rect -769 1811 -735 1845
rect -701 1811 -667 1845
rect -633 1811 -599 1845
rect -565 1811 -531 1845
rect -497 1811 -463 1845
rect -429 1811 -395 1845
rect -361 1811 -327 1845
rect -293 1811 -259 1845
rect -225 1811 -191 1845
rect -157 1811 -123 1845
rect -89 1811 -55 1845
rect -21 1811 13 1845
rect 47 1811 81 1845
rect 115 1811 149 1845
rect 183 1811 217 1845
rect 251 1811 285 1845
rect 319 1811 353 1845
rect 387 1811 421 1845
rect 455 1811 489 1845
rect 523 1811 557 1845
rect 591 1811 625 1845
rect 659 1811 693 1845
rect 727 1811 761 1845
rect 795 1811 829 1845
rect 863 1811 897 1845
rect 931 1811 965 1845
rect 999 1811 1033 1845
rect 1067 1811 1101 1845
rect 1135 1811 1169 1845
rect 1203 1811 1237 1845
rect 1271 1811 1305 1845
rect 1339 1811 1373 1845
rect 1407 1811 1441 1845
rect 1475 1811 1509 1845
rect 1543 1811 1577 1845
rect 1611 1811 1645 1845
rect 1679 1811 1713 1845
rect 1747 1811 1781 1845
rect 1815 1811 1849 1845
rect 1883 1811 1917 1845
rect 1951 1811 1985 1845
rect 2019 1811 2053 1845
rect 2087 1811 2121 1845
rect 2155 1811 2189 1845
rect 2223 1811 2257 1845
rect 2291 1811 2325 1845
rect 2359 1811 2393 1845
rect 2427 1811 2461 1845
rect 2495 1811 2529 1845
rect 2563 1811 2597 1845
rect 2631 1811 2665 1845
rect 2699 1811 2733 1845
rect 2767 1811 2801 1845
rect 2835 1811 2869 1845
rect 2903 1811 2937 1845
rect 2971 1811 3005 1845
rect 3039 1811 3073 1845
rect 3107 1811 3141 1845
rect 3175 1811 3209 1845
rect 3243 1811 3277 1845
rect 3311 1811 3345 1845
rect 3379 1811 3413 1845
rect 3447 1811 3481 1845
rect 3515 1811 3549 1845
rect 3583 1811 3617 1845
rect 3651 1811 3685 1845
rect 3719 1811 3753 1845
rect 3787 1811 3821 1845
rect 3855 1811 3889 1845
rect 3923 1811 3957 1845
rect 3991 1811 4025 1845
rect 4059 1811 4093 1845
rect 4127 1811 4161 1845
rect 4195 1811 4229 1845
rect 4263 1811 4297 1845
rect 4331 1811 4365 1845
rect 4399 1811 4433 1845
rect 4467 1811 4501 1845
rect 4535 1811 4569 1845
rect 4603 1811 4637 1845
rect 4671 1811 4705 1845
rect 4739 1811 4773 1845
rect 4807 1811 4841 1845
rect 4875 1811 4909 1845
rect 4943 1811 4977 1845
rect 5011 1811 5045 1845
rect 5079 1811 5113 1845
rect 5147 1811 5181 1845
rect 5215 1811 5249 1845
<< nsubdiffcont >>
rect -4849 10255 -4815 10289
rect -4781 10255 -4747 10289
rect -4713 10255 -4679 10289
rect -4645 10255 -4611 10289
rect -4577 10255 -4543 10289
rect -4509 10255 -4475 10289
rect -4441 10255 -4407 10289
rect -4373 10255 -4339 10289
rect -4305 10255 -4271 10289
rect -4237 10255 -4203 10289
rect -4169 10255 -4135 10289
rect -4101 10255 -4067 10289
rect -4033 10255 -3999 10289
rect -3965 10255 -3931 10289
rect -3897 10255 -3863 10289
rect -3829 10255 -3795 10289
rect -3761 10255 -3727 10289
rect -3693 10255 -3659 10289
rect -3625 10255 -3591 10289
rect -3557 10255 -3523 10289
rect -3489 10255 -3455 10289
rect -3421 10255 -3387 10289
rect -3353 10255 -3319 10289
rect -3285 10255 -3251 10289
rect -3217 10255 -3183 10289
rect -3149 10255 -3115 10289
rect -3081 10255 -3047 10289
rect -3013 10255 -2979 10289
rect -2945 10255 -2911 10289
rect -2877 10255 -2843 10289
rect -2809 10255 -2775 10289
rect -2741 10255 -2707 10289
rect -2673 10255 -2639 10289
rect -2605 10255 -2571 10289
rect -2537 10255 -2503 10289
rect -2469 10255 -2435 10289
rect -2401 10255 -2367 10289
rect -2333 10255 -2299 10289
rect -2265 10255 -2231 10289
rect -2197 10255 -2163 10289
rect -2129 10255 -2095 10289
rect -2061 10255 -2027 10289
rect -1993 10255 -1959 10289
rect -1925 10255 -1891 10289
rect -1857 10255 -1823 10289
rect -1789 10255 -1755 10289
rect -1721 10255 -1687 10289
rect -1653 10255 -1619 10289
rect -1585 10255 -1551 10289
rect -1517 10255 -1483 10289
rect -1449 10255 -1415 10289
rect -1381 10255 -1347 10289
rect -1313 10255 -1279 10289
rect -1245 10255 -1211 10289
rect -1177 10255 -1143 10289
rect -1109 10255 -1075 10289
rect -1041 10255 -1007 10289
rect -973 10255 -939 10289
rect -905 10255 -871 10289
rect -837 10255 -803 10289
rect -769 10255 -735 10289
rect -701 10255 -667 10289
rect -633 10255 -599 10289
rect -565 10255 -531 10289
rect -497 10255 -463 10289
rect -429 10255 -395 10289
rect -361 10255 -327 10289
rect -293 10255 -259 10289
rect -225 10255 -191 10289
rect -157 10255 -123 10289
rect -89 10255 -55 10289
rect -21 10255 13 10289
rect 47 10255 81 10289
rect 115 10255 149 10289
rect 183 10255 217 10289
rect 251 10255 285 10289
rect 319 10255 353 10289
rect 387 10255 421 10289
rect 455 10255 489 10289
rect 523 10255 557 10289
rect 591 10255 625 10289
rect 659 10255 693 10289
rect 727 10255 761 10289
rect 795 10255 829 10289
rect 863 10255 897 10289
rect 931 10255 965 10289
rect 999 10255 1033 10289
rect 1067 10255 1101 10289
rect 1135 10255 1169 10289
rect 1203 10255 1237 10289
rect 1271 10255 1305 10289
rect 1339 10255 1373 10289
rect 1407 10255 1441 10289
rect 1475 10255 1509 10289
rect 1543 10255 1577 10289
rect 1611 10255 1645 10289
rect 1679 10255 1713 10289
rect 1747 10255 1781 10289
rect 1815 10255 1849 10289
rect 1883 10255 1917 10289
rect 1951 10255 1985 10289
rect 2019 10255 2053 10289
rect 2087 10255 2121 10289
rect 2155 10255 2189 10289
rect 2223 10255 2257 10289
rect 2291 10255 2325 10289
rect 2359 10255 2393 10289
rect 2427 10255 2461 10289
rect 2495 10255 2529 10289
rect 2563 10255 2597 10289
rect 2631 10255 2665 10289
rect 2699 10255 2733 10289
rect 2767 10255 2801 10289
rect 2835 10255 2869 10289
rect 2903 10255 2937 10289
rect 2971 10255 3005 10289
rect 3039 10255 3073 10289
rect 3107 10255 3141 10289
rect 3175 10255 3209 10289
rect 3243 10255 3277 10289
rect 3311 10255 3345 10289
rect 3379 10255 3413 10289
rect 3447 10255 3481 10289
rect 3515 10255 3549 10289
rect 3583 10255 3617 10289
rect 3651 10255 3685 10289
rect 3719 10255 3753 10289
rect 3787 10255 3821 10289
rect 3855 10255 3889 10289
rect 3923 10255 3957 10289
rect 3991 10255 4025 10289
rect 4059 10255 4093 10289
rect 4127 10255 4161 10289
rect 4195 10255 4229 10289
rect 4263 10255 4297 10289
rect 4331 10255 4365 10289
rect 4399 10255 4433 10289
rect 4467 10255 4501 10289
rect 4535 10255 4569 10289
rect 4603 10255 4637 10289
rect 4671 10255 4705 10289
rect 4739 10255 4773 10289
rect 4807 10255 4841 10289
rect 4875 10255 4909 10289
rect 4943 10255 4977 10289
rect 5011 10255 5045 10289
rect 5079 10255 5113 10289
rect 5147 10255 5181 10289
rect 5215 10255 5249 10289
rect -4989 10103 -4955 10137
rect -4989 10035 -4955 10069
rect -4989 9967 -4955 10001
rect -4989 9899 -4955 9933
rect -4989 9831 -4955 9865
rect -4989 9763 -4955 9797
rect -4989 9695 -4955 9729
rect -4989 9627 -4955 9661
rect -4989 9559 -4955 9593
rect -4989 9491 -4955 9525
rect -4989 9423 -4955 9457
rect -4989 9355 -4955 9389
rect -4989 9287 -4955 9321
rect -4989 9219 -4955 9253
rect -4989 9151 -4955 9185
rect -4989 9083 -4955 9117
rect -4989 9015 -4955 9049
rect -4989 8947 -4955 8981
rect -4989 8879 -4955 8913
rect -4989 8811 -4955 8845
rect -4989 8743 -4955 8777
rect -4989 8675 -4955 8709
rect -4989 8607 -4955 8641
rect -4989 8539 -4955 8573
rect -4989 8471 -4955 8505
rect -4989 8403 -4955 8437
rect -4989 8335 -4955 8369
rect -4989 8267 -4955 8301
rect -4989 8199 -4955 8233
rect -4989 8131 -4955 8165
rect -4989 8063 -4955 8097
rect -4989 7995 -4955 8029
rect -4989 7927 -4955 7961
rect -4989 7859 -4955 7893
rect -4989 7791 -4955 7825
rect -4989 7723 -4955 7757
rect -4989 7655 -4955 7689
rect -4989 7587 -4955 7621
rect -4989 7519 -4955 7553
rect -4989 7451 -4955 7485
rect -4989 7383 -4955 7417
rect -4989 7315 -4955 7349
rect -4989 7247 -4955 7281
rect -4989 7179 -4955 7213
rect -4989 7111 -4955 7145
rect -4989 7043 -4955 7077
rect -4989 6975 -4955 7009
rect -4989 6907 -4955 6941
rect -4989 6839 -4955 6873
rect -4989 6771 -4955 6805
rect -4989 6703 -4955 6737
rect -4989 6635 -4955 6669
rect -4989 6567 -4955 6601
rect -4989 6499 -4955 6533
rect -4989 6431 -4955 6465
rect -4989 6363 -4955 6397
rect -4989 6295 -4955 6329
rect -4989 6227 -4955 6261
rect -4989 6159 -4955 6193
rect -4989 6091 -4955 6125
rect -4989 6023 -4955 6057
rect -4989 5955 -4955 5989
rect -4989 5887 -4955 5921
rect -4989 5819 -4955 5853
rect -4989 5751 -4955 5785
rect -4989 5683 -4955 5717
rect -4989 5615 -4955 5649
rect -4989 5547 -4955 5581
rect -4989 5479 -4955 5513
rect -4989 5411 -4955 5445
rect -4989 5343 -4955 5377
rect -4989 5275 -4955 5309
rect -4989 5207 -4955 5241
rect -4989 5139 -4955 5173
rect -4989 5071 -4955 5105
rect -4989 5003 -4955 5037
rect -4989 4935 -4955 4969
rect -4989 4867 -4955 4901
rect -4989 4799 -4955 4833
rect -4989 4731 -4955 4765
rect -4989 4663 -4955 4697
rect 5355 10103 5389 10137
rect 5355 10035 5389 10069
rect 5355 9967 5389 10001
rect 5355 9899 5389 9933
rect 5355 9831 5389 9865
rect 5355 9763 5389 9797
rect 5355 9695 5389 9729
rect 5355 9627 5389 9661
rect 5355 9559 5389 9593
rect 5355 9491 5389 9525
rect 5355 9423 5389 9457
rect 5355 9355 5389 9389
rect 5355 9287 5389 9321
rect 5355 9219 5389 9253
rect 5355 9151 5389 9185
rect 5355 9083 5389 9117
rect 5355 9015 5389 9049
rect 5355 8947 5389 8981
rect 5355 8879 5389 8913
rect 5355 8811 5389 8845
rect 5355 8743 5389 8777
rect 5355 8675 5389 8709
rect 5355 8607 5389 8641
rect 5355 8539 5389 8573
rect 5355 8471 5389 8505
rect 5355 8403 5389 8437
rect 5355 8335 5389 8369
rect 5355 8267 5389 8301
rect 5355 8199 5389 8233
rect 5355 8131 5389 8165
rect 5355 8063 5389 8097
rect 5355 7995 5389 8029
rect 5355 7927 5389 7961
rect 5355 7859 5389 7893
rect 5355 7791 5389 7825
rect 5355 7723 5389 7757
rect 5355 7655 5389 7689
rect 5355 7587 5389 7621
rect 5355 7519 5389 7553
rect 5355 7451 5389 7485
rect 5355 7383 5389 7417
rect 5355 7315 5389 7349
rect 5355 7247 5389 7281
rect 5355 7179 5389 7213
rect 5355 7111 5389 7145
rect 5355 7043 5389 7077
rect 5355 6975 5389 7009
rect 5355 6907 5389 6941
rect 5355 6839 5389 6873
rect 5355 6771 5389 6805
rect 5355 6703 5389 6737
rect 5355 6635 5389 6669
rect 5355 6567 5389 6601
rect 5355 6499 5389 6533
rect 5355 6431 5389 6465
rect 5355 6363 5389 6397
rect 5355 6295 5389 6329
rect 5355 6227 5389 6261
rect 5355 6159 5389 6193
rect 5355 6091 5389 6125
rect 5355 6023 5389 6057
rect 5355 5955 5389 5989
rect 5355 5887 5389 5921
rect 5355 5819 5389 5853
rect 5355 5751 5389 5785
rect 5355 5683 5389 5717
rect 5355 5615 5389 5649
rect 5355 5547 5389 5581
rect 5355 5479 5389 5513
rect 5355 5411 5389 5445
rect 5355 5343 5389 5377
rect 5355 5275 5389 5309
rect 5355 5207 5389 5241
rect 5355 5139 5389 5173
rect 5355 5071 5389 5105
rect 5355 5003 5389 5037
rect 5355 4935 5389 4969
rect 5355 4867 5389 4901
rect 5355 4799 5389 4833
rect 5355 4731 5389 4765
rect 5355 4663 5389 4697
rect -4849 4511 -4815 4545
rect -4781 4511 -4747 4545
rect -4713 4511 -4679 4545
rect -4645 4511 -4611 4545
rect -4577 4511 -4543 4545
rect -4509 4511 -4475 4545
rect -4441 4511 -4407 4545
rect -4373 4511 -4339 4545
rect -4305 4511 -4271 4545
rect -4237 4511 -4203 4545
rect -4169 4511 -4135 4545
rect -4101 4511 -4067 4545
rect -4033 4511 -3999 4545
rect -3965 4511 -3931 4545
rect -3897 4511 -3863 4545
rect -3829 4511 -3795 4545
rect -3761 4511 -3727 4545
rect -3693 4511 -3659 4545
rect -3625 4511 -3591 4545
rect -3557 4511 -3523 4545
rect -3489 4511 -3455 4545
rect -3421 4511 -3387 4545
rect -3353 4511 -3319 4545
rect -3285 4511 -3251 4545
rect -3217 4511 -3183 4545
rect -3149 4511 -3115 4545
rect -3081 4511 -3047 4545
rect -3013 4511 -2979 4545
rect -2945 4511 -2911 4545
rect -2877 4511 -2843 4545
rect -2809 4511 -2775 4545
rect -2741 4511 -2707 4545
rect -2673 4511 -2639 4545
rect -2605 4511 -2571 4545
rect -2537 4511 -2503 4545
rect -2469 4511 -2435 4545
rect -2401 4511 -2367 4545
rect -2333 4511 -2299 4545
rect -2265 4511 -2231 4545
rect -2197 4511 -2163 4545
rect -2129 4511 -2095 4545
rect -2061 4511 -2027 4545
rect -1993 4511 -1959 4545
rect -1925 4511 -1891 4545
rect -1857 4511 -1823 4545
rect -1789 4511 -1755 4545
rect -1721 4511 -1687 4545
rect -1653 4511 -1619 4545
rect -1585 4511 -1551 4545
rect -1517 4511 -1483 4545
rect -1449 4511 -1415 4545
rect -1381 4511 -1347 4545
rect -1313 4511 -1279 4545
rect -1245 4511 -1211 4545
rect -1177 4511 -1143 4545
rect -1109 4511 -1075 4545
rect -1041 4511 -1007 4545
rect -973 4511 -939 4545
rect -905 4511 -871 4545
rect -837 4511 -803 4545
rect -769 4511 -735 4545
rect -701 4511 -667 4545
rect -633 4511 -599 4545
rect -565 4511 -531 4545
rect -497 4511 -463 4545
rect -429 4511 -395 4545
rect -361 4511 -327 4545
rect -293 4511 -259 4545
rect -225 4511 -191 4545
rect -157 4511 -123 4545
rect -89 4511 -55 4545
rect -21 4511 13 4545
rect 47 4511 81 4545
rect 115 4511 149 4545
rect 183 4511 217 4545
rect 251 4511 285 4545
rect 319 4511 353 4545
rect 387 4511 421 4545
rect 455 4511 489 4545
rect 523 4511 557 4545
rect 591 4511 625 4545
rect 659 4511 693 4545
rect 727 4511 761 4545
rect 795 4511 829 4545
rect 863 4511 897 4545
rect 931 4511 965 4545
rect 999 4511 1033 4545
rect 1067 4511 1101 4545
rect 1135 4511 1169 4545
rect 1203 4511 1237 4545
rect 1271 4511 1305 4545
rect 1339 4511 1373 4545
rect 1407 4511 1441 4545
rect 1475 4511 1509 4545
rect 1543 4511 1577 4545
rect 1611 4511 1645 4545
rect 1679 4511 1713 4545
rect 1747 4511 1781 4545
rect 1815 4511 1849 4545
rect 1883 4511 1917 4545
rect 1951 4511 1985 4545
rect 2019 4511 2053 4545
rect 2087 4511 2121 4545
rect 2155 4511 2189 4545
rect 2223 4511 2257 4545
rect 2291 4511 2325 4545
rect 2359 4511 2393 4545
rect 2427 4511 2461 4545
rect 2495 4511 2529 4545
rect 2563 4511 2597 4545
rect 2631 4511 2665 4545
rect 2699 4511 2733 4545
rect 2767 4511 2801 4545
rect 2835 4511 2869 4545
rect 2903 4511 2937 4545
rect 2971 4511 3005 4545
rect 3039 4511 3073 4545
rect 3107 4511 3141 4545
rect 3175 4511 3209 4545
rect 3243 4511 3277 4545
rect 3311 4511 3345 4545
rect 3379 4511 3413 4545
rect 3447 4511 3481 4545
rect 3515 4511 3549 4545
rect 3583 4511 3617 4545
rect 3651 4511 3685 4545
rect 3719 4511 3753 4545
rect 3787 4511 3821 4545
rect 3855 4511 3889 4545
rect 3923 4511 3957 4545
rect 3991 4511 4025 4545
rect 4059 4511 4093 4545
rect 4127 4511 4161 4545
rect 4195 4511 4229 4545
rect 4263 4511 4297 4545
rect 4331 4511 4365 4545
rect 4399 4511 4433 4545
rect 4467 4511 4501 4545
rect 4535 4511 4569 4545
rect 4603 4511 4637 4545
rect 4671 4511 4705 4545
rect 4739 4511 4773 4545
rect 4807 4511 4841 4545
rect 4875 4511 4909 4545
rect 4943 4511 4977 4545
rect 5011 4511 5045 4545
rect 5079 4511 5113 4545
rect 5147 4511 5181 4545
rect 5215 4511 5249 4545
<< locali >>
rect -5022 10289 5422 10322
rect -5022 10255 -4893 10289
rect -4859 10255 -4849 10289
rect -4787 10255 -4781 10289
rect -4715 10255 -4713 10289
rect -4679 10255 -4677 10289
rect -4611 10255 -4605 10289
rect -4543 10255 -4533 10289
rect -4475 10255 -4461 10289
rect -4407 10255 -4389 10289
rect -4339 10255 -4317 10289
rect -4271 10255 -4245 10289
rect -4203 10255 -4173 10289
rect -4135 10255 -4101 10289
rect -4067 10255 -4033 10289
rect -3995 10255 -3965 10289
rect -3923 10255 -3897 10289
rect -3851 10255 -3829 10289
rect -3779 10255 -3761 10289
rect -3707 10255 -3693 10289
rect -3635 10255 -3625 10289
rect -3563 10255 -3557 10289
rect -3491 10255 -3489 10289
rect -3455 10255 -3453 10289
rect -3387 10255 -3381 10289
rect -3319 10255 -3309 10289
rect -3251 10255 -3237 10289
rect -3183 10255 -3165 10289
rect -3115 10255 -3093 10289
rect -3047 10255 -3021 10289
rect -2979 10255 -2949 10289
rect -2911 10255 -2877 10289
rect -2843 10255 -2809 10289
rect -2771 10255 -2741 10289
rect -2699 10255 -2673 10289
rect -2627 10255 -2605 10289
rect -2555 10255 -2537 10289
rect -2483 10255 -2469 10289
rect -2411 10255 -2401 10289
rect -2339 10255 -2333 10289
rect -2267 10255 -2265 10289
rect -2231 10255 -2229 10289
rect -2163 10255 -2157 10289
rect -2095 10255 -2085 10289
rect -2027 10255 -2013 10289
rect -1959 10255 -1941 10289
rect -1891 10255 -1869 10289
rect -1823 10255 -1797 10289
rect -1755 10255 -1725 10289
rect -1687 10255 -1653 10289
rect -1619 10255 -1585 10289
rect -1547 10255 -1517 10289
rect -1475 10255 -1449 10289
rect -1403 10255 -1381 10289
rect -1331 10255 -1313 10289
rect -1259 10255 -1245 10289
rect -1187 10255 -1177 10289
rect -1115 10255 -1109 10289
rect -1043 10255 -1041 10289
rect -1007 10255 -1005 10289
rect -939 10255 -933 10289
rect -871 10255 -861 10289
rect -803 10255 -789 10289
rect -735 10255 -717 10289
rect -667 10255 -645 10289
rect -599 10255 -573 10289
rect -531 10255 -501 10289
rect -463 10255 -429 10289
rect -395 10255 -361 10289
rect -323 10255 -293 10289
rect -251 10255 -225 10289
rect -179 10255 -157 10289
rect -107 10255 -89 10289
rect -35 10255 -21 10289
rect 37 10255 47 10289
rect 109 10255 115 10289
rect 181 10255 183 10289
rect 217 10255 219 10289
rect 285 10255 291 10289
rect 353 10255 363 10289
rect 421 10255 435 10289
rect 489 10255 507 10289
rect 557 10255 579 10289
rect 625 10255 651 10289
rect 693 10255 723 10289
rect 761 10255 795 10289
rect 829 10255 863 10289
rect 901 10255 931 10289
rect 973 10255 999 10289
rect 1045 10255 1067 10289
rect 1117 10255 1135 10289
rect 1189 10255 1203 10289
rect 1261 10255 1271 10289
rect 1333 10255 1339 10289
rect 1405 10255 1407 10289
rect 1441 10255 1443 10289
rect 1509 10255 1515 10289
rect 1577 10255 1587 10289
rect 1645 10255 1659 10289
rect 1713 10255 1731 10289
rect 1781 10255 1803 10289
rect 1849 10255 1875 10289
rect 1917 10255 1947 10289
rect 1985 10255 2019 10289
rect 2053 10255 2087 10289
rect 2125 10255 2155 10289
rect 2197 10255 2223 10289
rect 2269 10255 2291 10289
rect 2341 10255 2359 10289
rect 2413 10255 2427 10289
rect 2485 10255 2495 10289
rect 2557 10255 2563 10289
rect 2629 10255 2631 10289
rect 2665 10255 2667 10289
rect 2733 10255 2739 10289
rect 2801 10255 2811 10289
rect 2869 10255 2883 10289
rect 2937 10255 2955 10289
rect 3005 10255 3027 10289
rect 3073 10255 3099 10289
rect 3141 10255 3171 10289
rect 3209 10255 3243 10289
rect 3277 10255 3311 10289
rect 3349 10255 3379 10289
rect 3421 10255 3447 10289
rect 3493 10255 3515 10289
rect 3565 10255 3583 10289
rect 3637 10255 3651 10289
rect 3709 10255 3719 10289
rect 3781 10255 3787 10289
rect 3853 10255 3855 10289
rect 3889 10255 3891 10289
rect 3957 10255 3963 10289
rect 4025 10255 4035 10289
rect 4093 10255 4107 10289
rect 4161 10255 4179 10289
rect 4229 10255 4251 10289
rect 4297 10255 4323 10289
rect 4365 10255 4395 10289
rect 4433 10255 4467 10289
rect 4501 10255 4535 10289
rect 4573 10255 4603 10289
rect 4645 10255 4671 10289
rect 4717 10255 4739 10289
rect 4789 10255 4807 10289
rect 4861 10255 4875 10289
rect 4933 10255 4943 10289
rect 5005 10255 5011 10289
rect 5077 10255 5079 10289
rect 5113 10255 5115 10289
rect 5181 10255 5187 10289
rect 5249 10255 5259 10289
rect 5293 10255 5422 10289
rect -5022 10222 5422 10255
rect -5022 10137 -4922 10222
rect -5022 10103 -4989 10137
rect -4955 10103 -4922 10137
rect -5022 10069 -4922 10103
rect -5022 10035 -4989 10069
rect -4955 10035 -4922 10069
rect -5022 10001 -4922 10035
rect -5022 9967 -4989 10001
rect -4955 9967 -4922 10001
rect -5022 9933 -4922 9967
rect -5022 9885 -4989 9933
rect -4955 9885 -4922 9933
rect -5022 9865 -4922 9885
rect -5022 9813 -4989 9865
rect -4955 9813 -4922 9865
rect -5022 9797 -4922 9813
rect -5022 9741 -4989 9797
rect -4955 9741 -4922 9797
rect -5022 9729 -4922 9741
rect -5022 9669 -4989 9729
rect -4955 9669 -4922 9729
rect -5022 9661 -4922 9669
rect -5022 9597 -4989 9661
rect -4955 9597 -4922 9661
rect -5022 9593 -4922 9597
rect -5022 9491 -4989 9593
rect -4955 9491 -4922 9593
rect -5022 9487 -4922 9491
rect -5022 9423 -4989 9487
rect -4955 9423 -4922 9487
rect -5022 9415 -4922 9423
rect -5022 9355 -4989 9415
rect -4955 9355 -4922 9415
rect -5022 9343 -4922 9355
rect -5022 9287 -4989 9343
rect -4955 9287 -4922 9343
rect -5022 9271 -4922 9287
rect -5022 9219 -4989 9271
rect -4955 9219 -4922 9271
rect -5022 9199 -4922 9219
rect -5022 9151 -4989 9199
rect -4955 9151 -4922 9199
rect -5022 9127 -4922 9151
rect -5022 9083 -4989 9127
rect -4955 9083 -4922 9127
rect -5022 9055 -4922 9083
rect -5022 9015 -4989 9055
rect -4955 9015 -4922 9055
rect -5022 8983 -4922 9015
rect -5022 8947 -4989 8983
rect -4955 8947 -4922 8983
rect -5022 8913 -4922 8947
rect -5022 8877 -4989 8913
rect -4955 8877 -4922 8913
rect -5022 8845 -4922 8877
rect -5022 8805 -4989 8845
rect -4955 8805 -4922 8845
rect -5022 8777 -4922 8805
rect -5022 8733 -4989 8777
rect -4955 8733 -4922 8777
rect -5022 8709 -4922 8733
rect -5022 8661 -4989 8709
rect -4955 8661 -4922 8709
rect -5022 8641 -4922 8661
rect -5022 8589 -4989 8641
rect -4955 8589 -4922 8641
rect -5022 8573 -4922 8589
rect -5022 8517 -4989 8573
rect -4955 8517 -4922 8573
rect -5022 8505 -4922 8517
rect -5022 8445 -4989 8505
rect -4955 8445 -4922 8505
rect -5022 8437 -4922 8445
rect -5022 8373 -4989 8437
rect -4955 8373 -4922 8437
rect -5022 8369 -4922 8373
rect -5022 8267 -4989 8369
rect -4955 8267 -4922 8369
rect -5022 8263 -4922 8267
rect -5022 8199 -4989 8263
rect -4955 8199 -4922 8263
rect -5022 8191 -4922 8199
rect -5022 8131 -4989 8191
rect -4955 8131 -4922 8191
rect -5022 8119 -4922 8131
rect -5022 8063 -4989 8119
rect -4955 8063 -4922 8119
rect -5022 8047 -4922 8063
rect -5022 7995 -4989 8047
rect -4955 7995 -4922 8047
rect -5022 7975 -4922 7995
rect -5022 7927 -4989 7975
rect -4955 7927 -4922 7975
rect -5022 7903 -4922 7927
rect -5022 7859 -4989 7903
rect -4955 7859 -4922 7903
rect -5022 7831 -4922 7859
rect -5022 7791 -4989 7831
rect -4955 7791 -4922 7831
rect -5022 7759 -4922 7791
rect -5022 7723 -4989 7759
rect -4955 7723 -4922 7759
rect -5022 7689 -4922 7723
rect -5022 7653 -4989 7689
rect -4955 7653 -4922 7689
rect -5022 7621 -4922 7653
rect -5022 7581 -4989 7621
rect -4955 7581 -4922 7621
rect -5022 7553 -4922 7581
rect -5022 7509 -4989 7553
rect -4955 7509 -4922 7553
rect -5022 7485 -4922 7509
rect -5022 7437 -4989 7485
rect -4955 7437 -4922 7485
rect -5022 7417 -4922 7437
rect -5022 7365 -4989 7417
rect -4955 7365 -4922 7417
rect -5022 7349 -4922 7365
rect -5022 7293 -4989 7349
rect -4955 7293 -4922 7349
rect -5022 7281 -4922 7293
rect -5022 7221 -4989 7281
rect -4955 7221 -4922 7281
rect -5022 7213 -4922 7221
rect -5022 7149 -4989 7213
rect -4955 7149 -4922 7213
rect -5022 7145 -4922 7149
rect -5022 7043 -4989 7145
rect -4955 7043 -4922 7145
rect 5322 10137 5422 10222
rect 5322 10103 5355 10137
rect 5389 10103 5422 10137
rect 5322 10069 5422 10103
rect 5322 10035 5355 10069
rect 5389 10035 5422 10069
rect 5322 10001 5422 10035
rect 5322 9967 5355 10001
rect 5389 9967 5422 10001
rect 5322 9933 5422 9967
rect 5322 9885 5355 9933
rect 5389 9885 5422 9933
rect 5322 9865 5422 9885
rect 5322 9813 5355 9865
rect 5389 9813 5422 9865
rect 5322 9797 5422 9813
rect 5322 9741 5355 9797
rect 5389 9741 5422 9797
rect 5322 9729 5422 9741
rect 5322 9669 5355 9729
rect 5389 9669 5422 9729
rect 5322 9661 5422 9669
rect 5322 9597 5355 9661
rect 5389 9597 5422 9661
rect 5322 9593 5422 9597
rect 5322 9491 5355 9593
rect 5389 9491 5422 9593
rect 5322 9487 5422 9491
rect 5322 9423 5355 9487
rect 5389 9423 5422 9487
rect 5322 9415 5422 9423
rect 5322 9355 5355 9415
rect 5389 9355 5422 9415
rect 5322 9343 5422 9355
rect 5322 9287 5355 9343
rect 5389 9287 5422 9343
rect 5322 9271 5422 9287
rect 5322 9219 5355 9271
rect 5389 9219 5422 9271
rect 5322 9199 5422 9219
rect 5322 9151 5355 9199
rect 5389 9151 5422 9199
rect 5322 9127 5422 9151
rect 5322 9083 5355 9127
rect 5389 9083 5422 9127
rect 5322 9055 5422 9083
rect 5322 9015 5355 9055
rect 5389 9015 5422 9055
rect 5322 8983 5422 9015
rect 5322 8947 5355 8983
rect 5389 8947 5422 8983
rect 5322 8913 5422 8947
rect 5322 8877 5355 8913
rect 5389 8877 5422 8913
rect 5322 8845 5422 8877
rect 5322 8805 5355 8845
rect 5389 8805 5422 8845
rect 5322 8777 5422 8805
rect 5322 8733 5355 8777
rect 5389 8733 5422 8777
rect 5322 8709 5422 8733
rect 5322 8661 5355 8709
rect 5389 8661 5422 8709
rect 5322 8641 5422 8661
rect 5322 8589 5355 8641
rect 5389 8589 5422 8641
rect 5322 8573 5422 8589
rect 5322 8517 5355 8573
rect 5389 8517 5422 8573
rect 5322 8505 5422 8517
rect 5322 8445 5355 8505
rect 5389 8445 5422 8505
rect 5322 8437 5422 8445
rect 5322 8373 5355 8437
rect 5389 8373 5422 8437
rect 5322 8369 5422 8373
rect 5322 8267 5355 8369
rect 5389 8267 5422 8369
rect 5322 8263 5422 8267
rect 5322 8199 5355 8263
rect 5389 8199 5422 8263
rect 5322 8191 5422 8199
rect 5322 8131 5355 8191
rect 5389 8131 5422 8191
rect 5322 8119 5422 8131
rect 5322 8063 5355 8119
rect 5389 8063 5422 8119
rect 5322 8047 5422 8063
rect 5322 7995 5355 8047
rect 5389 7995 5422 8047
rect 5322 7975 5422 7995
rect 5322 7927 5355 7975
rect 5389 7927 5422 7975
rect 5322 7903 5422 7927
rect 5322 7859 5355 7903
rect 5389 7859 5422 7903
rect 5322 7831 5422 7859
rect 5322 7791 5355 7831
rect 5389 7791 5422 7831
rect 5322 7759 5422 7791
rect 5322 7723 5355 7759
rect 5389 7723 5422 7759
rect 5322 7689 5422 7723
rect 5322 7653 5355 7689
rect 5389 7653 5422 7689
rect 5322 7621 5422 7653
rect 5322 7581 5355 7621
rect 5389 7581 5422 7621
rect 5322 7553 5422 7581
rect 5322 7509 5355 7553
rect 5389 7509 5422 7553
rect 5322 7485 5422 7509
rect 5322 7437 5355 7485
rect 5389 7437 5422 7485
rect 5322 7417 5422 7437
rect 5322 7365 5355 7417
rect 5389 7365 5422 7417
rect 5322 7349 5422 7365
rect 5322 7293 5355 7349
rect 5389 7293 5422 7349
rect 5322 7281 5422 7293
rect 5322 7221 5355 7281
rect 5389 7221 5422 7281
rect 5322 7213 5422 7221
rect 5322 7149 5355 7213
rect 5389 7149 5422 7213
rect 5322 7145 5422 7149
rect -158 7099 362 7112
rect -158 7065 -145 7099
rect -111 7065 315 7099
rect 349 7065 362 7099
rect -158 7052 362 7065
rect -5022 7039 -4922 7043
rect -5022 6975 -4989 7039
rect -4955 6975 -4922 7039
rect -5022 6967 -4922 6975
rect -5022 6907 -4989 6967
rect -4955 6907 -4922 6967
rect -5022 6895 -4922 6907
rect -5022 6839 -4989 6895
rect -4955 6839 -4922 6895
rect -5022 6823 -4922 6839
rect -5022 6771 -4989 6823
rect -4955 6771 -4922 6823
rect -5022 6751 -4922 6771
rect -5022 6703 -4989 6751
rect -4955 6703 -4922 6751
rect -5022 6679 -4922 6703
rect -5022 6635 -4989 6679
rect -4955 6635 -4922 6679
rect -5022 6607 -4922 6635
rect -5022 6567 -4989 6607
rect -4955 6567 -4922 6607
rect -5022 6535 -4922 6567
rect -5022 6499 -4989 6535
rect -4955 6499 -4922 6535
rect -5022 6465 -4922 6499
rect -5022 6429 -4989 6465
rect -4955 6429 -4922 6465
rect -5022 6397 -4922 6429
rect -5022 6357 -4989 6397
rect -4955 6357 -4922 6397
rect -5022 6329 -4922 6357
rect -5022 6285 -4989 6329
rect -4955 6285 -4922 6329
rect -5022 6261 -4922 6285
rect -5022 6213 -4989 6261
rect -4955 6213 -4922 6261
rect -5022 6193 -4922 6213
rect -5022 6141 -4989 6193
rect -4955 6141 -4922 6193
rect -5022 6125 -4922 6141
rect -5022 6069 -4989 6125
rect -4955 6069 -4922 6125
rect -5022 6057 -4922 6069
rect -5022 5997 -4989 6057
rect -4955 5997 -4922 6057
rect -5022 5989 -4922 5997
rect -5022 5925 -4989 5989
rect -4955 5925 -4922 5989
rect -5022 5921 -4922 5925
rect -5022 5819 -4989 5921
rect -4955 5819 -4922 5921
rect -5022 5815 -4922 5819
rect -5022 5751 -4989 5815
rect -4955 5751 -4922 5815
rect -5022 5743 -4922 5751
rect -5022 5683 -4989 5743
rect -4955 5683 -4922 5743
rect -5022 5671 -4922 5683
rect -5022 5615 -4989 5671
rect -4955 5615 -4922 5671
rect -5022 5599 -4922 5615
rect -5022 5547 -4989 5599
rect -4955 5547 -4922 5599
rect -5022 5527 -4922 5547
rect -5022 5479 -4989 5527
rect -4955 5479 -4922 5527
rect -5022 5455 -4922 5479
rect -5022 5411 -4989 5455
rect -4955 5411 -4922 5455
rect -5022 5383 -4922 5411
rect -5022 5343 -4989 5383
rect -4955 5343 -4922 5383
rect -5022 5311 -4922 5343
rect -5022 5275 -4989 5311
rect -4955 5275 -4922 5311
rect -5022 5241 -4922 5275
rect -5022 5205 -4989 5241
rect -4955 5205 -4922 5241
rect -5022 5173 -4922 5205
rect -5022 5133 -4989 5173
rect -4955 5133 -4922 5173
rect -5022 5105 -4922 5133
rect -5022 5061 -4989 5105
rect -4955 5061 -4922 5105
rect -5022 5037 -4922 5061
rect -5022 4989 -4989 5037
rect -4955 4989 -4922 5037
rect -5022 4969 -4922 4989
rect -5022 4917 -4989 4969
rect -4955 4917 -4922 4969
rect -5022 4901 -4922 4917
rect -5022 4845 -4989 4901
rect -4955 4845 -4922 4901
rect -5022 4833 -4922 4845
rect -5022 4773 -4989 4833
rect -4955 4773 -4922 4833
rect -5022 4765 -4922 4773
rect -5022 4731 -4989 4765
rect -4955 4731 -4922 4765
rect -5022 4697 -4922 4731
rect -5022 4663 -4989 4697
rect -4955 4663 -4922 4697
rect -5022 4578 -4922 4663
rect 5322 7043 5355 7145
rect 5389 7043 5422 7145
rect 5322 7039 5422 7043
rect 5322 6975 5355 7039
rect 5389 6975 5422 7039
rect 5322 6967 5422 6975
rect 5322 6907 5355 6967
rect 5389 6907 5422 6967
rect 5322 6895 5422 6907
rect 5322 6839 5355 6895
rect 5389 6839 5422 6895
rect 5322 6823 5422 6839
rect 5322 6771 5355 6823
rect 5389 6771 5422 6823
rect 5322 6751 5422 6771
rect 5322 6703 5355 6751
rect 5389 6703 5422 6751
rect 5322 6679 5422 6703
rect 5322 6635 5355 6679
rect 5389 6635 5422 6679
rect 5322 6607 5422 6635
rect 5322 6567 5355 6607
rect 5389 6567 5422 6607
rect 5322 6535 5422 6567
rect 5322 6499 5355 6535
rect 5389 6499 5422 6535
rect 5322 6465 5422 6499
rect 5322 6429 5355 6465
rect 5389 6429 5422 6465
rect 5322 6397 5422 6429
rect 5322 6357 5355 6397
rect 5389 6357 5422 6397
rect 5322 6329 5422 6357
rect 5322 6285 5355 6329
rect 5389 6285 5422 6329
rect 5322 6261 5422 6285
rect 5322 6213 5355 6261
rect 5389 6213 5422 6261
rect 5322 6193 5422 6213
rect 5322 6141 5355 6193
rect 5389 6141 5422 6193
rect 5322 6125 5422 6141
rect 5322 6069 5355 6125
rect 5389 6069 5422 6125
rect 5322 6057 5422 6069
rect 5322 5997 5355 6057
rect 5389 5997 5422 6057
rect 5322 5989 5422 5997
rect 5322 5925 5355 5989
rect 5389 5925 5422 5989
rect 5322 5921 5422 5925
rect 5322 5819 5355 5921
rect 5389 5819 5422 5921
rect 5322 5815 5422 5819
rect 5322 5751 5355 5815
rect 5389 5751 5422 5815
rect 5322 5743 5422 5751
rect 5322 5683 5355 5743
rect 5389 5683 5422 5743
rect 5322 5671 5422 5683
rect 5322 5615 5355 5671
rect 5389 5615 5422 5671
rect 5322 5599 5422 5615
rect 5322 5547 5355 5599
rect 5389 5547 5422 5599
rect 5322 5527 5422 5547
rect 5322 5479 5355 5527
rect 5389 5479 5422 5527
rect 5322 5455 5422 5479
rect 5322 5411 5355 5455
rect 5389 5411 5422 5455
rect 5322 5383 5422 5411
rect 5322 5343 5355 5383
rect 5389 5343 5422 5383
rect 5322 5311 5422 5343
rect 5322 5275 5355 5311
rect 5389 5275 5422 5311
rect 5322 5241 5422 5275
rect 5322 5205 5355 5241
rect 5389 5205 5422 5241
rect 5322 5173 5422 5205
rect 5322 5133 5355 5173
rect 5389 5133 5422 5173
rect 5322 5105 5422 5133
rect 5322 5061 5355 5105
rect 5389 5061 5422 5105
rect 5322 5037 5422 5061
rect 5322 4989 5355 5037
rect 5389 4989 5422 5037
rect 5322 4969 5422 4989
rect 5322 4917 5355 4969
rect 5389 4917 5422 4969
rect 5322 4901 5422 4917
rect 5322 4845 5355 4901
rect 5389 4845 5422 4901
rect 5322 4833 5422 4845
rect 5322 4773 5355 4833
rect 5389 4773 5422 4833
rect 5322 4765 5422 4773
rect 5322 4731 5355 4765
rect 5389 4731 5422 4765
rect 5322 4697 5422 4731
rect 5322 4663 5355 4697
rect 5389 4663 5422 4697
rect 5322 4578 5422 4663
rect -5022 4545 5422 4578
rect -5022 4511 -4893 4545
rect -4859 4511 -4849 4545
rect -4787 4511 -4781 4545
rect -4715 4511 -4713 4545
rect -4679 4511 -4677 4545
rect -4611 4511 -4605 4545
rect -4543 4511 -4533 4545
rect -4475 4511 -4461 4545
rect -4407 4511 -4389 4545
rect -4339 4511 -4317 4545
rect -4271 4511 -4245 4545
rect -4203 4511 -4173 4545
rect -4135 4511 -4101 4545
rect -4067 4511 -4033 4545
rect -3995 4511 -3965 4545
rect -3923 4511 -3897 4545
rect -3851 4511 -3829 4545
rect -3779 4511 -3761 4545
rect -3707 4511 -3693 4545
rect -3635 4511 -3625 4545
rect -3563 4511 -3557 4545
rect -3491 4511 -3489 4545
rect -3455 4511 -3453 4545
rect -3387 4511 -3381 4545
rect -3319 4511 -3309 4545
rect -3251 4511 -3237 4545
rect -3183 4511 -3165 4545
rect -3115 4511 -3093 4545
rect -3047 4511 -3021 4545
rect -2979 4511 -2949 4545
rect -2911 4511 -2877 4545
rect -2843 4511 -2809 4545
rect -2771 4511 -2741 4545
rect -2699 4511 -2673 4545
rect -2627 4511 -2605 4545
rect -2555 4511 -2537 4545
rect -2483 4511 -2469 4545
rect -2411 4511 -2401 4545
rect -2339 4511 -2333 4545
rect -2267 4511 -2265 4545
rect -2231 4511 -2229 4545
rect -2163 4511 -2157 4545
rect -2095 4511 -2085 4545
rect -2027 4511 -2013 4545
rect -1959 4511 -1941 4545
rect -1891 4511 -1869 4545
rect -1823 4511 -1797 4545
rect -1755 4511 -1725 4545
rect -1687 4511 -1653 4545
rect -1619 4511 -1585 4545
rect -1547 4511 -1517 4545
rect -1475 4511 -1449 4545
rect -1403 4511 -1381 4545
rect -1331 4511 -1313 4545
rect -1259 4511 -1245 4545
rect -1187 4511 -1177 4545
rect -1115 4511 -1109 4545
rect -1043 4511 -1041 4545
rect -1007 4511 -1005 4545
rect -939 4511 -933 4545
rect -871 4511 -861 4545
rect -803 4511 -789 4545
rect -735 4511 -717 4545
rect -667 4511 -645 4545
rect -599 4511 -573 4545
rect -531 4511 -501 4545
rect -463 4511 -429 4545
rect -395 4511 -361 4545
rect -323 4511 -293 4545
rect -251 4511 -225 4545
rect -179 4511 -157 4545
rect -107 4511 -89 4545
rect -35 4511 -21 4545
rect 37 4511 47 4545
rect 109 4511 115 4545
rect 181 4511 183 4545
rect 217 4511 219 4545
rect 285 4511 291 4545
rect 353 4511 363 4545
rect 421 4511 435 4545
rect 489 4511 507 4545
rect 557 4511 579 4545
rect 625 4511 651 4545
rect 693 4511 723 4545
rect 761 4511 795 4545
rect 829 4511 863 4545
rect 901 4511 931 4545
rect 973 4511 999 4545
rect 1045 4511 1067 4545
rect 1117 4511 1135 4545
rect 1189 4511 1203 4545
rect 1261 4511 1271 4545
rect 1333 4511 1339 4545
rect 1405 4511 1407 4545
rect 1441 4511 1443 4545
rect 1509 4511 1515 4545
rect 1577 4511 1587 4545
rect 1645 4511 1659 4545
rect 1713 4511 1731 4545
rect 1781 4511 1803 4545
rect 1849 4511 1875 4545
rect 1917 4511 1947 4545
rect 1985 4511 2019 4545
rect 2053 4511 2087 4545
rect 2125 4511 2155 4545
rect 2197 4511 2223 4545
rect 2269 4511 2291 4545
rect 2341 4511 2359 4545
rect 2413 4511 2427 4545
rect 2485 4511 2495 4545
rect 2557 4511 2563 4545
rect 2629 4511 2631 4545
rect 2665 4511 2667 4545
rect 2733 4511 2739 4545
rect 2801 4511 2811 4545
rect 2869 4511 2883 4545
rect 2937 4511 2955 4545
rect 3005 4511 3027 4545
rect 3073 4511 3099 4545
rect 3141 4511 3171 4545
rect 3209 4511 3243 4545
rect 3277 4511 3311 4545
rect 3349 4511 3379 4545
rect 3421 4511 3447 4545
rect 3493 4511 3515 4545
rect 3565 4511 3583 4545
rect 3637 4511 3651 4545
rect 3709 4511 3719 4545
rect 3781 4511 3787 4545
rect 3853 4511 3855 4545
rect 3889 4511 3891 4545
rect 3957 4511 3963 4545
rect 4025 4511 4035 4545
rect 4093 4511 4107 4545
rect 4161 4511 4179 4545
rect 4229 4511 4251 4545
rect 4297 4511 4323 4545
rect 4365 4511 4395 4545
rect 4433 4511 4467 4545
rect 4501 4511 4535 4545
rect 4573 4511 4603 4545
rect 4645 4511 4671 4545
rect 4717 4511 4739 4545
rect 4789 4511 4807 4545
rect 4861 4511 4875 4545
rect 4933 4511 4943 4545
rect 5005 4511 5011 4545
rect 5077 4511 5079 4545
rect 5113 4511 5115 4545
rect 5181 4511 5187 4545
rect 5249 4511 5259 4545
rect 5293 4511 5422 4545
rect -5022 4478 5422 4511
rect -5022 4209 5422 4242
rect -5022 4175 -4893 4209
rect -4859 4175 -4849 4209
rect -4787 4175 -4781 4209
rect -4715 4175 -4713 4209
rect -4679 4175 -4677 4209
rect -4611 4175 -4605 4209
rect -4543 4175 -4533 4209
rect -4475 4175 -4461 4209
rect -4407 4175 -4389 4209
rect -4339 4175 -4317 4209
rect -4271 4175 -4245 4209
rect -4203 4175 -4173 4209
rect -4135 4175 -4101 4209
rect -4067 4175 -4033 4209
rect -3995 4175 -3965 4209
rect -3923 4175 -3897 4209
rect -3851 4175 -3829 4209
rect -3779 4175 -3761 4209
rect -3707 4175 -3693 4209
rect -3635 4175 -3625 4209
rect -3563 4175 -3557 4209
rect -3491 4175 -3489 4209
rect -3455 4175 -3453 4209
rect -3387 4175 -3381 4209
rect -3319 4175 -3309 4209
rect -3251 4175 -3237 4209
rect -3183 4175 -3165 4209
rect -3115 4175 -3093 4209
rect -3047 4175 -3021 4209
rect -2979 4175 -2949 4209
rect -2911 4175 -2877 4209
rect -2843 4175 -2809 4209
rect -2771 4175 -2741 4209
rect -2699 4175 -2673 4209
rect -2627 4175 -2605 4209
rect -2555 4175 -2537 4209
rect -2483 4175 -2469 4209
rect -2411 4175 -2401 4209
rect -2339 4175 -2333 4209
rect -2267 4175 -2265 4209
rect -2231 4175 -2229 4209
rect -2163 4175 -2157 4209
rect -2095 4175 -2085 4209
rect -2027 4175 -2013 4209
rect -1959 4175 -1941 4209
rect -1891 4175 -1869 4209
rect -1823 4175 -1797 4209
rect -1755 4175 -1725 4209
rect -1687 4175 -1653 4209
rect -1619 4175 -1585 4209
rect -1547 4175 -1517 4209
rect -1475 4175 -1449 4209
rect -1403 4175 -1381 4209
rect -1331 4175 -1313 4209
rect -1259 4175 -1245 4209
rect -1187 4175 -1177 4209
rect -1115 4175 -1109 4209
rect -1043 4175 -1041 4209
rect -1007 4175 -1005 4209
rect -939 4175 -933 4209
rect -871 4175 -861 4209
rect -803 4175 -789 4209
rect -735 4175 -717 4209
rect -667 4175 -645 4209
rect -599 4175 -573 4209
rect -531 4175 -501 4209
rect -463 4175 -429 4209
rect -395 4175 -361 4209
rect -323 4175 -293 4209
rect -251 4175 -225 4209
rect -179 4175 -157 4209
rect -107 4175 -89 4209
rect -35 4175 -21 4209
rect 37 4175 47 4209
rect 109 4175 115 4209
rect 181 4175 183 4209
rect 217 4175 219 4209
rect 285 4175 291 4209
rect 353 4175 363 4209
rect 421 4175 435 4209
rect 489 4175 507 4209
rect 557 4175 579 4209
rect 625 4175 651 4209
rect 693 4175 723 4209
rect 761 4175 795 4209
rect 829 4175 863 4209
rect 901 4175 931 4209
rect 973 4175 999 4209
rect 1045 4175 1067 4209
rect 1117 4175 1135 4209
rect 1189 4175 1203 4209
rect 1261 4175 1271 4209
rect 1333 4175 1339 4209
rect 1405 4175 1407 4209
rect 1441 4175 1443 4209
rect 1509 4175 1515 4209
rect 1577 4175 1587 4209
rect 1645 4175 1659 4209
rect 1713 4175 1731 4209
rect 1781 4175 1803 4209
rect 1849 4175 1875 4209
rect 1917 4175 1947 4209
rect 1985 4175 2019 4209
rect 2053 4175 2087 4209
rect 2125 4175 2155 4209
rect 2197 4175 2223 4209
rect 2269 4175 2291 4209
rect 2341 4175 2359 4209
rect 2413 4175 2427 4209
rect 2485 4175 2495 4209
rect 2557 4175 2563 4209
rect 2629 4175 2631 4209
rect 2665 4175 2667 4209
rect 2733 4175 2739 4209
rect 2801 4175 2811 4209
rect 2869 4175 2883 4209
rect 2937 4175 2955 4209
rect 3005 4175 3027 4209
rect 3073 4175 3099 4209
rect 3141 4175 3171 4209
rect 3209 4175 3243 4209
rect 3277 4175 3311 4209
rect 3349 4175 3379 4209
rect 3421 4175 3447 4209
rect 3493 4175 3515 4209
rect 3565 4175 3583 4209
rect 3637 4175 3651 4209
rect 3709 4175 3719 4209
rect 3781 4175 3787 4209
rect 3853 4175 3855 4209
rect 3889 4175 3891 4209
rect 3957 4175 3963 4209
rect 4025 4175 4035 4209
rect 4093 4175 4107 4209
rect 4161 4175 4179 4209
rect 4229 4175 4251 4209
rect 4297 4175 4323 4209
rect 4365 4175 4395 4209
rect 4433 4175 4467 4209
rect 4501 4175 4535 4209
rect 4573 4175 4603 4209
rect 4645 4175 4671 4209
rect 4717 4175 4739 4209
rect 4789 4175 4807 4209
rect 4861 4175 4875 4209
rect 4933 4175 4943 4209
rect 5005 4175 5011 4209
rect 5077 4175 5079 4209
rect 5113 4175 5115 4209
rect 5181 4175 5187 4209
rect 5249 4175 5259 4209
rect 5293 4175 5422 4209
rect -5022 4142 5422 4175
rect -5022 4047 -4922 4142
rect -5022 4013 -4989 4047
rect -4955 4013 -4922 4047
rect -5022 3999 -4922 4013
rect -5022 3945 -4989 3999
rect -4955 3945 -4922 3999
rect -5022 3927 -4922 3945
rect -5022 3877 -4989 3927
rect -4955 3877 -4922 3927
rect -5022 3855 -4922 3877
rect -5022 3809 -4989 3855
rect -4955 3809 -4922 3855
rect -5022 3783 -4922 3809
rect -5022 3741 -4989 3783
rect -4955 3741 -4922 3783
rect -5022 3711 -4922 3741
rect -5022 3673 -4989 3711
rect -4955 3673 -4922 3711
rect -5022 3639 -4922 3673
rect -5022 3605 -4989 3639
rect -4955 3605 -4922 3639
rect -5022 3571 -4922 3605
rect -5022 3533 -4989 3571
rect -4955 3533 -4922 3571
rect -5022 3503 -4922 3533
rect -5022 3461 -4989 3503
rect -4955 3461 -4922 3503
rect -5022 3435 -4922 3461
rect -5022 3389 -4989 3435
rect -4955 3389 -4922 3435
rect -5022 3367 -4922 3389
rect -5022 3317 -4989 3367
rect -4955 3317 -4922 3367
rect -5022 3299 -4922 3317
rect -5022 3245 -4989 3299
rect -4955 3245 -4922 3299
rect -5022 3231 -4922 3245
rect -5022 3173 -4989 3231
rect -4955 3173 -4922 3231
rect -5022 3163 -4922 3173
rect -5022 3101 -4989 3163
rect -4955 3101 -4922 3163
rect -5022 3095 -4922 3101
rect -5022 3029 -4989 3095
rect -4955 3029 -4922 3095
rect -5022 3027 -4922 3029
rect -5022 2993 -4989 3027
rect -4955 2993 -4922 3027
rect -5022 2991 -4922 2993
rect -5022 2925 -4989 2991
rect -4955 2925 -4922 2991
rect -5022 2919 -4922 2925
rect -5022 2857 -4989 2919
rect -4955 2857 -4922 2919
rect -5022 2847 -4922 2857
rect -5022 2789 -4989 2847
rect -4955 2789 -4922 2847
rect -5022 2775 -4922 2789
rect -5022 2721 -4989 2775
rect -4955 2721 -4922 2775
rect -5022 2703 -4922 2721
rect -5022 2653 -4989 2703
rect -4955 2653 -4922 2703
rect -5022 2631 -4922 2653
rect -5022 2585 -4989 2631
rect -4955 2585 -4922 2631
rect -5022 2559 -4922 2585
rect -5022 2517 -4989 2559
rect -4955 2517 -4922 2559
rect -5022 2487 -4922 2517
rect -5022 2449 -4989 2487
rect -4955 2449 -4922 2487
rect -5022 2415 -4922 2449
rect -5022 2381 -4989 2415
rect -4955 2381 -4922 2415
rect -5022 2347 -4922 2381
rect -5022 2309 -4989 2347
rect -4955 2309 -4922 2347
rect -5022 2279 -4922 2309
rect -5022 2237 -4989 2279
rect -4955 2237 -4922 2279
rect -5022 2211 -4922 2237
rect -5022 2165 -4989 2211
rect -4955 2165 -4922 2211
rect -5022 2143 -4922 2165
rect -5022 2093 -4989 2143
rect -4955 2093 -4922 2143
rect -5022 2075 -4922 2093
rect -5022 2021 -4989 2075
rect -4955 2021 -4922 2075
rect -5022 2007 -4922 2021
rect -5022 1973 -4989 2007
rect -4955 1973 -4922 2007
rect -5022 1878 -4922 1973
rect 5322 4047 5422 4142
rect 5322 4013 5355 4047
rect 5389 4013 5422 4047
rect 5322 3999 5422 4013
rect 5322 3945 5355 3999
rect 5389 3945 5422 3999
rect 5322 3927 5422 3945
rect 5322 3877 5355 3927
rect 5389 3877 5422 3927
rect 5322 3855 5422 3877
rect 5322 3809 5355 3855
rect 5389 3809 5422 3855
rect 5322 3783 5422 3809
rect 5322 3741 5355 3783
rect 5389 3741 5422 3783
rect 5322 3711 5422 3741
rect 5322 3673 5355 3711
rect 5389 3673 5422 3711
rect 5322 3639 5422 3673
rect 5322 3605 5355 3639
rect 5389 3605 5422 3639
rect 5322 3571 5422 3605
rect 5322 3533 5355 3571
rect 5389 3533 5422 3571
rect 5322 3503 5422 3533
rect 5322 3461 5355 3503
rect 5389 3461 5422 3503
rect 5322 3435 5422 3461
rect 5322 3389 5355 3435
rect 5389 3389 5422 3435
rect 5322 3367 5422 3389
rect 5322 3317 5355 3367
rect 5389 3317 5422 3367
rect 5322 3299 5422 3317
rect 5322 3245 5355 3299
rect 5389 3245 5422 3299
rect 5322 3231 5422 3245
rect 5322 3173 5355 3231
rect 5389 3173 5422 3231
rect 5322 3163 5422 3173
rect 5322 3101 5355 3163
rect 5389 3101 5422 3163
rect 5322 3095 5422 3101
rect 5322 3029 5355 3095
rect 5389 3029 5422 3095
rect 5322 3027 5422 3029
rect 5322 2993 5355 3027
rect 5389 2993 5422 3027
rect 5322 2991 5422 2993
rect 5322 2925 5355 2991
rect 5389 2925 5422 2991
rect 5322 2919 5422 2925
rect 5322 2857 5355 2919
rect 5389 2857 5422 2919
rect 5322 2847 5422 2857
rect 5322 2789 5355 2847
rect 5389 2789 5422 2847
rect 5322 2775 5422 2789
rect 5322 2721 5355 2775
rect 5389 2721 5422 2775
rect 5322 2703 5422 2721
rect 5322 2653 5355 2703
rect 5389 2653 5422 2703
rect 5322 2631 5422 2653
rect 5322 2585 5355 2631
rect 5389 2585 5422 2631
rect 5322 2559 5422 2585
rect 5322 2517 5355 2559
rect 5389 2517 5422 2559
rect 5322 2487 5422 2517
rect 5322 2449 5355 2487
rect 5389 2449 5422 2487
rect 5322 2415 5422 2449
rect 5322 2381 5355 2415
rect 5389 2381 5422 2415
rect 5322 2347 5422 2381
rect 5322 2309 5355 2347
rect 5389 2309 5422 2347
rect 5322 2279 5422 2309
rect 5322 2237 5355 2279
rect 5389 2237 5422 2279
rect 5322 2211 5422 2237
rect 5322 2165 5355 2211
rect 5389 2165 5422 2211
rect 5322 2143 5422 2165
rect 5322 2093 5355 2143
rect 5389 2093 5422 2143
rect 5322 2075 5422 2093
rect 5322 2021 5355 2075
rect 5389 2021 5422 2075
rect 5322 2007 5422 2021
rect 5322 1973 5355 2007
rect 5389 1973 5422 2007
rect 5322 1878 5422 1973
rect -5022 1845 5422 1878
rect -5022 1811 -4893 1845
rect -4859 1811 -4849 1845
rect -4787 1811 -4781 1845
rect -4715 1811 -4713 1845
rect -4679 1811 -4677 1845
rect -4611 1811 -4605 1845
rect -4543 1811 -4533 1845
rect -4475 1811 -4461 1845
rect -4407 1811 -4389 1845
rect -4339 1811 -4317 1845
rect -4271 1811 -4245 1845
rect -4203 1811 -4173 1845
rect -4135 1811 -4101 1845
rect -4067 1811 -4033 1845
rect -3995 1811 -3965 1845
rect -3923 1811 -3897 1845
rect -3851 1811 -3829 1845
rect -3779 1811 -3761 1845
rect -3707 1811 -3693 1845
rect -3635 1811 -3625 1845
rect -3563 1811 -3557 1845
rect -3491 1811 -3489 1845
rect -3455 1811 -3453 1845
rect -3387 1811 -3381 1845
rect -3319 1811 -3309 1845
rect -3251 1811 -3237 1845
rect -3183 1811 -3165 1845
rect -3115 1811 -3093 1845
rect -3047 1811 -3021 1845
rect -2979 1811 -2949 1845
rect -2911 1811 -2877 1845
rect -2843 1811 -2809 1845
rect -2771 1811 -2741 1845
rect -2699 1811 -2673 1845
rect -2627 1811 -2605 1845
rect -2555 1811 -2537 1845
rect -2483 1811 -2469 1845
rect -2411 1811 -2401 1845
rect -2339 1811 -2333 1845
rect -2267 1811 -2265 1845
rect -2231 1811 -2229 1845
rect -2163 1811 -2157 1845
rect -2095 1811 -2085 1845
rect -2027 1811 -2013 1845
rect -1959 1811 -1941 1845
rect -1891 1811 -1869 1845
rect -1823 1811 -1797 1845
rect -1755 1811 -1725 1845
rect -1687 1811 -1653 1845
rect -1619 1811 -1585 1845
rect -1547 1811 -1517 1845
rect -1475 1811 -1449 1845
rect -1403 1811 -1381 1845
rect -1331 1811 -1313 1845
rect -1259 1811 -1245 1845
rect -1187 1811 -1177 1845
rect -1115 1811 -1109 1845
rect -1043 1811 -1041 1845
rect -1007 1811 -1005 1845
rect -939 1811 -933 1845
rect -871 1811 -861 1845
rect -803 1811 -789 1845
rect -735 1811 -717 1845
rect -667 1811 -645 1845
rect -599 1811 -573 1845
rect -531 1811 -501 1845
rect -463 1811 -429 1845
rect -395 1811 -361 1845
rect -323 1811 -293 1845
rect -251 1811 -225 1845
rect -179 1811 -157 1845
rect -107 1811 -89 1845
rect -35 1811 -21 1845
rect 37 1811 47 1845
rect 109 1811 115 1845
rect 181 1811 183 1845
rect 217 1811 219 1845
rect 285 1811 291 1845
rect 353 1811 363 1845
rect 421 1811 435 1845
rect 489 1811 507 1845
rect 557 1811 579 1845
rect 625 1811 651 1845
rect 693 1811 723 1845
rect 761 1811 795 1845
rect 829 1811 863 1845
rect 901 1811 931 1845
rect 973 1811 999 1845
rect 1045 1811 1067 1845
rect 1117 1811 1135 1845
rect 1189 1811 1203 1845
rect 1261 1811 1271 1845
rect 1333 1811 1339 1845
rect 1405 1811 1407 1845
rect 1441 1811 1443 1845
rect 1509 1811 1515 1845
rect 1577 1811 1587 1845
rect 1645 1811 1659 1845
rect 1713 1811 1731 1845
rect 1781 1811 1803 1845
rect 1849 1811 1875 1845
rect 1917 1811 1947 1845
rect 1985 1811 2019 1845
rect 2053 1811 2087 1845
rect 2125 1811 2155 1845
rect 2197 1811 2223 1845
rect 2269 1811 2291 1845
rect 2341 1811 2359 1845
rect 2413 1811 2427 1845
rect 2485 1811 2495 1845
rect 2557 1811 2563 1845
rect 2629 1811 2631 1845
rect 2665 1811 2667 1845
rect 2733 1811 2739 1845
rect 2801 1811 2811 1845
rect 2869 1811 2883 1845
rect 2937 1811 2955 1845
rect 3005 1811 3027 1845
rect 3073 1811 3099 1845
rect 3141 1811 3171 1845
rect 3209 1811 3243 1845
rect 3277 1811 3311 1845
rect 3349 1811 3379 1845
rect 3421 1811 3447 1845
rect 3493 1811 3515 1845
rect 3565 1811 3583 1845
rect 3637 1811 3651 1845
rect 3709 1811 3719 1845
rect 3781 1811 3787 1845
rect 3853 1811 3855 1845
rect 3889 1811 3891 1845
rect 3957 1811 3963 1845
rect 4025 1811 4035 1845
rect 4093 1811 4107 1845
rect 4161 1811 4179 1845
rect 4229 1811 4251 1845
rect 4297 1811 4323 1845
rect 4365 1811 4395 1845
rect 4433 1811 4467 1845
rect 4501 1811 4535 1845
rect 4573 1811 4603 1845
rect 4645 1811 4671 1845
rect 4717 1811 4739 1845
rect 4789 1811 4807 1845
rect 4861 1811 4875 1845
rect 4933 1811 4943 1845
rect 5005 1811 5011 1845
rect 5077 1811 5079 1845
rect 5113 1811 5115 1845
rect 5181 1811 5187 1845
rect 5249 1811 5259 1845
rect 5293 1811 5422 1845
rect -5022 1778 5422 1811
<< viali >>
rect -4893 10255 -4859 10289
rect -4821 10255 -4815 10289
rect -4815 10255 -4787 10289
rect -4749 10255 -4747 10289
rect -4747 10255 -4715 10289
rect -4677 10255 -4645 10289
rect -4645 10255 -4643 10289
rect -4605 10255 -4577 10289
rect -4577 10255 -4571 10289
rect -4533 10255 -4509 10289
rect -4509 10255 -4499 10289
rect -4461 10255 -4441 10289
rect -4441 10255 -4427 10289
rect -4389 10255 -4373 10289
rect -4373 10255 -4355 10289
rect -4317 10255 -4305 10289
rect -4305 10255 -4283 10289
rect -4245 10255 -4237 10289
rect -4237 10255 -4211 10289
rect -4173 10255 -4169 10289
rect -4169 10255 -4139 10289
rect -4101 10255 -4067 10289
rect -4029 10255 -3999 10289
rect -3999 10255 -3995 10289
rect -3957 10255 -3931 10289
rect -3931 10255 -3923 10289
rect -3885 10255 -3863 10289
rect -3863 10255 -3851 10289
rect -3813 10255 -3795 10289
rect -3795 10255 -3779 10289
rect -3741 10255 -3727 10289
rect -3727 10255 -3707 10289
rect -3669 10255 -3659 10289
rect -3659 10255 -3635 10289
rect -3597 10255 -3591 10289
rect -3591 10255 -3563 10289
rect -3525 10255 -3523 10289
rect -3523 10255 -3491 10289
rect -3453 10255 -3421 10289
rect -3421 10255 -3419 10289
rect -3381 10255 -3353 10289
rect -3353 10255 -3347 10289
rect -3309 10255 -3285 10289
rect -3285 10255 -3275 10289
rect -3237 10255 -3217 10289
rect -3217 10255 -3203 10289
rect -3165 10255 -3149 10289
rect -3149 10255 -3131 10289
rect -3093 10255 -3081 10289
rect -3081 10255 -3059 10289
rect -3021 10255 -3013 10289
rect -3013 10255 -2987 10289
rect -2949 10255 -2945 10289
rect -2945 10255 -2915 10289
rect -2877 10255 -2843 10289
rect -2805 10255 -2775 10289
rect -2775 10255 -2771 10289
rect -2733 10255 -2707 10289
rect -2707 10255 -2699 10289
rect -2661 10255 -2639 10289
rect -2639 10255 -2627 10289
rect -2589 10255 -2571 10289
rect -2571 10255 -2555 10289
rect -2517 10255 -2503 10289
rect -2503 10255 -2483 10289
rect -2445 10255 -2435 10289
rect -2435 10255 -2411 10289
rect -2373 10255 -2367 10289
rect -2367 10255 -2339 10289
rect -2301 10255 -2299 10289
rect -2299 10255 -2267 10289
rect -2229 10255 -2197 10289
rect -2197 10255 -2195 10289
rect -2157 10255 -2129 10289
rect -2129 10255 -2123 10289
rect -2085 10255 -2061 10289
rect -2061 10255 -2051 10289
rect -2013 10255 -1993 10289
rect -1993 10255 -1979 10289
rect -1941 10255 -1925 10289
rect -1925 10255 -1907 10289
rect -1869 10255 -1857 10289
rect -1857 10255 -1835 10289
rect -1797 10255 -1789 10289
rect -1789 10255 -1763 10289
rect -1725 10255 -1721 10289
rect -1721 10255 -1691 10289
rect -1653 10255 -1619 10289
rect -1581 10255 -1551 10289
rect -1551 10255 -1547 10289
rect -1509 10255 -1483 10289
rect -1483 10255 -1475 10289
rect -1437 10255 -1415 10289
rect -1415 10255 -1403 10289
rect -1365 10255 -1347 10289
rect -1347 10255 -1331 10289
rect -1293 10255 -1279 10289
rect -1279 10255 -1259 10289
rect -1221 10255 -1211 10289
rect -1211 10255 -1187 10289
rect -1149 10255 -1143 10289
rect -1143 10255 -1115 10289
rect -1077 10255 -1075 10289
rect -1075 10255 -1043 10289
rect -1005 10255 -973 10289
rect -973 10255 -971 10289
rect -933 10255 -905 10289
rect -905 10255 -899 10289
rect -861 10255 -837 10289
rect -837 10255 -827 10289
rect -789 10255 -769 10289
rect -769 10255 -755 10289
rect -717 10255 -701 10289
rect -701 10255 -683 10289
rect -645 10255 -633 10289
rect -633 10255 -611 10289
rect -573 10255 -565 10289
rect -565 10255 -539 10289
rect -501 10255 -497 10289
rect -497 10255 -467 10289
rect -429 10255 -395 10289
rect -357 10255 -327 10289
rect -327 10255 -323 10289
rect -285 10255 -259 10289
rect -259 10255 -251 10289
rect -213 10255 -191 10289
rect -191 10255 -179 10289
rect -141 10255 -123 10289
rect -123 10255 -107 10289
rect -69 10255 -55 10289
rect -55 10255 -35 10289
rect 3 10255 13 10289
rect 13 10255 37 10289
rect 75 10255 81 10289
rect 81 10255 109 10289
rect 147 10255 149 10289
rect 149 10255 181 10289
rect 219 10255 251 10289
rect 251 10255 253 10289
rect 291 10255 319 10289
rect 319 10255 325 10289
rect 363 10255 387 10289
rect 387 10255 397 10289
rect 435 10255 455 10289
rect 455 10255 469 10289
rect 507 10255 523 10289
rect 523 10255 541 10289
rect 579 10255 591 10289
rect 591 10255 613 10289
rect 651 10255 659 10289
rect 659 10255 685 10289
rect 723 10255 727 10289
rect 727 10255 757 10289
rect 795 10255 829 10289
rect 867 10255 897 10289
rect 897 10255 901 10289
rect 939 10255 965 10289
rect 965 10255 973 10289
rect 1011 10255 1033 10289
rect 1033 10255 1045 10289
rect 1083 10255 1101 10289
rect 1101 10255 1117 10289
rect 1155 10255 1169 10289
rect 1169 10255 1189 10289
rect 1227 10255 1237 10289
rect 1237 10255 1261 10289
rect 1299 10255 1305 10289
rect 1305 10255 1333 10289
rect 1371 10255 1373 10289
rect 1373 10255 1405 10289
rect 1443 10255 1475 10289
rect 1475 10255 1477 10289
rect 1515 10255 1543 10289
rect 1543 10255 1549 10289
rect 1587 10255 1611 10289
rect 1611 10255 1621 10289
rect 1659 10255 1679 10289
rect 1679 10255 1693 10289
rect 1731 10255 1747 10289
rect 1747 10255 1765 10289
rect 1803 10255 1815 10289
rect 1815 10255 1837 10289
rect 1875 10255 1883 10289
rect 1883 10255 1909 10289
rect 1947 10255 1951 10289
rect 1951 10255 1981 10289
rect 2019 10255 2053 10289
rect 2091 10255 2121 10289
rect 2121 10255 2125 10289
rect 2163 10255 2189 10289
rect 2189 10255 2197 10289
rect 2235 10255 2257 10289
rect 2257 10255 2269 10289
rect 2307 10255 2325 10289
rect 2325 10255 2341 10289
rect 2379 10255 2393 10289
rect 2393 10255 2413 10289
rect 2451 10255 2461 10289
rect 2461 10255 2485 10289
rect 2523 10255 2529 10289
rect 2529 10255 2557 10289
rect 2595 10255 2597 10289
rect 2597 10255 2629 10289
rect 2667 10255 2699 10289
rect 2699 10255 2701 10289
rect 2739 10255 2767 10289
rect 2767 10255 2773 10289
rect 2811 10255 2835 10289
rect 2835 10255 2845 10289
rect 2883 10255 2903 10289
rect 2903 10255 2917 10289
rect 2955 10255 2971 10289
rect 2971 10255 2989 10289
rect 3027 10255 3039 10289
rect 3039 10255 3061 10289
rect 3099 10255 3107 10289
rect 3107 10255 3133 10289
rect 3171 10255 3175 10289
rect 3175 10255 3205 10289
rect 3243 10255 3277 10289
rect 3315 10255 3345 10289
rect 3345 10255 3349 10289
rect 3387 10255 3413 10289
rect 3413 10255 3421 10289
rect 3459 10255 3481 10289
rect 3481 10255 3493 10289
rect 3531 10255 3549 10289
rect 3549 10255 3565 10289
rect 3603 10255 3617 10289
rect 3617 10255 3637 10289
rect 3675 10255 3685 10289
rect 3685 10255 3709 10289
rect 3747 10255 3753 10289
rect 3753 10255 3781 10289
rect 3819 10255 3821 10289
rect 3821 10255 3853 10289
rect 3891 10255 3923 10289
rect 3923 10255 3925 10289
rect 3963 10255 3991 10289
rect 3991 10255 3997 10289
rect 4035 10255 4059 10289
rect 4059 10255 4069 10289
rect 4107 10255 4127 10289
rect 4127 10255 4141 10289
rect 4179 10255 4195 10289
rect 4195 10255 4213 10289
rect 4251 10255 4263 10289
rect 4263 10255 4285 10289
rect 4323 10255 4331 10289
rect 4331 10255 4357 10289
rect 4395 10255 4399 10289
rect 4399 10255 4429 10289
rect 4467 10255 4501 10289
rect 4539 10255 4569 10289
rect 4569 10255 4573 10289
rect 4611 10255 4637 10289
rect 4637 10255 4645 10289
rect 4683 10255 4705 10289
rect 4705 10255 4717 10289
rect 4755 10255 4773 10289
rect 4773 10255 4789 10289
rect 4827 10255 4841 10289
rect 4841 10255 4861 10289
rect 4899 10255 4909 10289
rect 4909 10255 4933 10289
rect 4971 10255 4977 10289
rect 4977 10255 5005 10289
rect 5043 10255 5045 10289
rect 5045 10255 5077 10289
rect 5115 10255 5147 10289
rect 5147 10255 5149 10289
rect 5187 10255 5215 10289
rect 5215 10255 5221 10289
rect 5259 10255 5293 10289
rect -4989 9899 -4955 9919
rect -4989 9885 -4955 9899
rect -4989 9831 -4955 9847
rect -4989 9813 -4955 9831
rect -4989 9763 -4955 9775
rect -4989 9741 -4955 9763
rect -4989 9695 -4955 9703
rect -4989 9669 -4955 9695
rect -4989 9627 -4955 9631
rect -4989 9597 -4955 9627
rect -4989 9525 -4955 9559
rect -4989 9457 -4955 9487
rect -4989 9453 -4955 9457
rect -4989 9389 -4955 9415
rect -4989 9381 -4955 9389
rect -4989 9321 -4955 9343
rect -4989 9309 -4955 9321
rect -4989 9253 -4955 9271
rect -4989 9237 -4955 9253
rect -4989 9185 -4955 9199
rect -4989 9165 -4955 9185
rect -4989 9117 -4955 9127
rect -4989 9093 -4955 9117
rect -4989 9049 -4955 9055
rect -4989 9021 -4955 9049
rect -4989 8981 -4955 8983
rect -4989 8949 -4955 8981
rect -4989 8879 -4955 8911
rect -4989 8877 -4955 8879
rect -4989 8811 -4955 8839
rect -4989 8805 -4955 8811
rect -4989 8743 -4955 8767
rect -4989 8733 -4955 8743
rect -4989 8675 -4955 8695
rect -4989 8661 -4955 8675
rect -4989 8607 -4955 8623
rect -4989 8589 -4955 8607
rect -4989 8539 -4955 8551
rect -4989 8517 -4955 8539
rect -4989 8471 -4955 8479
rect -4989 8445 -4955 8471
rect -4989 8403 -4955 8407
rect -4989 8373 -4955 8403
rect -4989 8301 -4955 8335
rect -4989 8233 -4955 8263
rect -4989 8229 -4955 8233
rect -4989 8165 -4955 8191
rect -4989 8157 -4955 8165
rect -4989 8097 -4955 8119
rect -4989 8085 -4955 8097
rect -4989 8029 -4955 8047
rect -4989 8013 -4955 8029
rect -4989 7961 -4955 7975
rect -4989 7941 -4955 7961
rect -4989 7893 -4955 7903
rect -4989 7869 -4955 7893
rect -4989 7825 -4955 7831
rect -4989 7797 -4955 7825
rect -4989 7757 -4955 7759
rect -4989 7725 -4955 7757
rect -4989 7655 -4955 7687
rect -4989 7653 -4955 7655
rect -4989 7587 -4955 7615
rect -4989 7581 -4955 7587
rect -4989 7519 -4955 7543
rect -4989 7509 -4955 7519
rect -4989 7451 -4955 7471
rect -4989 7437 -4955 7451
rect -4989 7383 -4955 7399
rect -4989 7365 -4955 7383
rect -4989 7315 -4955 7327
rect -4989 7293 -4955 7315
rect -4989 7247 -4955 7255
rect -4989 7221 -4955 7247
rect -4989 7179 -4955 7183
rect -4989 7149 -4955 7179
rect -4989 7077 -4955 7111
rect 5355 9899 5389 9919
rect 5355 9885 5389 9899
rect 5355 9831 5389 9847
rect 5355 9813 5389 9831
rect 5355 9763 5389 9775
rect 5355 9741 5389 9763
rect 5355 9695 5389 9703
rect 5355 9669 5389 9695
rect 5355 9627 5389 9631
rect 5355 9597 5389 9627
rect 5355 9525 5389 9559
rect 5355 9457 5389 9487
rect 5355 9453 5389 9457
rect 5355 9389 5389 9415
rect 5355 9381 5389 9389
rect 5355 9321 5389 9343
rect 5355 9309 5389 9321
rect 5355 9253 5389 9271
rect 5355 9237 5389 9253
rect 5355 9185 5389 9199
rect 5355 9165 5389 9185
rect 5355 9117 5389 9127
rect 5355 9093 5389 9117
rect 5355 9049 5389 9055
rect 5355 9021 5389 9049
rect 5355 8981 5389 8983
rect 5355 8949 5389 8981
rect 5355 8879 5389 8911
rect 5355 8877 5389 8879
rect 5355 8811 5389 8839
rect 5355 8805 5389 8811
rect 5355 8743 5389 8767
rect 5355 8733 5389 8743
rect 5355 8675 5389 8695
rect 5355 8661 5389 8675
rect 5355 8607 5389 8623
rect 5355 8589 5389 8607
rect 5355 8539 5389 8551
rect 5355 8517 5389 8539
rect 5355 8471 5389 8479
rect 5355 8445 5389 8471
rect 5355 8403 5389 8407
rect 5355 8373 5389 8403
rect 5355 8301 5389 8335
rect 5355 8233 5389 8263
rect 5355 8229 5389 8233
rect 5355 8165 5389 8191
rect 5355 8157 5389 8165
rect 5355 8097 5389 8119
rect 5355 8085 5389 8097
rect 5355 8029 5389 8047
rect 5355 8013 5389 8029
rect 5355 7961 5389 7975
rect 5355 7941 5389 7961
rect 5355 7893 5389 7903
rect 5355 7869 5389 7893
rect 5355 7825 5389 7831
rect 5355 7797 5389 7825
rect 5355 7757 5389 7759
rect 5355 7725 5389 7757
rect 5355 7655 5389 7687
rect 5355 7653 5389 7655
rect 5355 7587 5389 7615
rect 5355 7581 5389 7587
rect 5355 7519 5389 7543
rect 5355 7509 5389 7519
rect 5355 7451 5389 7471
rect 5355 7437 5389 7451
rect 5355 7383 5389 7399
rect 5355 7365 5389 7383
rect 5355 7315 5389 7327
rect 5355 7293 5389 7315
rect 5355 7247 5389 7255
rect 5355 7221 5389 7247
rect 5355 7179 5389 7183
rect 5355 7149 5389 7179
rect -145 7065 -111 7099
rect 315 7065 349 7099
rect -4989 7009 -4955 7039
rect -4989 7005 -4955 7009
rect -4989 6941 -4955 6967
rect -4989 6933 -4955 6941
rect -4989 6873 -4955 6895
rect -4989 6861 -4955 6873
rect -4989 6805 -4955 6823
rect -4989 6789 -4955 6805
rect -4989 6737 -4955 6751
rect -4989 6717 -4955 6737
rect -4989 6669 -4955 6679
rect -4989 6645 -4955 6669
rect -4989 6601 -4955 6607
rect -4989 6573 -4955 6601
rect -4989 6533 -4955 6535
rect -4989 6501 -4955 6533
rect -4989 6431 -4955 6463
rect -4989 6429 -4955 6431
rect -4989 6363 -4955 6391
rect -4989 6357 -4955 6363
rect -4989 6295 -4955 6319
rect -4989 6285 -4955 6295
rect -4989 6227 -4955 6247
rect -4989 6213 -4955 6227
rect -4989 6159 -4955 6175
rect -4989 6141 -4955 6159
rect -4989 6091 -4955 6103
rect -4989 6069 -4955 6091
rect -4989 6023 -4955 6031
rect -4989 5997 -4955 6023
rect -4989 5955 -4955 5959
rect -4989 5925 -4955 5955
rect -4989 5853 -4955 5887
rect -4989 5785 -4955 5815
rect -4989 5781 -4955 5785
rect -4989 5717 -4955 5743
rect -4989 5709 -4955 5717
rect -4989 5649 -4955 5671
rect -4989 5637 -4955 5649
rect -4989 5581 -4955 5599
rect -4989 5565 -4955 5581
rect -4989 5513 -4955 5527
rect -4989 5493 -4955 5513
rect -4989 5445 -4955 5455
rect -4989 5421 -4955 5445
rect -4989 5377 -4955 5383
rect -4989 5349 -4955 5377
rect -4989 5309 -4955 5311
rect -4989 5277 -4955 5309
rect -4989 5207 -4955 5239
rect -4989 5205 -4955 5207
rect -4989 5139 -4955 5167
rect -4989 5133 -4955 5139
rect -4989 5071 -4955 5095
rect -4989 5061 -4955 5071
rect -4989 5003 -4955 5023
rect -4989 4989 -4955 5003
rect -4989 4935 -4955 4951
rect -4989 4917 -4955 4935
rect -4989 4867 -4955 4879
rect -4989 4845 -4955 4867
rect -4989 4799 -4955 4807
rect -4989 4773 -4955 4799
rect 5355 7077 5389 7111
rect 5355 7009 5389 7039
rect 5355 7005 5389 7009
rect 5355 6941 5389 6967
rect 5355 6933 5389 6941
rect 5355 6873 5389 6895
rect 5355 6861 5389 6873
rect 5355 6805 5389 6823
rect 5355 6789 5389 6805
rect 5355 6737 5389 6751
rect 5355 6717 5389 6737
rect 5355 6669 5389 6679
rect 5355 6645 5389 6669
rect 5355 6601 5389 6607
rect 5355 6573 5389 6601
rect 5355 6533 5389 6535
rect 5355 6501 5389 6533
rect 5355 6431 5389 6463
rect 5355 6429 5389 6431
rect 5355 6363 5389 6391
rect 5355 6357 5389 6363
rect 5355 6295 5389 6319
rect 5355 6285 5389 6295
rect 5355 6227 5389 6247
rect 5355 6213 5389 6227
rect 5355 6159 5389 6175
rect 5355 6141 5389 6159
rect 5355 6091 5389 6103
rect 5355 6069 5389 6091
rect 5355 6023 5389 6031
rect 5355 5997 5389 6023
rect 5355 5955 5389 5959
rect 5355 5925 5389 5955
rect 5355 5853 5389 5887
rect 5355 5785 5389 5815
rect 5355 5781 5389 5785
rect 5355 5717 5389 5743
rect 5355 5709 5389 5717
rect 5355 5649 5389 5671
rect 5355 5637 5389 5649
rect 5355 5581 5389 5599
rect 5355 5565 5389 5581
rect 5355 5513 5389 5527
rect 5355 5493 5389 5513
rect 5355 5445 5389 5455
rect 5355 5421 5389 5445
rect 5355 5377 5389 5383
rect 5355 5349 5389 5377
rect 5355 5309 5389 5311
rect 5355 5277 5389 5309
rect 5355 5207 5389 5239
rect 5355 5205 5389 5207
rect 5355 5139 5389 5167
rect 5355 5133 5389 5139
rect 5355 5071 5389 5095
rect 5355 5061 5389 5071
rect 5355 5003 5389 5023
rect 5355 4989 5389 5003
rect 5355 4935 5389 4951
rect 5355 4917 5389 4935
rect 5355 4867 5389 4879
rect 5355 4845 5389 4867
rect 5355 4799 5389 4807
rect 5355 4773 5389 4799
rect -4893 4511 -4859 4545
rect -4821 4511 -4815 4545
rect -4815 4511 -4787 4545
rect -4749 4511 -4747 4545
rect -4747 4511 -4715 4545
rect -4677 4511 -4645 4545
rect -4645 4511 -4643 4545
rect -4605 4511 -4577 4545
rect -4577 4511 -4571 4545
rect -4533 4511 -4509 4545
rect -4509 4511 -4499 4545
rect -4461 4511 -4441 4545
rect -4441 4511 -4427 4545
rect -4389 4511 -4373 4545
rect -4373 4511 -4355 4545
rect -4317 4511 -4305 4545
rect -4305 4511 -4283 4545
rect -4245 4511 -4237 4545
rect -4237 4511 -4211 4545
rect -4173 4511 -4169 4545
rect -4169 4511 -4139 4545
rect -4101 4511 -4067 4545
rect -4029 4511 -3999 4545
rect -3999 4511 -3995 4545
rect -3957 4511 -3931 4545
rect -3931 4511 -3923 4545
rect -3885 4511 -3863 4545
rect -3863 4511 -3851 4545
rect -3813 4511 -3795 4545
rect -3795 4511 -3779 4545
rect -3741 4511 -3727 4545
rect -3727 4511 -3707 4545
rect -3669 4511 -3659 4545
rect -3659 4511 -3635 4545
rect -3597 4511 -3591 4545
rect -3591 4511 -3563 4545
rect -3525 4511 -3523 4545
rect -3523 4511 -3491 4545
rect -3453 4511 -3421 4545
rect -3421 4511 -3419 4545
rect -3381 4511 -3353 4545
rect -3353 4511 -3347 4545
rect -3309 4511 -3285 4545
rect -3285 4511 -3275 4545
rect -3237 4511 -3217 4545
rect -3217 4511 -3203 4545
rect -3165 4511 -3149 4545
rect -3149 4511 -3131 4545
rect -3093 4511 -3081 4545
rect -3081 4511 -3059 4545
rect -3021 4511 -3013 4545
rect -3013 4511 -2987 4545
rect -2949 4511 -2945 4545
rect -2945 4511 -2915 4545
rect -2877 4511 -2843 4545
rect -2805 4511 -2775 4545
rect -2775 4511 -2771 4545
rect -2733 4511 -2707 4545
rect -2707 4511 -2699 4545
rect -2661 4511 -2639 4545
rect -2639 4511 -2627 4545
rect -2589 4511 -2571 4545
rect -2571 4511 -2555 4545
rect -2517 4511 -2503 4545
rect -2503 4511 -2483 4545
rect -2445 4511 -2435 4545
rect -2435 4511 -2411 4545
rect -2373 4511 -2367 4545
rect -2367 4511 -2339 4545
rect -2301 4511 -2299 4545
rect -2299 4511 -2267 4545
rect -2229 4511 -2197 4545
rect -2197 4511 -2195 4545
rect -2157 4511 -2129 4545
rect -2129 4511 -2123 4545
rect -2085 4511 -2061 4545
rect -2061 4511 -2051 4545
rect -2013 4511 -1993 4545
rect -1993 4511 -1979 4545
rect -1941 4511 -1925 4545
rect -1925 4511 -1907 4545
rect -1869 4511 -1857 4545
rect -1857 4511 -1835 4545
rect -1797 4511 -1789 4545
rect -1789 4511 -1763 4545
rect -1725 4511 -1721 4545
rect -1721 4511 -1691 4545
rect -1653 4511 -1619 4545
rect -1581 4511 -1551 4545
rect -1551 4511 -1547 4545
rect -1509 4511 -1483 4545
rect -1483 4511 -1475 4545
rect -1437 4511 -1415 4545
rect -1415 4511 -1403 4545
rect -1365 4511 -1347 4545
rect -1347 4511 -1331 4545
rect -1293 4511 -1279 4545
rect -1279 4511 -1259 4545
rect -1221 4511 -1211 4545
rect -1211 4511 -1187 4545
rect -1149 4511 -1143 4545
rect -1143 4511 -1115 4545
rect -1077 4511 -1075 4545
rect -1075 4511 -1043 4545
rect -1005 4511 -973 4545
rect -973 4511 -971 4545
rect -933 4511 -905 4545
rect -905 4511 -899 4545
rect -861 4511 -837 4545
rect -837 4511 -827 4545
rect -789 4511 -769 4545
rect -769 4511 -755 4545
rect -717 4511 -701 4545
rect -701 4511 -683 4545
rect -645 4511 -633 4545
rect -633 4511 -611 4545
rect -573 4511 -565 4545
rect -565 4511 -539 4545
rect -501 4511 -497 4545
rect -497 4511 -467 4545
rect -429 4511 -395 4545
rect -357 4511 -327 4545
rect -327 4511 -323 4545
rect -285 4511 -259 4545
rect -259 4511 -251 4545
rect -213 4511 -191 4545
rect -191 4511 -179 4545
rect -141 4511 -123 4545
rect -123 4511 -107 4545
rect -69 4511 -55 4545
rect -55 4511 -35 4545
rect 3 4511 13 4545
rect 13 4511 37 4545
rect 75 4511 81 4545
rect 81 4511 109 4545
rect 147 4511 149 4545
rect 149 4511 181 4545
rect 219 4511 251 4545
rect 251 4511 253 4545
rect 291 4511 319 4545
rect 319 4511 325 4545
rect 363 4511 387 4545
rect 387 4511 397 4545
rect 435 4511 455 4545
rect 455 4511 469 4545
rect 507 4511 523 4545
rect 523 4511 541 4545
rect 579 4511 591 4545
rect 591 4511 613 4545
rect 651 4511 659 4545
rect 659 4511 685 4545
rect 723 4511 727 4545
rect 727 4511 757 4545
rect 795 4511 829 4545
rect 867 4511 897 4545
rect 897 4511 901 4545
rect 939 4511 965 4545
rect 965 4511 973 4545
rect 1011 4511 1033 4545
rect 1033 4511 1045 4545
rect 1083 4511 1101 4545
rect 1101 4511 1117 4545
rect 1155 4511 1169 4545
rect 1169 4511 1189 4545
rect 1227 4511 1237 4545
rect 1237 4511 1261 4545
rect 1299 4511 1305 4545
rect 1305 4511 1333 4545
rect 1371 4511 1373 4545
rect 1373 4511 1405 4545
rect 1443 4511 1475 4545
rect 1475 4511 1477 4545
rect 1515 4511 1543 4545
rect 1543 4511 1549 4545
rect 1587 4511 1611 4545
rect 1611 4511 1621 4545
rect 1659 4511 1679 4545
rect 1679 4511 1693 4545
rect 1731 4511 1747 4545
rect 1747 4511 1765 4545
rect 1803 4511 1815 4545
rect 1815 4511 1837 4545
rect 1875 4511 1883 4545
rect 1883 4511 1909 4545
rect 1947 4511 1951 4545
rect 1951 4511 1981 4545
rect 2019 4511 2053 4545
rect 2091 4511 2121 4545
rect 2121 4511 2125 4545
rect 2163 4511 2189 4545
rect 2189 4511 2197 4545
rect 2235 4511 2257 4545
rect 2257 4511 2269 4545
rect 2307 4511 2325 4545
rect 2325 4511 2341 4545
rect 2379 4511 2393 4545
rect 2393 4511 2413 4545
rect 2451 4511 2461 4545
rect 2461 4511 2485 4545
rect 2523 4511 2529 4545
rect 2529 4511 2557 4545
rect 2595 4511 2597 4545
rect 2597 4511 2629 4545
rect 2667 4511 2699 4545
rect 2699 4511 2701 4545
rect 2739 4511 2767 4545
rect 2767 4511 2773 4545
rect 2811 4511 2835 4545
rect 2835 4511 2845 4545
rect 2883 4511 2903 4545
rect 2903 4511 2917 4545
rect 2955 4511 2971 4545
rect 2971 4511 2989 4545
rect 3027 4511 3039 4545
rect 3039 4511 3061 4545
rect 3099 4511 3107 4545
rect 3107 4511 3133 4545
rect 3171 4511 3175 4545
rect 3175 4511 3205 4545
rect 3243 4511 3277 4545
rect 3315 4511 3345 4545
rect 3345 4511 3349 4545
rect 3387 4511 3413 4545
rect 3413 4511 3421 4545
rect 3459 4511 3481 4545
rect 3481 4511 3493 4545
rect 3531 4511 3549 4545
rect 3549 4511 3565 4545
rect 3603 4511 3617 4545
rect 3617 4511 3637 4545
rect 3675 4511 3685 4545
rect 3685 4511 3709 4545
rect 3747 4511 3753 4545
rect 3753 4511 3781 4545
rect 3819 4511 3821 4545
rect 3821 4511 3853 4545
rect 3891 4511 3923 4545
rect 3923 4511 3925 4545
rect 3963 4511 3991 4545
rect 3991 4511 3997 4545
rect 4035 4511 4059 4545
rect 4059 4511 4069 4545
rect 4107 4511 4127 4545
rect 4127 4511 4141 4545
rect 4179 4511 4195 4545
rect 4195 4511 4213 4545
rect 4251 4511 4263 4545
rect 4263 4511 4285 4545
rect 4323 4511 4331 4545
rect 4331 4511 4357 4545
rect 4395 4511 4399 4545
rect 4399 4511 4429 4545
rect 4467 4511 4501 4545
rect 4539 4511 4569 4545
rect 4569 4511 4573 4545
rect 4611 4511 4637 4545
rect 4637 4511 4645 4545
rect 4683 4511 4705 4545
rect 4705 4511 4717 4545
rect 4755 4511 4773 4545
rect 4773 4511 4789 4545
rect 4827 4511 4841 4545
rect 4841 4511 4861 4545
rect 4899 4511 4909 4545
rect 4909 4511 4933 4545
rect 4971 4511 4977 4545
rect 4977 4511 5005 4545
rect 5043 4511 5045 4545
rect 5045 4511 5077 4545
rect 5115 4511 5147 4545
rect 5147 4511 5149 4545
rect 5187 4511 5215 4545
rect 5215 4511 5221 4545
rect 5259 4511 5293 4545
rect -4893 4175 -4859 4209
rect -4821 4175 -4815 4209
rect -4815 4175 -4787 4209
rect -4749 4175 -4747 4209
rect -4747 4175 -4715 4209
rect -4677 4175 -4645 4209
rect -4645 4175 -4643 4209
rect -4605 4175 -4577 4209
rect -4577 4175 -4571 4209
rect -4533 4175 -4509 4209
rect -4509 4175 -4499 4209
rect -4461 4175 -4441 4209
rect -4441 4175 -4427 4209
rect -4389 4175 -4373 4209
rect -4373 4175 -4355 4209
rect -4317 4175 -4305 4209
rect -4305 4175 -4283 4209
rect -4245 4175 -4237 4209
rect -4237 4175 -4211 4209
rect -4173 4175 -4169 4209
rect -4169 4175 -4139 4209
rect -4101 4175 -4067 4209
rect -4029 4175 -3999 4209
rect -3999 4175 -3995 4209
rect -3957 4175 -3931 4209
rect -3931 4175 -3923 4209
rect -3885 4175 -3863 4209
rect -3863 4175 -3851 4209
rect -3813 4175 -3795 4209
rect -3795 4175 -3779 4209
rect -3741 4175 -3727 4209
rect -3727 4175 -3707 4209
rect -3669 4175 -3659 4209
rect -3659 4175 -3635 4209
rect -3597 4175 -3591 4209
rect -3591 4175 -3563 4209
rect -3525 4175 -3523 4209
rect -3523 4175 -3491 4209
rect -3453 4175 -3421 4209
rect -3421 4175 -3419 4209
rect -3381 4175 -3353 4209
rect -3353 4175 -3347 4209
rect -3309 4175 -3285 4209
rect -3285 4175 -3275 4209
rect -3237 4175 -3217 4209
rect -3217 4175 -3203 4209
rect -3165 4175 -3149 4209
rect -3149 4175 -3131 4209
rect -3093 4175 -3081 4209
rect -3081 4175 -3059 4209
rect -3021 4175 -3013 4209
rect -3013 4175 -2987 4209
rect -2949 4175 -2945 4209
rect -2945 4175 -2915 4209
rect -2877 4175 -2843 4209
rect -2805 4175 -2775 4209
rect -2775 4175 -2771 4209
rect -2733 4175 -2707 4209
rect -2707 4175 -2699 4209
rect -2661 4175 -2639 4209
rect -2639 4175 -2627 4209
rect -2589 4175 -2571 4209
rect -2571 4175 -2555 4209
rect -2517 4175 -2503 4209
rect -2503 4175 -2483 4209
rect -2445 4175 -2435 4209
rect -2435 4175 -2411 4209
rect -2373 4175 -2367 4209
rect -2367 4175 -2339 4209
rect -2301 4175 -2299 4209
rect -2299 4175 -2267 4209
rect -2229 4175 -2197 4209
rect -2197 4175 -2195 4209
rect -2157 4175 -2129 4209
rect -2129 4175 -2123 4209
rect -2085 4175 -2061 4209
rect -2061 4175 -2051 4209
rect -2013 4175 -1993 4209
rect -1993 4175 -1979 4209
rect -1941 4175 -1925 4209
rect -1925 4175 -1907 4209
rect -1869 4175 -1857 4209
rect -1857 4175 -1835 4209
rect -1797 4175 -1789 4209
rect -1789 4175 -1763 4209
rect -1725 4175 -1721 4209
rect -1721 4175 -1691 4209
rect -1653 4175 -1619 4209
rect -1581 4175 -1551 4209
rect -1551 4175 -1547 4209
rect -1509 4175 -1483 4209
rect -1483 4175 -1475 4209
rect -1437 4175 -1415 4209
rect -1415 4175 -1403 4209
rect -1365 4175 -1347 4209
rect -1347 4175 -1331 4209
rect -1293 4175 -1279 4209
rect -1279 4175 -1259 4209
rect -1221 4175 -1211 4209
rect -1211 4175 -1187 4209
rect -1149 4175 -1143 4209
rect -1143 4175 -1115 4209
rect -1077 4175 -1075 4209
rect -1075 4175 -1043 4209
rect -1005 4175 -973 4209
rect -973 4175 -971 4209
rect -933 4175 -905 4209
rect -905 4175 -899 4209
rect -861 4175 -837 4209
rect -837 4175 -827 4209
rect -789 4175 -769 4209
rect -769 4175 -755 4209
rect -717 4175 -701 4209
rect -701 4175 -683 4209
rect -645 4175 -633 4209
rect -633 4175 -611 4209
rect -573 4175 -565 4209
rect -565 4175 -539 4209
rect -501 4175 -497 4209
rect -497 4175 -467 4209
rect -429 4175 -395 4209
rect -357 4175 -327 4209
rect -327 4175 -323 4209
rect -285 4175 -259 4209
rect -259 4175 -251 4209
rect -213 4175 -191 4209
rect -191 4175 -179 4209
rect -141 4175 -123 4209
rect -123 4175 -107 4209
rect -69 4175 -55 4209
rect -55 4175 -35 4209
rect 3 4175 13 4209
rect 13 4175 37 4209
rect 75 4175 81 4209
rect 81 4175 109 4209
rect 147 4175 149 4209
rect 149 4175 181 4209
rect 219 4175 251 4209
rect 251 4175 253 4209
rect 291 4175 319 4209
rect 319 4175 325 4209
rect 363 4175 387 4209
rect 387 4175 397 4209
rect 435 4175 455 4209
rect 455 4175 469 4209
rect 507 4175 523 4209
rect 523 4175 541 4209
rect 579 4175 591 4209
rect 591 4175 613 4209
rect 651 4175 659 4209
rect 659 4175 685 4209
rect 723 4175 727 4209
rect 727 4175 757 4209
rect 795 4175 829 4209
rect 867 4175 897 4209
rect 897 4175 901 4209
rect 939 4175 965 4209
rect 965 4175 973 4209
rect 1011 4175 1033 4209
rect 1033 4175 1045 4209
rect 1083 4175 1101 4209
rect 1101 4175 1117 4209
rect 1155 4175 1169 4209
rect 1169 4175 1189 4209
rect 1227 4175 1237 4209
rect 1237 4175 1261 4209
rect 1299 4175 1305 4209
rect 1305 4175 1333 4209
rect 1371 4175 1373 4209
rect 1373 4175 1405 4209
rect 1443 4175 1475 4209
rect 1475 4175 1477 4209
rect 1515 4175 1543 4209
rect 1543 4175 1549 4209
rect 1587 4175 1611 4209
rect 1611 4175 1621 4209
rect 1659 4175 1679 4209
rect 1679 4175 1693 4209
rect 1731 4175 1747 4209
rect 1747 4175 1765 4209
rect 1803 4175 1815 4209
rect 1815 4175 1837 4209
rect 1875 4175 1883 4209
rect 1883 4175 1909 4209
rect 1947 4175 1951 4209
rect 1951 4175 1981 4209
rect 2019 4175 2053 4209
rect 2091 4175 2121 4209
rect 2121 4175 2125 4209
rect 2163 4175 2189 4209
rect 2189 4175 2197 4209
rect 2235 4175 2257 4209
rect 2257 4175 2269 4209
rect 2307 4175 2325 4209
rect 2325 4175 2341 4209
rect 2379 4175 2393 4209
rect 2393 4175 2413 4209
rect 2451 4175 2461 4209
rect 2461 4175 2485 4209
rect 2523 4175 2529 4209
rect 2529 4175 2557 4209
rect 2595 4175 2597 4209
rect 2597 4175 2629 4209
rect 2667 4175 2699 4209
rect 2699 4175 2701 4209
rect 2739 4175 2767 4209
rect 2767 4175 2773 4209
rect 2811 4175 2835 4209
rect 2835 4175 2845 4209
rect 2883 4175 2903 4209
rect 2903 4175 2917 4209
rect 2955 4175 2971 4209
rect 2971 4175 2989 4209
rect 3027 4175 3039 4209
rect 3039 4175 3061 4209
rect 3099 4175 3107 4209
rect 3107 4175 3133 4209
rect 3171 4175 3175 4209
rect 3175 4175 3205 4209
rect 3243 4175 3277 4209
rect 3315 4175 3345 4209
rect 3345 4175 3349 4209
rect 3387 4175 3413 4209
rect 3413 4175 3421 4209
rect 3459 4175 3481 4209
rect 3481 4175 3493 4209
rect 3531 4175 3549 4209
rect 3549 4175 3565 4209
rect 3603 4175 3617 4209
rect 3617 4175 3637 4209
rect 3675 4175 3685 4209
rect 3685 4175 3709 4209
rect 3747 4175 3753 4209
rect 3753 4175 3781 4209
rect 3819 4175 3821 4209
rect 3821 4175 3853 4209
rect 3891 4175 3923 4209
rect 3923 4175 3925 4209
rect 3963 4175 3991 4209
rect 3991 4175 3997 4209
rect 4035 4175 4059 4209
rect 4059 4175 4069 4209
rect 4107 4175 4127 4209
rect 4127 4175 4141 4209
rect 4179 4175 4195 4209
rect 4195 4175 4213 4209
rect 4251 4175 4263 4209
rect 4263 4175 4285 4209
rect 4323 4175 4331 4209
rect 4331 4175 4357 4209
rect 4395 4175 4399 4209
rect 4399 4175 4429 4209
rect 4467 4175 4501 4209
rect 4539 4175 4569 4209
rect 4569 4175 4573 4209
rect 4611 4175 4637 4209
rect 4637 4175 4645 4209
rect 4683 4175 4705 4209
rect 4705 4175 4717 4209
rect 4755 4175 4773 4209
rect 4773 4175 4789 4209
rect 4827 4175 4841 4209
rect 4841 4175 4861 4209
rect 4899 4175 4909 4209
rect 4909 4175 4933 4209
rect 4971 4175 4977 4209
rect 4977 4175 5005 4209
rect 5043 4175 5045 4209
rect 5045 4175 5077 4209
rect 5115 4175 5147 4209
rect 5147 4175 5149 4209
rect 5187 4175 5215 4209
rect 5215 4175 5221 4209
rect 5259 4175 5293 4209
rect -4989 3979 -4955 3999
rect -4989 3965 -4955 3979
rect -4989 3911 -4955 3927
rect -4989 3893 -4955 3911
rect -4989 3843 -4955 3855
rect -4989 3821 -4955 3843
rect -4989 3775 -4955 3783
rect -4989 3749 -4955 3775
rect -4989 3707 -4955 3711
rect -4989 3677 -4955 3707
rect -4989 3605 -4955 3639
rect -4989 3537 -4955 3567
rect -4989 3533 -4955 3537
rect -4989 3469 -4955 3495
rect -4989 3461 -4955 3469
rect -4989 3401 -4955 3423
rect -4989 3389 -4955 3401
rect -4989 3333 -4955 3351
rect -4989 3317 -4955 3333
rect -4989 3265 -4955 3279
rect -4989 3245 -4955 3265
rect -4989 3197 -4955 3207
rect -4989 3173 -4955 3197
rect -4989 3129 -4955 3135
rect -4989 3101 -4955 3129
rect -4989 3061 -4955 3063
rect -4989 3029 -4955 3061
rect -4989 2959 -4955 2991
rect -4989 2957 -4955 2959
rect -4989 2891 -4955 2919
rect -4989 2885 -4955 2891
rect -4989 2823 -4955 2847
rect -4989 2813 -4955 2823
rect -4989 2755 -4955 2775
rect -4989 2741 -4955 2755
rect -4989 2687 -4955 2703
rect -4989 2669 -4955 2687
rect -4989 2619 -4955 2631
rect -4989 2597 -4955 2619
rect -4989 2551 -4955 2559
rect -4989 2525 -4955 2551
rect -4989 2483 -4955 2487
rect -4989 2453 -4955 2483
rect -4989 2381 -4955 2415
rect -4989 2313 -4955 2343
rect -4989 2309 -4955 2313
rect -4989 2245 -4955 2271
rect -4989 2237 -4955 2245
rect -4989 2177 -4955 2199
rect -4989 2165 -4955 2177
rect -4989 2109 -4955 2127
rect -4989 2093 -4955 2109
rect -4989 2041 -4955 2055
rect -4989 2021 -4955 2041
rect 5355 3979 5389 3999
rect 5355 3965 5389 3979
rect 5355 3911 5389 3927
rect 5355 3893 5389 3911
rect 5355 3843 5389 3855
rect 5355 3821 5389 3843
rect 5355 3775 5389 3783
rect 5355 3749 5389 3775
rect 5355 3707 5389 3711
rect 5355 3677 5389 3707
rect 5355 3605 5389 3639
rect 5355 3537 5389 3567
rect 5355 3533 5389 3537
rect 5355 3469 5389 3495
rect 5355 3461 5389 3469
rect 5355 3401 5389 3423
rect 5355 3389 5389 3401
rect 5355 3333 5389 3351
rect 5355 3317 5389 3333
rect 5355 3265 5389 3279
rect 5355 3245 5389 3265
rect 5355 3197 5389 3207
rect 5355 3173 5389 3197
rect 5355 3129 5389 3135
rect 5355 3101 5389 3129
rect 5355 3061 5389 3063
rect 5355 3029 5389 3061
rect 5355 2959 5389 2991
rect 5355 2957 5389 2959
rect 5355 2891 5389 2919
rect 5355 2885 5389 2891
rect 5355 2823 5389 2847
rect 5355 2813 5389 2823
rect 5355 2755 5389 2775
rect 5355 2741 5389 2755
rect 5355 2687 5389 2703
rect 5355 2669 5389 2687
rect 5355 2619 5389 2631
rect 5355 2597 5389 2619
rect 5355 2551 5389 2559
rect 5355 2525 5389 2551
rect 5355 2483 5389 2487
rect 5355 2453 5389 2483
rect 5355 2381 5389 2415
rect 5355 2313 5389 2343
rect 5355 2309 5389 2313
rect 5355 2245 5389 2271
rect 5355 2237 5389 2245
rect 5355 2177 5389 2199
rect 5355 2165 5389 2177
rect 5355 2109 5389 2127
rect 5355 2093 5389 2109
rect 5355 2041 5389 2055
rect 5355 2021 5389 2041
rect -4893 1811 -4859 1845
rect -4821 1811 -4815 1845
rect -4815 1811 -4787 1845
rect -4749 1811 -4747 1845
rect -4747 1811 -4715 1845
rect -4677 1811 -4645 1845
rect -4645 1811 -4643 1845
rect -4605 1811 -4577 1845
rect -4577 1811 -4571 1845
rect -4533 1811 -4509 1845
rect -4509 1811 -4499 1845
rect -4461 1811 -4441 1845
rect -4441 1811 -4427 1845
rect -4389 1811 -4373 1845
rect -4373 1811 -4355 1845
rect -4317 1811 -4305 1845
rect -4305 1811 -4283 1845
rect -4245 1811 -4237 1845
rect -4237 1811 -4211 1845
rect -4173 1811 -4169 1845
rect -4169 1811 -4139 1845
rect -4101 1811 -4067 1845
rect -4029 1811 -3999 1845
rect -3999 1811 -3995 1845
rect -3957 1811 -3931 1845
rect -3931 1811 -3923 1845
rect -3885 1811 -3863 1845
rect -3863 1811 -3851 1845
rect -3813 1811 -3795 1845
rect -3795 1811 -3779 1845
rect -3741 1811 -3727 1845
rect -3727 1811 -3707 1845
rect -3669 1811 -3659 1845
rect -3659 1811 -3635 1845
rect -3597 1811 -3591 1845
rect -3591 1811 -3563 1845
rect -3525 1811 -3523 1845
rect -3523 1811 -3491 1845
rect -3453 1811 -3421 1845
rect -3421 1811 -3419 1845
rect -3381 1811 -3353 1845
rect -3353 1811 -3347 1845
rect -3309 1811 -3285 1845
rect -3285 1811 -3275 1845
rect -3237 1811 -3217 1845
rect -3217 1811 -3203 1845
rect -3165 1811 -3149 1845
rect -3149 1811 -3131 1845
rect -3093 1811 -3081 1845
rect -3081 1811 -3059 1845
rect -3021 1811 -3013 1845
rect -3013 1811 -2987 1845
rect -2949 1811 -2945 1845
rect -2945 1811 -2915 1845
rect -2877 1811 -2843 1845
rect -2805 1811 -2775 1845
rect -2775 1811 -2771 1845
rect -2733 1811 -2707 1845
rect -2707 1811 -2699 1845
rect -2661 1811 -2639 1845
rect -2639 1811 -2627 1845
rect -2589 1811 -2571 1845
rect -2571 1811 -2555 1845
rect -2517 1811 -2503 1845
rect -2503 1811 -2483 1845
rect -2445 1811 -2435 1845
rect -2435 1811 -2411 1845
rect -2373 1811 -2367 1845
rect -2367 1811 -2339 1845
rect -2301 1811 -2299 1845
rect -2299 1811 -2267 1845
rect -2229 1811 -2197 1845
rect -2197 1811 -2195 1845
rect -2157 1811 -2129 1845
rect -2129 1811 -2123 1845
rect -2085 1811 -2061 1845
rect -2061 1811 -2051 1845
rect -2013 1811 -1993 1845
rect -1993 1811 -1979 1845
rect -1941 1811 -1925 1845
rect -1925 1811 -1907 1845
rect -1869 1811 -1857 1845
rect -1857 1811 -1835 1845
rect -1797 1811 -1789 1845
rect -1789 1811 -1763 1845
rect -1725 1811 -1721 1845
rect -1721 1811 -1691 1845
rect -1653 1811 -1619 1845
rect -1581 1811 -1551 1845
rect -1551 1811 -1547 1845
rect -1509 1811 -1483 1845
rect -1483 1811 -1475 1845
rect -1437 1811 -1415 1845
rect -1415 1811 -1403 1845
rect -1365 1811 -1347 1845
rect -1347 1811 -1331 1845
rect -1293 1811 -1279 1845
rect -1279 1811 -1259 1845
rect -1221 1811 -1211 1845
rect -1211 1811 -1187 1845
rect -1149 1811 -1143 1845
rect -1143 1811 -1115 1845
rect -1077 1811 -1075 1845
rect -1075 1811 -1043 1845
rect -1005 1811 -973 1845
rect -973 1811 -971 1845
rect -933 1811 -905 1845
rect -905 1811 -899 1845
rect -861 1811 -837 1845
rect -837 1811 -827 1845
rect -789 1811 -769 1845
rect -769 1811 -755 1845
rect -717 1811 -701 1845
rect -701 1811 -683 1845
rect -645 1811 -633 1845
rect -633 1811 -611 1845
rect -573 1811 -565 1845
rect -565 1811 -539 1845
rect -501 1811 -497 1845
rect -497 1811 -467 1845
rect -429 1811 -395 1845
rect -357 1811 -327 1845
rect -327 1811 -323 1845
rect -285 1811 -259 1845
rect -259 1811 -251 1845
rect -213 1811 -191 1845
rect -191 1811 -179 1845
rect -141 1811 -123 1845
rect -123 1811 -107 1845
rect -69 1811 -55 1845
rect -55 1811 -35 1845
rect 3 1811 13 1845
rect 13 1811 37 1845
rect 75 1811 81 1845
rect 81 1811 109 1845
rect 147 1811 149 1845
rect 149 1811 181 1845
rect 219 1811 251 1845
rect 251 1811 253 1845
rect 291 1811 319 1845
rect 319 1811 325 1845
rect 363 1811 387 1845
rect 387 1811 397 1845
rect 435 1811 455 1845
rect 455 1811 469 1845
rect 507 1811 523 1845
rect 523 1811 541 1845
rect 579 1811 591 1845
rect 591 1811 613 1845
rect 651 1811 659 1845
rect 659 1811 685 1845
rect 723 1811 727 1845
rect 727 1811 757 1845
rect 795 1811 829 1845
rect 867 1811 897 1845
rect 897 1811 901 1845
rect 939 1811 965 1845
rect 965 1811 973 1845
rect 1011 1811 1033 1845
rect 1033 1811 1045 1845
rect 1083 1811 1101 1845
rect 1101 1811 1117 1845
rect 1155 1811 1169 1845
rect 1169 1811 1189 1845
rect 1227 1811 1237 1845
rect 1237 1811 1261 1845
rect 1299 1811 1305 1845
rect 1305 1811 1333 1845
rect 1371 1811 1373 1845
rect 1373 1811 1405 1845
rect 1443 1811 1475 1845
rect 1475 1811 1477 1845
rect 1515 1811 1543 1845
rect 1543 1811 1549 1845
rect 1587 1811 1611 1845
rect 1611 1811 1621 1845
rect 1659 1811 1679 1845
rect 1679 1811 1693 1845
rect 1731 1811 1747 1845
rect 1747 1811 1765 1845
rect 1803 1811 1815 1845
rect 1815 1811 1837 1845
rect 1875 1811 1883 1845
rect 1883 1811 1909 1845
rect 1947 1811 1951 1845
rect 1951 1811 1981 1845
rect 2019 1811 2053 1845
rect 2091 1811 2121 1845
rect 2121 1811 2125 1845
rect 2163 1811 2189 1845
rect 2189 1811 2197 1845
rect 2235 1811 2257 1845
rect 2257 1811 2269 1845
rect 2307 1811 2325 1845
rect 2325 1811 2341 1845
rect 2379 1811 2393 1845
rect 2393 1811 2413 1845
rect 2451 1811 2461 1845
rect 2461 1811 2485 1845
rect 2523 1811 2529 1845
rect 2529 1811 2557 1845
rect 2595 1811 2597 1845
rect 2597 1811 2629 1845
rect 2667 1811 2699 1845
rect 2699 1811 2701 1845
rect 2739 1811 2767 1845
rect 2767 1811 2773 1845
rect 2811 1811 2835 1845
rect 2835 1811 2845 1845
rect 2883 1811 2903 1845
rect 2903 1811 2917 1845
rect 2955 1811 2971 1845
rect 2971 1811 2989 1845
rect 3027 1811 3039 1845
rect 3039 1811 3061 1845
rect 3099 1811 3107 1845
rect 3107 1811 3133 1845
rect 3171 1811 3175 1845
rect 3175 1811 3205 1845
rect 3243 1811 3277 1845
rect 3315 1811 3345 1845
rect 3345 1811 3349 1845
rect 3387 1811 3413 1845
rect 3413 1811 3421 1845
rect 3459 1811 3481 1845
rect 3481 1811 3493 1845
rect 3531 1811 3549 1845
rect 3549 1811 3565 1845
rect 3603 1811 3617 1845
rect 3617 1811 3637 1845
rect 3675 1811 3685 1845
rect 3685 1811 3709 1845
rect 3747 1811 3753 1845
rect 3753 1811 3781 1845
rect 3819 1811 3821 1845
rect 3821 1811 3853 1845
rect 3891 1811 3923 1845
rect 3923 1811 3925 1845
rect 3963 1811 3991 1845
rect 3991 1811 3997 1845
rect 4035 1811 4059 1845
rect 4059 1811 4069 1845
rect 4107 1811 4127 1845
rect 4127 1811 4141 1845
rect 4179 1811 4195 1845
rect 4195 1811 4213 1845
rect 4251 1811 4263 1845
rect 4263 1811 4285 1845
rect 4323 1811 4331 1845
rect 4331 1811 4357 1845
rect 4395 1811 4399 1845
rect 4399 1811 4429 1845
rect 4467 1811 4501 1845
rect 4539 1811 4569 1845
rect 4569 1811 4573 1845
rect 4611 1811 4637 1845
rect 4637 1811 4645 1845
rect 4683 1811 4705 1845
rect 4705 1811 4717 1845
rect 4755 1811 4773 1845
rect 4773 1811 4789 1845
rect 4827 1811 4841 1845
rect 4841 1811 4861 1845
rect 4899 1811 4909 1845
rect 4909 1811 4933 1845
rect 4971 1811 4977 1845
rect 4977 1811 5005 1845
rect 5043 1811 5045 1845
rect 5045 1811 5077 1845
rect 5115 1811 5147 1845
rect 5147 1811 5149 1845
rect 5187 1811 5215 1845
rect 5215 1811 5221 1845
rect 5259 1811 5293 1845
<< metal1 >>
rect -5028 10289 5428 10328
rect -5028 10255 -4893 10289
rect -4859 10255 -4821 10289
rect -4787 10255 -4749 10289
rect -4715 10255 -4677 10289
rect -4643 10255 -4605 10289
rect -4571 10255 -4533 10289
rect -4499 10255 -4461 10289
rect -4427 10255 -4389 10289
rect -4355 10255 -4317 10289
rect -4283 10255 -4245 10289
rect -4211 10255 -4173 10289
rect -4139 10255 -4101 10289
rect -4067 10255 -4029 10289
rect -3995 10255 -3957 10289
rect -3923 10255 -3885 10289
rect -3851 10255 -3813 10289
rect -3779 10255 -3741 10289
rect -3707 10255 -3669 10289
rect -3635 10255 -3597 10289
rect -3563 10255 -3525 10289
rect -3491 10255 -3453 10289
rect -3419 10255 -3381 10289
rect -3347 10255 -3309 10289
rect -3275 10255 -3237 10289
rect -3203 10255 -3165 10289
rect -3131 10255 -3093 10289
rect -3059 10255 -3021 10289
rect -2987 10255 -2949 10289
rect -2915 10255 -2877 10289
rect -2843 10255 -2805 10289
rect -2771 10255 -2733 10289
rect -2699 10255 -2661 10289
rect -2627 10255 -2589 10289
rect -2555 10255 -2517 10289
rect -2483 10255 -2445 10289
rect -2411 10255 -2373 10289
rect -2339 10255 -2301 10289
rect -2267 10255 -2229 10289
rect -2195 10255 -2157 10289
rect -2123 10255 -2085 10289
rect -2051 10255 -2013 10289
rect -1979 10255 -1941 10289
rect -1907 10255 -1869 10289
rect -1835 10255 -1797 10289
rect -1763 10255 -1725 10289
rect -1691 10255 -1653 10289
rect -1619 10255 -1581 10289
rect -1547 10255 -1509 10289
rect -1475 10255 -1437 10289
rect -1403 10255 -1365 10289
rect -1331 10255 -1293 10289
rect -1259 10255 -1221 10289
rect -1187 10255 -1149 10289
rect -1115 10255 -1077 10289
rect -1043 10255 -1005 10289
rect -971 10255 -933 10289
rect -899 10255 -861 10289
rect -827 10255 -789 10289
rect -755 10255 -717 10289
rect -683 10255 -645 10289
rect -611 10255 -573 10289
rect -539 10255 -501 10289
rect -467 10255 -429 10289
rect -395 10255 -357 10289
rect -323 10255 -285 10289
rect -251 10255 -213 10289
rect -179 10255 -141 10289
rect -107 10255 -69 10289
rect -35 10255 3 10289
rect 37 10255 75 10289
rect 109 10255 147 10289
rect 181 10255 219 10289
rect 253 10255 291 10289
rect 325 10255 363 10289
rect 397 10255 435 10289
rect 469 10255 507 10289
rect 541 10255 579 10289
rect 613 10255 651 10289
rect 685 10255 723 10289
rect 757 10255 795 10289
rect 829 10255 867 10289
rect 901 10255 939 10289
rect 973 10255 1011 10289
rect 1045 10255 1083 10289
rect 1117 10255 1155 10289
rect 1189 10255 1227 10289
rect 1261 10255 1299 10289
rect 1333 10255 1371 10289
rect 1405 10255 1443 10289
rect 1477 10255 1515 10289
rect 1549 10255 1587 10289
rect 1621 10255 1659 10289
rect 1693 10255 1731 10289
rect 1765 10255 1803 10289
rect 1837 10255 1875 10289
rect 1909 10255 1947 10289
rect 1981 10255 2019 10289
rect 2053 10255 2091 10289
rect 2125 10255 2163 10289
rect 2197 10255 2235 10289
rect 2269 10255 2307 10289
rect 2341 10255 2379 10289
rect 2413 10255 2451 10289
rect 2485 10255 2523 10289
rect 2557 10255 2595 10289
rect 2629 10255 2667 10289
rect 2701 10255 2739 10289
rect 2773 10255 2811 10289
rect 2845 10255 2883 10289
rect 2917 10255 2955 10289
rect 2989 10255 3027 10289
rect 3061 10255 3099 10289
rect 3133 10255 3171 10289
rect 3205 10255 3243 10289
rect 3277 10255 3315 10289
rect 3349 10255 3387 10289
rect 3421 10255 3459 10289
rect 3493 10255 3531 10289
rect 3565 10255 3603 10289
rect 3637 10255 3675 10289
rect 3709 10255 3747 10289
rect 3781 10255 3819 10289
rect 3853 10255 3891 10289
rect 3925 10255 3963 10289
rect 3997 10255 4035 10289
rect 4069 10255 4107 10289
rect 4141 10255 4179 10289
rect 4213 10255 4251 10289
rect 4285 10255 4323 10289
rect 4357 10255 4395 10289
rect 4429 10255 4467 10289
rect 4501 10255 4539 10289
rect 4573 10255 4611 10289
rect 4645 10255 4683 10289
rect 4717 10255 4755 10289
rect 4789 10255 4827 10289
rect 4861 10255 4899 10289
rect 4933 10255 4971 10289
rect 5005 10255 5043 10289
rect 5077 10255 5115 10289
rect 5149 10255 5187 10289
rect 5221 10255 5259 10289
rect 5293 10255 5428 10289
rect -5028 10216 5428 10255
rect -5028 10188 -4306 10216
rect -5028 9944 -4898 10188
rect -4334 9944 -4306 10188
rect -5028 9919 -4306 9944
rect -5028 9885 -4989 9919
rect -4955 9916 -4306 9919
rect 4706 10188 5428 10216
rect 4706 9944 4734 10188
rect 5298 9944 5428 10188
rect 4706 9919 5428 9944
rect 4706 9916 5355 9919
rect -4955 9885 -4916 9916
rect -5028 9847 -4916 9885
rect -5028 9813 -4989 9847
rect -4955 9813 -4916 9847
rect -5028 9775 -4916 9813
rect -5028 9741 -4989 9775
rect -4955 9741 -4916 9775
rect 5316 9885 5355 9916
rect 5389 9885 5428 9919
rect 5316 9847 5428 9885
rect 5316 9813 5355 9847
rect 5389 9813 5428 9847
rect 5316 9775 5428 9813
rect -5028 9703 -4916 9741
rect -5028 9669 -4989 9703
rect -4955 9669 -4916 9703
rect -5028 9631 -4916 9669
rect -4078 9725 4278 9756
rect -4078 9673 -4042 9725
rect -3990 9673 -3442 9725
rect -3390 9673 -2842 9725
rect -2790 9673 -2242 9725
rect -2190 9673 -1642 9725
rect -1590 9673 -1042 9725
rect -990 9673 -442 9725
rect -390 9673 158 9725
rect 210 9673 758 9725
rect 810 9673 1358 9725
rect 1410 9673 1958 9725
rect 2010 9673 2558 9725
rect 2610 9673 3158 9725
rect 3210 9673 3758 9725
rect 3810 9673 4178 9725
rect 4230 9673 4278 9725
rect -4078 9646 4278 9673
rect 5316 9741 5355 9775
rect 5389 9741 5428 9775
rect 5316 9703 5428 9741
rect 5316 9669 5355 9703
rect 5389 9669 5428 9703
rect -5028 9597 -4989 9631
rect -4955 9597 -4916 9631
rect -5028 9559 -4916 9597
rect -5028 9525 -4989 9559
rect -4955 9525 -4916 9559
rect -5028 9487 -4916 9525
rect -5028 9453 -4989 9487
rect -4955 9453 -4916 9487
rect -5028 9415 -4916 9453
rect -5028 9381 -4989 9415
rect -4955 9381 -4916 9415
rect -5028 9343 -4916 9381
rect -5028 9309 -4989 9343
rect -4955 9309 -4916 9343
rect -5028 9271 -4916 9309
rect -5028 9237 -4989 9271
rect -4955 9237 -4916 9271
rect -5028 9199 -4916 9237
rect -5028 9165 -4989 9199
rect -4955 9165 -4916 9199
rect -5028 9127 -4916 9165
rect -5028 9093 -4989 9127
rect -4955 9093 -4916 9127
rect -5028 9055 -4916 9093
rect -5028 9021 -4989 9055
rect -4955 9021 -4916 9055
rect -5028 8983 -4916 9021
rect -5028 8949 -4989 8983
rect -4955 8949 -4916 8983
rect -5028 8911 -4916 8949
rect -5028 8877 -4989 8911
rect -4955 8877 -4916 8911
rect -5028 8839 -4916 8877
rect -5028 8805 -4989 8839
rect -4955 8805 -4916 8839
rect -4050 8826 -3990 9646
rect -3818 8918 -3758 9646
rect -5028 8767 -4916 8805
rect -3592 8794 -3532 9646
rect -2676 9392 2882 9452
rect -3366 9080 -3294 9084
rect -3366 9028 -3356 9080
rect -3304 9028 -3294 9080
rect -3366 9024 -3294 9028
rect -2910 9080 -2838 9084
rect -2910 9028 -2900 9080
rect -2848 9028 -2838 9080
rect -2910 9024 -2838 9028
rect -3360 8916 -3300 9024
rect -2904 8918 -2844 9024
rect -2676 8800 -2616 9392
rect -1760 9258 1962 9318
rect -2450 9080 -2378 9084
rect -2450 9028 -2440 9080
rect -2388 9028 -2378 9080
rect -2450 9024 -2378 9028
rect -1994 9080 -1922 9084
rect -1994 9028 -1984 9080
rect -1932 9028 -1922 9080
rect -1994 9024 -1922 9028
rect -2444 8912 -2384 9024
rect -1988 8918 -1928 9024
rect -1760 8798 -1700 9258
rect -844 9134 1046 9194
rect -1536 9080 -1464 9084
rect -1536 9028 -1526 9080
rect -1474 9028 -1464 9080
rect -1536 9024 -1464 9028
rect -1072 9080 -1000 9084
rect -1072 9028 -1062 9080
rect -1010 9028 -1000 9080
rect -1072 9024 -1000 9028
rect -1530 8918 -1470 9024
rect -1066 8914 -1006 9024
rect -844 8780 -784 9134
rect -622 9080 -550 9084
rect -622 9028 -612 9080
rect -560 9028 -550 9080
rect -622 9024 -550 9028
rect -166 9080 -94 9084
rect -166 9028 -156 9080
rect -104 9028 -94 9080
rect -166 9024 -94 9028
rect 302 9080 374 9084
rect 302 9028 312 9080
rect 364 9028 374 9080
rect 302 9024 374 9028
rect 760 9080 832 9084
rect 760 9028 770 9080
rect 822 9028 832 9080
rect 760 9024 832 9028
rect -616 8920 -556 9024
rect -160 8920 -100 9024
rect 308 8920 368 9024
rect 766 8924 826 9024
rect 986 8814 1046 9134
rect 1216 9080 1288 9084
rect 1216 9028 1226 9080
rect 1278 9028 1288 9080
rect 1216 9024 1288 9028
rect 1672 9080 1744 9084
rect 1672 9028 1682 9080
rect 1734 9028 1744 9080
rect 1672 9024 1744 9028
rect 1222 8918 1282 9024
rect 1678 8918 1738 9024
rect 1902 8800 1962 9258
rect 2128 9080 2200 9084
rect 2128 9028 2138 9080
rect 2190 9028 2200 9080
rect 2128 9024 2200 9028
rect 2584 9080 2656 9084
rect 2584 9028 2594 9080
rect 2646 9028 2656 9080
rect 2584 9024 2656 9028
rect 2134 8918 2194 9024
rect 2590 8922 2650 9024
rect 2822 8802 2882 9392
rect 3042 9080 3114 9084
rect 3042 9028 3052 9080
rect 3104 9028 3114 9080
rect 3042 9024 3114 9028
rect 3502 9080 3574 9084
rect 3502 9028 3512 9080
rect 3564 9028 3574 9080
rect 3502 9024 3574 9028
rect 3048 8918 3108 9024
rect 3508 8914 3568 9024
rect 3738 8782 3798 9646
rect 3968 8916 4028 9646
rect 4196 8788 4256 9646
rect 5316 9631 5428 9669
rect 5316 9597 5355 9631
rect 5389 9597 5428 9631
rect 5316 9559 5428 9597
rect 5316 9525 5355 9559
rect 5389 9525 5428 9559
rect 5316 9487 5428 9525
rect 5316 9453 5355 9487
rect 5389 9453 5428 9487
rect 5316 9415 5428 9453
rect 5316 9381 5355 9415
rect 5389 9381 5428 9415
rect 5316 9343 5428 9381
rect 5316 9309 5355 9343
rect 5389 9309 5428 9343
rect 5316 9271 5428 9309
rect 5316 9237 5355 9271
rect 5389 9237 5428 9271
rect 5316 9199 5428 9237
rect 5316 9165 5355 9199
rect 5389 9165 5428 9199
rect 5316 9127 5428 9165
rect 5316 9093 5355 9127
rect 5389 9093 5428 9127
rect 5316 9055 5428 9093
rect 5316 9021 5355 9055
rect 5389 9021 5428 9055
rect 5316 8983 5428 9021
rect 5316 8949 5355 8983
rect 5389 8949 5428 8983
rect 5316 8911 5428 8949
rect 5316 8877 5355 8911
rect 5389 8877 5428 8911
rect 5316 8839 5428 8877
rect 5316 8805 5355 8839
rect 5389 8805 5428 8839
rect -5028 8733 -4989 8767
rect -4955 8733 -4916 8767
rect -5028 8695 -4916 8733
rect -5028 8661 -4989 8695
rect -4955 8661 -4916 8695
rect -5028 8623 -4916 8661
rect -5028 8589 -4989 8623
rect -4955 8589 -4916 8623
rect -5028 8551 -4916 8589
rect -5028 8517 -4989 8551
rect -4955 8517 -4916 8551
rect -5028 8479 -4916 8517
rect -5028 8445 -4989 8479
rect -4955 8445 -4916 8479
rect -5028 8407 -4916 8445
rect -5028 8373 -4989 8407
rect -4955 8373 -4916 8407
rect -5028 8335 -4916 8373
rect -5028 8301 -4989 8335
rect -4955 8301 -4916 8335
rect -5028 8263 -4916 8301
rect -5028 8229 -4989 8263
rect -4955 8229 -4916 8263
rect -5028 8191 -4916 8229
rect -5028 8157 -4989 8191
rect -4955 8157 -4916 8191
rect -5028 8119 -4916 8157
rect -5028 8085 -4989 8119
rect -4955 8085 -4916 8119
rect -5028 8047 -4916 8085
rect -5028 8013 -4989 8047
rect -4955 8013 -4916 8047
rect -5028 7975 -4916 8013
rect -5028 7941 -4989 7975
rect -4955 7941 -4916 7975
rect -5028 7903 -4916 7941
rect -5028 7869 -4989 7903
rect -4955 7869 -4916 7903
rect -5028 7831 -4916 7869
rect -5028 7797 -4989 7831
rect -4955 7797 -4916 7831
rect -5028 7759 -4916 7797
rect -5028 7725 -4989 7759
rect -4955 7725 -4916 7759
rect -5028 7687 -4916 7725
rect -5028 7653 -4989 7687
rect -4955 7653 -4916 7687
rect -5028 7615 -4916 7653
rect -5028 7581 -4989 7615
rect -4955 7581 -4916 7615
rect -5028 7543 -4916 7581
rect -5028 7509 -4989 7543
rect -4955 7509 -4916 7543
rect -5028 7471 -4916 7509
rect -5028 7437 -4989 7471
rect -4955 7437 -4916 7471
rect -5028 7399 -4916 7437
rect -5028 7365 -4989 7399
rect -4955 7365 -4916 7399
rect 5316 8767 5428 8805
rect 5316 8733 5355 8767
rect 5389 8733 5428 8767
rect 5316 8695 5428 8733
rect 5316 8661 5355 8695
rect 5389 8661 5428 8695
rect 5316 8623 5428 8661
rect 5316 8589 5355 8623
rect 5389 8589 5428 8623
rect 5316 8551 5428 8589
rect 5316 8517 5355 8551
rect 5389 8517 5428 8551
rect 5316 8479 5428 8517
rect 5316 8445 5355 8479
rect 5389 8445 5428 8479
rect 5316 8407 5428 8445
rect 5316 8373 5355 8407
rect 5389 8373 5428 8407
rect 5316 8335 5428 8373
rect 5316 8301 5355 8335
rect 5389 8301 5428 8335
rect 5316 8263 5428 8301
rect 5316 8229 5355 8263
rect 5389 8229 5428 8263
rect 5316 8191 5428 8229
rect 5316 8157 5355 8191
rect 5389 8157 5428 8191
rect 5316 8119 5428 8157
rect 5316 8085 5355 8119
rect 5389 8085 5428 8119
rect 5316 8047 5428 8085
rect 5316 8013 5355 8047
rect 5389 8013 5428 8047
rect 5316 7975 5428 8013
rect 5316 7941 5355 7975
rect 5389 7941 5428 7975
rect 5316 7903 5428 7941
rect 5316 7869 5355 7903
rect 5389 7869 5428 7903
rect 5316 7831 5428 7869
rect 5316 7797 5355 7831
rect 5389 7797 5428 7831
rect 5316 7759 5428 7797
rect 5316 7725 5355 7759
rect 5389 7725 5428 7759
rect 5316 7687 5428 7725
rect 5316 7653 5355 7687
rect 5389 7653 5428 7687
rect 5316 7615 5428 7653
rect 5316 7581 5355 7615
rect 5389 7581 5428 7615
rect 5316 7543 5428 7581
rect 5316 7509 5355 7543
rect 5389 7509 5428 7543
rect 5316 7471 5428 7509
rect 5316 7437 5355 7471
rect 5389 7437 5428 7471
rect 5316 7399 5428 7437
rect -5028 7327 -4916 7365
rect -5028 7293 -4989 7327
rect -4955 7293 -4916 7327
rect -5028 7255 -4916 7293
rect -5028 7221 -4989 7255
rect -4955 7221 -4916 7255
rect -5028 7183 -4916 7221
rect -5028 7149 -4989 7183
rect -4955 7149 -4916 7183
rect -5028 7111 -4916 7149
rect -5028 7077 -4989 7111
rect -4955 7110 -4916 7111
rect -4048 7110 -3988 7342
rect -3820 7110 -3760 7226
rect -3594 7110 -3534 7326
rect -3364 7110 -3304 7218
rect -4955 7077 -3534 7110
rect -5028 7050 -3534 7077
rect -3370 7106 -3298 7110
rect -3370 7054 -3360 7106
rect -3308 7054 -3298 7106
rect -3370 7050 -3298 7054
rect -5028 7039 -4916 7050
rect -5028 7005 -4989 7039
rect -4955 7005 -4916 7039
rect -5028 6967 -4916 7005
rect -5028 6933 -4989 6967
rect -4955 6933 -4916 6967
rect -5028 6895 -4916 6933
rect -5028 6861 -4989 6895
rect -4955 6861 -4916 6895
rect -5028 6823 -4916 6861
rect -5028 6789 -4989 6823
rect -4955 6789 -4916 6823
rect -5028 6751 -4916 6789
rect -5028 6717 -4989 6751
rect -4955 6717 -4916 6751
rect -5028 6679 -4916 6717
rect -5028 6645 -4989 6679
rect -4955 6678 -4916 6679
rect -4048 6678 -3988 7050
rect -4955 6645 -3988 6678
rect -5028 6618 -3988 6645
rect -3136 6630 -3076 7366
rect 5316 7365 5355 7399
rect 5389 7365 5428 7399
rect -2908 7110 -2848 7216
rect -2448 7110 -2388 7222
rect -2914 7106 -2842 7110
rect -2914 7054 -2904 7106
rect -2852 7054 -2842 7106
rect -2914 7050 -2842 7054
rect -2454 7106 -2382 7110
rect -2454 7054 -2444 7106
rect -2392 7054 -2382 7106
rect -2454 7050 -2382 7054
rect -2218 6760 -2158 7360
rect -1992 7110 -1932 7216
rect -1534 7110 -1474 7216
rect -1998 7106 -1926 7110
rect -1998 7054 -1988 7106
rect -1936 7054 -1926 7106
rect -1998 7050 -1926 7054
rect -1540 7106 -1468 7110
rect -1540 7054 -1530 7106
rect -1478 7054 -1468 7106
rect -1540 7050 -1468 7054
rect -1310 6886 -1250 7354
rect -1070 7110 -1010 7220
rect -616 7110 -556 7222
rect -1076 7106 -1004 7110
rect -1076 7054 -1066 7106
rect -1014 7054 -1004 7106
rect -1076 7050 -1004 7054
rect -622 7106 -550 7110
rect -622 7054 -612 7106
rect -560 7054 -550 7106
rect -622 7050 -550 7054
rect -386 7002 -326 7362
rect -158 7112 -98 7220
rect 76 7118 136 7304
rect 302 7118 362 7228
rect -164 7106 -92 7112
rect -164 7054 -154 7106
rect -102 7054 -92 7106
rect 76 7066 80 7118
rect 132 7066 136 7118
rect 76 7056 136 7066
rect 290 7106 374 7118
rect -164 7050 -92 7054
rect 290 7054 306 7106
rect 358 7054 374 7106
rect 290 7046 374 7054
rect 532 7002 592 7310
rect 758 7110 818 7222
rect 1218 7110 1278 7216
rect 752 7106 824 7110
rect 752 7054 762 7106
rect 814 7054 824 7106
rect 752 7050 824 7054
rect 1212 7106 1284 7110
rect 1212 7054 1222 7106
rect 1274 7054 1284 7106
rect 1212 7050 1284 7054
rect -386 6942 592 7002
rect 1446 6886 1506 7314
rect 1674 7110 1734 7216
rect 2130 7110 2190 7216
rect 1668 7106 1740 7110
rect 1668 7054 1678 7106
rect 1730 7054 1740 7106
rect 1668 7050 1740 7054
rect 2124 7106 2196 7110
rect 2124 7054 2134 7106
rect 2186 7054 2196 7106
rect 2124 7050 2196 7054
rect -1310 6826 1506 6886
rect 2366 6760 2426 7350
rect 2586 7110 2646 7212
rect 3044 7110 3104 7216
rect 2580 7106 2652 7110
rect 2580 7054 2590 7106
rect 2642 7054 2652 7106
rect 2580 7050 2652 7054
rect 3038 7106 3110 7110
rect 3038 7054 3048 7106
rect 3100 7054 3110 7106
rect 3038 7050 3110 7054
rect -2218 6700 2426 6760
rect 3280 6630 3340 7342
rect 3504 7110 3564 7220
rect 3498 7106 3570 7110
rect 3498 7054 3508 7106
rect 3560 7054 3570 7106
rect 3498 7050 3570 7054
rect 3734 7108 3794 7344
rect 5316 7327 5428 7365
rect 3966 7108 4026 7224
rect 4192 7108 4252 7326
rect 5316 7293 5355 7327
rect 5389 7293 5428 7327
rect 5316 7255 5428 7293
rect 5316 7221 5355 7255
rect 5389 7221 5428 7255
rect 5316 7183 5428 7221
rect 5316 7149 5355 7183
rect 5389 7149 5428 7183
rect 5316 7111 5428 7149
rect 5316 7108 5355 7111
rect 3734 7077 5355 7108
rect 5389 7077 5428 7111
rect 3734 7048 5428 7077
rect -5028 6607 -4916 6618
rect -5028 6573 -4989 6607
rect -4955 6573 -4916 6607
rect -5028 6535 -4916 6573
rect -5028 6501 -4989 6535
rect -4955 6501 -4916 6535
rect -5028 6463 -4916 6501
rect -5028 6429 -4989 6463
rect -4955 6429 -4916 6463
rect -5028 6391 -4916 6429
rect -5028 6357 -4989 6391
rect -4955 6357 -4916 6391
rect -5028 6319 -4916 6357
rect -5028 6285 -4989 6319
rect -4955 6285 -4916 6319
rect -5028 6247 -4916 6285
rect -5028 6213 -4989 6247
rect -4955 6213 -4916 6247
rect -5028 6175 -4916 6213
rect -5028 6141 -4989 6175
rect -4955 6141 -4916 6175
rect -4608 6146 -4548 6618
rect -4380 6254 -4320 6618
rect -3136 6570 3340 6630
rect 4192 6614 4252 7048
rect 5316 7039 5428 7048
rect 5316 7005 5355 7039
rect 5389 7005 5428 7039
rect 5316 6967 5428 7005
rect 5316 6933 5355 6967
rect 5389 6933 5428 6967
rect 5316 6895 5428 6933
rect 5316 6861 5355 6895
rect 5389 6861 5428 6895
rect 5316 6823 5428 6861
rect 5316 6789 5355 6823
rect 5389 6789 5428 6823
rect 5316 6751 5428 6789
rect 5316 6717 5355 6751
rect 5389 6717 5428 6751
rect 5316 6679 5428 6717
rect 5316 6645 5355 6679
rect 5389 6645 5428 6679
rect 5316 6614 5428 6645
rect 4192 6607 5428 6614
rect 4192 6573 5355 6607
rect 5389 6573 5428 6607
rect 4192 6554 5428 6573
rect -4156 6520 -4084 6524
rect -4156 6468 -4146 6520
rect -4094 6468 -4084 6520
rect -4156 6464 -4084 6468
rect -5028 6103 -4916 6141
rect -4150 6126 -4090 6464
rect -3918 6362 -654 6422
rect -3918 6250 -3858 6362
rect -3456 6266 -3396 6362
rect -3002 6260 -2942 6362
rect -2540 6260 -2480 6362
rect -2086 6260 -2026 6362
rect -1636 6266 -1576 6362
rect -1170 6272 -1110 6362
rect -714 6266 -654 6362
rect -258 6344 910 6404
rect -258 6254 -198 6344
rect -28 6178 32 6344
rect 392 6172 452 6344
rect 624 6254 684 6344
rect 850 6150 910 6344
rect 1076 6362 4340 6422
rect 1076 6250 1136 6362
rect 1538 6266 1598 6362
rect 1992 6260 2052 6362
rect 2454 6260 2514 6362
rect 2908 6260 2968 6362
rect 3358 6266 3418 6362
rect 3824 6272 3884 6362
rect 4280 6266 4340 6362
rect 4742 6256 4802 6554
rect 4968 6140 5028 6554
rect 5316 6535 5428 6554
rect 5316 6501 5355 6535
rect 5389 6501 5428 6535
rect 5316 6463 5428 6501
rect 5316 6429 5355 6463
rect 5389 6429 5428 6463
rect 5316 6391 5428 6429
rect 5316 6357 5355 6391
rect 5389 6357 5428 6391
rect 5316 6319 5428 6357
rect 5316 6285 5355 6319
rect 5389 6285 5428 6319
rect 5316 6247 5428 6285
rect 5316 6213 5355 6247
rect 5389 6213 5428 6247
rect 5316 6175 5428 6213
rect 5316 6141 5355 6175
rect 5389 6141 5428 6175
rect -5028 6069 -4989 6103
rect -4955 6069 -4916 6103
rect -5028 6031 -4916 6069
rect -5028 5997 -4989 6031
rect -4955 5997 -4916 6031
rect -5028 5959 -4916 5997
rect -5028 5925 -4989 5959
rect -4955 5925 -4916 5959
rect -5028 5887 -4916 5925
rect -5028 5853 -4989 5887
rect -4955 5853 -4916 5887
rect -5028 5815 -4916 5853
rect -5028 5781 -4989 5815
rect -4955 5781 -4916 5815
rect -5028 5743 -4916 5781
rect -5028 5709 -4989 5743
rect -4955 5709 -4916 5743
rect -5028 5671 -4916 5709
rect -5028 5637 -4989 5671
rect -4955 5637 -4916 5671
rect -5028 5599 -4916 5637
rect -5028 5565 -4989 5599
rect -4955 5565 -4916 5599
rect -5028 5527 -4916 5565
rect -5028 5493 -4989 5527
rect -4955 5493 -4916 5527
rect -5028 5455 -4916 5493
rect -5028 5421 -4989 5455
rect -4955 5421 -4916 5455
rect -5028 5383 -4916 5421
rect -5028 5349 -4989 5383
rect -4955 5349 -4916 5383
rect -5028 5311 -4916 5349
rect -5028 5277 -4989 5311
rect -4955 5277 -4916 5311
rect -5028 5239 -4916 5277
rect -5028 5205 -4989 5239
rect -4955 5205 -4916 5239
rect -5028 5167 -4916 5205
rect -5028 5133 -4989 5167
rect -4955 5133 -4916 5167
rect -5028 5095 -4916 5133
rect -5028 5061 -4989 5095
rect -4955 5061 -4916 5095
rect 5316 6103 5428 6141
rect 5316 6069 5355 6103
rect 5389 6069 5428 6103
rect 5316 6031 5428 6069
rect 5316 5997 5355 6031
rect 5389 5997 5428 6031
rect 5316 5959 5428 5997
rect 5316 5925 5355 5959
rect 5389 5925 5428 5959
rect 5316 5887 5428 5925
rect 5316 5853 5355 5887
rect 5389 5853 5428 5887
rect 5316 5815 5428 5853
rect 5316 5781 5355 5815
rect 5389 5781 5428 5815
rect 5316 5743 5428 5781
rect 5316 5709 5355 5743
rect 5389 5709 5428 5743
rect 5316 5671 5428 5709
rect 5316 5637 5355 5671
rect 5389 5637 5428 5671
rect 5316 5599 5428 5637
rect 5316 5565 5355 5599
rect 5389 5565 5428 5599
rect 5316 5527 5428 5565
rect 5316 5493 5355 5527
rect 5389 5493 5428 5527
rect 5316 5455 5428 5493
rect 5316 5421 5355 5455
rect 5389 5421 5428 5455
rect 5316 5383 5428 5421
rect 5316 5349 5355 5383
rect 5389 5349 5428 5383
rect 5316 5311 5428 5349
rect 5316 5277 5355 5311
rect 5389 5277 5428 5311
rect 5316 5239 5428 5277
rect 5316 5205 5355 5239
rect 5389 5205 5428 5239
rect 5316 5167 5428 5205
rect 5316 5133 5355 5167
rect 5389 5133 5428 5167
rect 5316 5095 5428 5133
rect -5028 5023 -4916 5061
rect -5028 4989 -4989 5023
rect -4955 4989 -4916 5023
rect -5028 4951 -4916 4989
rect -5028 4917 -4989 4951
rect -4955 4917 -4916 4951
rect -5028 4879 -4916 4917
rect -5028 4845 -4989 4879
rect -4955 4845 -4916 4879
rect -5028 4807 -4916 4845
rect -5028 4773 -4989 4807
rect -4955 4773 -4916 4807
rect -5028 4584 -4916 4773
rect -4608 4584 -4548 5038
rect -4380 4584 -4320 4958
rect -3926 4850 -3866 4962
rect -3464 4850 -3404 4946
rect -3010 4850 -2950 4952
rect -2548 4850 -2488 4952
rect -2094 4850 -2034 4952
rect -1644 4850 -1584 4946
rect -1178 4850 -1118 4940
rect -722 4850 -662 4946
rect -3926 4846 -662 4850
rect -3926 4842 -3006 4846
rect -3926 4790 -3922 4842
rect -3870 4790 -3460 4842
rect -3408 4794 -3006 4842
rect -2954 4794 -2544 4846
rect -2492 4840 -1640 4846
rect -2492 4794 -2090 4840
rect -3408 4790 -2090 4794
rect -3926 4780 -3866 4790
rect -3464 4780 -3404 4790
rect -3010 4784 -2950 4790
rect -2548 4784 -2488 4790
rect -2094 4788 -2090 4790
rect -2038 4794 -1640 4840
rect -1588 4794 -1174 4846
rect -1122 4842 -662 4846
rect -1122 4794 -718 4842
rect -2038 4790 -718 4794
rect -666 4790 -662 4842
rect -2038 4788 -2034 4790
rect -2094 4778 -2034 4788
rect -1644 4784 -1584 4790
rect -1178 4784 -1118 4790
rect -722 4780 -662 4790
rect -488 4724 -428 5084
rect 5316 5061 5355 5095
rect 5389 5061 5428 5095
rect -494 4720 -422 4724
rect -494 4668 -484 4720
rect -432 4668 -422 4720
rect -494 4664 -422 4668
rect -258 4584 -198 4960
rect -30 4584 30 5052
rect 390 4584 450 5052
rect 618 4584 678 4956
rect 848 4584 908 5058
rect 1076 4850 1136 4962
rect 1538 4850 1598 4946
rect 1992 4850 2052 4952
rect 2454 4850 2514 4952
rect 2908 4850 2968 4952
rect 3358 4850 3418 4946
rect 3824 4850 3884 4940
rect 4280 4850 4340 4946
rect 1076 4842 1542 4850
rect 1076 4790 1080 4842
rect 1132 4798 1542 4842
rect 1594 4844 3362 4850
rect 1594 4798 1996 4844
rect 1132 4792 1996 4798
rect 2048 4792 2458 4844
rect 2510 4792 2912 4844
rect 2964 4798 3362 4844
rect 3414 4844 4340 4850
rect 3414 4798 3828 4844
rect 2964 4792 3828 4798
rect 3880 4792 4284 4844
rect 4336 4792 4340 4844
rect 1132 4790 4340 4792
rect 1076 4780 1136 4790
rect 1538 4788 1598 4790
rect 1992 4782 2052 4790
rect 2454 4782 2514 4790
rect 2908 4782 2968 4790
rect 3358 4788 3418 4790
rect 3824 4782 3884 4790
rect 4280 4782 4340 4790
rect 4512 4714 4572 5024
rect 4512 4662 4516 4714
rect 4568 4662 4572 4714
rect 4512 4652 4572 4662
rect 4742 4584 4802 4956
rect 4970 4584 5030 5050
rect 5316 5023 5428 5061
rect 5316 4989 5355 5023
rect 5389 4989 5428 5023
rect 5316 4951 5428 4989
rect 5316 4917 5355 4951
rect 5389 4917 5428 4951
rect 5316 4879 5428 4917
rect 5316 4845 5355 4879
rect 5389 4845 5428 4879
rect 5316 4807 5428 4845
rect 5316 4773 5355 4807
rect 5389 4773 5428 4807
rect 5316 4584 5428 4773
rect -5028 4545 5428 4584
rect -5028 4511 -4893 4545
rect -4859 4511 -4821 4545
rect -4787 4511 -4749 4545
rect -4715 4511 -4677 4545
rect -4643 4511 -4605 4545
rect -4571 4511 -4533 4545
rect -4499 4511 -4461 4545
rect -4427 4511 -4389 4545
rect -4355 4511 -4317 4545
rect -4283 4511 -4245 4545
rect -4211 4511 -4173 4545
rect -4139 4511 -4101 4545
rect -4067 4511 -4029 4545
rect -3995 4511 -3957 4545
rect -3923 4511 -3885 4545
rect -3851 4511 -3813 4545
rect -3779 4511 -3741 4545
rect -3707 4511 -3669 4545
rect -3635 4511 -3597 4545
rect -3563 4511 -3525 4545
rect -3491 4511 -3453 4545
rect -3419 4511 -3381 4545
rect -3347 4511 -3309 4545
rect -3275 4511 -3237 4545
rect -3203 4511 -3165 4545
rect -3131 4511 -3093 4545
rect -3059 4511 -3021 4545
rect -2987 4511 -2949 4545
rect -2915 4511 -2877 4545
rect -2843 4511 -2805 4545
rect -2771 4511 -2733 4545
rect -2699 4511 -2661 4545
rect -2627 4511 -2589 4545
rect -2555 4511 -2517 4545
rect -2483 4511 -2445 4545
rect -2411 4511 -2373 4545
rect -2339 4511 -2301 4545
rect -2267 4511 -2229 4545
rect -2195 4511 -2157 4545
rect -2123 4511 -2085 4545
rect -2051 4511 -2013 4545
rect -1979 4511 -1941 4545
rect -1907 4511 -1869 4545
rect -1835 4511 -1797 4545
rect -1763 4511 -1725 4545
rect -1691 4511 -1653 4545
rect -1619 4511 -1581 4545
rect -1547 4511 -1509 4545
rect -1475 4511 -1437 4545
rect -1403 4511 -1365 4545
rect -1331 4511 -1293 4545
rect -1259 4511 -1221 4545
rect -1187 4511 -1149 4545
rect -1115 4511 -1077 4545
rect -1043 4511 -1005 4545
rect -971 4511 -933 4545
rect -899 4511 -861 4545
rect -827 4511 -789 4545
rect -755 4511 -717 4545
rect -683 4511 -645 4545
rect -611 4511 -573 4545
rect -539 4511 -501 4545
rect -467 4511 -429 4545
rect -395 4511 -357 4545
rect -323 4511 -285 4545
rect -251 4511 -213 4545
rect -179 4511 -141 4545
rect -107 4511 -69 4545
rect -35 4511 3 4545
rect 37 4511 75 4545
rect 109 4511 147 4545
rect 181 4511 219 4545
rect 253 4511 291 4545
rect 325 4511 363 4545
rect 397 4511 435 4545
rect 469 4511 507 4545
rect 541 4511 579 4545
rect 613 4511 651 4545
rect 685 4511 723 4545
rect 757 4511 795 4545
rect 829 4511 867 4545
rect 901 4511 939 4545
rect 973 4511 1011 4545
rect 1045 4511 1083 4545
rect 1117 4511 1155 4545
rect 1189 4511 1227 4545
rect 1261 4511 1299 4545
rect 1333 4511 1371 4545
rect 1405 4511 1443 4545
rect 1477 4511 1515 4545
rect 1549 4511 1587 4545
rect 1621 4511 1659 4545
rect 1693 4511 1731 4545
rect 1765 4511 1803 4545
rect 1837 4511 1875 4545
rect 1909 4511 1947 4545
rect 1981 4511 2019 4545
rect 2053 4511 2091 4545
rect 2125 4511 2163 4545
rect 2197 4511 2235 4545
rect 2269 4511 2307 4545
rect 2341 4511 2379 4545
rect 2413 4511 2451 4545
rect 2485 4511 2523 4545
rect 2557 4511 2595 4545
rect 2629 4511 2667 4545
rect 2701 4511 2739 4545
rect 2773 4511 2811 4545
rect 2845 4511 2883 4545
rect 2917 4511 2955 4545
rect 2989 4511 3027 4545
rect 3061 4511 3099 4545
rect 3133 4511 3171 4545
rect 3205 4511 3243 4545
rect 3277 4511 3315 4545
rect 3349 4511 3387 4545
rect 3421 4511 3459 4545
rect 3493 4511 3531 4545
rect 3565 4511 3603 4545
rect 3637 4511 3675 4545
rect 3709 4511 3747 4545
rect 3781 4511 3819 4545
rect 3853 4511 3891 4545
rect 3925 4511 3963 4545
rect 3997 4511 4035 4545
rect 4069 4511 4107 4545
rect 4141 4511 4179 4545
rect 4213 4511 4251 4545
rect 4285 4511 4323 4545
rect 4357 4511 4395 4545
rect 4429 4511 4467 4545
rect 4501 4511 4539 4545
rect 4573 4511 4611 4545
rect 4645 4511 4683 4545
rect 4717 4511 4755 4545
rect 4789 4511 4827 4545
rect 4861 4511 4899 4545
rect 4933 4511 4971 4545
rect 5005 4511 5043 4545
rect 5077 4511 5115 4545
rect 5149 4511 5187 4545
rect 5221 4511 5259 4545
rect 5293 4511 5428 4545
rect -5028 4472 5428 4511
rect -5028 4209 5428 4248
rect -5028 4175 -4893 4209
rect -4859 4175 -4821 4209
rect -4787 4175 -4749 4209
rect -4715 4175 -4677 4209
rect -4643 4175 -4605 4209
rect -4571 4175 -4533 4209
rect -4499 4175 -4461 4209
rect -4427 4175 -4389 4209
rect -4355 4175 -4317 4209
rect -4283 4175 -4245 4209
rect -4211 4175 -4173 4209
rect -4139 4175 -4101 4209
rect -4067 4175 -4029 4209
rect -3995 4175 -3957 4209
rect -3923 4175 -3885 4209
rect -3851 4175 -3813 4209
rect -3779 4175 -3741 4209
rect -3707 4175 -3669 4209
rect -3635 4175 -3597 4209
rect -3563 4175 -3525 4209
rect -3491 4175 -3453 4209
rect -3419 4175 -3381 4209
rect -3347 4175 -3309 4209
rect -3275 4175 -3237 4209
rect -3203 4175 -3165 4209
rect -3131 4175 -3093 4209
rect -3059 4175 -3021 4209
rect -2987 4175 -2949 4209
rect -2915 4175 -2877 4209
rect -2843 4175 -2805 4209
rect -2771 4175 -2733 4209
rect -2699 4175 -2661 4209
rect -2627 4175 -2589 4209
rect -2555 4175 -2517 4209
rect -2483 4175 -2445 4209
rect -2411 4175 -2373 4209
rect -2339 4175 -2301 4209
rect -2267 4175 -2229 4209
rect -2195 4175 -2157 4209
rect -2123 4175 -2085 4209
rect -2051 4175 -2013 4209
rect -1979 4175 -1941 4209
rect -1907 4175 -1869 4209
rect -1835 4175 -1797 4209
rect -1763 4175 -1725 4209
rect -1691 4175 -1653 4209
rect -1619 4175 -1581 4209
rect -1547 4175 -1509 4209
rect -1475 4175 -1437 4209
rect -1403 4175 -1365 4209
rect -1331 4175 -1293 4209
rect -1259 4175 -1221 4209
rect -1187 4175 -1149 4209
rect -1115 4175 -1077 4209
rect -1043 4175 -1005 4209
rect -971 4175 -933 4209
rect -899 4175 -861 4209
rect -827 4175 -789 4209
rect -755 4175 -717 4209
rect -683 4175 -645 4209
rect -611 4175 -573 4209
rect -539 4175 -501 4209
rect -467 4175 -429 4209
rect -395 4175 -357 4209
rect -323 4175 -285 4209
rect -251 4175 -213 4209
rect -179 4175 -141 4209
rect -107 4175 -69 4209
rect -35 4175 3 4209
rect 37 4175 75 4209
rect 109 4175 147 4209
rect 181 4175 219 4209
rect 253 4175 291 4209
rect 325 4175 363 4209
rect 397 4175 435 4209
rect 469 4175 507 4209
rect 541 4175 579 4209
rect 613 4175 651 4209
rect 685 4175 723 4209
rect 757 4175 795 4209
rect 829 4175 867 4209
rect 901 4175 939 4209
rect 973 4175 1011 4209
rect 1045 4175 1083 4209
rect 1117 4175 1155 4209
rect 1189 4175 1227 4209
rect 1261 4175 1299 4209
rect 1333 4175 1371 4209
rect 1405 4175 1443 4209
rect 1477 4175 1515 4209
rect 1549 4175 1587 4209
rect 1621 4175 1659 4209
rect 1693 4175 1731 4209
rect 1765 4175 1803 4209
rect 1837 4175 1875 4209
rect 1909 4175 1947 4209
rect 1981 4175 2019 4209
rect 2053 4175 2091 4209
rect 2125 4175 2163 4209
rect 2197 4175 2235 4209
rect 2269 4175 2307 4209
rect 2341 4175 2379 4209
rect 2413 4175 2451 4209
rect 2485 4175 2523 4209
rect 2557 4175 2595 4209
rect 2629 4175 2667 4209
rect 2701 4175 2739 4209
rect 2773 4175 2811 4209
rect 2845 4175 2883 4209
rect 2917 4175 2955 4209
rect 2989 4175 3027 4209
rect 3061 4175 3099 4209
rect 3133 4175 3171 4209
rect 3205 4175 3243 4209
rect 3277 4175 3315 4209
rect 3349 4175 3387 4209
rect 3421 4175 3459 4209
rect 3493 4175 3531 4209
rect 3565 4175 3603 4209
rect 3637 4175 3675 4209
rect 3709 4175 3747 4209
rect 3781 4175 3819 4209
rect 3853 4175 3891 4209
rect 3925 4175 3963 4209
rect 3997 4175 4035 4209
rect 4069 4175 4107 4209
rect 4141 4175 4179 4209
rect 4213 4175 4251 4209
rect 4285 4175 4323 4209
rect 4357 4175 4395 4209
rect 4429 4175 4467 4209
rect 4501 4175 4539 4209
rect 4573 4175 4611 4209
rect 4645 4175 4683 4209
rect 4717 4175 4755 4209
rect 4789 4175 4827 4209
rect 4861 4175 4899 4209
rect 4933 4175 4971 4209
rect 5005 4175 5043 4209
rect 5077 4175 5115 4209
rect 5149 4175 5187 4209
rect 5221 4175 5259 4209
rect 5293 4175 5428 4209
rect -5028 4136 5428 4175
rect -5028 3999 -4916 4136
rect -5028 3965 -4989 3999
rect -4955 3965 -4916 3999
rect -5028 3927 -4916 3965
rect -5028 3893 -4989 3927
rect -4955 3893 -4916 3927
rect -5028 3855 -4916 3893
rect -5028 3821 -4989 3855
rect -4955 3821 -4916 3855
rect -5028 3783 -4916 3821
rect -5028 3749 -4989 3783
rect -4955 3749 -4916 3783
rect -5028 3711 -4916 3749
rect -5028 3677 -4989 3711
rect -4955 3677 -4916 3711
rect -5028 3639 -4916 3677
rect -4608 3660 -4548 4136
rect -4378 3748 -4318 4136
rect -488 4040 -428 4050
rect -488 3988 -484 4040
rect -432 3988 -428 4040
rect -3920 3912 -656 3916
rect -3920 3910 -3460 3912
rect -3932 3906 -3460 3910
rect -3932 3854 -3922 3906
rect -3870 3860 -3460 3906
rect -3408 3906 -2544 3912
rect -3408 3860 -3006 3906
rect -3870 3856 -3006 3860
rect -3870 3854 -3860 3856
rect -3932 3850 -3860 3854
rect -3926 3754 -3860 3850
rect -3920 3750 -3860 3754
rect -3464 3760 -3398 3856
rect -3016 3854 -3006 3856
rect -2954 3860 -2544 3906
rect -2492 3860 -2090 3912
rect -2038 3860 -1640 3912
rect -1588 3906 -718 3912
rect -1588 3860 -1174 3906
rect -2954 3856 -1174 3860
rect -2954 3854 -2944 3856
rect -3016 3850 -2944 3854
rect -3464 3752 -3404 3760
rect -3010 3758 -2944 3850
rect -3004 3754 -2944 3758
rect -2548 3754 -2482 3856
rect -2094 3758 -2028 3856
rect -2088 3754 -2028 3758
rect -1644 3760 -1578 3856
rect -1184 3854 -1174 3856
rect -1122 3860 -718 3906
rect -666 3860 -656 3912
rect -1122 3856 -656 3860
rect -1122 3854 -1112 3856
rect -1184 3850 -1112 3854
rect -1178 3766 -1112 3850
rect -1644 3748 -1584 3760
rect -1178 3748 -1118 3766
rect -722 3760 -656 3856
rect -722 3758 -662 3760
rect -488 3670 -428 3988
rect -260 3752 -200 4136
rect -28 3672 32 4136
rect 392 3664 452 4136
rect 626 3752 686 4136
rect -5028 3605 -4989 3639
rect -4955 3605 -4916 3639
rect 848 3636 908 4136
rect 4506 4052 4578 4056
rect 4506 4000 4516 4052
rect 4568 4000 4578 4052
rect 4506 3996 4578 4000
rect 3352 3916 3424 3920
rect 1070 3912 3362 3916
rect 1070 3860 1080 3912
rect 1132 3910 3362 3912
rect 1132 3860 1542 3910
rect 1070 3858 1542 3860
rect 1594 3858 1996 3910
rect 2048 3858 2458 3910
rect 2510 3858 2912 3910
rect 2964 3864 3362 3910
rect 3414 3912 4346 3916
rect 3414 3864 3828 3912
rect 2964 3860 3828 3864
rect 3880 3860 4284 3912
rect 4336 3860 4346 3912
rect 2964 3858 4346 3860
rect 1070 3856 4346 3858
rect 1076 3750 1140 3856
rect 1532 3854 1604 3856
rect 1986 3854 2058 3856
rect 2448 3854 2520 3856
rect 2902 3854 2974 3856
rect 1538 3760 1602 3854
rect 1538 3752 1598 3760
rect 1992 3754 2056 3854
rect 2454 3754 2518 3854
rect 2908 3754 2972 3854
rect 3358 3760 3422 3856
rect 3824 3766 3888 3856
rect 1076 3746 1136 3750
rect 1992 3746 2052 3754
rect 2454 3748 2514 3754
rect 2908 3748 2968 3754
rect 3358 3752 3418 3760
rect 3824 3752 3884 3766
rect 4280 3760 4344 3856
rect 4280 3748 4340 3760
rect 4512 3658 4572 3996
rect 4752 3754 4812 4136
rect 4970 3660 5030 4136
rect 5316 3999 5428 4136
rect 5316 3965 5355 3999
rect 5389 3965 5428 3999
rect 5316 3927 5428 3965
rect 5316 3893 5355 3927
rect 5389 3893 5428 3927
rect 5316 3855 5428 3893
rect 5316 3821 5355 3855
rect 5389 3821 5428 3855
rect 5316 3783 5428 3821
rect 5316 3749 5355 3783
rect 5389 3749 5428 3783
rect 5316 3711 5428 3749
rect 5316 3677 5355 3711
rect 5389 3677 5428 3711
rect 5316 3639 5428 3677
rect -5028 3567 -4916 3605
rect 5316 3605 5355 3639
rect 5389 3605 5428 3639
rect -5028 3533 -4989 3567
rect -4955 3533 -4916 3567
rect -5028 3495 -4916 3533
rect -5028 3461 -4989 3495
rect -4955 3461 -4916 3495
rect -5028 3423 -4916 3461
rect -5028 3389 -4989 3423
rect -4955 3389 -4916 3423
rect -5028 3351 -4916 3389
rect -5028 3317 -4989 3351
rect -4955 3317 -4916 3351
rect -5028 3279 -4916 3317
rect -5028 3245 -4989 3279
rect -4955 3245 -4916 3279
rect -5028 3207 -4916 3245
rect -5028 3173 -4989 3207
rect -4955 3173 -4916 3207
rect -5028 3135 -4916 3173
rect -5028 3101 -4989 3135
rect -4955 3101 -4916 3135
rect -5028 3063 -4916 3101
rect -5028 3029 -4989 3063
rect -4955 3029 -4916 3063
rect -5028 2991 -4916 3029
rect -4608 3308 -4548 3564
rect -4380 3308 -4320 3472
rect -4608 3248 -4320 3308
rect -4608 3012 -4548 3248
rect -4380 3082 -4320 3248
rect -4152 3004 -4092 3566
rect -3926 3368 -3866 3474
rect -3464 3368 -3404 3464
rect -3010 3368 -2950 3470
rect -2548 3368 -2488 3470
rect -2094 3368 -2034 3470
rect -1644 3368 -1584 3464
rect -1178 3368 -1118 3458
rect -722 3368 -662 3464
rect -3926 3308 -662 3368
rect -3920 3188 -656 3248
rect -3920 3082 -3860 3188
rect -3458 3092 -3398 3188
rect -3004 3086 -2944 3188
rect -2542 3086 -2482 3188
rect -2088 3086 -2028 3188
rect -1638 3092 -1578 3188
rect -1172 3098 -1112 3188
rect -716 3092 -656 3188
rect -260 3084 -200 3476
rect -5028 2957 -4989 2991
rect -4955 2957 -4916 2991
rect -5028 2919 -4916 2957
rect -5028 2885 -4989 2919
rect -4955 2885 -4916 2919
rect -5028 2847 -4916 2885
rect -5028 2813 -4989 2847
rect -4955 2813 -4916 2847
rect -5028 2775 -4916 2813
rect -5028 2741 -4989 2775
rect -4955 2741 -4916 2775
rect -5028 2703 -4916 2741
rect -5028 2669 -4989 2703
rect -4955 2669 -4916 2703
rect -5028 2631 -4916 2669
rect -5028 2597 -4989 2631
rect -4955 2597 -4916 2631
rect -5028 2559 -4916 2597
rect -5028 2525 -4989 2559
rect -4955 2525 -4916 2559
rect -5028 2487 -4916 2525
rect -5028 2453 -4989 2487
rect -4955 2453 -4916 2487
rect -4616 2476 -4556 2886
rect -4376 2476 -4316 2806
rect -3926 2700 -3866 2806
rect -3464 2700 -3404 2796
rect -3010 2700 -2950 2802
rect -2548 2700 -2488 2802
rect -2094 2700 -2034 2802
rect -1644 2700 -1584 2796
rect -1178 2700 -1118 2790
rect -722 2700 -662 2796
rect -3926 2640 -662 2700
rect -488 2476 -428 2884
rect -262 2476 -202 2808
rect -28 2476 32 3580
rect 388 3370 448 3560
rect 616 3370 676 3478
rect 848 3370 908 3568
rect 388 3310 908 3370
rect 388 2476 448 3310
rect 616 2476 676 3310
rect 848 2476 908 3310
rect 1074 3368 1134 3474
rect 1536 3368 1596 3464
rect 1990 3368 2050 3470
rect 2452 3368 2512 3470
rect 2906 3368 2966 3470
rect 3356 3368 3416 3464
rect 3822 3368 3882 3458
rect 4278 3368 4338 3464
rect 1074 3308 4338 3368
rect 4742 2476 4802 3474
rect 4968 2476 5028 3570
rect 5316 3567 5428 3605
rect 5316 3533 5355 3567
rect 5389 3533 5428 3567
rect 5316 3495 5428 3533
rect 5316 3461 5355 3495
rect 5389 3461 5428 3495
rect 5316 3423 5428 3461
rect 5316 3389 5355 3423
rect 5389 3389 5428 3423
rect 5316 3351 5428 3389
rect 5316 3317 5355 3351
rect 5389 3317 5428 3351
rect 5316 3279 5428 3317
rect 5316 3245 5355 3279
rect 5389 3245 5428 3279
rect 5316 3207 5428 3245
rect 5316 3173 5355 3207
rect 5389 3173 5428 3207
rect 5316 3135 5428 3173
rect 5316 3101 5355 3135
rect 5389 3101 5428 3135
rect 5316 3063 5428 3101
rect 5316 3029 5355 3063
rect 5389 3029 5428 3063
rect 5316 2991 5428 3029
rect 5316 2957 5355 2991
rect 5389 2957 5428 2991
rect 5316 2919 5428 2957
rect 5316 2885 5355 2919
rect 5389 2885 5428 2919
rect 5316 2847 5428 2885
rect 5316 2813 5355 2847
rect 5389 2813 5428 2847
rect 5316 2775 5428 2813
rect 5316 2741 5355 2775
rect 5389 2741 5428 2775
rect 5316 2703 5428 2741
rect 5316 2669 5355 2703
rect 5389 2669 5428 2703
rect 5316 2631 5428 2669
rect 5316 2597 5355 2631
rect 5389 2597 5428 2631
rect 5316 2559 5428 2597
rect 5316 2525 5355 2559
rect 5389 2525 5428 2559
rect 5316 2487 5428 2525
rect -5028 2415 -4916 2453
rect -5028 2381 -4989 2415
rect -4955 2381 -4916 2415
rect -5028 2343 -4916 2381
rect -5028 2309 -4989 2343
rect -4955 2309 -4916 2343
rect -4680 2431 5090 2476
rect -4680 2379 -4608 2431
rect -4556 2379 -4028 2431
rect -3976 2379 -3428 2431
rect -3376 2379 -2828 2431
rect -2776 2379 -2228 2431
rect -2176 2379 -1628 2431
rect -1576 2379 -1028 2431
rect -976 2379 -428 2431
rect -376 2379 172 2431
rect 224 2379 772 2431
rect 824 2379 1372 2431
rect 1424 2379 1972 2431
rect 2024 2379 2572 2431
rect 2624 2379 3172 2431
rect 3224 2379 3772 2431
rect 3824 2379 4372 2431
rect 4424 2379 4972 2431
rect 5024 2379 5090 2431
rect -4680 2332 5090 2379
rect 5316 2453 5355 2487
rect 5389 2453 5428 2487
rect 5316 2415 5428 2453
rect 5316 2381 5355 2415
rect 5389 2381 5428 2415
rect 5316 2343 5428 2381
rect -5028 2271 -4916 2309
rect -5028 2237 -4989 2271
rect -4955 2237 -4916 2271
rect -5028 2199 -4916 2237
rect -5028 2165 -4989 2199
rect -4955 2184 -4916 2199
rect 5316 2309 5355 2343
rect 5389 2309 5428 2343
rect 5316 2271 5428 2309
rect 5316 2237 5355 2271
rect 5389 2237 5428 2271
rect 5316 2199 5428 2237
rect 5316 2184 5355 2199
rect -4955 2165 -4306 2184
rect -5028 2156 -4306 2165
rect -5028 2127 -4898 2156
rect -5028 2093 -4989 2127
rect -4955 2093 -4898 2127
rect -5028 2055 -4898 2093
rect -5028 2021 -4989 2055
rect -4955 2021 -4898 2055
rect -5028 1912 -4898 2021
rect -4334 1912 -4306 2156
rect -5028 1884 -4306 1912
rect 4706 2165 5355 2184
rect 5389 2165 5428 2199
rect 4706 2156 5428 2165
rect 4706 1912 4734 2156
rect 5298 2127 5428 2156
rect 5298 2093 5355 2127
rect 5389 2093 5428 2127
rect 5298 2055 5428 2093
rect 5298 2021 5355 2055
rect 5389 2021 5428 2055
rect 5298 1912 5428 2021
rect 4706 1884 5428 1912
rect -5028 1845 5428 1884
rect -5028 1811 -4893 1845
rect -4859 1811 -4821 1845
rect -4787 1811 -4749 1845
rect -4715 1811 -4677 1845
rect -4643 1811 -4605 1845
rect -4571 1811 -4533 1845
rect -4499 1811 -4461 1845
rect -4427 1811 -4389 1845
rect -4355 1811 -4317 1845
rect -4283 1811 -4245 1845
rect -4211 1811 -4173 1845
rect -4139 1811 -4101 1845
rect -4067 1811 -4029 1845
rect -3995 1811 -3957 1845
rect -3923 1811 -3885 1845
rect -3851 1811 -3813 1845
rect -3779 1811 -3741 1845
rect -3707 1811 -3669 1845
rect -3635 1811 -3597 1845
rect -3563 1811 -3525 1845
rect -3491 1811 -3453 1845
rect -3419 1811 -3381 1845
rect -3347 1811 -3309 1845
rect -3275 1811 -3237 1845
rect -3203 1811 -3165 1845
rect -3131 1811 -3093 1845
rect -3059 1811 -3021 1845
rect -2987 1811 -2949 1845
rect -2915 1811 -2877 1845
rect -2843 1811 -2805 1845
rect -2771 1811 -2733 1845
rect -2699 1811 -2661 1845
rect -2627 1811 -2589 1845
rect -2555 1811 -2517 1845
rect -2483 1811 -2445 1845
rect -2411 1811 -2373 1845
rect -2339 1811 -2301 1845
rect -2267 1811 -2229 1845
rect -2195 1811 -2157 1845
rect -2123 1811 -2085 1845
rect -2051 1811 -2013 1845
rect -1979 1811 -1941 1845
rect -1907 1811 -1869 1845
rect -1835 1811 -1797 1845
rect -1763 1811 -1725 1845
rect -1691 1811 -1653 1845
rect -1619 1811 -1581 1845
rect -1547 1811 -1509 1845
rect -1475 1811 -1437 1845
rect -1403 1811 -1365 1845
rect -1331 1811 -1293 1845
rect -1259 1811 -1221 1845
rect -1187 1811 -1149 1845
rect -1115 1811 -1077 1845
rect -1043 1811 -1005 1845
rect -971 1811 -933 1845
rect -899 1811 -861 1845
rect -827 1811 -789 1845
rect -755 1811 -717 1845
rect -683 1811 -645 1845
rect -611 1811 -573 1845
rect -539 1811 -501 1845
rect -467 1811 -429 1845
rect -395 1811 -357 1845
rect -323 1811 -285 1845
rect -251 1811 -213 1845
rect -179 1811 -141 1845
rect -107 1811 -69 1845
rect -35 1811 3 1845
rect 37 1811 75 1845
rect 109 1811 147 1845
rect 181 1811 219 1845
rect 253 1811 291 1845
rect 325 1811 363 1845
rect 397 1811 435 1845
rect 469 1811 507 1845
rect 541 1811 579 1845
rect 613 1811 651 1845
rect 685 1811 723 1845
rect 757 1811 795 1845
rect 829 1811 867 1845
rect 901 1811 939 1845
rect 973 1811 1011 1845
rect 1045 1811 1083 1845
rect 1117 1811 1155 1845
rect 1189 1811 1227 1845
rect 1261 1811 1299 1845
rect 1333 1811 1371 1845
rect 1405 1811 1443 1845
rect 1477 1811 1515 1845
rect 1549 1811 1587 1845
rect 1621 1811 1659 1845
rect 1693 1811 1731 1845
rect 1765 1811 1803 1845
rect 1837 1811 1875 1845
rect 1909 1811 1947 1845
rect 1981 1811 2019 1845
rect 2053 1811 2091 1845
rect 2125 1811 2163 1845
rect 2197 1811 2235 1845
rect 2269 1811 2307 1845
rect 2341 1811 2379 1845
rect 2413 1811 2451 1845
rect 2485 1811 2523 1845
rect 2557 1811 2595 1845
rect 2629 1811 2667 1845
rect 2701 1811 2739 1845
rect 2773 1811 2811 1845
rect 2845 1811 2883 1845
rect 2917 1811 2955 1845
rect 2989 1811 3027 1845
rect 3061 1811 3099 1845
rect 3133 1811 3171 1845
rect 3205 1811 3243 1845
rect 3277 1811 3315 1845
rect 3349 1811 3387 1845
rect 3421 1811 3459 1845
rect 3493 1811 3531 1845
rect 3565 1811 3603 1845
rect 3637 1811 3675 1845
rect 3709 1811 3747 1845
rect 3781 1811 3819 1845
rect 3853 1811 3891 1845
rect 3925 1811 3963 1845
rect 3997 1811 4035 1845
rect 4069 1811 4107 1845
rect 4141 1811 4179 1845
rect 4213 1811 4251 1845
rect 4285 1811 4323 1845
rect 4357 1811 4395 1845
rect 4429 1811 4467 1845
rect 4501 1811 4539 1845
rect 4573 1811 4611 1845
rect 4645 1811 4683 1845
rect 4717 1811 4755 1845
rect 4789 1811 4827 1845
rect 4861 1811 4899 1845
rect 4933 1811 4971 1845
rect 5005 1811 5043 1845
rect 5077 1811 5115 1845
rect 5149 1811 5187 1845
rect 5221 1811 5259 1845
rect 5293 1811 5428 1845
rect -5028 1772 5428 1811
<< via1 >>
rect -4898 9944 -4334 10188
rect 4734 9944 5298 10188
rect -4042 9673 -3990 9725
rect -3442 9673 -3390 9725
rect -2842 9673 -2790 9725
rect -2242 9673 -2190 9725
rect -1642 9673 -1590 9725
rect -1042 9673 -990 9725
rect -442 9673 -390 9725
rect 158 9673 210 9725
rect 758 9673 810 9725
rect 1358 9673 1410 9725
rect 1958 9673 2010 9725
rect 2558 9673 2610 9725
rect 3158 9673 3210 9725
rect 3758 9673 3810 9725
rect 4178 9673 4230 9725
rect -3356 9028 -3304 9080
rect -2900 9028 -2848 9080
rect -2440 9028 -2388 9080
rect -1984 9028 -1932 9080
rect -1526 9028 -1474 9080
rect -1062 9028 -1010 9080
rect -612 9028 -560 9080
rect -156 9028 -104 9080
rect 312 9028 364 9080
rect 770 9028 822 9080
rect 1226 9028 1278 9080
rect 1682 9028 1734 9080
rect 2138 9028 2190 9080
rect 2594 9028 2646 9080
rect 3052 9028 3104 9080
rect 3512 9028 3564 9080
rect -3360 7054 -3308 7106
rect -2904 7054 -2852 7106
rect -2444 7054 -2392 7106
rect -1988 7054 -1936 7106
rect -1530 7054 -1478 7106
rect -1066 7054 -1014 7106
rect -612 7054 -560 7106
rect -154 7099 -102 7106
rect -154 7065 -145 7099
rect -145 7065 -111 7099
rect -111 7065 -102 7099
rect -154 7054 -102 7065
rect 80 7066 132 7118
rect 306 7099 358 7106
rect 306 7065 315 7099
rect 315 7065 349 7099
rect 349 7065 358 7099
rect 306 7054 358 7065
rect 762 7054 814 7106
rect 1222 7054 1274 7106
rect 1678 7054 1730 7106
rect 2134 7054 2186 7106
rect 2590 7054 2642 7106
rect 3048 7054 3100 7106
rect 3508 7054 3560 7106
rect -4146 6468 -4094 6520
rect -3922 4790 -3870 4842
rect -3460 4790 -3408 4842
rect -3006 4794 -2954 4846
rect -2544 4794 -2492 4846
rect -2090 4788 -2038 4840
rect -1640 4794 -1588 4846
rect -1174 4794 -1122 4846
rect -718 4790 -666 4842
rect -484 4668 -432 4720
rect 1080 4790 1132 4842
rect 1542 4798 1594 4850
rect 1996 4792 2048 4844
rect 2458 4792 2510 4844
rect 2912 4792 2964 4844
rect 3362 4798 3414 4850
rect 3828 4792 3880 4844
rect 4284 4792 4336 4844
rect 4516 4662 4568 4714
rect -484 3988 -432 4040
rect -3922 3854 -3870 3906
rect -3460 3860 -3408 3912
rect -3006 3854 -2954 3906
rect -2544 3860 -2492 3912
rect -2090 3860 -2038 3912
rect -1640 3860 -1588 3912
rect -1174 3854 -1122 3906
rect -718 3860 -666 3912
rect 4516 4000 4568 4052
rect 1080 3860 1132 3912
rect 1542 3858 1594 3910
rect 1996 3858 2048 3910
rect 2458 3858 2510 3910
rect 2912 3858 2964 3910
rect 3362 3864 3414 3916
rect 3828 3860 3880 3912
rect 4284 3860 4336 3912
rect -4608 2379 -4556 2431
rect -4028 2379 -3976 2431
rect -3428 2379 -3376 2431
rect -2828 2379 -2776 2431
rect -2228 2379 -2176 2431
rect -1628 2379 -1576 2431
rect -1028 2379 -976 2431
rect -428 2379 -376 2431
rect 172 2379 224 2431
rect 772 2379 824 2431
rect 1372 2379 1424 2431
rect 1972 2379 2024 2431
rect 2572 2379 2624 2431
rect 3172 2379 3224 2431
rect 3772 2379 3824 2431
rect 4372 2379 4424 2431
rect 4972 2379 5024 2431
rect -4898 1912 -4334 2156
rect 4734 1912 5298 2156
<< metal2 >>
rect -4916 10214 -4316 10226
rect -4916 10188 -4884 10214
rect -4348 10188 -4316 10214
rect -4916 9944 -4898 10188
rect -4334 9944 -4316 10188
rect -4916 9918 -4884 9944
rect -4348 9918 -4316 9944
rect -4916 9906 -4316 9918
rect 4716 10214 5316 10226
rect 4716 10188 4748 10214
rect 5284 10188 5316 10214
rect 4716 9944 4734 10188
rect 5298 9944 5316 10188
rect 4716 9918 4748 9944
rect 5284 9918 5316 9944
rect 4716 9906 5316 9918
rect -4078 9727 4278 9756
rect -4078 9671 -4044 9727
rect -3988 9671 -3444 9727
rect -3388 9671 -2844 9727
rect -2788 9671 -2244 9727
rect -2188 9671 -1644 9727
rect -1588 9671 -1044 9727
rect -988 9671 -444 9727
rect -388 9671 156 9727
rect 212 9671 756 9727
rect 812 9671 1356 9727
rect 1412 9671 1956 9727
rect 2012 9671 2556 9727
rect 2612 9671 3156 9727
rect 3212 9671 3756 9727
rect 3812 9671 4176 9727
rect 4232 9671 4278 9727
rect -4078 9646 4278 9671
rect -3360 9084 -3300 9090
rect -2904 9084 -2844 9090
rect -2444 9084 -2384 9090
rect -1988 9084 -1928 9090
rect -1530 9084 -1470 9090
rect -1066 9084 -1006 9090
rect -616 9084 -556 9090
rect -160 9084 -100 9090
rect 308 9084 368 9090
rect 766 9084 826 9090
rect 1222 9084 1282 9090
rect 1678 9084 1738 9090
rect 2134 9084 2194 9090
rect 2590 9084 2650 9090
rect 3048 9084 3108 9090
rect 3508 9084 3568 9090
rect -3360 9080 3568 9084
rect -3360 9028 -3356 9080
rect -3304 9028 -2900 9080
rect -2848 9028 -2440 9080
rect -2388 9028 -1984 9080
rect -1932 9028 -1526 9080
rect -1474 9028 -1062 9080
rect -1010 9028 -612 9080
rect -560 9028 -156 9080
rect -104 9028 312 9080
rect 364 9028 770 9080
rect 822 9028 1226 9080
rect 1278 9028 1682 9080
rect 1734 9028 2138 9080
rect 2190 9028 2594 9080
rect 2646 9028 3052 9080
rect 3104 9028 3512 9080
rect 3564 9028 3568 9080
rect -3360 9024 3568 9028
rect -3360 9018 -3300 9024
rect -2904 9018 -2844 9024
rect -2444 9018 -2384 9024
rect -1988 9018 -1928 9024
rect -1530 9018 -1470 9024
rect -1066 9018 -1006 9024
rect -616 9018 -556 9024
rect -160 9018 -100 9024
rect 308 9018 368 9024
rect 766 9018 826 9024
rect 1222 9018 1282 9024
rect 1678 9018 1738 9024
rect 2134 9018 2194 9024
rect 2590 9018 2650 9024
rect 3048 9018 3108 9024
rect 3508 9018 3568 9024
rect 70 7118 142 7122
rect -3364 7110 -3304 7116
rect -2908 7110 -2848 7116
rect -2448 7110 -2388 7116
rect -1992 7110 -1932 7116
rect -1534 7110 -1474 7116
rect -1070 7110 -1010 7116
rect -616 7110 -556 7116
rect -158 7110 -98 7116
rect -3364 7106 -98 7110
rect -3364 7054 -3360 7106
rect -3308 7054 -2904 7106
rect -2852 7054 -2444 7106
rect -2392 7054 -1988 7106
rect -1936 7054 -1530 7106
rect -1478 7054 -1066 7106
rect -1014 7054 -612 7106
rect -560 7054 -154 7106
rect -102 7054 -98 7106
rect 70 7066 80 7118
rect 132 7066 142 7118
rect 70 7062 142 7066
rect 302 7110 362 7116
rect 758 7110 818 7116
rect 1218 7110 1278 7116
rect 1674 7110 1734 7116
rect 2130 7110 2190 7116
rect 2586 7110 2646 7116
rect 3044 7110 3104 7116
rect 3504 7110 3564 7116
rect 302 7106 3564 7110
rect -3364 7050 -98 7054
rect -3364 7044 -3304 7050
rect -2908 7044 -2848 7050
rect -2448 7044 -2388 7050
rect -1992 7044 -1932 7050
rect -1534 7044 -1474 7050
rect -1070 7044 -1010 7050
rect -616 7044 -556 7050
rect -158 7044 -98 7050
rect -4150 6524 -4090 6530
rect 76 6524 136 7062
rect 302 7054 306 7106
rect 358 7054 762 7106
rect 814 7054 1222 7106
rect 1274 7054 1678 7106
rect 1730 7054 2134 7106
rect 2186 7054 2590 7106
rect 2642 7054 3048 7106
rect 3100 7054 3508 7106
rect 3560 7054 3564 7106
rect 302 7050 3564 7054
rect 302 7044 362 7050
rect 758 7044 818 7050
rect 1218 7044 1278 7050
rect 1674 7044 1734 7050
rect 2130 7044 2190 7050
rect 2586 7044 2646 7050
rect 3044 7044 3104 7050
rect 3504 7044 3564 7050
rect -4150 6520 136 6524
rect -4150 6468 -4146 6520
rect -4094 6468 136 6520
rect -4150 6464 136 6468
rect -4150 6458 -4090 6464
rect 1532 4850 1604 4854
rect -3016 4846 -2944 4850
rect -3932 4842 -3860 4846
rect -3932 4790 -3922 4842
rect -3870 4790 -3860 4842
rect -3932 4786 -3860 4790
rect -3470 4842 -3398 4846
rect -3470 4790 -3460 4842
rect -3408 4790 -3398 4842
rect -3016 4794 -3006 4846
rect -2954 4794 -2944 4846
rect -3016 4790 -2944 4794
rect -2554 4846 -2482 4850
rect -2554 4794 -2544 4846
rect -2492 4794 -2482 4846
rect -1650 4846 -1578 4850
rect -2554 4790 -2482 4794
rect -2100 4840 -2028 4844
rect -3470 4786 -3398 4790
rect -3926 4392 -3866 4786
rect -3464 4392 -3404 4786
rect -3010 4392 -2950 4790
rect -2548 4392 -2488 4790
rect -2100 4788 -2090 4840
rect -2038 4788 -2028 4840
rect -1650 4794 -1640 4846
rect -1588 4794 -1578 4846
rect -1650 4790 -1578 4794
rect -1184 4846 -1112 4850
rect -1184 4794 -1174 4846
rect -1122 4794 -1112 4846
rect -1184 4790 -1112 4794
rect -728 4842 -656 4846
rect -728 4790 -718 4842
rect -666 4790 -656 4842
rect -2100 4784 -2028 4788
rect -2094 4392 -2034 4784
rect -1644 4392 -1584 4790
rect -1178 4392 -1118 4790
rect -728 4786 -656 4790
rect 1070 4842 1142 4846
rect 1070 4790 1080 4842
rect 1132 4790 1142 4842
rect 1532 4798 1542 4850
rect 1594 4798 1604 4850
rect 3352 4850 3424 4854
rect 1532 4794 1604 4798
rect 1986 4844 2058 4848
rect 1070 4786 1142 4790
rect -722 4392 -662 4786
rect -3928 4332 -662 4392
rect -3926 3906 -3866 4332
rect -3926 3854 -3922 3906
rect -3870 3854 -3866 3906
rect -3926 3844 -3866 3854
rect -3464 3912 -3404 4332
rect -3464 3860 -3460 3912
rect -3408 3860 -3404 3912
rect -3464 3850 -3404 3860
rect -3010 3906 -2950 4332
rect -3010 3854 -3006 3906
rect -2954 3854 -2950 3906
rect -3010 3844 -2950 3854
rect -2548 3912 -2488 4332
rect -2548 3860 -2544 3912
rect -2492 3860 -2488 3912
rect -2548 3850 -2488 3860
rect -2094 3912 -2034 4332
rect -2094 3860 -2090 3912
rect -2038 3860 -2034 3912
rect -2094 3850 -2034 3860
rect -1644 3912 -1584 4332
rect -1644 3860 -1640 3912
rect -1588 3860 -1584 3912
rect -1644 3850 -1584 3860
rect -1178 3906 -1118 4332
rect -1178 3854 -1174 3906
rect -1122 3854 -1118 3906
rect -1178 3844 -1118 3854
rect -722 3912 -662 4332
rect -488 4720 -428 4730
rect -488 4668 -484 4720
rect -432 4668 -428 4720
rect -488 4386 -428 4668
rect 1076 4386 1136 4786
rect 1538 4386 1598 4794
rect 1986 4792 1996 4844
rect 2048 4792 2058 4844
rect 1986 4788 2058 4792
rect 2448 4844 2520 4848
rect 2448 4792 2458 4844
rect 2510 4792 2520 4844
rect 2448 4788 2520 4792
rect 2902 4844 2974 4848
rect 2902 4792 2912 4844
rect 2964 4792 2974 4844
rect 3352 4798 3362 4850
rect 3414 4798 3424 4850
rect 3352 4794 3424 4798
rect 3818 4844 3890 4848
rect 2902 4788 2974 4792
rect 1992 4386 2052 4788
rect 2454 4386 2514 4788
rect 2908 4386 2968 4788
rect 3358 4386 3418 4794
rect 3818 4792 3828 4844
rect 3880 4792 3890 4844
rect 3818 4788 3890 4792
rect 4274 4844 4346 4848
rect 4274 4792 4284 4844
rect 4336 4792 4346 4844
rect 4274 4788 4346 4792
rect 3824 4386 3884 4788
rect 4280 4386 4340 4788
rect 4506 4714 4578 4718
rect 4506 4662 4516 4714
rect 4568 4662 4578 4714
rect 4506 4658 4578 4662
rect -488 4326 4340 4386
rect -488 4044 -428 4326
rect -494 4040 -422 4044
rect -494 3988 -484 4040
rect -432 3988 -422 4040
rect -494 3984 -422 3988
rect -722 3860 -718 3912
rect -666 3860 -662 3912
rect -722 3850 -662 3860
rect 1076 3912 1136 4326
rect 1076 3860 1080 3912
rect 1132 3860 1136 3912
rect 1076 3850 1136 3860
rect 1538 3910 1598 4326
rect 1538 3858 1542 3910
rect 1594 3858 1598 3910
rect 1538 3848 1598 3858
rect 1992 3910 2052 4326
rect 1992 3858 1996 3910
rect 2048 3858 2052 3910
rect 1992 3848 2052 3858
rect 2454 3910 2514 4326
rect 2454 3858 2458 3910
rect 2510 3858 2514 3910
rect 2454 3848 2514 3858
rect 2908 3910 2968 4326
rect 2908 3858 2912 3910
rect 2964 3858 2968 3910
rect 2908 3848 2968 3858
rect 3358 3916 3418 4326
rect 3358 3864 3362 3916
rect 3414 3864 3418 3916
rect 3358 3854 3418 3864
rect 3824 3912 3884 4326
rect 3824 3860 3828 3912
rect 3880 3860 3884 3912
rect 3824 3850 3884 3860
rect 4280 3912 4340 4326
rect 4512 4382 4572 4658
rect 4512 4322 5598 4382
rect 4512 4052 4572 4322
rect 5498 4193 5598 4322
rect 5494 4176 5602 4193
rect 5494 4120 5520 4176
rect 5576 4120 5602 4176
rect 5494 4103 5602 4120
rect 5498 4098 5598 4103
rect 4512 4000 4516 4052
rect 4568 4000 4572 4052
rect 4512 3990 4572 4000
rect 4280 3860 4284 3912
rect 4336 3860 4340 3912
rect 4280 3850 4340 3860
rect -4680 2433 5090 2476
rect -4680 2377 -4610 2433
rect -4554 2377 -4030 2433
rect -3974 2377 -3430 2433
rect -3374 2377 -2830 2433
rect -2774 2377 -2230 2433
rect -2174 2377 -1630 2433
rect -1574 2377 -1030 2433
rect -974 2377 -430 2433
rect -374 2377 170 2433
rect 226 2377 770 2433
rect 826 2377 1370 2433
rect 1426 2377 1970 2433
rect 2026 2377 2570 2433
rect 2626 2377 3170 2433
rect 3226 2377 3770 2433
rect 3826 2377 4370 2433
rect 4426 2377 4970 2433
rect 5026 2377 5090 2433
rect -4680 2332 5090 2377
rect -4916 2182 -4316 2194
rect -4916 2156 -4884 2182
rect -4348 2156 -4316 2182
rect -4916 1912 -4898 2156
rect -4334 1912 -4316 2156
rect -4916 1886 -4884 1912
rect -4348 1886 -4316 1912
rect -4916 1874 -4316 1886
rect 4716 2182 5316 2194
rect 4716 2156 4748 2182
rect 5284 2156 5316 2182
rect 4716 1912 4734 2156
rect 5298 1912 5316 2156
rect 4716 1886 4748 1912
rect 5284 1886 5316 1912
rect 4716 1874 5316 1886
<< via2 >>
rect -4884 10188 -4348 10214
rect -4884 9944 -4348 10188
rect -4884 9918 -4348 9944
rect 4748 10188 5284 10214
rect 4748 9944 5284 10188
rect 4748 9918 5284 9944
rect -4044 9725 -3988 9727
rect -4044 9673 -4042 9725
rect -4042 9673 -3990 9725
rect -3990 9673 -3988 9725
rect -4044 9671 -3988 9673
rect -3444 9725 -3388 9727
rect -3444 9673 -3442 9725
rect -3442 9673 -3390 9725
rect -3390 9673 -3388 9725
rect -3444 9671 -3388 9673
rect -2844 9725 -2788 9727
rect -2844 9673 -2842 9725
rect -2842 9673 -2790 9725
rect -2790 9673 -2788 9725
rect -2844 9671 -2788 9673
rect -2244 9725 -2188 9727
rect -2244 9673 -2242 9725
rect -2242 9673 -2190 9725
rect -2190 9673 -2188 9725
rect -2244 9671 -2188 9673
rect -1644 9725 -1588 9727
rect -1644 9673 -1642 9725
rect -1642 9673 -1590 9725
rect -1590 9673 -1588 9725
rect -1644 9671 -1588 9673
rect -1044 9725 -988 9727
rect -1044 9673 -1042 9725
rect -1042 9673 -990 9725
rect -990 9673 -988 9725
rect -1044 9671 -988 9673
rect -444 9725 -388 9727
rect -444 9673 -442 9725
rect -442 9673 -390 9725
rect -390 9673 -388 9725
rect -444 9671 -388 9673
rect 156 9725 212 9727
rect 156 9673 158 9725
rect 158 9673 210 9725
rect 210 9673 212 9725
rect 156 9671 212 9673
rect 756 9725 812 9727
rect 756 9673 758 9725
rect 758 9673 810 9725
rect 810 9673 812 9725
rect 756 9671 812 9673
rect 1356 9725 1412 9727
rect 1356 9673 1358 9725
rect 1358 9673 1410 9725
rect 1410 9673 1412 9725
rect 1356 9671 1412 9673
rect 1956 9725 2012 9727
rect 1956 9673 1958 9725
rect 1958 9673 2010 9725
rect 2010 9673 2012 9725
rect 1956 9671 2012 9673
rect 2556 9725 2612 9727
rect 2556 9673 2558 9725
rect 2558 9673 2610 9725
rect 2610 9673 2612 9725
rect 2556 9671 2612 9673
rect 3156 9725 3212 9727
rect 3156 9673 3158 9725
rect 3158 9673 3210 9725
rect 3210 9673 3212 9725
rect 3156 9671 3212 9673
rect 3756 9725 3812 9727
rect 3756 9673 3758 9725
rect 3758 9673 3810 9725
rect 3810 9673 3812 9725
rect 3756 9671 3812 9673
rect 4176 9725 4232 9727
rect 4176 9673 4178 9725
rect 4178 9673 4230 9725
rect 4230 9673 4232 9725
rect 4176 9671 4232 9673
rect 5520 4120 5576 4176
rect -4610 2431 -4554 2433
rect -4610 2379 -4608 2431
rect -4608 2379 -4556 2431
rect -4556 2379 -4554 2431
rect -4610 2377 -4554 2379
rect -4030 2431 -3974 2433
rect -4030 2379 -4028 2431
rect -4028 2379 -3976 2431
rect -3976 2379 -3974 2431
rect -4030 2377 -3974 2379
rect -3430 2431 -3374 2433
rect -3430 2379 -3428 2431
rect -3428 2379 -3376 2431
rect -3376 2379 -3374 2431
rect -3430 2377 -3374 2379
rect -2830 2431 -2774 2433
rect -2830 2379 -2828 2431
rect -2828 2379 -2776 2431
rect -2776 2379 -2774 2431
rect -2830 2377 -2774 2379
rect -2230 2431 -2174 2433
rect -2230 2379 -2228 2431
rect -2228 2379 -2176 2431
rect -2176 2379 -2174 2431
rect -2230 2377 -2174 2379
rect -1630 2431 -1574 2433
rect -1630 2379 -1628 2431
rect -1628 2379 -1576 2431
rect -1576 2379 -1574 2431
rect -1630 2377 -1574 2379
rect -1030 2431 -974 2433
rect -1030 2379 -1028 2431
rect -1028 2379 -976 2431
rect -976 2379 -974 2431
rect -1030 2377 -974 2379
rect -430 2431 -374 2433
rect -430 2379 -428 2431
rect -428 2379 -376 2431
rect -376 2379 -374 2431
rect -430 2377 -374 2379
rect 170 2431 226 2433
rect 170 2379 172 2431
rect 172 2379 224 2431
rect 224 2379 226 2431
rect 170 2377 226 2379
rect 770 2431 826 2433
rect 770 2379 772 2431
rect 772 2379 824 2431
rect 824 2379 826 2431
rect 770 2377 826 2379
rect 1370 2431 1426 2433
rect 1370 2379 1372 2431
rect 1372 2379 1424 2431
rect 1424 2379 1426 2431
rect 1370 2377 1426 2379
rect 1970 2431 2026 2433
rect 1970 2379 1972 2431
rect 1972 2379 2024 2431
rect 2024 2379 2026 2431
rect 1970 2377 2026 2379
rect 2570 2431 2626 2433
rect 2570 2379 2572 2431
rect 2572 2379 2624 2431
rect 2624 2379 2626 2431
rect 2570 2377 2626 2379
rect 3170 2431 3226 2433
rect 3170 2379 3172 2431
rect 3172 2379 3224 2431
rect 3224 2379 3226 2431
rect 3170 2377 3226 2379
rect 3770 2431 3826 2433
rect 3770 2379 3772 2431
rect 3772 2379 3824 2431
rect 3824 2379 3826 2431
rect 3770 2377 3826 2379
rect 4370 2431 4426 2433
rect 4370 2379 4372 2431
rect 4372 2379 4424 2431
rect 4424 2379 4426 2431
rect 4370 2377 4426 2379
rect 4970 2431 5026 2433
rect 4970 2379 4972 2431
rect 4972 2379 5024 2431
rect 5024 2379 5026 2431
rect 4970 2377 5026 2379
rect -4884 2156 -4348 2182
rect -4884 1912 -4348 2156
rect -4884 1886 -4348 1912
rect 4748 2156 5284 2182
rect 4748 1912 5284 2156
rect 4748 1886 5284 1912
<< metal3 >>
rect -4926 10214 -4306 10221
rect -4926 10178 -4884 10214
rect -4348 10178 -4306 10214
rect -4926 9954 -4888 10178
rect -4344 9954 -4306 10178
rect -4926 9918 -4884 9954
rect -4348 9918 -4306 9954
rect -4926 9911 -4306 9918
rect 4706 10214 5326 10221
rect 4706 10178 4748 10214
rect 5284 10178 5326 10214
rect 4706 9954 4744 10178
rect 5288 9954 5326 10178
rect 4706 9918 4748 9954
rect 5284 9918 5326 9954
rect 4706 9911 5326 9918
rect -4078 9731 4278 9756
rect -4078 9667 -4048 9731
rect -3984 9667 -3448 9731
rect -3384 9667 -2848 9731
rect -2784 9667 -2248 9731
rect -2184 9667 -1648 9731
rect -1584 9667 -1048 9731
rect -984 9667 -448 9731
rect -384 9667 152 9731
rect 216 9667 752 9731
rect 816 9667 1352 9731
rect 1416 9667 1952 9731
rect 2016 9667 2552 9731
rect 2616 9667 3152 9731
rect 3216 9667 3752 9731
rect 3816 9667 4172 9731
rect 4236 9667 4278 9731
rect -4078 9646 4278 9667
rect 5498 4197 5598 4198
rect 5493 4180 5603 4197
rect 5493 4116 5516 4180
rect 5580 4116 5603 4180
rect 5493 4099 5603 4116
rect 5498 4098 5598 4099
rect -4680 2437 5090 2476
rect -4680 2373 -4614 2437
rect -4550 2373 -4034 2437
rect -3970 2373 -3434 2437
rect -3370 2373 -2834 2437
rect -2770 2373 -2234 2437
rect -2170 2373 -1634 2437
rect -1570 2373 -1034 2437
rect -970 2373 -434 2437
rect -370 2373 166 2437
rect 230 2373 766 2437
rect 830 2373 1366 2437
rect 1430 2373 1966 2437
rect 2030 2373 2566 2437
rect 2630 2373 3166 2437
rect 3230 2373 3766 2437
rect 3830 2373 4366 2437
rect 4430 2373 4966 2437
rect 5030 2373 5090 2437
rect -4680 2332 5090 2373
rect -4926 2182 -4306 2189
rect -4926 2146 -4884 2182
rect -4348 2146 -4306 2182
rect -4926 1922 -4888 2146
rect -4344 1922 -4306 2146
rect -4926 1886 -4884 1922
rect -4348 1886 -4306 1922
rect -4926 1879 -4306 1886
rect 4706 2182 5326 2189
rect 4706 2146 4748 2182
rect 5284 2146 5326 2182
rect 4706 1922 4744 2146
rect 5288 1922 5326 2146
rect 5698 2064 9326 5518
rect 4706 1886 4748 1922
rect 5284 1886 5326 1922
rect 4706 1879 5326 1886
<< via3 >>
rect -4888 9954 -4884 10178
rect -4884 9954 -4348 10178
rect -4348 9954 -4344 10178
rect 4744 9954 4748 10178
rect 4748 9954 5284 10178
rect 5284 9954 5288 10178
rect -4048 9727 -3984 9731
rect -4048 9671 -4044 9727
rect -4044 9671 -3988 9727
rect -3988 9671 -3984 9727
rect -4048 9667 -3984 9671
rect -3448 9727 -3384 9731
rect -3448 9671 -3444 9727
rect -3444 9671 -3388 9727
rect -3388 9671 -3384 9727
rect -3448 9667 -3384 9671
rect -2848 9727 -2784 9731
rect -2848 9671 -2844 9727
rect -2844 9671 -2788 9727
rect -2788 9671 -2784 9727
rect -2848 9667 -2784 9671
rect -2248 9727 -2184 9731
rect -2248 9671 -2244 9727
rect -2244 9671 -2188 9727
rect -2188 9671 -2184 9727
rect -2248 9667 -2184 9671
rect -1648 9727 -1584 9731
rect -1648 9671 -1644 9727
rect -1644 9671 -1588 9727
rect -1588 9671 -1584 9727
rect -1648 9667 -1584 9671
rect -1048 9727 -984 9731
rect -1048 9671 -1044 9727
rect -1044 9671 -988 9727
rect -988 9671 -984 9727
rect -1048 9667 -984 9671
rect -448 9727 -384 9731
rect -448 9671 -444 9727
rect -444 9671 -388 9727
rect -388 9671 -384 9727
rect -448 9667 -384 9671
rect 152 9727 216 9731
rect 152 9671 156 9727
rect 156 9671 212 9727
rect 212 9671 216 9727
rect 152 9667 216 9671
rect 752 9727 816 9731
rect 752 9671 756 9727
rect 756 9671 812 9727
rect 812 9671 816 9727
rect 752 9667 816 9671
rect 1352 9727 1416 9731
rect 1352 9671 1356 9727
rect 1356 9671 1412 9727
rect 1412 9671 1416 9727
rect 1352 9667 1416 9671
rect 1952 9727 2016 9731
rect 1952 9671 1956 9727
rect 1956 9671 2012 9727
rect 2012 9671 2016 9727
rect 1952 9667 2016 9671
rect 2552 9727 2616 9731
rect 2552 9671 2556 9727
rect 2556 9671 2612 9727
rect 2612 9671 2616 9727
rect 2552 9667 2616 9671
rect 3152 9727 3216 9731
rect 3152 9671 3156 9727
rect 3156 9671 3212 9727
rect 3212 9671 3216 9727
rect 3152 9667 3216 9671
rect 3752 9727 3816 9731
rect 3752 9671 3756 9727
rect 3756 9671 3812 9727
rect 3812 9671 3816 9727
rect 3752 9667 3816 9671
rect 4172 9727 4236 9731
rect 4172 9671 4176 9727
rect 4176 9671 4232 9727
rect 4232 9671 4236 9727
rect 4172 9667 4236 9671
rect 5516 4176 5580 4180
rect 5516 4120 5520 4176
rect 5520 4120 5576 4176
rect 5576 4120 5580 4176
rect 5516 4116 5580 4120
rect -4614 2433 -4550 2437
rect -4614 2377 -4610 2433
rect -4610 2377 -4554 2433
rect -4554 2377 -4550 2433
rect -4614 2373 -4550 2377
rect -4034 2433 -3970 2437
rect -4034 2377 -4030 2433
rect -4030 2377 -3974 2433
rect -3974 2377 -3970 2433
rect -4034 2373 -3970 2377
rect -3434 2433 -3370 2437
rect -3434 2377 -3430 2433
rect -3430 2377 -3374 2433
rect -3374 2377 -3370 2433
rect -3434 2373 -3370 2377
rect -2834 2433 -2770 2437
rect -2834 2377 -2830 2433
rect -2830 2377 -2774 2433
rect -2774 2377 -2770 2433
rect -2834 2373 -2770 2377
rect -2234 2433 -2170 2437
rect -2234 2377 -2230 2433
rect -2230 2377 -2174 2433
rect -2174 2377 -2170 2433
rect -2234 2373 -2170 2377
rect -1634 2433 -1570 2437
rect -1634 2377 -1630 2433
rect -1630 2377 -1574 2433
rect -1574 2377 -1570 2433
rect -1634 2373 -1570 2377
rect -1034 2433 -970 2437
rect -1034 2377 -1030 2433
rect -1030 2377 -974 2433
rect -974 2377 -970 2433
rect -1034 2373 -970 2377
rect -434 2433 -370 2437
rect -434 2377 -430 2433
rect -430 2377 -374 2433
rect -374 2377 -370 2433
rect -434 2373 -370 2377
rect 166 2433 230 2437
rect 166 2377 170 2433
rect 170 2377 226 2433
rect 226 2377 230 2433
rect 166 2373 230 2377
rect 766 2433 830 2437
rect 766 2377 770 2433
rect 770 2377 826 2433
rect 826 2377 830 2433
rect 766 2373 830 2377
rect 1366 2433 1430 2437
rect 1366 2377 1370 2433
rect 1370 2377 1426 2433
rect 1426 2377 1430 2433
rect 1366 2373 1430 2377
rect 1966 2433 2030 2437
rect 1966 2377 1970 2433
rect 1970 2377 2026 2433
rect 2026 2377 2030 2433
rect 1966 2373 2030 2377
rect 2566 2433 2630 2437
rect 2566 2377 2570 2433
rect 2570 2377 2626 2433
rect 2626 2377 2630 2433
rect 2566 2373 2630 2377
rect 3166 2433 3230 2437
rect 3166 2377 3170 2433
rect 3170 2377 3226 2433
rect 3226 2377 3230 2433
rect 3166 2373 3230 2377
rect 3766 2433 3830 2437
rect 3766 2377 3770 2433
rect 3770 2377 3826 2433
rect 3826 2377 3830 2433
rect 3766 2373 3830 2377
rect 4366 2433 4430 2437
rect 4366 2377 4370 2433
rect 4370 2377 4426 2433
rect 4426 2377 4430 2433
rect 4366 2373 4430 2377
rect 4966 2433 5030 2437
rect 4966 2377 4970 2433
rect 4970 2377 5026 2433
rect 5026 2377 5030 2433
rect 4966 2373 5030 2377
rect -4888 1922 -4884 2146
rect -4884 1922 -4348 2146
rect -4348 1922 -4344 2146
rect 4744 1922 4748 2146
rect 4748 1922 5284 2146
rect 5284 1922 5288 2146
<< metal4 >>
rect -5100 10178 9448 10400
rect -5100 9954 -4888 10178
rect -4344 9954 4744 10178
rect 5288 9954 9448 10178
rect -5100 9731 9448 9954
rect -5100 9667 -4048 9731
rect -3984 9667 -3448 9731
rect -3384 9667 -2848 9731
rect -2784 9667 -2248 9731
rect -2184 9667 -1648 9731
rect -1584 9667 -1048 9731
rect -984 9667 -448 9731
rect -384 9667 152 9731
rect 216 9667 752 9731
rect 816 9667 1352 9731
rect 1416 9667 1952 9731
rect 2016 9667 2552 9731
rect 2616 9667 3152 9731
rect 3216 9667 3752 9731
rect 3816 9667 4172 9731
rect 4236 9667 9448 9731
rect -5100 9600 9448 9667
rect 5974 5144 9288 5244
rect 5974 4554 6074 5144
rect 6310 4554 6410 5144
rect 5974 4454 6410 4554
rect 5974 4340 6074 4454
rect 6310 4340 6410 4454
rect 6688 4790 8232 4890
rect 6688 4198 6788 4790
rect 7408 4198 7508 4790
rect 8130 4198 8231 4790
rect 8476 4555 8578 5144
rect 8478 4550 8578 4555
rect 8850 4550 8950 5144
rect 9188 5089 9288 5144
rect 9188 4594 9291 5089
rect 9188 4550 9288 4594
rect 8478 4450 9288 4550
rect 8478 4300 8578 4450
rect 8850 4338 8950 4450
rect 9188 4300 9288 4450
rect 5498 4180 9450 4198
rect 5498 4116 5516 4180
rect 5580 4116 9450 4180
rect 5498 4098 9450 4116
rect 5974 3852 6074 3962
rect 6310 3852 6410 3962
rect 5974 3752 6410 3852
rect 5974 3146 6074 3752
rect 6310 3146 6410 3752
rect 5974 3046 6410 3146
rect 5974 2500 6074 3046
rect 6310 2500 6410 3046
rect 6688 3496 6788 4098
rect 7408 3496 7508 4098
rect 8130 3496 8231 4098
rect 6688 3396 8231 3496
rect 6688 2796 6788 3396
rect 7408 2796 7508 3396
rect 8130 2796 8231 3396
rect 8478 3846 8578 4000
rect 8850 3846 8950 3962
rect 9188 3846 9288 4000
rect 8478 3746 9288 3846
rect 8478 3154 8578 3746
rect 8850 3154 8950 3746
rect 9188 3154 9288 3746
rect 8478 3054 9288 3154
rect 8478 2995 8578 3054
rect 6688 2696 8232 2796
rect 8476 2500 8578 2995
rect 8850 2500 8950 3054
rect 9188 3035 9288 3054
rect 9188 2500 9291 3035
rect -5100 2437 9448 2500
rect -5100 2373 -4614 2437
rect -4550 2373 -4034 2437
rect -3970 2373 -3434 2437
rect -3370 2373 -2834 2437
rect -2770 2373 -2234 2437
rect -2170 2373 -1634 2437
rect -1570 2373 -1034 2437
rect -970 2373 -434 2437
rect -370 2373 166 2437
rect 230 2373 766 2437
rect 830 2373 1366 2437
rect 1430 2373 1966 2437
rect 2030 2373 2566 2437
rect 2630 2373 3166 2437
rect 3230 2373 3766 2437
rect 3830 2373 4366 2437
rect 4430 2373 4966 2437
rect 5030 2373 9448 2437
rect -5100 2146 9448 2373
rect -5100 1922 -4888 2146
rect -4344 1922 4744 2146
rect 5288 1922 9448 2146
rect -5100 1700 9448 1922
rect 8478 1696 8578 1700
use sky130_fd_pr__cap_mim_m3_1_FAR8MD  sky130_fd_pr__cap_mim_m3_1_FAR8MD_0
timestamp 1626486988
transform 1 0 7508 0 1 3800
box -1788 -1700 1787 1700
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_0
timestamp 1626486988
transform 1 0 2711 0 1 3612
box -2345 -188 2345 188
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_1
timestamp 1626486988
transform 1 0 -2289 0 1 3612
box -2345 -188 2345 188
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_2
timestamp 1626486988
transform 1 0 -2289 0 1 2944
box -2345 -188 2345 188
use sky130_fd_pr__pfet_01v8_hvt_GK2P2M  sky130_fd_pr__pfet_01v8_hvt_GK2P2M_0
timestamp 1626486988
transform 1 0 103 0 1 8070
box -4187 -900 4187 900
use sky130_fd_pr__pfet_01v8_hvt_8Q5PU3  sky130_fd_pr__pfet_01v8_hvt_8Q5PU3_0
timestamp 1626486988
transform 1 0 -2288 0 1 5605
box -2355 -700 2355 700
use sky130_fd_pr__pfet_01v8_hvt_8Q5PU3  sky130_fd_pr__pfet_01v8_hvt_8Q5PU3_1
timestamp 1626486988
transform 1 0 2712 0 1 5605
box -2355 -700 2355 700
<< labels >>
flabel metal4 s -2300 2102 -2280 2122 1 FreeSans 600 0 0 0 VSS
flabel metal4 s -2534 10006 -2500 10030 1 FreeSans 600 0 0 0 VDD
flabel metal2 s -3700 4356 -3686 4370 1 FreeSans 600 0 0 0 vin
flabel metal1 s -3698 2662 -3690 2672 1 FreeSans 600 0 0 0 vbiasn
flabel metal2 s -3228 7078 -3218 7084 1 FreeSans 600 0 0 0 vbiasp
flabel metal2 s 4126 4350 4138 4364 1 FreeSans 600 0 0 0 voutcs
flabel metal2 s 4532 4380 4544 4390 1 FreeSans 600 0 0 0 vout
flabel metal1 s -4134 3252 -4122 3270 1 FreeSans 600 0 0 0 csinvn
flabel metal2 s -3584 6480 -3574 6494 1 FreeSans 600 0 0 0 csinvp
<< properties >>
string FIXED_BBOX -4972 1328 5372 4032
<< end >>
