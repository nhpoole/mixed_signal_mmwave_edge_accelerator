magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -262 -1256 81981 3271
rect 114 -1260 81981 -1256
<< metal1 >>
rect 1500 1959 1530 2011
rect 1702 1959 1732 2011
rect 3996 1959 4026 2011
rect 4198 1959 4228 2011
rect 6492 1959 6522 2011
rect 6694 1959 6724 2011
rect 8988 1959 9018 2011
rect 9190 1959 9220 2011
rect 11484 1959 11514 2011
rect 11686 1959 11716 2011
rect 13980 1959 14010 2011
rect 14182 1959 14212 2011
rect 16476 1959 16506 2011
rect 16678 1959 16708 2011
rect 18972 1959 19002 2011
rect 19174 1959 19204 2011
rect 21468 1959 21498 2011
rect 21670 1959 21700 2011
rect 23964 1959 23994 2011
rect 24166 1959 24196 2011
rect 26460 1959 26490 2011
rect 26662 1959 26692 2011
rect 28956 1959 28986 2011
rect 29158 1959 29188 2011
rect 31452 1959 31482 2011
rect 31654 1959 31684 2011
rect 33948 1959 33978 2011
rect 34150 1959 34180 2011
rect 36444 1959 36474 2011
rect 36646 1959 36676 2011
rect 38940 1959 38970 2011
rect 39142 1959 39172 2011
rect 41436 1959 41466 2011
rect 41638 1959 41668 2011
rect 43932 1959 43962 2011
rect 44134 1959 44164 2011
rect 46428 1959 46458 2011
rect 46630 1959 46660 2011
rect 48924 1959 48954 2011
rect 49126 1959 49156 2011
rect 51420 1959 51450 2011
rect 51622 1959 51652 2011
rect 53916 1959 53946 2011
rect 54118 1959 54148 2011
rect 56412 1959 56442 2011
rect 56614 1959 56644 2011
rect 58908 1959 58938 2011
rect 59110 1959 59140 2011
rect 61404 1959 61434 2011
rect 61606 1959 61636 2011
rect 63900 1959 63930 2011
rect 64102 1959 64132 2011
rect 66396 1959 66426 2011
rect 66598 1959 66628 2011
rect 68892 1959 68922 2011
rect 69094 1959 69124 2011
rect 71388 1959 71418 2011
rect 71590 1959 71620 2011
rect 73884 1959 73914 2011
rect 74086 1959 74116 2011
rect 76380 1959 76410 2011
rect 76582 1959 76612 2011
rect 78876 1959 78906 2011
rect 79078 1959 79108 2011
rect 1473 94 20817 128
rect 21441 94 40785 128
rect 41409 94 60753 128
rect 61377 94 80721 128
rect 1629 4 1689 60
rect 4125 4 4185 60
rect 6621 4 6681 60
rect 9117 4 9177 60
rect 11613 4 11673 60
rect 14109 4 14169 60
rect 16605 4 16665 60
rect 19101 4 19161 60
rect 21597 4 21657 60
rect 24093 4 24153 60
rect 26589 4 26649 60
rect 29085 4 29145 60
rect 31581 4 31641 60
rect 34077 4 34137 60
rect 36573 4 36633 60
rect 39069 4 39129 60
rect 41565 4 41625 60
rect 44061 4 44121 60
rect 46557 4 46617 60
rect 49053 4 49113 60
rect 51549 4 51609 60
rect 54045 4 54105 60
rect 56541 4 56601 60
rect 59037 4 59097 60
rect 61533 4 61593 60
rect 64029 4 64089 60
rect 66525 4 66585 60
rect 69021 4 69081 60
rect 71517 4 71577 60
rect 74013 4 74073 60
rect 76509 4 76569 60
rect 79005 4 79065 60
<< metal2 >>
rect 1613 1554 1669 1602
rect 4109 1554 4165 1602
rect 6605 1554 6661 1602
rect 9101 1554 9157 1602
rect 11597 1554 11653 1602
rect 14093 1554 14149 1602
rect 16589 1554 16645 1602
rect 19085 1554 19141 1602
rect 21581 1554 21637 1602
rect 24077 1554 24133 1602
rect 26573 1554 26629 1602
rect 29069 1554 29125 1602
rect 31565 1554 31621 1602
rect 34061 1554 34117 1602
rect 36557 1554 36613 1602
rect 39053 1554 39109 1602
rect 41549 1554 41605 1602
rect 44045 1554 44101 1602
rect 46541 1554 46597 1602
rect 49037 1554 49093 1602
rect 51533 1554 51589 1602
rect 54029 1554 54085 1602
rect 56525 1554 56581 1602
rect 59021 1554 59077 1602
rect 61517 1554 61573 1602
rect 64013 1554 64069 1602
rect 66509 1554 66565 1602
rect 69005 1554 69061 1602
rect 71501 1554 71557 1602
rect 73997 1554 74053 1602
rect 76493 1554 76549 1602
rect 78989 1554 79045 1602
rect 1602 1117 1658 1165
rect 4098 1117 4154 1165
rect 6594 1117 6650 1165
rect 9090 1117 9146 1165
rect 11586 1117 11642 1165
rect 14082 1117 14138 1165
rect 16578 1117 16634 1165
rect 19074 1117 19130 1165
rect 21570 1117 21626 1165
rect 24066 1117 24122 1165
rect 26562 1117 26618 1165
rect 29058 1117 29114 1165
rect 31554 1117 31610 1165
rect 34050 1117 34106 1165
rect 36546 1117 36602 1165
rect 39042 1117 39098 1165
rect 41538 1117 41594 1165
rect 44034 1117 44090 1165
rect 46530 1117 46586 1165
rect 49026 1117 49082 1165
rect 51522 1117 51578 1165
rect 54018 1117 54074 1165
rect 56514 1117 56570 1165
rect 59010 1117 59066 1165
rect 61506 1117 61562 1165
rect 64002 1117 64058 1165
rect 66498 1117 66554 1165
rect 68994 1117 69050 1165
rect 71490 1117 71546 1165
rect 73986 1117 74042 1165
rect 76482 1117 76538 1165
rect 78978 1117 79034 1165
rect 1723 785 1779 833
rect 4219 785 4275 833
rect 6715 785 6771 833
rect 9211 785 9267 833
rect 11707 785 11763 833
rect 14203 785 14259 833
rect 16699 785 16755 833
rect 19195 785 19251 833
rect 21691 785 21747 833
rect 24187 785 24243 833
rect 26683 785 26739 833
rect 29179 785 29235 833
rect 31675 785 31731 833
rect 34171 785 34227 833
rect 36667 785 36723 833
rect 39163 785 39219 833
rect 41659 785 41715 833
rect 44155 785 44211 833
rect 46651 785 46707 833
rect 49147 785 49203 833
rect 51643 785 51699 833
rect 54139 785 54195 833
rect 56635 785 56691 833
rect 59131 785 59187 833
rect 61627 785 61683 833
rect 64123 785 64179 833
rect 66619 785 66675 833
rect 69115 785 69171 833
rect 71611 785 71667 833
rect 74107 785 74163 833
rect 76603 785 76659 833
rect 79099 785 79155 833
rect 1608 583 1664 631
rect 4104 583 4160 631
rect 6600 583 6656 631
rect 9096 583 9152 631
rect 11592 583 11648 631
rect 14088 583 14144 631
rect 16584 583 16640 631
rect 19080 583 19136 631
rect 21576 583 21632 631
rect 24072 583 24128 631
rect 26568 583 26624 631
rect 29064 583 29120 631
rect 31560 583 31616 631
rect 34056 583 34112 631
rect 36552 583 36608 631
rect 39048 583 39104 631
rect 41544 583 41600 631
rect 44040 583 44096 631
rect 46536 583 46592 631
rect 49032 583 49088 631
rect 51528 583 51584 631
rect 54024 583 54080 631
rect 56520 583 56576 631
rect 59016 583 59072 631
rect 61512 583 61568 631
rect 64008 583 64064 631
rect 66504 583 66560 631
rect 69000 583 69056 631
rect 71496 583 71552 631
rect 73992 583 74048 631
rect 76488 583 76544 631
rect 78984 583 79040 631
rect 1622 167 1678 215
rect 4118 167 4174 215
rect 6614 167 6670 215
rect 9110 167 9166 215
rect 11606 167 11662 215
rect 14102 167 14158 215
rect 16598 167 16654 215
rect 19094 167 19150 215
rect 21590 167 21646 215
rect 24086 167 24142 215
rect 26582 167 26638 215
rect 29078 167 29134 215
rect 31574 167 31630 215
rect 34070 167 34126 215
rect 36566 167 36622 215
rect 39062 167 39118 215
rect 41558 167 41614 215
rect 44054 167 44110 215
rect 46550 167 46606 215
rect 49046 167 49102 215
rect 51542 167 51598 215
rect 54038 167 54094 215
rect 56534 167 56590 215
rect 59030 167 59086 215
rect 61526 167 61582 215
rect 64022 167 64078 215
rect 66518 167 66574 215
rect 69014 167 69070 215
rect 71510 167 71566 215
rect 74006 167 74062 215
rect 76502 167 76558 215
rect 78998 167 79054 215
<< metal3 >>
rect 1592 1529 1690 1627
rect 4088 1529 4186 1627
rect 6584 1529 6682 1627
rect 9080 1529 9178 1627
rect 11576 1529 11674 1627
rect 14072 1529 14170 1627
rect 16568 1529 16666 1627
rect 19064 1529 19162 1627
rect 21560 1529 21658 1627
rect 24056 1529 24154 1627
rect 26552 1529 26650 1627
rect 29048 1529 29146 1627
rect 31544 1529 31642 1627
rect 34040 1529 34138 1627
rect 36536 1529 36634 1627
rect 39032 1529 39130 1627
rect 41528 1529 41626 1627
rect 44024 1529 44122 1627
rect 46520 1529 46618 1627
rect 49016 1529 49114 1627
rect 51512 1529 51610 1627
rect 54008 1529 54106 1627
rect 56504 1529 56602 1627
rect 59000 1529 59098 1627
rect 61496 1529 61594 1627
rect 63992 1529 64090 1627
rect 66488 1529 66586 1627
rect 68984 1529 69082 1627
rect 71480 1529 71578 1627
rect 73976 1529 74074 1627
rect 76472 1529 76570 1627
rect 78968 1529 79066 1627
rect 1581 1092 1679 1190
rect 4077 1092 4175 1190
rect 6573 1092 6671 1190
rect 9069 1092 9167 1190
rect 11565 1092 11663 1190
rect 14061 1092 14159 1190
rect 16557 1092 16655 1190
rect 19053 1092 19151 1190
rect 21549 1092 21647 1190
rect 24045 1092 24143 1190
rect 26541 1092 26639 1190
rect 29037 1092 29135 1190
rect 31533 1092 31631 1190
rect 34029 1092 34127 1190
rect 36525 1092 36623 1190
rect 39021 1092 39119 1190
rect 41517 1092 41615 1190
rect 44013 1092 44111 1190
rect 46509 1092 46607 1190
rect 49005 1092 49103 1190
rect 51501 1092 51599 1190
rect 53997 1092 54095 1190
rect 56493 1092 56591 1190
rect 58989 1092 59087 1190
rect 61485 1092 61583 1190
rect 63981 1092 64079 1190
rect 66477 1092 66575 1190
rect 68973 1092 69071 1190
rect 71469 1092 71567 1190
rect 73965 1092 74063 1190
rect 76461 1092 76559 1190
rect 78957 1092 79055 1190
rect 1702 760 1800 858
rect 4198 760 4296 858
rect 6694 760 6792 858
rect 9190 760 9288 858
rect 11686 760 11784 858
rect 14182 760 14280 858
rect 16678 760 16776 858
rect 19174 760 19272 858
rect 21670 760 21768 858
rect 24166 760 24264 858
rect 26662 760 26760 858
rect 29158 760 29256 858
rect 31654 760 31752 858
rect 34150 760 34248 858
rect 36646 760 36744 858
rect 39142 760 39240 858
rect 41638 760 41736 858
rect 44134 760 44232 858
rect 46630 760 46728 858
rect 49126 760 49224 858
rect 51622 760 51720 858
rect 54118 760 54216 858
rect 56614 760 56712 858
rect 59110 760 59208 858
rect 61606 760 61704 858
rect 64102 760 64200 858
rect 66598 760 66696 858
rect 69094 760 69192 858
rect 71590 760 71688 858
rect 74086 760 74184 858
rect 76582 760 76680 858
rect 79078 760 79176 858
rect 1587 558 1685 656
rect 4083 558 4181 656
rect 6579 558 6677 656
rect 9075 558 9173 656
rect 11571 558 11669 656
rect 14067 558 14165 656
rect 16563 558 16661 656
rect 19059 558 19157 656
rect 21555 558 21653 656
rect 24051 558 24149 656
rect 26547 558 26645 656
rect 29043 558 29141 656
rect 31539 558 31637 656
rect 34035 558 34133 656
rect 36531 558 36629 656
rect 39027 558 39125 656
rect 41523 558 41621 656
rect 44019 558 44117 656
rect 46515 558 46613 656
rect 49011 558 49109 656
rect 51507 558 51605 656
rect 54003 558 54101 656
rect 56499 558 56597 656
rect 58995 558 59093 656
rect 61491 558 61589 656
rect 63987 558 64085 656
rect 66483 558 66581 656
rect 68979 558 69077 656
rect 71475 558 71573 656
rect 73971 558 74069 656
rect 76467 558 76565 656
rect 78963 558 79061 656
rect 1601 142 1699 240
rect 4097 142 4195 240
rect 6593 142 6691 240
rect 9089 142 9187 240
rect 11585 142 11683 240
rect 14081 142 14179 240
rect 16577 142 16675 240
rect 19073 142 19171 240
rect 21569 142 21667 240
rect 24065 142 24163 240
rect 26561 142 26659 240
rect 29057 142 29155 240
rect 31553 142 31651 240
rect 34049 142 34147 240
rect 36545 142 36643 240
rect 39041 142 39139 240
rect 41537 142 41635 240
rect 44033 142 44131 240
rect 46529 142 46627 240
rect 49025 142 49123 240
rect 51521 142 51619 240
rect 54017 142 54115 240
rect 56513 142 56611 240
rect 59009 142 59107 240
rect 61505 142 61603 240
rect 64001 142 64099 240
rect 66497 142 66595 240
rect 68993 142 69091 240
rect 71489 142 71587 240
rect 73985 142 74083 240
rect 76481 142 76579 240
rect 78977 142 79075 240
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_159
timestamp 1626486988
transform 1 0 61521 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_158
timestamp 1626486988
transform 1 0 61501 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_157
timestamp 1626486988
transform 1 0 61507 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_156
timestamp 1626486988
transform 1 0 61622 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_155
timestamp 1626486988
transform 1 0 61512 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_154
timestamp 1626486988
transform 1 0 64017 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_153
timestamp 1626486988
transform 1 0 63997 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_152
timestamp 1626486988
transform 1 0 64003 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_151
timestamp 1626486988
transform 1 0 64118 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_150
timestamp 1626486988
transform 1 0 64008 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_149
timestamp 1626486988
transform 1 0 66513 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_148
timestamp 1626486988
transform 1 0 66493 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_147
timestamp 1626486988
transform 1 0 66499 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_146
timestamp 1626486988
transform 1 0 66614 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_145
timestamp 1626486988
transform 1 0 66504 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_144
timestamp 1626486988
transform 1 0 69009 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_143
timestamp 1626486988
transform 1 0 68989 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_142
timestamp 1626486988
transform 1 0 68995 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_141
timestamp 1626486988
transform 1 0 69110 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_140
timestamp 1626486988
transform 1 0 69000 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_139
timestamp 1626486988
transform 1 0 71505 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_138
timestamp 1626486988
transform 1 0 71485 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_137
timestamp 1626486988
transform 1 0 71491 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_136
timestamp 1626486988
transform 1 0 71606 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_135
timestamp 1626486988
transform 1 0 71496 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_134
timestamp 1626486988
transform 1 0 74001 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_133
timestamp 1626486988
transform 1 0 73981 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_132
timestamp 1626486988
transform 1 0 73987 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_131
timestamp 1626486988
transform 1 0 74102 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_130
timestamp 1626486988
transform 1 0 73992 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_129
timestamp 1626486988
transform 1 0 76497 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_128
timestamp 1626486988
transform 1 0 76477 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_127
timestamp 1626486988
transform 1 0 76483 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_126
timestamp 1626486988
transform 1 0 76598 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_125
timestamp 1626486988
transform 1 0 76488 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_124
timestamp 1626486988
transform 1 0 78993 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_123
timestamp 1626486988
transform 1 0 78973 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_122
timestamp 1626486988
transform 1 0 78979 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_121
timestamp 1626486988
transform 1 0 79094 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_120
timestamp 1626486988
transform 1 0 78984 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_119
timestamp 1626486988
transform 1 0 59005 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_118
timestamp 1626486988
transform 1 0 59011 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_117
timestamp 1626486988
transform 1 0 59126 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_116
timestamp 1626486988
transform 1 0 59016 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_115
timestamp 1626486988
transform 1 0 41553 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_114
timestamp 1626486988
transform 1 0 41533 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_113
timestamp 1626486988
transform 1 0 41539 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_112
timestamp 1626486988
transform 1 0 41654 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_111
timestamp 1626486988
transform 1 0 41544 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_110
timestamp 1626486988
transform 1 0 44049 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_109
timestamp 1626486988
transform 1 0 44029 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_108
timestamp 1626486988
transform 1 0 44035 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_107
timestamp 1626486988
transform 1 0 44150 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_106
timestamp 1626486988
transform 1 0 44040 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_105
timestamp 1626486988
transform 1 0 46545 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_104
timestamp 1626486988
transform 1 0 46525 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_103
timestamp 1626486988
transform 1 0 46531 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_102
timestamp 1626486988
transform 1 0 46646 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_101
timestamp 1626486988
transform 1 0 46536 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_100
timestamp 1626486988
transform 1 0 49041 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_99
timestamp 1626486988
transform 1 0 49021 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_98
timestamp 1626486988
transform 1 0 49027 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_97
timestamp 1626486988
transform 1 0 49142 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_96
timestamp 1626486988
transform 1 0 49032 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_95
timestamp 1626486988
transform 1 0 51537 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_94
timestamp 1626486988
transform 1 0 51517 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_93
timestamp 1626486988
transform 1 0 51523 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_92
timestamp 1626486988
transform 1 0 51638 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_91
timestamp 1626486988
transform 1 0 51528 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_90
timestamp 1626486988
transform 1 0 54033 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_89
timestamp 1626486988
transform 1 0 54013 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_88
timestamp 1626486988
transform 1 0 54019 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_87
timestamp 1626486988
transform 1 0 54134 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_86
timestamp 1626486988
transform 1 0 54024 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_85
timestamp 1626486988
transform 1 0 56529 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_84
timestamp 1626486988
transform 1 0 56509 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_83
timestamp 1626486988
transform 1 0 56515 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_82
timestamp 1626486988
transform 1 0 56630 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_81
timestamp 1626486988
transform 1 0 56520 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_80
timestamp 1626486988
transform 1 0 59025 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_79
timestamp 1626486988
transform 1 0 36547 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_78
timestamp 1626486988
transform 1 0 36662 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_77
timestamp 1626486988
transform 1 0 36552 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_76
timestamp 1626486988
transform 1 0 39057 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_75
timestamp 1626486988
transform 1 0 39037 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_74
timestamp 1626486988
transform 1 0 39043 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_73
timestamp 1626486988
transform 1 0 39158 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_72
timestamp 1626486988
transform 1 0 39048 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_71
timestamp 1626486988
transform 1 0 21585 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_70
timestamp 1626486988
transform 1 0 21565 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_69
timestamp 1626486988
transform 1 0 21571 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_68
timestamp 1626486988
transform 1 0 21686 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_67
timestamp 1626486988
transform 1 0 21576 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_66
timestamp 1626486988
transform 1 0 24081 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_65
timestamp 1626486988
transform 1 0 24061 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_64
timestamp 1626486988
transform 1 0 24067 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_63
timestamp 1626486988
transform 1 0 24182 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_62
timestamp 1626486988
transform 1 0 24072 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_61
timestamp 1626486988
transform 1 0 26577 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_60
timestamp 1626486988
transform 1 0 26557 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_59
timestamp 1626486988
transform 1 0 26563 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_58
timestamp 1626486988
transform 1 0 26678 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_57
timestamp 1626486988
transform 1 0 26568 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_56
timestamp 1626486988
transform 1 0 29073 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_55
timestamp 1626486988
transform 1 0 29053 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_54
timestamp 1626486988
transform 1 0 29059 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_53
timestamp 1626486988
transform 1 0 29174 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_52
timestamp 1626486988
transform 1 0 29064 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_51
timestamp 1626486988
transform 1 0 31569 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_50
timestamp 1626486988
transform 1 0 31549 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_49
timestamp 1626486988
transform 1 0 31555 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_48
timestamp 1626486988
transform 1 0 31670 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_47
timestamp 1626486988
transform 1 0 31560 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_46
timestamp 1626486988
transform 1 0 34065 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_45
timestamp 1626486988
transform 1 0 34045 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_44
timestamp 1626486988
transform 1 0 34051 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_43
timestamp 1626486988
transform 1 0 34166 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_42
timestamp 1626486988
transform 1 0 34056 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_41
timestamp 1626486988
transform 1 0 36561 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_40
timestamp 1626486988
transform 1 0 36541 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_39
timestamp 1626486988
transform 1 0 14198 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_38
timestamp 1626486988
transform 1 0 14088 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_37
timestamp 1626486988
transform 1 0 16593 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_36
timestamp 1626486988
transform 1 0 16573 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_35
timestamp 1626486988
transform 1 0 16579 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_34
timestamp 1626486988
transform 1 0 16694 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_33
timestamp 1626486988
transform 1 0 16584 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_32
timestamp 1626486988
transform 1 0 19089 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_31
timestamp 1626486988
transform 1 0 19069 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_30
timestamp 1626486988
transform 1 0 19075 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_29
timestamp 1626486988
transform 1 0 19190 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_28
timestamp 1626486988
transform 1 0 19080 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_27
timestamp 1626486988
transform 1 0 1617 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_26
timestamp 1626486988
transform 1 0 1597 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_25
timestamp 1626486988
transform 1 0 1603 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_24
timestamp 1626486988
transform 1 0 1718 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_23
timestamp 1626486988
transform 1 0 1608 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_22
timestamp 1626486988
transform 1 0 4113 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_21
timestamp 1626486988
transform 1 0 4093 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_20
timestamp 1626486988
transform 1 0 4099 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_19
timestamp 1626486988
transform 1 0 4214 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_18
timestamp 1626486988
transform 1 0 4104 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_17
timestamp 1626486988
transform 1 0 6609 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_16
timestamp 1626486988
transform 1 0 6589 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_15
timestamp 1626486988
transform 1 0 6595 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_14
timestamp 1626486988
transform 1 0 6710 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_13
timestamp 1626486988
transform 1 0 6600 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_12
timestamp 1626486988
transform 1 0 9105 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_11
timestamp 1626486988
transform 1 0 9085 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_10
timestamp 1626486988
transform 1 0 9091 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_9
timestamp 1626486988
transform 1 0 9206 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_8
timestamp 1626486988
transform 1 0 9096 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_7
timestamp 1626486988
transform 1 0 11601 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_6
timestamp 1626486988
transform 1 0 11581 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_5
timestamp 1626486988
transform 1 0 11587 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_4
timestamp 1626486988
transform 1 0 11702 0 1 772
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_3
timestamp 1626486988
transform 1 0 11592 0 1 1541
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_2
timestamp 1626486988
transform 1 0 14097 0 1 154
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_1
timestamp 1626486988
transform 1 0 14077 0 1 1104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_0
timestamp 1626486988
transform 1 0 14083 0 1 570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_159
timestamp 1626486988
transform 1 0 61528 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_158
timestamp 1626486988
transform 1 0 61508 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_157
timestamp 1626486988
transform 1 0 61514 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_156
timestamp 1626486988
transform 1 0 61629 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_155
timestamp 1626486988
transform 1 0 61519 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_154
timestamp 1626486988
transform 1 0 64024 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_153
timestamp 1626486988
transform 1 0 64004 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_152
timestamp 1626486988
transform 1 0 64010 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_151
timestamp 1626486988
transform 1 0 64125 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_150
timestamp 1626486988
transform 1 0 64015 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_149
timestamp 1626486988
transform 1 0 66520 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_148
timestamp 1626486988
transform 1 0 66500 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_147
timestamp 1626486988
transform 1 0 66506 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_146
timestamp 1626486988
transform 1 0 66621 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_145
timestamp 1626486988
transform 1 0 66511 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_144
timestamp 1626486988
transform 1 0 69016 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_143
timestamp 1626486988
transform 1 0 68996 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_142
timestamp 1626486988
transform 1 0 69002 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_141
timestamp 1626486988
transform 1 0 69117 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_140
timestamp 1626486988
transform 1 0 69007 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_139
timestamp 1626486988
transform 1 0 71512 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_138
timestamp 1626486988
transform 1 0 71492 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_137
timestamp 1626486988
transform 1 0 71498 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_136
timestamp 1626486988
transform 1 0 71613 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_135
timestamp 1626486988
transform 1 0 71503 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_134
timestamp 1626486988
transform 1 0 74008 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_133
timestamp 1626486988
transform 1 0 73988 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_132
timestamp 1626486988
transform 1 0 73994 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_131
timestamp 1626486988
transform 1 0 74109 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_130
timestamp 1626486988
transform 1 0 73999 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_129
timestamp 1626486988
transform 1 0 76504 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_128
timestamp 1626486988
transform 1 0 76484 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_127
timestamp 1626486988
transform 1 0 76490 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_126
timestamp 1626486988
transform 1 0 76605 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_125
timestamp 1626486988
transform 1 0 76495 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_124
timestamp 1626486988
transform 1 0 79000 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_123
timestamp 1626486988
transform 1 0 78980 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_122
timestamp 1626486988
transform 1 0 78986 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_121
timestamp 1626486988
transform 1 0 79101 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_120
timestamp 1626486988
transform 1 0 78991 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_119
timestamp 1626486988
transform 1 0 59012 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_118
timestamp 1626486988
transform 1 0 59018 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_117
timestamp 1626486988
transform 1 0 59133 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_116
timestamp 1626486988
transform 1 0 59023 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_115
timestamp 1626486988
transform 1 0 41560 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_114
timestamp 1626486988
transform 1 0 41540 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_113
timestamp 1626486988
transform 1 0 41546 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_112
timestamp 1626486988
transform 1 0 41661 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_111
timestamp 1626486988
transform 1 0 41551 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_110
timestamp 1626486988
transform 1 0 44056 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_109
timestamp 1626486988
transform 1 0 44036 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_108
timestamp 1626486988
transform 1 0 44042 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_107
timestamp 1626486988
transform 1 0 44157 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_106
timestamp 1626486988
transform 1 0 44047 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_105
timestamp 1626486988
transform 1 0 46552 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_104
timestamp 1626486988
transform 1 0 46532 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_103
timestamp 1626486988
transform 1 0 46538 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_102
timestamp 1626486988
transform 1 0 46653 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_101
timestamp 1626486988
transform 1 0 46543 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_100
timestamp 1626486988
transform 1 0 49048 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_99
timestamp 1626486988
transform 1 0 49028 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_98
timestamp 1626486988
transform 1 0 49034 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_97
timestamp 1626486988
transform 1 0 49149 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_96
timestamp 1626486988
transform 1 0 49039 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_95
timestamp 1626486988
transform 1 0 51544 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_94
timestamp 1626486988
transform 1 0 51524 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_93
timestamp 1626486988
transform 1 0 51530 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_92
timestamp 1626486988
transform 1 0 51645 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_91
timestamp 1626486988
transform 1 0 51535 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_90
timestamp 1626486988
transform 1 0 54040 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_89
timestamp 1626486988
transform 1 0 54020 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_88
timestamp 1626486988
transform 1 0 54026 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_87
timestamp 1626486988
transform 1 0 54141 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_86
timestamp 1626486988
transform 1 0 54031 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_85
timestamp 1626486988
transform 1 0 56536 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_84
timestamp 1626486988
transform 1 0 56516 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_83
timestamp 1626486988
transform 1 0 56522 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_82
timestamp 1626486988
transform 1 0 56637 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_81
timestamp 1626486988
transform 1 0 56527 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_80
timestamp 1626486988
transform 1 0 59032 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_79
timestamp 1626486988
transform 1 0 36554 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_78
timestamp 1626486988
transform 1 0 36669 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_77
timestamp 1626486988
transform 1 0 36559 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_76
timestamp 1626486988
transform 1 0 39064 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_75
timestamp 1626486988
transform 1 0 39044 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_74
timestamp 1626486988
transform 1 0 39050 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_73
timestamp 1626486988
transform 1 0 39165 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_72
timestamp 1626486988
transform 1 0 39055 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_71
timestamp 1626486988
transform 1 0 21592 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_70
timestamp 1626486988
transform 1 0 21572 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_69
timestamp 1626486988
transform 1 0 21578 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_68
timestamp 1626486988
transform 1 0 21693 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_67
timestamp 1626486988
transform 1 0 21583 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_66
timestamp 1626486988
transform 1 0 24088 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_65
timestamp 1626486988
transform 1 0 24068 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_64
timestamp 1626486988
transform 1 0 24074 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_63
timestamp 1626486988
transform 1 0 24189 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_62
timestamp 1626486988
transform 1 0 24079 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_61
timestamp 1626486988
transform 1 0 26584 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_60
timestamp 1626486988
transform 1 0 26564 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_59
timestamp 1626486988
transform 1 0 26570 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_58
timestamp 1626486988
transform 1 0 26685 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_57
timestamp 1626486988
transform 1 0 26575 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_56
timestamp 1626486988
transform 1 0 29080 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_55
timestamp 1626486988
transform 1 0 29060 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_54
timestamp 1626486988
transform 1 0 29066 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_53
timestamp 1626486988
transform 1 0 29181 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_52
timestamp 1626486988
transform 1 0 29071 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_51
timestamp 1626486988
transform 1 0 31576 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_50
timestamp 1626486988
transform 1 0 31556 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_49
timestamp 1626486988
transform 1 0 31562 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_48
timestamp 1626486988
transform 1 0 31677 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_47
timestamp 1626486988
transform 1 0 31567 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_46
timestamp 1626486988
transform 1 0 34072 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_45
timestamp 1626486988
transform 1 0 34052 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_44
timestamp 1626486988
transform 1 0 34058 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_43
timestamp 1626486988
transform 1 0 34173 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_42
timestamp 1626486988
transform 1 0 34063 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_41
timestamp 1626486988
transform 1 0 36568 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_40
timestamp 1626486988
transform 1 0 36548 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_39
timestamp 1626486988
transform 1 0 14205 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_38
timestamp 1626486988
transform 1 0 14095 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_37
timestamp 1626486988
transform 1 0 16600 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_36
timestamp 1626486988
transform 1 0 16580 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_35
timestamp 1626486988
transform 1 0 16586 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_34
timestamp 1626486988
transform 1 0 16701 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_33
timestamp 1626486988
transform 1 0 16591 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_32
timestamp 1626486988
transform 1 0 19096 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_31
timestamp 1626486988
transform 1 0 19076 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_30
timestamp 1626486988
transform 1 0 19082 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_29
timestamp 1626486988
transform 1 0 19197 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_28
timestamp 1626486988
transform 1 0 19087 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_27
timestamp 1626486988
transform 1 0 1624 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_26
timestamp 1626486988
transform 1 0 1604 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_25
timestamp 1626486988
transform 1 0 1610 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_24
timestamp 1626486988
transform 1 0 1725 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_23
timestamp 1626486988
transform 1 0 1615 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_22
timestamp 1626486988
transform 1 0 4120 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_21
timestamp 1626486988
transform 1 0 4100 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_20
timestamp 1626486988
transform 1 0 4106 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_19
timestamp 1626486988
transform 1 0 4221 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_18
timestamp 1626486988
transform 1 0 4111 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_17
timestamp 1626486988
transform 1 0 6616 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_16
timestamp 1626486988
transform 1 0 6596 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_15
timestamp 1626486988
transform 1 0 6602 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_14
timestamp 1626486988
transform 1 0 6717 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_13
timestamp 1626486988
transform 1 0 6607 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_12
timestamp 1626486988
transform 1 0 9112 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_11
timestamp 1626486988
transform 1 0 9092 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_10
timestamp 1626486988
transform 1 0 9098 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_9
timestamp 1626486988
transform 1 0 9213 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_8
timestamp 1626486988
transform 1 0 9103 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_7
timestamp 1626486988
transform 1 0 11608 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_6
timestamp 1626486988
transform 1 0 11588 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_5
timestamp 1626486988
transform 1 0 11594 0 1 575
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_4
timestamp 1626486988
transform 1 0 11709 0 1 778
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_3
timestamp 1626486988
transform 1 0 11599 0 1 1546
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_2
timestamp 1626486988
transform 1 0 14104 0 1 159
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_1
timestamp 1626486988
transform 1 0 14084 0 1 1109
box 0 0 52 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_0
timestamp 1626486988
transform 1 0 14090 0 1 575
box 0 0 52 64
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_31
timestamp 1626486988
transform 1 0 61278 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_30
timestamp 1626486988
transform 1 0 63774 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_29
timestamp 1626486988
transform 1 0 66270 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_28
timestamp 1626486988
transform 1 0 68766 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_27
timestamp 1626486988
transform 1 0 71262 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_26
timestamp 1626486988
transform 1 0 73758 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_25
timestamp 1626486988
transform 1 0 76254 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_24
timestamp 1626486988
transform 1 0 78750 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_23
timestamp 1626486988
transform 1 0 41310 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_22
timestamp 1626486988
transform 1 0 43806 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_21
timestamp 1626486988
transform 1 0 46302 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_20
timestamp 1626486988
transform 1 0 48798 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_19
timestamp 1626486988
transform 1 0 51294 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_18
timestamp 1626486988
transform 1 0 53790 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_17
timestamp 1626486988
transform 1 0 56286 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_16
timestamp 1626486988
transform 1 0 58782 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_15
timestamp 1626486988
transform 1 0 21342 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_14
timestamp 1626486988
transform 1 0 23838 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_13
timestamp 1626486988
transform 1 0 26334 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_12
timestamp 1626486988
transform 1 0 28830 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_11
timestamp 1626486988
transform 1 0 31326 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_10
timestamp 1626486988
transform 1 0 33822 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_9
timestamp 1626486988
transform 1 0 36318 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_8
timestamp 1626486988
transform 1 0 38814 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_7
timestamp 1626486988
transform 1 0 1374 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_6
timestamp 1626486988
transform 1 0 3870 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_5
timestamp 1626486988
transform 1 0 6366 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_4
timestamp 1626486988
transform 1 0 8862 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_3
timestamp 1626486988
transform 1 0 11358 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_2
timestamp 1626486988
transform 1 0 13854 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_1
timestamp 1626486988
transform 1 0 16350 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_0
timestamp 1626486988
transform 1 0 18846 0 1 0
box -376 4 880 2011
<< labels >>
rlabel metal3 s 46509 1092 46607 1190 4 vdd
rlabel metal3 s 49005 1092 49103 1190 4 vdd
rlabel metal3 s 71469 1092 71567 1190 4 vdd
rlabel metal3 s 68973 1092 69071 1190 4 vdd
rlabel metal3 s 53997 1092 54095 1190 4 vdd
rlabel metal3 s 66477 1092 66575 1190 4 vdd
rlabel metal3 s 51501 1092 51599 1190 4 vdd
rlabel metal3 s 73965 1092 74063 1190 4 vdd
rlabel metal3 s 41517 1092 41615 1190 4 vdd
rlabel metal3 s 58989 1092 59087 1190 4 vdd
rlabel metal3 s 61485 1092 61583 1190 4 vdd
rlabel metal3 s 78957 1092 79055 1190 4 vdd
rlabel metal3 s 44013 1092 44111 1190 4 vdd
rlabel metal3 s 56493 1092 56591 1190 4 vdd
rlabel metal3 s 63981 1092 64079 1190 4 vdd
rlabel metal3 s 76461 1092 76559 1190 4 vdd
rlabel metal3 s 49126 760 49224 858 4 gnd
rlabel metal3 s 61606 760 61704 858 4 gnd
rlabel metal3 s 79078 760 79176 858 4 gnd
rlabel metal3 s 59000 1529 59098 1627 4 gnd
rlabel metal3 s 69094 760 69192 858 4 gnd
rlabel metal3 s 41523 558 41621 656 4 gnd
rlabel metal3 s 66483 558 66581 656 4 gnd
rlabel metal3 s 76582 760 76680 858 4 gnd
rlabel metal3 s 63987 558 64085 656 4 gnd
rlabel metal3 s 71590 760 71688 858 4 gnd
rlabel metal3 s 51622 760 51720 858 4 gnd
rlabel metal3 s 51512 1529 51610 1627 4 gnd
rlabel metal3 s 68979 558 69077 656 4 gnd
rlabel metal3 s 54008 1529 54106 1627 4 gnd
rlabel metal3 s 66598 760 66696 858 4 gnd
rlabel metal3 s 76472 1529 76570 1627 4 gnd
rlabel metal3 s 56504 1529 56602 1627 4 gnd
rlabel metal3 s 41528 1529 41626 1627 4 gnd
rlabel metal3 s 54118 760 54216 858 4 gnd
rlabel metal3 s 73976 1529 74074 1627 4 gnd
rlabel metal3 s 49011 558 49109 656 4 gnd
rlabel metal3 s 59110 760 59208 858 4 gnd
rlabel metal3 s 64102 760 64200 858 4 gnd
rlabel metal3 s 74086 760 74184 858 4 gnd
rlabel metal3 s 68984 1529 69082 1627 4 gnd
rlabel metal3 s 58995 558 59093 656 4 gnd
rlabel metal3 s 46515 558 46613 656 4 gnd
rlabel metal3 s 49016 1529 49114 1627 4 gnd
rlabel metal3 s 73971 558 74069 656 4 gnd
rlabel metal3 s 44019 558 44117 656 4 gnd
rlabel metal3 s 71480 1529 71578 1627 4 gnd
rlabel metal3 s 61496 1529 61594 1627 4 gnd
rlabel metal3 s 76467 558 76565 656 4 gnd
rlabel metal3 s 63992 1529 64090 1627 4 gnd
rlabel metal3 s 78968 1529 79066 1627 4 gnd
rlabel metal3 s 44134 760 44232 858 4 gnd
rlabel metal3 s 78963 558 79061 656 4 gnd
rlabel metal3 s 46630 760 46728 858 4 gnd
rlabel metal3 s 46520 1529 46618 1627 4 gnd
rlabel metal3 s 66488 1529 66586 1627 4 gnd
rlabel metal3 s 61491 558 61589 656 4 gnd
rlabel metal3 s 56614 760 56712 858 4 gnd
rlabel metal3 s 54003 558 54101 656 4 gnd
rlabel metal3 s 56499 558 56597 656 4 gnd
rlabel metal3 s 41638 760 41736 858 4 gnd
rlabel metal3 s 44024 1529 44122 1627 4 gnd
rlabel metal3 s 51507 558 51605 656 4 gnd
rlabel metal3 s 71475 558 71573 656 4 gnd
rlabel metal3 s 34040 1529 34138 1627 4 gnd
rlabel metal3 s 1581 1092 1679 1190 4 vdd
rlabel metal3 s 16557 1092 16655 1190 4 vdd
rlabel metal3 s 16563 558 16661 656 4 gnd
rlabel metal3 s 31654 760 31752 858 4 gnd
rlabel metal3 s 29158 760 29256 858 4 gnd
rlabel metal3 s 4088 1529 4186 1627 4 gnd
rlabel metal3 s 14182 760 14280 858 4 gnd
rlabel metal3 s 6579 558 6677 656 4 gnd
rlabel metal3 s 11565 1092 11663 1190 4 vdd
rlabel metal3 s 14061 1092 14159 1190 4 vdd
rlabel metal3 s 6573 1092 6671 1190 4 vdd
rlabel metal3 s 26552 1529 26650 1627 4 gnd
rlabel metal3 s 1592 1529 1690 1627 4 gnd
rlabel metal3 s 16568 1529 16666 1627 4 gnd
rlabel metal3 s 11576 1529 11674 1627 4 gnd
rlabel metal3 s 36531 558 36629 656 4 gnd
rlabel metal3 s 36525 1092 36623 1190 4 vdd
rlabel metal3 s 9080 1529 9178 1627 4 gnd
rlabel metal3 s 16678 760 16776 858 4 gnd
rlabel metal3 s 39027 558 39125 656 4 gnd
rlabel metal3 s 24166 760 24264 858 4 gnd
rlabel metal3 s 21670 760 21768 858 4 gnd
rlabel metal3 s 29037 1092 29135 1190 4 vdd
rlabel metal3 s 4077 1092 4175 1190 4 vdd
rlabel metal3 s 9075 558 9173 656 4 gnd
rlabel metal3 s 24045 1092 24143 1190 4 vdd
rlabel metal3 s 14072 1529 14170 1627 4 gnd
rlabel metal3 s 4198 760 4296 858 4 gnd
rlabel metal3 s 39021 1092 39119 1190 4 vdd
rlabel metal3 s 21560 1529 21658 1627 4 gnd
rlabel metal3 s 31544 1529 31642 1627 4 gnd
rlabel metal3 s 19053 1092 19151 1190 4 vdd
rlabel metal3 s 39142 760 39240 858 4 gnd
rlabel metal3 s 21549 1092 21647 1190 4 vdd
rlabel metal3 s 34035 558 34133 656 4 gnd
rlabel metal3 s 11571 558 11669 656 4 gnd
rlabel metal3 s 31539 558 31637 656 4 gnd
rlabel metal3 s 31533 1092 31631 1190 4 vdd
rlabel metal3 s 26541 1092 26639 1190 4 vdd
rlabel metal3 s 24051 558 24149 656 4 gnd
rlabel metal3 s 36646 760 36744 858 4 gnd
rlabel metal3 s 11686 760 11784 858 4 gnd
rlabel metal3 s 4083 558 4181 656 4 gnd
rlabel metal3 s 19174 760 19272 858 4 gnd
rlabel metal3 s 9069 1092 9167 1190 4 vdd
rlabel metal3 s 9190 760 9288 858 4 gnd
rlabel metal3 s 21555 558 21653 656 4 gnd
rlabel metal3 s 6694 760 6792 858 4 gnd
rlabel metal3 s 19059 558 19157 656 4 gnd
rlabel metal3 s 6584 1529 6682 1627 4 gnd
rlabel metal3 s 1587 558 1685 656 4 gnd
rlabel metal3 s 26662 760 26760 858 4 gnd
rlabel metal3 s 14067 558 14165 656 4 gnd
rlabel metal3 s 1702 760 1800 858 4 gnd
rlabel metal3 s 36536 1529 36634 1627 4 gnd
rlabel metal3 s 29048 1529 29146 1627 4 gnd
rlabel metal3 s 34150 760 34248 858 4 gnd
rlabel metal3 s 24056 1529 24154 1627 4 gnd
rlabel metal3 s 29043 558 29141 656 4 gnd
rlabel metal3 s 34029 1092 34127 1190 4 vdd
rlabel metal3 s 26547 558 26645 656 4 gnd
rlabel metal3 s 39032 1529 39130 1627 4 gnd
rlabel metal3 s 19064 1529 19162 1627 4 gnd
rlabel metal3 s 34049 142 34147 240 4 vdd
rlabel metal3 s 16577 142 16675 240 4 vdd
rlabel metal3 s 14081 142 14179 240 4 vdd
rlabel metal3 s 1601 142 1699 240 4 vdd
rlabel metal3 s 39041 142 39139 240 4 vdd
rlabel metal3 s 21569 142 21667 240 4 vdd
rlabel metal3 s 36545 142 36643 240 4 vdd
rlabel metal3 s 26561 142 26659 240 4 vdd
rlabel metal3 s 9089 142 9187 240 4 vdd
rlabel metal3 s 19073 142 19171 240 4 vdd
rlabel metal3 s 31553 142 31651 240 4 vdd
rlabel metal3 s 29057 142 29155 240 4 vdd
rlabel metal3 s 11585 142 11683 240 4 vdd
rlabel metal3 s 4097 142 4195 240 4 vdd
rlabel metal3 s 24065 142 24163 240 4 vdd
rlabel metal3 s 6593 142 6691 240 4 vdd
rlabel metal3 s 46529 142 46627 240 4 vdd
rlabel metal3 s 71489 142 71587 240 4 vdd
rlabel metal3 s 41537 142 41635 240 4 vdd
rlabel metal3 s 76481 142 76579 240 4 vdd
rlabel metal3 s 68993 142 69091 240 4 vdd
rlabel metal3 s 73985 142 74083 240 4 vdd
rlabel metal3 s 61505 142 61603 240 4 vdd
rlabel metal3 s 56513 142 56611 240 4 vdd
rlabel metal3 s 66497 142 66595 240 4 vdd
rlabel metal3 s 51521 142 51619 240 4 vdd
rlabel metal3 s 64001 142 64099 240 4 vdd
rlabel metal3 s 49025 142 49123 240 4 vdd
rlabel metal3 s 78977 142 79075 240 4 vdd
rlabel metal3 s 44033 142 44131 240 4 vdd
rlabel metal3 s 54017 142 54115 240 4 vdd
rlabel metal3 s 59009 142 59107 240 4 vdd
rlabel metal1 s 1629 4 1689 60 4 data_0
rlabel metal1 s 1500 1959 1530 2011 4 bl_0
rlabel metal1 s 1702 1959 1732 2011 4 br_0
rlabel metal1 s 4125 4 4185 60 4 data_1
rlabel metal1 s 3996 1959 4026 2011 4 bl_1
rlabel metal1 s 4198 1959 4228 2011 4 br_1
rlabel metal1 s 6621 4 6681 60 4 data_2
rlabel metal1 s 6492 1959 6522 2011 4 bl_2
rlabel metal1 s 6694 1959 6724 2011 4 br_2
rlabel metal1 s 9117 4 9177 60 4 data_3
rlabel metal1 s 8988 1959 9018 2011 4 bl_3
rlabel metal1 s 9190 1959 9220 2011 4 br_3
rlabel metal1 s 11613 4 11673 60 4 data_4
rlabel metal1 s 11484 1959 11514 2011 4 bl_4
rlabel metal1 s 11686 1959 11716 2011 4 br_4
rlabel metal1 s 14109 4 14169 60 4 data_5
rlabel metal1 s 13980 1959 14010 2011 4 bl_5
rlabel metal1 s 14182 1959 14212 2011 4 br_5
rlabel metal1 s 16605 4 16665 60 4 data_6
rlabel metal1 s 16476 1959 16506 2011 4 bl_6
rlabel metal1 s 16678 1959 16708 2011 4 br_6
rlabel metal1 s 19101 4 19161 60 4 data_7
rlabel metal1 s 18972 1959 19002 2011 4 bl_7
rlabel metal1 s 19174 1959 19204 2011 4 br_7
rlabel metal1 s 21597 4 21657 60 4 data_8
rlabel metal1 s 21468 1959 21498 2011 4 bl_8
rlabel metal1 s 21670 1959 21700 2011 4 br_8
rlabel metal1 s 24093 4 24153 60 4 data_9
rlabel metal1 s 23964 1959 23994 2011 4 bl_9
rlabel metal1 s 24166 1959 24196 2011 4 br_9
rlabel metal1 s 26589 4 26649 60 4 data_10
rlabel metal1 s 26460 1959 26490 2011 4 bl_10
rlabel metal1 s 26662 1959 26692 2011 4 br_10
rlabel metal1 s 29085 4 29145 60 4 data_11
rlabel metal1 s 28956 1959 28986 2011 4 bl_11
rlabel metal1 s 29158 1959 29188 2011 4 br_11
rlabel metal1 s 31581 4 31641 60 4 data_12
rlabel metal1 s 31452 1959 31482 2011 4 bl_12
rlabel metal1 s 31654 1959 31684 2011 4 br_12
rlabel metal1 s 34077 4 34137 60 4 data_13
rlabel metal1 s 33948 1959 33978 2011 4 bl_13
rlabel metal1 s 34150 1959 34180 2011 4 br_13
rlabel metal1 s 36573 4 36633 60 4 data_14
rlabel metal1 s 36444 1959 36474 2011 4 bl_14
rlabel metal1 s 36646 1959 36676 2011 4 br_14
rlabel metal1 s 39069 4 39129 60 4 data_15
rlabel metal1 s 38940 1959 38970 2011 4 bl_15
rlabel metal1 s 39142 1959 39172 2011 4 br_15
rlabel metal1 s 41565 4 41625 60 4 data_16
rlabel metal1 s 41436 1959 41466 2011 4 bl_16
rlabel metal1 s 41638 1959 41668 2011 4 br_16
rlabel metal1 s 44061 4 44121 60 4 data_17
rlabel metal1 s 43932 1959 43962 2011 4 bl_17
rlabel metal1 s 44134 1959 44164 2011 4 br_17
rlabel metal1 s 46557 4 46617 60 4 data_18
rlabel metal1 s 46428 1959 46458 2011 4 bl_18
rlabel metal1 s 46630 1959 46660 2011 4 br_18
rlabel metal1 s 49053 4 49113 60 4 data_19
rlabel metal1 s 48924 1959 48954 2011 4 bl_19
rlabel metal1 s 49126 1959 49156 2011 4 br_19
rlabel metal1 s 51549 4 51609 60 4 data_20
rlabel metal1 s 51420 1959 51450 2011 4 bl_20
rlabel metal1 s 51622 1959 51652 2011 4 br_20
rlabel metal1 s 54045 4 54105 60 4 data_21
rlabel metal1 s 53916 1959 53946 2011 4 bl_21
rlabel metal1 s 54118 1959 54148 2011 4 br_21
rlabel metal1 s 56541 4 56601 60 4 data_22
rlabel metal1 s 56412 1959 56442 2011 4 bl_22
rlabel metal1 s 56614 1959 56644 2011 4 br_22
rlabel metal1 s 59037 4 59097 60 4 data_23
rlabel metal1 s 58908 1959 58938 2011 4 bl_23
rlabel metal1 s 59110 1959 59140 2011 4 br_23
rlabel metal1 s 61533 4 61593 60 4 data_24
rlabel metal1 s 61404 1959 61434 2011 4 bl_24
rlabel metal1 s 61606 1959 61636 2011 4 br_24
rlabel metal1 s 64029 4 64089 60 4 data_25
rlabel metal1 s 63900 1959 63930 2011 4 bl_25
rlabel metal1 s 64102 1959 64132 2011 4 br_25
rlabel metal1 s 66525 4 66585 60 4 data_26
rlabel metal1 s 66396 1959 66426 2011 4 bl_26
rlabel metal1 s 66598 1959 66628 2011 4 br_26
rlabel metal1 s 69021 4 69081 60 4 data_27
rlabel metal1 s 68892 1959 68922 2011 4 bl_27
rlabel metal1 s 69094 1959 69124 2011 4 br_27
rlabel metal1 s 71517 4 71577 60 4 data_28
rlabel metal1 s 71388 1959 71418 2011 4 bl_28
rlabel metal1 s 71590 1959 71620 2011 4 br_28
rlabel metal1 s 74013 4 74073 60 4 data_29
rlabel metal1 s 73884 1959 73914 2011 4 bl_29
rlabel metal1 s 74086 1959 74116 2011 4 br_29
rlabel metal1 s 76509 4 76569 60 4 data_30
rlabel metal1 s 76380 1959 76410 2011 4 bl_30
rlabel metal1 s 76582 1959 76612 2011 4 br_30
rlabel metal1 s 79005 4 79065 60 4 data_31
rlabel metal1 s 78876 1959 78906 2011 4 bl_31
rlabel metal1 s 79078 1959 79108 2011 4 br_31
rlabel metal1 s 1473 94 20817 128 4 en_0
rlabel metal1 s 21441 94 40785 128 4 en_1
rlabel metal1 s 41409 94 60753 128 4 en_2
rlabel metal1 s 61377 94 80721 128 4 en_3
<< properties >>
string FIXED_BBOX 0 0 79250 2011
<< end >>
