magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_s >>
rect 1422 679 1458 1471
<< locali >>
rect 0 1396 2518 1432
rect 0 -18 2518 18
<< metal1 >>
rect -32 1388 32 1440
rect -32 -26 32 26
<< metal2 >>
rect -28 1390 28 1438
rect 137 538 203 590
rect -28 -24 28 24
rect 369 0 397 1414
rect 1822 871 1850 899
rect 2328 489 2356 517
<< metal3 >>
rect -49 1365 49 1463
rect -49 -49 49 49
use dff_buf_0  dff_buf_0_0
timestamp 1624494425
transform 1 0 0 0 1 0
box -36 -43 2554 1471
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 -33 0 1 -37
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 -32 0 1 -32
box 0 0 64 64
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 -29 0 1 -33
box 0 0 58 66
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 -33 0 1 1377
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 -32 0 1 1382
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 -29 0 1 1381
box 0 0 58 66
<< labels >>
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal2 s 137 538 203 590 4 din_0
rlabel metal2 s 2328 489 2356 517 4 dout_0
rlabel metal2 s 1822 871 1850 899 4 dout_bar_0
rlabel metal2 s 369 0 397 1414 4 clk
<< properties >>
string FIXED_BBOX 0 0 2518 1414
<< end >>
