magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1309 -1260 83929 53400
<< metal1 >>
rect 972 0 1008 52140
rect 1044 0 1080 52140
rect 1116 51429 1152 51770
rect 1116 50639 1152 51271
rect 1116 49849 1152 50481
rect 1116 49059 1152 49691
rect 1116 48269 1152 48901
rect 1116 47479 1152 48111
rect 1116 46689 1152 47321
rect 1116 45899 1152 46531
rect 1116 45109 1152 45741
rect 1116 44319 1152 44951
rect 1116 43529 1152 44161
rect 1116 42739 1152 43371
rect 1116 41949 1152 42581
rect 1116 41159 1152 41791
rect 1116 40369 1152 41001
rect 1116 39579 1152 40211
rect 1116 38789 1152 39421
rect 1116 37999 1152 38631
rect 1116 37209 1152 37841
rect 1116 36419 1152 37051
rect 1116 35629 1152 36261
rect 1116 34839 1152 35471
rect 1116 34049 1152 34681
rect 1116 33259 1152 33891
rect 1116 32469 1152 33101
rect 1116 31679 1152 32311
rect 1116 30889 1152 31521
rect 1116 30099 1152 30731
rect 1116 29309 1152 29941
rect 1116 28519 1152 29151
rect 1116 27729 1152 28361
rect 1116 26939 1152 27571
rect 1116 26149 1152 26781
rect 1116 25359 1152 25991
rect 1116 24569 1152 25201
rect 1116 23779 1152 24411
rect 1116 22989 1152 23621
rect 1116 22199 1152 22831
rect 1116 21409 1152 22041
rect 1116 20619 1152 21251
rect 1116 19829 1152 20461
rect 1116 19039 1152 19671
rect 1116 18249 1152 18881
rect 1116 17459 1152 18091
rect 1116 16669 1152 17301
rect 1116 15879 1152 16511
rect 1116 15089 1152 15721
rect 1116 14299 1152 14931
rect 1116 13509 1152 14141
rect 1116 12719 1152 13351
rect 1116 11929 1152 12561
rect 1116 11139 1152 11771
rect 1116 10349 1152 10981
rect 1116 9559 1152 10191
rect 1116 8769 1152 9401
rect 1116 7979 1152 8611
rect 1116 7189 1152 7821
rect 1116 6399 1152 7031
rect 1116 5609 1152 6241
rect 1116 4819 1152 5451
rect 1116 4029 1152 4661
rect 1116 3239 1152 3871
rect 1116 2449 1152 3081
rect 1116 1659 1152 2291
rect 1116 869 1152 1501
rect 1116 370 1152 711
rect 1188 0 1224 52140
rect 1260 0 1296 52140
rect 1452 0 1488 52140
rect 1524 0 1560 52140
rect 1668 0 1704 52140
rect 1740 0 1776 52140
rect 2220 0 2256 52140
rect 2292 0 2328 52140
rect 2436 0 2472 52140
rect 2508 0 2544 52140
rect 2700 0 2736 52140
rect 2772 0 2808 52140
rect 2916 0 2952 52140
rect 2988 0 3024 52140
rect 3468 0 3504 52140
rect 3540 0 3576 52140
rect 3684 0 3720 52140
rect 3756 0 3792 52140
rect 3948 0 3984 52140
rect 4020 0 4056 52140
rect 4164 0 4200 52140
rect 4236 0 4272 52140
rect 4716 0 4752 52140
rect 4788 0 4824 52140
rect 4932 0 4968 52140
rect 5004 0 5040 52140
rect 5196 0 5232 52140
rect 5268 0 5304 52140
rect 5412 0 5448 52140
rect 5484 0 5520 52140
rect 5964 0 6000 52140
rect 6036 0 6072 52140
rect 6180 0 6216 52140
rect 6252 0 6288 52140
rect 6444 0 6480 52140
rect 6516 0 6552 52140
rect 6660 0 6696 52140
rect 6732 0 6768 52140
rect 7212 0 7248 52140
rect 7284 0 7320 52140
rect 7428 0 7464 52140
rect 7500 0 7536 52140
rect 7692 0 7728 52140
rect 7764 0 7800 52140
rect 7908 0 7944 52140
rect 7980 0 8016 52140
rect 8460 0 8496 52140
rect 8532 0 8568 52140
rect 8676 0 8712 52140
rect 8748 0 8784 52140
rect 8940 0 8976 52140
rect 9012 0 9048 52140
rect 9156 0 9192 52140
rect 9228 0 9264 52140
rect 9708 0 9744 52140
rect 9780 0 9816 52140
rect 9924 0 9960 52140
rect 9996 0 10032 52140
rect 10188 0 10224 52140
rect 10260 0 10296 52140
rect 10404 0 10440 52140
rect 10476 0 10512 52140
rect 10956 0 10992 52140
rect 11028 0 11064 52140
rect 11172 0 11208 52140
rect 11244 0 11280 52140
rect 11436 0 11472 52140
rect 11508 0 11544 52140
rect 11652 0 11688 52140
rect 11724 0 11760 52140
rect 12204 0 12240 52140
rect 12276 0 12312 52140
rect 12420 0 12456 52140
rect 12492 0 12528 52140
rect 12684 0 12720 52140
rect 12756 0 12792 52140
rect 12900 0 12936 52140
rect 12972 0 13008 52140
rect 13452 0 13488 52140
rect 13524 0 13560 52140
rect 13668 0 13704 52140
rect 13740 0 13776 52140
rect 13932 0 13968 52140
rect 14004 0 14040 52140
rect 14148 0 14184 52140
rect 14220 0 14256 52140
rect 14700 0 14736 52140
rect 14772 0 14808 52140
rect 14916 0 14952 52140
rect 14988 0 15024 52140
rect 15180 0 15216 52140
rect 15252 0 15288 52140
rect 15396 0 15432 52140
rect 15468 0 15504 52140
rect 15948 0 15984 52140
rect 16020 0 16056 52140
rect 16164 0 16200 52140
rect 16236 0 16272 52140
rect 16428 0 16464 52140
rect 16500 0 16536 52140
rect 16644 0 16680 52140
rect 16716 0 16752 52140
rect 17196 0 17232 52140
rect 17268 0 17304 52140
rect 17412 0 17448 52140
rect 17484 0 17520 52140
rect 17676 0 17712 52140
rect 17748 0 17784 52140
rect 17892 0 17928 52140
rect 17964 0 18000 52140
rect 18444 0 18480 52140
rect 18516 0 18552 52140
rect 18660 0 18696 52140
rect 18732 0 18768 52140
rect 18924 0 18960 52140
rect 18996 0 19032 52140
rect 19140 0 19176 52140
rect 19212 0 19248 52140
rect 19692 0 19728 52140
rect 19764 0 19800 52140
rect 19908 0 19944 52140
rect 19980 0 20016 52140
rect 20172 0 20208 52140
rect 20244 0 20280 52140
rect 20388 0 20424 52140
rect 20460 0 20496 52140
rect 20940 0 20976 52140
rect 21012 0 21048 52140
rect 21156 0 21192 52140
rect 21228 0 21264 52140
rect 21420 0 21456 52140
rect 21492 0 21528 52140
rect 21636 0 21672 52140
rect 21708 0 21744 52140
rect 22188 0 22224 52140
rect 22260 0 22296 52140
rect 22404 0 22440 52140
rect 22476 0 22512 52140
rect 22668 0 22704 52140
rect 22740 0 22776 52140
rect 22884 0 22920 52140
rect 22956 0 22992 52140
rect 23436 0 23472 52140
rect 23508 0 23544 52140
rect 23652 0 23688 52140
rect 23724 0 23760 52140
rect 23916 0 23952 52140
rect 23988 0 24024 52140
rect 24132 0 24168 52140
rect 24204 0 24240 52140
rect 24684 0 24720 52140
rect 24756 0 24792 52140
rect 24900 0 24936 52140
rect 24972 0 25008 52140
rect 25164 0 25200 52140
rect 25236 0 25272 52140
rect 25380 0 25416 52140
rect 25452 0 25488 52140
rect 25932 0 25968 52140
rect 26004 0 26040 52140
rect 26148 0 26184 52140
rect 26220 0 26256 52140
rect 26412 0 26448 52140
rect 26484 0 26520 52140
rect 26628 0 26664 52140
rect 26700 0 26736 52140
rect 27180 0 27216 52140
rect 27252 0 27288 52140
rect 27396 0 27432 52140
rect 27468 0 27504 52140
rect 27660 0 27696 52140
rect 27732 0 27768 52140
rect 27876 0 27912 52140
rect 27948 0 27984 52140
rect 28428 0 28464 52140
rect 28500 0 28536 52140
rect 28644 0 28680 52140
rect 28716 0 28752 52140
rect 28908 0 28944 52140
rect 28980 0 29016 52140
rect 29124 0 29160 52140
rect 29196 0 29232 52140
rect 29676 0 29712 52140
rect 29748 0 29784 52140
rect 29892 0 29928 52140
rect 29964 0 30000 52140
rect 30156 0 30192 52140
rect 30228 0 30264 52140
rect 30372 0 30408 52140
rect 30444 0 30480 52140
rect 30924 0 30960 52140
rect 30996 0 31032 52140
rect 31140 0 31176 52140
rect 31212 0 31248 52140
rect 31404 0 31440 52140
rect 31476 0 31512 52140
rect 31620 0 31656 52140
rect 31692 0 31728 52140
rect 32172 0 32208 52140
rect 32244 0 32280 52140
rect 32388 0 32424 52140
rect 32460 0 32496 52140
rect 32652 0 32688 52140
rect 32724 0 32760 52140
rect 32868 0 32904 52140
rect 32940 0 32976 52140
rect 33420 0 33456 52140
rect 33492 0 33528 52140
rect 33636 0 33672 52140
rect 33708 0 33744 52140
rect 33900 0 33936 52140
rect 33972 0 34008 52140
rect 34116 0 34152 52140
rect 34188 0 34224 52140
rect 34668 0 34704 52140
rect 34740 0 34776 52140
rect 34884 0 34920 52140
rect 34956 0 34992 52140
rect 35148 0 35184 52140
rect 35220 0 35256 52140
rect 35364 0 35400 52140
rect 35436 0 35472 52140
rect 35916 0 35952 52140
rect 35988 0 36024 52140
rect 36132 0 36168 52140
rect 36204 0 36240 52140
rect 36396 0 36432 52140
rect 36468 0 36504 52140
rect 36612 0 36648 52140
rect 36684 0 36720 52140
rect 37164 0 37200 52140
rect 37236 0 37272 52140
rect 37380 0 37416 52140
rect 37452 0 37488 52140
rect 37644 0 37680 52140
rect 37716 0 37752 52140
rect 37860 0 37896 52140
rect 37932 0 37968 52140
rect 38412 0 38448 52140
rect 38484 0 38520 52140
rect 38628 0 38664 52140
rect 38700 0 38736 52140
rect 38892 0 38928 52140
rect 38964 0 39000 52140
rect 39108 0 39144 52140
rect 39180 0 39216 52140
rect 39660 0 39696 52140
rect 39732 0 39768 52140
rect 39876 0 39912 52140
rect 39948 0 39984 52140
rect 40140 0 40176 52140
rect 40212 0 40248 52140
rect 40356 0 40392 52140
rect 40428 0 40464 52140
rect 40908 0 40944 52140
rect 40980 0 41016 52140
rect 41124 0 41160 52140
rect 41196 0 41232 52140
rect 41388 0 41424 52140
rect 41460 0 41496 52140
rect 41604 0 41640 52140
rect 41676 0 41712 52140
rect 42156 0 42192 52140
rect 42228 0 42264 52140
rect 42372 0 42408 52140
rect 42444 0 42480 52140
rect 42636 0 42672 52140
rect 42708 0 42744 52140
rect 42852 0 42888 52140
rect 42924 0 42960 52140
rect 43404 0 43440 52140
rect 43476 0 43512 52140
rect 43620 0 43656 52140
rect 43692 0 43728 52140
rect 43884 0 43920 52140
rect 43956 0 43992 52140
rect 44100 0 44136 52140
rect 44172 0 44208 52140
rect 44652 0 44688 52140
rect 44724 0 44760 52140
rect 44868 0 44904 52140
rect 44940 0 44976 52140
rect 45132 0 45168 52140
rect 45204 0 45240 52140
rect 45348 0 45384 52140
rect 45420 0 45456 52140
rect 45900 0 45936 52140
rect 45972 0 46008 52140
rect 46116 0 46152 52140
rect 46188 0 46224 52140
rect 46380 0 46416 52140
rect 46452 0 46488 52140
rect 46596 0 46632 52140
rect 46668 0 46704 52140
rect 47148 0 47184 52140
rect 47220 0 47256 52140
rect 47364 0 47400 52140
rect 47436 0 47472 52140
rect 47628 0 47664 52140
rect 47700 0 47736 52140
rect 47844 0 47880 52140
rect 47916 0 47952 52140
rect 48396 0 48432 52140
rect 48468 0 48504 52140
rect 48612 0 48648 52140
rect 48684 0 48720 52140
rect 48876 0 48912 52140
rect 48948 0 48984 52140
rect 49092 0 49128 52140
rect 49164 0 49200 52140
rect 49644 0 49680 52140
rect 49716 0 49752 52140
rect 49860 0 49896 52140
rect 49932 0 49968 52140
rect 50124 0 50160 52140
rect 50196 0 50232 52140
rect 50340 0 50376 52140
rect 50412 0 50448 52140
rect 50892 0 50928 52140
rect 50964 0 51000 52140
rect 51108 0 51144 52140
rect 51180 0 51216 52140
rect 51372 0 51408 52140
rect 51444 0 51480 52140
rect 51588 0 51624 52140
rect 51660 0 51696 52140
rect 52140 0 52176 52140
rect 52212 0 52248 52140
rect 52356 0 52392 52140
rect 52428 0 52464 52140
rect 52620 0 52656 52140
rect 52692 0 52728 52140
rect 52836 0 52872 52140
rect 52908 0 52944 52140
rect 53388 0 53424 52140
rect 53460 0 53496 52140
rect 53604 0 53640 52140
rect 53676 0 53712 52140
rect 53868 0 53904 52140
rect 53940 0 53976 52140
rect 54084 0 54120 52140
rect 54156 0 54192 52140
rect 54636 0 54672 52140
rect 54708 0 54744 52140
rect 54852 0 54888 52140
rect 54924 0 54960 52140
rect 55116 0 55152 52140
rect 55188 0 55224 52140
rect 55332 0 55368 52140
rect 55404 0 55440 52140
rect 55884 0 55920 52140
rect 55956 0 55992 52140
rect 56100 0 56136 52140
rect 56172 0 56208 52140
rect 56364 0 56400 52140
rect 56436 0 56472 52140
rect 56580 0 56616 52140
rect 56652 0 56688 52140
rect 57132 0 57168 52140
rect 57204 0 57240 52140
rect 57348 0 57384 52140
rect 57420 0 57456 52140
rect 57612 0 57648 52140
rect 57684 0 57720 52140
rect 57828 0 57864 52140
rect 57900 0 57936 52140
rect 58380 0 58416 52140
rect 58452 0 58488 52140
rect 58596 0 58632 52140
rect 58668 0 58704 52140
rect 58860 0 58896 52140
rect 58932 0 58968 52140
rect 59076 0 59112 52140
rect 59148 0 59184 52140
rect 59628 0 59664 52140
rect 59700 0 59736 52140
rect 59844 0 59880 52140
rect 59916 0 59952 52140
rect 60108 0 60144 52140
rect 60180 0 60216 52140
rect 60324 0 60360 52140
rect 60396 0 60432 52140
rect 60876 0 60912 52140
rect 60948 0 60984 52140
rect 61092 0 61128 52140
rect 61164 0 61200 52140
rect 61356 0 61392 52140
rect 61428 0 61464 52140
rect 61572 0 61608 52140
rect 61644 0 61680 52140
rect 62124 0 62160 52140
rect 62196 0 62232 52140
rect 62340 0 62376 52140
rect 62412 0 62448 52140
rect 62604 0 62640 52140
rect 62676 0 62712 52140
rect 62820 0 62856 52140
rect 62892 0 62928 52140
rect 63372 0 63408 52140
rect 63444 0 63480 52140
rect 63588 0 63624 52140
rect 63660 0 63696 52140
rect 63852 0 63888 52140
rect 63924 0 63960 52140
rect 64068 0 64104 52140
rect 64140 0 64176 52140
rect 64620 0 64656 52140
rect 64692 0 64728 52140
rect 64836 0 64872 52140
rect 64908 0 64944 52140
rect 65100 0 65136 52140
rect 65172 0 65208 52140
rect 65316 0 65352 52140
rect 65388 0 65424 52140
rect 65868 0 65904 52140
rect 65940 0 65976 52140
rect 66084 0 66120 52140
rect 66156 0 66192 52140
rect 66348 0 66384 52140
rect 66420 0 66456 52140
rect 66564 0 66600 52140
rect 66636 0 66672 52140
rect 67116 0 67152 52140
rect 67188 0 67224 52140
rect 67332 0 67368 52140
rect 67404 0 67440 52140
rect 67596 0 67632 52140
rect 67668 0 67704 52140
rect 67812 0 67848 52140
rect 67884 0 67920 52140
rect 68364 0 68400 52140
rect 68436 0 68472 52140
rect 68580 0 68616 52140
rect 68652 0 68688 52140
rect 68844 0 68880 52140
rect 68916 0 68952 52140
rect 69060 0 69096 52140
rect 69132 0 69168 52140
rect 69612 0 69648 52140
rect 69684 0 69720 52140
rect 69828 0 69864 52140
rect 69900 0 69936 52140
rect 70092 0 70128 52140
rect 70164 0 70200 52140
rect 70308 0 70344 52140
rect 70380 0 70416 52140
rect 70860 0 70896 52140
rect 70932 0 70968 52140
rect 71076 0 71112 52140
rect 71148 0 71184 52140
rect 71340 0 71376 52140
rect 71412 0 71448 52140
rect 71556 0 71592 52140
rect 71628 0 71664 52140
rect 72108 0 72144 52140
rect 72180 0 72216 52140
rect 72324 0 72360 52140
rect 72396 0 72432 52140
rect 72588 0 72624 52140
rect 72660 0 72696 52140
rect 72804 0 72840 52140
rect 72876 0 72912 52140
rect 73356 0 73392 52140
rect 73428 0 73464 52140
rect 73572 0 73608 52140
rect 73644 0 73680 52140
rect 73836 0 73872 52140
rect 73908 0 73944 52140
rect 74052 0 74088 52140
rect 74124 0 74160 52140
rect 74604 0 74640 52140
rect 74676 0 74712 52140
rect 74820 0 74856 52140
rect 74892 0 74928 52140
rect 75084 0 75120 52140
rect 75156 0 75192 52140
rect 75300 0 75336 52140
rect 75372 0 75408 52140
rect 75852 0 75888 52140
rect 75924 0 75960 52140
rect 76068 0 76104 52140
rect 76140 0 76176 52140
rect 76332 0 76368 52140
rect 76404 0 76440 52140
rect 76548 0 76584 52140
rect 76620 0 76656 52140
rect 77100 0 77136 52140
rect 77172 0 77208 52140
rect 77316 0 77352 52140
rect 77388 0 77424 52140
rect 77580 0 77616 52140
rect 77652 0 77688 52140
rect 77796 0 77832 52140
rect 77868 0 77904 52140
rect 78348 0 78384 52140
rect 78420 0 78456 52140
rect 78564 0 78600 52140
rect 78636 0 78672 52140
rect 78828 0 78864 52140
rect 78900 0 78936 52140
rect 79044 0 79080 52140
rect 79116 0 79152 52140
rect 79596 0 79632 52140
rect 79668 0 79704 52140
rect 79812 0 79848 52140
rect 79884 0 79920 52140
rect 80076 0 80112 52140
rect 80148 0 80184 52140
rect 80292 0 80328 52140
rect 80364 0 80400 52140
rect 80844 0 80880 52140
rect 80916 0 80952 52140
rect 81060 0 81096 52140
rect 81132 0 81168 52140
rect 81324 0 81360 52140
rect 81396 0 81432 52140
rect 81468 51429 81504 51770
rect 81468 50639 81504 51271
rect 81468 49849 81504 50481
rect 81468 49059 81504 49691
rect 81468 48269 81504 48901
rect 81468 47479 81504 48111
rect 81468 46689 81504 47321
rect 81468 45899 81504 46531
rect 81468 45109 81504 45741
rect 81468 44319 81504 44951
rect 81468 43529 81504 44161
rect 81468 42739 81504 43371
rect 81468 41949 81504 42581
rect 81468 41159 81504 41791
rect 81468 40369 81504 41001
rect 81468 39579 81504 40211
rect 81468 38789 81504 39421
rect 81468 37999 81504 38631
rect 81468 37209 81504 37841
rect 81468 36419 81504 37051
rect 81468 35629 81504 36261
rect 81468 34839 81504 35471
rect 81468 34049 81504 34681
rect 81468 33259 81504 33891
rect 81468 32469 81504 33101
rect 81468 31679 81504 32311
rect 81468 30889 81504 31521
rect 81468 30099 81504 30731
rect 81468 29309 81504 29941
rect 81468 28519 81504 29151
rect 81468 27729 81504 28361
rect 81468 26939 81504 27571
rect 81468 26149 81504 26781
rect 81468 25359 81504 25991
rect 81468 24569 81504 25201
rect 81468 23779 81504 24411
rect 81468 22989 81504 23621
rect 81468 22199 81504 22831
rect 81468 21409 81504 22041
rect 81468 20619 81504 21251
rect 81468 19829 81504 20461
rect 81468 19039 81504 19671
rect 81468 18249 81504 18881
rect 81468 17459 81504 18091
rect 81468 16669 81504 17301
rect 81468 15879 81504 16511
rect 81468 15089 81504 15721
rect 81468 14299 81504 14931
rect 81468 13509 81504 14141
rect 81468 12719 81504 13351
rect 81468 11929 81504 12561
rect 81468 11139 81504 11771
rect 81468 10349 81504 10981
rect 81468 9559 81504 10191
rect 81468 8769 81504 9401
rect 81468 7979 81504 8611
rect 81468 7189 81504 7821
rect 81468 6399 81504 7031
rect 81468 5609 81504 6241
rect 81468 4819 81504 5451
rect 81468 4029 81504 4661
rect 81468 3239 81504 3871
rect 81468 2449 81504 3081
rect 81468 1659 81504 2291
rect 81468 869 81504 1501
rect 81468 370 81504 711
rect 81540 0 81576 52140
rect 81612 0 81648 52140
<< metal2 >>
rect 0 51716 82620 51721
rect -37 51679 82657 51716
rect 0 51673 82620 51679
rect 1080 51549 1188 51625
rect 81432 51549 81540 51625
rect 0 51453 82620 51501
rect 1080 51295 1188 51405
rect 81432 51295 81540 51405
rect 0 51199 82620 51247
rect 1080 51075 1188 51151
rect 81432 51075 81540 51151
rect 0 50979 82620 51027
rect 0 50883 82620 50931
rect 1080 50759 1188 50835
rect 81432 50759 81540 50835
rect 0 50663 82620 50711
rect 1080 50505 1188 50615
rect 81432 50505 81540 50615
rect 0 50409 82620 50457
rect 1080 50285 1188 50361
rect 81432 50285 81540 50361
rect 0 50189 82620 50237
rect 0 50093 82620 50141
rect 1080 49969 1188 50045
rect 81432 49969 81540 50045
rect 0 49873 82620 49921
rect 1080 49715 1188 49825
rect 81432 49715 81540 49825
rect 0 49619 82620 49667
rect 1080 49495 1188 49571
rect 81432 49495 81540 49571
rect 0 49399 82620 49447
rect 0 49303 82620 49351
rect 1080 49179 1188 49255
rect 81432 49179 81540 49255
rect 0 49083 82620 49131
rect 1080 48925 1188 49035
rect 81432 48925 81540 49035
rect 0 48829 82620 48877
rect 1080 48705 1188 48781
rect 81432 48705 81540 48781
rect 0 48609 82620 48657
rect 0 48513 82620 48561
rect 1080 48389 1188 48465
rect 81432 48389 81540 48465
rect 0 48293 82620 48341
rect 1080 48135 1188 48245
rect 81432 48135 81540 48245
rect 0 48039 82620 48087
rect 1080 47915 1188 47991
rect 81432 47915 81540 47991
rect 0 47819 82620 47867
rect 0 47723 82620 47771
rect 1080 47599 1188 47675
rect 81432 47599 81540 47675
rect 0 47503 82620 47551
rect 1080 47345 1188 47455
rect 81432 47345 81540 47455
rect 0 47249 82620 47297
rect 1080 47125 1188 47201
rect 81432 47125 81540 47201
rect 0 47029 82620 47077
rect 0 46933 82620 46981
rect 1080 46809 1188 46885
rect 81432 46809 81540 46885
rect 0 46713 82620 46761
rect 1080 46555 1188 46665
rect 81432 46555 81540 46665
rect 0 46459 82620 46507
rect 1080 46335 1188 46411
rect 81432 46335 81540 46411
rect 0 46239 82620 46287
rect 0 46143 82620 46191
rect 1080 46019 1188 46095
rect 81432 46019 81540 46095
rect 0 45923 82620 45971
rect 1080 45765 1188 45875
rect 81432 45765 81540 45875
rect 0 45669 82620 45717
rect 1080 45545 1188 45621
rect 81432 45545 81540 45621
rect 0 45449 82620 45497
rect 0 45353 82620 45401
rect 1080 45229 1188 45305
rect 81432 45229 81540 45305
rect 0 45133 82620 45181
rect 1080 44975 1188 45085
rect 81432 44975 81540 45085
rect 0 44879 82620 44927
rect 1080 44755 1188 44831
rect 81432 44755 81540 44831
rect 0 44659 82620 44707
rect 0 44563 82620 44611
rect 1080 44439 1188 44515
rect 81432 44439 81540 44515
rect 0 44343 82620 44391
rect 1080 44185 1188 44295
rect 81432 44185 81540 44295
rect 0 44089 82620 44137
rect 1080 43965 1188 44041
rect 81432 43965 81540 44041
rect 0 43869 82620 43917
rect 0 43773 82620 43821
rect 1080 43649 1188 43725
rect 81432 43649 81540 43725
rect 0 43553 82620 43601
rect 1080 43395 1188 43505
rect 81432 43395 81540 43505
rect 0 43299 82620 43347
rect 1080 43175 1188 43251
rect 81432 43175 81540 43251
rect 0 43079 82620 43127
rect 0 42983 82620 43031
rect 1080 42859 1188 42935
rect 81432 42859 81540 42935
rect 0 42763 82620 42811
rect 1080 42605 1188 42715
rect 81432 42605 81540 42715
rect 0 42509 82620 42557
rect 1080 42385 1188 42461
rect 81432 42385 81540 42461
rect 0 42289 82620 42337
rect 0 42193 82620 42241
rect 1080 42069 1188 42145
rect 81432 42069 81540 42145
rect 0 41973 82620 42021
rect 1080 41815 1188 41925
rect 81432 41815 81540 41925
rect 0 41719 82620 41767
rect 1080 41595 1188 41671
rect 81432 41595 81540 41671
rect 0 41499 82620 41547
rect 0 41403 82620 41451
rect 1080 41279 1188 41355
rect 81432 41279 81540 41355
rect 0 41183 82620 41231
rect 1080 41025 1188 41135
rect 81432 41025 81540 41135
rect 0 40929 82620 40977
rect 1080 40805 1188 40881
rect 81432 40805 81540 40881
rect 0 40709 82620 40757
rect 0 40613 82620 40661
rect 1080 40489 1188 40565
rect 81432 40489 81540 40565
rect 0 40393 82620 40441
rect 1080 40235 1188 40345
rect 81432 40235 81540 40345
rect 0 40139 82620 40187
rect 1080 40015 1188 40091
rect 81432 40015 81540 40091
rect 0 39919 82620 39967
rect 0 39823 82620 39871
rect 1080 39699 1188 39775
rect 81432 39699 81540 39775
rect 0 39603 82620 39651
rect 1080 39445 1188 39555
rect 81432 39445 81540 39555
rect 0 39349 82620 39397
rect 1080 39225 1188 39301
rect 81432 39225 81540 39301
rect 0 39129 82620 39177
rect 0 39033 82620 39081
rect 1080 38909 1188 38985
rect 81432 38909 81540 38985
rect 0 38813 82620 38861
rect 1080 38655 1188 38765
rect 81432 38655 81540 38765
rect 0 38559 82620 38607
rect 1080 38435 1188 38511
rect 81432 38435 81540 38511
rect 0 38339 82620 38387
rect 0 38243 82620 38291
rect 1080 38119 1188 38195
rect 81432 38119 81540 38195
rect 0 38023 82620 38071
rect 1080 37865 1188 37975
rect 81432 37865 81540 37975
rect 0 37769 82620 37817
rect 1080 37645 1188 37721
rect 81432 37645 81540 37721
rect 0 37549 82620 37597
rect 0 37453 82620 37501
rect 1080 37329 1188 37405
rect 81432 37329 81540 37405
rect 0 37233 82620 37281
rect 1080 37075 1188 37185
rect 81432 37075 81540 37185
rect 0 36979 82620 37027
rect 1080 36855 1188 36931
rect 81432 36855 81540 36931
rect 0 36759 82620 36807
rect 0 36663 82620 36711
rect 1080 36539 1188 36615
rect 81432 36539 81540 36615
rect 0 36443 82620 36491
rect 1080 36285 1188 36395
rect 81432 36285 81540 36395
rect 0 36189 82620 36237
rect 1080 36065 1188 36141
rect 81432 36065 81540 36141
rect 0 35969 82620 36017
rect 0 35873 82620 35921
rect 1080 35749 1188 35825
rect 81432 35749 81540 35825
rect 0 35653 82620 35701
rect 1080 35495 1188 35605
rect 81432 35495 81540 35605
rect 0 35399 82620 35447
rect 1080 35275 1188 35351
rect 81432 35275 81540 35351
rect 0 35179 82620 35227
rect 0 35083 82620 35131
rect 1080 34959 1188 35035
rect 81432 34959 81540 35035
rect 0 34863 82620 34911
rect 1080 34705 1188 34815
rect 81432 34705 81540 34815
rect 0 34609 82620 34657
rect 1080 34485 1188 34561
rect 81432 34485 81540 34561
rect 0 34389 82620 34437
rect 0 34293 82620 34341
rect 1080 34169 1188 34245
rect 81432 34169 81540 34245
rect 0 34073 82620 34121
rect 1080 33915 1188 34025
rect 81432 33915 81540 34025
rect 0 33819 82620 33867
rect 1080 33695 1188 33771
rect 81432 33695 81540 33771
rect 0 33599 82620 33647
rect 0 33503 82620 33551
rect 1080 33379 1188 33455
rect 81432 33379 81540 33455
rect 0 33283 82620 33331
rect 1080 33125 1188 33235
rect 81432 33125 81540 33235
rect 0 33029 82620 33077
rect 1080 32905 1188 32981
rect 81432 32905 81540 32981
rect 0 32809 82620 32857
rect 0 32713 82620 32761
rect 1080 32589 1188 32665
rect 81432 32589 81540 32665
rect 0 32493 82620 32541
rect 1080 32335 1188 32445
rect 81432 32335 81540 32445
rect 0 32239 82620 32287
rect 1080 32115 1188 32191
rect 81432 32115 81540 32191
rect 0 32019 82620 32067
rect 0 31923 82620 31971
rect 1080 31799 1188 31875
rect 81432 31799 81540 31875
rect 0 31703 82620 31751
rect 1080 31545 1188 31655
rect 81432 31545 81540 31655
rect 0 31449 82620 31497
rect 1080 31325 1188 31401
rect 81432 31325 81540 31401
rect 0 31229 82620 31277
rect 0 31133 82620 31181
rect 1080 31009 1188 31085
rect 81432 31009 81540 31085
rect 0 30913 82620 30961
rect 1080 30755 1188 30865
rect 81432 30755 81540 30865
rect 0 30659 82620 30707
rect 1080 30535 1188 30611
rect 81432 30535 81540 30611
rect 0 30439 82620 30487
rect 0 30343 82620 30391
rect 1080 30219 1188 30295
rect 81432 30219 81540 30295
rect 0 30123 82620 30171
rect 1080 29965 1188 30075
rect 81432 29965 81540 30075
rect 0 29869 82620 29917
rect 1080 29745 1188 29821
rect 81432 29745 81540 29821
rect 0 29649 82620 29697
rect 0 29553 82620 29601
rect 1080 29429 1188 29505
rect 81432 29429 81540 29505
rect 0 29333 82620 29381
rect 1080 29175 1188 29285
rect 81432 29175 81540 29285
rect 0 29079 82620 29127
rect 1080 28955 1188 29031
rect 81432 28955 81540 29031
rect 0 28859 82620 28907
rect 0 28763 82620 28811
rect 1080 28639 1188 28715
rect 81432 28639 81540 28715
rect 0 28543 82620 28591
rect 1080 28385 1188 28495
rect 81432 28385 81540 28495
rect 0 28289 82620 28337
rect 1080 28165 1188 28241
rect 81432 28165 81540 28241
rect 0 28069 82620 28117
rect 0 27973 82620 28021
rect 1080 27849 1188 27925
rect 81432 27849 81540 27925
rect 0 27753 82620 27801
rect 1080 27595 1188 27705
rect 81432 27595 81540 27705
rect 0 27499 82620 27547
rect 1080 27375 1188 27451
rect 81432 27375 81540 27451
rect 0 27279 82620 27327
rect 0 27183 82620 27231
rect 1080 27059 1188 27135
rect 81432 27059 81540 27135
rect 0 26963 82620 27011
rect 1080 26805 1188 26915
rect 81432 26805 81540 26915
rect 0 26709 82620 26757
rect 1080 26585 1188 26661
rect 81432 26585 81540 26661
rect 0 26489 82620 26537
rect 0 26393 82620 26441
rect 1080 26269 1188 26345
rect 81432 26269 81540 26345
rect 0 26173 82620 26221
rect 1080 26015 1188 26125
rect 81432 26015 81540 26125
rect 0 25919 82620 25967
rect 1080 25795 1188 25871
rect 81432 25795 81540 25871
rect 0 25699 82620 25747
rect 0 25603 82620 25651
rect 1080 25479 1188 25555
rect 81432 25479 81540 25555
rect 0 25383 82620 25431
rect 1080 25225 1188 25335
rect 81432 25225 81540 25335
rect 0 25129 82620 25177
rect 1080 25005 1188 25081
rect 81432 25005 81540 25081
rect 0 24909 82620 24957
rect 0 24813 82620 24861
rect 1080 24689 1188 24765
rect 81432 24689 81540 24765
rect 0 24593 82620 24641
rect 1080 24435 1188 24545
rect 81432 24435 81540 24545
rect 0 24339 82620 24387
rect 1080 24215 1188 24291
rect 81432 24215 81540 24291
rect 0 24119 82620 24167
rect 0 24023 82620 24071
rect 1080 23899 1188 23975
rect 81432 23899 81540 23975
rect 0 23803 82620 23851
rect 1080 23645 1188 23755
rect 81432 23645 81540 23755
rect 0 23549 82620 23597
rect 1080 23425 1188 23501
rect 81432 23425 81540 23501
rect 0 23329 82620 23377
rect 0 23233 82620 23281
rect 1080 23109 1188 23185
rect 81432 23109 81540 23185
rect 0 23013 82620 23061
rect 1080 22855 1188 22965
rect 81432 22855 81540 22965
rect 0 22759 82620 22807
rect 1080 22635 1188 22711
rect 81432 22635 81540 22711
rect 0 22539 82620 22587
rect 0 22443 82620 22491
rect 1080 22319 1188 22395
rect 81432 22319 81540 22395
rect 0 22223 82620 22271
rect 1080 22065 1188 22175
rect 81432 22065 81540 22175
rect 0 21969 82620 22017
rect 1080 21845 1188 21921
rect 81432 21845 81540 21921
rect 0 21749 82620 21797
rect 0 21653 82620 21701
rect 1080 21529 1188 21605
rect 81432 21529 81540 21605
rect 0 21433 82620 21481
rect 1080 21275 1188 21385
rect 81432 21275 81540 21385
rect 0 21179 82620 21227
rect 1080 21055 1188 21131
rect 81432 21055 81540 21131
rect 0 20959 82620 21007
rect 0 20863 82620 20911
rect 1080 20739 1188 20815
rect 81432 20739 81540 20815
rect 0 20643 82620 20691
rect 1080 20485 1188 20595
rect 81432 20485 81540 20595
rect 0 20389 82620 20437
rect 1080 20265 1188 20341
rect 81432 20265 81540 20341
rect 0 20169 82620 20217
rect 0 20073 82620 20121
rect 1080 19949 1188 20025
rect 81432 19949 81540 20025
rect 0 19853 82620 19901
rect 1080 19695 1188 19805
rect 81432 19695 81540 19805
rect 0 19599 82620 19647
rect 1080 19475 1188 19551
rect 81432 19475 81540 19551
rect 0 19379 82620 19427
rect 0 19283 82620 19331
rect 1080 19159 1188 19235
rect 81432 19159 81540 19235
rect 0 19063 82620 19111
rect 1080 18905 1188 19015
rect 81432 18905 81540 19015
rect 0 18809 82620 18857
rect 1080 18685 1188 18761
rect 81432 18685 81540 18761
rect 0 18589 82620 18637
rect 0 18493 82620 18541
rect 1080 18369 1188 18445
rect 81432 18369 81540 18445
rect 0 18273 82620 18321
rect 1080 18115 1188 18225
rect 81432 18115 81540 18225
rect 0 18019 82620 18067
rect 1080 17895 1188 17971
rect 81432 17895 81540 17971
rect 0 17799 82620 17847
rect 0 17703 82620 17751
rect 1080 17579 1188 17655
rect 81432 17579 81540 17655
rect 0 17483 82620 17531
rect 1080 17325 1188 17435
rect 81432 17325 81540 17435
rect 0 17229 82620 17277
rect 1080 17105 1188 17181
rect 81432 17105 81540 17181
rect 0 17009 82620 17057
rect 0 16913 82620 16961
rect 1080 16789 1188 16865
rect 81432 16789 81540 16865
rect 0 16693 82620 16741
rect 1080 16535 1188 16645
rect 81432 16535 81540 16645
rect 0 16439 82620 16487
rect 1080 16315 1188 16391
rect 81432 16315 81540 16391
rect 0 16219 82620 16267
rect 0 16123 82620 16171
rect 1080 15999 1188 16075
rect 81432 15999 81540 16075
rect 0 15903 82620 15951
rect 1080 15745 1188 15855
rect 81432 15745 81540 15855
rect 0 15649 82620 15697
rect 1080 15525 1188 15601
rect 81432 15525 81540 15601
rect 0 15429 82620 15477
rect 0 15333 82620 15381
rect 1080 15209 1188 15285
rect 81432 15209 81540 15285
rect 0 15113 82620 15161
rect 1080 14955 1188 15065
rect 81432 14955 81540 15065
rect 0 14859 82620 14907
rect 1080 14735 1188 14811
rect 81432 14735 81540 14811
rect 0 14639 82620 14687
rect 0 14543 82620 14591
rect 1080 14419 1188 14495
rect 81432 14419 81540 14495
rect 0 14323 82620 14371
rect 1080 14165 1188 14275
rect 81432 14165 81540 14275
rect 0 14069 82620 14117
rect 1080 13945 1188 14021
rect 81432 13945 81540 14021
rect 0 13849 82620 13897
rect 0 13753 82620 13801
rect 1080 13629 1188 13705
rect 81432 13629 81540 13705
rect 0 13533 82620 13581
rect 1080 13375 1188 13485
rect 81432 13375 81540 13485
rect 0 13279 82620 13327
rect 1080 13155 1188 13231
rect 81432 13155 81540 13231
rect 0 13059 82620 13107
rect 0 12963 82620 13011
rect 1080 12839 1188 12915
rect 81432 12839 81540 12915
rect 0 12743 82620 12791
rect 1080 12585 1188 12695
rect 81432 12585 81540 12695
rect 0 12489 82620 12537
rect 1080 12365 1188 12441
rect 81432 12365 81540 12441
rect 0 12269 82620 12317
rect 0 12173 82620 12221
rect 1080 12049 1188 12125
rect 81432 12049 81540 12125
rect 0 11953 82620 12001
rect 1080 11795 1188 11905
rect 81432 11795 81540 11905
rect 0 11699 82620 11747
rect 1080 11575 1188 11651
rect 81432 11575 81540 11651
rect 0 11479 82620 11527
rect 0 11383 82620 11431
rect 1080 11259 1188 11335
rect 81432 11259 81540 11335
rect 0 11163 82620 11211
rect 1080 11005 1188 11115
rect 81432 11005 81540 11115
rect 0 10909 82620 10957
rect 1080 10785 1188 10861
rect 81432 10785 81540 10861
rect 0 10689 82620 10737
rect 0 10593 82620 10641
rect 1080 10469 1188 10545
rect 81432 10469 81540 10545
rect 0 10373 82620 10421
rect 1080 10215 1188 10325
rect 81432 10215 81540 10325
rect 0 10119 82620 10167
rect 1080 9995 1188 10071
rect 81432 9995 81540 10071
rect 0 9899 82620 9947
rect 0 9803 82620 9851
rect 1080 9679 1188 9755
rect 81432 9679 81540 9755
rect 0 9583 82620 9631
rect 1080 9425 1188 9535
rect 81432 9425 81540 9535
rect 0 9329 82620 9377
rect 1080 9205 1188 9281
rect 81432 9205 81540 9281
rect 0 9109 82620 9157
rect 0 9013 82620 9061
rect 1080 8889 1188 8965
rect 81432 8889 81540 8965
rect 0 8793 82620 8841
rect 1080 8635 1188 8745
rect 81432 8635 81540 8745
rect 0 8539 82620 8587
rect 1080 8415 1188 8491
rect 81432 8415 81540 8491
rect 0 8319 82620 8367
rect 0 8223 82620 8271
rect 1080 8099 1188 8175
rect 81432 8099 81540 8175
rect 0 8003 82620 8051
rect 1080 7845 1188 7955
rect 81432 7845 81540 7955
rect 0 7749 82620 7797
rect 1080 7625 1188 7701
rect 81432 7625 81540 7701
rect 0 7529 82620 7577
rect 0 7433 82620 7481
rect 1080 7309 1188 7385
rect 81432 7309 81540 7385
rect 0 7213 82620 7261
rect 1080 7055 1188 7165
rect 81432 7055 81540 7165
rect 0 6959 82620 7007
rect 1080 6835 1188 6911
rect 81432 6835 81540 6911
rect 0 6739 82620 6787
rect 0 6643 82620 6691
rect 1080 6519 1188 6595
rect 81432 6519 81540 6595
rect 0 6423 82620 6471
rect 1080 6265 1188 6375
rect 81432 6265 81540 6375
rect 0 6169 82620 6217
rect 1080 6045 1188 6121
rect 81432 6045 81540 6121
rect 0 5949 82620 5997
rect 0 5853 82620 5901
rect 1080 5729 1188 5805
rect 81432 5729 81540 5805
rect 0 5633 82620 5681
rect 1080 5475 1188 5585
rect 81432 5475 81540 5585
rect 0 5379 82620 5427
rect 1080 5255 1188 5331
rect 81432 5255 81540 5331
rect 0 5159 82620 5207
rect 0 5063 82620 5111
rect 1080 4939 1188 5015
rect 81432 4939 81540 5015
rect 0 4843 82620 4891
rect 1080 4685 1188 4795
rect 81432 4685 81540 4795
rect 0 4589 82620 4637
rect 1080 4465 1188 4541
rect 81432 4465 81540 4541
rect 0 4369 82620 4417
rect 0 4273 82620 4321
rect 1080 4149 1188 4225
rect 81432 4149 81540 4225
rect 0 4053 82620 4101
rect 1080 3895 1188 4005
rect 81432 3895 81540 4005
rect 0 3799 82620 3847
rect 1080 3675 1188 3751
rect 81432 3675 81540 3751
rect 0 3579 82620 3627
rect 0 3483 82620 3531
rect 1080 3359 1188 3435
rect 81432 3359 81540 3435
rect 0 3263 82620 3311
rect 1080 3105 1188 3215
rect 81432 3105 81540 3215
rect 0 3009 82620 3057
rect 1080 2885 1188 2961
rect 81432 2885 81540 2961
rect 0 2789 82620 2837
rect 0 2693 82620 2741
rect 1080 2569 1188 2645
rect 81432 2569 81540 2645
rect 0 2473 82620 2521
rect 1080 2315 1188 2425
rect 81432 2315 81540 2425
rect 0 2219 82620 2267
rect 1080 2095 1188 2171
rect 81432 2095 81540 2171
rect 0 1999 82620 2047
rect 0 1903 82620 1951
rect 1080 1779 1188 1855
rect 81432 1779 81540 1855
rect 0 1683 82620 1731
rect 1080 1525 1188 1635
rect 81432 1525 81540 1635
rect 0 1429 82620 1477
rect 1080 1305 1188 1381
rect 81432 1305 81540 1381
rect 0 1209 82620 1257
rect 0 1113 82620 1161
rect 1080 989 1188 1065
rect 81432 989 81540 1065
rect 0 893 82620 941
rect 1080 735 1188 845
rect 81432 735 81540 845
rect 0 682 82620 687
rect -37 645 82657 682
rect 0 639 82620 645
rect 1080 515 1188 591
rect 81432 515 81540 591
rect 0 419 82620 467
<< metal3 >>
rect 1013 51862 1111 51960
rect 1637 51862 1735 51960
rect 2261 51862 2359 51960
rect 2885 51862 2983 51960
rect 3509 51862 3607 51960
rect 4133 51862 4231 51960
rect 4757 51862 4855 51960
rect 5381 51862 5479 51960
rect 6005 51862 6103 51960
rect 6629 51862 6727 51960
rect 7253 51862 7351 51960
rect 7877 51862 7975 51960
rect 8501 51862 8599 51960
rect 9125 51862 9223 51960
rect 9749 51862 9847 51960
rect 10373 51862 10471 51960
rect 10997 51862 11095 51960
rect 11621 51862 11719 51960
rect 12245 51862 12343 51960
rect 12869 51862 12967 51960
rect 13493 51862 13591 51960
rect 14117 51862 14215 51960
rect 14741 51862 14839 51960
rect 15365 51862 15463 51960
rect 15989 51862 16087 51960
rect 16613 51862 16711 51960
rect 17237 51862 17335 51960
rect 17861 51862 17959 51960
rect 18485 51862 18583 51960
rect 19109 51862 19207 51960
rect 19733 51862 19831 51960
rect 20357 51862 20455 51960
rect 20981 51862 21079 51960
rect 21605 51862 21703 51960
rect 22229 51862 22327 51960
rect 22853 51862 22951 51960
rect 23477 51862 23575 51960
rect 24101 51862 24199 51960
rect 24725 51862 24823 51960
rect 25349 51862 25447 51960
rect 25973 51862 26071 51960
rect 26597 51862 26695 51960
rect 27221 51862 27319 51960
rect 27845 51862 27943 51960
rect 28469 51862 28567 51960
rect 29093 51862 29191 51960
rect 29717 51862 29815 51960
rect 30341 51862 30439 51960
rect 30965 51862 31063 51960
rect 31589 51862 31687 51960
rect 32213 51862 32311 51960
rect 32837 51862 32935 51960
rect 33461 51862 33559 51960
rect 34085 51862 34183 51960
rect 34709 51862 34807 51960
rect 35333 51862 35431 51960
rect 35957 51862 36055 51960
rect 36581 51862 36679 51960
rect 37205 51862 37303 51960
rect 37829 51862 37927 51960
rect 38453 51862 38551 51960
rect 39077 51862 39175 51960
rect 39701 51862 39799 51960
rect 40325 51862 40423 51960
rect 40949 51862 41047 51960
rect 41573 51862 41671 51960
rect 42197 51862 42295 51960
rect 42821 51862 42919 51960
rect 43445 51862 43543 51960
rect 44069 51862 44167 51960
rect 44693 51862 44791 51960
rect 45317 51862 45415 51960
rect 45941 51862 46039 51960
rect 46565 51862 46663 51960
rect 47189 51862 47287 51960
rect 47813 51862 47911 51960
rect 48437 51862 48535 51960
rect 49061 51862 49159 51960
rect 49685 51862 49783 51960
rect 50309 51862 50407 51960
rect 50933 51862 51031 51960
rect 51557 51862 51655 51960
rect 52181 51862 52279 51960
rect 52805 51862 52903 51960
rect 53429 51862 53527 51960
rect 54053 51862 54151 51960
rect 54677 51862 54775 51960
rect 55301 51862 55399 51960
rect 55925 51862 56023 51960
rect 56549 51862 56647 51960
rect 57173 51862 57271 51960
rect 57797 51862 57895 51960
rect 58421 51862 58519 51960
rect 59045 51862 59143 51960
rect 59669 51862 59767 51960
rect 60293 51862 60391 51960
rect 60917 51862 61015 51960
rect 61541 51862 61639 51960
rect 62165 51862 62263 51960
rect 62789 51862 62887 51960
rect 63413 51862 63511 51960
rect 64037 51862 64135 51960
rect 64661 51862 64759 51960
rect 65285 51862 65383 51960
rect 65909 51862 66007 51960
rect 66533 51862 66631 51960
rect 67157 51862 67255 51960
rect 67781 51862 67879 51960
rect 68405 51862 68503 51960
rect 69029 51862 69127 51960
rect 69653 51862 69751 51960
rect 70277 51862 70375 51960
rect 70901 51862 70999 51960
rect 71525 51862 71623 51960
rect 72149 51862 72247 51960
rect 72773 51862 72871 51960
rect 73397 51862 73495 51960
rect 74021 51862 74119 51960
rect 74645 51862 74743 51960
rect 75269 51862 75367 51960
rect 75893 51862 75991 51960
rect 76517 51862 76615 51960
rect 77141 51862 77239 51960
rect 77765 51862 77863 51960
rect 78389 51862 78487 51960
rect 79013 51862 79111 51960
rect 79637 51862 79735 51960
rect 80261 51862 80359 51960
rect 80885 51862 80983 51960
rect 81509 51862 81607 51960
rect -49 51648 49 51746
rect 82571 51648 82669 51746
rect 317 51301 415 51399
rect 82205 51301 82303 51399
rect 317 51064 415 51162
rect 82205 51064 82303 51162
rect 317 50748 415 50846
rect 82205 50748 82303 50846
rect 317 50511 415 50609
rect 82205 50511 82303 50609
rect 317 50274 415 50372
rect 82205 50274 82303 50372
rect 317 49958 415 50056
rect 82205 49958 82303 50056
rect 317 49721 415 49819
rect 82205 49721 82303 49819
rect 317 49484 415 49582
rect 82205 49484 82303 49582
rect 317 49168 415 49266
rect 82205 49168 82303 49266
rect 317 48931 415 49029
rect 82205 48931 82303 49029
rect 317 48694 415 48792
rect 82205 48694 82303 48792
rect 317 48378 415 48476
rect 82205 48378 82303 48476
rect 317 48141 415 48239
rect 82205 48141 82303 48239
rect 317 47904 415 48002
rect 82205 47904 82303 48002
rect 317 47588 415 47686
rect 82205 47588 82303 47686
rect 317 47351 415 47449
rect 82205 47351 82303 47449
rect 317 47114 415 47212
rect 82205 47114 82303 47212
rect 317 46798 415 46896
rect 82205 46798 82303 46896
rect 317 46561 415 46659
rect 82205 46561 82303 46659
rect 317 46324 415 46422
rect 82205 46324 82303 46422
rect 317 46008 415 46106
rect 82205 46008 82303 46106
rect 317 45771 415 45869
rect 82205 45771 82303 45869
rect 317 45534 415 45632
rect 82205 45534 82303 45632
rect 317 45218 415 45316
rect 82205 45218 82303 45316
rect 317 44981 415 45079
rect 82205 44981 82303 45079
rect 317 44744 415 44842
rect 82205 44744 82303 44842
rect 317 44428 415 44526
rect 82205 44428 82303 44526
rect 317 44191 415 44289
rect 82205 44191 82303 44289
rect 317 43954 415 44052
rect 82205 43954 82303 44052
rect 317 43638 415 43736
rect 82205 43638 82303 43736
rect 317 43401 415 43499
rect 82205 43401 82303 43499
rect 317 43164 415 43262
rect 82205 43164 82303 43262
rect 317 42848 415 42946
rect 82205 42848 82303 42946
rect 317 42611 415 42709
rect 82205 42611 82303 42709
rect 317 42374 415 42472
rect 82205 42374 82303 42472
rect 317 42058 415 42156
rect 82205 42058 82303 42156
rect 317 41821 415 41919
rect 82205 41821 82303 41919
rect 317 41584 415 41682
rect 82205 41584 82303 41682
rect 317 41268 415 41366
rect 82205 41268 82303 41366
rect 317 41031 415 41129
rect 82205 41031 82303 41129
rect 317 40794 415 40892
rect 82205 40794 82303 40892
rect 317 40478 415 40576
rect 82205 40478 82303 40576
rect 317 40241 415 40339
rect 82205 40241 82303 40339
rect 317 40004 415 40102
rect 82205 40004 82303 40102
rect 317 39688 415 39786
rect 82205 39688 82303 39786
rect 317 39451 415 39549
rect 82205 39451 82303 39549
rect 317 39214 415 39312
rect 82205 39214 82303 39312
rect 317 38898 415 38996
rect 82205 38898 82303 38996
rect 317 38661 415 38759
rect 82205 38661 82303 38759
rect 317 38424 415 38522
rect 82205 38424 82303 38522
rect 317 38108 415 38206
rect 82205 38108 82303 38206
rect 317 37871 415 37969
rect 82205 37871 82303 37969
rect 317 37634 415 37732
rect 82205 37634 82303 37732
rect 317 37318 415 37416
rect 82205 37318 82303 37416
rect 317 37081 415 37179
rect 82205 37081 82303 37179
rect 317 36844 415 36942
rect 82205 36844 82303 36942
rect 317 36528 415 36626
rect 82205 36528 82303 36626
rect 317 36291 415 36389
rect 82205 36291 82303 36389
rect 317 36054 415 36152
rect 82205 36054 82303 36152
rect 317 35738 415 35836
rect 82205 35738 82303 35836
rect 317 35501 415 35599
rect 82205 35501 82303 35599
rect 317 35264 415 35362
rect 82205 35264 82303 35362
rect 317 34948 415 35046
rect 82205 34948 82303 35046
rect 317 34711 415 34809
rect 82205 34711 82303 34809
rect 317 34474 415 34572
rect 82205 34474 82303 34572
rect 317 34158 415 34256
rect 82205 34158 82303 34256
rect 317 33921 415 34019
rect 82205 33921 82303 34019
rect 317 33684 415 33782
rect 82205 33684 82303 33782
rect 317 33368 415 33466
rect 82205 33368 82303 33466
rect 317 33131 415 33229
rect 82205 33131 82303 33229
rect 317 32894 415 32992
rect 82205 32894 82303 32992
rect 317 32578 415 32676
rect 82205 32578 82303 32676
rect 317 32341 415 32439
rect 82205 32341 82303 32439
rect 317 32104 415 32202
rect 82205 32104 82303 32202
rect 317 31788 415 31886
rect 82205 31788 82303 31886
rect 317 31551 415 31649
rect 82205 31551 82303 31649
rect 317 31314 415 31412
rect 82205 31314 82303 31412
rect 317 30998 415 31096
rect 82205 30998 82303 31096
rect 317 30761 415 30859
rect 82205 30761 82303 30859
rect 317 30524 415 30622
rect 82205 30524 82303 30622
rect 317 30208 415 30306
rect 82205 30208 82303 30306
rect 317 29971 415 30069
rect 82205 29971 82303 30069
rect 317 29734 415 29832
rect 82205 29734 82303 29832
rect 317 29418 415 29516
rect 82205 29418 82303 29516
rect 317 29181 415 29279
rect 82205 29181 82303 29279
rect 317 28944 415 29042
rect 82205 28944 82303 29042
rect 317 28628 415 28726
rect 82205 28628 82303 28726
rect 317 28391 415 28489
rect 82205 28391 82303 28489
rect 317 28154 415 28252
rect 82205 28154 82303 28252
rect 317 27838 415 27936
rect 82205 27838 82303 27936
rect 317 27601 415 27699
rect 82205 27601 82303 27699
rect 317 27364 415 27462
rect 82205 27364 82303 27462
rect 317 27048 415 27146
rect 82205 27048 82303 27146
rect 317 26811 415 26909
rect 82205 26811 82303 26909
rect 317 26574 415 26672
rect 82205 26574 82303 26672
rect 317 26258 415 26356
rect 82205 26258 82303 26356
rect 317 26021 415 26119
rect 82205 26021 82303 26119
rect 317 25784 415 25882
rect 82205 25784 82303 25882
rect 317 25468 415 25566
rect 82205 25468 82303 25566
rect 317 25231 415 25329
rect 82205 25231 82303 25329
rect 317 24994 415 25092
rect 82205 24994 82303 25092
rect 317 24678 415 24776
rect 82205 24678 82303 24776
rect 317 24441 415 24539
rect 82205 24441 82303 24539
rect 317 24204 415 24302
rect 82205 24204 82303 24302
rect 317 23888 415 23986
rect 82205 23888 82303 23986
rect 317 23651 415 23749
rect 82205 23651 82303 23749
rect 317 23414 415 23512
rect 82205 23414 82303 23512
rect 317 23098 415 23196
rect 82205 23098 82303 23196
rect 317 22861 415 22959
rect 82205 22861 82303 22959
rect 317 22624 415 22722
rect 82205 22624 82303 22722
rect 317 22308 415 22406
rect 82205 22308 82303 22406
rect 317 22071 415 22169
rect 82205 22071 82303 22169
rect 317 21834 415 21932
rect 82205 21834 82303 21932
rect 317 21518 415 21616
rect 82205 21518 82303 21616
rect 317 21281 415 21379
rect 82205 21281 82303 21379
rect 317 21044 415 21142
rect 82205 21044 82303 21142
rect 317 20728 415 20826
rect 82205 20728 82303 20826
rect 317 20491 415 20589
rect 82205 20491 82303 20589
rect 317 20254 415 20352
rect 82205 20254 82303 20352
rect 317 19938 415 20036
rect 82205 19938 82303 20036
rect 317 19701 415 19799
rect 82205 19701 82303 19799
rect 317 19464 415 19562
rect 82205 19464 82303 19562
rect 317 19148 415 19246
rect 82205 19148 82303 19246
rect 317 18911 415 19009
rect 82205 18911 82303 19009
rect 317 18674 415 18772
rect 82205 18674 82303 18772
rect 317 18358 415 18456
rect 82205 18358 82303 18456
rect 317 18121 415 18219
rect 82205 18121 82303 18219
rect 317 17884 415 17982
rect 82205 17884 82303 17982
rect 317 17568 415 17666
rect 82205 17568 82303 17666
rect 317 17331 415 17429
rect 82205 17331 82303 17429
rect 317 17094 415 17192
rect 82205 17094 82303 17192
rect 317 16778 415 16876
rect 82205 16778 82303 16876
rect 317 16541 415 16639
rect 82205 16541 82303 16639
rect 317 16304 415 16402
rect 82205 16304 82303 16402
rect 317 15988 415 16086
rect 82205 15988 82303 16086
rect 317 15751 415 15849
rect 82205 15751 82303 15849
rect 317 15514 415 15612
rect 82205 15514 82303 15612
rect 317 15198 415 15296
rect 82205 15198 82303 15296
rect 317 14961 415 15059
rect 82205 14961 82303 15059
rect 317 14724 415 14822
rect 82205 14724 82303 14822
rect 317 14408 415 14506
rect 82205 14408 82303 14506
rect 317 14171 415 14269
rect 82205 14171 82303 14269
rect 317 13934 415 14032
rect 82205 13934 82303 14032
rect 317 13618 415 13716
rect 82205 13618 82303 13716
rect 317 13381 415 13479
rect 82205 13381 82303 13479
rect 317 13144 415 13242
rect 82205 13144 82303 13242
rect 317 12828 415 12926
rect 82205 12828 82303 12926
rect 317 12591 415 12689
rect 82205 12591 82303 12689
rect 317 12354 415 12452
rect 82205 12354 82303 12452
rect 317 12038 415 12136
rect 82205 12038 82303 12136
rect 317 11801 415 11899
rect 82205 11801 82303 11899
rect 317 11564 415 11662
rect 82205 11564 82303 11662
rect 317 11248 415 11346
rect 82205 11248 82303 11346
rect 317 11011 415 11109
rect 82205 11011 82303 11109
rect 317 10774 415 10872
rect 82205 10774 82303 10872
rect 317 10458 415 10556
rect 82205 10458 82303 10556
rect 317 10221 415 10319
rect 82205 10221 82303 10319
rect 317 9984 415 10082
rect 82205 9984 82303 10082
rect 317 9668 415 9766
rect 82205 9668 82303 9766
rect 317 9431 415 9529
rect 82205 9431 82303 9529
rect 317 9194 415 9292
rect 82205 9194 82303 9292
rect 317 8878 415 8976
rect 82205 8878 82303 8976
rect 317 8641 415 8739
rect 82205 8641 82303 8739
rect 317 8404 415 8502
rect 82205 8404 82303 8502
rect 317 8088 415 8186
rect 82205 8088 82303 8186
rect 317 7851 415 7949
rect 82205 7851 82303 7949
rect 317 7614 415 7712
rect 82205 7614 82303 7712
rect 317 7298 415 7396
rect 82205 7298 82303 7396
rect 317 7061 415 7159
rect 82205 7061 82303 7159
rect 317 6824 415 6922
rect 82205 6824 82303 6922
rect 317 6508 415 6606
rect 82205 6508 82303 6606
rect 317 6271 415 6369
rect 82205 6271 82303 6369
rect 317 6034 415 6132
rect 82205 6034 82303 6132
rect 317 5718 415 5816
rect 82205 5718 82303 5816
rect 317 5481 415 5579
rect 82205 5481 82303 5579
rect 317 5244 415 5342
rect 82205 5244 82303 5342
rect 317 4928 415 5026
rect 82205 4928 82303 5026
rect 317 4691 415 4789
rect 82205 4691 82303 4789
rect 317 4454 415 4552
rect 82205 4454 82303 4552
rect 317 4138 415 4236
rect 82205 4138 82303 4236
rect 317 3901 415 3999
rect 82205 3901 82303 3999
rect 317 3664 415 3762
rect 82205 3664 82303 3762
rect 317 3348 415 3446
rect 82205 3348 82303 3446
rect 317 3111 415 3209
rect 82205 3111 82303 3209
rect 317 2874 415 2972
rect 82205 2874 82303 2972
rect 317 2558 415 2656
rect 82205 2558 82303 2656
rect 317 2321 415 2419
rect 82205 2321 82303 2419
rect 317 2084 415 2182
rect 82205 2084 82303 2182
rect 317 1768 415 1866
rect 82205 1768 82303 1866
rect 317 1531 415 1629
rect 82205 1531 82303 1629
rect 317 1294 415 1392
rect 82205 1294 82303 1392
rect 317 978 415 1076
rect 82205 978 82303 1076
rect 317 741 415 839
rect 82205 741 82303 839
rect -49 614 49 712
rect 82571 614 82669 712
rect 1013 180 1111 278
rect 1637 180 1735 278
rect 2261 180 2359 278
rect 2885 180 2983 278
rect 3509 180 3607 278
rect 4133 180 4231 278
rect 4757 180 4855 278
rect 5381 180 5479 278
rect 6005 180 6103 278
rect 6629 180 6727 278
rect 7253 180 7351 278
rect 7877 180 7975 278
rect 8501 180 8599 278
rect 9125 180 9223 278
rect 9749 180 9847 278
rect 10373 180 10471 278
rect 10997 180 11095 278
rect 11621 180 11719 278
rect 12245 180 12343 278
rect 12869 180 12967 278
rect 13493 180 13591 278
rect 14117 180 14215 278
rect 14741 180 14839 278
rect 15365 180 15463 278
rect 15989 180 16087 278
rect 16613 180 16711 278
rect 17237 180 17335 278
rect 17861 180 17959 278
rect 18485 180 18583 278
rect 19109 180 19207 278
rect 19733 180 19831 278
rect 20357 180 20455 278
rect 20981 180 21079 278
rect 21605 180 21703 278
rect 22229 180 22327 278
rect 22853 180 22951 278
rect 23477 180 23575 278
rect 24101 180 24199 278
rect 24725 180 24823 278
rect 25349 180 25447 278
rect 25973 180 26071 278
rect 26597 180 26695 278
rect 27221 180 27319 278
rect 27845 180 27943 278
rect 28469 180 28567 278
rect 29093 180 29191 278
rect 29717 180 29815 278
rect 30341 180 30439 278
rect 30965 180 31063 278
rect 31589 180 31687 278
rect 32213 180 32311 278
rect 32837 180 32935 278
rect 33461 180 33559 278
rect 34085 180 34183 278
rect 34709 180 34807 278
rect 35333 180 35431 278
rect 35957 180 36055 278
rect 36581 180 36679 278
rect 37205 180 37303 278
rect 37829 180 37927 278
rect 38453 180 38551 278
rect 39077 180 39175 278
rect 39701 180 39799 278
rect 40325 180 40423 278
rect 40949 180 41047 278
rect 41573 180 41671 278
rect 42197 180 42295 278
rect 42821 180 42919 278
rect 43445 180 43543 278
rect 44069 180 44167 278
rect 44693 180 44791 278
rect 45317 180 45415 278
rect 45941 180 46039 278
rect 46565 180 46663 278
rect 47189 180 47287 278
rect 47813 180 47911 278
rect 48437 180 48535 278
rect 49061 180 49159 278
rect 49685 180 49783 278
rect 50309 180 50407 278
rect 50933 180 51031 278
rect 51557 180 51655 278
rect 52181 180 52279 278
rect 52805 180 52903 278
rect 53429 180 53527 278
rect 54053 180 54151 278
rect 54677 180 54775 278
rect 55301 180 55399 278
rect 55925 180 56023 278
rect 56549 180 56647 278
rect 57173 180 57271 278
rect 57797 180 57895 278
rect 58421 180 58519 278
rect 59045 180 59143 278
rect 59669 180 59767 278
rect 60293 180 60391 278
rect 60917 180 61015 278
rect 61541 180 61639 278
rect 62165 180 62263 278
rect 62789 180 62887 278
rect 63413 180 63511 278
rect 64037 180 64135 278
rect 64661 180 64759 278
rect 65285 180 65383 278
rect 65909 180 66007 278
rect 66533 180 66631 278
rect 67157 180 67255 278
rect 67781 180 67879 278
rect 68405 180 68503 278
rect 69029 180 69127 278
rect 69653 180 69751 278
rect 70277 180 70375 278
rect 70901 180 70999 278
rect 71525 180 71623 278
rect 72149 180 72247 278
rect 72773 180 72871 278
rect 73397 180 73495 278
rect 74021 180 74119 278
rect 74645 180 74743 278
rect 75269 180 75367 278
rect 75893 180 75991 278
rect 76517 180 76615 278
rect 77141 180 77239 278
rect 77765 180 77863 278
rect 78389 180 78487 278
rect 79013 180 79111 278
rect 79637 180 79735 278
rect 80261 180 80359 278
rect 80885 180 80983 278
rect 81509 180 81607 278
use sky130_sram_2kbyte_1rw1r_32x512_8_row_cap_array  sky130_sram_2kbyte_1rw1r_32x512_8_row_cap_array_0
timestamp 1626065694
transform 1 0 126 0 1 0
box -42 419 624 51721
use sky130_sram_2kbyte_1rw1r_32x512_8_row_cap_array_0  sky130_sram_2kbyte_1rw1r_32x512_8_row_cap_array_0_0
timestamp 1626065694
transform 1 0 81870 0 1 0
box 0 419 666 51721
use sky130_sram_2kbyte_1rw1r_32x512_8_col_cap_array_0  sky130_sram_2kbyte_1rw1r_32x512_8_col_cap_array_0_0
timestamp 1626065694
transform 1 0 1374 0 1 0
box 0 0 79872 474
use sky130_sram_2kbyte_1rw1r_32x512_8_col_cap_array  sky130_sram_2kbyte_1rw1r_32x512_8_col_cap_array_0
timestamp 1626065694
transform 1 0 1374 0 -1 52140
box 0 0 79872 474
use sky130_sram_2kbyte_1rw1r_32x512_8_dummy_array  sky130_sram_2kbyte_1rw1r_32x512_8_dummy_array_1
timestamp 1626065694
transform 1 0 1374 0 -1 790
box -42 -105 79914 421
use sky130_sram_2kbyte_1rw1r_32x512_8_dummy_array  sky130_sram_2kbyte_1rw1r_32x512_8_dummy_array_0
timestamp 1626065694
transform 1 0 1374 0 1 51350
box -42 -105 79914 421
use sky130_sram_2kbyte_1rw1r_32x512_8_replica_column  sky130_sram_2kbyte_1rw1r_32x512_8_replica_column_0
timestamp 1626065694
transform 1 0 750 0 1 0
box -26 0 666 52140
use sky130_sram_2kbyte_1rw1r_32x512_8_replica_column_0  sky130_sram_2kbyte_1rw1r_32x512_8_replica_column_0_0
timestamp 1626065694
transform 1 0 81246 0 1 0
box -42 0 650 52140
use sky130_sram_2kbyte_1rw1r_32x512_8_bitcell_array  sky130_sram_2kbyte_1rw1r_32x512_8_bitcell_array_0
timestamp 1626065694
transform 1 0 1374 0 1 790
box -42 -105 79914 50665
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_9  sky130_sram_2kbyte_1rw1r_32x512_8_contact_9_3
timestamp 1626065694
transform 1 0 -37 0 1 630
box 0 0 74 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_9  sky130_sram_2kbyte_1rw1r_32x512_8_contact_9_2
timestamp 1626065694
transform 1 0 82583 0 1 630
box 0 0 74 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_9  sky130_sram_2kbyte_1rw1r_32x512_8_contact_9_1
timestamp 1626065694
transform 1 0 -37 0 1 51664
box 0 0 74 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_9  sky130_sram_2kbyte_1rw1r_32x512_8_contact_9_0
timestamp 1626065694
transform 1 0 82583 0 1 51664
box 0 0 74 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_8  sky130_sram_2kbyte_1rw1r_32x512_8_contact_8_3
timestamp 1626065694
transform 1 0 -32 0 1 637
box 0 0 64 52
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_8  sky130_sram_2kbyte_1rw1r_32x512_8_contact_8_2
timestamp 1626065694
transform 1 0 82588 0 1 637
box 0 0 64 52
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_8  sky130_sram_2kbyte_1rw1r_32x512_8_contact_8_1
timestamp 1626065694
transform 1 0 -32 0 1 51671
box 0 0 64 52
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_8  sky130_sram_2kbyte_1rw1r_32x512_8_contact_8_0
timestamp 1626065694
transform 1 0 82588 0 1 51671
box 0 0 64 52
<< labels >>
rlabel metal3 s 80885 51862 80983 51960 4 vdd
rlabel metal3 s 74021 51862 74119 51960 4 vdd
rlabel metal3 s 75269 51862 75367 51960 4 vdd
rlabel metal3 s 66533 51862 66631 51960 4 vdd
rlabel metal3 s 79013 51862 79111 51960 4 vdd
rlabel metal3 s 64661 51862 64759 51960 4 vdd
rlabel metal3 s 63413 51862 63511 51960 4 vdd
rlabel metal3 s 67157 51862 67255 51960 4 vdd
rlabel metal3 s 62165 51862 62263 51960 4 vdd
rlabel metal3 s 73397 51862 73495 51960 4 vdd
rlabel metal3 s 71525 51862 71623 51960 4 vdd
rlabel metal3 s 67781 51862 67879 51960 4 vdd
rlabel metal3 s 72773 51862 72871 51960 4 vdd
rlabel metal3 s 77141 51862 77239 51960 4 vdd
rlabel metal3 s 62789 51862 62887 51960 4 vdd
rlabel metal3 s 64037 51862 64135 51960 4 vdd
rlabel metal3 s 72149 51862 72247 51960 4 vdd
rlabel metal3 s 70901 51862 70999 51960 4 vdd
rlabel metal3 s 81509 51862 81607 51960 4 vdd
rlabel metal3 s 77765 51862 77863 51960 4 vdd
rlabel metal3 s 69029 51862 69127 51960 4 vdd
rlabel metal3 s 74645 51862 74743 51960 4 vdd
rlabel metal3 s 69653 51862 69751 51960 4 vdd
rlabel metal3 s 76517 51862 76615 51960 4 vdd
rlabel metal3 s 80261 51862 80359 51960 4 vdd
rlabel metal3 s 65909 51862 66007 51960 4 vdd
rlabel metal3 s 79637 51862 79735 51960 4 vdd
rlabel metal3 s 65285 51862 65383 51960 4 vdd
rlabel metal3 s 78389 51862 78487 51960 4 vdd
rlabel metal3 s 75893 51862 75991 51960 4 vdd
rlabel metal3 s 70277 51862 70375 51960 4 vdd
rlabel metal3 s 68405 51862 68503 51960 4 vdd
rlabel metal3 s 82205 49721 82303 49819 4 gnd
rlabel metal3 s 82205 41821 82303 41919 4 gnd
rlabel metal3 s 82205 46561 82303 46659 4 gnd
rlabel metal3 s 82205 49958 82303 50056 4 gnd
rlabel metal3 s 82205 43164 82303 43262 4 gnd
rlabel metal3 s 82205 45771 82303 45869 4 gnd
rlabel metal3 s 82205 40478 82303 40576 4 gnd
rlabel metal3 s 82205 47351 82303 47449 4 gnd
rlabel metal3 s 82205 42058 82303 42156 4 gnd
rlabel metal3 s 82205 50511 82303 50609 4 gnd
rlabel metal3 s 82205 41268 82303 41366 4 gnd
rlabel metal3 s 82205 51064 82303 51162 4 gnd
rlabel metal3 s 82205 45218 82303 45316 4 gnd
rlabel metal3 s 82205 47588 82303 47686 4 gnd
rlabel metal3 s 82205 46798 82303 46896 4 gnd
rlabel metal3 s 82205 48141 82303 48239 4 gnd
rlabel metal3 s 82205 42848 82303 42946 4 gnd
rlabel metal3 s 82205 39451 82303 39549 4 gnd
rlabel metal3 s 82205 44428 82303 44526 4 gnd
rlabel metal3 s 82205 44981 82303 45079 4 gnd
rlabel metal3 s 82205 46324 82303 46422 4 gnd
rlabel metal3 s 82205 48694 82303 48792 4 gnd
rlabel metal3 s 82205 40241 82303 40339 4 gnd
rlabel metal3 s 82205 47114 82303 47212 4 gnd
rlabel metal3 s 82205 50748 82303 50846 4 gnd
rlabel metal3 s 82205 46008 82303 46106 4 gnd
rlabel metal3 s 82205 45534 82303 45632 4 gnd
rlabel metal3 s 82205 42611 82303 42709 4 gnd
rlabel metal3 s 82205 39688 82303 39786 4 gnd
rlabel metal3 s 82205 40004 82303 40102 4 gnd
rlabel metal3 s 82205 47904 82303 48002 4 gnd
rlabel metal3 s 82205 40794 82303 40892 4 gnd
rlabel metal3 s 82205 43954 82303 44052 4 gnd
rlabel metal3 s 82205 44744 82303 44842 4 gnd
rlabel metal3 s 82205 48378 82303 48476 4 gnd
rlabel metal3 s 82205 41031 82303 41129 4 gnd
rlabel metal3 s 82205 42374 82303 42472 4 gnd
rlabel metal3 s 82205 49168 82303 49266 4 gnd
rlabel metal3 s 82205 48931 82303 49029 4 gnd
rlabel metal3 s 82205 39214 82303 39312 4 gnd
rlabel metal3 s 82205 44191 82303 44289 4 gnd
rlabel metal3 s 82205 51301 82303 51399 4 gnd
rlabel metal3 s 82205 50274 82303 50372 4 gnd
rlabel metal3 s 82205 49484 82303 49582 4 gnd
rlabel metal3 s 82571 51648 82669 51746 4 gnd
rlabel metal3 s 82205 43638 82303 43736 4 gnd
rlabel metal3 s 82205 43401 82303 43499 4 gnd
rlabel metal3 s 82205 41584 82303 41682 4 gnd
rlabel metal3 s 52805 51862 52903 51960 4 vdd
rlabel metal3 s 42821 51862 42919 51960 4 vdd
rlabel metal3 s 59669 51862 59767 51960 4 vdd
rlabel metal3 s 49061 51862 49159 51960 4 vdd
rlabel metal3 s 61541 51862 61639 51960 4 vdd
rlabel metal3 s 51557 51862 51655 51960 4 vdd
rlabel metal3 s 42197 51862 42295 51960 4 vdd
rlabel metal3 s 47189 51862 47287 51960 4 vdd
rlabel metal3 s 48437 51862 48535 51960 4 vdd
rlabel metal3 s 54053 51862 54151 51960 4 vdd
rlabel metal3 s 53429 51862 53527 51960 4 vdd
rlabel metal3 s 58421 51862 58519 51960 4 vdd
rlabel metal3 s 50309 51862 50407 51960 4 vdd
rlabel metal3 s 57173 51862 57271 51960 4 vdd
rlabel metal3 s 57797 51862 57895 51960 4 vdd
rlabel metal3 s 45941 51862 46039 51960 4 vdd
rlabel metal3 s 50933 51862 51031 51960 4 vdd
rlabel metal3 s 44693 51862 44791 51960 4 vdd
rlabel metal3 s 54677 51862 54775 51960 4 vdd
rlabel metal3 s 44069 51862 44167 51960 4 vdd
rlabel metal3 s 49685 51862 49783 51960 4 vdd
rlabel metal3 s 45317 51862 45415 51960 4 vdd
rlabel metal3 s 55301 51862 55399 51960 4 vdd
rlabel metal3 s 60917 51862 61015 51960 4 vdd
rlabel metal3 s 59045 51862 59143 51960 4 vdd
rlabel metal3 s 41573 51862 41671 51960 4 vdd
rlabel metal3 s 46565 51862 46663 51960 4 vdd
rlabel metal3 s 43445 51862 43543 51960 4 vdd
rlabel metal3 s 47813 51862 47911 51960 4 vdd
rlabel metal3 s 60293 51862 60391 51960 4 vdd
rlabel metal3 s 52181 51862 52279 51960 4 vdd
rlabel metal3 s 56549 51862 56647 51960 4 vdd
rlabel metal3 s 55925 51862 56023 51960 4 vdd
rlabel metal3 s 82205 31314 82303 31412 4 gnd
rlabel metal3 s 82205 35501 82303 35599 4 gnd
rlabel metal3 s 82205 37318 82303 37416 4 gnd
rlabel metal3 s 82205 28391 82303 28489 4 gnd
rlabel metal3 s 82205 36528 82303 36626 4 gnd
rlabel metal3 s 82205 37871 82303 37969 4 gnd
rlabel metal3 s 82205 38661 82303 38759 4 gnd
rlabel metal3 s 82205 26811 82303 26909 4 gnd
rlabel metal3 s 82205 27048 82303 27146 4 gnd
rlabel metal3 s 82205 28944 82303 29042 4 gnd
rlabel metal3 s 82205 29971 82303 30069 4 gnd
rlabel metal3 s 82205 37081 82303 37179 4 gnd
rlabel metal3 s 82205 27364 82303 27462 4 gnd
rlabel metal3 s 82205 30208 82303 30306 4 gnd
rlabel metal3 s 82205 30998 82303 31096 4 gnd
rlabel metal3 s 82205 32104 82303 32202 4 gnd
rlabel metal3 s 82205 29418 82303 29516 4 gnd
rlabel metal3 s 82205 34474 82303 34572 4 gnd
rlabel metal3 s 82205 29181 82303 29279 4 gnd
rlabel metal3 s 82205 30761 82303 30859 4 gnd
rlabel metal3 s 82205 33131 82303 33229 4 gnd
rlabel metal3 s 82205 32578 82303 32676 4 gnd
rlabel metal3 s 82205 34948 82303 35046 4 gnd
rlabel metal3 s 82205 33368 82303 33466 4 gnd
rlabel metal3 s 82205 28628 82303 28726 4 gnd
rlabel metal3 s 82205 36054 82303 36152 4 gnd
rlabel metal3 s 82205 27601 82303 27699 4 gnd
rlabel metal3 s 82205 26574 82303 26672 4 gnd
rlabel metal3 s 82205 36844 82303 36942 4 gnd
rlabel metal3 s 82205 28154 82303 28252 4 gnd
rlabel metal3 s 82205 38424 82303 38522 4 gnd
rlabel metal3 s 82205 37634 82303 37732 4 gnd
rlabel metal3 s 82205 30524 82303 30622 4 gnd
rlabel metal3 s 82205 34158 82303 34256 4 gnd
rlabel metal3 s 82205 38898 82303 38996 4 gnd
rlabel metal3 s 82205 35264 82303 35362 4 gnd
rlabel metal3 s 82205 36291 82303 36389 4 gnd
rlabel metal3 s 82205 29734 82303 29832 4 gnd
rlabel metal3 s 82205 38108 82303 38206 4 gnd
rlabel metal3 s 82205 34711 82303 34809 4 gnd
rlabel metal3 s 82205 27838 82303 27936 4 gnd
rlabel metal3 s 82205 33921 82303 34019 4 gnd
rlabel metal3 s 82205 31788 82303 31886 4 gnd
rlabel metal3 s 82205 32341 82303 32439 4 gnd
rlabel metal3 s 82205 35738 82303 35836 4 gnd
rlabel metal3 s 82205 26258 82303 26356 4 gnd
rlabel metal3 s 82205 33684 82303 33782 4 gnd
rlabel metal3 s 82205 32894 82303 32992 4 gnd
rlabel metal3 s 82205 31551 82303 31649 4 gnd
rlabel metal3 s 31589 51862 31687 51960 4 vdd
rlabel metal3 s 30965 51862 31063 51960 4 vdd
rlabel metal3 s 37205 51862 37303 51960 4 vdd
rlabel metal3 s 21605 51862 21703 51960 4 vdd
rlabel metal3 s 36581 51862 36679 51960 4 vdd
rlabel metal3 s 39077 51862 39175 51960 4 vdd
rlabel metal3 s 32837 51862 32935 51960 4 vdd
rlabel metal3 s 30341 51862 30439 51960 4 vdd
rlabel metal3 s 27845 51862 27943 51960 4 vdd
rlabel metal3 s 29093 51862 29191 51960 4 vdd
rlabel metal3 s 24101 51862 24199 51960 4 vdd
rlabel metal3 s 25973 51862 26071 51960 4 vdd
rlabel metal3 s 39701 51862 39799 51960 4 vdd
rlabel metal3 s 28469 51862 28567 51960 4 vdd
rlabel metal3 s 35957 51862 36055 51960 4 vdd
rlabel metal3 s 38453 51862 38551 51960 4 vdd
rlabel metal3 s 24725 51862 24823 51960 4 vdd
rlabel metal3 s 40949 51862 41047 51960 4 vdd
rlabel metal3 s 33461 51862 33559 51960 4 vdd
rlabel metal3 s 26597 51862 26695 51960 4 vdd
rlabel metal3 s 35333 51862 35431 51960 4 vdd
rlabel metal3 s 22853 51862 22951 51960 4 vdd
rlabel metal3 s 40325 51862 40423 51960 4 vdd
rlabel metal3 s 27221 51862 27319 51960 4 vdd
rlabel metal3 s 23477 51862 23575 51960 4 vdd
rlabel metal3 s 34709 51862 34807 51960 4 vdd
rlabel metal3 s 25349 51862 25447 51960 4 vdd
rlabel metal3 s 32213 51862 32311 51960 4 vdd
rlabel metal3 s 20981 51862 21079 51960 4 vdd
rlabel metal3 s 29717 51862 29815 51960 4 vdd
rlabel metal3 s 34085 51862 34183 51960 4 vdd
rlabel metal3 s 37829 51862 37927 51960 4 vdd
rlabel metal3 s 22229 51862 22327 51960 4 vdd
rlabel metal3 s 317 43638 415 43736 4 gnd
rlabel metal3 s 12869 51862 12967 51960 4 vdd
rlabel metal3 s 317 43164 415 43262 4 gnd
rlabel metal3 s 317 48694 415 48792 4 gnd
rlabel metal3 s 317 44191 415 44289 4 gnd
rlabel metal3 s 317 40794 415 40892 4 gnd
rlabel metal3 s 317 39451 415 39549 4 gnd
rlabel metal3 s 2261 51862 2359 51960 4 vdd
rlabel metal3 s 317 41584 415 41682 4 gnd
rlabel metal3 s 317 45771 415 45869 4 gnd
rlabel metal3 s 3509 51862 3607 51960 4 vdd
rlabel metal3 s 317 49484 415 49582 4 gnd
rlabel metal3 s 7877 51862 7975 51960 4 vdd
rlabel metal3 s -49 51648 49 51746 4 gnd
rlabel metal3 s 11621 51862 11719 51960 4 vdd
rlabel metal3 s 317 44428 415 44526 4 gnd
rlabel metal3 s 18485 51862 18583 51960 4 vdd
rlabel metal3 s 15365 51862 15463 51960 4 vdd
rlabel metal3 s 317 46798 415 46896 4 gnd
rlabel metal3 s 317 46561 415 46659 4 gnd
rlabel metal3 s 1637 51862 1735 51960 4 vdd
rlabel metal3 s 13493 51862 13591 51960 4 vdd
rlabel metal3 s 317 50511 415 50609 4 gnd
rlabel metal3 s 6629 51862 6727 51960 4 vdd
rlabel metal3 s 19109 51862 19207 51960 4 vdd
rlabel metal3 s 317 42611 415 42709 4 gnd
rlabel metal3 s 8501 51862 8599 51960 4 vdd
rlabel metal3 s 4757 51862 4855 51960 4 vdd
rlabel metal3 s 14741 51862 14839 51960 4 vdd
rlabel metal3 s 14117 51862 14215 51960 4 vdd
rlabel metal3 s 10997 51862 11095 51960 4 vdd
rlabel metal3 s 317 39214 415 39312 4 gnd
rlabel metal3 s 17237 51862 17335 51960 4 vdd
rlabel metal3 s 15989 51862 16087 51960 4 vdd
rlabel metal3 s 16613 51862 16711 51960 4 vdd
rlabel metal3 s 317 45218 415 45316 4 gnd
rlabel metal3 s 9749 51862 9847 51960 4 vdd
rlabel metal3 s 7253 51862 7351 51960 4 vdd
rlabel metal3 s 317 46324 415 46422 4 gnd
rlabel metal3 s 317 40478 415 40576 4 gnd
rlabel metal3 s 317 41821 415 41919 4 gnd
rlabel metal3 s 317 43954 415 44052 4 gnd
rlabel metal3 s 317 49168 415 49266 4 gnd
rlabel metal3 s 12245 51862 12343 51960 4 vdd
rlabel metal3 s 317 44981 415 45079 4 gnd
rlabel metal3 s 317 49721 415 49819 4 gnd
rlabel metal3 s 317 47351 415 47449 4 gnd
rlabel metal3 s 317 41268 415 41366 4 gnd
rlabel metal3 s 317 48141 415 48239 4 gnd
rlabel metal3 s 317 41031 415 41129 4 gnd
rlabel metal3 s 317 49958 415 50056 4 gnd
rlabel metal3 s 17861 51862 17959 51960 4 vdd
rlabel metal3 s 317 44744 415 44842 4 gnd
rlabel metal3 s 20357 51862 20455 51960 4 vdd
rlabel metal3 s 2885 51862 2983 51960 4 vdd
rlabel metal3 s 317 39688 415 39786 4 gnd
rlabel metal3 s 5381 51862 5479 51960 4 vdd
rlabel metal3 s 317 51064 415 51162 4 gnd
rlabel metal3 s 317 42058 415 42156 4 gnd
rlabel metal3 s 317 48931 415 49029 4 gnd
rlabel metal3 s 317 45534 415 45632 4 gnd
rlabel metal3 s 317 46008 415 46106 4 gnd
rlabel metal3 s 317 47904 415 48002 4 gnd
rlabel metal3 s 317 51301 415 51399 4 gnd
rlabel metal3 s 10373 51862 10471 51960 4 vdd
rlabel metal3 s 317 40241 415 40339 4 gnd
rlabel metal3 s 19733 51862 19831 51960 4 vdd
rlabel metal3 s 6005 51862 6103 51960 4 vdd
rlabel metal3 s 317 47114 415 47212 4 gnd
rlabel metal3 s 4133 51862 4231 51960 4 vdd
rlabel metal3 s 317 42374 415 42472 4 gnd
rlabel metal3 s 317 42848 415 42946 4 gnd
rlabel metal3 s 317 48378 415 48476 4 gnd
rlabel metal3 s 317 50274 415 50372 4 gnd
rlabel metal3 s 317 40004 415 40102 4 gnd
rlabel metal3 s 317 43401 415 43499 4 gnd
rlabel metal3 s 317 47588 415 47686 4 gnd
rlabel metal3 s 317 50748 415 50846 4 gnd
rlabel metal3 s 9125 51862 9223 51960 4 vdd
rlabel metal3 s 1013 51862 1111 51960 4 vdd
rlabel metal3 s 317 37871 415 37969 4 gnd
rlabel metal3 s 317 29971 415 30069 4 gnd
rlabel metal3 s 317 30998 415 31096 4 gnd
rlabel metal3 s 317 29734 415 29832 4 gnd
rlabel metal3 s 317 32341 415 32439 4 gnd
rlabel metal3 s 317 32894 415 32992 4 gnd
rlabel metal3 s 317 37634 415 37732 4 gnd
rlabel metal3 s 317 29181 415 29279 4 gnd
rlabel metal3 s 317 32578 415 32676 4 gnd
rlabel metal3 s 317 34474 415 34572 4 gnd
rlabel metal3 s 317 29418 415 29516 4 gnd
rlabel metal3 s 317 37081 415 37179 4 gnd
rlabel metal3 s 317 35501 415 35599 4 gnd
rlabel metal3 s 317 35738 415 35836 4 gnd
rlabel metal3 s 317 28944 415 29042 4 gnd
rlabel metal3 s 317 36528 415 36626 4 gnd
rlabel metal3 s 317 36291 415 36389 4 gnd
rlabel metal3 s 317 28391 415 28489 4 gnd
rlabel metal3 s 317 28154 415 28252 4 gnd
rlabel metal3 s 317 30524 415 30622 4 gnd
rlabel metal3 s 317 27048 415 27146 4 gnd
rlabel metal3 s 317 34711 415 34809 4 gnd
rlabel metal3 s 317 32104 415 32202 4 gnd
rlabel metal3 s 317 38898 415 38996 4 gnd
rlabel metal3 s 317 27601 415 27699 4 gnd
rlabel metal3 s 317 36054 415 36152 4 gnd
rlabel metal3 s 317 33921 415 34019 4 gnd
rlabel metal3 s 317 35264 415 35362 4 gnd
rlabel metal3 s 317 37318 415 37416 4 gnd
rlabel metal3 s 317 26258 415 26356 4 gnd
rlabel metal3 s 317 34948 415 35046 4 gnd
rlabel metal3 s 317 31551 415 31649 4 gnd
rlabel metal3 s 317 38661 415 38759 4 gnd
rlabel metal3 s 317 31314 415 31412 4 gnd
rlabel metal3 s 317 33684 415 33782 4 gnd
rlabel metal3 s 317 30208 415 30306 4 gnd
rlabel metal3 s 317 28628 415 28726 4 gnd
rlabel metal3 s 317 30761 415 30859 4 gnd
rlabel metal3 s 317 38424 415 38522 4 gnd
rlabel metal3 s 317 33131 415 33229 4 gnd
rlabel metal3 s 317 26574 415 26672 4 gnd
rlabel metal3 s 317 36844 415 36942 4 gnd
rlabel metal3 s 317 31788 415 31886 4 gnd
rlabel metal3 s 317 26811 415 26909 4 gnd
rlabel metal3 s 317 27364 415 27462 4 gnd
rlabel metal3 s 317 27838 415 27936 4 gnd
rlabel metal3 s 317 33368 415 33466 4 gnd
rlabel metal3 s 317 34158 415 34256 4 gnd
rlabel metal3 s 317 38108 415 38206 4 gnd
rlabel metal3 s 317 24204 415 24302 4 gnd
rlabel metal3 s 317 13934 415 14032 4 gnd
rlabel metal3 s 317 13144 415 13242 4 gnd
rlabel metal3 s 317 24678 415 24776 4 gnd
rlabel metal3 s 317 18911 415 19009 4 gnd
rlabel metal3 s 317 16778 415 16876 4 gnd
rlabel metal3 s 317 18121 415 18219 4 gnd
rlabel metal3 s 317 19938 415 20036 4 gnd
rlabel metal3 s 317 13381 415 13479 4 gnd
rlabel metal3 s 317 20254 415 20352 4 gnd
rlabel metal3 s 317 14961 415 15059 4 gnd
rlabel metal3 s 317 26021 415 26119 4 gnd
rlabel metal3 s 317 22071 415 22169 4 gnd
rlabel metal3 s 317 24441 415 24539 4 gnd
rlabel metal3 s 317 22308 415 22406 4 gnd
rlabel metal3 s 317 16304 415 16402 4 gnd
rlabel metal3 s 317 15514 415 15612 4 gnd
rlabel metal3 s 317 23414 415 23512 4 gnd
rlabel metal3 s 317 23888 415 23986 4 gnd
rlabel metal3 s 317 19701 415 19799 4 gnd
rlabel metal3 s 317 20491 415 20589 4 gnd
rlabel metal3 s 317 15988 415 16086 4 gnd
rlabel metal3 s 317 23098 415 23196 4 gnd
rlabel metal3 s 317 25231 415 25329 4 gnd
rlabel metal3 s 317 21834 415 21932 4 gnd
rlabel metal3 s 317 25784 415 25882 4 gnd
rlabel metal3 s 317 17331 415 17429 4 gnd
rlabel metal3 s 317 17884 415 17982 4 gnd
rlabel metal3 s 317 22861 415 22959 4 gnd
rlabel metal3 s 317 17094 415 17192 4 gnd
rlabel metal3 s 317 15198 415 15296 4 gnd
rlabel metal3 s 317 21281 415 21379 4 gnd
rlabel metal3 s 317 18358 415 18456 4 gnd
rlabel metal3 s 317 15751 415 15849 4 gnd
rlabel metal3 s 317 24994 415 25092 4 gnd
rlabel metal3 s 317 14408 415 14506 4 gnd
rlabel metal3 s 317 16541 415 16639 4 gnd
rlabel metal3 s 317 21518 415 21616 4 gnd
rlabel metal3 s 317 17568 415 17666 4 gnd
rlabel metal3 s 317 21044 415 21142 4 gnd
rlabel metal3 s 317 18674 415 18772 4 gnd
rlabel metal3 s 317 23651 415 23749 4 gnd
rlabel metal3 s 317 25468 415 25566 4 gnd
rlabel metal3 s 317 19464 415 19562 4 gnd
rlabel metal3 s 317 14724 415 14822 4 gnd
rlabel metal3 s 317 19148 415 19246 4 gnd
rlabel metal3 s 317 20728 415 20826 4 gnd
rlabel metal3 s 317 22624 415 22722 4 gnd
rlabel metal3 s 317 13618 415 13716 4 gnd
rlabel metal3 s 317 14171 415 14269 4 gnd
rlabel metal3 s 20357 180 20455 278 4 vdd
rlabel metal3 s 317 5244 415 5342 4 gnd
rlabel metal3 s 16613 180 16711 278 4 vdd
rlabel metal3 s 317 4138 415 4236 4 gnd
rlabel metal3 s 12869 180 12967 278 4 vdd
rlabel metal3 s 10997 180 11095 278 4 vdd
rlabel metal3 s 317 12591 415 12689 4 gnd
rlabel metal3 s 14117 180 14215 278 4 vdd
rlabel metal3 s 15989 180 16087 278 4 vdd
rlabel metal3 s 15365 180 15463 278 4 vdd
rlabel metal3 s 317 9431 415 9529 4 gnd
rlabel metal3 s 317 2874 415 2972 4 gnd
rlabel metal3 s 317 12038 415 12136 4 gnd
rlabel metal3 s 317 7614 415 7712 4 gnd
rlabel metal3 s 1637 180 1735 278 4 vdd
rlabel metal3 s 317 6508 415 6606 4 gnd
rlabel metal3 s 4757 180 4855 278 4 vdd
rlabel metal3 s 10373 180 10471 278 4 vdd
rlabel metal3 s 317 6034 415 6132 4 gnd
rlabel metal3 s 317 3111 415 3209 4 gnd
rlabel metal3 s 317 2084 415 2182 4 gnd
rlabel metal3 s 19109 180 19207 278 4 vdd
rlabel metal3 s 13493 180 13591 278 4 vdd
rlabel metal3 s 317 1294 415 1392 4 gnd
rlabel metal3 s 317 1768 415 1866 4 gnd
rlabel metal3 s 4133 180 4231 278 4 vdd
rlabel metal3 s 317 4454 415 4552 4 gnd
rlabel metal3 s 6005 180 6103 278 4 vdd
rlabel metal3 s 5381 180 5479 278 4 vdd
rlabel metal3 s 317 10774 415 10872 4 gnd
rlabel metal3 s 9125 180 9223 278 4 vdd
rlabel metal3 s 317 10458 415 10556 4 gnd
rlabel metal3 s 317 8878 415 8976 4 gnd
rlabel metal3 s 317 6824 415 6922 4 gnd
rlabel metal3 s 317 3901 415 3999 4 gnd
rlabel metal3 s 7877 180 7975 278 4 vdd
rlabel metal3 s 317 6271 415 6369 4 gnd
rlabel metal3 s 3509 180 3607 278 4 vdd
rlabel metal3 s 7253 180 7351 278 4 vdd
rlabel metal3 s 19733 180 19831 278 4 vdd
rlabel metal3 s 317 4691 415 4789 4 gnd
rlabel metal3 s 317 8404 415 8502 4 gnd
rlabel metal3 s 317 12828 415 12926 4 gnd
rlabel metal3 s 317 8088 415 8186 4 gnd
rlabel metal3 s 8501 180 8599 278 4 vdd
rlabel metal3 s 317 2558 415 2656 4 gnd
rlabel metal3 s 317 5718 415 5816 4 gnd
rlabel metal3 s 11621 180 11719 278 4 vdd
rlabel metal3 s 317 11248 415 11346 4 gnd
rlabel metal3 s 317 2321 415 2419 4 gnd
rlabel metal3 s 317 741 415 839 4 gnd
rlabel metal3 s 317 7298 415 7396 4 gnd
rlabel metal3 s 317 11801 415 11899 4 gnd
rlabel metal3 s 17861 180 17959 278 4 vdd
rlabel metal3 s 317 7851 415 7949 4 gnd
rlabel metal3 s 317 10221 415 10319 4 gnd
rlabel metal3 s 317 11564 415 11662 4 gnd
rlabel metal3 s 317 3664 415 3762 4 gnd
rlabel metal3 s 12245 180 12343 278 4 vdd
rlabel metal3 s 317 8641 415 8739 4 gnd
rlabel metal3 s 2885 180 2983 278 4 vdd
rlabel metal3 s 17237 180 17335 278 4 vdd
rlabel metal3 s 317 11011 415 11109 4 gnd
rlabel metal3 s 317 7061 415 7159 4 gnd
rlabel metal3 s 317 1531 415 1629 4 gnd
rlabel metal3 s 317 4928 415 5026 4 gnd
rlabel metal3 s 317 5481 415 5579 4 gnd
rlabel metal3 s 317 12354 415 12452 4 gnd
rlabel metal3 s 317 9668 415 9766 4 gnd
rlabel metal3 s 317 3348 415 3446 4 gnd
rlabel metal3 s 2261 180 2359 278 4 vdd
rlabel metal3 s 317 9984 415 10082 4 gnd
rlabel metal3 s 1013 180 1111 278 4 vdd
rlabel metal3 s 18485 180 18583 278 4 vdd
rlabel metal3 s 9749 180 9847 278 4 vdd
rlabel metal3 s 317 9194 415 9292 4 gnd
rlabel metal3 s 6629 180 6727 278 4 vdd
rlabel metal3 s -49 614 49 712 4 gnd
rlabel metal3 s 317 978 415 1076 4 gnd
rlabel metal3 s 14741 180 14839 278 4 vdd
rlabel metal3 s 23477 180 23575 278 4 vdd
rlabel metal3 s 26597 180 26695 278 4 vdd
rlabel metal3 s 20981 180 21079 278 4 vdd
rlabel metal3 s 37205 180 37303 278 4 vdd
rlabel metal3 s 40949 180 41047 278 4 vdd
rlabel metal3 s 27221 180 27319 278 4 vdd
rlabel metal3 s 35957 180 36055 278 4 vdd
rlabel metal3 s 34085 180 34183 278 4 vdd
rlabel metal3 s 39701 180 39799 278 4 vdd
rlabel metal3 s 30341 180 30439 278 4 vdd
rlabel metal3 s 29717 180 29815 278 4 vdd
rlabel metal3 s 30965 180 31063 278 4 vdd
rlabel metal3 s 37829 180 37927 278 4 vdd
rlabel metal3 s 24725 180 24823 278 4 vdd
rlabel metal3 s 31589 180 31687 278 4 vdd
rlabel metal3 s 21605 180 21703 278 4 vdd
rlabel metal3 s 22229 180 22327 278 4 vdd
rlabel metal3 s 25973 180 26071 278 4 vdd
rlabel metal3 s 35333 180 35431 278 4 vdd
rlabel metal3 s 38453 180 38551 278 4 vdd
rlabel metal3 s 36581 180 36679 278 4 vdd
rlabel metal3 s 29093 180 29191 278 4 vdd
rlabel metal3 s 27845 180 27943 278 4 vdd
rlabel metal3 s 33461 180 33559 278 4 vdd
rlabel metal3 s 25349 180 25447 278 4 vdd
rlabel metal3 s 32837 180 32935 278 4 vdd
rlabel metal3 s 34709 180 34807 278 4 vdd
rlabel metal3 s 40325 180 40423 278 4 vdd
rlabel metal3 s 24101 180 24199 278 4 vdd
rlabel metal3 s 39077 180 39175 278 4 vdd
rlabel metal3 s 32213 180 32311 278 4 vdd
rlabel metal3 s 28469 180 28567 278 4 vdd
rlabel metal3 s 22853 180 22951 278 4 vdd
rlabel metal3 s 82205 14961 82303 15059 4 gnd
rlabel metal3 s 82205 13144 82303 13242 4 gnd
rlabel metal3 s 82205 23414 82303 23512 4 gnd
rlabel metal3 s 82205 13934 82303 14032 4 gnd
rlabel metal3 s 82205 19701 82303 19799 4 gnd
rlabel metal3 s 82205 15198 82303 15296 4 gnd
rlabel metal3 s 82205 15751 82303 15849 4 gnd
rlabel metal3 s 82205 14171 82303 14269 4 gnd
rlabel metal3 s 82205 24204 82303 24302 4 gnd
rlabel metal3 s 82205 22308 82303 22406 4 gnd
rlabel metal3 s 82205 18358 82303 18456 4 gnd
rlabel metal3 s 82205 16778 82303 16876 4 gnd
rlabel metal3 s 82205 13381 82303 13479 4 gnd
rlabel metal3 s 82205 21044 82303 21142 4 gnd
rlabel metal3 s 82205 18911 82303 19009 4 gnd
rlabel metal3 s 82205 25784 82303 25882 4 gnd
rlabel metal3 s 82205 14724 82303 14822 4 gnd
rlabel metal3 s 82205 17568 82303 17666 4 gnd
rlabel metal3 s 82205 23651 82303 23749 4 gnd
rlabel metal3 s 82205 15514 82303 15612 4 gnd
rlabel metal3 s 82205 23888 82303 23986 4 gnd
rlabel metal3 s 82205 16541 82303 16639 4 gnd
rlabel metal3 s 82205 21834 82303 21932 4 gnd
rlabel metal3 s 82205 17884 82303 17982 4 gnd
rlabel metal3 s 82205 17331 82303 17429 4 gnd
rlabel metal3 s 82205 21281 82303 21379 4 gnd
rlabel metal3 s 82205 24441 82303 24539 4 gnd
rlabel metal3 s 82205 20254 82303 20352 4 gnd
rlabel metal3 s 82205 24678 82303 24776 4 gnd
rlabel metal3 s 82205 18121 82303 18219 4 gnd
rlabel metal3 s 82205 22861 82303 22959 4 gnd
rlabel metal3 s 82205 14408 82303 14506 4 gnd
rlabel metal3 s 82205 20728 82303 20826 4 gnd
rlabel metal3 s 82205 13618 82303 13716 4 gnd
rlabel metal3 s 82205 21518 82303 21616 4 gnd
rlabel metal3 s 82205 20491 82303 20589 4 gnd
rlabel metal3 s 82205 15988 82303 16086 4 gnd
rlabel metal3 s 82205 16304 82303 16402 4 gnd
rlabel metal3 s 82205 24994 82303 25092 4 gnd
rlabel metal3 s 82205 25468 82303 25566 4 gnd
rlabel metal3 s 82205 17094 82303 17192 4 gnd
rlabel metal3 s 82205 26021 82303 26119 4 gnd
rlabel metal3 s 82205 18674 82303 18772 4 gnd
rlabel metal3 s 82205 22071 82303 22169 4 gnd
rlabel metal3 s 82205 19148 82303 19246 4 gnd
rlabel metal3 s 82205 25231 82303 25329 4 gnd
rlabel metal3 s 82205 23098 82303 23196 4 gnd
rlabel metal3 s 82205 19464 82303 19562 4 gnd
rlabel metal3 s 82205 19938 82303 20036 4 gnd
rlabel metal3 s 82205 22624 82303 22722 4 gnd
rlabel metal3 s 52805 180 52903 278 4 vdd
rlabel metal3 s 54053 180 54151 278 4 vdd
rlabel metal3 s 45317 180 45415 278 4 vdd
rlabel metal3 s 57797 180 57895 278 4 vdd
rlabel metal3 s 50933 180 51031 278 4 vdd
rlabel metal3 s 59669 180 59767 278 4 vdd
rlabel metal3 s 44693 180 44791 278 4 vdd
rlabel metal3 s 55301 180 55399 278 4 vdd
rlabel metal3 s 60917 180 61015 278 4 vdd
rlabel metal3 s 53429 180 53527 278 4 vdd
rlabel metal3 s 49685 180 49783 278 4 vdd
rlabel metal3 s 46565 180 46663 278 4 vdd
rlabel metal3 s 56549 180 56647 278 4 vdd
rlabel metal3 s 50309 180 50407 278 4 vdd
rlabel metal3 s 58421 180 58519 278 4 vdd
rlabel metal3 s 47189 180 47287 278 4 vdd
rlabel metal3 s 61541 180 61639 278 4 vdd
rlabel metal3 s 54677 180 54775 278 4 vdd
rlabel metal3 s 59045 180 59143 278 4 vdd
rlabel metal3 s 45941 180 46039 278 4 vdd
rlabel metal3 s 55925 180 56023 278 4 vdd
rlabel metal3 s 44069 180 44167 278 4 vdd
rlabel metal3 s 51557 180 51655 278 4 vdd
rlabel metal3 s 48437 180 48535 278 4 vdd
rlabel metal3 s 43445 180 43543 278 4 vdd
rlabel metal3 s 41573 180 41671 278 4 vdd
rlabel metal3 s 52181 180 52279 278 4 vdd
rlabel metal3 s 57173 180 57271 278 4 vdd
rlabel metal3 s 42197 180 42295 278 4 vdd
rlabel metal3 s 47813 180 47911 278 4 vdd
rlabel metal3 s 42821 180 42919 278 4 vdd
rlabel metal3 s 49061 180 49159 278 4 vdd
rlabel metal3 s 60293 180 60391 278 4 vdd
rlabel metal3 s 82205 10221 82303 10319 4 gnd
rlabel metal3 s 82205 7614 82303 7712 4 gnd
rlabel metal3 s 72773 180 72871 278 4 vdd
rlabel metal3 s 77141 180 77239 278 4 vdd
rlabel metal3 s 66533 180 66631 278 4 vdd
rlabel metal3 s 82205 2321 82303 2419 4 gnd
rlabel metal3 s 65285 180 65383 278 4 vdd
rlabel metal3 s 68405 180 68503 278 4 vdd
rlabel metal3 s 80261 180 80359 278 4 vdd
rlabel metal3 s 82205 7061 82303 7159 4 gnd
rlabel metal3 s 82205 6508 82303 6606 4 gnd
rlabel metal3 s 65909 180 66007 278 4 vdd
rlabel metal3 s 75893 180 75991 278 4 vdd
rlabel metal3 s 67157 180 67255 278 4 vdd
rlabel metal3 s 72149 180 72247 278 4 vdd
rlabel metal3 s 82205 1531 82303 1629 4 gnd
rlabel metal3 s 73397 180 73495 278 4 vdd
rlabel metal3 s 82205 1768 82303 1866 4 gnd
rlabel metal3 s 82205 11564 82303 11662 4 gnd
rlabel metal3 s 82571 614 82669 712 4 gnd
rlabel metal3 s 82205 9668 82303 9766 4 gnd
rlabel metal3 s 82205 6034 82303 6132 4 gnd
rlabel metal3 s 82205 9194 82303 9292 4 gnd
rlabel metal3 s 67781 180 67879 278 4 vdd
rlabel metal3 s 82205 2874 82303 2972 4 gnd
rlabel metal3 s 81509 180 81607 278 4 vdd
rlabel metal3 s 82205 7298 82303 7396 4 gnd
rlabel metal3 s 82205 8088 82303 8186 4 gnd
rlabel metal3 s 82205 12354 82303 12452 4 gnd
rlabel metal3 s 70277 180 70375 278 4 vdd
rlabel metal3 s 82205 4454 82303 4552 4 gnd
rlabel metal3 s 78389 180 78487 278 4 vdd
rlabel metal3 s 69029 180 69127 278 4 vdd
rlabel metal3 s 82205 9431 82303 9529 4 gnd
rlabel metal3 s 64037 180 64135 278 4 vdd
rlabel metal3 s 82205 3664 82303 3762 4 gnd
rlabel metal3 s 80885 180 80983 278 4 vdd
rlabel metal3 s 82205 3111 82303 3209 4 gnd
rlabel metal3 s 82205 10774 82303 10872 4 gnd
rlabel metal3 s 82205 9984 82303 10082 4 gnd
rlabel metal3 s 82205 5244 82303 5342 4 gnd
rlabel metal3 s 82205 741 82303 839 4 gnd
rlabel metal3 s 62789 180 62887 278 4 vdd
rlabel metal3 s 82205 978 82303 1076 4 gnd
rlabel metal3 s 69653 180 69751 278 4 vdd
rlabel metal3 s 70901 180 70999 278 4 vdd
rlabel metal3 s 82205 6824 82303 6922 4 gnd
rlabel metal3 s 82205 12591 82303 12689 4 gnd
rlabel metal3 s 62165 180 62263 278 4 vdd
rlabel metal3 s 82205 7851 82303 7949 4 gnd
rlabel metal3 s 71525 180 71623 278 4 vdd
rlabel metal3 s 82205 10458 82303 10556 4 gnd
rlabel metal3 s 82205 6271 82303 6369 4 gnd
rlabel metal3 s 79637 180 79735 278 4 vdd
rlabel metal3 s 82205 12828 82303 12926 4 gnd
rlabel metal3 s 82205 2084 82303 2182 4 gnd
rlabel metal3 s 82205 3901 82303 3999 4 gnd
rlabel metal3 s 82205 4928 82303 5026 4 gnd
rlabel metal3 s 82205 4138 82303 4236 4 gnd
rlabel metal3 s 82205 5718 82303 5816 4 gnd
rlabel metal3 s 82205 2558 82303 2656 4 gnd
rlabel metal3 s 82205 3348 82303 3446 4 gnd
rlabel metal3 s 75269 180 75367 278 4 vdd
rlabel metal3 s 63413 180 63511 278 4 vdd
rlabel metal3 s 74021 180 74119 278 4 vdd
rlabel metal3 s 82205 4691 82303 4789 4 gnd
rlabel metal3 s 82205 12038 82303 12136 4 gnd
rlabel metal3 s 76517 180 76615 278 4 vdd
rlabel metal3 s 82205 5481 82303 5579 4 gnd
rlabel metal3 s 82205 1294 82303 1392 4 gnd
rlabel metal3 s 82205 8641 82303 8739 4 gnd
rlabel metal3 s 82205 11801 82303 11899 4 gnd
rlabel metal3 s 79013 180 79111 278 4 vdd
rlabel metal3 s 82205 8404 82303 8502 4 gnd
rlabel metal3 s 64661 180 64759 278 4 vdd
rlabel metal3 s 82205 11248 82303 11346 4 gnd
rlabel metal3 s 82205 8878 82303 8976 4 gnd
rlabel metal3 s 77765 180 77863 278 4 vdd
rlabel metal3 s 74645 180 74743 278 4 vdd
rlabel metal3 s 82205 11011 82303 11109 4 gnd
rlabel metal2 s 81432 31009 81540 31085 4 gnd
rlabel metal2 s 81432 42069 81540 42145 4 gnd
rlabel metal2 s 81432 34705 81540 34815 4 gnd
rlabel metal2 s 81432 51295 81540 51405 4 gnd
rlabel metal2 s 81432 42385 81540 42461 4 gnd
rlabel metal2 s 81432 48389 81540 48465 4 gnd
rlabel metal2 s 81432 27849 81540 27925 4 gnd
rlabel metal2 s 81432 29429 81540 29505 4 gnd
rlabel metal2 s 81432 30535 81540 30611 4 gnd
rlabel metal2 s 81432 43649 81540 43725 4 gnd
rlabel metal2 s 81432 48705 81540 48781 4 gnd
rlabel metal2 s 81432 29175 81540 29285 4 gnd
rlabel metal2 s 81432 46019 81540 46095 4 gnd
rlabel metal2 s 81432 48925 81540 49035 4 gnd
rlabel metal2 s 81432 44185 81540 44295 4 gnd
rlabel metal2 s 81432 28639 81540 28715 4 gnd
rlabel metal2 s 81432 30219 81540 30295 4 gnd
rlabel metal2 s 81432 34169 81540 34245 4 gnd
rlabel metal2 s 81432 27059 81540 27135 4 gnd
rlabel metal2 s 81432 32115 81540 32191 4 gnd
rlabel metal2 s 81432 42859 81540 42935 4 gnd
rlabel metal2 s 81432 41595 81540 41671 4 gnd
rlabel metal2 s 81432 50505 81540 50615 4 gnd
rlabel metal2 s 81432 45545 81540 45621 4 gnd
rlabel metal2 s 81432 49969 81540 50045 4 gnd
rlabel metal2 s 81432 44755 81540 44831 4 gnd
rlabel metal2 s 81432 28385 81540 28495 4 gnd
rlabel metal2 s 81432 46809 81540 46885 4 gnd
rlabel metal2 s 81432 27595 81540 27705 4 gnd
rlabel metal2 s 81432 45229 81540 45305 4 gnd
rlabel metal2 s 81432 40015 81540 40091 4 gnd
rlabel metal2 s 81432 33379 81540 33455 4 gnd
rlabel metal2 s 81432 40235 81540 40345 4 gnd
rlabel metal2 s 81432 43175 81540 43251 4 gnd
rlabel metal2 s 81432 33125 81540 33235 4 gnd
rlabel metal2 s 81432 43395 81540 43505 4 gnd
rlabel metal2 s 81432 36539 81540 36615 4 gnd
rlabel metal2 s 81432 31545 81540 31655 4 gnd
rlabel metal2 s 81432 50759 81540 50835 4 gnd
rlabel metal2 s 81432 47345 81540 47455 4 gnd
rlabel metal2 s 81432 39225 81540 39301 4 gnd
rlabel metal2 s 81432 48135 81540 48245 4 gnd
rlabel metal2 s 81432 41815 81540 41925 4 gnd
rlabel metal2 s 81432 36285 81540 36395 4 gnd
rlabel metal2 s 81432 34959 81540 35035 4 gnd
rlabel metal2 s 81432 39699 81540 39775 4 gnd
rlabel metal2 s 81432 26805 81540 26915 4 gnd
rlabel metal2 s 81432 49179 81540 49255 4 gnd
rlabel metal2 s 81432 32335 81540 32445 4 gnd
rlabel metal2 s 81432 38655 81540 38765 4 gnd
rlabel metal2 s 81432 47599 81540 47675 4 gnd
rlabel metal2 s 81432 44975 81540 45085 4 gnd
rlabel metal2 s 81432 32905 81540 32981 4 gnd
rlabel metal2 s 81432 47125 81540 47201 4 gnd
rlabel metal2 s 81432 38119 81540 38195 4 gnd
rlabel metal2 s 81432 35495 81540 35605 4 gnd
rlabel metal2 s 81432 29965 81540 30075 4 gnd
rlabel metal2 s 81432 40805 81540 40881 4 gnd
rlabel metal2 s 81432 35275 81540 35351 4 gnd
rlabel metal2 s 81432 46555 81540 46665 4 gnd
rlabel metal2 s 81432 33695 81540 33771 4 gnd
rlabel metal2 s 81432 50285 81540 50361 4 gnd
rlabel metal2 s 81432 45765 81540 45875 4 gnd
rlabel metal2 s 81432 51549 81540 51625 4 gnd
rlabel metal2 s 81432 31325 81540 31401 4 gnd
rlabel metal2 s 81432 41025 81540 41135 4 gnd
rlabel metal2 s 81432 31799 81540 31875 4 gnd
rlabel metal2 s 81432 38435 81540 38511 4 gnd
rlabel metal2 s 81432 33915 81540 34025 4 gnd
rlabel metal2 s 81432 47915 81540 47991 4 gnd
rlabel metal2 s 81432 49495 81540 49571 4 gnd
rlabel metal2 s 81432 28165 81540 28241 4 gnd
rlabel metal2 s 81432 37329 81540 37405 4 gnd
rlabel metal2 s 81432 26585 81540 26661 4 gnd
rlabel metal2 s 81432 43965 81540 44041 4 gnd
rlabel metal2 s 81432 44439 81540 44515 4 gnd
rlabel metal2 s 81432 46335 81540 46411 4 gnd
rlabel metal2 s 81432 41279 81540 41355 4 gnd
rlabel metal2 s 81432 32589 81540 32665 4 gnd
rlabel metal2 s 81432 37075 81540 37185 4 gnd
rlabel metal2 s 81432 28955 81540 29031 4 gnd
rlabel metal2 s 81432 35749 81540 35825 4 gnd
rlabel metal2 s 81432 38909 81540 38985 4 gnd
rlabel metal2 s 81432 40489 81540 40565 4 gnd
rlabel metal2 s 81432 36065 81540 36141 4 gnd
rlabel metal2 s 81432 42605 81540 42715 4 gnd
rlabel metal2 s 81432 29745 81540 29821 4 gnd
rlabel metal2 s 81432 49715 81540 49825 4 gnd
rlabel metal2 s 81432 39445 81540 39555 4 gnd
rlabel metal2 s 81432 37865 81540 37975 4 gnd
rlabel metal2 s 81432 26269 81540 26345 4 gnd
rlabel metal2 s 81432 27375 81540 27451 4 gnd
rlabel metal2 s 81432 34485 81540 34561 4 gnd
rlabel metal2 s 81432 51075 81540 51151 4 gnd
rlabel metal2 s 81432 37645 81540 37721 4 gnd
rlabel metal2 s 81432 36855 81540 36931 4 gnd
rlabel metal2 s 81432 30755 81540 30865 4 gnd
rlabel metal2 s 81432 26015 81540 26125 4 gnd
rlabel metal2 s 0 45449 82620 45497 4 wl_0_113
rlabel metal2 s 0 45669 82620 45717 4 wl_1_113
rlabel metal2 s 0 46143 82620 46191 4 wl_0_114
rlabel metal2 s 0 45923 82620 45971 4 wl_1_114
rlabel metal2 s 0 46239 82620 46287 4 wl_0_115
rlabel metal2 s 0 46459 82620 46507 4 wl_1_115
rlabel metal2 s 0 46933 82620 46981 4 wl_0_116
rlabel metal2 s 0 46713 82620 46761 4 wl_1_116
rlabel metal2 s 0 47029 82620 47077 4 wl_0_117
rlabel metal2 s 0 47249 82620 47297 4 wl_1_117
rlabel metal2 s 0 47723 82620 47771 4 wl_0_118
rlabel metal2 s 0 47503 82620 47551 4 wl_1_118
rlabel metal2 s 0 47819 82620 47867 4 wl_0_119
rlabel metal2 s 0 48039 82620 48087 4 wl_1_119
rlabel metal2 s 0 48513 82620 48561 4 wl_0_120
rlabel metal2 s 0 48293 82620 48341 4 wl_1_120
rlabel metal2 s 0 48609 82620 48657 4 wl_0_121
rlabel metal2 s 0 48829 82620 48877 4 wl_1_121
rlabel metal2 s 0 49303 82620 49351 4 wl_0_122
rlabel metal2 s 0 49083 82620 49131 4 wl_1_122
rlabel metal2 s 0 49399 82620 49447 4 wl_0_123
rlabel metal2 s 0 49619 82620 49667 4 wl_1_123
rlabel metal2 s 0 50093 82620 50141 4 wl_0_124
rlabel metal2 s 0 49873 82620 49921 4 wl_1_124
rlabel metal2 s 0 50189 82620 50237 4 wl_0_125
rlabel metal2 s 0 50409 82620 50457 4 wl_1_125
rlabel metal2 s 0 50883 82620 50931 4 wl_0_126
rlabel metal2 s 0 50663 82620 50711 4 wl_1_126
rlabel metal2 s 0 50979 82620 51027 4 wl_0_127
rlabel metal2 s 0 51199 82620 51247 4 wl_1_127
rlabel metal2 s 0 51453 82620 51501 4 rbl_wl_1_1
rlabel metal2 s 0 39033 82620 39081 4 wl_0_96
rlabel metal2 s 0 38813 82620 38861 4 wl_1_96
rlabel metal2 s 0 39129 82620 39177 4 wl_0_97
rlabel metal2 s 0 39349 82620 39397 4 wl_1_97
rlabel metal2 s 0 39823 82620 39871 4 wl_0_98
rlabel metal2 s 0 39603 82620 39651 4 wl_1_98
rlabel metal2 s 0 39919 82620 39967 4 wl_0_99
rlabel metal2 s 0 40139 82620 40187 4 wl_1_99
rlabel metal2 s 0 40613 82620 40661 4 wl_0_100
rlabel metal2 s 0 40393 82620 40441 4 wl_1_100
rlabel metal2 s 0 40709 82620 40757 4 wl_0_101
rlabel metal2 s 0 40929 82620 40977 4 wl_1_101
rlabel metal2 s 0 41403 82620 41451 4 wl_0_102
rlabel metal2 s 0 41183 82620 41231 4 wl_1_102
rlabel metal2 s 0 41499 82620 41547 4 wl_0_103
rlabel metal2 s 0 41719 82620 41767 4 wl_1_103
rlabel metal2 s 0 42193 82620 42241 4 wl_0_104
rlabel metal2 s 0 41973 82620 42021 4 wl_1_104
rlabel metal2 s 0 42289 82620 42337 4 wl_0_105
rlabel metal2 s 0 42509 82620 42557 4 wl_1_105
rlabel metal2 s 0 42983 82620 43031 4 wl_0_106
rlabel metal2 s 0 42763 82620 42811 4 wl_1_106
rlabel metal2 s 0 43079 82620 43127 4 wl_0_107
rlabel metal2 s 0 43299 82620 43347 4 wl_1_107
rlabel metal2 s 0 43773 82620 43821 4 wl_0_108
rlabel metal2 s 0 43553 82620 43601 4 wl_1_108
rlabel metal2 s 0 43869 82620 43917 4 wl_0_109
rlabel metal2 s 0 44089 82620 44137 4 wl_1_109
rlabel metal2 s 0 44563 82620 44611 4 wl_0_110
rlabel metal2 s 0 44343 82620 44391 4 wl_1_110
rlabel metal2 s 0 44659 82620 44707 4 wl_0_111
rlabel metal2 s 0 44879 82620 44927 4 wl_1_111
rlabel metal2 s 0 45353 82620 45401 4 wl_0_112
rlabel metal2 s 0 45133 82620 45181 4 wl_1_112
rlabel metal2 s 1080 41595 1188 41671 4 gnd
rlabel metal2 s 1080 43175 1188 43251 4 gnd
rlabel metal2 s 1080 39445 1188 39555 4 gnd
rlabel metal2 s 1080 49969 1188 50045 4 gnd
rlabel metal2 s 1080 49179 1188 49255 4 gnd
rlabel metal2 s 1080 48389 1188 48465 4 gnd
rlabel metal2 s 1080 44975 1188 45085 4 gnd
rlabel metal2 s 1080 47125 1188 47201 4 gnd
rlabel metal2 s 1080 45545 1188 45621 4 gnd
rlabel metal2 s 1080 44755 1188 44831 4 gnd
rlabel metal2 s 1080 46809 1188 46885 4 gnd
rlabel metal2 s 1080 38909 1188 38985 4 gnd
rlabel metal2 s 1080 41815 1188 41925 4 gnd
rlabel metal2 s 1080 48925 1188 49035 4 gnd
rlabel metal2 s 1080 46555 1188 46665 4 gnd
rlabel metal2 s 1080 50759 1188 50835 4 gnd
rlabel metal2 s 1080 44185 1188 44295 4 gnd
rlabel metal2 s 1080 39225 1188 39301 4 gnd
rlabel metal2 s 1080 43649 1188 43725 4 gnd
rlabel metal2 s 1080 46019 1188 46095 4 gnd
rlabel metal2 s 1080 49495 1188 49571 4 gnd
rlabel metal2 s 1080 47915 1188 47991 4 gnd
rlabel metal2 s 1080 40805 1188 40881 4 gnd
rlabel metal2 s 1080 44439 1188 44515 4 gnd
rlabel metal2 s 1080 51075 1188 51151 4 gnd
rlabel metal2 s 1080 45765 1188 45875 4 gnd
rlabel metal2 s 1080 48705 1188 48781 4 gnd
rlabel metal2 s 1080 40489 1188 40565 4 gnd
rlabel metal2 s 1080 43395 1188 43505 4 gnd
rlabel metal2 s 1080 42069 1188 42145 4 gnd
rlabel metal2 s 1080 45229 1188 45305 4 gnd
rlabel metal2 s 1080 42385 1188 42461 4 gnd
rlabel metal2 s 1080 41279 1188 41355 4 gnd
rlabel metal2 s 1080 46335 1188 46411 4 gnd
rlabel metal2 s 1080 40235 1188 40345 4 gnd
rlabel metal2 s 1080 42605 1188 42715 4 gnd
rlabel metal2 s 1080 51295 1188 51405 4 gnd
rlabel metal2 s 1080 43965 1188 44041 4 gnd
rlabel metal2 s 1080 40015 1188 40091 4 gnd
rlabel metal2 s 1080 50285 1188 50361 4 gnd
rlabel metal2 s 1080 39699 1188 39775 4 gnd
rlabel metal2 s 1080 48135 1188 48245 4 gnd
rlabel metal2 s 1080 41025 1188 41135 4 gnd
rlabel metal2 s 1080 50505 1188 50615 4 gnd
rlabel metal2 s 1080 51549 1188 51625 4 gnd
rlabel metal2 s 1080 47599 1188 47675 4 gnd
rlabel metal2 s 1080 49715 1188 49825 4 gnd
rlabel metal2 s 1080 42859 1188 42935 4 gnd
rlabel metal2 s 1080 47345 1188 47455 4 gnd
rlabel metal2 s 1080 32115 1188 32191 4 gnd
rlabel metal2 s 1080 38435 1188 38511 4 gnd
rlabel metal2 s 1080 35749 1188 35825 4 gnd
rlabel metal2 s 1080 26015 1188 26125 4 gnd
rlabel metal2 s 1080 27595 1188 27705 4 gnd
rlabel metal2 s 1080 36285 1188 36395 4 gnd
rlabel metal2 s 1080 36065 1188 36141 4 gnd
rlabel metal2 s 1080 26805 1188 26915 4 gnd
rlabel metal2 s 1080 34485 1188 34561 4 gnd
rlabel metal2 s 1080 33125 1188 33235 4 gnd
rlabel metal2 s 1080 33915 1188 34025 4 gnd
rlabel metal2 s 1080 31799 1188 31875 4 gnd
rlabel metal2 s 1080 33379 1188 33455 4 gnd
rlabel metal2 s 1080 35275 1188 35351 4 gnd
rlabel metal2 s 1080 28165 1188 28241 4 gnd
rlabel metal2 s 1080 30535 1188 30611 4 gnd
rlabel metal2 s 1080 31009 1188 31085 4 gnd
rlabel metal2 s 1080 26269 1188 26345 4 gnd
rlabel metal2 s 1080 29429 1188 29505 4 gnd
rlabel metal2 s 1080 38655 1188 38765 4 gnd
rlabel metal2 s 1080 28385 1188 28495 4 gnd
rlabel metal2 s 1080 31545 1188 31655 4 gnd
rlabel metal2 s 1080 36855 1188 36931 4 gnd
rlabel metal2 s 1080 32335 1188 32445 4 gnd
rlabel metal2 s 1080 26585 1188 26661 4 gnd
rlabel metal2 s 1080 27059 1188 27135 4 gnd
rlabel metal2 s 1080 30755 1188 30865 4 gnd
rlabel metal2 s 1080 29175 1188 29285 4 gnd
rlabel metal2 s 1080 38119 1188 38195 4 gnd
rlabel metal2 s 1080 28639 1188 28715 4 gnd
rlabel metal2 s 1080 34959 1188 35035 4 gnd
rlabel metal2 s 1080 36539 1188 36615 4 gnd
rlabel metal2 s 1080 35495 1188 35605 4 gnd
rlabel metal2 s 1080 33695 1188 33771 4 gnd
rlabel metal2 s 1080 31325 1188 31401 4 gnd
rlabel metal2 s 1080 37075 1188 37185 4 gnd
rlabel metal2 s 1080 37329 1188 37405 4 gnd
rlabel metal2 s 1080 32905 1188 32981 4 gnd
rlabel metal2 s 1080 34169 1188 34245 4 gnd
rlabel metal2 s 1080 37865 1188 37975 4 gnd
rlabel metal2 s 1080 30219 1188 30295 4 gnd
rlabel metal2 s 1080 29965 1188 30075 4 gnd
rlabel metal2 s 1080 28955 1188 29031 4 gnd
rlabel metal2 s 1080 37645 1188 37721 4 gnd
rlabel metal2 s 1080 34705 1188 34815 4 gnd
rlabel metal2 s 1080 27849 1188 27925 4 gnd
rlabel metal2 s 1080 32589 1188 32665 4 gnd
rlabel metal2 s 1080 29745 1188 29821 4 gnd
rlabel metal2 s 1080 27375 1188 27451 4 gnd
rlabel metal2 s 0 32809 82620 32857 4 wl_0_81
rlabel metal2 s 0 27499 82620 27547 4 wl_1_67
rlabel metal2 s 0 33029 82620 33077 4 wl_1_81
rlabel metal2 s 0 33503 82620 33551 4 wl_0_82
rlabel metal2 s 0 33283 82620 33331 4 wl_1_82
rlabel metal2 s 0 33599 82620 33647 4 wl_0_83
rlabel metal2 s 0 27973 82620 28021 4 wl_0_68
rlabel metal2 s 0 26173 82620 26221 4 wl_1_64
rlabel metal2 s 0 33819 82620 33867 4 wl_1_83
rlabel metal2 s 0 34293 82620 34341 4 wl_0_84
rlabel metal2 s 0 34073 82620 34121 4 wl_1_84
rlabel metal2 s 0 34389 82620 34437 4 wl_0_85
rlabel metal2 s 0 34609 82620 34657 4 wl_1_85
rlabel metal2 s 0 35083 82620 35131 4 wl_0_86
rlabel metal2 s 0 27753 82620 27801 4 wl_1_68
rlabel metal2 s 0 28069 82620 28117 4 wl_0_69
rlabel metal2 s 0 34863 82620 34911 4 wl_1_86
rlabel metal2 s 0 35179 82620 35227 4 wl_0_87
rlabel metal2 s 0 26709 82620 26757 4 wl_1_65
rlabel metal2 s 0 35399 82620 35447 4 wl_1_87
rlabel metal2 s 0 28289 82620 28337 4 wl_1_69
rlabel metal2 s 0 35873 82620 35921 4 wl_0_88
rlabel metal2 s 0 28763 82620 28811 4 wl_0_70
rlabel metal2 s 0 35653 82620 35701 4 wl_1_88
rlabel metal2 s 0 28543 82620 28591 4 wl_1_70
rlabel metal2 s 0 35969 82620 36017 4 wl_0_89
rlabel metal2 s 0 36189 82620 36237 4 wl_1_89
rlabel metal2 s 0 30123 82620 30171 4 wl_1_74
rlabel metal2 s 0 36663 82620 36711 4 wl_0_90
rlabel metal2 s 0 30439 82620 30487 4 wl_0_75
rlabel metal2 s 0 36443 82620 36491 4 wl_1_90
rlabel metal2 s 0 36759 82620 36807 4 wl_0_91
rlabel metal2 s 0 36979 82620 37027 4 wl_1_91
rlabel metal2 s 0 26489 82620 26537 4 wl_0_65
rlabel metal2 s 0 37453 82620 37501 4 wl_0_92
rlabel metal2 s 0 30659 82620 30707 4 wl_1_75
rlabel metal2 s 0 31133 82620 31181 4 wl_0_76
rlabel metal2 s 0 37233 82620 37281 4 wl_1_92
rlabel metal2 s 0 37549 82620 37597 4 wl_0_93
rlabel metal2 s 0 37769 82620 37817 4 wl_1_93
rlabel metal2 s 0 30913 82620 30961 4 wl_1_76
rlabel metal2 s 0 38243 82620 38291 4 wl_0_94
rlabel metal2 s 0 31229 82620 31277 4 wl_0_77
rlabel metal2 s 0 38023 82620 38071 4 wl_1_94
rlabel metal2 s 0 28859 82620 28907 4 wl_0_71
rlabel metal2 s 0 27183 82620 27231 4 wl_0_66
rlabel metal2 s 0 38339 82620 38387 4 wl_0_95
rlabel metal2 s 0 29079 82620 29127 4 wl_1_71
rlabel metal2 s 0 38559 82620 38607 4 wl_1_95
rlabel metal2 s 0 29553 82620 29601 4 wl_0_72
rlabel metal2 s 0 31449 82620 31497 4 wl_1_77
rlabel metal2 s 0 31923 82620 31971 4 wl_0_78
rlabel metal2 s 0 31703 82620 31751 4 wl_1_78
rlabel metal2 s 0 32019 82620 32067 4 wl_0_79
rlabel metal2 s 0 29333 82620 29381 4 wl_1_72
rlabel metal2 s 0 29649 82620 29697 4 wl_0_73
rlabel metal2 s 0 29869 82620 29917 4 wl_1_73
rlabel metal2 s 0 30343 82620 30391 4 wl_0_74
rlabel metal2 s 0 26963 82620 27011 4 wl_1_66
rlabel metal2 s 0 26393 82620 26441 4 wl_0_64
rlabel metal2 s 0 27279 82620 27327 4 wl_0_67
rlabel metal2 s 0 32239 82620 32287 4 wl_1_79
rlabel metal2 s 0 32713 82620 32761 4 wl_0_80
rlabel metal2 s 0 32493 82620 32541 4 wl_1_80
rlabel metal2 s 0 13279 82620 13327 4 wl_1_31
rlabel metal2 s 0 13753 82620 13801 4 wl_0_32
rlabel metal2 s 0 13533 82620 13581 4 wl_1_32
rlabel metal2 s 0 13849 82620 13897 4 wl_0_33
rlabel metal2 s 0 14069 82620 14117 4 wl_1_33
rlabel metal2 s 0 14543 82620 14591 4 wl_0_34
rlabel metal2 s 0 14323 82620 14371 4 wl_1_34
rlabel metal2 s 0 14639 82620 14687 4 wl_0_35
rlabel metal2 s 0 14859 82620 14907 4 wl_1_35
rlabel metal2 s 0 15333 82620 15381 4 wl_0_36
rlabel metal2 s 0 15113 82620 15161 4 wl_1_36
rlabel metal2 s 0 15429 82620 15477 4 wl_0_37
rlabel metal2 s 0 15649 82620 15697 4 wl_1_37
rlabel metal2 s 0 16123 82620 16171 4 wl_0_38
rlabel metal2 s 0 15903 82620 15951 4 wl_1_38
rlabel metal2 s 0 16219 82620 16267 4 wl_0_39
rlabel metal2 s 0 16439 82620 16487 4 wl_1_39
rlabel metal2 s 0 16913 82620 16961 4 wl_0_40
rlabel metal2 s 0 16693 82620 16741 4 wl_1_40
rlabel metal2 s 0 17009 82620 17057 4 wl_0_41
rlabel metal2 s 0 17229 82620 17277 4 wl_1_41
rlabel metal2 s 0 17703 82620 17751 4 wl_0_42
rlabel metal2 s 0 17483 82620 17531 4 wl_1_42
rlabel metal2 s 0 17799 82620 17847 4 wl_0_43
rlabel metal2 s 0 18019 82620 18067 4 wl_1_43
rlabel metal2 s 0 18493 82620 18541 4 wl_0_44
rlabel metal2 s 0 18273 82620 18321 4 wl_1_44
rlabel metal2 s 0 18589 82620 18637 4 wl_0_45
rlabel metal2 s 0 18809 82620 18857 4 wl_1_45
rlabel metal2 s 0 19283 82620 19331 4 wl_0_46
rlabel metal2 s 0 19063 82620 19111 4 wl_1_46
rlabel metal2 s 0 19379 82620 19427 4 wl_0_47
rlabel metal2 s 0 19599 82620 19647 4 wl_1_47
rlabel metal2 s 0 20073 82620 20121 4 wl_0_48
rlabel metal2 s 0 19853 82620 19901 4 wl_1_48
rlabel metal2 s 0 20169 82620 20217 4 wl_0_49
rlabel metal2 s 0 20389 82620 20437 4 wl_1_49
rlabel metal2 s 0 20863 82620 20911 4 wl_0_50
rlabel metal2 s 0 20643 82620 20691 4 wl_1_50
rlabel metal2 s 0 20959 82620 21007 4 wl_0_51
rlabel metal2 s 0 21179 82620 21227 4 wl_1_51
rlabel metal2 s 0 21653 82620 21701 4 wl_0_52
rlabel metal2 s 0 21433 82620 21481 4 wl_1_52
rlabel metal2 s 0 21749 82620 21797 4 wl_0_53
rlabel metal2 s 0 21969 82620 22017 4 wl_1_53
rlabel metal2 s 0 22443 82620 22491 4 wl_0_54
rlabel metal2 s 0 22223 82620 22271 4 wl_1_54
rlabel metal2 s 0 22539 82620 22587 4 wl_0_55
rlabel metal2 s 0 22759 82620 22807 4 wl_1_55
rlabel metal2 s 0 23233 82620 23281 4 wl_0_56
rlabel metal2 s 0 23013 82620 23061 4 wl_1_56
rlabel metal2 s 0 23329 82620 23377 4 wl_0_57
rlabel metal2 s 0 23549 82620 23597 4 wl_1_57
rlabel metal2 s 0 24023 82620 24071 4 wl_0_58
rlabel metal2 s 0 23803 82620 23851 4 wl_1_58
rlabel metal2 s 0 24119 82620 24167 4 wl_0_59
rlabel metal2 s 0 24339 82620 24387 4 wl_1_59
rlabel metal2 s 0 24813 82620 24861 4 wl_0_60
rlabel metal2 s 0 24593 82620 24641 4 wl_1_60
rlabel metal2 s 0 24909 82620 24957 4 wl_0_61
rlabel metal2 s 0 25129 82620 25177 4 wl_1_61
rlabel metal2 s 0 25603 82620 25651 4 wl_0_62
rlabel metal2 s 0 25383 82620 25431 4 wl_1_62
rlabel metal2 s 0 25699 82620 25747 4 wl_0_63
rlabel metal2 s 0 25919 82620 25967 4 wl_1_63
rlabel metal2 s 1080 25479 1188 25555 4 gnd
rlabel metal2 s 1080 14419 1188 14495 4 gnd
rlabel metal2 s 1080 18369 1188 18445 4 gnd
rlabel metal2 s 1080 13945 1188 14021 4 gnd
rlabel metal2 s 1080 23899 1188 23975 4 gnd
rlabel metal2 s 1080 22065 1188 22175 4 gnd
rlabel metal2 s 1080 19159 1188 19235 4 gnd
rlabel metal2 s 1080 18685 1188 18761 4 gnd
rlabel metal2 s 1080 25795 1188 25871 4 gnd
rlabel metal2 s 1080 17895 1188 17971 4 gnd
rlabel metal2 s 1080 24215 1188 24291 4 gnd
rlabel metal2 s 1080 24435 1188 24545 4 gnd
rlabel metal2 s 1080 20739 1188 20815 4 gnd
rlabel metal2 s 1080 16789 1188 16865 4 gnd
rlabel metal2 s 1080 21055 1188 21131 4 gnd
rlabel metal2 s 1080 13375 1188 13485 4 gnd
rlabel metal2 s 1080 19475 1188 19551 4 gnd
rlabel metal2 s 1080 23425 1188 23501 4 gnd
rlabel metal2 s 1080 18115 1188 18225 4 gnd
rlabel metal2 s 1080 15999 1188 16075 4 gnd
rlabel metal2 s 1080 22855 1188 22965 4 gnd
rlabel metal2 s 1080 25225 1188 25335 4 gnd
rlabel metal2 s 1080 24689 1188 24765 4 gnd
rlabel metal2 s 1080 21529 1188 21605 4 gnd
rlabel metal2 s 1080 19949 1188 20025 4 gnd
rlabel metal2 s 1080 16315 1188 16391 4 gnd
rlabel metal2 s 1080 14165 1188 14275 4 gnd
rlabel metal2 s 1080 20265 1188 20341 4 gnd
rlabel metal2 s 1080 17105 1188 17181 4 gnd
rlabel metal2 s 1080 15209 1188 15285 4 gnd
rlabel metal2 s 1080 20485 1188 20595 4 gnd
rlabel metal2 s 1080 16535 1188 16645 4 gnd
rlabel metal2 s 1080 22319 1188 22395 4 gnd
rlabel metal2 s 1080 21845 1188 21921 4 gnd
rlabel metal2 s 1080 23109 1188 23185 4 gnd
rlabel metal2 s 1080 14955 1188 15065 4 gnd
rlabel metal2 s 1080 22635 1188 22711 4 gnd
rlabel metal2 s 1080 15525 1188 15601 4 gnd
rlabel metal2 s 1080 15745 1188 15855 4 gnd
rlabel metal2 s 1080 25005 1188 25081 4 gnd
rlabel metal2 s 1080 17325 1188 17435 4 gnd
rlabel metal2 s 1080 18905 1188 19015 4 gnd
rlabel metal2 s 1080 13629 1188 13705 4 gnd
rlabel metal2 s 1080 17579 1188 17655 4 gnd
rlabel metal2 s 1080 14735 1188 14811 4 gnd
rlabel metal2 s 1080 23645 1188 23755 4 gnd
rlabel metal2 s 1080 19695 1188 19805 4 gnd
rlabel metal2 s 1080 21275 1188 21385 4 gnd
rlabel metal2 s 1080 12049 1188 12125 4 gnd
rlabel metal2 s 1080 8889 1188 8965 4 gnd
rlabel metal2 s 1080 7845 1188 7955 4 gnd
rlabel metal2 s 1080 3675 1188 3751 4 gnd
rlabel metal2 s 1080 7055 1188 7165 4 gnd
rlabel metal2 s 1080 3359 1188 3435 4 gnd
rlabel metal2 s 1080 12839 1188 12915 4 gnd
rlabel metal2 s 1080 4685 1188 4795 4 gnd
rlabel metal2 s 1080 2569 1188 2645 4 gnd
rlabel metal2 s 1080 7309 1188 7385 4 gnd
rlabel metal2 s 1080 6835 1188 6911 4 gnd
rlabel metal2 s 1080 11259 1188 11335 4 gnd
rlabel metal2 s 1080 9205 1188 9281 4 gnd
rlabel metal2 s 1080 10469 1188 10545 4 gnd
rlabel metal2 s 1080 11005 1188 11115 4 gnd
rlabel metal2 s 1080 5475 1188 5585 4 gnd
rlabel metal2 s 1080 2095 1188 2171 4 gnd
rlabel metal2 s 1080 9425 1188 9535 4 gnd
rlabel metal2 s 1080 8635 1188 8745 4 gnd
rlabel metal2 s 1080 515 1188 591 4 gnd
rlabel metal2 s 1080 3895 1188 4005 4 gnd
rlabel metal2 s 1080 8099 1188 8175 4 gnd
rlabel metal2 s 1080 11575 1188 11651 4 gnd
rlabel metal2 s 1080 5729 1188 5805 4 gnd
rlabel metal2 s 1080 13155 1188 13231 4 gnd
rlabel metal2 s 1080 4939 1188 5015 4 gnd
rlabel metal2 s 1080 8415 1188 8491 4 gnd
rlabel metal2 s 1080 2315 1188 2425 4 gnd
rlabel metal2 s 1080 2885 1188 2961 4 gnd
rlabel metal2 s 1080 12365 1188 12441 4 gnd
rlabel metal2 s 1080 10785 1188 10861 4 gnd
rlabel metal2 s 1080 11795 1188 11905 4 gnd
rlabel metal2 s 1080 12585 1188 12695 4 gnd
rlabel metal2 s 1080 1779 1188 1855 4 gnd
rlabel metal2 s 1080 1525 1188 1635 4 gnd
rlabel metal2 s 1080 6045 1188 6121 4 gnd
rlabel metal2 s 1080 5255 1188 5331 4 gnd
rlabel metal2 s 1080 1305 1188 1381 4 gnd
rlabel metal2 s 1080 989 1188 1065 4 gnd
rlabel metal2 s 1080 4149 1188 4225 4 gnd
rlabel metal2 s 1080 10215 1188 10325 4 gnd
rlabel metal2 s 1080 4465 1188 4541 4 gnd
rlabel metal2 s 1080 735 1188 845 4 gnd
rlabel metal2 s 1080 6265 1188 6375 4 gnd
rlabel metal2 s 1080 9995 1188 10071 4 gnd
rlabel metal2 s 1080 3105 1188 3215 4 gnd
rlabel metal2 s 1080 7625 1188 7701 4 gnd
rlabel metal2 s 1080 9679 1188 9755 4 gnd
rlabel metal2 s 1080 6519 1188 6595 4 gnd
rlabel metal2 s 0 10373 82620 10421 4 wl_1_24
rlabel metal2 s 0 4369 82620 4417 4 wl_0_9
rlabel metal2 s 0 4589 82620 4637 4 wl_1_9
rlabel metal2 s 0 5063 82620 5111 4 wl_0_10
rlabel metal2 s 0 4843 82620 4891 4 wl_1_10
rlabel metal2 s 0 5159 82620 5207 4 wl_0_11
rlabel metal2 s 0 893 82620 941 4 wl_1_0
rlabel metal2 s 0 5379 82620 5427 4 wl_1_11
rlabel metal2 s 0 11699 82620 11747 4 wl_1_27
rlabel metal2 s 0 1209 82620 1257 4 wl_0_1
rlabel metal2 s 0 12173 82620 12221 4 wl_0_28
rlabel metal2 s 0 5853 82620 5901 4 wl_0_12
rlabel metal2 s 0 5633 82620 5681 4 wl_1_12
rlabel metal2 s 0 5949 82620 5997 4 wl_0_13
rlabel metal2 s 0 1429 82620 1477 4 wl_1_1
rlabel metal2 s 0 1903 82620 1951 4 wl_0_2
rlabel metal2 s 0 9899 82620 9947 4 wl_0_23
rlabel metal2 s 0 6169 82620 6217 4 wl_1_13
rlabel metal2 s 0 6643 82620 6691 4 wl_0_14
rlabel metal2 s 0 6423 82620 6471 4 wl_1_14
rlabel metal2 s 0 1683 82620 1731 4 wl_1_2
rlabel metal2 s 0 6739 82620 6787 4 wl_0_15
rlabel metal2 s 0 1999 82620 2047 4 wl_0_3
rlabel metal2 s 0 6959 82620 7007 4 wl_1_15
rlabel metal2 s 0 2219 82620 2267 4 wl_1_3
rlabel metal2 s 0 11953 82620 12001 4 wl_1_28
rlabel metal2 s 0 10689 82620 10737 4 wl_0_25
rlabel metal2 s 0 12269 82620 12317 4 wl_0_29
rlabel metal2 s 0 2693 82620 2741 4 wl_0_4
rlabel metal2 s 0 7433 82620 7481 4 wl_0_16
rlabel metal2 s 0 12489 82620 12537 4 wl_1_29
rlabel metal2 s 0 2473 82620 2521 4 wl_1_4
rlabel metal2 s 0 2789 82620 2837 4 wl_0_5
rlabel metal2 s 0 3009 82620 3057 4 wl_1_5
rlabel metal2 s 0 12963 82620 13011 4 wl_0_30
rlabel metal2 s 0 7213 82620 7261 4 wl_1_16
rlabel metal2 s 0 7529 82620 7577 4 wl_0_17
rlabel metal2 s 0 7749 82620 7797 4 wl_1_17
rlabel metal2 s 0 8223 82620 8271 4 wl_0_18
rlabel metal2 s 0 8003 82620 8051 4 wl_1_18
rlabel metal2 s 0 3483 82620 3531 4 wl_0_6
rlabel metal2 s 0 3263 82620 3311 4 wl_1_6
rlabel metal2 s 0 3579 82620 3627 4 wl_0_7
rlabel metal2 s 0 3799 82620 3847 4 wl_1_7
rlabel metal2 s 0 10909 82620 10957 4 wl_1_25
rlabel metal2 s 0 12743 82620 12791 4 wl_1_30
rlabel metal2 s 0 13059 82620 13107 4 wl_0_31
rlabel metal2 s 0 4273 82620 4321 4 wl_0_8
rlabel metal2 s 0 8319 82620 8367 4 wl_0_19
rlabel metal2 s 0 8539 82620 8587 4 wl_1_19
rlabel metal2 s 0 9583 82620 9631 4 wl_1_22
rlabel metal2 s 0 10119 82620 10167 4 wl_1_23
rlabel metal2 s 0 10593 82620 10641 4 wl_0_24
rlabel metal2 s 0 11383 82620 11431 4 wl_0_26
rlabel metal2 s 0 9013 82620 9061 4 wl_0_20
rlabel metal2 s 0 8793 82620 8841 4 wl_1_20
rlabel metal2 s 0 419 82620 467 4 rbl_wl_0_0
rlabel metal2 s 0 9109 82620 9157 4 wl_0_21
rlabel metal2 s 0 9329 82620 9377 4 wl_1_21
rlabel metal2 s 0 11163 82620 11211 4 wl_1_26
rlabel metal2 s 0 1113 82620 1161 4 wl_0_0
rlabel metal2 s 0 11479 82620 11527 4 wl_0_27
rlabel metal2 s 0 4053 82620 4101 4 wl_1_8
rlabel metal2 s 0 9803 82620 9851 4 wl_0_22
rlabel metal2 s 81432 22635 81540 22711 4 gnd
rlabel metal2 s 81432 8635 81540 8745 4 gnd
rlabel metal2 s 81432 19695 81540 19805 4 gnd
rlabel metal2 s 81432 19949 81540 20025 4 gnd
rlabel metal2 s 81432 23425 81540 23501 4 gnd
rlabel metal2 s 81432 11795 81540 11905 4 gnd
rlabel metal2 s 81432 23109 81540 23185 4 gnd
rlabel metal2 s 81432 15999 81540 16075 4 gnd
rlabel metal2 s 81432 7055 81540 7165 4 gnd
rlabel metal2 s 81432 16789 81540 16865 4 gnd
rlabel metal2 s 81432 9425 81540 9535 4 gnd
rlabel metal2 s 81432 20485 81540 20595 4 gnd
rlabel metal2 s 81432 16535 81540 16645 4 gnd
rlabel metal2 s 81432 13375 81540 13485 4 gnd
rlabel metal2 s 81432 9205 81540 9281 4 gnd
rlabel metal2 s 81432 2885 81540 2961 4 gnd
rlabel metal2 s 81432 5255 81540 5331 4 gnd
rlabel metal2 s 81432 11005 81540 11115 4 gnd
rlabel metal2 s 81432 6265 81540 6375 4 gnd
rlabel metal2 s 81432 7845 81540 7955 4 gnd
rlabel metal2 s 81432 7309 81540 7385 4 gnd
rlabel metal2 s 81432 25225 81540 25335 4 gnd
rlabel metal2 s 81432 2095 81540 2171 4 gnd
rlabel metal2 s 81432 6045 81540 6121 4 gnd
rlabel metal2 s 81432 3895 81540 4005 4 gnd
rlabel metal2 s 81432 4149 81540 4225 4 gnd
rlabel metal2 s 81432 22855 81540 22965 4 gnd
rlabel metal2 s 81432 12365 81540 12441 4 gnd
rlabel metal2 s 81432 7625 81540 7701 4 gnd
rlabel metal2 s 81432 515 81540 591 4 gnd
rlabel metal2 s 81432 20739 81540 20815 4 gnd
rlabel metal2 s 81432 8415 81540 8491 4 gnd
rlabel metal2 s 81432 17105 81540 17181 4 gnd
rlabel metal2 s 81432 22065 81540 22175 4 gnd
rlabel metal2 s 81432 15209 81540 15285 4 gnd
rlabel metal2 s 81432 735 81540 845 4 gnd
rlabel metal2 s 81432 5729 81540 5805 4 gnd
rlabel metal2 s 81432 18115 81540 18225 4 gnd
rlabel metal2 s 81432 4465 81540 4541 4 gnd
rlabel metal2 s 81432 25479 81540 25555 4 gnd
rlabel metal2 s 81432 18685 81540 18761 4 gnd
rlabel metal2 s 81432 13629 81540 13705 4 gnd
rlabel metal2 s 81432 25005 81540 25081 4 gnd
rlabel metal2 s 81432 21055 81540 21131 4 gnd
rlabel metal2 s 81432 1305 81540 1381 4 gnd
rlabel metal2 s 81432 18369 81540 18445 4 gnd
rlabel metal2 s 81432 989 81540 1065 4 gnd
rlabel metal2 s 81432 14419 81540 14495 4 gnd
rlabel metal2 s 81432 13155 81540 13231 4 gnd
rlabel metal2 s 81432 15525 81540 15601 4 gnd
rlabel metal2 s 81432 10469 81540 10545 4 gnd
rlabel metal2 s 81432 14735 81540 14811 4 gnd
rlabel metal2 s 81432 11575 81540 11651 4 gnd
rlabel metal2 s 81432 3675 81540 3751 4 gnd
rlabel metal2 s 81432 11259 81540 11335 4 gnd
rlabel metal2 s 81432 8889 81540 8965 4 gnd
rlabel metal2 s 81432 17579 81540 17655 4 gnd
rlabel metal2 s 81432 14165 81540 14275 4 gnd
rlabel metal2 s 81432 24435 81540 24545 4 gnd
rlabel metal2 s 81432 18905 81540 19015 4 gnd
rlabel metal2 s 81432 17325 81540 17435 4 gnd
rlabel metal2 s 81432 6835 81540 6911 4 gnd
rlabel metal2 s 81432 21275 81540 21385 4 gnd
rlabel metal2 s 81432 23645 81540 23755 4 gnd
rlabel metal2 s 81432 12049 81540 12125 4 gnd
rlabel metal2 s 81432 8099 81540 8175 4 gnd
rlabel metal2 s 81432 12585 81540 12695 4 gnd
rlabel metal2 s 81432 10785 81540 10861 4 gnd
rlabel metal2 s 81432 22319 81540 22395 4 gnd
rlabel metal2 s 81432 6519 81540 6595 4 gnd
rlabel metal2 s 81432 14955 81540 15065 4 gnd
rlabel metal2 s 81432 3359 81540 3435 4 gnd
rlabel metal2 s 81432 2569 81540 2645 4 gnd
rlabel metal2 s 81432 16315 81540 16391 4 gnd
rlabel metal2 s 81432 19159 81540 19235 4 gnd
rlabel metal2 s 81432 13945 81540 14021 4 gnd
rlabel metal2 s 81432 10215 81540 10325 4 gnd
rlabel metal2 s 81432 24689 81540 24765 4 gnd
rlabel metal2 s 81432 1525 81540 1635 4 gnd
rlabel metal2 s 81432 24215 81540 24291 4 gnd
rlabel metal2 s 81432 9679 81540 9755 4 gnd
rlabel metal2 s 81432 20265 81540 20341 4 gnd
rlabel metal2 s 81432 19475 81540 19551 4 gnd
rlabel metal2 s 81432 21845 81540 21921 4 gnd
rlabel metal2 s 81432 3105 81540 3215 4 gnd
rlabel metal2 s 81432 21529 81540 21605 4 gnd
rlabel metal2 s 81432 12839 81540 12915 4 gnd
rlabel metal2 s 81432 25795 81540 25871 4 gnd
rlabel metal2 s 81432 5475 81540 5585 4 gnd
rlabel metal2 s 81432 2315 81540 2425 4 gnd
rlabel metal2 s 81432 4939 81540 5015 4 gnd
rlabel metal2 s 81432 9995 81540 10071 4 gnd
rlabel metal2 s 81432 15745 81540 15855 4 gnd
rlabel metal2 s 81432 23899 81540 23975 4 gnd
rlabel metal2 s 81432 1779 81540 1855 4 gnd
rlabel metal2 s 81432 4685 81540 4795 4 gnd
rlabel metal2 s 81432 17895 81540 17971 4 gnd
rlabel metal1 s 81468 39579 81504 39920 4 vdd
rlabel metal1 s 81468 26440 81504 26781 4 vdd
rlabel metal1 s 81468 35920 81504 36261 4 vdd
rlabel metal1 s 81468 38789 81504 39130 4 vdd
rlabel metal1 s 81468 28519 81504 28860 4 vdd
rlabel metal1 s 81468 31180 81504 31521 4 vdd
rlabel metal1 s 81468 42240 81504 42581 4 vdd
rlabel metal1 s 81468 28020 81504 28361 4 vdd
rlabel metal1 s 81468 41949 81504 42290 4 vdd
rlabel metal1 s 81468 47479 81504 47820 4 vdd
rlabel metal1 s 81468 41159 81504 41500 4 vdd
rlabel metal1 s 81468 32760 81504 33101 4 vdd
rlabel metal1 s 81468 27230 81504 27571 4 vdd
rlabel metal1 s 81468 27729 81504 28070 4 vdd
rlabel metal1 s 81468 44319 81504 44660 4 vdd
rlabel metal1 s 81468 37999 81504 38340 4 vdd
rlabel metal1 s 81468 34049 81504 34390 4 vdd
rlabel metal1 s 81468 35130 81504 35471 4 vdd
rlabel metal1 s 81468 34340 81504 34681 4 vdd
rlabel metal1 s 81468 46190 81504 46531 4 vdd
rlabel metal1 s 81468 26939 81504 27280 4 vdd
rlabel metal1 s 81468 36710 81504 37051 4 vdd
rlabel metal1 s 81468 30099 81504 30440 4 vdd
rlabel metal1 s 81468 33550 81504 33891 4 vdd
rlabel metal1 s 81468 41450 81504 41791 4 vdd
rlabel metal1 s 81468 37500 81504 37841 4 vdd
rlabel metal1 s 81468 42739 81504 43080 4 vdd
rlabel metal1 s 81468 39080 81504 39421 4 vdd
rlabel metal1 s 81468 34839 81504 35180 4 vdd
rlabel metal1 s 81468 31679 81504 32020 4 vdd
rlabel metal1 s 81468 33259 81504 33600 4 vdd
rlabel metal1 s 81468 30390 81504 30731 4 vdd
rlabel metal1 s 81468 32469 81504 32810 4 vdd
rlabel metal1 s 81468 43820 81504 44161 4 vdd
rlabel metal1 s 81468 40660 81504 41001 4 vdd
rlabel metal1 s 81468 38290 81504 38631 4 vdd
rlabel metal1 s 81468 45109 81504 45450 4 vdd
rlabel metal1 s 81468 50639 81504 50980 4 vdd
rlabel metal1 s 81468 36419 81504 36760 4 vdd
rlabel metal1 s 81468 29600 81504 29941 4 vdd
rlabel metal1 s 81468 39870 81504 40211 4 vdd
rlabel metal1 s 81468 29309 81504 29650 4 vdd
rlabel metal1 s 81468 50930 81504 51271 4 vdd
rlabel metal1 s 81468 45400 81504 45741 4 vdd
rlabel metal1 s 81468 45899 81504 46240 4 vdd
rlabel metal1 s 81468 40369 81504 40710 4 vdd
rlabel metal1 s 81468 43030 81504 43371 4 vdd
rlabel metal1 s 81468 46980 81504 47321 4 vdd
rlabel metal1 s 81468 35629 81504 35970 4 vdd
rlabel metal1 s 81468 49350 81504 49691 4 vdd
rlabel metal1 s 81468 50140 81504 50481 4 vdd
rlabel metal1 s 81468 44610 81504 44951 4 vdd
rlabel metal1 s 81468 43529 81504 43870 4 vdd
rlabel metal1 s 81468 49849 81504 50190 4 vdd
rlabel metal1 s 81468 49059 81504 49400 4 vdd
rlabel metal1 s 81468 46689 81504 47030 4 vdd
rlabel metal1 s 81468 48269 81504 48610 4 vdd
rlabel metal1 s 81468 26149 81504 26490 4 vdd
rlabel metal1 s 81468 28810 81504 29151 4 vdd
rlabel metal1 s 81468 48560 81504 48901 4 vdd
rlabel metal1 s 81468 30889 81504 31230 4 vdd
rlabel metal1 s 81468 47770 81504 48111 4 vdd
rlabel metal1 s 81468 37209 81504 37550 4 vdd
rlabel metal1 s 81468 31970 81504 32311 4 vdd
rlabel metal1 s 81468 51429 81504 51770 4 vdd
rlabel metal1 s 1116 50140 1152 50481 4 vdd
rlabel metal1 s 1116 36419 1152 36760 4 vdd
rlabel metal1 s 1116 27729 1152 28070 4 vdd
rlabel metal1 s 1116 41949 1152 42290 4 vdd
rlabel metal1 s 1116 41450 1152 41791 4 vdd
rlabel metal1 s 1116 40369 1152 40710 4 vdd
rlabel metal1 s 1116 50639 1152 50980 4 vdd
rlabel metal1 s 1116 28020 1152 28361 4 vdd
rlabel metal1 s 1116 37209 1152 37550 4 vdd
rlabel metal1 s 1116 31970 1152 32311 4 vdd
rlabel metal1 s 1116 45109 1152 45450 4 vdd
rlabel metal1 s 1116 30889 1152 31230 4 vdd
rlabel metal1 s 1116 35920 1152 36261 4 vdd
rlabel metal1 s 1116 41159 1152 41500 4 vdd
rlabel metal1 s 1116 28810 1152 29151 4 vdd
rlabel metal1 s 1116 49350 1152 49691 4 vdd
rlabel metal1 s 1116 47770 1152 48111 4 vdd
rlabel metal1 s 1116 30390 1152 30731 4 vdd
rlabel metal1 s 1116 37500 1152 37841 4 vdd
rlabel metal1 s 1116 31180 1152 31521 4 vdd
rlabel metal1 s 1116 49059 1152 49400 4 vdd
rlabel metal1 s 1116 35629 1152 35970 4 vdd
rlabel metal1 s 1116 34839 1152 35180 4 vdd
rlabel metal1 s 1116 32760 1152 33101 4 vdd
rlabel metal1 s 1116 43030 1152 43371 4 vdd
rlabel metal1 s 1116 30099 1152 30440 4 vdd
rlabel metal1 s 1116 45899 1152 46240 4 vdd
rlabel metal1 s 1116 33550 1152 33891 4 vdd
rlabel metal1 s 1116 32469 1152 32810 4 vdd
rlabel metal1 s 1116 29600 1152 29941 4 vdd
rlabel metal1 s 1116 42240 1152 42581 4 vdd
rlabel metal1 s 1116 48269 1152 48610 4 vdd
rlabel metal1 s 1116 42739 1152 43080 4 vdd
rlabel metal1 s 1116 26440 1152 26781 4 vdd
rlabel metal1 s 1116 40660 1152 41001 4 vdd
rlabel metal1 s 1116 34340 1152 34681 4 vdd
rlabel metal1 s 1116 35130 1152 35471 4 vdd
rlabel metal1 s 1116 44610 1152 44951 4 vdd
rlabel metal1 s 1116 29309 1152 29650 4 vdd
rlabel metal1 s 1116 43820 1152 44161 4 vdd
rlabel metal1 s 1116 39080 1152 39421 4 vdd
rlabel metal1 s 1116 31679 1152 32020 4 vdd
rlabel metal1 s 1116 43529 1152 43870 4 vdd
rlabel metal1 s 1116 37999 1152 38340 4 vdd
rlabel metal1 s 1116 27230 1152 27571 4 vdd
rlabel metal1 s 1116 26149 1152 26490 4 vdd
rlabel metal1 s 1116 46980 1152 47321 4 vdd
rlabel metal1 s 1116 44319 1152 44660 4 vdd
rlabel metal1 s 1116 47479 1152 47820 4 vdd
rlabel metal1 s 1116 46190 1152 46531 4 vdd
rlabel metal1 s 1116 34049 1152 34390 4 vdd
rlabel metal1 s 1116 50930 1152 51271 4 vdd
rlabel metal1 s 1116 33259 1152 33600 4 vdd
rlabel metal1 s 1116 48560 1152 48901 4 vdd
rlabel metal1 s 1116 51429 1152 51770 4 vdd
rlabel metal1 s 1116 26939 1152 27280 4 vdd
rlabel metal1 s 1116 36710 1152 37051 4 vdd
rlabel metal1 s 1116 38290 1152 38631 4 vdd
rlabel metal1 s 1116 39579 1152 39920 4 vdd
rlabel metal1 s 1116 38789 1152 39130 4 vdd
rlabel metal1 s 1116 46689 1152 47030 4 vdd
rlabel metal1 s 1116 28519 1152 28860 4 vdd
rlabel metal1 s 1116 45400 1152 45741 4 vdd
rlabel metal1 s 1116 39870 1152 40211 4 vdd
rlabel metal1 s 1116 49849 1152 50190 4 vdd
rlabel metal1 s 31404 0 31440 52140 4 bl_0_48
rlabel metal1 s 31620 0 31656 52140 4 bl_1_48
rlabel metal1 s 31476 0 31512 52140 4 br_0_48
rlabel metal1 s 31692 0 31728 52140 4 br_1_48
rlabel metal1 s 32460 0 32496 52140 4 bl_0_49
rlabel metal1 s 32244 0 32280 52140 4 bl_1_49
rlabel metal1 s 32388 0 32424 52140 4 br_0_49
rlabel metal1 s 32172 0 32208 52140 4 br_1_49
rlabel metal1 s 32652 0 32688 52140 4 bl_0_50
rlabel metal1 s 32868 0 32904 52140 4 bl_1_50
rlabel metal1 s 32724 0 32760 52140 4 br_0_50
rlabel metal1 s 32940 0 32976 52140 4 br_1_50
rlabel metal1 s 33708 0 33744 52140 4 bl_0_51
rlabel metal1 s 33492 0 33528 52140 4 bl_1_51
rlabel metal1 s 33636 0 33672 52140 4 br_0_51
rlabel metal1 s 33420 0 33456 52140 4 br_1_51
rlabel metal1 s 33900 0 33936 52140 4 bl_0_52
rlabel metal1 s 34116 0 34152 52140 4 bl_1_52
rlabel metal1 s 33972 0 34008 52140 4 br_0_52
rlabel metal1 s 34188 0 34224 52140 4 br_1_52
rlabel metal1 s 34956 0 34992 52140 4 bl_0_53
rlabel metal1 s 34740 0 34776 52140 4 bl_1_53
rlabel metal1 s 34884 0 34920 52140 4 br_0_53
rlabel metal1 s 34668 0 34704 52140 4 br_1_53
rlabel metal1 s 35148 0 35184 52140 4 bl_0_54
rlabel metal1 s 35364 0 35400 52140 4 bl_1_54
rlabel metal1 s 35220 0 35256 52140 4 br_0_54
rlabel metal1 s 35436 0 35472 52140 4 br_1_54
rlabel metal1 s 36204 0 36240 52140 4 bl_0_55
rlabel metal1 s 35988 0 36024 52140 4 bl_1_55
rlabel metal1 s 36132 0 36168 52140 4 br_0_55
rlabel metal1 s 35916 0 35952 52140 4 br_1_55
rlabel metal1 s 36396 0 36432 52140 4 bl_0_56
rlabel metal1 s 36612 0 36648 52140 4 bl_1_56
rlabel metal1 s 36468 0 36504 52140 4 br_0_56
rlabel metal1 s 36684 0 36720 52140 4 br_1_56
rlabel metal1 s 37452 0 37488 52140 4 bl_0_57
rlabel metal1 s 37236 0 37272 52140 4 bl_1_57
rlabel metal1 s 37380 0 37416 52140 4 br_0_57
rlabel metal1 s 37164 0 37200 52140 4 br_1_57
rlabel metal1 s 37644 0 37680 52140 4 bl_0_58
rlabel metal1 s 37860 0 37896 52140 4 bl_1_58
rlabel metal1 s 37716 0 37752 52140 4 br_0_58
rlabel metal1 s 37932 0 37968 52140 4 br_1_58
rlabel metal1 s 38700 0 38736 52140 4 bl_0_59
rlabel metal1 s 38484 0 38520 52140 4 bl_1_59
rlabel metal1 s 38628 0 38664 52140 4 br_0_59
rlabel metal1 s 38412 0 38448 52140 4 br_1_59
rlabel metal1 s 38892 0 38928 52140 4 bl_0_60
rlabel metal1 s 39108 0 39144 52140 4 bl_1_60
rlabel metal1 s 38964 0 39000 52140 4 br_0_60
rlabel metal1 s 39180 0 39216 52140 4 br_1_60
rlabel metal1 s 39948 0 39984 52140 4 bl_0_61
rlabel metal1 s 39732 0 39768 52140 4 bl_1_61
rlabel metal1 s 39876 0 39912 52140 4 br_0_61
rlabel metal1 s 39660 0 39696 52140 4 br_1_61
rlabel metal1 s 40140 0 40176 52140 4 bl_0_62
rlabel metal1 s 40356 0 40392 52140 4 bl_1_62
rlabel metal1 s 40212 0 40248 52140 4 br_0_62
rlabel metal1 s 40428 0 40464 52140 4 br_1_62
rlabel metal1 s 41196 0 41232 52140 4 bl_0_63
rlabel metal1 s 40980 0 41016 52140 4 bl_1_63
rlabel metal1 s 41124 0 41160 52140 4 br_0_63
rlabel metal1 s 40908 0 40944 52140 4 br_1_63
rlabel metal1 s 22476 0 22512 52140 4 bl_0_33
rlabel metal1 s 22260 0 22296 52140 4 bl_1_33
rlabel metal1 s 22404 0 22440 52140 4 br_0_33
rlabel metal1 s 22188 0 22224 52140 4 br_1_33
rlabel metal1 s 22668 0 22704 52140 4 bl_0_34
rlabel metal1 s 22884 0 22920 52140 4 bl_1_34
rlabel metal1 s 22740 0 22776 52140 4 br_0_34
rlabel metal1 s 22956 0 22992 52140 4 br_1_34
rlabel metal1 s 23724 0 23760 52140 4 bl_0_35
rlabel metal1 s 23508 0 23544 52140 4 bl_1_35
rlabel metal1 s 23652 0 23688 52140 4 br_0_35
rlabel metal1 s 23436 0 23472 52140 4 br_1_35
rlabel metal1 s 23916 0 23952 52140 4 bl_0_36
rlabel metal1 s 24132 0 24168 52140 4 bl_1_36
rlabel metal1 s 23988 0 24024 52140 4 br_0_36
rlabel metal1 s 24204 0 24240 52140 4 br_1_36
rlabel metal1 s 24972 0 25008 52140 4 bl_0_37
rlabel metal1 s 24756 0 24792 52140 4 bl_1_37
rlabel metal1 s 24900 0 24936 52140 4 br_0_37
rlabel metal1 s 24684 0 24720 52140 4 br_1_37
rlabel metal1 s 25164 0 25200 52140 4 bl_0_38
rlabel metal1 s 25380 0 25416 52140 4 bl_1_38
rlabel metal1 s 25236 0 25272 52140 4 br_0_38
rlabel metal1 s 25452 0 25488 52140 4 br_1_38
rlabel metal1 s 26220 0 26256 52140 4 bl_0_39
rlabel metal1 s 26004 0 26040 52140 4 bl_1_39
rlabel metal1 s 26148 0 26184 52140 4 br_0_39
rlabel metal1 s 25932 0 25968 52140 4 br_1_39
rlabel metal1 s 26412 0 26448 52140 4 bl_0_40
rlabel metal1 s 26628 0 26664 52140 4 bl_1_40
rlabel metal1 s 26484 0 26520 52140 4 br_0_40
rlabel metal1 s 26700 0 26736 52140 4 br_1_40
rlabel metal1 s 27468 0 27504 52140 4 bl_0_41
rlabel metal1 s 27252 0 27288 52140 4 bl_1_41
rlabel metal1 s 27396 0 27432 52140 4 br_0_41
rlabel metal1 s 27180 0 27216 52140 4 br_1_41
rlabel metal1 s 27660 0 27696 52140 4 bl_0_42
rlabel metal1 s 27876 0 27912 52140 4 bl_1_42
rlabel metal1 s 27732 0 27768 52140 4 br_0_42
rlabel metal1 s 27948 0 27984 52140 4 br_1_42
rlabel metal1 s 28716 0 28752 52140 4 bl_0_43
rlabel metal1 s 28500 0 28536 52140 4 bl_1_43
rlabel metal1 s 28644 0 28680 52140 4 br_0_43
rlabel metal1 s 28428 0 28464 52140 4 br_1_43
rlabel metal1 s 28908 0 28944 52140 4 bl_0_44
rlabel metal1 s 29124 0 29160 52140 4 bl_1_44
rlabel metal1 s 28980 0 29016 52140 4 br_0_44
rlabel metal1 s 29196 0 29232 52140 4 br_1_44
rlabel metal1 s 29964 0 30000 52140 4 bl_0_45
rlabel metal1 s 29748 0 29784 52140 4 bl_1_45
rlabel metal1 s 29892 0 29928 52140 4 br_0_45
rlabel metal1 s 29676 0 29712 52140 4 br_1_45
rlabel metal1 s 30156 0 30192 52140 4 bl_0_46
rlabel metal1 s 30372 0 30408 52140 4 bl_1_46
rlabel metal1 s 30228 0 30264 52140 4 br_0_46
rlabel metal1 s 30444 0 30480 52140 4 br_1_46
rlabel metal1 s 31212 0 31248 52140 4 bl_0_47
rlabel metal1 s 30996 0 31032 52140 4 bl_1_47
rlabel metal1 s 31140 0 31176 52140 4 br_0_47
rlabel metal1 s 30924 0 30960 52140 4 br_1_47
rlabel metal1 s 21492 0 21528 52140 4 br_0_32
rlabel metal1 s 21708 0 21744 52140 4 br_1_32
rlabel metal1 s 21228 0 21264 52140 4 bl_0_31
rlabel metal1 s 21156 0 21192 52140 4 br_0_31
rlabel metal1 s 21420 0 21456 52140 4 bl_0_32
rlabel metal1 s 21636 0 21672 52140 4 bl_1_32
rlabel metal1 s 11244 0 11280 52140 4 bl_0_15
rlabel metal1 s 11172 0 11208 52140 4 br_0_15
rlabel metal1 s 11436 0 11472 52140 4 bl_0_16
rlabel metal1 s 11652 0 11688 52140 4 bl_1_16
rlabel metal1 s 11508 0 11544 52140 4 br_0_16
rlabel metal1 s 11724 0 11760 52140 4 br_1_16
rlabel metal1 s 12492 0 12528 52140 4 bl_0_17
rlabel metal1 s 12276 0 12312 52140 4 bl_1_17
rlabel metal1 s 12420 0 12456 52140 4 br_0_17
rlabel metal1 s 12204 0 12240 52140 4 br_1_17
rlabel metal1 s 12684 0 12720 52140 4 bl_0_18
rlabel metal1 s 12900 0 12936 52140 4 bl_1_18
rlabel metal1 s 12756 0 12792 52140 4 br_0_18
rlabel metal1 s 12972 0 13008 52140 4 br_1_18
rlabel metal1 s 13740 0 13776 52140 4 bl_0_19
rlabel metal1 s 13524 0 13560 52140 4 bl_1_19
rlabel metal1 s 13668 0 13704 52140 4 br_0_19
rlabel metal1 s 13452 0 13488 52140 4 br_1_19
rlabel metal1 s 13932 0 13968 52140 4 bl_0_20
rlabel metal1 s 14148 0 14184 52140 4 bl_1_20
rlabel metal1 s 14004 0 14040 52140 4 br_0_20
rlabel metal1 s 14220 0 14256 52140 4 br_1_20
rlabel metal1 s 14988 0 15024 52140 4 bl_0_21
rlabel metal1 s 14772 0 14808 52140 4 bl_1_21
rlabel metal1 s 14916 0 14952 52140 4 br_0_21
rlabel metal1 s 14700 0 14736 52140 4 br_1_21
rlabel metal1 s 15180 0 15216 52140 4 bl_0_22
rlabel metal1 s 15396 0 15432 52140 4 bl_1_22
rlabel metal1 s 15252 0 15288 52140 4 br_0_22
rlabel metal1 s 15468 0 15504 52140 4 br_1_22
rlabel metal1 s 16236 0 16272 52140 4 bl_0_23
rlabel metal1 s 16020 0 16056 52140 4 bl_1_23
rlabel metal1 s 16164 0 16200 52140 4 br_0_23
rlabel metal1 s 15948 0 15984 52140 4 br_1_23
rlabel metal1 s 16428 0 16464 52140 4 bl_0_24
rlabel metal1 s 16644 0 16680 52140 4 bl_1_24
rlabel metal1 s 16500 0 16536 52140 4 br_0_24
rlabel metal1 s 16716 0 16752 52140 4 br_1_24
rlabel metal1 s 17484 0 17520 52140 4 bl_0_25
rlabel metal1 s 17268 0 17304 52140 4 bl_1_25
rlabel metal1 s 17412 0 17448 52140 4 br_0_25
rlabel metal1 s 17196 0 17232 52140 4 br_1_25
rlabel metal1 s 17676 0 17712 52140 4 bl_0_26
rlabel metal1 s 17892 0 17928 52140 4 bl_1_26
rlabel metal1 s 17748 0 17784 52140 4 br_0_26
rlabel metal1 s 17964 0 18000 52140 4 br_1_26
rlabel metal1 s 18732 0 18768 52140 4 bl_0_27
rlabel metal1 s 18516 0 18552 52140 4 bl_1_27
rlabel metal1 s 18660 0 18696 52140 4 br_0_27
rlabel metal1 s 18444 0 18480 52140 4 br_1_27
rlabel metal1 s 18924 0 18960 52140 4 bl_0_28
rlabel metal1 s 19140 0 19176 52140 4 bl_1_28
rlabel metal1 s 18996 0 19032 52140 4 br_0_28
rlabel metal1 s 19212 0 19248 52140 4 br_1_28
rlabel metal1 s 19980 0 20016 52140 4 bl_0_29
rlabel metal1 s 19764 0 19800 52140 4 bl_1_29
rlabel metal1 s 19908 0 19944 52140 4 br_0_29
rlabel metal1 s 19692 0 19728 52140 4 br_1_29
rlabel metal1 s 20172 0 20208 52140 4 bl_0_30
rlabel metal1 s 20388 0 20424 52140 4 bl_1_30
rlabel metal1 s 20244 0 20280 52140 4 br_0_30
rlabel metal1 s 20460 0 20496 52140 4 br_1_30
rlabel metal1 s 21012 0 21048 52140 4 bl_1_31
rlabel metal1 s 20940 0 20976 52140 4 br_1_31
rlabel metal1 s 1452 0 1488 52140 4 bl_0_0
rlabel metal1 s 11028 0 11064 52140 4 bl_1_15
rlabel metal1 s 1668 0 1704 52140 4 bl_1_0
rlabel metal1 s 10956 0 10992 52140 4 br_1_15
rlabel metal1 s 1524 0 1560 52140 4 br_0_0
rlabel metal1 s 1116 20619 1152 20960 4 vdd
rlabel metal1 s 1740 0 1776 52140 4 br_1_0
rlabel metal1 s 2508 0 2544 52140 4 bl_0_1
rlabel metal1 s 2292 0 2328 52140 4 bl_1_1
rlabel metal1 s 2436 0 2472 52140 4 br_0_1
rlabel metal1 s 2220 0 2256 52140 4 br_1_1
rlabel metal1 s 2700 0 2736 52140 4 bl_0_2
rlabel metal1 s 2916 0 2952 52140 4 bl_1_2
rlabel metal1 s 2772 0 2808 52140 4 br_0_2
rlabel metal1 s 2988 0 3024 52140 4 br_1_2
rlabel metal1 s 3756 0 3792 52140 4 bl_0_3
rlabel metal1 s 3540 0 3576 52140 4 bl_1_3
rlabel metal1 s 3684 0 3720 52140 4 br_0_3
rlabel metal1 s 1116 22199 1152 22540 4 vdd
rlabel metal1 s 3468 0 3504 52140 4 br_1_3
rlabel metal1 s 3948 0 3984 52140 4 bl_0_4
rlabel metal1 s 4164 0 4200 52140 4 bl_1_4
rlabel metal1 s 4020 0 4056 52140 4 br_0_4
rlabel metal1 s 1116 22490 1152 22831 4 vdd
rlabel metal1 s 1116 24070 1152 24411 4 vdd
rlabel metal1 s 4236 0 4272 52140 4 br_1_4
rlabel metal1 s 1116 20120 1152 20461 4 vdd
rlabel metal1 s 5004 0 5040 52140 4 bl_0_5
rlabel metal1 s 4788 0 4824 52140 4 bl_1_5
rlabel metal1 s 4932 0 4968 52140 4 br_0_5
rlabel metal1 s 1116 25650 1152 25991 4 vdd
rlabel metal1 s 4716 0 4752 52140 4 br_1_5
rlabel metal1 s 5196 0 5232 52140 4 bl_0_6
rlabel metal1 s 5412 0 5448 52140 4 bl_1_6
rlabel metal1 s 1116 21409 1152 21750 4 vdd
rlabel metal1 s 5268 0 5304 52140 4 br_0_6
rlabel metal1 s 1116 20910 1152 21251 4 vdd
rlabel metal1 s 1116 22989 1152 23330 4 vdd
rlabel metal1 s 5484 0 5520 52140 4 br_1_6
rlabel metal1 s 6252 0 6288 52140 4 bl_0_7
rlabel metal1 s 6036 0 6072 52140 4 bl_1_7
rlabel metal1 s 6180 0 6216 52140 4 br_0_7
rlabel metal1 s 5964 0 6000 52140 4 br_1_7
rlabel metal1 s 6444 0 6480 52140 4 bl_0_8
rlabel metal1 s 1116 19829 1152 20170 4 vdd
rlabel metal1 s 6660 0 6696 52140 4 bl_1_8
rlabel metal1 s 1116 23280 1152 23621 4 vdd
rlabel metal1 s 6516 0 6552 52140 4 br_0_8
rlabel metal1 s 1116 23779 1152 24120 4 vdd
rlabel metal1 s 6732 0 6768 52140 4 br_1_8
rlabel metal1 s 7500 0 7536 52140 4 bl_0_9
rlabel metal1 s 7284 0 7320 52140 4 bl_1_9
rlabel metal1 s 7428 0 7464 52140 4 br_0_9
rlabel metal1 s 7212 0 7248 52140 4 br_1_9
rlabel metal1 s 1116 24569 1152 24910 4 vdd
rlabel metal1 s 1116 25359 1152 25700 4 vdd
rlabel metal1 s 7692 0 7728 52140 4 bl_0_10
rlabel metal1 s 1116 24860 1152 25201 4 vdd
rlabel metal1 s 7908 0 7944 52140 4 bl_1_10
rlabel metal1 s 7764 0 7800 52140 4 br_0_10
rlabel metal1 s 7980 0 8016 52140 4 br_1_10
rlabel metal1 s 8748 0 8784 52140 4 bl_0_11
rlabel metal1 s 8532 0 8568 52140 4 bl_1_11
rlabel metal1 s 8676 0 8712 52140 4 br_0_11
rlabel metal1 s 8460 0 8496 52140 4 br_1_11
rlabel metal1 s 8940 0 8976 52140 4 bl_0_12
rlabel metal1 s 9156 0 9192 52140 4 bl_1_12
rlabel metal1 s 9012 0 9048 52140 4 br_0_12
rlabel metal1 s 9228 0 9264 52140 4 br_1_12
rlabel metal1 s 9996 0 10032 52140 4 bl_0_13
rlabel metal1 s 9780 0 9816 52140 4 bl_1_13
rlabel metal1 s 9924 0 9960 52140 4 br_0_13
rlabel metal1 s 9708 0 9744 52140 4 br_1_13
rlabel metal1 s 10188 0 10224 52140 4 bl_0_14
rlabel metal1 s 10404 0 10440 52140 4 bl_1_14
rlabel metal1 s 1260 0 1296 52140 4 rbl_bl_0_0
rlabel metal1 s 10260 0 10296 52140 4 br_0_14
rlabel metal1 s 1116 21700 1152 22041 4 vdd
rlabel metal1 s 1044 0 1080 52140 4 rbl_bl_1_0
rlabel metal1 s 10476 0 10512 52140 4 br_1_14
rlabel metal1 s 1188 0 1224 52140 4 rbl_br_0_0
rlabel metal1 s 972 0 1008 52140 4 rbl_br_1_0
rlabel metal1 s 1116 14590 1152 14931 4 vdd
rlabel metal1 s 1116 13800 1152 14141 4 vdd
rlabel metal1 s 1116 17750 1152 18091 4 vdd
rlabel metal1 s 1116 16170 1152 16511 4 vdd
rlabel metal1 s 1116 14299 1152 14640 4 vdd
rlabel metal1 s 1116 19039 1152 19380 4 vdd
rlabel metal1 s 1116 16669 1152 17010 4 vdd
rlabel metal1 s 1116 16960 1152 17301 4 vdd
rlabel metal1 s 1116 13509 1152 13850 4 vdd
rlabel metal1 s 1116 18249 1152 18590 4 vdd
rlabel metal1 s 1116 15380 1152 15721 4 vdd
rlabel metal1 s 1116 15089 1152 15430 4 vdd
rlabel metal1 s 1116 17459 1152 17800 4 vdd
rlabel metal1 s 1116 19330 1152 19671 4 vdd
rlabel metal1 s 1116 18540 1152 18881 4 vdd
rlabel metal1 s 1116 15879 1152 16220 4 vdd
rlabel metal1 s 1116 5609 1152 5950 4 vdd
rlabel metal1 s 1116 3239 1152 3580 4 vdd
rlabel metal1 s 1116 3530 1152 3871 4 vdd
rlabel metal1 s 1116 1659 1152 2000 4 vdd
rlabel metal1 s 1116 5900 1152 6241 4 vdd
rlabel metal1 s 1116 4320 1152 4661 4 vdd
rlabel metal1 s 1116 1950 1152 2291 4 vdd
rlabel metal1 s 1116 2740 1152 3081 4 vdd
rlabel metal1 s 1116 869 1152 1210 4 vdd
rlabel metal1 s 1116 10640 1152 10981 4 vdd
rlabel metal1 s 1116 4029 1152 4370 4 vdd
rlabel metal1 s 1116 5110 1152 5451 4 vdd
rlabel metal1 s 1116 1160 1152 1501 4 vdd
rlabel metal1 s 1116 13010 1152 13351 4 vdd
rlabel metal1 s 1116 8769 1152 9110 4 vdd
rlabel metal1 s 1116 10349 1152 10690 4 vdd
rlabel metal1 s 1116 7979 1152 8320 4 vdd
rlabel metal1 s 1116 9850 1152 10191 4 vdd
rlabel metal1 s 1116 11430 1152 11771 4 vdd
rlabel metal1 s 1116 11929 1152 12270 4 vdd
rlabel metal1 s 1116 7189 1152 7530 4 vdd
rlabel metal1 s 1116 12220 1152 12561 4 vdd
rlabel metal1 s 1116 11139 1152 11480 4 vdd
rlabel metal1 s 1116 370 1152 711 4 vdd
rlabel metal1 s 1116 4819 1152 5160 4 vdd
rlabel metal1 s 1116 7480 1152 7821 4 vdd
rlabel metal1 s 1116 9559 1152 9900 4 vdd
rlabel metal1 s 1116 2449 1152 2790 4 vdd
rlabel metal1 s 1116 12719 1152 13060 4 vdd
rlabel metal1 s 1116 9060 1152 9401 4 vdd
rlabel metal1 s 1116 6399 1152 6740 4 vdd
rlabel metal1 s 1116 6690 1152 7031 4 vdd
rlabel metal1 s 1116 8270 1152 8611 4 vdd
rlabel metal1 s 72108 0 72144 52140 4 br_1_113
rlabel metal1 s 72588 0 72624 52140 4 bl_0_114
rlabel metal1 s 72804 0 72840 52140 4 bl_1_114
rlabel metal1 s 72660 0 72696 52140 4 br_0_114
rlabel metal1 s 72876 0 72912 52140 4 br_1_114
rlabel metal1 s 73644 0 73680 52140 4 bl_0_115
rlabel metal1 s 73428 0 73464 52140 4 bl_1_115
rlabel metal1 s 73572 0 73608 52140 4 br_0_115
rlabel metal1 s 73356 0 73392 52140 4 br_1_115
rlabel metal1 s 73836 0 73872 52140 4 bl_0_116
rlabel metal1 s 74052 0 74088 52140 4 bl_1_116
rlabel metal1 s 73908 0 73944 52140 4 br_0_116
rlabel metal1 s 74124 0 74160 52140 4 br_1_116
rlabel metal1 s 74892 0 74928 52140 4 bl_0_117
rlabel metal1 s 74676 0 74712 52140 4 bl_1_117
rlabel metal1 s 74820 0 74856 52140 4 br_0_117
rlabel metal1 s 74604 0 74640 52140 4 br_1_117
rlabel metal1 s 75084 0 75120 52140 4 bl_0_118
rlabel metal1 s 75300 0 75336 52140 4 bl_1_118
rlabel metal1 s 75156 0 75192 52140 4 br_0_118
rlabel metal1 s 75372 0 75408 52140 4 br_1_118
rlabel metal1 s 76140 0 76176 52140 4 bl_0_119
rlabel metal1 s 75924 0 75960 52140 4 bl_1_119
rlabel metal1 s 76068 0 76104 52140 4 br_0_119
rlabel metal1 s 75852 0 75888 52140 4 br_1_119
rlabel metal1 s 76332 0 76368 52140 4 bl_0_120
rlabel metal1 s 76548 0 76584 52140 4 bl_1_120
rlabel metal1 s 76404 0 76440 52140 4 br_0_120
rlabel metal1 s 76620 0 76656 52140 4 br_1_120
rlabel metal1 s 77388 0 77424 52140 4 bl_0_121
rlabel metal1 s 77172 0 77208 52140 4 bl_1_121
rlabel metal1 s 77316 0 77352 52140 4 br_0_121
rlabel metal1 s 77100 0 77136 52140 4 br_1_121
rlabel metal1 s 77580 0 77616 52140 4 bl_0_122
rlabel metal1 s 77796 0 77832 52140 4 bl_1_122
rlabel metal1 s 77652 0 77688 52140 4 br_0_122
rlabel metal1 s 77868 0 77904 52140 4 br_1_122
rlabel metal1 s 78636 0 78672 52140 4 bl_0_123
rlabel metal1 s 78420 0 78456 52140 4 bl_1_123
rlabel metal1 s 78564 0 78600 52140 4 br_0_123
rlabel metal1 s 78348 0 78384 52140 4 br_1_123
rlabel metal1 s 78828 0 78864 52140 4 bl_0_124
rlabel metal1 s 79044 0 79080 52140 4 bl_1_124
rlabel metal1 s 78900 0 78936 52140 4 br_0_124
rlabel metal1 s 79116 0 79152 52140 4 br_1_124
rlabel metal1 s 79884 0 79920 52140 4 bl_0_125
rlabel metal1 s 79668 0 79704 52140 4 bl_1_125
rlabel metal1 s 79812 0 79848 52140 4 br_0_125
rlabel metal1 s 79596 0 79632 52140 4 br_1_125
rlabel metal1 s 80076 0 80112 52140 4 bl_0_126
rlabel metal1 s 80292 0 80328 52140 4 bl_1_126
rlabel metal1 s 80148 0 80184 52140 4 br_0_126
rlabel metal1 s 80364 0 80400 52140 4 br_1_126
rlabel metal1 s 81132 0 81168 52140 4 bl_0_127
rlabel metal1 s 80916 0 80952 52140 4 bl_1_127
rlabel metal1 s 81060 0 81096 52140 4 br_0_127
rlabel metal1 s 80844 0 80880 52140 4 br_1_127
rlabel metal1 s 81324 0 81360 52140 4 rbl_bl_0_1
rlabel metal1 s 81540 0 81576 52140 4 rbl_bl_1_1
rlabel metal1 s 81396 0 81432 52140 4 rbl_br_0_1
rlabel metal1 s 81612 0 81648 52140 4 rbl_br_1_1
rlabel metal1 s 81468 19829 81504 20170 4 vdd
rlabel metal1 s 81468 23280 81504 23621 4 vdd
rlabel metal1 s 81468 21409 81504 21750 4 vdd
rlabel metal1 s 81468 20910 81504 21251 4 vdd
rlabel metal1 s 81468 22490 81504 22831 4 vdd
rlabel metal1 s 81468 21700 81504 22041 4 vdd
rlabel metal1 s 81468 23779 81504 24120 4 vdd
rlabel metal1 s 81468 20619 81504 20960 4 vdd
rlabel metal1 s 81468 22199 81504 22540 4 vdd
rlabel metal1 s 81468 24070 81504 24411 4 vdd
rlabel metal1 s 81468 22989 81504 23330 4 vdd
rlabel metal1 s 81468 25359 81504 25700 4 vdd
rlabel metal1 s 81468 24860 81504 25201 4 vdd
rlabel metal1 s 81468 20120 81504 20461 4 vdd
rlabel metal1 s 81468 25650 81504 25991 4 vdd
rlabel metal1 s 71556 0 71592 52140 4 bl_1_112
rlabel metal1 s 81468 24569 81504 24910 4 vdd
rlabel metal1 s 71628 0 71664 52140 4 br_1_112
rlabel metal1 s 72396 0 72432 52140 4 bl_0_113
rlabel metal1 s 72180 0 72216 52140 4 bl_1_113
rlabel metal1 s 72324 0 72360 52140 4 br_0_113
rlabel metal1 s 63660 0 63696 52140 4 bl_0_99
rlabel metal1 s 63444 0 63480 52140 4 bl_1_99
rlabel metal1 s 63588 0 63624 52140 4 br_0_99
rlabel metal1 s 63372 0 63408 52140 4 br_1_99
rlabel metal1 s 63852 0 63888 52140 4 bl_0_100
rlabel metal1 s 64068 0 64104 52140 4 bl_1_100
rlabel metal1 s 63924 0 63960 52140 4 br_0_100
rlabel metal1 s 64140 0 64176 52140 4 br_1_100
rlabel metal1 s 64908 0 64944 52140 4 bl_0_101
rlabel metal1 s 64692 0 64728 52140 4 bl_1_101
rlabel metal1 s 64836 0 64872 52140 4 br_0_101
rlabel metal1 s 64620 0 64656 52140 4 br_1_101
rlabel metal1 s 65100 0 65136 52140 4 bl_0_102
rlabel metal1 s 65316 0 65352 52140 4 bl_1_102
rlabel metal1 s 65172 0 65208 52140 4 br_0_102
rlabel metal1 s 65388 0 65424 52140 4 br_1_102
rlabel metal1 s 66156 0 66192 52140 4 bl_0_103
rlabel metal1 s 65940 0 65976 52140 4 bl_1_103
rlabel metal1 s 66084 0 66120 52140 4 br_0_103
rlabel metal1 s 61572 0 61608 52140 4 bl_1_96
rlabel metal1 s 65868 0 65904 52140 4 br_1_103
rlabel metal1 s 66348 0 66384 52140 4 bl_0_104
rlabel metal1 s 66564 0 66600 52140 4 bl_1_104
rlabel metal1 s 66420 0 66456 52140 4 br_0_104
rlabel metal1 s 66636 0 66672 52140 4 br_1_104
rlabel metal1 s 67404 0 67440 52140 4 bl_0_105
rlabel metal1 s 67188 0 67224 52140 4 bl_1_105
rlabel metal1 s 67332 0 67368 52140 4 br_0_105
rlabel metal1 s 67116 0 67152 52140 4 br_1_105
rlabel metal1 s 67596 0 67632 52140 4 bl_0_106
rlabel metal1 s 61644 0 61680 52140 4 br_1_96
rlabel metal1 s 67812 0 67848 52140 4 bl_1_106
rlabel metal1 s 62412 0 62448 52140 4 bl_0_97
rlabel metal1 s 67668 0 67704 52140 4 br_0_106
rlabel metal1 s 67884 0 67920 52140 4 br_1_106
rlabel metal1 s 68652 0 68688 52140 4 bl_0_107
rlabel metal1 s 68436 0 68472 52140 4 bl_1_107
rlabel metal1 s 68580 0 68616 52140 4 br_0_107
rlabel metal1 s 68364 0 68400 52140 4 br_1_107
rlabel metal1 s 68844 0 68880 52140 4 bl_0_108
rlabel metal1 s 69060 0 69096 52140 4 bl_1_108
rlabel metal1 s 68916 0 68952 52140 4 br_0_108
rlabel metal1 s 69132 0 69168 52140 4 br_1_108
rlabel metal1 s 69900 0 69936 52140 4 bl_0_109
rlabel metal1 s 69684 0 69720 52140 4 bl_1_109
rlabel metal1 s 69828 0 69864 52140 4 br_0_109
rlabel metal1 s 69612 0 69648 52140 4 br_1_109
rlabel metal1 s 70092 0 70128 52140 4 bl_0_110
rlabel metal1 s 70308 0 70344 52140 4 bl_1_110
rlabel metal1 s 70164 0 70200 52140 4 br_0_110
rlabel metal1 s 62196 0 62232 52140 4 bl_1_97
rlabel metal1 s 70380 0 70416 52140 4 br_1_110
rlabel metal1 s 71148 0 71184 52140 4 bl_0_111
rlabel metal1 s 70932 0 70968 52140 4 bl_1_111
rlabel metal1 s 71076 0 71112 52140 4 br_0_111
rlabel metal1 s 70860 0 70896 52140 4 br_1_111
rlabel metal1 s 71340 0 71376 52140 4 bl_0_112
rlabel metal1 s 62340 0 62376 52140 4 br_0_97
rlabel metal1 s 62124 0 62160 52140 4 br_1_97
rlabel metal1 s 71412 0 71448 52140 4 br_0_112
rlabel metal1 s 62604 0 62640 52140 4 bl_0_98
rlabel metal1 s 62820 0 62856 52140 4 bl_1_98
rlabel metal1 s 62676 0 62712 52140 4 br_0_98
rlabel metal1 s 62892 0 62928 52140 4 br_1_98
rlabel metal1 s 81468 18249 81504 18590 4 vdd
rlabel metal1 s 81468 13509 81504 13850 4 vdd
rlabel metal1 s 81468 13800 81504 14141 4 vdd
rlabel metal1 s 81468 19039 81504 19380 4 vdd
rlabel metal1 s 81468 17459 81504 17800 4 vdd
rlabel metal1 s 81468 15089 81504 15430 4 vdd
rlabel metal1 s 81468 16960 81504 17301 4 vdd
rlabel metal1 s 81468 15380 81504 15721 4 vdd
rlabel metal1 s 81468 14299 81504 14640 4 vdd
rlabel metal1 s 81468 18540 81504 18881 4 vdd
rlabel metal1 s 81468 16669 81504 17010 4 vdd
rlabel metal1 s 81468 15879 81504 16220 4 vdd
rlabel metal1 s 81468 16170 81504 16511 4 vdd
rlabel metal1 s 81468 14590 81504 14931 4 vdd
rlabel metal1 s 81468 19330 81504 19671 4 vdd
rlabel metal1 s 81468 17750 81504 18091 4 vdd
rlabel metal1 s 54924 0 54960 52140 4 bl_0_85
rlabel metal1 s 54708 0 54744 52140 4 bl_1_85
rlabel metal1 s 54852 0 54888 52140 4 br_0_85
rlabel metal1 s 54636 0 54672 52140 4 br_1_85
rlabel metal1 s 55116 0 55152 52140 4 bl_0_86
rlabel metal1 s 55332 0 55368 52140 4 bl_1_86
rlabel metal1 s 55188 0 55224 52140 4 br_0_86
rlabel metal1 s 55404 0 55440 52140 4 br_1_86
rlabel metal1 s 56172 0 56208 52140 4 bl_0_87
rlabel metal1 s 55956 0 55992 52140 4 bl_1_87
rlabel metal1 s 56100 0 56136 52140 4 br_0_87
rlabel metal1 s 55884 0 55920 52140 4 br_1_87
rlabel metal1 s 56364 0 56400 52140 4 bl_0_88
rlabel metal1 s 56580 0 56616 52140 4 bl_1_88
rlabel metal1 s 56436 0 56472 52140 4 br_0_88
rlabel metal1 s 56652 0 56688 52140 4 br_1_88
rlabel metal1 s 57420 0 57456 52140 4 bl_0_89
rlabel metal1 s 57204 0 57240 52140 4 bl_1_89
rlabel metal1 s 57348 0 57384 52140 4 br_0_89
rlabel metal1 s 57132 0 57168 52140 4 br_1_89
rlabel metal1 s 57612 0 57648 52140 4 bl_0_90
rlabel metal1 s 57828 0 57864 52140 4 bl_1_90
rlabel metal1 s 57684 0 57720 52140 4 br_0_90
rlabel metal1 s 57900 0 57936 52140 4 br_1_90
rlabel metal1 s 58668 0 58704 52140 4 bl_0_91
rlabel metal1 s 58452 0 58488 52140 4 bl_1_91
rlabel metal1 s 58596 0 58632 52140 4 br_0_91
rlabel metal1 s 58380 0 58416 52140 4 br_1_91
rlabel metal1 s 58860 0 58896 52140 4 bl_0_92
rlabel metal1 s 59076 0 59112 52140 4 bl_1_92
rlabel metal1 s 58932 0 58968 52140 4 br_0_92
rlabel metal1 s 59148 0 59184 52140 4 br_1_92
rlabel metal1 s 59916 0 59952 52140 4 bl_0_93
rlabel metal1 s 59700 0 59736 52140 4 bl_1_93
rlabel metal1 s 59844 0 59880 52140 4 br_0_93
rlabel metal1 s 59628 0 59664 52140 4 br_1_93
rlabel metal1 s 60108 0 60144 52140 4 bl_0_94
rlabel metal1 s 60324 0 60360 52140 4 bl_1_94
rlabel metal1 s 60180 0 60216 52140 4 br_0_94
rlabel metal1 s 60396 0 60432 52140 4 br_1_94
rlabel metal1 s 61164 0 61200 52140 4 bl_0_95
rlabel metal1 s 60948 0 60984 52140 4 bl_1_95
rlabel metal1 s 61092 0 61128 52140 4 br_0_95
rlabel metal1 s 60876 0 60912 52140 4 br_1_95
rlabel metal1 s 61356 0 61392 52140 4 bl_0_96
rlabel metal1 s 61428 0 61464 52140 4 br_0_96
rlabel metal1 s 51588 0 51624 52140 4 bl_1_80
rlabel metal1 s 51444 0 51480 52140 4 br_0_80
rlabel metal1 s 51660 0 51696 52140 4 br_1_80
rlabel metal1 s 52428 0 52464 52140 4 bl_0_81
rlabel metal1 s 52212 0 52248 52140 4 bl_1_81
rlabel metal1 s 52356 0 52392 52140 4 br_0_81
rlabel metal1 s 52140 0 52176 52140 4 br_1_81
rlabel metal1 s 52620 0 52656 52140 4 bl_0_82
rlabel metal1 s 52836 0 52872 52140 4 bl_1_82
rlabel metal1 s 52692 0 52728 52140 4 br_0_82
rlabel metal1 s 52908 0 52944 52140 4 br_1_82
rlabel metal1 s 53676 0 53712 52140 4 bl_0_83
rlabel metal1 s 53460 0 53496 52140 4 bl_1_83
rlabel metal1 s 53604 0 53640 52140 4 br_0_83
rlabel metal1 s 53388 0 53424 52140 4 br_1_83
rlabel metal1 s 53868 0 53904 52140 4 bl_0_84
rlabel metal1 s 54084 0 54120 52140 4 bl_1_84
rlabel metal1 s 53940 0 53976 52140 4 br_0_84
rlabel metal1 s 54156 0 54192 52140 4 br_1_84
rlabel metal1 s 45420 0 45456 52140 4 br_1_70
rlabel metal1 s 46188 0 46224 52140 4 bl_0_71
rlabel metal1 s 45972 0 46008 52140 4 bl_1_71
rlabel metal1 s 42852 0 42888 52140 4 bl_1_66
rlabel metal1 s 46116 0 46152 52140 4 br_0_71
rlabel metal1 s 45900 0 45936 52140 4 br_1_71
rlabel metal1 s 46380 0 46416 52140 4 bl_0_72
rlabel metal1 s 46596 0 46632 52140 4 bl_1_72
rlabel metal1 s 46452 0 46488 52140 4 br_0_72
rlabel metal1 s 46668 0 46704 52140 4 br_1_72
rlabel metal1 s 47436 0 47472 52140 4 bl_0_73
rlabel metal1 s 47220 0 47256 52140 4 bl_1_73
rlabel metal1 s 47364 0 47400 52140 4 br_0_73
rlabel metal1 s 47148 0 47184 52140 4 br_1_73
rlabel metal1 s 47628 0 47664 52140 4 bl_0_74
rlabel metal1 s 47844 0 47880 52140 4 bl_1_74
rlabel metal1 s 47700 0 47736 52140 4 br_0_74
rlabel metal1 s 41388 0 41424 52140 4 bl_0_64
rlabel metal1 s 47916 0 47952 52140 4 br_1_74
rlabel metal1 s 48684 0 48720 52140 4 bl_0_75
rlabel metal1 s 48468 0 48504 52140 4 bl_1_75
rlabel metal1 s 41604 0 41640 52140 4 bl_1_64
rlabel metal1 s 48612 0 48648 52140 4 br_0_75
rlabel metal1 s 48396 0 48432 52140 4 br_1_75
rlabel metal1 s 48876 0 48912 52140 4 bl_0_76
rlabel metal1 s 49092 0 49128 52140 4 bl_1_76
rlabel metal1 s 42708 0 42744 52140 4 br_0_66
rlabel metal1 s 42924 0 42960 52140 4 br_1_66
rlabel metal1 s 48948 0 48984 52140 4 br_0_76
rlabel metal1 s 49164 0 49200 52140 4 br_1_76
rlabel metal1 s 49932 0 49968 52140 4 bl_0_77
rlabel metal1 s 49716 0 49752 52140 4 bl_1_77
rlabel metal1 s 49860 0 49896 52140 4 br_0_77
rlabel metal1 s 43692 0 43728 52140 4 bl_0_67
rlabel metal1 s 49644 0 49680 52140 4 br_1_77
rlabel metal1 s 50124 0 50160 52140 4 bl_0_78
rlabel metal1 s 50340 0 50376 52140 4 bl_1_78
rlabel metal1 s 43476 0 43512 52140 4 bl_1_67
rlabel metal1 s 50196 0 50232 52140 4 br_0_78
rlabel metal1 s 50412 0 50448 52140 4 br_1_78
rlabel metal1 s 51180 0 51216 52140 4 bl_0_79
rlabel metal1 s 50964 0 51000 52140 4 bl_1_79
rlabel metal1 s 51108 0 51144 52140 4 br_0_79
rlabel metal1 s 50892 0 50928 52140 4 br_1_79
rlabel metal1 s 51372 0 51408 52140 4 bl_0_80
rlabel metal1 s 44100 0 44136 52140 4 bl_1_68
rlabel metal1 s 43404 0 43440 52140 4 br_1_67
rlabel metal1 s 42444 0 42480 52140 4 bl_0_65
rlabel metal1 s 43884 0 43920 52140 4 bl_0_68
rlabel metal1 s 41676 0 41712 52140 4 br_1_64
rlabel metal1 s 42228 0 42264 52140 4 bl_1_65
rlabel metal1 s 43956 0 43992 52140 4 br_0_68
rlabel metal1 s 41460 0 41496 52140 4 br_0_64
rlabel metal1 s 43620 0 43656 52140 4 br_0_67
rlabel metal1 s 44172 0 44208 52140 4 br_1_68
rlabel metal1 s 42372 0 42408 52140 4 br_0_65
rlabel metal1 s 44940 0 44976 52140 4 bl_0_69
rlabel metal1 s 44724 0 44760 52140 4 bl_1_69
rlabel metal1 s 44868 0 44904 52140 4 br_0_69
rlabel metal1 s 44652 0 44688 52140 4 br_1_69
rlabel metal1 s 42156 0 42192 52140 4 br_1_65
rlabel metal1 s 45132 0 45168 52140 4 bl_0_70
rlabel metal1 s 45348 0 45384 52140 4 bl_1_70
rlabel metal1 s 45204 0 45240 52140 4 br_0_70
rlabel metal1 s 42636 0 42672 52140 4 bl_0_66
rlabel metal1 s 81468 869 81504 1210 4 vdd
rlabel metal1 s 81468 7979 81504 8320 4 vdd
rlabel metal1 s 81468 370 81504 711 4 vdd
rlabel metal1 s 81468 9060 81504 9401 4 vdd
rlabel metal1 s 81468 7480 81504 7821 4 vdd
rlabel metal1 s 81468 1950 81504 2291 4 vdd
rlabel metal1 s 81468 12220 81504 12561 4 vdd
rlabel metal1 s 81468 8769 81504 9110 4 vdd
rlabel metal1 s 81468 1659 81504 2000 4 vdd
rlabel metal1 s 81468 3530 81504 3871 4 vdd
rlabel metal1 s 81468 9850 81504 10191 4 vdd
rlabel metal1 s 81468 4819 81504 5160 4 vdd
rlabel metal1 s 81468 7189 81504 7530 4 vdd
rlabel metal1 s 81468 1160 81504 1501 4 vdd
rlabel metal1 s 81468 6690 81504 7031 4 vdd
rlabel metal1 s 81468 5900 81504 6241 4 vdd
rlabel metal1 s 81468 12719 81504 13060 4 vdd
rlabel metal1 s 81468 11139 81504 11480 4 vdd
rlabel metal1 s 81468 10349 81504 10690 4 vdd
rlabel metal1 s 81468 8270 81504 8611 4 vdd
rlabel metal1 s 81468 5609 81504 5950 4 vdd
rlabel metal1 s 81468 9559 81504 9900 4 vdd
rlabel metal1 s 81468 5110 81504 5451 4 vdd
rlabel metal1 s 81468 6399 81504 6740 4 vdd
rlabel metal1 s 81468 11430 81504 11771 4 vdd
rlabel metal1 s 81468 4320 81504 4661 4 vdd
rlabel metal1 s 81468 2449 81504 2790 4 vdd
rlabel metal1 s 81468 11929 81504 12270 4 vdd
rlabel metal1 s 81468 10640 81504 10981 4 vdd
rlabel metal1 s 81468 3239 81504 3580 4 vdd
rlabel metal1 s 81468 4029 81504 4370 4 vdd
rlabel metal1 s 81468 2740 81504 3081 4 vdd
rlabel metal1 s 81468 13010 81504 13351 4 vdd
<< properties >>
string FIXED_BBOX 0 0 82620 52140
<< end >>
