* Clock divider test

vclk clk 0 pulse(0 1.8 50p 2p 2p 50p 100p)
vvdd vdd 0 dc 1.8

Aadc [clk] [clk_digital] myadc
.model myadc adc_bridge(in_low = 0.9 in_high = 0.9 rise_delay = 10e-12 fall_delay = 10e-12)

Adiv clk_digital clk_div_digital myclkdiv
.model myclkdiv d_fdiv(div_factor = 16 high_cycles = 8 rise_delay = 10e-12 fall_delay = 10e-12)

Adac [clk_div_digital] [clk_div] mydac
.model mydac dac_bridge(out_low = 0 out_high = 1.8 t_rise = 10e-12 t_fall = 10e-12)

cout clk_div 0 1e-12

.control
save all
tran 1p 2n
write clk_divider_test_tran.raw
.endc