magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< metal3 >>
rect -1550 194 1549 300
rect -1550 -272 1465 194
rect 1529 -272 1549 194
rect -1550 -300 1549 -272
<< via3 >>
rect 1465 -272 1529 194
<< mimcap >>
rect -1450 160 1350 200
rect -1450 -160 -1410 160
rect 1310 -160 1350 160
rect -1450 -200 1350 -160
<< mimcapcontact >>
rect -1410 -160 1310 160
<< metal4 >>
rect 1449 194 1545 234
rect -1411 160 1311 161
rect -1411 -160 -1410 160
rect 1310 -160 1311 160
rect -1411 -161 1311 -160
rect 1449 -272 1465 194
rect 1529 -272 1545 194
rect 1449 -288 1545 -272
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1550 -300 1450 300
string parameters w 14.00 l 2.00 val 62.08 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
