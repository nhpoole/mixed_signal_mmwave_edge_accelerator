magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -646 -646 646 646
<< metal1 >>
rect -13 13 13 16
rect -13 -16 13 -13
<< via1 >>
rect -13 -13 13 13
<< metal2 >>
rect -16 -13 -13 13
rect 13 -13 16 13
<< end >>
