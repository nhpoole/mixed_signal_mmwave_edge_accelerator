magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1302 -841 1884 52981
<< metal2 >>
rect 0 51199 28 51247
rect 0 50979 28 51027
rect 0 50883 28 50931
rect 0 50663 28 50711
rect 0 50409 28 50457
rect 0 50189 28 50237
rect 0 50093 28 50141
rect 0 49873 28 49921
rect 0 49619 28 49667
rect 0 49399 28 49447
rect 0 49303 28 49351
rect 0 49083 28 49131
rect 0 48829 28 48877
rect 0 48609 28 48657
rect 0 48513 28 48561
rect 0 48293 28 48341
rect 0 48039 28 48087
rect 0 47819 28 47867
rect 0 47723 28 47771
rect 0 47503 28 47551
rect 0 47249 28 47297
rect 0 47029 28 47077
rect 0 46933 28 46981
rect 0 46713 28 46761
rect 0 46459 28 46507
rect 0 46239 28 46287
rect 0 46143 28 46191
rect 0 45923 28 45971
rect 0 45669 28 45717
rect 0 45449 28 45497
rect 0 45353 28 45401
rect 0 45133 28 45181
rect 0 44879 28 44927
rect 0 44659 28 44707
rect 0 44563 28 44611
rect 0 44343 28 44391
rect 0 44089 28 44137
rect 0 43869 28 43917
rect 0 43773 28 43821
rect 0 43553 28 43601
rect 0 43299 28 43347
rect 0 43079 28 43127
rect 0 42983 28 43031
rect 0 42763 28 42811
rect 0 42509 28 42557
rect 0 42289 28 42337
rect 0 42193 28 42241
rect 0 41973 28 42021
rect 0 41719 28 41767
rect 0 41499 28 41547
rect 0 41403 28 41451
rect 0 41183 28 41231
rect 0 40929 28 40977
rect 0 40709 28 40757
rect 0 40613 28 40661
rect 0 40393 28 40441
rect 0 40139 28 40187
rect 0 39919 28 39967
rect 0 39823 28 39871
rect 0 39603 28 39651
rect 0 39349 28 39397
rect 0 39129 28 39177
rect 0 39033 28 39081
rect 0 38813 28 38861
rect 0 38559 28 38607
rect 0 38339 28 38387
rect 0 38243 28 38291
rect 0 38023 28 38071
rect 0 37769 28 37817
rect 0 37549 28 37597
rect 0 37453 28 37501
rect 0 37233 28 37281
rect 0 36979 28 37027
rect 0 36759 28 36807
rect 0 36663 28 36711
rect 0 36443 28 36491
rect 0 36189 28 36237
rect 0 35969 28 36017
rect 0 35873 28 35921
rect 0 35653 28 35701
rect 0 35399 28 35447
rect 0 35179 28 35227
rect 0 35083 28 35131
rect 0 34863 28 34911
rect 0 34609 28 34657
rect 0 34389 28 34437
rect 0 34293 28 34341
rect 0 34073 28 34121
rect 0 33819 28 33867
rect 0 33599 28 33647
rect 0 33503 28 33551
rect 0 33283 28 33331
rect 0 33029 28 33077
rect 0 32809 28 32857
rect 0 32713 28 32761
rect 0 32493 28 32541
rect 0 32239 28 32287
rect 0 32019 28 32067
rect 0 31923 28 31971
rect 0 31703 28 31751
rect 0 31449 28 31497
rect 0 31229 28 31277
rect 0 31133 28 31181
rect 0 30913 28 30961
rect 0 30659 28 30707
rect 0 30439 28 30487
rect 0 30343 28 30391
rect 0 30123 28 30171
rect 0 29869 28 29917
rect 0 29649 28 29697
rect 0 29553 28 29601
rect 0 29333 28 29381
rect 0 29079 28 29127
rect 0 28859 28 28907
rect 0 28763 28 28811
rect 0 28543 28 28591
rect 0 28289 28 28337
rect 0 28069 28 28117
rect 0 27973 28 28021
rect 0 27753 28 27801
rect 0 27499 28 27547
rect 0 27279 28 27327
rect 0 27183 28 27231
rect 0 26963 28 27011
rect 0 26709 28 26757
rect 0 26489 28 26537
rect 0 26393 28 26441
rect 0 26173 28 26221
rect 0 25919 28 25967
rect 0 25699 28 25747
rect 0 25603 28 25651
rect 0 25383 28 25431
rect 0 25129 28 25177
rect 0 24909 28 24957
rect 0 24813 28 24861
rect 0 24593 28 24641
rect 0 24339 28 24387
rect 0 24119 28 24167
rect 0 24023 28 24071
rect 0 23803 28 23851
rect 0 23549 28 23597
rect 0 23329 28 23377
rect 0 23233 28 23281
rect 0 23013 28 23061
rect 0 22759 28 22807
rect 0 22539 28 22587
rect 0 22443 28 22491
rect 0 22223 28 22271
rect 0 21969 28 22017
rect 0 21749 28 21797
rect 0 21653 28 21701
rect 0 21433 28 21481
rect 0 21179 28 21227
rect 0 20959 28 21007
rect 0 20863 28 20911
rect 0 20643 28 20691
rect 0 20389 28 20437
rect 0 20169 28 20217
rect 0 20073 28 20121
rect 0 19853 28 19901
rect 0 19599 28 19647
rect 0 19379 28 19427
rect 0 19283 28 19331
rect 0 19063 28 19111
rect 0 18809 28 18857
rect 0 18589 28 18637
rect 0 18493 28 18541
rect 0 18273 28 18321
rect 0 18019 28 18067
rect 0 17799 28 17847
rect 0 17703 28 17751
rect 0 17483 28 17531
rect 0 17229 28 17277
rect 0 17009 28 17057
rect 0 16913 28 16961
rect 0 16693 28 16741
rect 0 16439 28 16487
rect 0 16219 28 16267
rect 0 16123 28 16171
rect 0 15903 28 15951
rect 0 15649 28 15697
rect 0 15429 28 15477
rect 0 15333 28 15381
rect 0 15113 28 15161
rect 0 14859 28 14907
rect 0 14639 28 14687
rect 0 14543 28 14591
rect 0 14323 28 14371
rect 0 14069 28 14117
rect 0 13849 28 13897
rect 0 13753 28 13801
rect 0 13533 28 13581
rect 0 13279 28 13327
rect 0 13059 28 13107
rect 0 12963 28 13011
rect 0 12743 28 12791
rect 0 12489 28 12537
rect 0 12269 28 12317
rect 0 12173 28 12221
rect 0 11953 28 12001
rect 0 11699 28 11747
rect 0 11479 28 11527
rect 0 11383 28 11431
rect 0 11163 28 11211
rect 0 10909 28 10957
rect 0 10689 28 10737
rect 0 10593 28 10641
rect 0 10373 28 10421
rect 0 10119 28 10167
rect 0 9899 28 9947
rect 0 9803 28 9851
rect 0 9583 28 9631
rect 0 9329 28 9377
rect 0 9109 28 9157
rect 0 9013 28 9061
rect 0 8793 28 8841
rect 0 8539 28 8587
rect 0 8319 28 8367
rect 0 8223 28 8271
rect 0 8003 28 8051
rect 0 7749 28 7797
rect 0 7529 28 7577
rect 0 7433 28 7481
rect 0 7213 28 7261
rect 0 6959 28 7007
rect 0 6739 28 6787
rect 0 6643 28 6691
rect 0 6423 28 6471
rect 0 6169 28 6217
rect 0 5949 28 5997
rect 0 5853 28 5901
rect 0 5633 28 5681
rect 0 5379 28 5427
rect 0 5159 28 5207
rect 0 5063 28 5111
rect 0 4843 28 4891
rect 0 4589 28 4637
rect 0 4369 28 4417
rect 0 4273 28 4321
rect 0 4053 28 4101
rect 0 3799 28 3847
rect 0 3579 28 3627
rect 0 3483 28 3531
rect 0 3263 28 3311
rect 0 3009 28 3057
rect 0 2789 28 2837
rect 0 2693 28 2741
rect 0 2473 28 2521
rect 0 2219 28 2267
rect 0 1999 28 2047
rect 0 1903 28 1951
rect 0 1683 28 1731
rect 0 1429 28 1477
rect 0 1209 28 1257
rect 0 1113 28 1161
rect 0 893 28 941
<< metal3 >>
rect 191 51301 289 51399
rect 191 51064 289 51162
rect 191 50748 289 50846
rect 191 50511 289 50609
rect 191 50274 289 50372
rect 191 49958 289 50056
rect 191 49721 289 49819
rect 191 49484 289 49582
rect 191 49168 289 49266
rect 191 48931 289 49029
rect 191 48694 289 48792
rect 191 48378 289 48476
rect 191 48141 289 48239
rect 191 47904 289 48002
rect 191 47588 289 47686
rect 191 47351 289 47449
rect 191 47114 289 47212
rect 191 46798 289 46896
rect 191 46561 289 46659
rect 191 46324 289 46422
rect 191 46008 289 46106
rect 191 45771 289 45869
rect 191 45534 289 45632
rect 191 45218 289 45316
rect 191 44981 289 45079
rect 191 44744 289 44842
rect 191 44428 289 44526
rect 191 44191 289 44289
rect 191 43954 289 44052
rect 191 43638 289 43736
rect 191 43401 289 43499
rect 191 43164 289 43262
rect 191 42848 289 42946
rect 191 42611 289 42709
rect 191 42374 289 42472
rect 191 42058 289 42156
rect 191 41821 289 41919
rect 191 41584 289 41682
rect 191 41268 289 41366
rect 191 41031 289 41129
rect 191 40794 289 40892
rect 191 40478 289 40576
rect 191 40241 289 40339
rect 191 40004 289 40102
rect 191 39688 289 39786
rect 191 39451 289 39549
rect 191 39214 289 39312
rect 191 38898 289 38996
rect 191 38661 289 38759
rect 191 38424 289 38522
rect 191 38108 289 38206
rect 191 37871 289 37969
rect 191 37634 289 37732
rect 191 37318 289 37416
rect 191 37081 289 37179
rect 191 36844 289 36942
rect 191 36528 289 36626
rect 191 36291 289 36389
rect 191 36054 289 36152
rect 191 35738 289 35836
rect 191 35501 289 35599
rect 191 35264 289 35362
rect 191 34948 289 35046
rect 191 34711 289 34809
rect 191 34474 289 34572
rect 191 34158 289 34256
rect 191 33921 289 34019
rect 191 33684 289 33782
rect 191 33368 289 33466
rect 191 33131 289 33229
rect 191 32894 289 32992
rect 191 32578 289 32676
rect 191 32341 289 32439
rect 191 32104 289 32202
rect 191 31788 289 31886
rect 191 31551 289 31649
rect 191 31314 289 31412
rect 191 30998 289 31096
rect 191 30761 289 30859
rect 191 30524 289 30622
rect 191 30208 289 30306
rect 191 29971 289 30069
rect 191 29734 289 29832
rect 191 29418 289 29516
rect 191 29181 289 29279
rect 191 28944 289 29042
rect 191 28628 289 28726
rect 191 28391 289 28489
rect 191 28154 289 28252
rect 191 27838 289 27936
rect 191 27601 289 27699
rect 191 27364 289 27462
rect 191 27048 289 27146
rect 191 26811 289 26909
rect 191 26574 289 26672
rect 191 26258 289 26356
rect 191 26021 289 26119
rect 191 25784 289 25882
rect 191 25468 289 25566
rect 191 25231 289 25329
rect 191 24994 289 25092
rect 191 24678 289 24776
rect 191 24441 289 24539
rect 191 24204 289 24302
rect 191 23888 289 23986
rect 191 23651 289 23749
rect 191 23414 289 23512
rect 191 23098 289 23196
rect 191 22861 289 22959
rect 191 22624 289 22722
rect 191 22308 289 22406
rect 191 22071 289 22169
rect 191 21834 289 21932
rect 191 21518 289 21616
rect 191 21281 289 21379
rect 191 21044 289 21142
rect 191 20728 289 20826
rect 191 20491 289 20589
rect 191 20254 289 20352
rect 191 19938 289 20036
rect 191 19701 289 19799
rect 191 19464 289 19562
rect 191 19148 289 19246
rect 191 18911 289 19009
rect 191 18674 289 18772
rect 191 18358 289 18456
rect 191 18121 289 18219
rect 191 17884 289 17982
rect 191 17568 289 17666
rect 191 17331 289 17429
rect 191 17094 289 17192
rect 191 16778 289 16876
rect 191 16541 289 16639
rect 191 16304 289 16402
rect 191 15988 289 16086
rect 191 15751 289 15849
rect 191 15514 289 15612
rect 191 15198 289 15296
rect 191 14961 289 15059
rect 191 14724 289 14822
rect 191 14408 289 14506
rect 191 14171 289 14269
rect 191 13934 289 14032
rect 191 13618 289 13716
rect 191 13381 289 13479
rect 191 13144 289 13242
rect 191 12828 289 12926
rect 191 12591 289 12689
rect 191 12354 289 12452
rect 191 12038 289 12136
rect 191 11801 289 11899
rect 191 11564 289 11662
rect 191 11248 289 11346
rect 191 11011 289 11109
rect 191 10774 289 10872
rect 191 10458 289 10556
rect 191 10221 289 10319
rect 191 9984 289 10082
rect 191 9668 289 9766
rect 191 9431 289 9529
rect 191 9194 289 9292
rect 191 8878 289 8976
rect 191 8641 289 8739
rect 191 8404 289 8502
rect 191 8088 289 8186
rect 191 7851 289 7949
rect 191 7614 289 7712
rect 191 7298 289 7396
rect 191 7061 289 7159
rect 191 6824 289 6922
rect 191 6508 289 6606
rect 191 6271 289 6369
rect 191 6034 289 6132
rect 191 5718 289 5816
rect 191 5481 289 5579
rect 191 5244 289 5342
rect 191 4928 289 5026
rect 191 4691 289 4789
rect 191 4454 289 4552
rect 191 4138 289 4236
rect 191 3901 289 3999
rect 191 3664 289 3762
rect 191 3348 289 3446
rect 191 3111 289 3209
rect 191 2874 289 2972
rect 191 2558 289 2656
rect 191 2321 289 2419
rect 191 2084 289 2182
rect 191 1768 289 1866
rect 191 1531 289 1629
rect 191 1294 289 1392
rect 191 978 289 1076
rect 191 741 289 839
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1626486988
transform 1 0 207 0 1 753
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_3
timestamp 1626486988
transform 1 0 0 0 1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_4
timestamp 1626486988
transform 1 0 0 0 -1 790
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1626486988
transform 1 0 207 0 1 990
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_6
timestamp 1626486988
transform 1 0 0 0 -1 1580
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1626486988
transform 1 0 207 0 1 1306
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1626486988
transform 1 0 207 0 1 1543
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1626486988
transform 1 0 207 0 1 1543
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_5
timestamp 1626486988
transform 1 0 0 0 1 1580
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1626486988
transform 1 0 207 0 1 1780
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1626486988
transform 1 0 207 0 1 2096
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_2
timestamp 1626486988
transform 1 0 0 0 -1 2370
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1626486988
transform 1 0 207 0 1 2333
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1626486988
transform 1 0 207 0 1 2333
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_1
timestamp 1626486988
transform 1 0 0 0 1 2370
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1626486988
transform 1 0 207 0 1 2570
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1626486988
transform 1 0 207 0 1 2886
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_0
timestamp 1626486988
transform 1 0 0 0 -1 3160
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1626486988
transform 1 0 207 0 1 3123
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1626486988
transform 1 0 207 0 1 3360
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1626486988
transform 1 0 207 0 1 3123
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_31
timestamp 1626486988
transform 1 0 0 0 1 3160
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1626486988
transform 1 0 207 0 1 3676
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_30
timestamp 1626486988
transform 1 0 0 0 -1 3950
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1626486988
transform 1 0 207 0 1 3913
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1626486988
transform 1 0 207 0 1 4150
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1626486988
transform 1 0 207 0 1 3913
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_29
timestamp 1626486988
transform 1 0 0 0 1 3950
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1626486988
transform 1 0 207 0 1 4466
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_27
timestamp 1626486988
transform 1 0 0 0 1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_28
timestamp 1626486988
transform 1 0 0 0 -1 4740
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1626486988
transform 1 0 207 0 1 4703
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1626486988
transform 1 0 207 0 1 4940
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1626486988
transform 1 0 207 0 1 4703
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1626486988
transform 1 0 207 0 1 5256
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1626486988
transform 1 0 207 0 1 5493
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1626486988
transform 1 0 207 0 1 5493
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_25
timestamp 1626486988
transform 1 0 0 0 1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_26
timestamp 1626486988
transform 1 0 0 0 -1 5530
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1626486988
transform 1 0 207 0 1 5730
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_24
timestamp 1626486988
transform 1 0 0 0 -1 6320
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1626486988
transform 1 0 207 0 1 6046
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1626486988
transform 1 0 207 0 1 6283
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1626486988
transform 1 0 207 0 1 6283
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_23
timestamp 1626486988
transform 1 0 0 0 1 6320
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1626486988
transform 1 0 207 0 1 6520
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_22
timestamp 1626486988
transform 1 0 0 0 -1 7110
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1626486988
transform 1 0 207 0 1 6836
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1626486988
transform 1 0 207 0 1 7073
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1626486988
transform 1 0 207 0 1 7073
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_21
timestamp 1626486988
transform 1 0 0 0 1 7110
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1626486988
transform 1 0 207 0 1 7310
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1626486988
transform 1 0 207 0 1 7626
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_20
timestamp 1626486988
transform 1 0 0 0 -1 7900
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1626486988
transform 1 0 207 0 1 7863
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1626486988
transform 1 0 207 0 1 8100
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1626486988
transform 1 0 207 0 1 7863
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_19
timestamp 1626486988
transform 1 0 0 0 1 7900
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1626486988
transform 1 0 207 0 1 8416
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_18
timestamp 1626486988
transform 1 0 0 0 -1 8690
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1626486988
transform 1 0 207 0 1 8653
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1626486988
transform 1 0 207 0 1 8890
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1626486988
transform 1 0 207 0 1 8653
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_17
timestamp 1626486988
transform 1 0 0 0 1 8690
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1626486988
transform 1 0 207 0 1 9206
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_16
timestamp 1626486988
transform 1 0 0 0 -1 9480
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1626486988
transform 1 0 207 0 1 9443
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1626486988
transform 1 0 207 0 1 9680
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626486988
transform 1 0 207 0 1 9443
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_15
timestamp 1626486988
transform 1 0 0 0 1 9480
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626486988
transform 1 0 207 0 1 9996
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626486988
transform 1 0 207 0 1 10233
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626486988
transform 1 0 207 0 1 10233
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_13
timestamp 1626486988
transform 1 0 0 0 1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_14
timestamp 1626486988
transform 1 0 0 0 -1 10270
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626486988
transform 1 0 207 0 1 10470
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626486988
transform 1 0 207 0 1 10786
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626486988
transform 1 0 207 0 1 11023
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626486988
transform 1 0 207 0 1 11023
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_11
timestamp 1626486988
transform 1 0 0 0 1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_12
timestamp 1626486988
transform 1 0 0 0 -1 11060
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626486988
transform 1 0 207 0 1 11260
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_10
timestamp 1626486988
transform 1 0 0 0 -1 11850
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626486988
transform 1 0 207 0 1 11576
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626486988
transform 1 0 207 0 1 11813
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626486988
transform 1 0 207 0 1 11813
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_9
timestamp 1626486988
transform 1 0 0 0 1 11850
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626486988
transform 1 0 207 0 1 12050
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626486988
transform 1 0 207 0 1 12366
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_8
timestamp 1626486988
transform 1 0 0 0 -1 12640
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626486988
transform 1 0 207 0 1 12603
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626486988
transform 1 0 207 0 1 12603
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_7
timestamp 1626486988
transform 1 0 0 0 1 12640
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1626486988
transform 1 0 207 0 1 13156
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626486988
transform 1 0 207 0 1 12840
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_63
timestamp 1626486988
transform 1 0 0 0 -1 13430
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1626486988
transform 1 0 207 0 1 13393
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1626486988
transform 1 0 207 0 1 13393
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1626486988
transform 1 0 207 0 1 13630
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_62
timestamp 1626486988
transform 1 0 0 0 1 13430
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1626486988
transform 1 0 207 0 1 13946
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_61
timestamp 1626486988
transform 1 0 0 0 -1 14220
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1626486988
transform 1 0 207 0 1 14183
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1626486988
transform 1 0 207 0 1 14420
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1626486988
transform 1 0 207 0 1 14183
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_60
timestamp 1626486988
transform 1 0 0 0 1 14220
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1626486988
transform 1 0 207 0 1 14736
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_59
timestamp 1626486988
transform 1 0 0 0 -1 15010
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1626486988
transform 1 0 207 0 1 14973
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1626486988
transform 1 0 207 0 1 15210
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1626486988
transform 1 0 207 0 1 14973
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_58
timestamp 1626486988
transform 1 0 0 0 1 15010
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1626486988
transform 1 0 207 0 1 15526
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1626486988
transform 1 0 207 0 1 15763
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1626486988
transform 1 0 207 0 1 15763
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_56
timestamp 1626486988
transform 1 0 0 0 1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_57
timestamp 1626486988
transform 1 0 0 0 -1 15800
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1626486988
transform 1 0 207 0 1 16000
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1626486988
transform 1 0 207 0 1 16316
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1626486988
transform 1 0 207 0 1 16553
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1626486988
transform 1 0 207 0 1 16553
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_54
timestamp 1626486988
transform 1 0 0 0 1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_55
timestamp 1626486988
transform 1 0 0 0 -1 16590
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1626486988
transform 1 0 207 0 1 16790
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_53
timestamp 1626486988
transform 1 0 0 0 -1 17380
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1626486988
transform 1 0 207 0 1 17106
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1626486988
transform 1 0 207 0 1 17343
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1626486988
transform 1 0 207 0 1 17343
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_52
timestamp 1626486988
transform 1 0 0 0 1 17380
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1626486988
transform 1 0 207 0 1 17580
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1626486988
transform 1 0 207 0 1 17896
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_51
timestamp 1626486988
transform 1 0 0 0 -1 18170
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1626486988
transform 1 0 207 0 1 18133
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1626486988
transform 1 0 207 0 1 18133
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_50
timestamp 1626486988
transform 1 0 0 0 1 18170
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1626486988
transform 1 0 207 0 1 18370
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1626486988
transform 1 0 207 0 1 18686
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_49
timestamp 1626486988
transform 1 0 0 0 -1 18960
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1626486988
transform 1 0 207 0 1 18923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1626486988
transform 1 0 207 0 1 19160
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1626486988
transform 1 0 207 0 1 18923
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_48
timestamp 1626486988
transform 1 0 0 0 1 18960
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1626486988
transform 1 0 207 0 1 19476
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_47
timestamp 1626486988
transform 1 0 0 0 -1 19750
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1626486988
transform 1 0 207 0 1 19713
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1626486988
transform 1 0 207 0 1 19950
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1626486988
transform 1 0 207 0 1 19713
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_46
timestamp 1626486988
transform 1 0 0 0 1 19750
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1626486988
transform 1 0 207 0 1 20266
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_44
timestamp 1626486988
transform 1 0 0 0 1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_45
timestamp 1626486988
transform 1 0 0 0 -1 20540
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1626486988
transform 1 0 207 0 1 20503
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1626486988
transform 1 0 207 0 1 20740
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1626486988
transform 1 0 207 0 1 20503
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1626486988
transform 1 0 207 0 1 21056
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1626486988
transform 1 0 207 0 1 21293
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1626486988
transform 1 0 207 0 1 21293
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_42
timestamp 1626486988
transform 1 0 0 0 1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_43
timestamp 1626486988
transform 1 0 0 0 -1 21330
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1626486988
transform 1 0 207 0 1 21530
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_41
timestamp 1626486988
transform 1 0 0 0 -1 22120
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1626486988
transform 1 0 207 0 1 21846
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1626486988
transform 1 0 207 0 1 22083
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1626486988
transform 1 0 207 0 1 22083
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_40
timestamp 1626486988
transform 1 0 0 0 1 22120
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1626486988
transform 1 0 207 0 1 22320
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_39
timestamp 1626486988
transform 1 0 0 0 -1 22910
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1626486988
transform 1 0 207 0 1 22636
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1626486988
transform 1 0 207 0 1 22873
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1626486988
transform 1 0 207 0 1 22873
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_38
timestamp 1626486988
transform 1 0 0 0 1 22910
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1626486988
transform 1 0 207 0 1 23110
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1626486988
transform 1 0 207 0 1 23426
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_37
timestamp 1626486988
transform 1 0 0 0 -1 23700
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1626486988
transform 1 0 207 0 1 23663
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1626486988
transform 1 0 207 0 1 23900
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1626486988
transform 1 0 207 0 1 23663
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_36
timestamp 1626486988
transform 1 0 0 0 1 23700
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1626486988
transform 1 0 207 0 1 24216
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_35
timestamp 1626486988
transform 1 0 0 0 -1 24490
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1626486988
transform 1 0 207 0 1 24453
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1626486988
transform 1 0 207 0 1 24690
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1626486988
transform 1 0 207 0 1 24453
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_34
timestamp 1626486988
transform 1 0 0 0 1 24490
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1626486988
transform 1 0 207 0 1 25006
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_33
timestamp 1626486988
transform 1 0 0 0 -1 25280
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1626486988
transform 1 0 207 0 1 25243
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1626486988
transform 1 0 207 0 1 25480
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1626486988
transform 1 0 207 0 1 25243
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_32
timestamp 1626486988
transform 1 0 0 0 1 25280
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_255
timestamp 1626486988
transform 1 0 207 0 1 26033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_254
timestamp 1626486988
transform 1 0 207 0 1 26033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1626486988
transform 1 0 207 0 1 25796
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_128
timestamp 1626486988
transform 1 0 0 0 1 26070
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_129
timestamp 1626486988
transform 1 0 0 0 -1 26070
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_158
timestamp 1626486988
transform 1 0 207 0 1 26270
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_157
timestamp 1626486988
transform 1 0 207 0 1 26586
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_156
timestamp 1626486988
transform 1 0 207 0 1 26823
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_154
timestamp 1626486988
transform 1 0 207 0 1 26823
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_64
timestamp 1626486988
transform 1 0 0 0 1 26860
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_65
timestamp 1626486988
transform 1 0 0 0 -1 26860
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_155
timestamp 1626486988
transform 1 0 207 0 1 27060
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_69
timestamp 1626486988
transform 1 0 0 0 -1 27650
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_153
timestamp 1626486988
transform 1 0 207 0 1 27376
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_152
timestamp 1626486988
transform 1 0 207 0 1 27613
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_150
timestamp 1626486988
transform 1 0 207 0 1 27613
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_68
timestamp 1626486988
transform 1 0 0 0 1 27650
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_151
timestamp 1626486988
transform 1 0 207 0 1 27850
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_149
timestamp 1626486988
transform 1 0 207 0 1 28166
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_67
timestamp 1626486988
transform 1 0 0 0 -1 28440
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_148
timestamp 1626486988
transform 1 0 207 0 1 28403
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_146
timestamp 1626486988
transform 1 0 207 0 1 28403
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_66
timestamp 1626486988
transform 1 0 0 0 1 28440
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_147
timestamp 1626486988
transform 1 0 207 0 1 28640
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_145
timestamp 1626486988
transform 1 0 207 0 1 28956
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_94
timestamp 1626486988
transform 1 0 0 0 -1 29230
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_144
timestamp 1626486988
transform 1 0 207 0 1 29193
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_143
timestamp 1626486988
transform 1 0 207 0 1 29430
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_142
timestamp 1626486988
transform 1 0 207 0 1 29193
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_93
timestamp 1626486988
transform 1 0 0 0 1 29230
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_141
timestamp 1626486988
transform 1 0 207 0 1 29746
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_92
timestamp 1626486988
transform 1 0 0 0 -1 30020
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_140
timestamp 1626486988
transform 1 0 207 0 1 29983
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_139
timestamp 1626486988
transform 1 0 207 0 1 30220
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_138
timestamp 1626486988
transform 1 0 207 0 1 29983
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_91
timestamp 1626486988
transform 1 0 0 0 1 30020
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_137
timestamp 1626486988
transform 1 0 207 0 1 30536
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_90
timestamp 1626486988
transform 1 0 0 0 -1 30810
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_136
timestamp 1626486988
transform 1 0 207 0 1 30773
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_135
timestamp 1626486988
transform 1 0 207 0 1 31010
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_134
timestamp 1626486988
transform 1 0 207 0 1 30773
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_89
timestamp 1626486988
transform 1 0 0 0 1 30810
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_133
timestamp 1626486988
transform 1 0 207 0 1 31326
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_132
timestamp 1626486988
transform 1 0 207 0 1 31563
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_130
timestamp 1626486988
transform 1 0 207 0 1 31563
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_87
timestamp 1626486988
transform 1 0 0 0 1 31600
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_88
timestamp 1626486988
transform 1 0 0 0 -1 31600
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_131
timestamp 1626486988
transform 1 0 207 0 1 31800
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_190
timestamp 1626486988
transform 1 0 207 0 1 32353
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_129
timestamp 1626486988
transform 1 0 207 0 1 32116
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_128
timestamp 1626486988
transform 1 0 207 0 1 32353
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_85
timestamp 1626486988
transform 1 0 0 0 1 32390
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_86
timestamp 1626486988
transform 1 0 0 0 -1 32390
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1626486988
transform 1 0 207 0 1 32590
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_84
timestamp 1626486988
transform 1 0 0 0 -1 33180
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_189
timestamp 1626486988
transform 1 0 207 0 1 32906
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_188
timestamp 1626486988
transform 1 0 207 0 1 33143
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_186
timestamp 1626486988
transform 1 0 207 0 1 33143
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_83
timestamp 1626486988
transform 1 0 0 0 1 33180
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_187
timestamp 1626486988
transform 1 0 207 0 1 33380
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_185
timestamp 1626486988
transform 1 0 207 0 1 33696
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_82
timestamp 1626486988
transform 1 0 0 0 -1 33970
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_184
timestamp 1626486988
transform 1 0 207 0 1 33933
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_182
timestamp 1626486988
transform 1 0 207 0 1 33933
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_81
timestamp 1626486988
transform 1 0 0 0 1 33970
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_183
timestamp 1626486988
transform 1 0 207 0 1 34170
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_181
timestamp 1626486988
transform 1 0 207 0 1 34486
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_80
timestamp 1626486988
transform 1 0 0 0 -1 34760
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_180
timestamp 1626486988
transform 1 0 207 0 1 34723
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_179
timestamp 1626486988
transform 1 0 207 0 1 34960
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_178
timestamp 1626486988
transform 1 0 207 0 1 34723
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_79
timestamp 1626486988
transform 1 0 0 0 1 34760
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_177
timestamp 1626486988
transform 1 0 207 0 1 35276
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_78
timestamp 1626486988
transform 1 0 0 0 -1 35550
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_176
timestamp 1626486988
transform 1 0 207 0 1 35513
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_175
timestamp 1626486988
transform 1 0 207 0 1 35750
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_174
timestamp 1626486988
transform 1 0 207 0 1 35513
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_77
timestamp 1626486988
transform 1 0 0 0 1 35550
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_173
timestamp 1626486988
transform 1 0 207 0 1 36066
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_75
timestamp 1626486988
transform 1 0 0 0 1 36340
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_76
timestamp 1626486988
transform 1 0 0 0 -1 36340
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_172
timestamp 1626486988
transform 1 0 207 0 1 36303
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_171
timestamp 1626486988
transform 1 0 207 0 1 36540
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_170
timestamp 1626486988
transform 1 0 207 0 1 36303
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_169
timestamp 1626486988
transform 1 0 207 0 1 36856
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_168
timestamp 1626486988
transform 1 0 207 0 1 37093
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_166
timestamp 1626486988
transform 1 0 207 0 1 37093
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_73
timestamp 1626486988
transform 1 0 0 0 1 37130
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_74
timestamp 1626486988
transform 1 0 0 0 -1 37130
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_167
timestamp 1626486988
transform 1 0 207 0 1 37330
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_72
timestamp 1626486988
transform 1 0 0 0 -1 37920
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_165
timestamp 1626486988
transform 1 0 207 0 1 37646
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_164
timestamp 1626486988
transform 1 0 207 0 1 37883
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_162
timestamp 1626486988
transform 1 0 207 0 1 37883
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_71
timestamp 1626486988
transform 1 0 0 0 1 37920
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_163
timestamp 1626486988
transform 1 0 207 0 1 38120
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_70
timestamp 1626486988
transform 1 0 0 0 -1 38710
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_161
timestamp 1626486988
transform 1 0 207 0 1 38436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_160
timestamp 1626486988
transform 1 0 207 0 1 38673
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_159
timestamp 1626486988
transform 1 0 207 0 1 38673
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_127
timestamp 1626486988
transform 1 0 0 0 1 38710
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_253
timestamp 1626486988
transform 1 0 207 0 1 38910
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_252
timestamp 1626486988
transform 1 0 207 0 1 39226
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_95
timestamp 1626486988
transform 1 0 0 0 -1 39500
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_251
timestamp 1626486988
transform 1 0 207 0 1 39463
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_250
timestamp 1626486988
transform 1 0 207 0 1 39700
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_249
timestamp 1626486988
transform 1 0 207 0 1 39463
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_126
timestamp 1626486988
transform 1 0 0 0 1 39500
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_248
timestamp 1626486988
transform 1 0 207 0 1 40016
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_125
timestamp 1626486988
transform 1 0 0 0 -1 40290
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_247
timestamp 1626486988
transform 1 0 207 0 1 40253
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_246
timestamp 1626486988
transform 1 0 207 0 1 40490
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_245
timestamp 1626486988
transform 1 0 207 0 1 40253
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_124
timestamp 1626486988
transform 1 0 0 0 1 40290
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_244
timestamp 1626486988
transform 1 0 207 0 1 40806
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_123
timestamp 1626486988
transform 1 0 0 0 -1 41080
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_243
timestamp 1626486988
transform 1 0 207 0 1 41043
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_242
timestamp 1626486988
transform 1 0 207 0 1 41280
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_241
timestamp 1626486988
transform 1 0 207 0 1 41043
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_122
timestamp 1626486988
transform 1 0 0 0 1 41080
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_240
timestamp 1626486988
transform 1 0 207 0 1 41596
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_239
timestamp 1626486988
transform 1 0 207 0 1 41833
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_237
timestamp 1626486988
transform 1 0 207 0 1 41833
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_120
timestamp 1626486988
transform 1 0 0 0 1 41870
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_121
timestamp 1626486988
transform 1 0 0 0 -1 41870
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_238
timestamp 1626486988
transform 1 0 207 0 1 42070
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_236
timestamp 1626486988
transform 1 0 207 0 1 42386
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_235
timestamp 1626486988
transform 1 0 207 0 1 42623
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_233
timestamp 1626486988
transform 1 0 207 0 1 42623
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_118
timestamp 1626486988
transform 1 0 0 0 1 42660
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_119
timestamp 1626486988
transform 1 0 0 0 -1 42660
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_234
timestamp 1626486988
transform 1 0 207 0 1 42860
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_117
timestamp 1626486988
transform 1 0 0 0 -1 43450
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_232
timestamp 1626486988
transform 1 0 207 0 1 43176
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_231
timestamp 1626486988
transform 1 0 207 0 1 43413
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_229
timestamp 1626486988
transform 1 0 207 0 1 43413
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_116
timestamp 1626486988
transform 1 0 0 0 1 43450
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_230
timestamp 1626486988
transform 1 0 207 0 1 43650
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_228
timestamp 1626486988
transform 1 0 207 0 1 43966
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_115
timestamp 1626486988
transform 1 0 0 0 -1 44240
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_227
timestamp 1626486988
transform 1 0 207 0 1 44203
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_225
timestamp 1626486988
transform 1 0 207 0 1 44203
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_114
timestamp 1626486988
transform 1 0 0 0 1 44240
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_226
timestamp 1626486988
transform 1 0 207 0 1 44440
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_224
timestamp 1626486988
transform 1 0 207 0 1 44756
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_113
timestamp 1626486988
transform 1 0 0 0 -1 45030
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_223
timestamp 1626486988
transform 1 0 207 0 1 44993
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_222
timestamp 1626486988
transform 1 0 207 0 1 45230
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_221
timestamp 1626486988
transform 1 0 207 0 1 44993
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_112
timestamp 1626486988
transform 1 0 0 0 1 45030
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_220
timestamp 1626486988
transform 1 0 207 0 1 45546
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_111
timestamp 1626486988
transform 1 0 0 0 -1 45820
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_219
timestamp 1626486988
transform 1 0 207 0 1 45783
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_218
timestamp 1626486988
transform 1 0 207 0 1 46020
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_217
timestamp 1626486988
transform 1 0 207 0 1 45783
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_110
timestamp 1626486988
transform 1 0 0 0 1 45820
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_216
timestamp 1626486988
transform 1 0 207 0 1 46336
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_109
timestamp 1626486988
transform 1 0 0 0 -1 46610
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_215
timestamp 1626486988
transform 1 0 207 0 1 46573
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_214
timestamp 1626486988
transform 1 0 207 0 1 46810
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_213
timestamp 1626486988
transform 1 0 207 0 1 46573
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_108
timestamp 1626486988
transform 1 0 0 0 1 46610
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_212
timestamp 1626486988
transform 1 0 207 0 1 47126
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_211
timestamp 1626486988
transform 1 0 207 0 1 47363
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_209
timestamp 1626486988
transform 1 0 207 0 1 47363
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_106
timestamp 1626486988
transform 1 0 0 0 1 47400
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_107
timestamp 1626486988
transform 1 0 0 0 -1 47400
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_210
timestamp 1626486988
transform 1 0 207 0 1 47600
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_208
timestamp 1626486988
transform 1 0 207 0 1 47916
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_207
timestamp 1626486988
transform 1 0 207 0 1 48153
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_205
timestamp 1626486988
transform 1 0 207 0 1 48153
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_104
timestamp 1626486988
transform 1 0 0 0 1 48190
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_105
timestamp 1626486988
transform 1 0 0 0 -1 48190
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_206
timestamp 1626486988
transform 1 0 207 0 1 48390
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_103
timestamp 1626486988
transform 1 0 0 0 -1 48980
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_204
timestamp 1626486988
transform 1 0 207 0 1 48706
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_203
timestamp 1626486988
transform 1 0 207 0 1 48943
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_201
timestamp 1626486988
transform 1 0 207 0 1 48943
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_102
timestamp 1626486988
transform 1 0 0 0 1 48980
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_202
timestamp 1626486988
transform 1 0 207 0 1 49180
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_200
timestamp 1626486988
transform 1 0 207 0 1 49496
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_101
timestamp 1626486988
transform 1 0 0 0 -1 49770
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_199
timestamp 1626486988
transform 1 0 207 0 1 49733
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_197
timestamp 1626486988
transform 1 0 207 0 1 49733
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_100
timestamp 1626486988
transform 1 0 0 0 1 49770
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_198
timestamp 1626486988
transform 1 0 207 0 1 49970
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_196
timestamp 1626486988
transform 1 0 207 0 1 50286
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_99
timestamp 1626486988
transform 1 0 0 0 -1 50560
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_195
timestamp 1626486988
transform 1 0 207 0 1 50523
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_194
timestamp 1626486988
transform 1 0 207 0 1 50760
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_193
timestamp 1626486988
transform 1 0 207 0 1 50523
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_98
timestamp 1626486988
transform 1 0 0 0 1 50560
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_192
timestamp 1626486988
transform 1 0 207 0 1 51076
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_97
timestamp 1626486988
transform 1 0 0 0 -1 51350
box -42 -55 624 371
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_191
timestamp 1626486988
transform 1 0 207 0 1 51313
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_96
timestamp 1626486988
transform 1 0 0 0 1 51350
box -42 -55 624 371
<< labels >>
rlabel metal3 s 191 35738 289 35836 4 gnd
rlabel metal3 s 191 39688 289 39786 4 gnd
rlabel metal3 s 191 34711 289 34809 4 gnd
rlabel metal3 s 191 28154 289 28252 4 gnd
rlabel metal3 s 191 35501 289 35599 4 gnd
rlabel metal3 s 191 42848 289 42946 4 gnd
rlabel metal3 s 191 47114 289 47212 4 gnd
rlabel metal3 s 191 46008 289 46106 4 gnd
rlabel metal3 s 191 28628 289 28726 4 gnd
rlabel metal3 s 191 42058 289 42156 4 gnd
rlabel metal3 s 191 44191 289 44289 4 gnd
rlabel metal3 s 191 32578 289 32676 4 gnd
rlabel metal3 s 191 38898 289 38996 4 gnd
rlabel metal3 s 191 44428 289 44526 4 gnd
rlabel metal3 s 191 30761 289 30859 4 gnd
rlabel metal3 s 191 51064 289 51162 4 gnd
rlabel metal3 s 191 30208 289 30306 4 gnd
rlabel metal3 s 191 38424 289 38522 4 gnd
rlabel metal3 s 191 50748 289 50846 4 gnd
rlabel metal3 s 191 39214 289 39312 4 gnd
rlabel metal3 s 191 31788 289 31886 4 gnd
rlabel metal3 s 191 36291 289 36389 4 gnd
rlabel metal3 s 191 40004 289 40102 4 gnd
rlabel metal3 s 191 49721 289 49819 4 gnd
rlabel metal3 s 191 34948 289 35046 4 gnd
rlabel metal3 s 191 48931 289 49029 4 gnd
rlabel metal3 s 191 40241 289 40339 4 gnd
rlabel metal3 s 191 29418 289 29516 4 gnd
rlabel metal3 s 191 31314 289 31412 4 gnd
rlabel metal3 s 191 47904 289 48002 4 gnd
rlabel metal3 s 191 38661 289 38759 4 gnd
rlabel metal3 s 191 28391 289 28489 4 gnd
rlabel metal3 s 191 33684 289 33782 4 gnd
rlabel metal3 s 191 41268 289 41366 4 gnd
rlabel metal3 s 191 30998 289 31096 4 gnd
rlabel metal3 s 191 46324 289 46422 4 gnd
rlabel metal3 s 191 49168 289 49266 4 gnd
rlabel metal3 s 191 49958 289 50056 4 gnd
rlabel metal3 s 191 37634 289 37732 4 gnd
rlabel metal3 s 191 49484 289 49582 4 gnd
rlabel metal3 s 191 38108 289 38206 4 gnd
rlabel metal3 s 191 47351 289 47449 4 gnd
rlabel metal3 s 191 29971 289 30069 4 gnd
rlabel metal3 s 191 40478 289 40576 4 gnd
rlabel metal3 s 191 33131 289 33229 4 gnd
rlabel metal3 s 191 47588 289 47686 4 gnd
rlabel metal3 s 191 48378 289 48476 4 gnd
rlabel metal3 s 191 26258 289 26356 4 gnd
rlabel metal3 s 191 31551 289 31649 4 gnd
rlabel metal3 s 191 41584 289 41682 4 gnd
rlabel metal3 s 191 48694 289 48792 4 gnd
rlabel metal3 s 191 29734 289 29832 4 gnd
rlabel metal3 s 191 43401 289 43499 4 gnd
rlabel metal3 s 191 32894 289 32992 4 gnd
rlabel metal3 s 191 36054 289 36152 4 gnd
rlabel metal3 s 191 33921 289 34019 4 gnd
rlabel metal3 s 191 26574 289 26672 4 gnd
rlabel metal3 s 191 50274 289 50372 4 gnd
rlabel metal3 s 191 30524 289 30622 4 gnd
rlabel metal3 s 191 33368 289 33466 4 gnd
rlabel metal3 s 191 36528 289 36626 4 gnd
rlabel metal3 s 191 46798 289 46896 4 gnd
rlabel metal3 s 191 37871 289 37969 4 gnd
rlabel metal3 s 191 45534 289 45632 4 gnd
rlabel metal3 s 191 42611 289 42709 4 gnd
rlabel metal3 s 191 42374 289 42472 4 gnd
rlabel metal3 s 191 43164 289 43262 4 gnd
rlabel metal3 s 191 35264 289 35362 4 gnd
rlabel metal3 s 191 32341 289 32439 4 gnd
rlabel metal3 s 191 43638 289 43736 4 gnd
rlabel metal3 s 191 45218 289 45316 4 gnd
rlabel metal3 s 191 36844 289 36942 4 gnd
rlabel metal3 s 191 46561 289 46659 4 gnd
rlabel metal3 s 191 27048 289 27146 4 gnd
rlabel metal3 s 191 26811 289 26909 4 gnd
rlabel metal3 s 191 40794 289 40892 4 gnd
rlabel metal3 s 191 41821 289 41919 4 gnd
rlabel metal3 s 191 37318 289 37416 4 gnd
rlabel metal3 s 191 51301 289 51399 4 gnd
rlabel metal3 s 191 29181 289 29279 4 gnd
rlabel metal3 s 191 39451 289 39549 4 gnd
rlabel metal3 s 191 43954 289 44052 4 gnd
rlabel metal3 s 191 45771 289 45869 4 gnd
rlabel metal3 s 191 41031 289 41129 4 gnd
rlabel metal3 s 191 28944 289 29042 4 gnd
rlabel metal3 s 191 34474 289 34572 4 gnd
rlabel metal3 s 191 27601 289 27699 4 gnd
rlabel metal3 s 191 37081 289 37179 4 gnd
rlabel metal3 s 191 34158 289 34256 4 gnd
rlabel metal3 s 191 44744 289 44842 4 gnd
rlabel metal3 s 191 48141 289 48239 4 gnd
rlabel metal3 s 191 44981 289 45079 4 gnd
rlabel metal3 s 191 27364 289 27462 4 gnd
rlabel metal3 s 191 50511 289 50609 4 gnd
rlabel metal3 s 191 32104 289 32202 4 gnd
rlabel metal3 s 191 27838 289 27936 4 gnd
rlabel metal3 s 191 16778 289 16876 4 gnd
rlabel metal3 s 191 8404 289 8502 4 gnd
rlabel metal3 s 191 2558 289 2656 4 gnd
rlabel metal3 s 191 8878 289 8976 4 gnd
rlabel metal3 s 191 25468 289 25566 4 gnd
rlabel metal3 s 191 13618 289 13716 4 gnd
rlabel metal3 s 191 5244 289 5342 4 gnd
rlabel metal3 s 191 19701 289 19799 4 gnd
rlabel metal3 s 191 2874 289 2972 4 gnd
rlabel metal3 s 191 12591 289 12689 4 gnd
rlabel metal3 s 191 19938 289 20036 4 gnd
rlabel metal3 s 191 14171 289 14269 4 gnd
rlabel metal3 s 191 24441 289 24539 4 gnd
rlabel metal3 s 191 6824 289 6922 4 gnd
rlabel metal3 s 191 6034 289 6132 4 gnd
rlabel metal3 s 191 8641 289 8739 4 gnd
rlabel metal3 s 191 2084 289 2182 4 gnd
rlabel metal3 s 191 11248 289 11346 4 gnd
rlabel metal3 s 191 3664 289 3762 4 gnd
rlabel metal3 s 191 18674 289 18772 4 gnd
rlabel metal3 s 191 7851 289 7949 4 gnd
rlabel metal3 s 191 10774 289 10872 4 gnd
rlabel metal3 s 191 11801 289 11899 4 gnd
rlabel metal3 s 191 9431 289 9529 4 gnd
rlabel metal3 s 191 3901 289 3999 4 gnd
rlabel metal3 s 191 7614 289 7712 4 gnd
rlabel metal3 s 191 13381 289 13479 4 gnd
rlabel metal3 s 191 17568 289 17666 4 gnd
rlabel metal3 s 191 15751 289 15849 4 gnd
rlabel metal3 s 191 1768 289 1866 4 gnd
rlabel metal3 s 191 3348 289 3446 4 gnd
rlabel metal3 s 191 22861 289 22959 4 gnd
rlabel metal3 s 191 15514 289 15612 4 gnd
rlabel metal3 s 191 10458 289 10556 4 gnd
rlabel metal3 s 191 1531 289 1629 4 gnd
rlabel metal3 s 191 21281 289 21379 4 gnd
rlabel metal3 s 191 14724 289 14822 4 gnd
rlabel metal3 s 191 9668 289 9766 4 gnd
rlabel metal3 s 191 4138 289 4236 4 gnd
rlabel metal3 s 191 11564 289 11662 4 gnd
rlabel metal3 s 191 24678 289 24776 4 gnd
rlabel metal3 s 191 978 289 1076 4 gnd
rlabel metal3 s 191 17884 289 17982 4 gnd
rlabel metal3 s 191 13144 289 13242 4 gnd
rlabel metal3 s 191 23098 289 23196 4 gnd
rlabel metal3 s 191 6271 289 6369 4 gnd
rlabel metal3 s 191 11011 289 11109 4 gnd
rlabel metal3 s 191 18121 289 18219 4 gnd
rlabel metal3 s 191 12354 289 12452 4 gnd
rlabel metal3 s 191 1294 289 1392 4 gnd
rlabel metal3 s 191 741 289 839 4 gnd
rlabel metal3 s 191 25784 289 25882 4 gnd
rlabel metal3 s 191 21518 289 21616 4 gnd
rlabel metal3 s 191 21834 289 21932 4 gnd
rlabel metal3 s 191 26021 289 26119 4 gnd
rlabel metal3 s 191 14408 289 14506 4 gnd
rlabel metal3 s 191 7061 289 7159 4 gnd
rlabel metal3 s 191 8088 289 8186 4 gnd
rlabel metal3 s 191 12038 289 12136 4 gnd
rlabel metal3 s 191 4691 289 4789 4 gnd
rlabel metal3 s 191 20491 289 20589 4 gnd
rlabel metal3 s 191 6508 289 6606 4 gnd
rlabel metal3 s 191 16541 289 16639 4 gnd
rlabel metal3 s 191 17331 289 17429 4 gnd
rlabel metal3 s 191 22624 289 22722 4 gnd
rlabel metal3 s 191 24994 289 25092 4 gnd
rlabel metal3 s 191 23414 289 23512 4 gnd
rlabel metal3 s 191 13934 289 14032 4 gnd
rlabel metal3 s 191 16304 289 16402 4 gnd
rlabel metal3 s 191 4928 289 5026 4 gnd
rlabel metal3 s 191 15988 289 16086 4 gnd
rlabel metal3 s 191 18911 289 19009 4 gnd
rlabel metal3 s 191 14961 289 15059 4 gnd
rlabel metal3 s 191 22071 289 22169 4 gnd
rlabel metal3 s 191 25231 289 25329 4 gnd
rlabel metal3 s 191 17094 289 17192 4 gnd
rlabel metal3 s 191 20254 289 20352 4 gnd
rlabel metal3 s 191 21044 289 21142 4 gnd
rlabel metal3 s 191 23651 289 23749 4 gnd
rlabel metal3 s 191 3111 289 3209 4 gnd
rlabel metal3 s 191 15198 289 15296 4 gnd
rlabel metal3 s 191 19148 289 19246 4 gnd
rlabel metal3 s 191 7298 289 7396 4 gnd
rlabel metal3 s 191 5718 289 5816 4 gnd
rlabel metal3 s 191 4454 289 4552 4 gnd
rlabel metal3 s 191 19464 289 19562 4 gnd
rlabel metal3 s 191 22308 289 22406 4 gnd
rlabel metal3 s 191 9984 289 10082 4 gnd
rlabel metal3 s 191 20728 289 20826 4 gnd
rlabel metal3 s 191 10221 289 10319 4 gnd
rlabel metal3 s 191 9194 289 9292 4 gnd
rlabel metal3 s 191 5481 289 5579 4 gnd
rlabel metal3 s 191 24204 289 24302 4 gnd
rlabel metal3 s 191 18358 289 18456 4 gnd
rlabel metal3 s 191 12828 289 12926 4 gnd
rlabel metal3 s 191 2321 289 2419 4 gnd
rlabel metal3 s 191 23888 289 23986 4 gnd
rlabel metal2 s 0 39033 28 39081 4 wl0_97
rlabel metal2 s 0 38813 28 38861 4 wl1_97
rlabel metal2 s 0 39129 28 39177 4 wl0_98
rlabel metal2 s 0 39349 28 39397 4 wl1_98
rlabel metal2 s 0 39823 28 39871 4 wl0_99
rlabel metal2 s 0 39603 28 39651 4 wl1_99
rlabel metal2 s 0 39919 28 39967 4 wl0_100
rlabel metal2 s 0 40139 28 40187 4 wl1_100
rlabel metal2 s 0 40613 28 40661 4 wl0_101
rlabel metal2 s 0 40393 28 40441 4 wl1_101
rlabel metal2 s 0 40709 28 40757 4 wl0_102
rlabel metal2 s 0 40929 28 40977 4 wl1_102
rlabel metal2 s 0 41403 28 41451 4 wl0_103
rlabel metal2 s 0 41183 28 41231 4 wl1_103
rlabel metal2 s 0 41499 28 41547 4 wl0_104
rlabel metal2 s 0 41719 28 41767 4 wl1_104
rlabel metal2 s 0 42193 28 42241 4 wl0_105
rlabel metal2 s 0 41973 28 42021 4 wl1_105
rlabel metal2 s 0 42289 28 42337 4 wl0_106
rlabel metal2 s 0 42509 28 42557 4 wl1_106
rlabel metal2 s 0 42983 28 43031 4 wl0_107
rlabel metal2 s 0 42763 28 42811 4 wl1_107
rlabel metal2 s 0 43079 28 43127 4 wl0_108
rlabel metal2 s 0 43299 28 43347 4 wl1_108
rlabel metal2 s 0 43773 28 43821 4 wl0_109
rlabel metal2 s 0 43553 28 43601 4 wl1_109
rlabel metal2 s 0 43869 28 43917 4 wl0_110
rlabel metal2 s 0 44089 28 44137 4 wl1_110
rlabel metal2 s 0 44563 28 44611 4 wl0_111
rlabel metal2 s 0 44343 28 44391 4 wl1_111
rlabel metal2 s 0 44659 28 44707 4 wl0_112
rlabel metal2 s 0 44879 28 44927 4 wl1_112
rlabel metal2 s 0 45353 28 45401 4 wl0_113
rlabel metal2 s 0 45133 28 45181 4 wl1_113
rlabel metal2 s 0 45449 28 45497 4 wl0_114
rlabel metal2 s 0 45669 28 45717 4 wl1_114
rlabel metal2 s 0 46143 28 46191 4 wl0_115
rlabel metal2 s 0 45923 28 45971 4 wl1_115
rlabel metal2 s 0 46239 28 46287 4 wl0_116
rlabel metal2 s 0 46459 28 46507 4 wl1_116
rlabel metal2 s 0 46933 28 46981 4 wl0_117
rlabel metal2 s 0 46713 28 46761 4 wl1_117
rlabel metal2 s 0 47029 28 47077 4 wl0_118
rlabel metal2 s 0 47249 28 47297 4 wl1_118
rlabel metal2 s 0 47723 28 47771 4 wl0_119
rlabel metal2 s 0 47503 28 47551 4 wl1_119
rlabel metal2 s 0 47819 28 47867 4 wl0_120
rlabel metal2 s 0 48039 28 48087 4 wl1_120
rlabel metal2 s 0 48513 28 48561 4 wl0_121
rlabel metal2 s 0 48293 28 48341 4 wl1_121
rlabel metal2 s 0 48609 28 48657 4 wl0_122
rlabel metal2 s 0 48829 28 48877 4 wl1_122
rlabel metal2 s 0 49303 28 49351 4 wl0_123
rlabel metal2 s 0 49083 28 49131 4 wl1_123
rlabel metal2 s 0 49399 28 49447 4 wl0_124
rlabel metal2 s 0 49619 28 49667 4 wl1_124
rlabel metal2 s 0 50093 28 50141 4 wl0_125
rlabel metal2 s 0 49873 28 49921 4 wl1_125
rlabel metal2 s 0 50189 28 50237 4 wl0_126
rlabel metal2 s 0 50409 28 50457 4 wl1_126
rlabel metal2 s 0 50883 28 50931 4 wl0_127
rlabel metal2 s 0 50663 28 50711 4 wl1_127
rlabel metal2 s 0 50979 28 51027 4 wl0_128
rlabel metal2 s 0 51199 28 51247 4 wl1_128
rlabel metal2 s 0 26393 28 26441 4 wl0_65
rlabel metal2 s 0 26173 28 26221 4 wl1_65
rlabel metal2 s 0 26489 28 26537 4 wl0_66
rlabel metal2 s 0 26709 28 26757 4 wl1_66
rlabel metal2 s 0 27183 28 27231 4 wl0_67
rlabel metal2 s 0 26963 28 27011 4 wl1_67
rlabel metal2 s 0 27279 28 27327 4 wl0_68
rlabel metal2 s 0 27499 28 27547 4 wl1_68
rlabel metal2 s 0 27973 28 28021 4 wl0_69
rlabel metal2 s 0 27753 28 27801 4 wl1_69
rlabel metal2 s 0 28069 28 28117 4 wl0_70
rlabel metal2 s 0 28289 28 28337 4 wl1_70
rlabel metal2 s 0 28763 28 28811 4 wl0_71
rlabel metal2 s 0 28543 28 28591 4 wl1_71
rlabel metal2 s 0 28859 28 28907 4 wl0_72
rlabel metal2 s 0 29079 28 29127 4 wl1_72
rlabel metal2 s 0 29553 28 29601 4 wl0_73
rlabel metal2 s 0 29333 28 29381 4 wl1_73
rlabel metal2 s 0 29649 28 29697 4 wl0_74
rlabel metal2 s 0 29869 28 29917 4 wl1_74
rlabel metal2 s 0 30343 28 30391 4 wl0_75
rlabel metal2 s 0 30123 28 30171 4 wl1_75
rlabel metal2 s 0 30439 28 30487 4 wl0_76
rlabel metal2 s 0 30659 28 30707 4 wl1_76
rlabel metal2 s 0 31133 28 31181 4 wl0_77
rlabel metal2 s 0 30913 28 30961 4 wl1_77
rlabel metal2 s 0 31229 28 31277 4 wl0_78
rlabel metal2 s 0 31449 28 31497 4 wl1_78
rlabel metal2 s 0 31923 28 31971 4 wl0_79
rlabel metal2 s 0 31703 28 31751 4 wl1_79
rlabel metal2 s 0 32019 28 32067 4 wl0_80
rlabel metal2 s 0 32239 28 32287 4 wl1_80
rlabel metal2 s 0 32713 28 32761 4 wl0_81
rlabel metal2 s 0 32493 28 32541 4 wl1_81
rlabel metal2 s 0 32809 28 32857 4 wl0_82
rlabel metal2 s 0 33029 28 33077 4 wl1_82
rlabel metal2 s 0 33503 28 33551 4 wl0_83
rlabel metal2 s 0 33283 28 33331 4 wl1_83
rlabel metal2 s 0 33599 28 33647 4 wl0_84
rlabel metal2 s 0 33819 28 33867 4 wl1_84
rlabel metal2 s 0 34293 28 34341 4 wl0_85
rlabel metal2 s 0 34073 28 34121 4 wl1_85
rlabel metal2 s 0 34389 28 34437 4 wl0_86
rlabel metal2 s 0 34609 28 34657 4 wl1_86
rlabel metal2 s 0 35083 28 35131 4 wl0_87
rlabel metal2 s 0 34863 28 34911 4 wl1_87
rlabel metal2 s 0 35179 28 35227 4 wl0_88
rlabel metal2 s 0 35399 28 35447 4 wl1_88
rlabel metal2 s 0 35873 28 35921 4 wl0_89
rlabel metal2 s 0 35653 28 35701 4 wl1_89
rlabel metal2 s 0 35969 28 36017 4 wl0_90
rlabel metal2 s 0 36189 28 36237 4 wl1_90
rlabel metal2 s 0 36663 28 36711 4 wl0_91
rlabel metal2 s 0 36443 28 36491 4 wl1_91
rlabel metal2 s 0 36759 28 36807 4 wl0_92
rlabel metal2 s 0 36979 28 37027 4 wl1_92
rlabel metal2 s 0 37453 28 37501 4 wl0_93
rlabel metal2 s 0 37233 28 37281 4 wl1_93
rlabel metal2 s 0 37549 28 37597 4 wl0_94
rlabel metal2 s 0 37769 28 37817 4 wl1_94
rlabel metal2 s 0 38243 28 38291 4 wl0_95
rlabel metal2 s 0 38023 28 38071 4 wl1_95
rlabel metal2 s 0 38339 28 38387 4 wl0_96
rlabel metal2 s 0 38559 28 38607 4 wl1_96
rlabel metal2 s 0 13753 28 13801 4 wl0_33
rlabel metal2 s 0 13533 28 13581 4 wl1_33
rlabel metal2 s 0 13849 28 13897 4 wl0_34
rlabel metal2 s 0 14069 28 14117 4 wl1_34
rlabel metal2 s 0 14543 28 14591 4 wl0_35
rlabel metal2 s 0 14323 28 14371 4 wl1_35
rlabel metal2 s 0 14639 28 14687 4 wl0_36
rlabel metal2 s 0 14859 28 14907 4 wl1_36
rlabel metal2 s 0 15333 28 15381 4 wl0_37
rlabel metal2 s 0 15113 28 15161 4 wl1_37
rlabel metal2 s 0 15429 28 15477 4 wl0_38
rlabel metal2 s 0 15649 28 15697 4 wl1_38
rlabel metal2 s 0 16123 28 16171 4 wl0_39
rlabel metal2 s 0 15903 28 15951 4 wl1_39
rlabel metal2 s 0 16219 28 16267 4 wl0_40
rlabel metal2 s 0 16439 28 16487 4 wl1_40
rlabel metal2 s 0 16913 28 16961 4 wl0_41
rlabel metal2 s 0 16693 28 16741 4 wl1_41
rlabel metal2 s 0 17009 28 17057 4 wl0_42
rlabel metal2 s 0 17229 28 17277 4 wl1_42
rlabel metal2 s 0 17703 28 17751 4 wl0_43
rlabel metal2 s 0 17483 28 17531 4 wl1_43
rlabel metal2 s 0 17799 28 17847 4 wl0_44
rlabel metal2 s 0 18019 28 18067 4 wl1_44
rlabel metal2 s 0 18493 28 18541 4 wl0_45
rlabel metal2 s 0 18273 28 18321 4 wl1_45
rlabel metal2 s 0 18589 28 18637 4 wl0_46
rlabel metal2 s 0 18809 28 18857 4 wl1_46
rlabel metal2 s 0 19283 28 19331 4 wl0_47
rlabel metal2 s 0 19063 28 19111 4 wl1_47
rlabel metal2 s 0 19379 28 19427 4 wl0_48
rlabel metal2 s 0 19599 28 19647 4 wl1_48
rlabel metal2 s 0 20073 28 20121 4 wl0_49
rlabel metal2 s 0 19853 28 19901 4 wl1_49
rlabel metal2 s 0 20169 28 20217 4 wl0_50
rlabel metal2 s 0 20389 28 20437 4 wl1_50
rlabel metal2 s 0 20863 28 20911 4 wl0_51
rlabel metal2 s 0 20643 28 20691 4 wl1_51
rlabel metal2 s 0 20959 28 21007 4 wl0_52
rlabel metal2 s 0 21179 28 21227 4 wl1_52
rlabel metal2 s 0 21653 28 21701 4 wl0_53
rlabel metal2 s 0 21433 28 21481 4 wl1_53
rlabel metal2 s 0 21749 28 21797 4 wl0_54
rlabel metal2 s 0 21969 28 22017 4 wl1_54
rlabel metal2 s 0 22443 28 22491 4 wl0_55
rlabel metal2 s 0 22223 28 22271 4 wl1_55
rlabel metal2 s 0 22539 28 22587 4 wl0_56
rlabel metal2 s 0 22759 28 22807 4 wl1_56
rlabel metal2 s 0 23233 28 23281 4 wl0_57
rlabel metal2 s 0 23013 28 23061 4 wl1_57
rlabel metal2 s 0 23329 28 23377 4 wl0_58
rlabel metal2 s 0 23549 28 23597 4 wl1_58
rlabel metal2 s 0 24023 28 24071 4 wl0_59
rlabel metal2 s 0 23803 28 23851 4 wl1_59
rlabel metal2 s 0 24119 28 24167 4 wl0_60
rlabel metal2 s 0 24339 28 24387 4 wl1_60
rlabel metal2 s 0 24813 28 24861 4 wl0_61
rlabel metal2 s 0 24593 28 24641 4 wl1_61
rlabel metal2 s 0 24909 28 24957 4 wl0_62
rlabel metal2 s 0 25129 28 25177 4 wl1_62
rlabel metal2 s 0 25603 28 25651 4 wl0_63
rlabel metal2 s 0 25383 28 25431 4 wl1_63
rlabel metal2 s 0 25699 28 25747 4 wl0_64
rlabel metal2 s 0 25919 28 25967 4 wl1_64
rlabel metal2 s 0 1113 28 1161 4 wl0_1
rlabel metal2 s 0 893 28 941 4 wl1_1
rlabel metal2 s 0 1209 28 1257 4 wl0_2
rlabel metal2 s 0 1429 28 1477 4 wl1_2
rlabel metal2 s 0 1903 28 1951 4 wl0_3
rlabel metal2 s 0 1683 28 1731 4 wl1_3
rlabel metal2 s 0 1999 28 2047 4 wl0_4
rlabel metal2 s 0 2219 28 2267 4 wl1_4
rlabel metal2 s 0 2693 28 2741 4 wl0_5
rlabel metal2 s 0 2473 28 2521 4 wl1_5
rlabel metal2 s 0 2789 28 2837 4 wl0_6
rlabel metal2 s 0 3009 28 3057 4 wl1_6
rlabel metal2 s 0 3483 28 3531 4 wl0_7
rlabel metal2 s 0 3263 28 3311 4 wl1_7
rlabel metal2 s 0 3579 28 3627 4 wl0_8
rlabel metal2 s 0 3799 28 3847 4 wl1_8
rlabel metal2 s 0 4273 28 4321 4 wl0_9
rlabel metal2 s 0 4053 28 4101 4 wl1_9
rlabel metal2 s 0 4369 28 4417 4 wl0_10
rlabel metal2 s 0 4589 28 4637 4 wl1_10
rlabel metal2 s 0 5063 28 5111 4 wl0_11
rlabel metal2 s 0 4843 28 4891 4 wl1_11
rlabel metal2 s 0 5159 28 5207 4 wl0_12
rlabel metal2 s 0 5379 28 5427 4 wl1_12
rlabel metal2 s 0 5853 28 5901 4 wl0_13
rlabel metal2 s 0 5633 28 5681 4 wl1_13
rlabel metal2 s 0 5949 28 5997 4 wl0_14
rlabel metal2 s 0 6169 28 6217 4 wl1_14
rlabel metal2 s 0 6643 28 6691 4 wl0_15
rlabel metal2 s 0 6423 28 6471 4 wl1_15
rlabel metal2 s 0 6739 28 6787 4 wl0_16
rlabel metal2 s 0 6959 28 7007 4 wl1_16
rlabel metal2 s 0 7433 28 7481 4 wl0_17
rlabel metal2 s 0 7213 28 7261 4 wl1_17
rlabel metal2 s 0 7529 28 7577 4 wl0_18
rlabel metal2 s 0 7749 28 7797 4 wl1_18
rlabel metal2 s 0 8223 28 8271 4 wl0_19
rlabel metal2 s 0 8003 28 8051 4 wl1_19
rlabel metal2 s 0 8319 28 8367 4 wl0_20
rlabel metal2 s 0 8539 28 8587 4 wl1_20
rlabel metal2 s 0 9013 28 9061 4 wl0_21
rlabel metal2 s 0 8793 28 8841 4 wl1_21
rlabel metal2 s 0 9109 28 9157 4 wl0_22
rlabel metal2 s 0 9329 28 9377 4 wl1_22
rlabel metal2 s 0 9803 28 9851 4 wl0_23
rlabel metal2 s 0 9583 28 9631 4 wl1_23
rlabel metal2 s 0 9899 28 9947 4 wl0_24
rlabel metal2 s 0 10119 28 10167 4 wl1_24
rlabel metal2 s 0 10593 28 10641 4 wl0_25
rlabel metal2 s 0 10373 28 10421 4 wl1_25
rlabel metal2 s 0 10689 28 10737 4 wl0_26
rlabel metal2 s 0 10909 28 10957 4 wl1_26
rlabel metal2 s 0 11383 28 11431 4 wl0_27
rlabel metal2 s 0 11163 28 11211 4 wl1_27
rlabel metal2 s 0 11479 28 11527 4 wl0_28
rlabel metal2 s 0 11699 28 11747 4 wl1_28
rlabel metal2 s 0 12173 28 12221 4 wl0_29
rlabel metal2 s 0 11953 28 12001 4 wl1_29
rlabel metal2 s 0 12269 28 12317 4 wl0_30
rlabel metal2 s 0 12489 28 12537 4 wl1_30
rlabel metal2 s 0 12963 28 13011 4 wl0_31
rlabel metal2 s 0 12743 28 12791 4 wl1_31
rlabel metal2 s 0 13059 28 13107 4 wl0_32
rlabel metal2 s 0 13279 28 13327 4 wl1_32
<< properties >>
string FIXED_BBOX 0 0 624 51745
<< end >>
