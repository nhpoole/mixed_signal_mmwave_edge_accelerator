magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal1 >>
rect 3283 -5276 5663 -5248
rect 2115 -5378 5539 -5350
<< metal2 >>
rect 2101 -6379 2129 -5364
rect 3269 -6379 3297 -5262
rect 5525 -5364 5553 2850
rect 5649 -5262 5677 4340
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 3251 0 1 -5294
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 5631 0 1 4308
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 5631 0 1 -5294
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 2083 0 1 -5396
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 5507 0 1 2818
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 5507 0 1 -5396
box 0 0 64 64
<< properties >>
string FIXED_BBOX 2083 -6379 5695 4372
<< end >>
