magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal2 >>
rect 14312 1401 14368 1449
rect 16808 1401 16864 1449
rect 19304 1401 19360 1449
rect 21800 1401 21856 1449
rect 24296 1401 24352 1449
rect 26792 1401 26848 1449
rect 29288 1401 29344 1449
rect 31784 1401 31840 1449
rect 34280 1401 34336 1449
rect 36776 1401 36832 1449
rect 39272 1401 39328 1449
rect 41768 1401 41824 1449
rect 44264 1401 44320 1449
rect 46760 1401 46816 1449
rect 49256 1401 49312 1449
rect 51752 1401 51808 1449
rect 54248 1401 54304 1449
rect 56744 1401 56800 1449
rect 59240 1401 59296 1449
rect 61736 1401 61792 1449
rect 64232 1401 64288 1449
rect 66728 1401 66784 1449
rect 69224 1401 69280 1449
rect 71720 1401 71776 1449
rect 74216 1401 74272 1449
rect 76712 1401 76768 1449
rect 79208 1401 79264 1449
rect 81704 1401 81760 1449
rect 84200 1401 84256 1449
rect 86696 1401 86752 1449
rect 89192 1401 89248 1449
rect 91688 1401 91744 1449
<< metal3 >>
rect 14265 1393 14415 1457
rect 16761 1393 16911 1457
rect 19257 1393 19407 1457
rect 21753 1393 21903 1457
rect 24249 1393 24399 1457
rect 26745 1393 26895 1457
rect 29241 1393 29391 1457
rect 31737 1393 31887 1457
rect 34233 1393 34383 1457
rect 36729 1393 36879 1457
rect 39225 1393 39375 1457
rect 41721 1393 41871 1457
rect 44217 1393 44367 1457
rect 46713 1393 46863 1457
rect 49209 1393 49359 1457
rect 51705 1393 51855 1457
rect 54201 1393 54351 1457
rect 56697 1393 56847 1457
rect 59193 1393 59343 1457
rect 61689 1393 61839 1457
rect 64185 1393 64335 1457
rect 66681 1393 66831 1457
rect 69177 1393 69327 1457
rect 71673 1393 71823 1457
rect 74169 1393 74319 1457
rect 76665 1393 76815 1457
rect 79161 1393 79311 1457
rect 81657 1393 81807 1457
rect 84153 1393 84303 1457
rect 86649 1393 86799 1457
rect 89145 1393 89295 1457
rect 91641 1393 91791 1457
rect 13980 273 14130 337
rect 33948 273 34098 337
rect 53916 273 54066 337
rect 73884 273 74034 337
rect 23139 -514 44292 -454
rect 45331 -514 91716 -454
rect 12627 -758 21828 -698
rect 44163 -758 89220 -698
rect 21971 -1002 41796 -942
rect 42995 -1002 86724 -942
rect 41827 -1246 84228 -1186
rect 20803 -1490 39300 -1430
rect 40659 -1490 81732 -1430
rect 39491 -1734 79236 -1674
rect 38323 -1978 76740 -1918
rect 33651 -2222 66756 -2162
rect 31315 -2466 61764 -2406
rect 28979 -2710 56772 -2650
rect 14963 -2954 26820 -2894
rect 27811 -2954 54276 -2894
rect 26643 -3198 51780 -3138
rect 19635 -3442 36804 -3382
rect 37155 -3442 74244 -3382
rect 13795 -3686 24324 -3626
rect 25475 -3686 49284 -3626
rect 11459 -3930 19332 -3870
rect 24307 -3930 46788 -3870
rect 10291 -4174 16836 -4114
rect 18467 -4174 34308 -4114
rect 35987 -4174 71748 -4114
rect 9123 -4418 14340 -4358
rect 17299 -4418 31812 -4358
rect 32483 -4418 64260 -4358
rect 7955 -4662 73959 -4602
rect 6787 -4906 53991 -4846
rect 5619 -5150 34023 -5090
rect 34819 -5150 69252 -5090
rect 4451 -5394 14055 -5334
rect 16131 -5394 29316 -5334
rect 30147 -5394 59268 -5334
rect 4376 -6397 4526 -6333
rect 5544 -6397 5694 -6333
rect 6712 -6397 6862 -6333
rect 7880 -6397 8030 -6333
rect 9048 -6397 9198 -6333
rect 10216 -6397 10366 -6333
rect 11384 -6397 11534 -6333
rect 12552 -6397 12702 -6333
rect 13720 -6397 13870 -6333
rect 14888 -6397 15038 -6333
rect 16056 -6397 16206 -6333
rect 17224 -6397 17374 -6333
rect 18392 -6397 18542 -6333
rect 19560 -6397 19710 -6333
rect 20728 -6397 20878 -6333
rect 21896 -6397 22046 -6333
rect 23064 -6397 23214 -6333
rect 24232 -6397 24382 -6333
rect 25400 -6397 25550 -6333
rect 26568 -6397 26718 -6333
rect 27736 -6397 27886 -6333
rect 28904 -6397 29054 -6333
rect 30072 -6397 30222 -6333
rect 31240 -6397 31390 -6333
rect 32408 -6397 32558 -6333
rect 33576 -6397 33726 -6333
rect 34744 -6397 34894 -6333
rect 35912 -6397 36062 -6333
rect 37080 -6397 37230 -6333
rect 38248 -6397 38398 -6333
rect 39416 -6397 39566 -6333
rect 40584 -6397 40734 -6333
rect 41752 -6397 41902 -6333
rect 42920 -6397 43070 -6333
rect 44088 -6397 44238 -6333
rect 45256 -6397 45406 -6333
<< metal4 >>
rect 4421 -6365 4481 -5364
rect 5589 -6365 5649 -5120
rect 6757 -6365 6817 -4876
rect 7925 -6365 7985 -4632
rect 9093 -6365 9153 -4388
rect 10261 -6365 10321 -4144
rect 11429 -6365 11489 -3900
rect 12597 -6365 12657 -728
rect 13765 -6365 13825 -3656
rect 14025 -5364 14085 305
rect 14310 -4388 14370 1425
rect 14933 -6365 14993 -2924
rect 16806 -4144 16866 1425
rect 19302 -3900 19362 1425
rect 21798 -728 21858 1425
rect 16101 -6365 16161 -5364
rect 17269 -6365 17329 -4388
rect 18437 -6365 18497 -4144
rect 19605 -6365 19665 -3412
rect 20773 -6365 20833 -1460
rect 21941 -6365 22001 -972
rect 23109 -6365 23169 -484
rect 24294 -3656 24354 1425
rect 26790 -2924 26850 1425
rect 24277 -6365 24337 -3900
rect 25445 -6365 25505 -3656
rect 26613 -6365 26673 -3168
rect 27781 -6365 27841 -2924
rect 28949 -6365 29009 -2680
rect 29286 -5364 29346 1425
rect 30117 -6365 30177 -5364
rect 31285 -6365 31345 -2436
rect 31782 -4388 31842 1425
rect 32453 -6365 32513 -4388
rect 33621 -6365 33681 -2192
rect 33993 -5120 34053 305
rect 34278 -4144 34338 1425
rect 36774 -3412 36834 1425
rect 39270 -1460 39330 1425
rect 41766 -972 41826 1425
rect 44262 -484 44322 1425
rect 34789 -6365 34849 -5120
rect 35957 -6365 36017 -4144
rect 37125 -6365 37185 -3412
rect 38293 -6365 38353 -1948
rect 39461 -6365 39521 -1704
rect 40629 -6365 40689 -1460
rect 41797 -6365 41857 -1216
rect 42965 -6365 43025 -972
rect 44133 -6365 44193 -728
rect 45301 -6365 45361 -484
rect 46758 -3900 46818 1425
rect 49254 -3656 49314 1425
rect 51750 -3168 51810 1425
rect 53961 -4876 54021 305
rect 54246 -2924 54306 1425
rect 56742 -2680 56802 1425
rect 59238 -5364 59298 1425
rect 61734 -2436 61794 1425
rect 64230 -4388 64290 1425
rect 66726 -2192 66786 1425
rect 69222 -5120 69282 1425
rect 71718 -4144 71778 1425
rect 73929 -4632 73989 305
rect 74214 -3412 74274 1425
rect 76710 -1948 76770 1425
rect 79206 -1704 79266 1425
rect 81702 -1460 81762 1425
rect 84198 -1216 84258 1425
rect 86694 -972 86754 1425
rect 89190 -728 89250 1425
rect 91686 -484 91746 1425
use contact_32  contact_32_141
timestamp 1624494425
transform 1 0 4413 0 1 -5397
box 0 0 76 66
use contact_9  contact_9_70
timestamp 1624494425
transform 1 0 4418 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_140
timestamp 1624494425
transform 1 0 4413 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_129
timestamp 1624494425
transform 1 0 5581 0 1 -5153
box 0 0 76 66
use contact_9  contact_9_64
timestamp 1624494425
transform 1 0 5586 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_128
timestamp 1624494425
transform 1 0 5581 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_121
timestamp 1624494425
transform 1 0 6749 0 1 -4909
box 0 0 76 66
use contact_9  contact_9_60
timestamp 1624494425
transform 1 0 6754 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_120
timestamp 1624494425
transform 1 0 6749 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_58
timestamp 1624494425
transform 1 0 7922 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_116
timestamp 1624494425
transform 1 0 7917 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_56
timestamp 1624494425
transform 1 0 9090 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_112
timestamp 1624494425
transform 1 0 9085 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_50
timestamp 1624494425
transform 1 0 10258 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_100
timestamp 1624494425
transform 1 0 10253 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_44
timestamp 1624494425
transform 1 0 11426 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_88
timestamp 1624494425
transform 1 0 11421 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 12594 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_12
timestamp 1624494425
transform 1 0 12589 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_143
timestamp 1624494425
transform 1 0 14017 0 1 -5397
box 0 0 76 66
use contact_9  contact_9_40
timestamp 1624494425
transform 1 0 13762 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_80
timestamp 1624494425
transform 1 0 13757 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_30
timestamp 1624494425
transform 1 0 14930 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_60
timestamp 1624494425
transform 1 0 14925 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_137
timestamp 1624494425
transform 1 0 16093 0 1 -5397
box 0 0 76 66
use contact_9  contact_9_68
timestamp 1624494425
transform 1 0 16098 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_136
timestamp 1624494425
transform 1 0 16093 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_54
timestamp 1624494425
transform 1 0 17266 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_108
timestamp 1624494425
transform 1 0 17261 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_48
timestamp 1624494425
transform 1 0 18434 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_96
timestamp 1624494425
transform 1 0 18429 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_36
timestamp 1624494425
transform 1 0 19602 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_72
timestamp 1624494425
transform 1 0 19597 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 20770 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_32
timestamp 1624494425
transform 1 0 20765 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 21938 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_20
timestamp 1624494425
transform 1 0 21933 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_42
timestamp 1624494425
transform 1 0 24274 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_84
timestamp 1624494425
transform 1 0 24269 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 23106 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_4
timestamp 1624494425
transform 1 0 23101 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_38
timestamp 1624494425
transform 1 0 25442 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_76
timestamp 1624494425
transform 1 0 25437 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_32
timestamp 1624494425
transform 1 0 26610 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_64
timestamp 1624494425
transform 1 0 26605 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_139
timestamp 1624494425
transform 1 0 29278 0 1 -5397
box 0 0 76 66
use contact_9  contact_9_28
timestamp 1624494425
transform 1 0 27778 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_56
timestamp 1624494425
transform 1 0 27773 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_26
timestamp 1624494425
transform 1 0 28946 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_52
timestamp 1624494425
transform 1 0 28941 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_133
timestamp 1624494425
transform 1 0 30109 0 1 -5397
box 0 0 76 66
use contact_9  contact_9_66
timestamp 1624494425
transform 1 0 30114 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_132
timestamp 1624494425
transform 1 0 30109 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_52
timestamp 1624494425
transform 1 0 32450 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_104
timestamp 1624494425
transform 1 0 32445 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_24
timestamp 1624494425
transform 1 0 31282 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_48
timestamp 1624494425
transform 1 0 31277 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_131
timestamp 1624494425
transform 1 0 33985 0 1 -5153
box 0 0 76 66
use contact_9  contact_9_22
timestamp 1624494425
transform 1 0 33618 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_44
timestamp 1624494425
transform 1 0 33613 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_125
timestamp 1624494425
transform 1 0 34781 0 1 -5153
box 0 0 76 66
use contact_9  contact_9_62
timestamp 1624494425
transform 1 0 34786 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_124
timestamp 1624494425
transform 1 0 34781 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_46
timestamp 1624494425
transform 1 0 35954 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_92
timestamp 1624494425
transform 1 0 35949 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_34
timestamp 1624494425
transform 1 0 37122 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_68
timestamp 1624494425
transform 1 0 37117 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 38290 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_40
timestamp 1624494425
transform 1 0 38285 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 39458 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_36
timestamp 1624494425
transform 1 0 39453 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 40626 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_28
timestamp 1624494425
transform 1 0 40621 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 41794 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_24
timestamp 1624494425
transform 1 0 41789 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 42962 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_16
timestamp 1624494425
transform 1 0 42957 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 44130 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_8
timestamp 1624494425
transform 1 0 44125 0 1 -6398
box 0 0 76 66
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 45298 0 1 -6402
box 0 0 66 74
use contact_32  contact_32_0
timestamp 1624494425
transform 1 0 45293 0 1 -6398
box 0 0 76 66
use contact_32  contact_32_123
timestamp 1624494425
transform 1 0 53953 0 1 -4909
box 0 0 76 66
use contact_32  contact_32_135
timestamp 1624494425
transform 1 0 59230 0 1 -5397
box 0 0 76 66
use contact_32  contact_32_127
timestamp 1624494425
transform 1 0 69214 0 1 -5153
box 0 0 76 66
use contact_32  contact_32_117
timestamp 1624494425
transform 1 0 7917 0 1 -4665
box 0 0 76 66
use contact_32  contact_32_113
timestamp 1624494425
transform 1 0 9085 0 1 -4421
box 0 0 76 66
use contact_32  contact_32_101
timestamp 1624494425
transform 1 0 10253 0 1 -4177
box 0 0 76 66
use contact_32  contact_32_89
timestamp 1624494425
transform 1 0 11421 0 1 -3933
box 0 0 76 66
use contact_32  contact_32_115
timestamp 1624494425
transform 1 0 14302 0 1 -4421
box 0 0 76 66
use contact_32  contact_32_81
timestamp 1624494425
transform 1 0 13757 0 1 -3689
box 0 0 76 66
use contact_32  contact_32_109
timestamp 1624494425
transform 1 0 17261 0 1 -4421
box 0 0 76 66
use contact_32  contact_32_103
timestamp 1624494425
transform 1 0 16798 0 1 -4177
box 0 0 76 66
use contact_32  contact_32_97
timestamp 1624494425
transform 1 0 18429 0 1 -4177
box 0 0 76 66
use contact_32  contact_32_91
timestamp 1624494425
transform 1 0 19294 0 1 -3933
box 0 0 76 66
use contact_32  contact_32_73
timestamp 1624494425
transform 1 0 19597 0 1 -3445
box 0 0 76 66
use contact_32  contact_32_85
timestamp 1624494425
transform 1 0 24269 0 1 -3933
box 0 0 76 66
use contact_32  contact_32_83
timestamp 1624494425
transform 1 0 24286 0 1 -3689
box 0 0 76 66
use contact_32  contact_32_77
timestamp 1624494425
transform 1 0 25437 0 1 -3689
box 0 0 76 66
use contact_32  contact_32_65
timestamp 1624494425
transform 1 0 26605 0 1 -3201
box 0 0 76 66
use contact_32  contact_32_111
timestamp 1624494425
transform 1 0 31774 0 1 -4421
box 0 0 76 66
use contact_32  contact_32_105
timestamp 1624494425
transform 1 0 32445 0 1 -4421
box 0 0 76 66
use contact_32  contact_32_99
timestamp 1624494425
transform 1 0 34270 0 1 -4177
box 0 0 76 66
use contact_32  contact_32_93
timestamp 1624494425
transform 1 0 35949 0 1 -4177
box 0 0 76 66
use contact_32  contact_32_75
timestamp 1624494425
transform 1 0 36766 0 1 -3445
box 0 0 76 66
use contact_32  contact_32_69
timestamp 1624494425
transform 1 0 37117 0 1 -3445
box 0 0 76 66
use contact_32  contact_32_87
timestamp 1624494425
transform 1 0 46750 0 1 -3933
box 0 0 76 66
use contact_32  contact_32_79
timestamp 1624494425
transform 1 0 49246 0 1 -3689
box 0 0 76 66
use contact_32  contact_32_67
timestamp 1624494425
transform 1 0 51742 0 1 -3201
box 0 0 76 66
use contact_32  contact_32_107
timestamp 1624494425
transform 1 0 64222 0 1 -4421
box 0 0 76 66
use contact_32  contact_32_95
timestamp 1624494425
transform 1 0 71710 0 1 -4177
box 0 0 76 66
use contact_32  contact_32_119
timestamp 1624494425
transform 1 0 73921 0 1 -4665
box 0 0 76 66
use contact_32  contact_32_71
timestamp 1624494425
transform 1 0 74206 0 1 -3445
box 0 0 76 66
use contact_32  contact_32_61
timestamp 1624494425
transform 1 0 14925 0 1 -2957
box 0 0 76 66
use contact_32  contact_32_33
timestamp 1624494425
transform 1 0 20765 0 1 -1493
box 0 0 76 66
use contact_32  contact_32_63
timestamp 1624494425
transform 1 0 26782 0 1 -2957
box 0 0 76 66
use contact_32  contact_32_57
timestamp 1624494425
transform 1 0 27773 0 1 -2957
box 0 0 76 66
use contact_32  contact_32_53
timestamp 1624494425
transform 1 0 28941 0 1 -2713
box 0 0 76 66
use contact_32  contact_32_49
timestamp 1624494425
transform 1 0 31277 0 1 -2469
box 0 0 76 66
use contact_32  contact_32_45
timestamp 1624494425
transform 1 0 33613 0 1 -2225
box 0 0 76 66
use contact_32  contact_32_41
timestamp 1624494425
transform 1 0 38285 0 1 -1981
box 0 0 76 66
use contact_32  contact_32_35
timestamp 1624494425
transform 1 0 39262 0 1 -1493
box 0 0 76 66
use contact_32  contact_32_37
timestamp 1624494425
transform 1 0 39453 0 1 -1737
box 0 0 76 66
use contact_32  contact_32_29
timestamp 1624494425
transform 1 0 40621 0 1 -1493
box 0 0 76 66
use contact_32  contact_32_59
timestamp 1624494425
transform 1 0 54238 0 1 -2957
box 0 0 76 66
use contact_32  contact_32_55
timestamp 1624494425
transform 1 0 56734 0 1 -2713
box 0 0 76 66
use contact_32  contact_32_51
timestamp 1624494425
transform 1 0 61726 0 1 -2469
box 0 0 76 66
use contact_32  contact_32_47
timestamp 1624494425
transform 1 0 66718 0 1 -2225
box 0 0 76 66
use contact_32  contact_32_43
timestamp 1624494425
transform 1 0 76702 0 1 -1981
box 0 0 76 66
use contact_32  contact_32_39
timestamp 1624494425
transform 1 0 79198 0 1 -1737
box 0 0 76 66
use contact_32  contact_32_31
timestamp 1624494425
transform 1 0 81694 0 1 -1493
box 0 0 76 66
use contact_32  contact_32_13
timestamp 1624494425
transform 1 0 12589 0 1 -761
box 0 0 76 66
use contact_32  contact_32_21
timestamp 1624494425
transform 1 0 21933 0 1 -1005
box 0 0 76 66
use contact_32  contact_32_15
timestamp 1624494425
transform 1 0 21790 0 1 -761
box 0 0 76 66
use contact_32  contact_32_5
timestamp 1624494425
transform 1 0 23101 0 1 -517
box 0 0 76 66
use contact_32  contact_32_25
timestamp 1624494425
transform 1 0 41789 0 1 -1249
box 0 0 76 66
use contact_32  contact_32_23
timestamp 1624494425
transform 1 0 41758 0 1 -1005
box 0 0 76 66
use contact_32  contact_32_17
timestamp 1624494425
transform 1 0 42957 0 1 -1005
box 0 0 76 66
use contact_32  contact_32_9
timestamp 1624494425
transform 1 0 44125 0 1 -761
box 0 0 76 66
use contact_32  contact_32_7
timestamp 1624494425
transform 1 0 44254 0 1 -517
box 0 0 76 66
use contact_32  contact_32_1
timestamp 1624494425
transform 1 0 45293 0 1 -517
box 0 0 76 66
use contact_32  contact_32_27
timestamp 1624494425
transform 1 0 84190 0 1 -1249
box 0 0 76 66
use contact_32  contact_32_19
timestamp 1624494425
transform 1 0 86686 0 1 -1005
box 0 0 76 66
use contact_32  contact_32_11
timestamp 1624494425
transform 1 0 89182 0 1 -761
box 0 0 76 66
use contact_32  contact_32_3
timestamp 1624494425
transform 1 0 91678 0 1 -517
box 0 0 76 66
use contact_9  contact_9_71
timestamp 1624494425
transform 1 0 14022 0 1 268
box 0 0 66 74
use contact_32  contact_32_142
timestamp 1624494425
transform 1 0 14017 0 1 272
box 0 0 76 66
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 14308 0 1 1393
box 0 0 64 64
use contact_9  contact_9_57
timestamp 1624494425
transform 1 0 14307 0 1 1388
box 0 0 66 74
use contact_32  contact_32_114
timestamp 1624494425
transform 1 0 14302 0 1 1392
box 0 0 76 66
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 16804 0 1 1393
box 0 0 64 64
use contact_9  contact_9_51
timestamp 1624494425
transform 1 0 16803 0 1 1388
box 0 0 66 74
use contact_32  contact_32_102
timestamp 1624494425
transform 1 0 16798 0 1 1392
box 0 0 76 66
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 19300 0 1 1393
box 0 0 64 64
use contact_9  contact_9_45
timestamp 1624494425
transform 1 0 19299 0 1 1388
box 0 0 66 74
use contact_32  contact_32_90
timestamp 1624494425
transform 1 0 19294 0 1 1392
box 0 0 76 66
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 21796 0 1 1393
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 21795 0 1 1388
box 0 0 66 74
use contact_32  contact_32_14
timestamp 1624494425
transform 1 0 21790 0 1 1392
box 0 0 76 66
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 24292 0 1 1393
box 0 0 64 64
use contact_9  contact_9_41
timestamp 1624494425
transform 1 0 24291 0 1 1388
box 0 0 66 74
use contact_32  contact_32_82
timestamp 1624494425
transform 1 0 24286 0 1 1392
box 0 0 76 66
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 26788 0 1 1393
box 0 0 64 64
use contact_9  contact_9_31
timestamp 1624494425
transform 1 0 26787 0 1 1388
box 0 0 66 74
use contact_32  contact_32_62
timestamp 1624494425
transform 1 0 26782 0 1 1392
box 0 0 76 66
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 29284 0 1 1393
box 0 0 64 64
use contact_9  contact_9_69
timestamp 1624494425
transform 1 0 29283 0 1 1388
box 0 0 66 74
use contact_32  contact_32_138
timestamp 1624494425
transform 1 0 29278 0 1 1392
box 0 0 76 66
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 31780 0 1 1393
box 0 0 64 64
use contact_9  contact_9_55
timestamp 1624494425
transform 1 0 31779 0 1 1388
box 0 0 66 74
use contact_32  contact_32_110
timestamp 1624494425
transform 1 0 31774 0 1 1392
box 0 0 76 66
use contact_9  contact_9_65
timestamp 1624494425
transform 1 0 33990 0 1 268
box 0 0 66 74
use contact_32  contact_32_130
timestamp 1624494425
transform 1 0 33985 0 1 272
box 0 0 76 66
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 34276 0 1 1393
box 0 0 64 64
use contact_9  contact_9_49
timestamp 1624494425
transform 1 0 34275 0 1 1388
box 0 0 66 74
use contact_32  contact_32_98
timestamp 1624494425
transform 1 0 34270 0 1 1392
box 0 0 76 66
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 36772 0 1 1393
box 0 0 64 64
use contact_9  contact_9_37
timestamp 1624494425
transform 1 0 36771 0 1 1388
box 0 0 66 74
use contact_32  contact_32_74
timestamp 1624494425
transform 1 0 36766 0 1 1392
box 0 0 76 66
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 39268 0 1 1393
box 0 0 64 64
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 39267 0 1 1388
box 0 0 66 74
use contact_32  contact_32_34
timestamp 1624494425
transform 1 0 39262 0 1 1392
box 0 0 76 66
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 41764 0 1 1393
box 0 0 64 64
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 41763 0 1 1388
box 0 0 66 74
use contact_32  contact_32_22
timestamp 1624494425
transform 1 0 41758 0 1 1392
box 0 0 76 66
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 44260 0 1 1393
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 44259 0 1 1388
box 0 0 66 74
use contact_32  contact_32_6
timestamp 1624494425
transform 1 0 44254 0 1 1392
box 0 0 76 66
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 46756 0 1 1393
box 0 0 64 64
use contact_9  contact_9_43
timestamp 1624494425
transform 1 0 46755 0 1 1388
box 0 0 66 74
use contact_32  contact_32_86
timestamp 1624494425
transform 1 0 46750 0 1 1392
box 0 0 76 66
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 49252 0 1 1393
box 0 0 64 64
use contact_9  contact_9_39
timestamp 1624494425
transform 1 0 49251 0 1 1388
box 0 0 66 74
use contact_32  contact_32_78
timestamp 1624494425
transform 1 0 49246 0 1 1392
box 0 0 76 66
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 51748 0 1 1393
box 0 0 64 64
use contact_9  contact_9_33
timestamp 1624494425
transform 1 0 51747 0 1 1388
box 0 0 66 74
use contact_32  contact_32_66
timestamp 1624494425
transform 1 0 51742 0 1 1392
box 0 0 76 66
use contact_9  contact_9_61
timestamp 1624494425
transform 1 0 53958 0 1 268
box 0 0 66 74
use contact_32  contact_32_122
timestamp 1624494425
transform 1 0 53953 0 1 272
box 0 0 76 66
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 54244 0 1 1393
box 0 0 64 64
use contact_9  contact_9_29
timestamp 1624494425
transform 1 0 54243 0 1 1388
box 0 0 66 74
use contact_32  contact_32_58
timestamp 1624494425
transform 1 0 54238 0 1 1392
box 0 0 76 66
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 56740 0 1 1393
box 0 0 64 64
use contact_9  contact_9_27
timestamp 1624494425
transform 1 0 56739 0 1 1388
box 0 0 66 74
use contact_32  contact_32_54
timestamp 1624494425
transform 1 0 56734 0 1 1392
box 0 0 76 66
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 59236 0 1 1393
box 0 0 64 64
use contact_9  contact_9_67
timestamp 1624494425
transform 1 0 59235 0 1 1388
box 0 0 66 74
use contact_32  contact_32_134
timestamp 1624494425
transform 1 0 59230 0 1 1392
box 0 0 76 66
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 61732 0 1 1393
box 0 0 64 64
use contact_9  contact_9_25
timestamp 1624494425
transform 1 0 61731 0 1 1388
box 0 0 66 74
use contact_32  contact_32_50
timestamp 1624494425
transform 1 0 61726 0 1 1392
box 0 0 76 66
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 64228 0 1 1393
box 0 0 64 64
use contact_9  contact_9_53
timestamp 1624494425
transform 1 0 64227 0 1 1388
box 0 0 66 74
use contact_32  contact_32_106
timestamp 1624494425
transform 1 0 64222 0 1 1392
box 0 0 76 66
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 66724 0 1 1393
box 0 0 64 64
use contact_9  contact_9_23
timestamp 1624494425
transform 1 0 66723 0 1 1388
box 0 0 66 74
use contact_32  contact_32_46
timestamp 1624494425
transform 1 0 66718 0 1 1392
box 0 0 76 66
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 69220 0 1 1393
box 0 0 64 64
use contact_9  contact_9_63
timestamp 1624494425
transform 1 0 69219 0 1 1388
box 0 0 66 74
use contact_32  contact_32_126
timestamp 1624494425
transform 1 0 69214 0 1 1392
box 0 0 76 66
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 71716 0 1 1393
box 0 0 64 64
use contact_9  contact_9_47
timestamp 1624494425
transform 1 0 71715 0 1 1388
box 0 0 66 74
use contact_32  contact_32_94
timestamp 1624494425
transform 1 0 71710 0 1 1392
box 0 0 76 66
use contact_9  contact_9_59
timestamp 1624494425
transform 1 0 73926 0 1 268
box 0 0 66 74
use contact_32  contact_32_118
timestamp 1624494425
transform 1 0 73921 0 1 272
box 0 0 76 66
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 74212 0 1 1393
box 0 0 64 64
use contact_9  contact_9_35
timestamp 1624494425
transform 1 0 74211 0 1 1388
box 0 0 66 74
use contact_32  contact_32_70
timestamp 1624494425
transform 1 0 74206 0 1 1392
box 0 0 76 66
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 76708 0 1 1393
box 0 0 64 64
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 76707 0 1 1388
box 0 0 66 74
use contact_32  contact_32_42
timestamp 1624494425
transform 1 0 76702 0 1 1392
box 0 0 76 66
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 79204 0 1 1393
box 0 0 64 64
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 79203 0 1 1388
box 0 0 66 74
use contact_32  contact_32_38
timestamp 1624494425
transform 1 0 79198 0 1 1392
box 0 0 76 66
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 81700 0 1 1393
box 0 0 64 64
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 81699 0 1 1388
box 0 0 66 74
use contact_32  contact_32_30
timestamp 1624494425
transform 1 0 81694 0 1 1392
box 0 0 76 66
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 84196 0 1 1393
box 0 0 64 64
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 84195 0 1 1388
box 0 0 66 74
use contact_32  contact_32_26
timestamp 1624494425
transform 1 0 84190 0 1 1392
box 0 0 76 66
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 86692 0 1 1393
box 0 0 64 64
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 86691 0 1 1388
box 0 0 66 74
use contact_32  contact_32_18
timestamp 1624494425
transform 1 0 86686 0 1 1392
box 0 0 76 66
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 89188 0 1 1393
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 89187 0 1 1388
box 0 0 66 74
use contact_32  contact_32_10
timestamp 1624494425
transform 1 0 89182 0 1 1392
box 0 0 76 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 91684 0 1 1393
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 91683 0 1 1388
box 0 0 66 74
use contact_32  contact_32_2
timestamp 1624494425
transform 1 0 91678 0 1 1392
box 0 0 76 66
<< properties >>
string FIXED_BBOX 4376 -6402 91791 1462
<< end >>
