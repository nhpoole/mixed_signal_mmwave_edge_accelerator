magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2003 -1602 2003 1604
<< nwell >>
rect -731 248 743 344
rect -743 -342 743 248
<< pmoslvt >>
rect -547 -100 -477 100
rect -419 -100 -349 100
rect -291 -100 -221 100
rect -163 -100 -93 100
rect -35 -100 35 100
rect 93 -100 163 100
rect 221 -100 291 100
rect 349 -100 419 100
rect 477 -100 547 100
<< pdiff >>
rect -605 85 -547 100
rect -605 51 -593 85
rect -559 51 -547 85
rect -605 17 -547 51
rect -605 -17 -593 17
rect -559 -17 -547 17
rect -605 -51 -547 -17
rect -605 -85 -593 -51
rect -559 -85 -547 -51
rect -605 -100 -547 -85
rect -477 85 -419 100
rect -477 51 -465 85
rect -431 51 -419 85
rect -477 17 -419 51
rect -477 -17 -465 17
rect -431 -17 -419 17
rect -477 -51 -419 -17
rect -477 -85 -465 -51
rect -431 -85 -419 -51
rect -477 -100 -419 -85
rect -349 85 -291 100
rect -349 51 -337 85
rect -303 51 -291 85
rect -349 17 -291 51
rect -349 -17 -337 17
rect -303 -17 -291 17
rect -349 -51 -291 -17
rect -349 -85 -337 -51
rect -303 -85 -291 -51
rect -349 -100 -291 -85
rect -221 85 -163 100
rect -221 51 -209 85
rect -175 51 -163 85
rect -221 17 -163 51
rect -221 -17 -209 17
rect -175 -17 -163 17
rect -221 -51 -163 -17
rect -221 -85 -209 -51
rect -175 -85 -163 -51
rect -221 -100 -163 -85
rect -93 85 -35 100
rect -93 51 -81 85
rect -47 51 -35 85
rect -93 17 -35 51
rect -93 -17 -81 17
rect -47 -17 -35 17
rect -93 -51 -35 -17
rect -93 -85 -81 -51
rect -47 -85 -35 -51
rect -93 -100 -35 -85
rect 35 85 93 100
rect 35 51 47 85
rect 81 51 93 85
rect 35 17 93 51
rect 35 -17 47 17
rect 81 -17 93 17
rect 35 -51 93 -17
rect 35 -85 47 -51
rect 81 -85 93 -51
rect 35 -100 93 -85
rect 163 85 221 100
rect 163 51 175 85
rect 209 51 221 85
rect 163 17 221 51
rect 163 -17 175 17
rect 209 -17 221 17
rect 163 -51 221 -17
rect 163 -85 175 -51
rect 209 -85 221 -51
rect 163 -100 221 -85
rect 291 85 349 100
rect 291 51 303 85
rect 337 51 349 85
rect 291 17 349 51
rect 291 -17 303 17
rect 337 -17 349 17
rect 291 -51 349 -17
rect 291 -85 303 -51
rect 337 -85 349 -51
rect 291 -100 349 -85
rect 419 85 477 100
rect 419 51 431 85
rect 465 51 477 85
rect 419 17 477 51
rect 419 -17 431 17
rect 465 -17 477 17
rect 419 -51 477 -17
rect 419 -85 431 -51
rect 465 -85 477 -51
rect 419 -100 477 -85
rect 547 85 605 100
rect 547 51 559 85
rect 593 51 605 85
rect 547 17 605 51
rect 547 -17 559 17
rect 593 -17 605 17
rect 547 -51 605 -17
rect 547 -85 559 -51
rect 593 -85 605 -51
rect 547 -100 605 -85
<< pdiffc >>
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -465 51 -431 85
rect -465 -17 -431 17
rect -465 -85 -431 -51
rect -337 51 -303 85
rect -337 -17 -303 17
rect -337 -85 -303 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -81 51 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -51
rect 47 51 81 85
rect 47 -17 81 17
rect 47 -85 81 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 303 51 337 85
rect 303 -17 337 17
rect 303 -85 337 -51
rect 431 51 465 85
rect 431 -17 465 17
rect 431 -85 465 -51
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
<< nsubdiff >>
rect -707 276 -595 310
rect -561 276 -527 310
rect -493 276 -459 310
rect -425 276 -391 310
rect -357 276 -323 310
rect -289 276 -255 310
rect -221 276 -187 310
rect -153 276 -119 310
rect -85 276 -51 310
rect -17 276 17 310
rect 51 276 85 310
rect 119 276 153 310
rect 187 276 221 310
rect 255 276 289 310
rect 323 276 357 310
rect 391 276 425 310
rect 459 276 493 310
rect 527 276 561 310
rect 595 276 707 310
rect -707 85 -673 276
rect -707 17 -673 51
rect -707 -51 -673 -17
rect -707 -272 -673 -85
rect 673 85 707 276
rect 673 17 707 51
rect 673 -51 707 -17
rect 673 -272 707 -85
rect -707 -306 -595 -272
rect -561 -306 -527 -272
rect -493 -306 -459 -272
rect -425 -306 -391 -272
rect -357 -306 -323 -272
rect -289 -306 -255 -272
rect -221 -306 -187 -272
rect -153 -306 -119 -272
rect -85 -306 -51 -272
rect -17 -306 17 -272
rect 51 -306 85 -272
rect 119 -306 153 -272
rect 187 -306 221 -272
rect 255 -306 289 -272
rect 323 -306 357 -272
rect 391 -306 425 -272
rect 459 -306 493 -272
rect 527 -306 561 -272
rect 595 -306 707 -272
<< nsubdiffcont >>
rect -595 276 -561 310
rect -527 276 -493 310
rect -459 276 -425 310
rect -391 276 -357 310
rect -323 276 -289 310
rect -255 276 -221 310
rect -187 276 -153 310
rect -119 276 -85 310
rect -51 276 -17 310
rect 17 276 51 310
rect 85 276 119 310
rect 153 276 187 310
rect 221 276 255 310
rect 289 276 323 310
rect 357 276 391 310
rect 425 276 459 310
rect 493 276 527 310
rect 561 276 595 310
rect -707 51 -673 85
rect -707 -17 -673 17
rect -707 -85 -673 -51
rect 673 51 707 85
rect 673 -17 707 17
rect 673 -85 707 -51
rect -595 -306 -561 -272
rect -527 -306 -493 -272
rect -459 -306 -425 -272
rect -391 -306 -357 -272
rect -323 -306 -289 -272
rect -255 -306 -221 -272
rect -187 -306 -153 -272
rect -119 -306 -85 -272
rect -51 -306 -17 -272
rect 17 -306 51 -272
rect 85 -306 119 -272
rect 153 -306 187 -272
rect 221 -306 255 -272
rect 289 -306 323 -272
rect 357 -306 391 -272
rect 425 -306 459 -272
rect 493 -306 527 -272
rect 561 -306 595 -272
<< poly >>
rect -547 100 -477 126
rect -419 100 -349 126
rect -291 100 -221 126
rect -163 100 -93 126
rect -35 100 35 126
rect 93 100 163 126
rect 221 100 291 126
rect 349 100 419 126
rect 477 100 547 126
rect -547 -126 -477 -100
rect -419 -126 -349 -100
rect -291 -126 -221 -100
rect -163 -126 -93 -100
rect -35 -126 35 -100
rect 93 -126 163 -100
rect 221 -126 291 -100
rect 349 -126 419 -100
rect 477 -126 547 -100
<< locali >>
rect -707 276 -595 310
rect -561 276 -527 310
rect -493 276 -459 310
rect -425 276 -391 310
rect -357 276 -323 310
rect -289 276 -255 310
rect -221 276 -187 310
rect -153 276 -119 310
rect -85 276 -51 310
rect -17 276 17 310
rect 51 276 85 310
rect 119 276 153 310
rect 187 276 221 310
rect 255 276 289 310
rect 323 276 357 310
rect 391 276 425 310
rect 459 276 493 310
rect 527 276 561 310
rect 595 276 707 310
rect -707 85 -673 276
rect -707 17 -673 51
rect -707 -51 -673 -17
rect -707 -272 -673 -85
rect -593 85 -559 104
rect -593 17 -559 19
rect -593 -19 -559 -17
rect -593 -104 -559 -85
rect -465 85 -431 104
rect -465 17 -431 19
rect -465 -19 -431 -17
rect -465 -104 -431 -85
rect -337 85 -303 104
rect -337 17 -303 19
rect -337 -19 -303 -17
rect -337 -104 -303 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -81 85 -47 104
rect -81 17 -47 19
rect -81 -19 -47 -17
rect -81 -104 -47 -85
rect 47 85 81 104
rect 47 17 81 19
rect 47 -19 81 -17
rect 47 -104 81 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 303 85 337 104
rect 303 17 337 19
rect 303 -19 337 -17
rect 303 -104 337 -85
rect 431 85 465 104
rect 431 17 465 19
rect 431 -19 465 -17
rect 431 -104 465 -85
rect 559 85 593 104
rect 559 17 593 19
rect 559 -19 593 -17
rect 559 -104 593 -85
rect 673 85 707 276
rect 673 17 707 51
rect 673 -51 707 -17
rect 673 -272 707 -85
rect -707 -306 -595 -272
rect -561 -306 -527 -272
rect -493 -306 -459 -272
rect -425 -306 -391 -272
rect -357 -306 -323 -272
rect -289 -306 -255 -272
rect -221 -306 -187 -272
rect -153 -306 -119 -272
rect -85 -306 -51 -272
rect -17 -306 17 -272
rect 51 -306 85 -272
rect 119 -306 153 -272
rect 187 -306 221 -272
rect 255 -306 289 -272
rect 323 -306 357 -272
rect 391 -306 425 -272
rect 459 -306 493 -272
rect 527 -306 561 -272
rect 595 -306 707 -272
<< viali >>
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -465 51 -431 53
rect -465 19 -431 51
rect -465 -51 -431 -19
rect -465 -53 -431 -51
rect -337 51 -303 53
rect -337 19 -303 51
rect -337 -51 -303 -19
rect -337 -53 -303 -51
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -81 51 -47 53
rect -81 19 -47 51
rect -81 -51 -47 -19
rect -81 -53 -47 -51
rect 47 51 81 53
rect 47 19 81 51
rect 47 -51 81 -19
rect 47 -53 81 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 303 51 337 53
rect 303 19 337 51
rect 303 -51 337 -19
rect 303 -53 337 -51
rect 431 51 465 53
rect 431 19 465 51
rect 431 -51 465 -19
rect 431 -53 465 -51
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
<< metal1 >>
rect -599 53 -553 100
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -100 -553 -53
rect -471 53 -425 100
rect -471 19 -465 53
rect -431 19 -425 53
rect -471 -19 -425 19
rect -471 -53 -465 -19
rect -431 -53 -425 -19
rect -471 -100 -425 -53
rect -343 53 -297 100
rect -343 19 -337 53
rect -303 19 -297 53
rect -343 -19 -297 19
rect -343 -53 -337 -19
rect -303 -53 -297 -19
rect -343 -100 -297 -53
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -87 53 -41 100
rect -87 19 -81 53
rect -47 19 -41 53
rect -87 -19 -41 19
rect -87 -53 -81 -19
rect -47 -53 -41 -19
rect -87 -100 -41 -53
rect 41 53 87 100
rect 41 19 47 53
rect 81 19 87 53
rect 41 -19 87 19
rect 41 -53 47 -19
rect 81 -53 87 -19
rect 41 -100 87 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect 297 53 343 100
rect 297 19 303 53
rect 337 19 343 53
rect 297 -19 343 19
rect 297 -53 303 -19
rect 337 -53 343 -19
rect 297 -100 343 -53
rect 425 53 471 100
rect 425 19 431 53
rect 465 19 471 53
rect 425 -19 471 19
rect 425 -53 431 -19
rect 465 -53 471 -19
rect 425 -100 471 -53
rect 553 53 599 100
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -100 599 -53
<< properties >>
string FIXED_BBOX -690 -195 690 195
<< end >>
