magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< nwell >>
rect -398 -7578 12658 2958
<< pwell >>
rect -398 -10858 12658 -7742
<< psubdiff >>
rect -362 -7878 -200 -7778
rect 12460 -7878 12622 -7778
rect -362 -7940 -262 -7878
rect -362 -10722 -262 -10660
rect 12522 -7940 12622 -7878
rect 12522 -10722 12622 -10660
rect -362 -10822 -200 -10722
rect 12460 -10822 12622 -10722
<< nsubdiff >>
rect -362 2822 -200 2922
rect 12460 2822 12622 2922
rect -362 2760 -262 2822
rect -362 -7442 -262 -7380
rect 12522 2760 12622 2822
rect 12522 -7442 12622 -7380
rect -362 -7542 -200 -7442
rect 12460 -7542 12622 -7442
<< psubdiffcont >>
rect -200 -7878 12460 -7778
rect -362 -10660 -262 -7940
rect 12522 -10660 12622 -7940
rect -200 -10822 12460 -10722
<< nsubdiffcont >>
rect -200 2822 12460 2922
rect -362 -7380 -262 2760
rect 12522 -7380 12622 2760
rect -200 -7542 12460 -7442
<< locali >>
rect -362 2760 -262 2922
rect -362 -7542 -262 -7380
rect 12522 2760 12622 2922
rect 12522 -7542 12622 -7380
rect -362 -7940 -262 -7778
rect -362 -10822 -262 -10660
rect 12522 -7940 12622 -7778
rect 12522 -10822 12622 -10660
<< viali >>
rect -262 2822 -200 2922
rect -200 2822 12460 2922
rect 12460 2822 12522 2922
rect -362 -7119 -262 2299
rect 12522 -7119 12622 2299
rect -262 -7542 -200 -7442
rect -200 -7542 12460 -7442
rect 12460 -7542 12522 -7442
rect -262 -7878 -200 -7778
rect -200 -7878 12460 -7778
rect 12460 -7878 12522 -7778
rect -362 -10570 -262 -7982
rect 12522 -10570 12622 -7982
rect -262 -10822 -200 -10722
rect -200 -10822 12460 -10722
rect 12460 -10822 12522 -10722
<< metal1 >>
rect -368 2922 12628 2928
rect -368 2822 -262 2922
rect 12522 2822 12628 2922
rect -368 2816 12628 2822
rect -368 2299 -256 2816
rect 344 2516 354 2816
rect 11906 2516 11916 2816
rect -368 -7119 -362 2299
rect -262 2108 -256 2299
rect 110 2396 12310 2438
rect 110 2232 158 2396
rect 12268 2232 12310 2396
rect 110 2192 12310 2232
rect 12516 2299 12628 2816
rect 172 2110 232 2192
rect 596 2110 656 2192
rect 1032 2110 1092 2192
rect 2746 2110 2806 2192
rect 4466 2110 4526 2192
rect 6174 2110 6234 2192
rect 7894 2110 7954 2192
rect 9608 2110 9668 2192
rect 11326 2110 11386 2192
rect 11754 2110 11814 2192
rect 12186 2110 12246 2192
rect 166 2108 172 2110
rect -262 2050 172 2108
rect 232 2050 238 2110
rect 590 2050 596 2110
rect 656 2050 662 2110
rect 1026 2050 1032 2110
rect 1092 2050 1098 2110
rect 2740 2050 2746 2110
rect 2806 2050 2812 2110
rect 4460 2050 4466 2110
rect 4526 2050 4532 2110
rect 6168 2050 6174 2110
rect 6234 2050 6240 2110
rect 7888 2050 7894 2110
rect 7954 2050 7960 2110
rect 9602 2050 9608 2110
rect 9668 2050 9674 2110
rect 11320 2050 11326 2110
rect 11386 2050 11392 2110
rect 11748 2050 11754 2110
rect 11814 2050 11820 2110
rect 12180 2050 12186 2110
rect 12246 2108 12252 2110
rect 12516 2108 12522 2299
rect 12246 2050 12522 2108
rect -262 2048 232 2050
rect -262 -5150 -256 2048
rect -98 1786 -92 1846
rect -32 1786 -26 1846
rect -92 -50 -32 1786
rect 44 1658 50 1718
rect 110 1658 116 1718
rect 50 56 110 1658
rect 172 1414 232 2048
rect 596 1550 656 2050
rect 1032 1414 1092 2050
rect 1452 1922 1458 1982
rect 1518 1922 1524 1982
rect 2306 1922 2312 1982
rect 2372 1922 2378 1982
rect 1458 1550 1518 1922
rect 2312 1556 2372 1922
rect 2746 1422 2806 2050
rect 3166 1922 3172 1982
rect 3232 1922 3238 1982
rect 4026 1922 4032 1982
rect 4092 1922 4098 1982
rect 3172 1556 3232 1922
rect 4032 1556 4092 1922
rect 4466 1436 4526 2050
rect 4886 1922 4892 1982
rect 4952 1922 4958 1982
rect 5746 1922 5752 1982
rect 5812 1922 5818 1982
rect 4892 1556 4952 1922
rect 5752 1556 5812 1922
rect 6174 1436 6234 2050
rect 6606 1922 6612 1982
rect 6672 1922 6678 1982
rect 7466 1922 7472 1982
rect 7532 1922 7538 1982
rect 6612 1556 6672 1922
rect 7472 1556 7532 1922
rect 7894 1416 7954 2050
rect 8326 1922 8332 1982
rect 8392 1922 8398 1982
rect 9166 1922 9172 1982
rect 9232 1922 9238 1982
rect 8332 1556 8392 1922
rect 8746 1658 8752 1718
rect 8812 1658 8818 1718
rect 8752 1342 8812 1658
rect 9172 1556 9232 1922
rect 9608 1414 9668 2050
rect 10024 1922 10030 1982
rect 10090 1922 10096 1982
rect 10886 1922 10892 1982
rect 10952 1922 10958 1982
rect 10030 1548 10090 1922
rect 10462 1786 10468 1846
rect 10528 1786 10534 1846
rect 10468 1356 10528 1786
rect 10892 1548 10952 1922
rect 11326 1432 11386 2050
rect 11754 1544 11814 2050
rect 12186 2048 12522 2050
rect 12186 1418 12246 2048
rect 170 62 230 394
rect 600 62 660 252
rect 1030 62 1090 396
rect 44 -4 50 56
rect 110 -4 116 56
rect 170 -6 1090 62
rect -98 -110 -92 -50
rect -32 -110 -26 -50
rect -98 -1640 -92 -1580
rect -32 -1640 -26 -1580
rect -92 -3530 -32 -1640
rect 170 -1682 230 -6
rect 600 -195 660 -6
rect 600 -1682 660 -1482
rect 1030 -1682 1090 -6
rect 1460 -195 1520 252
rect 1888 156 1948 454
rect 1882 96 1888 156
rect 1948 96 1954 156
rect 1884 -110 1890 -50
rect 1950 -110 1956 -50
rect 1890 -298 1950 -110
rect 2320 -195 2380 252
rect 1460 -1678 1520 -1482
rect 170 -1742 1090 -1682
rect 44 -1846 50 -1786
rect 110 -1846 116 -1786
rect 50 -3424 110 -1846
rect 170 -3424 230 -1742
rect 600 -1929 660 -1742
rect 600 -3424 660 -3222
rect 1030 -3424 1090 -1742
rect 1458 -1684 1520 -1678
rect 1518 -1744 1520 -1684
rect 1458 -1750 1520 -1744
rect 1460 -1929 1520 -1750
rect 2320 -1684 2380 -1482
rect 2320 -1929 2380 -1744
rect 44 -3484 50 -3424
rect 110 -3484 116 -3424
rect 170 -3484 1090 -3424
rect -98 -3590 -92 -3530
rect -32 -3590 -26 -3530
rect 170 -5150 230 -3484
rect 600 -3669 660 -3484
rect 600 -5150 660 -4964
rect 1030 -5150 1090 -3484
rect 1460 -3669 1520 -3222
rect 1888 -3324 1948 -3026
rect 1882 -3384 1888 -3324
rect 1948 -3384 1954 -3324
rect 1884 -3590 1890 -3530
rect 1950 -3590 1956 -3530
rect 1890 -3778 1950 -3590
rect 2320 -3669 2380 -3222
rect 1460 -5050 1520 -4964
rect 2320 -5050 2380 -4964
rect 1454 -5110 1460 -5050
rect 1520 -5110 1526 -5050
rect -262 -5210 1090 -5150
rect -262 -7076 -256 -5210
rect 170 -7070 230 -5210
rect 600 -5411 660 -5210
rect 1030 -5542 1090 -5210
rect 1460 -5411 1520 -5110
rect 1882 -5328 1888 -5268
rect 1948 -5328 1954 -5268
rect 1888 -5580 1948 -5328
rect 2320 -5411 2380 -5110
rect 590 -7070 650 -6700
rect 1030 -7070 1090 -6548
rect 1456 -6926 1516 -6700
rect 2326 -6926 2386 -6697
rect 1450 -6986 1456 -6926
rect 1516 -6986 1522 -6926
rect 2320 -6986 2326 -6926
rect 2386 -6986 2392 -6926
rect 2748 -7070 2808 388
rect 3180 -195 3240 252
rect 3464 -4 3470 56
rect 3530 -4 3536 56
rect 3604 54 3664 360
rect 3470 -48 3530 -4
rect 3598 -6 3604 54
rect 3664 -6 3670 54
rect 3470 -108 3664 -48
rect 3604 -312 3664 -108
rect 4040 -195 4100 252
rect 3180 -1678 3240 -1482
rect 3180 -1684 3242 -1678
rect 3180 -1744 3182 -1684
rect 3180 -1750 3242 -1744
rect 4040 -1684 4100 -1482
rect 3180 -1929 3240 -1750
rect 4040 -1929 4100 -1744
rect 3180 -3669 3240 -3222
rect 3464 -3484 3470 -3424
rect 3530 -3484 3536 -3424
rect 3604 -3426 3664 -3120
rect 3470 -3528 3530 -3484
rect 3598 -3486 3604 -3426
rect 3664 -3486 3670 -3426
rect 3470 -3588 3664 -3528
rect 3604 -3792 3664 -3588
rect 4040 -3669 4100 -3222
rect 4462 -3532 4522 386
rect 4900 -195 4960 252
rect 5318 54 5378 420
rect 7038 156 7098 368
rect 7038 96 7226 156
rect 5318 -6 7096 54
rect 5314 -110 5320 -50
rect 5380 -110 5386 -50
rect 5320 -406 5380 -110
rect 7036 -112 7096 -6
rect 7166 -50 7226 96
rect 7160 -110 7166 -50
rect 7226 -110 7232 -50
rect 7036 -280 7098 -112
rect 7480 -195 7540 252
rect 7038 -294 7098 -280
rect 4900 -1684 4960 -1482
rect 4900 -1929 4960 -1744
rect 5744 -1684 5804 -1485
rect 5744 -1936 5804 -1744
rect 3180 -5044 3240 -4964
rect 3176 -5050 3240 -5044
rect 3236 -5110 3240 -5050
rect 3176 -5116 3240 -5110
rect 3180 -5411 3240 -5116
rect 4040 -5044 4100 -4964
rect 4040 -5050 4102 -5044
rect 4040 -5110 4042 -5050
rect 4040 -5116 4102 -5110
rect 3600 -5214 3606 -5154
rect 3666 -5214 3672 -5154
rect 3606 -5520 3666 -5214
rect 4040 -5411 4100 -5116
rect 3184 -6926 3244 -6697
rect 4042 -6926 4102 -6697
rect 3178 -6986 3184 -6926
rect 3244 -6986 3250 -6926
rect 4036 -6986 4042 -6926
rect 4102 -6986 4108 -6926
rect 4462 -7070 4522 -3592
rect 4900 -3669 4960 -3222
rect 5318 -3426 5378 -3060
rect 6180 -3196 6240 -332
rect 6614 -1684 6674 -1481
rect 6614 -1932 6674 -1744
rect 7480 -1684 7540 -1482
rect 7480 -1929 7540 -1744
rect 6180 -3262 6240 -3256
rect 7038 -3324 7098 -3112
rect 7038 -3384 7226 -3324
rect 5318 -3486 7096 -3426
rect 5314 -3590 5320 -3530
rect 5380 -3590 5386 -3530
rect 5320 -3886 5380 -3590
rect 7036 -3592 7096 -3486
rect 7166 -3530 7226 -3384
rect 7160 -3590 7166 -3530
rect 7226 -3590 7232 -3530
rect 7036 -3760 7098 -3592
rect 7480 -3669 7540 -3222
rect 7894 -3530 7954 384
rect 8336 -195 8396 252
rect 8750 -6 8756 54
rect 8816 -6 8822 54
rect 8756 -340 8816 -6
rect 9192 -195 9252 252
rect 8336 -1684 8396 -1482
rect 8336 -1929 8396 -1744
rect 9192 -1684 9252 -1482
rect 8746 -1846 8752 -1786
rect 8812 -1846 8818 -1786
rect 8752 -2138 8812 -1846
rect 9192 -1929 9252 -1744
rect 7038 -3774 7098 -3760
rect 4900 -5044 4960 -4964
rect 4898 -5050 4960 -5044
rect 4958 -5110 4960 -5050
rect 4898 -5116 4960 -5110
rect 4900 -5411 4960 -5116
rect 5742 -5044 5802 -4967
rect 5742 -5050 5806 -5044
rect 5742 -5110 5746 -5050
rect 5742 -5116 5806 -5110
rect 5742 -5418 5802 -5116
rect 4900 -6926 4960 -6697
rect 5320 -6800 5380 -6540
rect 5314 -6860 5320 -6800
rect 5380 -6860 5386 -6800
rect 5758 -6926 5818 -6697
rect 4894 -6986 4900 -6926
rect 4960 -6986 4966 -6926
rect 5752 -6986 5758 -6926
rect 5818 -6986 5824 -6926
rect 6180 -7070 6240 -3788
rect 6602 -5044 6662 -4959
rect 6600 -5050 6662 -5044
rect 6660 -5110 6662 -5050
rect 6600 -5116 6662 -5110
rect 6602 -5410 6662 -5116
rect 7480 -5050 7540 -4964
rect 7480 -5411 7540 -5110
rect 6616 -6926 6676 -6697
rect 7038 -6800 7098 -6602
rect 7032 -6860 7038 -6800
rect 7098 -6860 7104 -6800
rect 7474 -6926 7534 -6697
rect 6610 -6986 6616 -6926
rect 6676 -6986 6682 -6926
rect 7468 -6986 7474 -6926
rect 7534 -6986 7540 -6926
rect 7894 -7070 7954 -3590
rect 8336 -3669 8396 -3222
rect 8750 -3486 8756 -3426
rect 8816 -3486 8822 -3426
rect 8756 -3820 8816 -3486
rect 9192 -3669 9252 -3222
rect 8336 -5044 8396 -4964
rect 8334 -5050 8396 -5044
rect 8394 -5110 8396 -5050
rect 8334 -5116 8396 -5110
rect 8336 -5411 8396 -5116
rect 9192 -5054 9252 -4964
rect 8746 -5214 8752 -5154
rect 8812 -5214 8818 -5154
rect 8752 -5518 8812 -5214
rect 9192 -5411 9252 -5114
rect 8332 -6926 8392 -6697
rect 9190 -6926 9250 -6697
rect 8326 -6986 8332 -6926
rect 8392 -6986 8398 -6926
rect 9184 -6986 9190 -6926
rect 9250 -6986 9256 -6926
rect 9608 -7070 9668 390
rect 10048 -195 10108 252
rect 10464 96 10470 156
rect 10530 96 10536 156
rect 10470 -304 10530 96
rect 10904 -190 10964 252
rect 11326 66 11386 406
rect 11750 66 11810 255
rect 12184 66 12244 394
rect 12516 66 12522 2048
rect 11326 6 12522 66
rect 10048 -1678 10108 -1482
rect 10462 -1640 10468 -1580
rect 10528 -1640 10534 -1580
rect 10046 -1684 10108 -1678
rect 10106 -1744 10108 -1684
rect 10046 -1750 10108 -1744
rect 10048 -1929 10108 -1750
rect 10468 -2124 10528 -1640
rect 10904 -1684 10964 -1482
rect 11326 -1680 11386 6
rect 11750 -196 11810 6
rect 11754 -1680 11814 -1481
rect 12184 -1680 12244 6
rect 12516 -1680 12522 6
rect 10898 -1744 10904 -1684
rect 10964 -1744 10970 -1684
rect 11326 -1740 12522 -1680
rect 10904 -1929 10964 -1744
rect 10048 -3669 10108 -3222
rect 10464 -3384 10470 -3324
rect 10530 -3384 10536 -3324
rect 10470 -3784 10530 -3384
rect 10904 -3669 10964 -3222
rect 11326 -3412 11386 -1740
rect 11754 -1932 11814 -1740
rect 11750 -3412 11810 -3223
rect 12184 -3412 12244 -1740
rect 12516 -3412 12522 -1740
rect 11326 -3472 12522 -3412
rect 10048 -5050 10108 -4964
rect 10048 -5411 10108 -5110
rect 10904 -5044 10964 -4964
rect 10904 -5050 10966 -5044
rect 10904 -5110 10906 -5050
rect 10904 -5116 10966 -5110
rect 10464 -5328 10470 -5268
rect 10530 -5328 10536 -5268
rect 10470 -5518 10530 -5328
rect 10904 -5411 10964 -5116
rect 11326 -5154 11386 -3472
rect 11750 -3674 11810 -3472
rect 11754 -5154 11814 -4959
rect 12184 -5154 12244 -3472
rect 12516 -5154 12522 -3472
rect 11326 -5214 12522 -5154
rect 11326 -5572 11386 -5214
rect 11754 -5410 11814 -5214
rect 12184 -5568 12244 -5214
rect 10048 -6926 10108 -6697
rect 10904 -6926 10964 -6700
rect 10042 -6986 10048 -6926
rect 10108 -6986 10114 -6926
rect 10898 -6986 10904 -6926
rect 10964 -6986 10970 -6926
rect 11324 -7070 11384 -6594
rect 11750 -7070 11810 -6704
rect 12184 -7070 12244 -6588
rect 164 -7076 170 -7070
rect -262 -7119 170 -7076
rect -368 -7130 170 -7119
rect 230 -7130 236 -7070
rect 584 -7130 590 -7070
rect 650 -7130 656 -7070
rect 1024 -7130 1030 -7070
rect 1090 -7130 1096 -7070
rect 2742 -7130 2748 -7070
rect 2808 -7130 2814 -7070
rect 4456 -7130 4462 -7070
rect 4522 -7130 4528 -7070
rect 6174 -7130 6180 -7070
rect 6240 -7130 6246 -7070
rect 7888 -7130 7894 -7070
rect 7954 -7130 7960 -7070
rect 9602 -7130 9608 -7070
rect 9668 -7130 9674 -7070
rect 11318 -7130 11324 -7070
rect 11384 -7130 11390 -7070
rect 11744 -7130 11750 -7070
rect 11810 -7130 11816 -7070
rect 12178 -7130 12184 -7070
rect 12244 -7072 12250 -7070
rect 12516 -7072 12522 -5214
rect 12244 -7119 12522 -7072
rect 12622 -7119 12628 2299
rect 12244 -7130 12628 -7119
rect -368 -7136 230 -7130
rect -368 -7436 -256 -7136
rect 170 -7436 230 -7136
rect 590 -7436 650 -7130
rect 1030 -7436 1090 -7130
rect 2748 -7436 2808 -7130
rect 4462 -7436 4522 -7130
rect 6180 -7436 6240 -7130
rect 7894 -7436 7954 -7130
rect 9608 -7436 9668 -7130
rect 11324 -7436 11384 -7130
rect 11750 -7436 11810 -7130
rect 12184 -7132 12628 -7130
rect 12184 -7436 12244 -7132
rect 12516 -7436 12628 -7132
rect -368 -7442 12628 -7436
rect -368 -7542 -262 -7442
rect 12522 -7542 12628 -7442
rect -368 -7548 12628 -7542
rect -368 -7778 12628 -7772
rect -368 -7878 -262 -7778
rect 12522 -7878 12628 -7778
rect -368 -7884 12628 -7878
rect -368 -7982 -256 -7884
rect -368 -10570 -362 -7982
rect -262 -10570 -256 -7982
rect 4792 -8222 4798 -8162
rect 4858 -8222 4864 -8162
rect 4798 -9092 4858 -8222
rect 4896 -8272 4956 -7884
rect 5124 -8272 5184 -7884
rect 4896 -8332 5184 -8272
rect 5576 -8330 5582 -8270
rect 5642 -8330 5648 -8270
rect 4896 -9032 4956 -8332
rect 5124 -8420 5184 -8332
rect 5582 -8424 5642 -8330
rect 5124 -9032 5184 -8892
rect 5356 -8978 5416 -8826
rect 4896 -9092 5184 -9032
rect 5350 -9038 5356 -8978
rect 5416 -9038 5422 -8978
rect 4792 -9152 4798 -9092
rect 4858 -9152 4864 -9092
rect 4896 -9794 4956 -9092
rect 5124 -9228 5184 -9092
rect 5350 -9152 5356 -9092
rect 5416 -9152 5422 -9092
rect 5356 -9316 5416 -9152
rect 5584 -9224 5644 -8898
rect 5124 -9794 5184 -9696
rect 5584 -9792 5644 -9690
rect 4896 -9854 5184 -9794
rect 5578 -9852 5584 -9792
rect 5644 -9852 5650 -9792
rect 4896 -10100 4956 -9854
rect 5124 -10100 5184 -9854
rect 5814 -9918 5874 -7884
rect 6264 -8222 6270 -8162
rect 6330 -8222 6336 -8162
rect 6036 -8330 6042 -8270
rect 6102 -8330 6108 -8270
rect 6042 -8424 6102 -8330
rect 6270 -8494 6330 -8222
rect 6498 -8330 6504 -8270
rect 6564 -8330 6570 -8270
rect 6504 -8424 6564 -8330
rect 6044 -9228 6104 -8892
rect 6264 -9038 6270 -8978
rect 6330 -9038 6336 -8978
rect 6270 -9324 6330 -9038
rect 6504 -9228 6564 -8892
rect 6044 -9792 6104 -9698
rect 6504 -9792 6564 -9696
rect 6038 -9852 6044 -9792
rect 6104 -9852 6110 -9792
rect 6498 -9852 6504 -9792
rect 6564 -9852 6570 -9792
rect 6728 -9918 6788 -7884
rect 7422 -8268 7482 -7884
rect 7646 -8268 7706 -7884
rect 6954 -8330 6960 -8270
rect 7020 -8330 7026 -8270
rect 7422 -8328 7706 -8268
rect 6960 -8424 7020 -8330
rect 7422 -8416 7482 -8328
rect 6964 -9228 7024 -8892
rect 7186 -8978 7246 -8804
rect 7180 -9038 7186 -8978
rect 7246 -9038 7252 -8978
rect 7424 -9034 7484 -8892
rect 7646 -9034 7706 -8328
rect 7180 -9152 7186 -9092
rect 7246 -9152 7252 -9092
rect 7424 -9094 7706 -9034
rect 7186 -9314 7246 -9152
rect 7424 -9228 7484 -9094
rect 6958 -9792 7018 -9694
rect 7422 -9790 7482 -9698
rect 7646 -9790 7706 -9094
rect 6952 -9852 6958 -9792
rect 7018 -9852 7024 -9792
rect 7422 -9850 7706 -9790
rect 5808 -9978 5814 -9918
rect 5874 -9978 5880 -9918
rect 6722 -9978 6728 -9918
rect 6788 -9978 6794 -9918
rect 5814 -10100 5874 -9978
rect 6728 -10100 6788 -9978
rect 7422 -10100 7482 -9850
rect 7646 -10100 7706 -9850
rect 12516 -7982 12628 -7884
rect 4664 -10168 7854 -10100
rect -368 -10716 -256 -10570
rect 344 -10716 354 -10416
rect 4664 -10594 4734 -10168
rect 7798 -10594 7854 -10168
rect 4664 -10646 7854 -10594
rect 11906 -10716 11916 -10416
rect 12516 -10570 12522 -7982
rect 12622 -10570 12628 -7982
rect 12516 -10716 12628 -10570
rect -368 -10722 12628 -10716
rect -368 -10822 -262 -10722
rect 12522 -10822 12628 -10722
rect -368 -10828 12628 -10822
<< via1 >>
rect -256 2516 344 2816
rect 11916 2516 12516 2816
rect 158 2232 12268 2396
rect 172 2050 232 2110
rect 596 2050 656 2110
rect 1032 2050 1092 2110
rect 2746 2050 2806 2110
rect 4466 2050 4526 2110
rect 6174 2050 6234 2110
rect 7894 2050 7954 2110
rect 9608 2050 9668 2110
rect 11326 2050 11386 2110
rect 11754 2050 11814 2110
rect 12186 2050 12246 2110
rect -92 1786 -32 1846
rect 50 1658 110 1718
rect 1458 1922 1518 1982
rect 2312 1922 2372 1982
rect 3172 1922 3232 1982
rect 4032 1922 4092 1982
rect 4892 1922 4952 1982
rect 5752 1922 5812 1982
rect 6612 1922 6672 1982
rect 7472 1922 7532 1982
rect 8332 1922 8392 1982
rect 9172 1922 9232 1982
rect 8752 1658 8812 1718
rect 10030 1922 10090 1982
rect 10892 1922 10952 1982
rect 10468 1786 10528 1846
rect 50 -4 110 56
rect -92 -110 -32 -50
rect -92 -1640 -32 -1580
rect 1888 96 1948 156
rect 1890 -110 1950 -50
rect 50 -1846 110 -1786
rect 1458 -1744 1518 -1684
rect 2320 -1744 2380 -1684
rect 50 -3484 110 -3424
rect -92 -3590 -32 -3530
rect 1888 -3384 1948 -3324
rect 1890 -3590 1950 -3530
rect 1460 -5110 1520 -5050
rect 2320 -5110 2380 -5050
rect 1888 -5328 1948 -5268
rect 1456 -6986 1516 -6926
rect 2326 -6986 2386 -6926
rect 3470 -4 3530 56
rect 3604 -6 3664 54
rect 3182 -1744 3242 -1684
rect 4040 -1744 4100 -1684
rect 3470 -3484 3530 -3424
rect 3604 -3486 3664 -3426
rect 5320 -110 5380 -50
rect 7166 -110 7226 -50
rect 4900 -1744 4960 -1684
rect 5744 -1744 5804 -1684
rect 4462 -3592 4522 -3532
rect 3176 -5110 3236 -5050
rect 4042 -5110 4102 -5050
rect 3606 -5214 3666 -5154
rect 3184 -6986 3244 -6926
rect 4042 -6986 4102 -6926
rect 6614 -1744 6674 -1684
rect 7480 -1744 7540 -1684
rect 6180 -3256 6240 -3196
rect 5320 -3590 5380 -3530
rect 7166 -3590 7226 -3530
rect 8756 -6 8816 54
rect 8336 -1744 8396 -1684
rect 9192 -1744 9252 -1684
rect 8752 -1846 8812 -1786
rect 7894 -3590 7954 -3530
rect 4898 -5110 4958 -5050
rect 5746 -5110 5806 -5050
rect 5320 -6860 5380 -6800
rect 4900 -6986 4960 -6926
rect 5758 -6986 5818 -6926
rect 6600 -5110 6660 -5050
rect 7480 -5110 7540 -5050
rect 7038 -6860 7098 -6800
rect 6616 -6986 6676 -6926
rect 7474 -6986 7534 -6926
rect 8756 -3486 8816 -3426
rect 8334 -5110 8394 -5050
rect 9192 -5114 9252 -5054
rect 8752 -5214 8812 -5154
rect 8332 -6986 8392 -6926
rect 9190 -6986 9250 -6926
rect 10470 96 10530 156
rect 10468 -1640 10528 -1580
rect 10046 -1744 10106 -1684
rect 10904 -1744 10964 -1684
rect 10470 -3384 10530 -3324
rect 10048 -5110 10108 -5050
rect 10906 -5110 10966 -5050
rect 10470 -5328 10530 -5268
rect 10048 -6986 10108 -6926
rect 10904 -6986 10964 -6926
rect 170 -7130 230 -7070
rect 590 -7130 650 -7070
rect 1030 -7130 1090 -7070
rect 2748 -7130 2808 -7070
rect 4462 -7130 4522 -7070
rect 6180 -7130 6240 -7070
rect 7894 -7130 7954 -7070
rect 9608 -7130 9668 -7070
rect 11324 -7130 11384 -7070
rect 11750 -7130 11810 -7070
rect 12184 -7130 12244 -7070
rect 4798 -8222 4858 -8162
rect 5582 -8330 5642 -8270
rect 5356 -9038 5416 -8978
rect 4798 -9152 4858 -9092
rect 5356 -9152 5416 -9092
rect 5584 -9852 5644 -9792
rect 6270 -8222 6330 -8162
rect 6042 -8330 6102 -8270
rect 6504 -8330 6564 -8270
rect 6270 -9038 6330 -8978
rect 6044 -9852 6104 -9792
rect 6504 -9852 6564 -9792
rect 6960 -8330 7020 -8270
rect 7186 -9038 7246 -8978
rect 7186 -9152 7246 -9092
rect 6958 -9852 7018 -9792
rect 5814 -9978 5874 -9918
rect 6728 -9978 6788 -9918
rect -256 -10716 344 -10416
rect 4734 -10594 7798 -10168
rect 11916 -10716 12516 -10416
<< metal2 >>
rect -256 2816 344 2826
rect -256 2506 344 2516
rect 11916 2816 12516 2826
rect 11916 2506 12516 2516
rect 110 2396 12310 2438
rect 110 2232 158 2396
rect 12268 2232 12310 2396
rect 110 2192 12310 2232
rect 172 2110 232 2116
rect 596 2110 656 2116
rect 1032 2110 1092 2116
rect 2746 2110 2806 2116
rect 4466 2110 4526 2116
rect 6174 2110 6234 2116
rect 7894 2110 7954 2116
rect 9608 2110 9668 2116
rect 11326 2110 11386 2116
rect 11754 2110 11814 2116
rect 12186 2110 12246 2116
rect 232 2050 596 2110
rect 656 2050 1032 2110
rect 1092 2050 2746 2110
rect 2806 2050 4466 2110
rect 4526 2050 6174 2110
rect 6234 2050 7894 2110
rect 7954 2050 9608 2110
rect 9668 2050 11326 2110
rect 11386 2050 11754 2110
rect 11814 2050 12186 2110
rect 172 2044 232 2050
rect 596 2044 656 2050
rect 1032 2044 1092 2050
rect 2746 2044 2806 2050
rect 4466 2044 4526 2050
rect 6174 2044 6234 2050
rect 7894 2044 7954 2050
rect 9608 2044 9668 2050
rect 11326 2044 11386 2050
rect 11754 2044 11814 2050
rect 12186 2044 12246 2050
rect 1458 1982 1518 1988
rect 2312 1982 2372 1988
rect 3172 1982 3232 1988
rect 4032 1982 4092 1988
rect 4892 1982 4952 1988
rect 5752 1982 5812 1988
rect 6612 1982 6672 1988
rect 7472 1982 7532 1988
rect 8332 1982 8392 1988
rect 9172 1982 9232 1988
rect 10030 1982 10090 1988
rect 10892 1982 10952 1988
rect 1518 1922 2312 1982
rect 2372 1922 3172 1982
rect 3232 1922 4032 1982
rect 4092 1922 4892 1982
rect 4952 1922 5752 1982
rect 5812 1922 6612 1982
rect 6672 1922 7472 1982
rect 7532 1922 8332 1982
rect 8392 1922 9172 1982
rect 9232 1922 10030 1982
rect 10090 1922 10892 1982
rect 1458 1916 1518 1922
rect 2312 1916 2372 1922
rect 3172 1916 3232 1922
rect 4032 1916 4092 1922
rect 4892 1916 4952 1922
rect 5752 1916 5812 1922
rect 6612 1916 6672 1922
rect 7472 1916 7532 1922
rect 8332 1916 8392 1922
rect 9172 1916 9232 1922
rect 10030 1916 10090 1922
rect 10892 1916 10952 1922
rect -92 1846 -32 1852
rect 10468 1846 10528 1852
rect -32 1786 10468 1846
rect -92 1780 -32 1786
rect 10468 1780 10528 1786
rect 50 1718 110 1724
rect 8752 1718 8812 1724
rect 110 1658 8752 1718
rect 50 1652 110 1658
rect 8752 1652 8812 1658
rect 1888 156 1948 162
rect 10470 156 10530 162
rect 1948 96 10470 156
rect 1888 90 1948 96
rect 10470 90 10530 96
rect 50 56 110 62
rect 3470 56 3530 62
rect 110 -4 3470 56
rect 50 -10 110 -4
rect 3470 -10 3530 -4
rect 3604 54 3664 60
rect 8756 54 8816 60
rect 3664 -6 8756 54
rect 3604 -12 3664 -6
rect 8756 -12 8816 -6
rect -92 -50 -32 -44
rect 1890 -50 1950 -44
rect -32 -110 1890 -50
rect -92 -116 -32 -110
rect 1890 -116 1950 -110
rect 5320 -50 5380 -44
rect 7166 -50 7226 -44
rect 5380 -110 7166 -50
rect 5320 -116 5380 -110
rect 7166 -116 7226 -110
rect -92 -1580 -32 -1574
rect 10468 -1580 10528 -1574
rect -32 -1640 10468 -1580
rect -92 -1646 -32 -1640
rect 10468 -1646 10528 -1640
rect 10904 -1684 10964 -1678
rect 1452 -1744 1458 -1684
rect 1518 -1744 2320 -1684
rect 2380 -1744 3182 -1684
rect 3242 -1744 4040 -1684
rect 4100 -1744 4900 -1684
rect 4960 -1744 5744 -1684
rect 5804 -1744 6614 -1684
rect 6674 -1744 7480 -1684
rect 7540 -1744 8336 -1684
rect 8396 -1744 9192 -1684
rect 9252 -1744 10046 -1684
rect 10106 -1744 10904 -1684
rect 10904 -1750 10964 -1744
rect 50 -1786 110 -1780
rect 8752 -1786 8812 -1780
rect 110 -1846 8752 -1786
rect 50 -1852 110 -1846
rect 8752 -1852 8812 -1846
rect 6180 -3196 6240 -3187
rect 6174 -3256 6180 -3196
rect 6240 -3256 6246 -3196
rect 6180 -3265 6240 -3256
rect 1888 -3324 1948 -3318
rect 10470 -3324 10530 -3318
rect 1948 -3384 10470 -3324
rect 1888 -3390 1948 -3384
rect 10470 -3390 10530 -3384
rect 50 -3424 110 -3418
rect 3470 -3424 3530 -3418
rect 110 -3484 3470 -3424
rect 50 -3490 110 -3484
rect 3470 -3490 3530 -3484
rect 3604 -3426 3664 -3420
rect 8756 -3426 8816 -3420
rect 3664 -3486 8756 -3426
rect 3604 -3492 3664 -3486
rect 8756 -3492 8816 -3486
rect -92 -3530 -32 -3524
rect 1890 -3530 1950 -3524
rect -32 -3590 1890 -3530
rect 4462 -3532 4522 -3523
rect 5320 -3530 5380 -3524
rect 7166 -3530 7226 -3524
rect 7894 -3530 7954 -3521
rect -92 -3596 -32 -3590
rect 1890 -3596 1950 -3590
rect 4456 -3592 4462 -3532
rect 4522 -3592 4528 -3532
rect 5380 -3590 7166 -3530
rect 7888 -3590 7894 -3530
rect 7954 -3590 7960 -3530
rect 4462 -3601 4522 -3592
rect 5320 -3596 5380 -3590
rect 7166 -3596 7226 -3590
rect 7894 -3599 7954 -3590
rect 1460 -5050 1520 -5044
rect 1520 -5110 2320 -5050
rect 2380 -5110 3176 -5050
rect 3236 -5110 4042 -5050
rect 4102 -5110 4898 -5050
rect 4958 -5110 5746 -5050
rect 5806 -5110 6600 -5050
rect 6660 -5110 7480 -5050
rect 7540 -5110 8334 -5050
rect 8394 -5054 10048 -5050
rect 8394 -5110 9192 -5054
rect 1460 -5116 1520 -5110
rect 9186 -5114 9192 -5110
rect 9252 -5110 10048 -5054
rect 10108 -5110 10906 -5050
rect 10966 -5110 10972 -5050
rect 9252 -5114 9258 -5110
rect 3606 -5154 3666 -5148
rect 8752 -5154 8812 -5148
rect 3666 -5214 8752 -5154
rect 3606 -5220 3666 -5214
rect 8752 -5220 8812 -5214
rect 1888 -5268 1948 -5262
rect 10470 -5268 10530 -5262
rect 1948 -5328 10470 -5268
rect 1888 -5334 1948 -5328
rect 10470 -5334 10530 -5328
rect 5320 -6800 5380 -6794
rect 7038 -6800 7098 -6794
rect 5380 -6860 7038 -6800
rect 5320 -6866 5380 -6860
rect 7038 -6866 7098 -6860
rect 1456 -6926 1516 -6920
rect 2326 -6926 2386 -6920
rect 3184 -6926 3244 -6920
rect 4042 -6926 4102 -6920
rect 4900 -6926 4960 -6920
rect 5758 -6926 5818 -6920
rect 6616 -6926 6676 -6920
rect 7474 -6926 7534 -6920
rect 8332 -6926 8392 -6920
rect 9190 -6926 9250 -6920
rect 10048 -6926 10108 -6920
rect 10904 -6926 10964 -6920
rect 1516 -6986 2326 -6926
rect 2386 -6986 3184 -6926
rect 3244 -6986 4042 -6926
rect 4102 -6986 4900 -6926
rect 4960 -6986 5758 -6926
rect 5818 -6986 6616 -6926
rect 6676 -6986 7474 -6926
rect 7534 -6986 8332 -6926
rect 8392 -6986 9190 -6926
rect 9250 -6986 10048 -6926
rect 10108 -6986 10904 -6926
rect 1456 -6992 1516 -6986
rect 2326 -6992 2386 -6986
rect 3184 -6992 3244 -6986
rect 4042 -6992 4102 -6986
rect 4900 -6992 4960 -6986
rect 5758 -6992 5818 -6986
rect 6616 -6992 6676 -6986
rect 7474 -6992 7534 -6986
rect 8332 -6992 8392 -6986
rect 9190 -6992 9250 -6986
rect 10048 -6992 10108 -6986
rect 10904 -6992 10964 -6986
rect 170 -7070 230 -7064
rect 590 -7070 650 -7064
rect 1030 -7070 1090 -7064
rect 2748 -7070 2808 -7064
rect 4462 -7070 4522 -7064
rect 6180 -7070 6240 -7064
rect 7894 -7070 7954 -7064
rect 9608 -7070 9668 -7064
rect 11324 -7070 11384 -7064
rect 11750 -7070 11810 -7064
rect 12184 -7070 12244 -7064
rect 230 -7130 590 -7070
rect 650 -7130 1030 -7070
rect 1090 -7130 2748 -7070
rect 2808 -7130 4462 -7070
rect 4522 -7130 6180 -7070
rect 6240 -7130 7894 -7070
rect 7954 -7130 9608 -7070
rect 9668 -7130 11324 -7070
rect 11384 -7130 11750 -7070
rect 11810 -7130 12184 -7070
rect 170 -7136 230 -7130
rect 590 -7136 650 -7130
rect 1030 -7136 1090 -7130
rect 2748 -7136 2808 -7130
rect 4462 -7136 4522 -7130
rect 6180 -7136 6240 -7130
rect 7894 -7136 7954 -7130
rect 9608 -7136 9668 -7130
rect 11324 -7136 11384 -7130
rect 11750 -7136 11810 -7130
rect 12184 -7136 12244 -7130
rect 4798 -8162 4858 -8156
rect 6270 -8162 6330 -8156
rect 4858 -8222 6270 -8162
rect 4798 -8228 4858 -8222
rect 6270 -8228 6330 -8222
rect 5582 -8270 5642 -8264
rect 6042 -8270 6102 -8264
rect 6504 -8270 6564 -8264
rect 6960 -8270 7020 -8264
rect 5642 -8330 6042 -8270
rect 6102 -8330 6504 -8270
rect 6564 -8330 6960 -8270
rect 5582 -8336 5642 -8330
rect 6042 -8336 6102 -8330
rect 6504 -8336 6564 -8330
rect 6960 -8336 7020 -8330
rect 5356 -8978 5416 -8972
rect 6270 -8978 6330 -8972
rect 7186 -8978 7246 -8972
rect 5416 -9038 6270 -8978
rect 6330 -9038 7186 -8978
rect 5356 -9044 5416 -9038
rect 6270 -9044 6330 -9038
rect 7186 -9044 7246 -9038
rect 4798 -9092 4858 -9086
rect 5356 -9092 5416 -9086
rect 7186 -9092 7246 -9086
rect 4858 -9152 5356 -9092
rect 5416 -9152 7186 -9092
rect 4798 -9158 4858 -9152
rect 5356 -9158 5416 -9152
rect 7186 -9158 7246 -9152
rect 5584 -9792 5644 -9786
rect 6044 -9792 6104 -9786
rect 6504 -9792 6564 -9786
rect 6958 -9792 7018 -9786
rect 5644 -9852 6044 -9792
rect 6104 -9852 6504 -9792
rect 6564 -9852 6958 -9792
rect 5584 -9858 5644 -9852
rect 6044 -9858 6104 -9852
rect 6504 -9858 6564 -9852
rect 6958 -9858 7018 -9852
rect 5814 -9918 5874 -9912
rect 6728 -9918 6788 -9912
rect 5874 -9978 6728 -9918
rect 5814 -9984 5874 -9978
rect 6728 -9984 6788 -9978
rect 4664 -10168 7854 -10100
rect -256 -10416 344 -10406
rect 4664 -10594 4734 -10168
rect 7798 -10594 7854 -10168
rect 4664 -10646 7854 -10594
rect 11916 -10416 12516 -10406
rect -256 -10726 344 -10716
rect 11916 -10726 12516 -10716
<< via2 >>
rect -256 2516 344 2816
rect 11916 2516 12516 2816
rect 158 2232 12268 2396
rect 6180 -3256 6240 -3196
rect 4462 -3592 4522 -3532
rect 7894 -3590 7954 -3530
rect -256 -10716 344 -10416
rect 4734 -10594 7798 -10168
rect 11916 -10716 12516 -10416
<< metal3 >>
rect -266 2816 354 2821
rect -266 2516 -256 2816
rect 344 2516 354 2816
rect -266 2511 354 2516
rect 11906 2816 12526 2821
rect 11906 2516 11916 2816
rect 12516 2516 12526 2816
rect 11906 2511 12526 2516
rect 110 2396 12310 2438
rect 110 2232 158 2396
rect 12268 2232 12310 2396
rect 110 2192 12310 2232
rect 6158 -3196 6258 -3176
rect 6158 -3256 6180 -3196
rect 6240 -3256 6258 -3196
rect 6158 -3512 6258 -3256
rect 4434 -3530 7988 -3512
rect 4434 -3532 7894 -3530
rect 4434 -3592 4462 -3532
rect 4522 -3590 7894 -3532
rect 7954 -3590 7988 -3530
rect 4522 -3592 7988 -3590
rect 4434 -3612 7988 -3592
rect 4664 -10168 7854 -10100
rect -266 -10416 354 -10411
rect -266 -10716 -256 -10416
rect 344 -10716 354 -10416
rect 4664 -10594 4734 -10168
rect 7798 -10594 7854 -10168
rect 4664 -10646 7854 -10594
rect 11906 -10416 12526 -10411
rect -266 -10721 354 -10716
rect 11906 -10716 11916 -10416
rect 12516 -10716 12526 -10416
rect 11906 -10721 12526 -10716
<< via3 >>
rect -256 2516 344 2816
rect 11916 2516 12516 2816
rect 158 2232 12268 2396
rect -256 -10716 344 -10416
rect 4734 -10594 7798 -10168
rect 11916 -10716 12516 -10416
<< metal4 >>
rect -440 2816 12700 3000
rect -440 2516 -256 2816
rect 344 2516 11916 2816
rect 12516 2516 12700 2816
rect -440 2396 12700 2516
rect -440 2232 158 2396
rect 12268 2232 12700 2396
rect -440 2200 12700 2232
rect -440 -10168 12700 -10100
rect -440 -10416 4734 -10168
rect -440 -10716 -256 -10416
rect 344 -10594 4734 -10416
rect 7798 -10416 12700 -10168
rect 7798 -10594 11916 -10416
rect 344 -10716 11916 -10594
rect 12516 -10716 12700 -10416
rect -440 -10900 12700 -10716
use sky130_fd_pr__nfet_01v8_C5Q2Z6  sky130_fd_pr__nfet_01v8_C5Q2Z6_0
timestamp 1624477805
transform 1 0 6301 0 1 -8660
box -1403 -288 1403 288
use sky130_fd_pr__nfet_01v8_C5Q2Z6  sky130_fd_pr__nfet_01v8_C5Q2Z6_1
timestamp 1624477805
transform 1 0 6301 0 1 -9460
box -1403 -288 1403 288
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_4
timestamp 1624477805
transform 1 0 6209 0 1 -6056
box -6071 -700 6071 700
use ntap  ntap_66 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/ntap
timestamp 1624477805
transform 1 0 266 0 1 -5512
box 250 218 480 436
use ntap  ntap_67
timestamp 1624477805
transform 1 0 1124 0 1 -5512
box 250 218 480 436
use ntap  ntap_69
timestamp 1624477805
transform 1 0 1982 0 1 -5512
box 250 218 480 436
use ntap  ntap_68
timestamp 1624477805
transform 1 0 2840 0 1 -5512
box 250 218 480 436
use ntap  ntap_56
timestamp 1624477805
transform 1 0 3698 0 1 -5512
box 250 218 480 436
use ntap  ntap_57
timestamp 1624477805
transform 1 0 4556 0 1 -5512
box 250 218 480 436
use ntap  ntap_58
timestamp 1624477805
transform 1 0 5414 0 1 -5512
box 250 218 480 436
use ntap  ntap_59
timestamp 1624477805
transform 1 0 6272 0 1 -5512
box 250 218 480 436
use ntap  ntap_60
timestamp 1624477805
transform 1 0 7130 0 1 -5512
box 250 218 480 436
use ntap  ntap_61
timestamp 1624477805
transform 1 0 7988 0 1 -5512
box 250 218 480 436
use ntap  ntap_62
timestamp 1624477805
transform 1 0 8846 0 1 -5512
box 250 218 480 436
use ntap  ntap_63
timestamp 1624477805
transform 1 0 9704 0 1 -5512
box 250 218 480 436
use ntap  ntap_64
timestamp 1624477805
transform 1 0 10562 0 1 -5512
box 250 218 480 436
use ntap  ntap_65
timestamp 1624477805
transform 1 0 11420 0 1 -5512
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_3
timestamp 1624477805
transform 1 0 6209 0 1 -4316
box -6071 -700 6071 700
use ntap  ntap_52
timestamp 1624477805
transform 1 0 278 0 1 -3768
box 250 218 480 436
use ntap  ntap_53
timestamp 1624477805
transform 1 0 1136 0 1 -3768
box 250 218 480 436
use ntap  ntap_55
timestamp 1624477805
transform 1 0 1994 0 1 -3768
box 250 218 480 436
use ntap  ntap_54
timestamp 1624477805
transform 1 0 2852 0 1 -3768
box 250 218 480 436
use ntap  ntap_42
timestamp 1624477805
transform 1 0 3710 0 1 -3768
box 250 218 480 436
use ntap  ntap_43
timestamp 1624477805
transform 1 0 4568 0 1 -3768
box 250 218 480 436
use ntap  ntap_44
timestamp 1624477805
transform 1 0 5426 0 1 -3768
box 250 218 480 436
use ntap  ntap_45
timestamp 1624477805
transform 1 0 6284 0 1 -3768
box 250 218 480 436
use ntap  ntap_46
timestamp 1624477805
transform 1 0 7142 0 1 -3768
box 250 218 480 436
use ntap  ntap_47
timestamp 1624477805
transform 1 0 8000 0 1 -3768
box 250 218 480 436
use ntap  ntap_48
timestamp 1624477805
transform 1 0 8858 0 1 -3768
box 250 218 480 436
use ntap  ntap_49
timestamp 1624477805
transform 1 0 9716 0 1 -3768
box 250 218 480 436
use ntap  ntap_50
timestamp 1624477805
transform 1 0 10574 0 1 -3768
box 250 218 480 436
use ntap  ntap_51
timestamp 1624477805
transform 1 0 11432 0 1 -3768
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_2
timestamp 1624477805
transform 1 0 6209 0 1 -2576
box -6071 -700 6071 700
use ntap  ntap_38
timestamp 1624477805
transform 1 0 278 0 1 -2032
box 250 218 480 436
use ntap  ntap_39
timestamp 1624477805
transform 1 0 1136 0 1 -2032
box 250 218 480 436
use ntap  ntap_41
timestamp 1624477805
transform 1 0 1994 0 1 -2032
box 250 218 480 436
use ntap  ntap_40
timestamp 1624477805
transform 1 0 2852 0 1 -2032
box 250 218 480 436
use ntap  ntap_28
timestamp 1624477805
transform 1 0 3710 0 1 -2032
box 250 218 480 436
use ntap  ntap_29
timestamp 1624477805
transform 1 0 4568 0 1 -2032
box 250 218 480 436
use ntap  ntap_30
timestamp 1624477805
transform 1 0 5426 0 1 -2032
box 250 218 480 436
use ntap  ntap_31
timestamp 1624477805
transform 1 0 6284 0 1 -2032
box 250 218 480 436
use ntap  ntap_32
timestamp 1624477805
transform 1 0 7142 0 1 -2032
box 250 218 480 436
use ntap  ntap_33
timestamp 1624477805
transform 1 0 8000 0 1 -2032
box 250 218 480 436
use ntap  ntap_34
timestamp 1624477805
transform 1 0 8858 0 1 -2032
box 250 218 480 436
use ntap  ntap_35
timestamp 1624477805
transform 1 0 9716 0 1 -2032
box 250 218 480 436
use ntap  ntap_36
timestamp 1624477805
transform 1 0 10574 0 1 -2032
box 250 218 480 436
use ntap  ntap_37
timestamp 1624477805
transform 1 0 11432 0 1 -2032
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_1
timestamp 1624477805
transform 1 0 6209 0 1 -836
box -6071 -700 6071 700
use ntap  ntap_24
timestamp 1624477805
transform 1 0 282 0 1 -290
box 250 218 480 436
use ntap  ntap_25
timestamp 1624477805
transform 1 0 1140 0 1 -290
box 250 218 480 436
use ntap  ntap_27
timestamp 1624477805
transform 1 0 1998 0 1 -290
box 250 218 480 436
use ntap  ntap_26
timestamp 1624477805
transform 1 0 2856 0 1 -290
box 250 218 480 436
use ntap  ntap_14
timestamp 1624477805
transform 1 0 3714 0 1 -290
box 250 218 480 436
use ntap  ntap_15
timestamp 1624477805
transform 1 0 4572 0 1 -290
box 250 218 480 436
use ntap  ntap_16
timestamp 1624477805
transform 1 0 5430 0 1 -290
box 250 218 480 436
use ntap  ntap_17
timestamp 1624477805
transform 1 0 6288 0 1 -290
box 250 218 480 436
use ntap  ntap_18
timestamp 1624477805
transform 1 0 7146 0 1 -290
box 250 218 480 436
use ntap  ntap_19
timestamp 1624477805
transform 1 0 8004 0 1 -290
box 250 218 480 436
use ntap  ntap_20
timestamp 1624477805
transform 1 0 8862 0 1 -290
box 250 218 480 436
use ntap  ntap_21
timestamp 1624477805
transform 1 0 9720 0 1 -290
box 250 218 480 436
use ntap  ntap_22
timestamp 1624477805
transform 1 0 10578 0 1 -290
box 250 218 480 436
use ntap  ntap_23
timestamp 1624477805
transform 1 0 11436 0 1 -290
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_0
timestamp 1624477805
transform 1 0 6209 0 1 904
box -6071 -700 6071 700
use ntap  ntap_0
timestamp 1624477805
transform 1 0 266 0 1 1474
box 250 218 480 436
use ntap  ntap_1
timestamp 1624477805
transform 1 0 1124 0 1 1474
box 250 218 480 436
use ntap  ntap_2
timestamp 1624477805
transform 1 0 1982 0 1 1474
box 250 218 480 436
use ntap  ntap_3
timestamp 1624477805
transform 1 0 2840 0 1 1474
box 250 218 480 436
use ntap  ntap_4
timestamp 1624477805
transform 1 0 3698 0 1 1474
box 250 218 480 436
use ntap  ntap_5
timestamp 1624477805
transform 1 0 4556 0 1 1474
box 250 218 480 436
use ntap  ntap_6
timestamp 1624477805
transform 1 0 5414 0 1 1474
box 250 218 480 436
use ntap  ntap_7
timestamp 1624477805
transform 1 0 6272 0 1 1474
box 250 218 480 436
use ntap  ntap_8
timestamp 1624477805
transform 1 0 7130 0 1 1474
box 250 218 480 436
use ntap  ntap_9
timestamp 1624477805
transform 1 0 7988 0 1 1474
box 250 218 480 436
use ntap  ntap_10
timestamp 1624477805
transform 1 0 8846 0 1 1474
box 250 218 480 436
use ntap  ntap_11
timestamp 1624477805
transform 1 0 9704 0 1 1474
box 250 218 480 436
use ntap  ntap_12
timestamp 1624477805
transform 1 0 10562 0 1 1474
box 250 218 480 436
use ntap  ntap_13
timestamp 1624477805
transform 1 0 11420 0 1 1474
box 250 218 480 436
<< labels >>
flabel metal2 2170 120 2190 138 1 FreeSans 480 0 0 0 low_freq_pll_ibiasn
flabel metal2 1436 -74 1454 -64 1 FreeSans 480 0 0 0 comparator_ibiasn
flabel metal2 3796 12 3814 26 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn4
flabel metal1 5340 180 5354 186 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn3
flabel metal2 5890 -90 5904 -74 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn2
flabel metal2 2212 16 2228 34 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn1
flabel metal2 1210 -3580 1234 -3554 1 FreeSans 480 0 0 0 sample_and_hold_ibiasn_A
flabel metal2 1524 -3460 1542 -3444 1 FreeSans 480 0 0 0 peak_detector_ibiasn2
flabel metal2 6342 -3576 6354 -3558 1 FreeSans 480 0 0 0 peak_detector_ibiasn1
flabel metal1 5342 -3304 5356 -3294 1 FreeSans 480 0 0 0 diff_to_se_converter_ibiasn
flabel metal2 3948 -3460 3954 -3444 1 FreeSans 480 0 0 0 input_amplifier_ibiasn2
flabel metal2 3240 -3356 3256 -3342 1 FreeSans 480 0 0 0 input_amplifier_ibiasn1
flabel metal2 6058 -6832 6082 -6816 1 FreeSans 480 0 0 0 dac_8bit_ibiasn_B
flabel metal2 4048 -5194 4060 -5174 1 FreeSans 480 0 0 0 sample_and_hold_ibiasn_B
flabel metal2 2324 -5298 2344 -5282 1 FreeSans 480 0 0 0 dac_8bit_ibiasn_A
flabel metal2 3562 -6966 3574 -6948 1 FreeSans 480 0 0 0 vbiasp
flabel metal4 -414 2968 -398 2984 1 FreeSans 480 0 0 0 VDD
flabel metal2 6620 -9826 6626 -9814 1 FreeSans 480 0 0 0 vbiasn
flabel metal2 5934 -9020 5950 -9006 1 FreeSans 480 0 0 0 dac_8bit_ibiasp_A
flabel metal2 5264 -9132 5274 -9118 1 FreeSans 480 0 0 0 dac_8bit_ibiasp_B
flabel metal4 -398 -10890 -382 -10872 1 FreeSans 480 0 0 0 VSS
<< properties >>
string FIXED_BBOX -312 -11172 12572 -8028
<< end >>
