magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_s >>
rect 79 421 91 424
rect 38 420 91 421
rect 101 420 113 424
rect 151 420 163 424
rect 173 420 185 424
rect 38 412 80 420
rect 38 395 113 412
rect 114 400 125 412
rect 139 400 150 412
rect 30 383 38 395
rect 42 378 76 395
rect 79 378 113 395
rect -25 262 25 264
rect -8 253 17 261
rect 25 253 27 262
rect -12 246 38 253
rect 71 251 80 279
rect -12 245 34 246
rect -12 241 8 245
rect 0 229 8 241
rect 17 229 34 245
rect 0 228 34 229
rect 0 221 38 228
rect 25 212 27 221
rect 69 213 80 251
rect 144 241 148 395
rect 151 378 156 412
rect 180 378 185 412
rect 186 400 197 412
rect 400 395 442 421
rect 806 395 848 421
rect 1063 420 1075 424
rect 1085 420 1097 424
rect 1135 420 1147 424
rect 1157 421 1169 424
rect 1327 421 1339 424
rect 1157 420 1210 421
rect 1168 412 1210 420
rect 1051 400 1062 412
rect 332 341 336 395
rect 392 387 438 395
rect 392 383 408 387
rect 400 380 408 383
rect 434 380 438 387
rect 442 383 450 395
rect 798 383 806 395
rect 810 387 844 395
rect 810 380 814 387
rect 840 380 844 387
rect 848 383 856 395
rect 388 379 454 380
rect 794 379 860 380
rect 400 371 404 379
rect 454 365 504 367
rect 744 365 794 367
rect 494 361 548 365
rect 700 361 754 365
rect 494 356 514 361
rect 734 356 754 361
rect 504 341 506 356
rect 332 261 336 329
rect 400 305 404 341
rect 498 331 506 341
rect 514 331 515 351
rect 504 315 506 331
rect 525 322 528 356
rect 547 331 548 351
rect 557 331 564 341
rect 684 331 691 341
rect 700 331 701 351
rect 720 322 723 356
rect 733 331 734 351
rect 743 331 750 341
rect 514 315 530 321
rect 532 315 548 321
rect 700 315 716 321
rect 718 315 734 321
rect 794 315 796 365
rect 337 267 373 295
rect 337 261 351 267
rect 107 207 119 241
rect 129 207 149 241
rect 42 94 76 98
rect 42 79 46 94
rect 72 79 76 94
rect 38 61 80 79
rect 16 55 102 61
rect 144 55 148 207
rect 174 183 181 211
rect 332 183 336 251
rect 341 233 351 261
rect 361 261 375 267
rect 400 261 411 305
rect 837 267 848 305
rect 875 267 911 295
rect 912 267 916 395
rect 1063 378 1068 412
rect 1092 378 1097 412
rect 1098 400 1109 412
rect 1123 400 1134 412
rect 1135 395 1210 412
rect 1286 420 1339 421
rect 1349 420 1361 424
rect 1399 420 1411 424
rect 1421 420 1433 424
rect 1286 412 1328 420
rect 1286 395 1361 412
rect 1362 400 1373 412
rect 1387 400 1398 412
rect 1100 341 1104 395
rect 1135 378 1206 395
rect 1210 383 1218 395
rect 1278 383 1286 395
rect 1290 378 1324 395
rect 1327 378 1361 395
rect 1168 371 1172 378
rect 562 262 612 264
rect 636 262 686 264
rect 361 233 381 261
rect 400 233 409 261
rect 463 253 497 261
rect 442 246 497 253
rect 463 245 497 246
rect 565 253 596 261
rect 565 245 599 253
rect 400 213 404 233
rect 596 229 599 245
rect 463 228 497 229
rect 442 221 497 228
rect 565 221 599 229
rect 612 212 614 262
rect 652 253 683 261
rect 686 253 688 262
rect 875 261 887 267
rect 652 245 688 253
rect 751 253 785 261
rect 751 246 806 253
rect 751 245 785 246
rect 683 229 688 245
rect 877 233 887 261
rect 897 233 917 267
rect 1100 261 1104 329
rect 1168 291 1172 341
rect 1168 251 1177 279
rect 1264 264 1274 291
rect 1223 262 1274 264
rect 1264 261 1275 262
rect 1231 253 1265 261
rect 1273 253 1275 261
rect 652 221 688 229
rect 751 228 785 229
rect 751 221 806 228
rect 686 212 688 221
rect 332 103 336 171
rect 400 133 404 183
rect 454 159 504 161
rect 744 159 794 161
rect 504 143 506 159
rect 514 153 530 159
rect 532 153 548 159
rect 700 153 716 159
rect 718 153 734 159
rect 525 143 548 152
rect 700 143 723 152
rect 498 133 506 143
rect 504 109 506 133
rect 514 123 515 143
rect 525 118 528 143
rect 547 123 548 143
rect 557 133 564 143
rect 684 133 691 143
rect 700 123 701 143
rect 720 118 723 143
rect 733 123 734 143
rect 743 133 750 143
rect 514 109 548 113
rect 700 109 734 113
rect 794 109 796 159
rect 400 103 442 104
rect 806 103 848 104
rect 400 96 404 103
rect 295 62 300 96
rect 324 62 329 96
rect 367 79 438 96
rect 810 79 844 96
rect 847 79 881 96
rect 367 62 442 79
rect 400 61 442 62
rect 806 62 881 79
rect 806 61 848 62
rect 378 55 464 61
rect 784 55 870 61
rect 912 55 916 233
rect 1100 183 1104 251
rect 1109 207 1119 241
rect 1129 213 1149 241
rect 1129 207 1143 213
rect 1168 207 1179 251
rect 1210 246 1286 253
rect 1319 251 1328 279
rect 1231 228 1265 246
rect 1273 228 1275 246
rect 1210 221 1286 228
rect 1273 213 1275 221
rect 1317 213 1328 251
rect 1392 241 1396 395
rect 1399 378 1404 412
rect 1428 378 1433 412
rect 1434 400 1445 412
rect 1648 395 1690 421
rect 2054 395 2096 421
rect 2311 420 2323 424
rect 2333 420 2345 424
rect 2383 420 2395 424
rect 2405 421 2417 424
rect 2575 421 2587 424
rect 2405 420 2458 421
rect 2416 412 2458 420
rect 2299 400 2310 412
rect 1580 341 1584 395
rect 1640 387 1686 395
rect 1640 383 1656 387
rect 1648 380 1656 383
rect 1682 380 1686 387
rect 1690 383 1698 395
rect 2046 383 2054 395
rect 2058 387 2092 395
rect 2058 380 2062 387
rect 2088 380 2092 387
rect 2096 383 2104 395
rect 1636 379 1702 380
rect 2042 379 2108 380
rect 1648 371 1652 379
rect 1702 365 1752 367
rect 1992 365 2042 367
rect 1742 361 1796 365
rect 1948 361 2002 365
rect 1742 356 1762 361
rect 1982 356 2002 361
rect 1752 341 1754 356
rect 1580 261 1584 329
rect 1648 305 1652 341
rect 1746 331 1754 341
rect 1762 331 1763 351
rect 1752 315 1754 331
rect 1773 322 1776 356
rect 1795 331 1796 351
rect 1805 331 1812 341
rect 1932 331 1939 341
rect 1948 331 1949 351
rect 1968 322 1971 356
rect 1981 331 1982 351
rect 1991 331 1998 341
rect 1762 315 1778 321
rect 1780 315 1796 321
rect 1948 315 1964 321
rect 1966 315 1982 321
rect 2042 315 2044 365
rect 1585 267 1621 295
rect 1585 261 1599 267
rect 1264 212 1275 213
rect 1109 183 1116 207
rect 1264 183 1274 212
rect 1355 207 1367 241
rect 1377 207 1397 241
rect 1100 103 1104 171
rect 1168 133 1172 183
rect 1168 98 1172 103
rect 919 62 924 96
rect 948 62 953 96
rect 1168 94 1206 98
rect 1168 79 1176 94
rect 1202 79 1206 94
rect 1290 94 1324 98
rect 1290 79 1294 94
rect 1320 79 1324 94
rect 1168 61 1210 79
rect 1286 61 1328 79
rect 1146 55 1232 61
rect 1264 55 1350 61
rect 1392 55 1396 207
rect 1422 183 1429 211
rect 1580 183 1584 251
rect 1589 233 1599 261
rect 1609 261 1623 267
rect 1648 261 1659 305
rect 2085 267 2096 305
rect 2123 267 2159 295
rect 2160 267 2164 395
rect 2311 378 2316 412
rect 2340 378 2345 412
rect 2346 400 2357 412
rect 2371 400 2382 412
rect 2383 395 2458 412
rect 2534 420 2587 421
rect 2597 420 2609 424
rect 2647 420 2659 424
rect 2669 420 2681 424
rect 2534 412 2576 420
rect 2534 395 2609 412
rect 2610 400 2621 412
rect 2635 400 2646 412
rect 2348 341 2352 395
rect 2383 378 2454 395
rect 2458 383 2466 395
rect 2526 383 2534 395
rect 2538 378 2572 395
rect 2575 378 2609 395
rect 2416 371 2420 378
rect 1810 262 1860 264
rect 1884 262 1934 264
rect 1609 233 1629 261
rect 1648 233 1657 261
rect 1711 253 1745 261
rect 1690 246 1745 253
rect 1711 245 1745 246
rect 1813 253 1844 261
rect 1813 245 1847 253
rect 1648 213 1652 233
rect 1844 229 1847 245
rect 1711 228 1745 229
rect 1690 221 1745 228
rect 1813 221 1847 229
rect 1860 212 1862 262
rect 1900 253 1931 261
rect 1934 253 1936 262
rect 2123 261 2135 267
rect 1900 245 1936 253
rect 1999 253 2033 261
rect 1999 246 2054 253
rect 1999 245 2033 246
rect 1931 229 1936 245
rect 2125 233 2135 261
rect 2145 233 2165 267
rect 2348 261 2352 329
rect 2416 291 2420 341
rect 2416 251 2425 279
rect 2512 264 2522 291
rect 2471 262 2522 264
rect 2512 261 2523 262
rect 2479 253 2513 261
rect 2521 253 2523 261
rect 1900 221 1936 229
rect 1999 228 2033 229
rect 1999 221 2054 228
rect 1934 212 1936 221
rect 1580 103 1584 171
rect 1648 133 1652 183
rect 1702 159 1752 161
rect 1992 159 2042 161
rect 1752 143 1754 159
rect 1762 153 1778 159
rect 1780 153 1796 159
rect 1948 153 1964 159
rect 1966 153 1982 159
rect 1773 143 1796 152
rect 1948 143 1971 152
rect 1746 133 1754 143
rect 1752 109 1754 133
rect 1762 123 1763 143
rect 1773 118 1776 143
rect 1795 123 1796 143
rect 1805 133 1812 143
rect 1932 133 1939 143
rect 1948 123 1949 143
rect 1968 118 1971 143
rect 1981 123 1982 143
rect 1991 133 1998 143
rect 1762 109 1796 113
rect 1948 109 1982 113
rect 2042 109 2044 159
rect 1648 103 1690 104
rect 2054 103 2096 104
rect 1648 96 1652 103
rect 1543 62 1548 96
rect 1572 62 1577 96
rect 1615 79 1686 96
rect 2058 79 2092 96
rect 2095 79 2129 96
rect 1615 62 1690 79
rect 1648 61 1690 62
rect 2054 62 2129 79
rect 2054 61 2096 62
rect 1626 55 1712 61
rect 2032 55 2118 61
rect 2160 55 2164 233
rect 2348 183 2352 251
rect 2357 207 2367 241
rect 2377 213 2397 241
rect 2377 207 2391 213
rect 2416 207 2427 251
rect 2458 246 2534 253
rect 2567 251 2576 279
rect 2479 228 2513 246
rect 2521 228 2523 246
rect 2458 221 2534 228
rect 2521 213 2523 221
rect 2565 213 2576 251
rect 2640 241 2644 395
rect 2647 378 2652 412
rect 2676 378 2681 412
rect 2682 400 2693 412
rect 2896 395 2938 421
rect 3302 395 3344 421
rect 3559 420 3571 424
rect 3581 420 3593 424
rect 3631 420 3643 424
rect 3653 421 3665 424
rect 3823 421 3835 424
rect 3653 420 3706 421
rect 3664 412 3706 420
rect 3547 400 3558 412
rect 2828 341 2832 395
rect 2888 387 2934 395
rect 2888 383 2904 387
rect 2896 380 2904 383
rect 2930 380 2934 387
rect 2938 383 2946 395
rect 3294 383 3302 395
rect 3306 387 3340 395
rect 3306 380 3310 387
rect 3336 380 3340 387
rect 3344 383 3352 395
rect 2884 379 2950 380
rect 3290 379 3356 380
rect 2896 371 2900 379
rect 2950 365 3000 367
rect 3240 365 3290 367
rect 2990 361 3044 365
rect 3196 361 3250 365
rect 2990 356 3010 361
rect 3230 356 3250 361
rect 3000 341 3002 356
rect 2828 261 2832 329
rect 2896 305 2900 341
rect 2994 331 3002 341
rect 3010 331 3011 351
rect 3000 315 3002 331
rect 3021 322 3024 356
rect 3043 331 3044 351
rect 3053 331 3060 341
rect 3180 331 3187 341
rect 3196 331 3197 351
rect 3216 322 3219 356
rect 3229 331 3230 351
rect 3239 331 3246 341
rect 3010 315 3026 321
rect 3028 315 3044 321
rect 3196 315 3212 321
rect 3214 315 3230 321
rect 3290 315 3292 365
rect 2833 267 2869 295
rect 2833 261 2847 267
rect 2512 212 2523 213
rect 2357 183 2364 207
rect 2512 183 2522 212
rect 2603 207 2615 241
rect 2625 207 2645 241
rect 2348 103 2352 171
rect 2416 133 2420 183
rect 2416 98 2420 103
rect 2167 62 2172 96
rect 2196 62 2201 96
rect 2416 94 2454 98
rect 2416 79 2424 94
rect 2450 79 2454 94
rect 2538 94 2572 98
rect 2538 79 2542 94
rect 2568 79 2572 94
rect 2416 61 2458 79
rect 2534 61 2576 79
rect 2394 55 2480 61
rect 2512 55 2598 61
rect 2640 55 2644 207
rect 2670 183 2677 211
rect 2828 183 2832 251
rect 2837 233 2847 261
rect 2857 261 2871 267
rect 2896 261 2907 305
rect 3333 267 3344 305
rect 3371 267 3407 295
rect 3408 267 3412 395
rect 3559 378 3564 412
rect 3588 378 3593 412
rect 3594 400 3605 412
rect 3619 400 3630 412
rect 3631 395 3706 412
rect 3782 420 3835 421
rect 3845 420 3857 424
rect 3895 420 3907 424
rect 3917 420 3929 424
rect 3782 412 3824 420
rect 3782 395 3857 412
rect 3858 400 3869 412
rect 3883 400 3894 412
rect 3596 341 3600 395
rect 3631 378 3702 395
rect 3706 383 3714 395
rect 3774 383 3782 395
rect 3786 378 3820 395
rect 3823 378 3857 395
rect 3664 371 3668 378
rect 3058 262 3108 264
rect 3132 262 3182 264
rect 2857 233 2877 261
rect 2896 233 2905 261
rect 2959 253 2993 261
rect 2938 246 2993 253
rect 2959 245 2993 246
rect 3061 253 3092 261
rect 3061 245 3095 253
rect 2896 213 2900 233
rect 3092 229 3095 245
rect 2959 228 2993 229
rect 2938 221 2993 228
rect 3061 221 3095 229
rect 3108 212 3110 262
rect 3148 253 3179 261
rect 3182 253 3184 262
rect 3371 261 3383 267
rect 3148 245 3184 253
rect 3247 253 3281 261
rect 3247 246 3302 253
rect 3247 245 3281 246
rect 3179 229 3184 245
rect 3373 233 3383 261
rect 3393 233 3413 267
rect 3596 261 3600 329
rect 3664 291 3668 341
rect 3664 251 3673 279
rect 3760 264 3770 291
rect 3719 262 3770 264
rect 3760 261 3771 262
rect 3727 253 3761 261
rect 3769 253 3771 261
rect 3148 221 3184 229
rect 3247 228 3281 229
rect 3247 221 3302 228
rect 3182 212 3184 221
rect 2828 103 2832 171
rect 2896 133 2900 183
rect 2950 159 3000 161
rect 3240 159 3290 161
rect 3000 143 3002 159
rect 3010 153 3026 159
rect 3028 153 3044 159
rect 3196 153 3212 159
rect 3214 153 3230 159
rect 3021 143 3044 152
rect 3196 143 3219 152
rect 2994 133 3002 143
rect 3000 109 3002 133
rect 3010 123 3011 143
rect 3021 118 3024 143
rect 3043 123 3044 143
rect 3053 133 3060 143
rect 3180 133 3187 143
rect 3196 123 3197 143
rect 3216 118 3219 143
rect 3229 123 3230 143
rect 3239 133 3246 143
rect 3010 109 3044 113
rect 3196 109 3230 113
rect 3290 109 3292 159
rect 2896 103 2938 104
rect 3302 103 3344 104
rect 2896 96 2900 103
rect 2791 62 2796 96
rect 2820 62 2825 96
rect 2863 79 2934 96
rect 3306 79 3340 96
rect 3343 79 3377 96
rect 2863 62 2938 79
rect 2896 61 2938 62
rect 3302 62 3377 79
rect 3302 61 3344 62
rect 2874 55 2960 61
rect 3280 55 3366 61
rect 3408 55 3412 233
rect 3596 183 3600 251
rect 3605 207 3615 241
rect 3625 213 3645 241
rect 3625 207 3639 213
rect 3664 207 3675 251
rect 3706 246 3782 253
rect 3815 251 3824 279
rect 3727 228 3761 246
rect 3769 228 3771 246
rect 3706 221 3782 228
rect 3769 213 3771 221
rect 3813 213 3824 251
rect 3888 241 3892 395
rect 3895 378 3900 412
rect 3924 378 3929 412
rect 3930 400 3941 412
rect 4144 395 4186 421
rect 4550 395 4592 421
rect 4807 420 4819 424
rect 4829 420 4841 424
rect 4879 420 4891 424
rect 4901 421 4913 424
rect 5071 421 5083 424
rect 4901 420 4954 421
rect 4912 412 4954 420
rect 4795 400 4806 412
rect 4076 341 4080 395
rect 4136 387 4182 395
rect 4136 383 4152 387
rect 4144 380 4152 383
rect 4178 380 4182 387
rect 4186 383 4194 395
rect 4542 383 4550 395
rect 4554 387 4588 395
rect 4554 380 4558 387
rect 4584 380 4588 387
rect 4592 383 4600 395
rect 4132 379 4198 380
rect 4538 379 4604 380
rect 4144 371 4148 379
rect 4198 365 4248 367
rect 4488 365 4538 367
rect 4238 361 4292 365
rect 4444 361 4498 365
rect 4238 356 4258 361
rect 4478 356 4498 361
rect 4248 341 4250 356
rect 4076 261 4080 329
rect 4144 305 4148 341
rect 4242 331 4250 341
rect 4258 331 4259 351
rect 4248 315 4250 331
rect 4269 322 4272 356
rect 4291 331 4292 351
rect 4301 331 4308 341
rect 4428 331 4435 341
rect 4444 331 4445 351
rect 4464 322 4467 356
rect 4477 331 4478 351
rect 4487 331 4494 341
rect 4258 315 4274 321
rect 4276 315 4292 321
rect 4444 315 4460 321
rect 4462 315 4478 321
rect 4538 315 4540 365
rect 4081 267 4117 295
rect 4081 261 4095 267
rect 3760 212 3771 213
rect 3605 183 3612 207
rect 3760 183 3770 212
rect 3851 207 3863 241
rect 3873 207 3893 241
rect 3596 103 3600 171
rect 3664 133 3668 183
rect 3664 98 3668 103
rect 3415 62 3420 96
rect 3444 62 3449 96
rect 3664 94 3702 98
rect 3664 79 3672 94
rect 3698 79 3702 94
rect 3786 94 3820 98
rect 3786 79 3790 94
rect 3816 79 3820 94
rect 3664 61 3706 79
rect 3782 61 3824 79
rect 3642 55 3728 61
rect 3760 55 3846 61
rect 3888 55 3892 207
rect 3918 183 3925 211
rect 4076 183 4080 251
rect 4085 233 4095 261
rect 4105 261 4119 267
rect 4144 261 4155 305
rect 4581 267 4592 305
rect 4619 267 4655 295
rect 4656 267 4660 395
rect 4807 378 4812 412
rect 4836 378 4841 412
rect 4842 400 4853 412
rect 4867 400 4878 412
rect 4879 395 4954 412
rect 5030 420 5083 421
rect 5093 420 5105 424
rect 5143 420 5155 424
rect 5165 420 5177 424
rect 5030 412 5072 420
rect 5030 395 5105 412
rect 5106 400 5117 412
rect 5131 400 5142 412
rect 4844 341 4848 395
rect 4879 378 4950 395
rect 4954 383 4962 395
rect 5022 383 5030 395
rect 5034 378 5068 395
rect 5071 378 5105 395
rect 4912 371 4916 378
rect 4306 262 4356 264
rect 4380 262 4430 264
rect 4105 233 4125 261
rect 4144 233 4153 261
rect 4207 253 4241 261
rect 4186 246 4241 253
rect 4207 245 4241 246
rect 4309 253 4340 261
rect 4309 245 4343 253
rect 4144 213 4148 233
rect 4340 229 4343 245
rect 4207 228 4241 229
rect 4186 221 4241 228
rect 4309 221 4343 229
rect 4356 212 4358 262
rect 4396 253 4427 261
rect 4430 253 4432 262
rect 4619 261 4631 267
rect 4396 245 4432 253
rect 4495 253 4529 261
rect 4495 246 4550 253
rect 4495 245 4529 246
rect 4427 229 4432 245
rect 4621 233 4631 261
rect 4641 233 4661 267
rect 4844 261 4848 329
rect 4912 291 4916 341
rect 4912 251 4921 279
rect 5008 264 5018 291
rect 4967 262 5018 264
rect 5008 261 5019 262
rect 4975 253 5009 261
rect 5017 253 5019 261
rect 4396 221 4432 229
rect 4495 228 4529 229
rect 4495 221 4550 228
rect 4430 212 4432 221
rect 4076 103 4080 171
rect 4144 133 4148 183
rect 4198 159 4248 161
rect 4488 159 4538 161
rect 4248 143 4250 159
rect 4258 153 4274 159
rect 4276 153 4292 159
rect 4444 153 4460 159
rect 4462 153 4478 159
rect 4269 143 4292 152
rect 4444 143 4467 152
rect 4242 133 4250 143
rect 4248 109 4250 133
rect 4258 123 4259 143
rect 4269 118 4272 143
rect 4291 123 4292 143
rect 4301 133 4308 143
rect 4428 133 4435 143
rect 4444 123 4445 143
rect 4464 118 4467 143
rect 4477 123 4478 143
rect 4487 133 4494 143
rect 4258 109 4292 113
rect 4444 109 4478 113
rect 4538 109 4540 159
rect 4144 103 4186 104
rect 4550 103 4592 104
rect 4144 96 4148 103
rect 4039 62 4044 96
rect 4068 62 4073 96
rect 4111 79 4182 96
rect 4554 79 4588 96
rect 4591 79 4625 96
rect 4111 62 4186 79
rect 4144 61 4186 62
rect 4550 62 4625 79
rect 4550 61 4592 62
rect 4122 55 4208 61
rect 4528 55 4614 61
rect 4656 55 4660 233
rect 4844 183 4848 251
rect 4853 207 4863 241
rect 4873 213 4893 241
rect 4873 207 4887 213
rect 4912 207 4923 251
rect 4954 246 5030 253
rect 5063 251 5072 279
rect 4975 228 5009 246
rect 5017 228 5019 246
rect 4954 221 5030 228
rect 5017 213 5019 221
rect 5061 213 5072 251
rect 5136 241 5140 395
rect 5143 378 5148 412
rect 5172 378 5177 412
rect 5178 400 5189 412
rect 5392 395 5434 421
rect 5798 395 5840 421
rect 6055 420 6067 424
rect 6077 420 6089 424
rect 6127 420 6139 424
rect 6149 421 6161 424
rect 6319 421 6331 424
rect 6149 420 6202 421
rect 6160 412 6202 420
rect 6043 400 6054 412
rect 5324 341 5328 395
rect 5384 387 5430 395
rect 5384 383 5400 387
rect 5392 380 5400 383
rect 5426 380 5430 387
rect 5434 383 5442 395
rect 5790 383 5798 395
rect 5802 387 5836 395
rect 5802 380 5806 387
rect 5832 380 5836 387
rect 5840 383 5848 395
rect 5380 379 5446 380
rect 5786 379 5852 380
rect 5392 371 5396 379
rect 5446 365 5496 367
rect 5736 365 5786 367
rect 5486 361 5540 365
rect 5692 361 5746 365
rect 5486 356 5506 361
rect 5726 356 5746 361
rect 5496 341 5498 356
rect 5324 261 5328 329
rect 5392 305 5396 341
rect 5490 331 5498 341
rect 5506 331 5507 351
rect 5496 315 5498 331
rect 5517 322 5520 356
rect 5539 331 5540 351
rect 5549 331 5556 341
rect 5676 331 5683 341
rect 5692 331 5693 351
rect 5712 322 5715 356
rect 5725 331 5726 351
rect 5735 331 5742 341
rect 5506 315 5522 321
rect 5524 315 5540 321
rect 5692 315 5708 321
rect 5710 315 5726 321
rect 5786 315 5788 365
rect 5329 267 5365 295
rect 5329 261 5343 267
rect 5008 212 5019 213
rect 4853 183 4860 207
rect 5008 183 5018 212
rect 5099 207 5111 241
rect 5121 207 5141 241
rect 4844 103 4848 171
rect 4912 133 4916 183
rect 4912 98 4916 103
rect 4663 62 4668 96
rect 4692 62 4697 96
rect 4912 94 4950 98
rect 4912 79 4920 94
rect 4946 79 4950 94
rect 5034 94 5068 98
rect 5034 79 5038 94
rect 5064 79 5068 94
rect 4912 61 4954 79
rect 5030 61 5072 79
rect 4890 55 4976 61
rect 5008 55 5094 61
rect 5136 55 5140 207
rect 5166 183 5173 211
rect 5324 183 5328 251
rect 5333 233 5343 261
rect 5353 261 5367 267
rect 5392 261 5403 305
rect 5829 267 5840 305
rect 5867 267 5903 295
rect 5904 267 5908 395
rect 6055 378 6060 412
rect 6084 378 6089 412
rect 6090 400 6101 412
rect 6115 400 6126 412
rect 6127 395 6202 412
rect 6278 420 6331 421
rect 6341 420 6353 424
rect 6391 420 6403 424
rect 6413 420 6425 424
rect 6278 412 6320 420
rect 6278 395 6353 412
rect 6354 400 6365 412
rect 6379 400 6390 412
rect 6092 341 6096 395
rect 6127 378 6198 395
rect 6202 383 6210 395
rect 6270 383 6278 395
rect 6282 378 6316 395
rect 6319 378 6353 395
rect 6160 371 6164 378
rect 5554 262 5604 264
rect 5628 262 5678 264
rect 5353 233 5373 261
rect 5392 233 5401 261
rect 5455 253 5489 261
rect 5434 246 5489 253
rect 5455 245 5489 246
rect 5557 253 5588 261
rect 5557 245 5591 253
rect 5392 213 5396 233
rect 5588 229 5591 245
rect 5455 228 5489 229
rect 5434 221 5489 228
rect 5557 221 5591 229
rect 5604 212 5606 262
rect 5644 253 5675 261
rect 5678 253 5680 262
rect 5867 261 5879 267
rect 5644 245 5680 253
rect 5743 253 5777 261
rect 5743 246 5798 253
rect 5743 245 5777 246
rect 5675 229 5680 245
rect 5869 233 5879 261
rect 5889 233 5909 267
rect 6092 261 6096 329
rect 6160 291 6164 341
rect 6160 251 6169 279
rect 6256 264 6266 291
rect 6215 262 6266 264
rect 6256 261 6267 262
rect 6223 253 6257 261
rect 6265 253 6267 261
rect 5644 221 5680 229
rect 5743 228 5777 229
rect 5743 221 5798 228
rect 5678 212 5680 221
rect 5324 103 5328 171
rect 5392 133 5396 183
rect 5446 159 5496 161
rect 5736 159 5786 161
rect 5496 143 5498 159
rect 5506 153 5522 159
rect 5524 153 5540 159
rect 5692 153 5708 159
rect 5710 153 5726 159
rect 5517 143 5540 152
rect 5692 143 5715 152
rect 5490 133 5498 143
rect 5496 109 5498 133
rect 5506 123 5507 143
rect 5517 118 5520 143
rect 5539 123 5540 143
rect 5549 133 5556 143
rect 5676 133 5683 143
rect 5692 123 5693 143
rect 5712 118 5715 143
rect 5725 123 5726 143
rect 5735 133 5742 143
rect 5506 109 5540 113
rect 5692 109 5726 113
rect 5786 109 5788 159
rect 5392 103 5434 104
rect 5798 103 5840 104
rect 5392 96 5396 103
rect 5287 62 5292 96
rect 5316 62 5321 96
rect 5359 79 5430 96
rect 5802 79 5836 96
rect 5839 79 5873 96
rect 5359 62 5434 79
rect 5392 61 5434 62
rect 5798 62 5873 79
rect 5798 61 5840 62
rect 5370 55 5456 61
rect 5776 55 5862 61
rect 5904 55 5908 233
rect 6092 183 6096 251
rect 6101 207 6111 241
rect 6121 213 6141 241
rect 6121 207 6135 213
rect 6160 207 6171 251
rect 6202 246 6278 253
rect 6311 251 6320 279
rect 6223 228 6257 246
rect 6265 228 6267 246
rect 6202 221 6278 228
rect 6265 213 6267 221
rect 6309 213 6320 251
rect 6384 241 6388 395
rect 6391 378 6396 412
rect 6420 378 6425 412
rect 6426 400 6437 412
rect 6640 395 6682 421
rect 7046 395 7088 421
rect 7303 420 7315 424
rect 7325 420 7337 424
rect 7375 420 7387 424
rect 7397 421 7409 424
rect 7567 421 7579 424
rect 7397 420 7450 421
rect 7408 412 7450 420
rect 7291 400 7302 412
rect 6572 341 6576 395
rect 6632 387 6678 395
rect 6632 383 6648 387
rect 6640 380 6648 383
rect 6674 380 6678 387
rect 6682 383 6690 395
rect 7038 383 7046 395
rect 7050 387 7084 395
rect 7050 380 7054 387
rect 7080 380 7084 387
rect 7088 383 7096 395
rect 6628 379 6694 380
rect 7034 379 7100 380
rect 6640 371 6644 379
rect 6694 365 6744 367
rect 6984 365 7034 367
rect 6734 361 6788 365
rect 6940 361 6994 365
rect 6734 356 6754 361
rect 6974 356 6994 361
rect 6744 341 6746 356
rect 6572 261 6576 329
rect 6640 305 6644 341
rect 6738 331 6746 341
rect 6754 331 6755 351
rect 6744 315 6746 331
rect 6765 322 6768 356
rect 6787 331 6788 351
rect 6797 331 6804 341
rect 6924 331 6931 341
rect 6940 331 6941 351
rect 6960 322 6963 356
rect 6973 331 6974 351
rect 6983 331 6990 341
rect 6754 315 6770 321
rect 6772 315 6788 321
rect 6940 315 6956 321
rect 6958 315 6974 321
rect 7034 315 7036 365
rect 6577 267 6613 295
rect 6577 261 6591 267
rect 6256 212 6267 213
rect 6101 183 6108 207
rect 6256 183 6266 212
rect 6347 207 6359 241
rect 6369 207 6389 241
rect 6092 103 6096 171
rect 6160 133 6164 183
rect 6160 98 6164 103
rect 5911 62 5916 96
rect 5940 62 5945 96
rect 6160 94 6198 98
rect 6160 79 6168 94
rect 6194 79 6198 94
rect 6282 94 6316 98
rect 6282 79 6286 94
rect 6312 79 6316 94
rect 6160 61 6202 79
rect 6278 61 6320 79
rect 6138 55 6224 61
rect 6256 55 6342 61
rect 6384 55 6388 207
rect 6414 183 6421 211
rect 6572 183 6576 251
rect 6581 233 6591 261
rect 6601 261 6615 267
rect 6640 261 6651 305
rect 7077 267 7088 305
rect 7115 267 7151 295
rect 7152 267 7156 395
rect 7303 378 7308 412
rect 7332 378 7337 412
rect 7338 400 7349 412
rect 7363 400 7374 412
rect 7375 395 7450 412
rect 7526 420 7579 421
rect 7589 420 7601 424
rect 7639 420 7651 424
rect 7661 420 7673 424
rect 7526 412 7568 420
rect 7526 395 7601 412
rect 7602 400 7613 412
rect 7627 400 7638 412
rect 7340 341 7344 395
rect 7375 378 7446 395
rect 7450 383 7458 395
rect 7518 383 7526 395
rect 7530 378 7564 395
rect 7567 378 7601 395
rect 7408 371 7412 378
rect 6802 262 6852 264
rect 6876 262 6926 264
rect 6601 233 6621 261
rect 6640 233 6649 261
rect 6703 253 6737 261
rect 6682 246 6737 253
rect 6703 245 6737 246
rect 6805 253 6836 261
rect 6805 245 6839 253
rect 6640 213 6644 233
rect 6836 229 6839 245
rect 6703 228 6737 229
rect 6682 221 6737 228
rect 6805 221 6839 229
rect 6852 212 6854 262
rect 6892 253 6923 261
rect 6926 253 6928 262
rect 7115 261 7127 267
rect 6892 245 6928 253
rect 6991 253 7025 261
rect 6991 246 7046 253
rect 6991 245 7025 246
rect 6923 229 6928 245
rect 7117 233 7127 261
rect 7137 233 7157 267
rect 7340 261 7344 329
rect 7408 291 7412 341
rect 7408 251 7417 279
rect 7504 264 7514 291
rect 7463 262 7514 264
rect 7504 261 7515 262
rect 7471 253 7505 261
rect 7513 253 7515 261
rect 6892 221 6928 229
rect 6991 228 7025 229
rect 6991 221 7046 228
rect 6926 212 6928 221
rect 6572 103 6576 171
rect 6640 133 6644 183
rect 6694 159 6744 161
rect 6984 159 7034 161
rect 6744 143 6746 159
rect 6754 153 6770 159
rect 6772 153 6788 159
rect 6940 153 6956 159
rect 6958 153 6974 159
rect 6765 143 6788 152
rect 6940 143 6963 152
rect 6738 133 6746 143
rect 6744 109 6746 133
rect 6754 123 6755 143
rect 6765 118 6768 143
rect 6787 123 6788 143
rect 6797 133 6804 143
rect 6924 133 6931 143
rect 6940 123 6941 143
rect 6960 118 6963 143
rect 6973 123 6974 143
rect 6983 133 6990 143
rect 6754 109 6788 113
rect 6940 109 6974 113
rect 7034 109 7036 159
rect 6640 103 6682 104
rect 7046 103 7088 104
rect 6640 96 6644 103
rect 6535 62 6540 96
rect 6564 62 6569 96
rect 6607 79 6678 96
rect 7050 79 7084 96
rect 7087 79 7121 96
rect 6607 62 6682 79
rect 6640 61 6682 62
rect 7046 62 7121 79
rect 7046 61 7088 62
rect 6618 55 6704 61
rect 7024 55 7110 61
rect 7152 55 7156 233
rect 7340 183 7344 251
rect 7349 207 7359 241
rect 7369 213 7389 241
rect 7369 207 7383 213
rect 7408 207 7419 251
rect 7450 246 7526 253
rect 7559 251 7568 279
rect 7471 228 7505 246
rect 7513 228 7515 246
rect 7450 221 7526 228
rect 7513 213 7515 221
rect 7557 213 7568 251
rect 7632 241 7636 395
rect 7639 378 7644 412
rect 7668 378 7673 412
rect 7674 400 7685 412
rect 7888 395 7930 421
rect 8294 395 8336 421
rect 8551 420 8563 424
rect 8573 420 8585 424
rect 8623 420 8635 424
rect 8645 421 8657 424
rect 8815 421 8827 424
rect 8645 420 8698 421
rect 8656 412 8698 420
rect 8539 400 8550 412
rect 7820 341 7824 395
rect 7880 387 7926 395
rect 7880 383 7896 387
rect 7888 380 7896 383
rect 7922 380 7926 387
rect 7930 383 7938 395
rect 8286 383 8294 395
rect 8298 387 8332 395
rect 8298 380 8302 387
rect 8328 380 8332 387
rect 8336 383 8344 395
rect 7876 379 7942 380
rect 8282 379 8348 380
rect 7888 371 7892 379
rect 7942 365 7992 367
rect 8232 365 8282 367
rect 7982 361 8036 365
rect 8188 361 8242 365
rect 7982 356 8002 361
rect 8222 356 8242 361
rect 7992 341 7994 356
rect 7820 261 7824 329
rect 7888 305 7892 341
rect 7986 331 7994 341
rect 8002 331 8003 351
rect 7992 315 7994 331
rect 8013 322 8016 356
rect 8035 331 8036 351
rect 8045 331 8052 341
rect 8172 331 8179 341
rect 8188 331 8189 351
rect 8208 322 8211 356
rect 8221 331 8222 351
rect 8231 331 8238 341
rect 8002 315 8018 321
rect 8020 315 8036 321
rect 8188 315 8204 321
rect 8206 315 8222 321
rect 8282 315 8284 365
rect 7825 267 7861 295
rect 7825 261 7839 267
rect 7504 212 7515 213
rect 7349 183 7356 207
rect 7504 183 7514 212
rect 7595 207 7607 241
rect 7617 207 7637 241
rect 7340 103 7344 171
rect 7408 133 7412 183
rect 7408 98 7412 103
rect 7159 62 7164 96
rect 7188 62 7193 96
rect 7408 94 7446 98
rect 7408 79 7416 94
rect 7442 79 7446 94
rect 7530 94 7564 98
rect 7530 79 7534 94
rect 7560 79 7564 94
rect 7408 61 7450 79
rect 7526 61 7568 79
rect 7386 55 7472 61
rect 7504 55 7590 61
rect 7632 55 7636 207
rect 7662 183 7669 211
rect 7820 183 7824 251
rect 7829 233 7839 261
rect 7849 261 7863 267
rect 7888 261 7899 305
rect 8325 267 8336 305
rect 8363 267 8399 295
rect 8400 267 8404 395
rect 8551 378 8556 412
rect 8580 378 8585 412
rect 8586 400 8597 412
rect 8611 400 8622 412
rect 8623 395 8698 412
rect 8774 420 8827 421
rect 8837 420 8849 424
rect 8887 420 8899 424
rect 8909 420 8921 424
rect 8774 412 8816 420
rect 8774 395 8849 412
rect 8850 400 8861 412
rect 8875 400 8886 412
rect 8588 341 8592 395
rect 8623 378 8694 395
rect 8698 383 8706 395
rect 8766 383 8774 395
rect 8778 378 8812 395
rect 8815 378 8849 395
rect 8656 371 8660 378
rect 8050 262 8100 264
rect 8124 262 8174 264
rect 7849 233 7869 261
rect 7888 233 7897 261
rect 7951 253 7985 261
rect 7930 246 7985 253
rect 7951 245 7985 246
rect 8053 253 8084 261
rect 8053 245 8087 253
rect 7888 213 7892 233
rect 8084 229 8087 245
rect 7951 228 7985 229
rect 7930 221 7985 228
rect 8053 221 8087 229
rect 8100 212 8102 262
rect 8140 253 8171 261
rect 8174 253 8176 262
rect 8363 261 8375 267
rect 8140 245 8176 253
rect 8239 253 8273 261
rect 8239 246 8294 253
rect 8239 245 8273 246
rect 8171 229 8176 245
rect 8365 233 8375 261
rect 8385 233 8405 267
rect 8588 261 8592 329
rect 8656 291 8660 341
rect 8656 251 8665 279
rect 8752 264 8762 291
rect 8711 262 8762 264
rect 8752 261 8763 262
rect 8719 253 8753 261
rect 8761 253 8763 261
rect 8140 221 8176 229
rect 8239 228 8273 229
rect 8239 221 8294 228
rect 8174 212 8176 221
rect 7820 103 7824 171
rect 7888 133 7892 183
rect 7942 159 7992 161
rect 8232 159 8282 161
rect 7992 143 7994 159
rect 8002 153 8018 159
rect 8020 153 8036 159
rect 8188 153 8204 159
rect 8206 153 8222 159
rect 8013 143 8036 152
rect 8188 143 8211 152
rect 7986 133 7994 143
rect 7992 109 7994 133
rect 8002 123 8003 143
rect 8013 118 8016 143
rect 8035 123 8036 143
rect 8045 133 8052 143
rect 8172 133 8179 143
rect 8188 123 8189 143
rect 8208 118 8211 143
rect 8221 123 8222 143
rect 8231 133 8238 143
rect 8002 109 8036 113
rect 8188 109 8222 113
rect 8282 109 8284 159
rect 7888 103 7930 104
rect 8294 103 8336 104
rect 7888 96 7892 103
rect 7783 62 7788 96
rect 7812 62 7817 96
rect 7855 79 7926 96
rect 8298 79 8332 96
rect 8335 79 8369 96
rect 7855 62 7930 79
rect 7888 61 7930 62
rect 8294 62 8369 79
rect 8294 61 8336 62
rect 7866 55 7952 61
rect 8272 55 8358 61
rect 8400 55 8404 233
rect 8588 183 8592 251
rect 8597 207 8607 241
rect 8617 213 8637 241
rect 8617 207 8631 213
rect 8656 207 8667 251
rect 8698 246 8774 253
rect 8807 251 8816 279
rect 8719 228 8753 246
rect 8761 228 8763 246
rect 8698 221 8774 228
rect 8761 213 8763 221
rect 8805 213 8816 251
rect 8880 241 8884 395
rect 8887 378 8892 412
rect 8916 378 8921 412
rect 8922 400 8933 412
rect 9136 395 9178 421
rect 9542 395 9584 421
rect 9799 420 9811 424
rect 9821 420 9833 424
rect 9871 420 9883 424
rect 9893 421 9905 424
rect 10063 421 10075 424
rect 9893 420 9946 421
rect 9904 412 9946 420
rect 9787 400 9798 412
rect 9068 341 9072 395
rect 9128 387 9174 395
rect 9128 383 9144 387
rect 9136 380 9144 383
rect 9170 380 9174 387
rect 9178 383 9186 395
rect 9534 383 9542 395
rect 9546 387 9580 395
rect 9546 380 9550 387
rect 9576 380 9580 387
rect 9584 383 9592 395
rect 9124 379 9190 380
rect 9530 379 9596 380
rect 9136 371 9140 379
rect 9190 365 9240 367
rect 9480 365 9530 367
rect 9230 361 9284 365
rect 9436 361 9490 365
rect 9230 356 9250 361
rect 9470 356 9490 361
rect 9240 341 9242 356
rect 9068 261 9072 329
rect 9136 305 9140 341
rect 9234 331 9242 341
rect 9250 331 9251 351
rect 9240 315 9242 331
rect 9261 322 9264 356
rect 9283 331 9284 351
rect 9293 331 9300 341
rect 9420 331 9427 341
rect 9436 331 9437 351
rect 9456 322 9459 356
rect 9469 331 9470 351
rect 9479 331 9486 341
rect 9250 315 9266 321
rect 9268 315 9284 321
rect 9436 315 9452 321
rect 9454 315 9470 321
rect 9530 315 9532 365
rect 9073 267 9109 295
rect 9073 261 9087 267
rect 8752 212 8763 213
rect 8597 183 8604 207
rect 8752 183 8762 212
rect 8843 207 8855 241
rect 8865 207 8885 241
rect 8588 103 8592 171
rect 8656 133 8660 183
rect 8656 98 8660 103
rect 8407 62 8412 96
rect 8436 62 8441 96
rect 8656 94 8694 98
rect 8656 79 8664 94
rect 8690 79 8694 94
rect 8778 94 8812 98
rect 8778 79 8782 94
rect 8808 79 8812 94
rect 8656 61 8698 79
rect 8774 61 8816 79
rect 8634 55 8720 61
rect 8752 55 8838 61
rect 8880 55 8884 207
rect 8910 183 8917 211
rect 9068 183 9072 251
rect 9077 233 9087 261
rect 9097 261 9111 267
rect 9136 261 9147 305
rect 9573 267 9584 305
rect 9611 267 9647 295
rect 9648 267 9652 395
rect 9799 378 9804 412
rect 9828 378 9833 412
rect 9834 400 9845 412
rect 9859 400 9870 412
rect 9871 395 9946 412
rect 10022 420 10075 421
rect 10085 420 10097 424
rect 10135 420 10147 424
rect 10157 420 10169 424
rect 10022 412 10064 420
rect 10022 395 10097 412
rect 10098 400 10109 412
rect 10123 400 10134 412
rect 9836 341 9840 395
rect 9871 378 9942 395
rect 9946 383 9954 395
rect 10014 383 10022 395
rect 10026 378 10060 395
rect 10063 378 10097 395
rect 9904 371 9908 378
rect 9298 262 9348 264
rect 9372 262 9422 264
rect 9097 233 9117 261
rect 9136 233 9145 261
rect 9199 253 9233 261
rect 9178 246 9233 253
rect 9199 245 9233 246
rect 9301 253 9332 261
rect 9301 245 9335 253
rect 9136 213 9140 233
rect 9332 229 9335 245
rect 9199 228 9233 229
rect 9178 221 9233 228
rect 9301 221 9335 229
rect 9348 212 9350 262
rect 9388 253 9419 261
rect 9422 253 9424 262
rect 9611 261 9623 267
rect 9388 245 9424 253
rect 9487 253 9521 261
rect 9487 246 9542 253
rect 9487 245 9521 246
rect 9419 229 9424 245
rect 9613 233 9623 261
rect 9633 233 9653 267
rect 9836 261 9840 329
rect 9904 291 9908 341
rect 9904 251 9913 279
rect 10000 264 10010 291
rect 9959 262 10010 264
rect 10000 261 10011 262
rect 9967 253 10001 261
rect 10009 253 10011 261
rect 9388 221 9424 229
rect 9487 228 9521 229
rect 9487 221 9542 228
rect 9422 212 9424 221
rect 9068 103 9072 171
rect 9136 133 9140 183
rect 9190 159 9240 161
rect 9480 159 9530 161
rect 9240 143 9242 159
rect 9250 153 9266 159
rect 9268 153 9284 159
rect 9436 153 9452 159
rect 9454 153 9470 159
rect 9261 143 9284 152
rect 9436 143 9459 152
rect 9234 133 9242 143
rect 9240 109 9242 133
rect 9250 123 9251 143
rect 9261 118 9264 143
rect 9283 123 9284 143
rect 9293 133 9300 143
rect 9420 133 9427 143
rect 9436 123 9437 143
rect 9456 118 9459 143
rect 9469 123 9470 143
rect 9479 133 9486 143
rect 9250 109 9284 113
rect 9436 109 9470 113
rect 9530 109 9532 159
rect 9136 103 9178 104
rect 9542 103 9584 104
rect 9136 96 9140 103
rect 9031 62 9036 96
rect 9060 62 9065 96
rect 9103 79 9174 96
rect 9546 79 9580 96
rect 9583 79 9617 96
rect 9103 62 9178 79
rect 9136 61 9178 62
rect 9542 62 9617 79
rect 9542 61 9584 62
rect 9114 55 9200 61
rect 9520 55 9606 61
rect 9648 55 9652 233
rect 9836 183 9840 251
rect 9845 207 9855 241
rect 9865 213 9885 241
rect 9865 207 9879 213
rect 9904 207 9915 251
rect 9946 246 10022 253
rect 10055 251 10064 279
rect 9967 228 10001 246
rect 10009 228 10011 246
rect 9946 221 10022 228
rect 10009 213 10011 221
rect 10053 213 10064 251
rect 10128 241 10132 395
rect 10135 378 10140 412
rect 10164 378 10169 412
rect 10170 400 10181 412
rect 10384 395 10426 421
rect 10790 395 10832 421
rect 11047 420 11059 424
rect 11069 420 11081 424
rect 11119 420 11131 424
rect 11141 421 11153 424
rect 11311 421 11323 424
rect 11141 420 11194 421
rect 11152 412 11194 420
rect 11035 400 11046 412
rect 10316 341 10320 395
rect 10376 387 10422 395
rect 10376 383 10392 387
rect 10384 380 10392 383
rect 10418 380 10422 387
rect 10426 383 10434 395
rect 10782 383 10790 395
rect 10794 387 10828 395
rect 10794 380 10798 387
rect 10824 380 10828 387
rect 10832 383 10840 395
rect 10372 379 10438 380
rect 10778 379 10844 380
rect 10384 371 10388 379
rect 10438 365 10488 367
rect 10728 365 10778 367
rect 10478 361 10532 365
rect 10684 361 10738 365
rect 10478 356 10498 361
rect 10718 356 10738 361
rect 10488 341 10490 356
rect 10316 261 10320 329
rect 10384 305 10388 341
rect 10482 331 10490 341
rect 10498 331 10499 351
rect 10488 315 10490 331
rect 10509 322 10512 356
rect 10531 331 10532 351
rect 10541 331 10548 341
rect 10668 331 10675 341
rect 10684 331 10685 351
rect 10704 322 10707 356
rect 10717 331 10718 351
rect 10727 331 10734 341
rect 10498 315 10514 321
rect 10516 315 10532 321
rect 10684 315 10700 321
rect 10702 315 10718 321
rect 10778 315 10780 365
rect 10321 267 10357 295
rect 10321 261 10335 267
rect 10000 212 10011 213
rect 9845 183 9852 207
rect 10000 183 10010 212
rect 10091 207 10103 241
rect 10113 207 10133 241
rect 9836 103 9840 171
rect 9904 133 9908 183
rect 9904 98 9908 103
rect 9655 62 9660 96
rect 9684 62 9689 96
rect 9904 94 9942 98
rect 9904 79 9912 94
rect 9938 79 9942 94
rect 10026 94 10060 98
rect 10026 79 10030 94
rect 10056 79 10060 94
rect 9904 61 9946 79
rect 10022 61 10064 79
rect 9882 55 9968 61
rect 10000 55 10086 61
rect 10128 55 10132 207
rect 10158 183 10165 211
rect 10316 183 10320 251
rect 10325 233 10335 261
rect 10345 261 10359 267
rect 10384 261 10395 305
rect 10821 267 10832 305
rect 10859 267 10895 295
rect 10896 267 10900 395
rect 11047 378 11052 412
rect 11076 378 11081 412
rect 11082 400 11093 412
rect 11107 400 11118 412
rect 11119 395 11194 412
rect 11270 420 11323 421
rect 11333 420 11345 424
rect 11383 420 11395 424
rect 11405 420 11417 424
rect 11270 412 11312 420
rect 11270 395 11345 412
rect 11346 400 11357 412
rect 11371 400 11382 412
rect 11084 341 11088 395
rect 11119 378 11190 395
rect 11194 383 11202 395
rect 11262 383 11270 395
rect 11274 378 11308 395
rect 11311 378 11345 395
rect 11152 371 11156 378
rect 10546 262 10596 264
rect 10620 262 10670 264
rect 10345 233 10365 261
rect 10384 233 10393 261
rect 10447 253 10481 261
rect 10426 246 10481 253
rect 10447 245 10481 246
rect 10549 253 10580 261
rect 10549 245 10583 253
rect 10384 213 10388 233
rect 10580 229 10583 245
rect 10447 228 10481 229
rect 10426 221 10481 228
rect 10549 221 10583 229
rect 10596 212 10598 262
rect 10636 253 10667 261
rect 10670 253 10672 262
rect 10859 261 10871 267
rect 10636 245 10672 253
rect 10735 253 10769 261
rect 10735 246 10790 253
rect 10735 245 10769 246
rect 10667 229 10672 245
rect 10861 233 10871 261
rect 10881 233 10901 267
rect 11084 261 11088 329
rect 11152 291 11156 341
rect 11152 251 11161 279
rect 11248 264 11258 291
rect 11207 262 11258 264
rect 11248 261 11259 262
rect 11215 253 11249 261
rect 11257 253 11259 261
rect 10636 221 10672 229
rect 10735 228 10769 229
rect 10735 221 10790 228
rect 10670 212 10672 221
rect 10316 103 10320 171
rect 10384 133 10388 183
rect 10438 159 10488 161
rect 10728 159 10778 161
rect 10488 143 10490 159
rect 10498 153 10514 159
rect 10516 153 10532 159
rect 10684 153 10700 159
rect 10702 153 10718 159
rect 10509 143 10532 152
rect 10684 143 10707 152
rect 10482 133 10490 143
rect 10488 109 10490 133
rect 10498 123 10499 143
rect 10509 118 10512 143
rect 10531 123 10532 143
rect 10541 133 10548 143
rect 10668 133 10675 143
rect 10684 123 10685 143
rect 10704 118 10707 143
rect 10717 123 10718 143
rect 10727 133 10734 143
rect 10498 109 10532 113
rect 10684 109 10718 113
rect 10778 109 10780 159
rect 10384 103 10426 104
rect 10790 103 10832 104
rect 10384 96 10388 103
rect 10279 62 10284 96
rect 10308 62 10313 96
rect 10351 79 10422 96
rect 10794 79 10828 96
rect 10831 79 10865 96
rect 10351 62 10426 79
rect 10384 61 10426 62
rect 10790 62 10865 79
rect 10790 61 10832 62
rect 10362 55 10448 61
rect 10768 55 10854 61
rect 10896 55 10900 233
rect 11084 183 11088 251
rect 11093 207 11103 241
rect 11113 213 11133 241
rect 11113 207 11127 213
rect 11152 207 11163 251
rect 11194 246 11270 253
rect 11303 251 11312 279
rect 11215 228 11249 246
rect 11257 228 11259 246
rect 11194 221 11270 228
rect 11257 213 11259 221
rect 11301 213 11312 251
rect 11376 241 11380 395
rect 11383 378 11388 412
rect 11412 378 11417 412
rect 11418 400 11429 412
rect 11632 395 11674 421
rect 12038 395 12080 421
rect 12295 420 12307 424
rect 12317 420 12329 424
rect 12367 420 12379 424
rect 12389 421 12401 424
rect 12559 421 12571 424
rect 12389 420 12442 421
rect 12400 412 12442 420
rect 12283 400 12294 412
rect 11564 341 11568 395
rect 11624 387 11670 395
rect 11624 383 11640 387
rect 11632 380 11640 383
rect 11666 380 11670 387
rect 11674 383 11682 395
rect 12030 383 12038 395
rect 12042 387 12076 395
rect 12042 380 12046 387
rect 12072 380 12076 387
rect 12080 383 12088 395
rect 11620 379 11686 380
rect 12026 379 12092 380
rect 11632 371 11636 379
rect 11686 365 11736 367
rect 11976 365 12026 367
rect 11726 361 11780 365
rect 11932 361 11986 365
rect 11726 356 11746 361
rect 11966 356 11986 361
rect 11736 341 11738 356
rect 11564 261 11568 329
rect 11632 305 11636 341
rect 11730 331 11738 341
rect 11746 331 11747 351
rect 11736 315 11738 331
rect 11757 322 11760 356
rect 11779 331 11780 351
rect 11789 331 11796 341
rect 11916 331 11923 341
rect 11932 331 11933 351
rect 11952 322 11955 356
rect 11965 331 11966 351
rect 11975 331 11982 341
rect 11746 315 11762 321
rect 11764 315 11780 321
rect 11932 315 11948 321
rect 11950 315 11966 321
rect 12026 315 12028 365
rect 11569 267 11605 295
rect 11569 261 11583 267
rect 11248 212 11259 213
rect 11093 183 11100 207
rect 11248 183 11258 212
rect 11339 207 11351 241
rect 11361 207 11381 241
rect 11084 103 11088 171
rect 11152 133 11156 183
rect 11152 98 11156 103
rect 10903 62 10908 96
rect 10932 62 10937 96
rect 11152 94 11190 98
rect 11152 79 11160 94
rect 11186 79 11190 94
rect 11274 94 11308 98
rect 11274 79 11278 94
rect 11304 79 11308 94
rect 11152 61 11194 79
rect 11270 61 11312 79
rect 11130 55 11216 61
rect 11248 55 11334 61
rect 11376 55 11380 207
rect 11406 183 11413 211
rect 11564 183 11568 251
rect 11573 233 11583 261
rect 11593 261 11607 267
rect 11632 261 11643 305
rect 12069 267 12080 305
rect 12107 267 12143 295
rect 12144 267 12148 395
rect 12295 378 12300 412
rect 12324 378 12329 412
rect 12330 400 12341 412
rect 12355 400 12366 412
rect 12367 395 12442 412
rect 12518 420 12571 421
rect 12581 420 12593 424
rect 12631 420 12643 424
rect 12653 420 12665 424
rect 12518 412 12560 420
rect 12518 395 12593 412
rect 12594 400 12605 412
rect 12619 400 12630 412
rect 12332 341 12336 395
rect 12367 378 12438 395
rect 12442 383 12450 395
rect 12510 383 12518 395
rect 12522 378 12556 395
rect 12559 378 12593 395
rect 12400 371 12404 378
rect 11794 262 11844 264
rect 11868 262 11918 264
rect 11593 233 11613 261
rect 11632 233 11641 261
rect 11695 253 11729 261
rect 11674 246 11729 253
rect 11695 245 11729 246
rect 11797 253 11828 261
rect 11797 245 11831 253
rect 11632 213 11636 233
rect 11828 229 11831 245
rect 11695 228 11729 229
rect 11674 221 11729 228
rect 11797 221 11831 229
rect 11844 212 11846 262
rect 11884 253 11915 261
rect 11918 253 11920 262
rect 12107 261 12119 267
rect 11884 245 11920 253
rect 11983 253 12017 261
rect 11983 246 12038 253
rect 11983 245 12017 246
rect 11915 229 11920 245
rect 12109 233 12119 261
rect 12129 233 12149 267
rect 12332 261 12336 329
rect 12400 291 12404 341
rect 12400 251 12409 279
rect 12496 264 12506 291
rect 12455 262 12506 264
rect 12496 261 12507 262
rect 12463 253 12497 261
rect 12505 253 12507 261
rect 11884 221 11920 229
rect 11983 228 12017 229
rect 11983 221 12038 228
rect 11918 212 11920 221
rect 11564 103 11568 171
rect 11632 133 11636 183
rect 11686 159 11736 161
rect 11976 159 12026 161
rect 11736 143 11738 159
rect 11746 153 11762 159
rect 11764 153 11780 159
rect 11932 153 11948 159
rect 11950 153 11966 159
rect 11757 143 11780 152
rect 11932 143 11955 152
rect 11730 133 11738 143
rect 11736 109 11738 133
rect 11746 123 11747 143
rect 11757 118 11760 143
rect 11779 123 11780 143
rect 11789 133 11796 143
rect 11916 133 11923 143
rect 11932 123 11933 143
rect 11952 118 11955 143
rect 11965 123 11966 143
rect 11975 133 11982 143
rect 11746 109 11780 113
rect 11932 109 11966 113
rect 12026 109 12028 159
rect 11632 103 11674 104
rect 12038 103 12080 104
rect 11632 96 11636 103
rect 11527 62 11532 96
rect 11556 62 11561 96
rect 11599 79 11670 96
rect 12042 79 12076 96
rect 12079 79 12113 96
rect 11599 62 11674 79
rect 11632 61 11674 62
rect 12038 62 12113 79
rect 12038 61 12080 62
rect 11610 55 11696 61
rect 12016 55 12102 61
rect 12144 55 12148 233
rect 12332 183 12336 251
rect 12341 207 12351 241
rect 12361 213 12381 241
rect 12361 207 12375 213
rect 12400 207 12411 251
rect 12442 246 12518 253
rect 12551 251 12560 279
rect 12463 228 12497 246
rect 12505 228 12507 246
rect 12442 221 12518 228
rect 12505 213 12507 221
rect 12549 213 12560 251
rect 12624 241 12628 395
rect 12631 378 12636 412
rect 12660 378 12665 412
rect 12666 400 12677 412
rect 12880 395 12922 421
rect 13286 395 13328 421
rect 13543 420 13555 424
rect 13565 420 13577 424
rect 13615 420 13627 424
rect 13637 421 13649 424
rect 13807 421 13819 424
rect 13637 420 13690 421
rect 13648 412 13690 420
rect 13531 400 13542 412
rect 12812 341 12816 395
rect 12872 387 12918 395
rect 12872 383 12888 387
rect 12880 380 12888 383
rect 12914 380 12918 387
rect 12922 383 12930 395
rect 13278 383 13286 395
rect 13290 387 13324 395
rect 13290 380 13294 387
rect 13320 380 13324 387
rect 13328 383 13336 395
rect 12868 379 12934 380
rect 13274 379 13340 380
rect 12880 371 12884 379
rect 12934 365 12984 367
rect 13224 365 13274 367
rect 12974 361 13028 365
rect 13180 361 13234 365
rect 12974 356 12994 361
rect 13214 356 13234 361
rect 12984 341 12986 356
rect 12812 261 12816 329
rect 12880 305 12884 341
rect 12978 331 12986 341
rect 12994 331 12995 351
rect 12984 315 12986 331
rect 13005 322 13008 356
rect 13027 331 13028 351
rect 13037 331 13044 341
rect 13164 331 13171 341
rect 13180 331 13181 351
rect 13200 322 13203 356
rect 13213 331 13214 351
rect 13223 331 13230 341
rect 12994 315 13010 321
rect 13012 315 13028 321
rect 13180 315 13196 321
rect 13198 315 13214 321
rect 13274 315 13276 365
rect 12817 267 12853 295
rect 12817 261 12831 267
rect 12496 212 12507 213
rect 12341 183 12348 207
rect 12496 183 12506 212
rect 12587 207 12599 241
rect 12609 207 12629 241
rect 12332 103 12336 171
rect 12400 133 12404 183
rect 12400 98 12404 103
rect 12151 62 12156 96
rect 12180 62 12185 96
rect 12400 94 12438 98
rect 12400 79 12408 94
rect 12434 79 12438 94
rect 12522 94 12556 98
rect 12522 79 12526 94
rect 12552 79 12556 94
rect 12400 61 12442 79
rect 12518 61 12560 79
rect 12378 55 12464 61
rect 12496 55 12582 61
rect 12624 55 12628 207
rect 12654 183 12661 211
rect 12812 183 12816 251
rect 12821 233 12831 261
rect 12841 261 12855 267
rect 12880 261 12891 305
rect 13317 267 13328 305
rect 13355 267 13391 295
rect 13392 267 13396 395
rect 13543 378 13548 412
rect 13572 378 13577 412
rect 13578 400 13589 412
rect 13603 400 13614 412
rect 13615 395 13690 412
rect 13766 420 13819 421
rect 13829 420 13841 424
rect 13879 420 13891 424
rect 13901 420 13913 424
rect 13766 412 13808 420
rect 13766 395 13841 412
rect 13842 400 13853 412
rect 13867 400 13878 412
rect 13580 341 13584 395
rect 13615 378 13686 395
rect 13690 383 13698 395
rect 13758 383 13766 395
rect 13770 378 13804 395
rect 13807 378 13841 395
rect 13648 371 13652 378
rect 13042 262 13092 264
rect 13116 262 13166 264
rect 12841 233 12861 261
rect 12880 233 12889 261
rect 12943 253 12977 261
rect 12922 246 12977 253
rect 12943 245 12977 246
rect 13045 253 13076 261
rect 13045 245 13079 253
rect 12880 213 12884 233
rect 13076 229 13079 245
rect 12943 228 12977 229
rect 12922 221 12977 228
rect 13045 221 13079 229
rect 13092 212 13094 262
rect 13132 253 13163 261
rect 13166 253 13168 262
rect 13355 261 13367 267
rect 13132 245 13168 253
rect 13231 253 13265 261
rect 13231 246 13286 253
rect 13231 245 13265 246
rect 13163 229 13168 245
rect 13357 233 13367 261
rect 13377 233 13397 267
rect 13580 261 13584 329
rect 13648 291 13652 341
rect 13648 251 13657 279
rect 13744 264 13754 291
rect 13703 262 13754 264
rect 13744 261 13755 262
rect 13711 253 13745 261
rect 13753 253 13755 261
rect 13132 221 13168 229
rect 13231 228 13265 229
rect 13231 221 13286 228
rect 13166 212 13168 221
rect 12812 103 12816 171
rect 12880 133 12884 183
rect 12934 159 12984 161
rect 13224 159 13274 161
rect 12984 143 12986 159
rect 12994 153 13010 159
rect 13012 153 13028 159
rect 13180 153 13196 159
rect 13198 153 13214 159
rect 13005 143 13028 152
rect 13180 143 13203 152
rect 12978 133 12986 143
rect 12984 109 12986 133
rect 12994 123 12995 143
rect 13005 118 13008 143
rect 13027 123 13028 143
rect 13037 133 13044 143
rect 13164 133 13171 143
rect 13180 123 13181 143
rect 13200 118 13203 143
rect 13213 123 13214 143
rect 13223 133 13230 143
rect 12994 109 13028 113
rect 13180 109 13214 113
rect 13274 109 13276 159
rect 12880 103 12922 104
rect 13286 103 13328 104
rect 12880 96 12884 103
rect 12775 62 12780 96
rect 12804 62 12809 96
rect 12847 79 12918 96
rect 13290 79 13324 96
rect 13327 79 13361 96
rect 12847 62 12922 79
rect 12880 61 12922 62
rect 13286 62 13361 79
rect 13286 61 13328 62
rect 12858 55 12944 61
rect 13264 55 13350 61
rect 13392 55 13396 233
rect 13580 183 13584 251
rect 13589 207 13599 241
rect 13609 213 13629 241
rect 13609 207 13623 213
rect 13648 207 13659 251
rect 13690 246 13766 253
rect 13799 251 13808 279
rect 13711 228 13745 246
rect 13753 228 13755 246
rect 13690 221 13766 228
rect 13753 213 13755 221
rect 13797 213 13808 251
rect 13872 241 13876 395
rect 13879 378 13884 412
rect 13908 378 13913 412
rect 13914 400 13925 412
rect 14128 395 14170 421
rect 14534 395 14576 421
rect 14791 420 14803 424
rect 14813 420 14825 424
rect 14863 420 14875 424
rect 14885 421 14897 424
rect 15055 421 15067 424
rect 14885 420 14938 421
rect 14896 412 14938 420
rect 14779 400 14790 412
rect 14060 341 14064 395
rect 14120 387 14166 395
rect 14120 383 14136 387
rect 14128 380 14136 383
rect 14162 380 14166 387
rect 14170 383 14178 395
rect 14526 383 14534 395
rect 14538 387 14572 395
rect 14538 380 14542 387
rect 14568 380 14572 387
rect 14576 383 14584 395
rect 14116 379 14182 380
rect 14522 379 14588 380
rect 14128 371 14132 379
rect 14182 365 14232 367
rect 14472 365 14522 367
rect 14222 361 14276 365
rect 14428 361 14482 365
rect 14222 356 14242 361
rect 14462 356 14482 361
rect 14232 341 14234 356
rect 14060 261 14064 329
rect 14128 305 14132 341
rect 14226 331 14234 341
rect 14242 331 14243 351
rect 14232 315 14234 331
rect 14253 322 14256 356
rect 14275 331 14276 351
rect 14285 331 14292 341
rect 14412 331 14419 341
rect 14428 331 14429 351
rect 14448 322 14451 356
rect 14461 331 14462 351
rect 14471 331 14478 341
rect 14242 315 14258 321
rect 14260 315 14276 321
rect 14428 315 14444 321
rect 14446 315 14462 321
rect 14522 315 14524 365
rect 14065 267 14101 295
rect 14065 261 14079 267
rect 13744 212 13755 213
rect 13589 183 13596 207
rect 13744 183 13754 212
rect 13835 207 13847 241
rect 13857 207 13877 241
rect 13580 103 13584 171
rect 13648 133 13652 183
rect 13648 98 13652 103
rect 13399 62 13404 96
rect 13428 62 13433 96
rect 13648 94 13686 98
rect 13648 79 13656 94
rect 13682 79 13686 94
rect 13770 94 13804 98
rect 13770 79 13774 94
rect 13800 79 13804 94
rect 13648 61 13690 79
rect 13766 61 13808 79
rect 13626 55 13712 61
rect 13744 55 13830 61
rect 13872 55 13876 207
rect 13902 183 13909 211
rect 14060 183 14064 251
rect 14069 233 14079 261
rect 14089 261 14103 267
rect 14128 261 14139 305
rect 14565 267 14576 305
rect 14603 267 14639 295
rect 14640 267 14644 395
rect 14791 378 14796 412
rect 14820 378 14825 412
rect 14826 400 14837 412
rect 14851 400 14862 412
rect 14863 395 14938 412
rect 15014 420 15067 421
rect 15077 420 15089 424
rect 15127 420 15139 424
rect 15149 420 15161 424
rect 15014 412 15056 420
rect 15014 395 15089 412
rect 15090 400 15101 412
rect 15115 400 15126 412
rect 14828 341 14832 395
rect 14863 378 14934 395
rect 14938 383 14946 395
rect 15006 383 15014 395
rect 15018 378 15052 395
rect 15055 378 15089 395
rect 14896 371 14900 378
rect 14290 262 14340 264
rect 14364 262 14414 264
rect 14089 233 14109 261
rect 14128 233 14137 261
rect 14191 253 14225 261
rect 14170 246 14225 253
rect 14191 245 14225 246
rect 14293 253 14324 261
rect 14293 245 14327 253
rect 14128 213 14132 233
rect 14324 229 14327 245
rect 14191 228 14225 229
rect 14170 221 14225 228
rect 14293 221 14327 229
rect 14340 212 14342 262
rect 14380 253 14411 261
rect 14414 253 14416 262
rect 14603 261 14615 267
rect 14380 245 14416 253
rect 14479 253 14513 261
rect 14479 246 14534 253
rect 14479 245 14513 246
rect 14411 229 14416 245
rect 14605 233 14615 261
rect 14625 233 14645 267
rect 14828 261 14832 329
rect 14896 291 14900 341
rect 14896 251 14905 279
rect 14992 264 15002 291
rect 14951 262 15002 264
rect 14992 261 15003 262
rect 14959 253 14993 261
rect 15001 253 15003 261
rect 14380 221 14416 229
rect 14479 228 14513 229
rect 14479 221 14534 228
rect 14414 212 14416 221
rect 14060 103 14064 171
rect 14128 133 14132 183
rect 14182 159 14232 161
rect 14472 159 14522 161
rect 14232 143 14234 159
rect 14242 153 14258 159
rect 14260 153 14276 159
rect 14428 153 14444 159
rect 14446 153 14462 159
rect 14253 143 14276 152
rect 14428 143 14451 152
rect 14226 133 14234 143
rect 14232 109 14234 133
rect 14242 123 14243 143
rect 14253 118 14256 143
rect 14275 123 14276 143
rect 14285 133 14292 143
rect 14412 133 14419 143
rect 14428 123 14429 143
rect 14448 118 14451 143
rect 14461 123 14462 143
rect 14471 133 14478 143
rect 14242 109 14276 113
rect 14428 109 14462 113
rect 14522 109 14524 159
rect 14128 103 14170 104
rect 14534 103 14576 104
rect 14128 96 14132 103
rect 14023 62 14028 96
rect 14052 62 14057 96
rect 14095 79 14166 96
rect 14538 79 14572 96
rect 14575 79 14609 96
rect 14095 62 14170 79
rect 14128 61 14170 62
rect 14534 62 14609 79
rect 14534 61 14576 62
rect 14106 55 14192 61
rect 14512 55 14598 61
rect 14640 55 14644 233
rect 14828 183 14832 251
rect 14837 207 14847 241
rect 14857 213 14877 241
rect 14857 207 14871 213
rect 14896 207 14907 251
rect 14938 246 15014 253
rect 15047 251 15056 279
rect 14959 228 14993 246
rect 15001 228 15003 246
rect 14938 221 15014 228
rect 15001 213 15003 221
rect 15045 213 15056 251
rect 15120 241 15124 395
rect 15127 378 15132 412
rect 15156 378 15161 412
rect 15162 400 15173 412
rect 15376 395 15418 421
rect 15782 395 15824 421
rect 16039 420 16051 424
rect 16061 420 16073 424
rect 16111 420 16123 424
rect 16133 421 16145 424
rect 16303 421 16315 424
rect 16133 420 16186 421
rect 16144 412 16186 420
rect 16027 400 16038 412
rect 15308 341 15312 395
rect 15368 387 15414 395
rect 15368 383 15384 387
rect 15376 380 15384 383
rect 15410 380 15414 387
rect 15418 383 15426 395
rect 15774 383 15782 395
rect 15786 387 15820 395
rect 15786 380 15790 387
rect 15816 380 15820 387
rect 15824 383 15832 395
rect 15364 379 15430 380
rect 15770 379 15836 380
rect 15376 371 15380 379
rect 15430 365 15480 367
rect 15720 365 15770 367
rect 15470 361 15524 365
rect 15676 361 15730 365
rect 15470 356 15490 361
rect 15710 356 15730 361
rect 15480 341 15482 356
rect 15308 261 15312 329
rect 15376 305 15380 341
rect 15474 331 15482 341
rect 15490 331 15491 351
rect 15480 315 15482 331
rect 15501 322 15504 356
rect 15523 331 15524 351
rect 15533 331 15540 341
rect 15660 331 15667 341
rect 15676 331 15677 351
rect 15696 322 15699 356
rect 15709 331 15710 351
rect 15719 331 15726 341
rect 15490 315 15506 321
rect 15508 315 15524 321
rect 15676 315 15692 321
rect 15694 315 15710 321
rect 15770 315 15772 365
rect 15313 267 15349 295
rect 15313 261 15327 267
rect 14992 212 15003 213
rect 14837 183 14844 207
rect 14992 183 15002 212
rect 15083 207 15095 241
rect 15105 207 15125 241
rect 14828 103 14832 171
rect 14896 133 14900 183
rect 14896 98 14900 103
rect 14647 62 14652 96
rect 14676 62 14681 96
rect 14896 94 14934 98
rect 14896 79 14904 94
rect 14930 79 14934 94
rect 15018 94 15052 98
rect 15018 79 15022 94
rect 15048 79 15052 94
rect 14896 61 14938 79
rect 15014 61 15056 79
rect 14874 55 14960 61
rect 14992 55 15078 61
rect 15120 55 15124 207
rect 15150 183 15157 211
rect 15308 183 15312 251
rect 15317 233 15327 261
rect 15337 261 15351 267
rect 15376 261 15387 305
rect 15813 267 15824 305
rect 15851 267 15887 295
rect 15888 267 15892 395
rect 16039 378 16044 412
rect 16068 378 16073 412
rect 16074 400 16085 412
rect 16099 400 16110 412
rect 16111 395 16186 412
rect 16262 420 16315 421
rect 16325 420 16337 424
rect 16375 420 16387 424
rect 16397 420 16409 424
rect 16262 412 16304 420
rect 16262 395 16337 412
rect 16338 400 16349 412
rect 16363 400 16374 412
rect 16076 341 16080 395
rect 16111 378 16182 395
rect 16186 383 16194 395
rect 16254 383 16262 395
rect 16266 378 16300 395
rect 16303 378 16337 395
rect 16144 371 16148 378
rect 15538 262 15588 264
rect 15612 262 15662 264
rect 15337 233 15357 261
rect 15376 233 15385 261
rect 15439 253 15473 261
rect 15418 246 15473 253
rect 15439 245 15473 246
rect 15541 253 15572 261
rect 15541 245 15575 253
rect 15376 213 15380 233
rect 15572 229 15575 245
rect 15439 228 15473 229
rect 15418 221 15473 228
rect 15541 221 15575 229
rect 15588 212 15590 262
rect 15628 253 15659 261
rect 15662 253 15664 262
rect 15851 261 15863 267
rect 15628 245 15664 253
rect 15727 253 15761 261
rect 15727 246 15782 253
rect 15727 245 15761 246
rect 15659 229 15664 245
rect 15853 233 15863 261
rect 15873 233 15893 267
rect 16076 261 16080 329
rect 16144 291 16148 341
rect 16144 251 16153 279
rect 16240 264 16250 291
rect 16199 262 16250 264
rect 16240 261 16251 262
rect 16207 253 16241 261
rect 16249 253 16251 261
rect 15628 221 15664 229
rect 15727 228 15761 229
rect 15727 221 15782 228
rect 15662 212 15664 221
rect 15308 103 15312 171
rect 15376 133 15380 183
rect 15430 159 15480 161
rect 15720 159 15770 161
rect 15480 143 15482 159
rect 15490 153 15506 159
rect 15508 153 15524 159
rect 15676 153 15692 159
rect 15694 153 15710 159
rect 15501 143 15524 152
rect 15676 143 15699 152
rect 15474 133 15482 143
rect 15480 109 15482 133
rect 15490 123 15491 143
rect 15501 118 15504 143
rect 15523 123 15524 143
rect 15533 133 15540 143
rect 15660 133 15667 143
rect 15676 123 15677 143
rect 15696 118 15699 143
rect 15709 123 15710 143
rect 15719 133 15726 143
rect 15490 109 15524 113
rect 15676 109 15710 113
rect 15770 109 15772 159
rect 15376 103 15418 104
rect 15782 103 15824 104
rect 15376 96 15380 103
rect 15271 62 15276 96
rect 15300 62 15305 96
rect 15343 79 15414 96
rect 15786 79 15820 96
rect 15823 79 15857 96
rect 15343 62 15418 79
rect 15376 61 15418 62
rect 15782 62 15857 79
rect 15782 61 15824 62
rect 15354 55 15440 61
rect 15760 55 15846 61
rect 15888 55 15892 233
rect 16076 183 16080 251
rect 16085 207 16095 241
rect 16105 213 16125 241
rect 16105 207 16119 213
rect 16144 207 16155 251
rect 16186 246 16262 253
rect 16295 251 16304 279
rect 16207 228 16241 246
rect 16249 228 16251 246
rect 16186 221 16262 228
rect 16249 213 16251 221
rect 16293 213 16304 251
rect 16368 241 16372 395
rect 16375 378 16380 412
rect 16404 378 16409 412
rect 16410 400 16421 412
rect 16624 395 16666 421
rect 17030 395 17072 421
rect 17287 420 17299 424
rect 17309 420 17321 424
rect 17359 420 17371 424
rect 17381 421 17393 424
rect 17551 421 17563 424
rect 17381 420 17434 421
rect 17392 412 17434 420
rect 17275 400 17286 412
rect 16556 341 16560 395
rect 16616 387 16662 395
rect 16616 383 16632 387
rect 16624 380 16632 383
rect 16658 380 16662 387
rect 16666 383 16674 395
rect 17022 383 17030 395
rect 17034 387 17068 395
rect 17034 380 17038 387
rect 17064 380 17068 387
rect 17072 383 17080 395
rect 16612 379 16678 380
rect 17018 379 17084 380
rect 16624 371 16628 379
rect 16678 365 16728 367
rect 16968 365 17018 367
rect 16718 361 16772 365
rect 16924 361 16978 365
rect 16718 356 16738 361
rect 16958 356 16978 361
rect 16728 341 16730 356
rect 16556 261 16560 329
rect 16624 305 16628 341
rect 16722 331 16730 341
rect 16738 331 16739 351
rect 16728 315 16730 331
rect 16749 322 16752 356
rect 16771 331 16772 351
rect 16781 331 16788 341
rect 16908 331 16915 341
rect 16924 331 16925 351
rect 16944 322 16947 356
rect 16957 331 16958 351
rect 16967 331 16974 341
rect 16738 315 16754 321
rect 16756 315 16772 321
rect 16924 315 16940 321
rect 16942 315 16958 321
rect 17018 315 17020 365
rect 16561 267 16597 295
rect 16561 261 16575 267
rect 16240 212 16251 213
rect 16085 183 16092 207
rect 16240 183 16250 212
rect 16331 207 16343 241
rect 16353 207 16373 241
rect 16076 103 16080 171
rect 16144 133 16148 183
rect 16144 98 16148 103
rect 15895 62 15900 96
rect 15924 62 15929 96
rect 16144 94 16182 98
rect 16144 79 16152 94
rect 16178 79 16182 94
rect 16266 94 16300 98
rect 16266 79 16270 94
rect 16296 79 16300 94
rect 16144 61 16186 79
rect 16262 61 16304 79
rect 16122 55 16208 61
rect 16240 55 16326 61
rect 16368 55 16372 207
rect 16398 183 16405 211
rect 16556 183 16560 251
rect 16565 233 16575 261
rect 16585 261 16599 267
rect 16624 261 16635 305
rect 17061 267 17072 305
rect 17099 267 17135 295
rect 17136 267 17140 395
rect 17287 378 17292 412
rect 17316 378 17321 412
rect 17322 400 17333 412
rect 17347 400 17358 412
rect 17359 395 17434 412
rect 17510 420 17563 421
rect 17573 420 17585 424
rect 17623 420 17635 424
rect 17645 420 17657 424
rect 17510 412 17552 420
rect 17510 395 17585 412
rect 17586 400 17597 412
rect 17611 400 17622 412
rect 17324 341 17328 395
rect 17359 378 17430 395
rect 17434 383 17442 395
rect 17502 383 17510 395
rect 17514 378 17548 395
rect 17551 378 17585 395
rect 17392 371 17396 378
rect 16786 262 16836 264
rect 16860 262 16910 264
rect 16585 233 16605 261
rect 16624 233 16633 261
rect 16687 253 16721 261
rect 16666 246 16721 253
rect 16687 245 16721 246
rect 16789 253 16820 261
rect 16789 245 16823 253
rect 16624 213 16628 233
rect 16820 229 16823 245
rect 16687 228 16721 229
rect 16666 221 16721 228
rect 16789 221 16823 229
rect 16836 212 16838 262
rect 16876 253 16907 261
rect 16910 253 16912 262
rect 17099 261 17111 267
rect 16876 245 16912 253
rect 16975 253 17009 261
rect 16975 246 17030 253
rect 16975 245 17009 246
rect 16907 229 16912 245
rect 17101 233 17111 261
rect 17121 233 17141 267
rect 17324 261 17328 329
rect 17392 291 17396 341
rect 17392 251 17401 279
rect 17488 264 17498 291
rect 17447 262 17498 264
rect 17488 261 17499 262
rect 17455 253 17489 261
rect 17497 253 17499 261
rect 16876 221 16912 229
rect 16975 228 17009 229
rect 16975 221 17030 228
rect 16910 212 16912 221
rect 16556 103 16560 171
rect 16624 133 16628 183
rect 16678 159 16728 161
rect 16968 159 17018 161
rect 16728 143 16730 159
rect 16738 153 16754 159
rect 16756 153 16772 159
rect 16924 153 16940 159
rect 16942 153 16958 159
rect 16749 143 16772 152
rect 16924 143 16947 152
rect 16722 133 16730 143
rect 16728 109 16730 133
rect 16738 123 16739 143
rect 16749 118 16752 143
rect 16771 123 16772 143
rect 16781 133 16788 143
rect 16908 133 16915 143
rect 16924 123 16925 143
rect 16944 118 16947 143
rect 16957 123 16958 143
rect 16967 133 16974 143
rect 16738 109 16772 113
rect 16924 109 16958 113
rect 17018 109 17020 159
rect 16624 103 16666 104
rect 17030 103 17072 104
rect 16624 96 16628 103
rect 16519 62 16524 96
rect 16548 62 16553 96
rect 16591 79 16662 96
rect 17034 79 17068 96
rect 17071 79 17105 96
rect 16591 62 16666 79
rect 16624 61 16666 62
rect 17030 62 17105 79
rect 17030 61 17072 62
rect 16602 55 16688 61
rect 17008 55 17094 61
rect 17136 55 17140 233
rect 17324 183 17328 251
rect 17333 207 17343 241
rect 17353 213 17373 241
rect 17353 207 17367 213
rect 17392 207 17403 251
rect 17434 246 17510 253
rect 17543 251 17552 279
rect 17455 228 17489 246
rect 17497 228 17499 246
rect 17434 221 17510 228
rect 17497 213 17499 221
rect 17541 213 17552 251
rect 17616 241 17620 395
rect 17623 378 17628 412
rect 17652 378 17657 412
rect 17658 400 17669 412
rect 17872 395 17914 421
rect 18278 395 18320 421
rect 18535 420 18547 424
rect 18557 420 18569 424
rect 18607 420 18619 424
rect 18629 421 18641 424
rect 18799 421 18811 424
rect 18629 420 18682 421
rect 18640 412 18682 420
rect 18523 400 18534 412
rect 17804 341 17808 395
rect 17864 387 17910 395
rect 17864 383 17880 387
rect 17872 380 17880 383
rect 17906 380 17910 387
rect 17914 383 17922 395
rect 18270 383 18278 395
rect 18282 387 18316 395
rect 18282 380 18286 387
rect 18312 380 18316 387
rect 18320 383 18328 395
rect 17860 379 17926 380
rect 18266 379 18332 380
rect 17872 371 17876 379
rect 17926 365 17976 367
rect 18216 365 18266 367
rect 17966 361 18020 365
rect 18172 361 18226 365
rect 17966 356 17986 361
rect 18206 356 18226 361
rect 17976 341 17978 356
rect 17804 261 17808 329
rect 17872 305 17876 341
rect 17970 331 17978 341
rect 17986 331 17987 351
rect 17976 315 17978 331
rect 17997 322 18000 356
rect 18019 331 18020 351
rect 18029 331 18036 341
rect 18156 331 18163 341
rect 18172 331 18173 351
rect 18192 322 18195 356
rect 18205 331 18206 351
rect 18215 331 18222 341
rect 17986 315 18002 321
rect 18004 315 18020 321
rect 18172 315 18188 321
rect 18190 315 18206 321
rect 18266 315 18268 365
rect 17809 267 17845 295
rect 17809 261 17823 267
rect 17488 212 17499 213
rect 17333 183 17340 207
rect 17488 183 17498 212
rect 17579 207 17591 241
rect 17601 207 17621 241
rect 17324 103 17328 171
rect 17392 133 17396 183
rect 17392 98 17396 103
rect 17143 62 17148 96
rect 17172 62 17177 96
rect 17392 94 17430 98
rect 17392 79 17400 94
rect 17426 79 17430 94
rect 17514 94 17548 98
rect 17514 79 17518 94
rect 17544 79 17548 94
rect 17392 61 17434 79
rect 17510 61 17552 79
rect 17370 55 17456 61
rect 17488 55 17574 61
rect 17616 55 17620 207
rect 17646 183 17653 211
rect 17804 183 17808 251
rect 17813 233 17823 261
rect 17833 261 17847 267
rect 17872 261 17883 305
rect 18309 267 18320 305
rect 18347 267 18383 295
rect 18384 267 18388 395
rect 18535 378 18540 412
rect 18564 378 18569 412
rect 18570 400 18581 412
rect 18595 400 18606 412
rect 18607 395 18682 412
rect 18758 420 18811 421
rect 18821 420 18833 424
rect 18871 420 18883 424
rect 18893 420 18905 424
rect 18758 412 18800 420
rect 18758 395 18833 412
rect 18834 400 18845 412
rect 18859 400 18870 412
rect 18572 341 18576 395
rect 18607 378 18678 395
rect 18682 383 18690 395
rect 18750 383 18758 395
rect 18762 378 18796 395
rect 18799 378 18833 395
rect 18640 371 18644 378
rect 18034 262 18084 264
rect 18108 262 18158 264
rect 17833 233 17853 261
rect 17872 233 17881 261
rect 17935 253 17969 261
rect 17914 246 17969 253
rect 17935 245 17969 246
rect 18037 253 18068 261
rect 18037 245 18071 253
rect 17872 213 17876 233
rect 18068 229 18071 245
rect 17935 228 17969 229
rect 17914 221 17969 228
rect 18037 221 18071 229
rect 18084 212 18086 262
rect 18124 253 18155 261
rect 18158 253 18160 262
rect 18347 261 18359 267
rect 18124 245 18160 253
rect 18223 253 18257 261
rect 18223 246 18278 253
rect 18223 245 18257 246
rect 18155 229 18160 245
rect 18349 233 18359 261
rect 18369 233 18389 267
rect 18572 261 18576 329
rect 18640 291 18644 341
rect 18640 251 18649 279
rect 18736 264 18746 291
rect 18695 262 18746 264
rect 18736 261 18747 262
rect 18703 253 18737 261
rect 18745 253 18747 261
rect 18124 221 18160 229
rect 18223 228 18257 229
rect 18223 221 18278 228
rect 18158 212 18160 221
rect 17804 103 17808 171
rect 17872 133 17876 183
rect 17926 159 17976 161
rect 18216 159 18266 161
rect 17976 143 17978 159
rect 17986 153 18002 159
rect 18004 153 18020 159
rect 18172 153 18188 159
rect 18190 153 18206 159
rect 17997 143 18020 152
rect 18172 143 18195 152
rect 17970 133 17978 143
rect 17976 109 17978 133
rect 17986 123 17987 143
rect 17997 118 18000 143
rect 18019 123 18020 143
rect 18029 133 18036 143
rect 18156 133 18163 143
rect 18172 123 18173 143
rect 18192 118 18195 143
rect 18205 123 18206 143
rect 18215 133 18222 143
rect 17986 109 18020 113
rect 18172 109 18206 113
rect 18266 109 18268 159
rect 17872 103 17914 104
rect 18278 103 18320 104
rect 17872 96 17876 103
rect 17767 62 17772 96
rect 17796 62 17801 96
rect 17839 79 17910 96
rect 18282 79 18316 96
rect 18319 79 18353 96
rect 17839 62 17914 79
rect 17872 61 17914 62
rect 18278 62 18353 79
rect 18278 61 18320 62
rect 17850 55 17936 61
rect 18256 55 18342 61
rect 18384 55 18388 233
rect 18572 183 18576 251
rect 18581 207 18591 241
rect 18601 213 18621 241
rect 18601 207 18615 213
rect 18640 207 18651 251
rect 18682 246 18758 253
rect 18791 251 18800 279
rect 18703 228 18737 246
rect 18745 228 18747 246
rect 18682 221 18758 228
rect 18745 213 18747 221
rect 18789 213 18800 251
rect 18864 241 18868 395
rect 18871 378 18876 412
rect 18900 378 18905 412
rect 18906 400 18917 412
rect 19120 395 19162 421
rect 19526 395 19568 421
rect 19783 420 19795 424
rect 19805 420 19817 424
rect 19855 420 19867 424
rect 19877 421 19889 424
rect 20047 421 20059 424
rect 19877 420 19930 421
rect 19888 412 19930 420
rect 19771 400 19782 412
rect 19052 341 19056 395
rect 19112 387 19158 395
rect 19112 383 19128 387
rect 19120 380 19128 383
rect 19154 380 19158 387
rect 19162 383 19170 395
rect 19518 383 19526 395
rect 19530 387 19564 395
rect 19530 380 19534 387
rect 19560 380 19564 387
rect 19568 383 19576 395
rect 19108 379 19174 380
rect 19514 379 19580 380
rect 19120 371 19124 379
rect 19174 365 19224 367
rect 19464 365 19514 367
rect 19214 361 19268 365
rect 19420 361 19474 365
rect 19214 356 19234 361
rect 19454 356 19474 361
rect 19224 341 19226 356
rect 19052 261 19056 329
rect 19120 305 19124 341
rect 19218 331 19226 341
rect 19234 331 19235 351
rect 19224 315 19226 331
rect 19245 322 19248 356
rect 19267 331 19268 351
rect 19277 331 19284 341
rect 19404 331 19411 341
rect 19420 331 19421 351
rect 19440 322 19443 356
rect 19453 331 19454 351
rect 19463 331 19470 341
rect 19234 315 19250 321
rect 19252 315 19268 321
rect 19420 315 19436 321
rect 19438 315 19454 321
rect 19514 315 19516 365
rect 19057 267 19093 295
rect 19057 261 19071 267
rect 18736 212 18747 213
rect 18581 183 18588 207
rect 18736 183 18746 212
rect 18827 207 18839 241
rect 18849 207 18869 241
rect 18572 103 18576 171
rect 18640 133 18644 183
rect 18640 98 18644 103
rect 18391 62 18396 96
rect 18420 62 18425 96
rect 18640 94 18678 98
rect 18640 79 18648 94
rect 18674 79 18678 94
rect 18762 94 18796 98
rect 18762 79 18766 94
rect 18792 79 18796 94
rect 18640 61 18682 79
rect 18758 61 18800 79
rect 18618 55 18704 61
rect 18736 55 18822 61
rect 18864 55 18868 207
rect 18894 183 18901 211
rect 19052 183 19056 251
rect 19061 233 19071 261
rect 19081 261 19095 267
rect 19120 261 19131 305
rect 19557 267 19568 305
rect 19595 267 19631 295
rect 19632 267 19636 395
rect 19783 378 19788 412
rect 19812 378 19817 412
rect 19818 400 19829 412
rect 19843 400 19854 412
rect 19855 395 19930 412
rect 20006 420 20059 421
rect 20069 420 20081 424
rect 20119 420 20131 424
rect 20141 420 20153 424
rect 20006 412 20048 420
rect 20006 395 20081 412
rect 20082 400 20093 412
rect 20107 400 20118 412
rect 19820 341 19824 395
rect 19855 378 19926 395
rect 19930 383 19938 395
rect 19998 383 20006 395
rect 20010 378 20044 395
rect 20047 378 20081 395
rect 19888 371 19892 378
rect 19282 262 19332 264
rect 19356 262 19406 264
rect 19081 233 19101 261
rect 19120 233 19129 261
rect 19183 253 19217 261
rect 19162 246 19217 253
rect 19183 245 19217 246
rect 19285 253 19316 261
rect 19285 245 19319 253
rect 19120 213 19124 233
rect 19316 229 19319 245
rect 19183 228 19217 229
rect 19162 221 19217 228
rect 19285 221 19319 229
rect 19332 212 19334 262
rect 19372 253 19403 261
rect 19406 253 19408 262
rect 19595 261 19607 267
rect 19372 245 19408 253
rect 19471 253 19505 261
rect 19471 246 19526 253
rect 19471 245 19505 246
rect 19403 229 19408 245
rect 19597 233 19607 261
rect 19617 233 19637 267
rect 19820 261 19824 329
rect 19888 291 19892 341
rect 19888 251 19897 279
rect 19984 264 19994 291
rect 19943 262 19994 264
rect 19984 261 19995 262
rect 19951 253 19985 261
rect 19993 253 19995 261
rect 19372 221 19408 229
rect 19471 228 19505 229
rect 19471 221 19526 228
rect 19406 212 19408 221
rect 19052 103 19056 171
rect 19120 133 19124 183
rect 19174 159 19224 161
rect 19464 159 19514 161
rect 19224 143 19226 159
rect 19234 153 19250 159
rect 19252 153 19268 159
rect 19420 153 19436 159
rect 19438 153 19454 159
rect 19245 143 19268 152
rect 19420 143 19443 152
rect 19218 133 19226 143
rect 19224 109 19226 133
rect 19234 123 19235 143
rect 19245 118 19248 143
rect 19267 123 19268 143
rect 19277 133 19284 143
rect 19404 133 19411 143
rect 19420 123 19421 143
rect 19440 118 19443 143
rect 19453 123 19454 143
rect 19463 133 19470 143
rect 19234 109 19268 113
rect 19420 109 19454 113
rect 19514 109 19516 159
rect 19120 103 19162 104
rect 19526 103 19568 104
rect 19120 96 19124 103
rect 19015 62 19020 96
rect 19044 62 19049 96
rect 19087 79 19158 96
rect 19530 79 19564 96
rect 19567 79 19601 96
rect 19087 62 19162 79
rect 19120 61 19162 62
rect 19526 62 19601 79
rect 19526 61 19568 62
rect 19098 55 19184 61
rect 19504 55 19590 61
rect 19632 55 19636 233
rect 19820 183 19824 251
rect 19829 207 19839 241
rect 19849 213 19869 241
rect 19849 207 19863 213
rect 19888 207 19899 251
rect 19930 246 20006 253
rect 20039 251 20048 279
rect 19951 228 19985 246
rect 19993 228 19995 246
rect 19930 221 20006 228
rect 19993 213 19995 221
rect 20037 213 20048 251
rect 20112 241 20116 395
rect 20119 378 20124 412
rect 20148 378 20153 412
rect 20154 400 20165 412
rect 20368 395 20410 421
rect 20774 395 20816 421
rect 21031 420 21043 424
rect 21053 420 21065 424
rect 21103 420 21115 424
rect 21125 421 21137 424
rect 21295 421 21307 424
rect 21125 420 21178 421
rect 21136 412 21178 420
rect 21019 400 21030 412
rect 20300 341 20304 395
rect 20360 387 20406 395
rect 20360 383 20376 387
rect 20368 380 20376 383
rect 20402 380 20406 387
rect 20410 383 20418 395
rect 20766 383 20774 395
rect 20778 387 20812 395
rect 20778 380 20782 387
rect 20808 380 20812 387
rect 20816 383 20824 395
rect 20356 379 20422 380
rect 20762 379 20828 380
rect 20368 371 20372 379
rect 20422 365 20472 367
rect 20712 365 20762 367
rect 20462 361 20516 365
rect 20668 361 20722 365
rect 20462 356 20482 361
rect 20702 356 20722 361
rect 20472 341 20474 356
rect 20300 261 20304 329
rect 20368 305 20372 341
rect 20466 331 20474 341
rect 20482 331 20483 351
rect 20472 315 20474 331
rect 20493 322 20496 356
rect 20515 331 20516 351
rect 20525 331 20532 341
rect 20652 331 20659 341
rect 20668 331 20669 351
rect 20688 322 20691 356
rect 20701 331 20702 351
rect 20711 331 20718 341
rect 20482 315 20498 321
rect 20500 315 20516 321
rect 20668 315 20684 321
rect 20686 315 20702 321
rect 20762 315 20764 365
rect 20305 267 20341 295
rect 20305 261 20319 267
rect 19984 212 19995 213
rect 19829 183 19836 207
rect 19984 183 19994 212
rect 20075 207 20087 241
rect 20097 207 20117 241
rect 19820 103 19824 171
rect 19888 133 19892 183
rect 19888 98 19892 103
rect 19639 62 19644 96
rect 19668 62 19673 96
rect 19888 94 19926 98
rect 19888 79 19896 94
rect 19922 79 19926 94
rect 20010 94 20044 98
rect 20010 79 20014 94
rect 20040 79 20044 94
rect 19888 61 19930 79
rect 20006 61 20048 79
rect 19866 55 19952 61
rect 19984 55 20070 61
rect 20112 55 20116 207
rect 20142 183 20149 211
rect 20300 183 20304 251
rect 20309 233 20319 261
rect 20329 261 20343 267
rect 20368 261 20379 305
rect 20805 267 20816 305
rect 20843 267 20879 295
rect 20880 267 20884 395
rect 21031 378 21036 412
rect 21060 378 21065 412
rect 21066 400 21077 412
rect 21091 400 21102 412
rect 21103 395 21178 412
rect 21254 420 21307 421
rect 21317 420 21329 424
rect 21367 420 21379 424
rect 21389 420 21401 424
rect 21254 412 21296 420
rect 21254 395 21329 412
rect 21330 400 21341 412
rect 21355 400 21366 412
rect 21068 341 21072 395
rect 21103 378 21174 395
rect 21178 383 21186 395
rect 21246 383 21254 395
rect 21258 378 21292 395
rect 21295 378 21329 395
rect 21136 371 21140 378
rect 20530 262 20580 264
rect 20604 262 20654 264
rect 20329 233 20349 261
rect 20368 233 20377 261
rect 20431 253 20465 261
rect 20410 246 20465 253
rect 20431 245 20465 246
rect 20533 253 20564 261
rect 20533 245 20567 253
rect 20368 213 20372 233
rect 20564 229 20567 245
rect 20431 228 20465 229
rect 20410 221 20465 228
rect 20533 221 20567 229
rect 20580 212 20582 262
rect 20620 253 20651 261
rect 20654 253 20656 262
rect 20843 261 20855 267
rect 20620 245 20656 253
rect 20719 253 20753 261
rect 20719 246 20774 253
rect 20719 245 20753 246
rect 20651 229 20656 245
rect 20845 233 20855 261
rect 20865 233 20885 267
rect 21068 261 21072 329
rect 21136 291 21140 341
rect 21136 251 21145 279
rect 21232 264 21242 291
rect 21191 262 21242 264
rect 21232 261 21243 262
rect 21199 253 21233 261
rect 21241 253 21243 261
rect 20620 221 20656 229
rect 20719 228 20753 229
rect 20719 221 20774 228
rect 20654 212 20656 221
rect 20300 103 20304 171
rect 20368 133 20372 183
rect 20422 159 20472 161
rect 20712 159 20762 161
rect 20472 143 20474 159
rect 20482 153 20498 159
rect 20500 153 20516 159
rect 20668 153 20684 159
rect 20686 153 20702 159
rect 20493 143 20516 152
rect 20668 143 20691 152
rect 20466 133 20474 143
rect 20472 109 20474 133
rect 20482 123 20483 143
rect 20493 118 20496 143
rect 20515 123 20516 143
rect 20525 133 20532 143
rect 20652 133 20659 143
rect 20668 123 20669 143
rect 20688 118 20691 143
rect 20701 123 20702 143
rect 20711 133 20718 143
rect 20482 109 20516 113
rect 20668 109 20702 113
rect 20762 109 20764 159
rect 20368 103 20410 104
rect 20774 103 20816 104
rect 20368 96 20372 103
rect 20263 62 20268 96
rect 20292 62 20297 96
rect 20335 79 20406 96
rect 20778 79 20812 96
rect 20815 79 20849 96
rect 20335 62 20410 79
rect 20368 61 20410 62
rect 20774 62 20849 79
rect 20774 61 20816 62
rect 20346 55 20432 61
rect 20752 55 20838 61
rect 20880 55 20884 233
rect 21068 183 21072 251
rect 21077 207 21087 241
rect 21097 213 21117 241
rect 21097 207 21111 213
rect 21136 207 21147 251
rect 21178 246 21254 253
rect 21287 251 21296 279
rect 21199 228 21233 246
rect 21241 228 21243 246
rect 21178 221 21254 228
rect 21241 213 21243 221
rect 21285 213 21296 251
rect 21360 241 21364 395
rect 21367 378 21372 412
rect 21396 378 21401 412
rect 21402 400 21413 412
rect 21616 395 21658 421
rect 22022 395 22064 421
rect 22279 420 22291 424
rect 22301 420 22313 424
rect 22351 420 22363 424
rect 22373 421 22385 424
rect 22543 421 22555 424
rect 22373 420 22426 421
rect 22384 412 22426 420
rect 22267 400 22278 412
rect 21548 341 21552 395
rect 21608 387 21654 395
rect 21608 383 21624 387
rect 21616 380 21624 383
rect 21650 380 21654 387
rect 21658 383 21666 395
rect 22014 383 22022 395
rect 22026 387 22060 395
rect 22026 380 22030 387
rect 22056 380 22060 387
rect 22064 383 22072 395
rect 21604 379 21670 380
rect 22010 379 22076 380
rect 21616 371 21620 379
rect 21670 365 21720 367
rect 21960 365 22010 367
rect 21710 361 21764 365
rect 21916 361 21970 365
rect 21710 356 21730 361
rect 21950 356 21970 361
rect 21720 341 21722 356
rect 21548 261 21552 329
rect 21616 305 21620 341
rect 21714 331 21722 341
rect 21730 331 21731 351
rect 21720 315 21722 331
rect 21741 322 21744 356
rect 21763 331 21764 351
rect 21773 331 21780 341
rect 21900 331 21907 341
rect 21916 331 21917 351
rect 21936 322 21939 356
rect 21949 331 21950 351
rect 21959 331 21966 341
rect 21730 315 21746 321
rect 21748 315 21764 321
rect 21916 315 21932 321
rect 21934 315 21950 321
rect 22010 315 22012 365
rect 21553 267 21589 295
rect 21553 261 21567 267
rect 21232 212 21243 213
rect 21077 183 21084 207
rect 21232 183 21242 212
rect 21323 207 21335 241
rect 21345 207 21365 241
rect 21068 103 21072 171
rect 21136 133 21140 183
rect 21136 98 21140 103
rect 20887 62 20892 96
rect 20916 62 20921 96
rect 21136 94 21174 98
rect 21136 79 21144 94
rect 21170 79 21174 94
rect 21258 94 21292 98
rect 21258 79 21262 94
rect 21288 79 21292 94
rect 21136 61 21178 79
rect 21254 61 21296 79
rect 21114 55 21200 61
rect 21232 55 21318 61
rect 21360 55 21364 207
rect 21390 183 21397 211
rect 21548 183 21552 251
rect 21557 233 21567 261
rect 21577 261 21591 267
rect 21616 261 21627 305
rect 22053 267 22064 305
rect 22091 267 22127 295
rect 22128 267 22132 395
rect 22279 378 22284 412
rect 22308 378 22313 412
rect 22314 400 22325 412
rect 22339 400 22350 412
rect 22351 395 22426 412
rect 22502 420 22555 421
rect 22565 420 22577 424
rect 22615 420 22627 424
rect 22637 420 22649 424
rect 22502 412 22544 420
rect 22502 395 22577 412
rect 22578 400 22589 412
rect 22603 400 22614 412
rect 22316 341 22320 395
rect 22351 378 22422 395
rect 22426 383 22434 395
rect 22494 383 22502 395
rect 22506 378 22540 395
rect 22543 378 22577 395
rect 22384 371 22388 378
rect 21778 262 21828 264
rect 21852 262 21902 264
rect 21577 233 21597 261
rect 21616 233 21625 261
rect 21679 253 21713 261
rect 21658 246 21713 253
rect 21679 245 21713 246
rect 21781 253 21812 261
rect 21781 245 21815 253
rect 21616 213 21620 233
rect 21812 229 21815 245
rect 21679 228 21713 229
rect 21658 221 21713 228
rect 21781 221 21815 229
rect 21828 212 21830 262
rect 21868 253 21899 261
rect 21902 253 21904 262
rect 22091 261 22103 267
rect 21868 245 21904 253
rect 21967 253 22001 261
rect 21967 246 22022 253
rect 21967 245 22001 246
rect 21899 229 21904 245
rect 22093 233 22103 261
rect 22113 233 22133 267
rect 22316 261 22320 329
rect 22384 291 22388 341
rect 22384 251 22393 279
rect 22480 264 22490 291
rect 22439 262 22490 264
rect 22480 261 22491 262
rect 22447 253 22481 261
rect 22489 253 22491 261
rect 21868 221 21904 229
rect 21967 228 22001 229
rect 21967 221 22022 228
rect 21902 212 21904 221
rect 21548 103 21552 171
rect 21616 133 21620 183
rect 21670 159 21720 161
rect 21960 159 22010 161
rect 21720 143 21722 159
rect 21730 153 21746 159
rect 21748 153 21764 159
rect 21916 153 21932 159
rect 21934 153 21950 159
rect 21741 143 21764 152
rect 21916 143 21939 152
rect 21714 133 21722 143
rect 21720 109 21722 133
rect 21730 123 21731 143
rect 21741 118 21744 143
rect 21763 123 21764 143
rect 21773 133 21780 143
rect 21900 133 21907 143
rect 21916 123 21917 143
rect 21936 118 21939 143
rect 21949 123 21950 143
rect 21959 133 21966 143
rect 21730 109 21764 113
rect 21916 109 21950 113
rect 22010 109 22012 159
rect 21616 103 21658 104
rect 22022 103 22064 104
rect 21616 96 21620 103
rect 21511 62 21516 96
rect 21540 62 21545 96
rect 21583 79 21654 96
rect 22026 79 22060 96
rect 22063 79 22097 96
rect 21583 62 21658 79
rect 21616 61 21658 62
rect 22022 62 22097 79
rect 22022 61 22064 62
rect 21594 55 21680 61
rect 22000 55 22086 61
rect 22128 55 22132 233
rect 22316 183 22320 251
rect 22325 207 22335 241
rect 22345 213 22365 241
rect 22345 207 22359 213
rect 22384 207 22395 251
rect 22426 246 22502 253
rect 22535 251 22544 279
rect 22447 228 22481 246
rect 22489 228 22491 246
rect 22426 221 22502 228
rect 22489 213 22491 221
rect 22533 213 22544 251
rect 22608 241 22612 395
rect 22615 378 22620 412
rect 22644 378 22649 412
rect 22650 400 22661 412
rect 22864 395 22906 421
rect 23270 395 23312 421
rect 23527 420 23539 424
rect 23549 420 23561 424
rect 23599 420 23611 424
rect 23621 421 23633 424
rect 23791 421 23803 424
rect 23621 420 23674 421
rect 23632 412 23674 420
rect 23515 400 23526 412
rect 22796 341 22800 395
rect 22856 387 22902 395
rect 22856 383 22872 387
rect 22864 380 22872 383
rect 22898 380 22902 387
rect 22906 383 22914 395
rect 23262 383 23270 395
rect 23274 387 23308 395
rect 23274 380 23278 387
rect 23304 380 23308 387
rect 23312 383 23320 395
rect 22852 379 22918 380
rect 23258 379 23324 380
rect 22864 371 22868 379
rect 22918 365 22968 367
rect 23208 365 23258 367
rect 22958 361 23012 365
rect 23164 361 23218 365
rect 22958 356 22978 361
rect 23198 356 23218 361
rect 22968 341 22970 356
rect 22796 261 22800 329
rect 22864 305 22868 341
rect 22962 331 22970 341
rect 22978 331 22979 351
rect 22968 315 22970 331
rect 22989 322 22992 356
rect 23011 331 23012 351
rect 23021 331 23028 341
rect 23148 331 23155 341
rect 23164 331 23165 351
rect 23184 322 23187 356
rect 23197 331 23198 351
rect 23207 331 23214 341
rect 22978 315 22994 321
rect 22996 315 23012 321
rect 23164 315 23180 321
rect 23182 315 23198 321
rect 23258 315 23260 365
rect 22801 267 22837 295
rect 22801 261 22815 267
rect 22480 212 22491 213
rect 22325 183 22332 207
rect 22480 183 22490 212
rect 22571 207 22583 241
rect 22593 207 22613 241
rect 22316 103 22320 171
rect 22384 133 22388 183
rect 22384 98 22388 103
rect 22135 62 22140 96
rect 22164 62 22169 96
rect 22384 94 22422 98
rect 22384 79 22392 94
rect 22418 79 22422 94
rect 22506 94 22540 98
rect 22506 79 22510 94
rect 22536 79 22540 94
rect 22384 61 22426 79
rect 22502 61 22544 79
rect 22362 55 22448 61
rect 22480 55 22566 61
rect 22608 55 22612 207
rect 22638 183 22645 211
rect 22796 183 22800 251
rect 22805 233 22815 261
rect 22825 261 22839 267
rect 22864 261 22875 305
rect 23301 267 23312 305
rect 23339 267 23375 295
rect 23376 267 23380 395
rect 23527 378 23532 412
rect 23556 378 23561 412
rect 23562 400 23573 412
rect 23587 400 23598 412
rect 23599 395 23674 412
rect 23750 420 23803 421
rect 23813 420 23825 424
rect 23863 420 23875 424
rect 23885 420 23897 424
rect 23750 412 23792 420
rect 23750 395 23825 412
rect 23826 400 23837 412
rect 23851 400 23862 412
rect 23564 341 23568 395
rect 23599 378 23670 395
rect 23674 383 23682 395
rect 23742 383 23750 395
rect 23754 378 23788 395
rect 23791 378 23825 395
rect 23632 371 23636 378
rect 23026 262 23076 264
rect 23100 262 23150 264
rect 22825 233 22845 261
rect 22864 233 22873 261
rect 22927 253 22961 261
rect 22906 246 22961 253
rect 22927 245 22961 246
rect 23029 253 23060 261
rect 23029 245 23063 253
rect 22864 213 22868 233
rect 23060 229 23063 245
rect 22927 228 22961 229
rect 22906 221 22961 228
rect 23029 221 23063 229
rect 23076 212 23078 262
rect 23116 253 23147 261
rect 23150 253 23152 262
rect 23339 261 23351 267
rect 23116 245 23152 253
rect 23215 253 23249 261
rect 23215 246 23270 253
rect 23215 245 23249 246
rect 23147 229 23152 245
rect 23341 233 23351 261
rect 23361 233 23381 267
rect 23564 261 23568 329
rect 23632 291 23636 341
rect 23632 251 23641 279
rect 23728 264 23738 291
rect 23687 262 23738 264
rect 23728 261 23739 262
rect 23695 253 23729 261
rect 23737 253 23739 261
rect 23116 221 23152 229
rect 23215 228 23249 229
rect 23215 221 23270 228
rect 23150 212 23152 221
rect 22796 103 22800 171
rect 22864 133 22868 183
rect 22918 159 22968 161
rect 23208 159 23258 161
rect 22968 143 22970 159
rect 22978 153 22994 159
rect 22996 153 23012 159
rect 23164 153 23180 159
rect 23182 153 23198 159
rect 22989 143 23012 152
rect 23164 143 23187 152
rect 22962 133 22970 143
rect 22968 109 22970 133
rect 22978 123 22979 143
rect 22989 118 22992 143
rect 23011 123 23012 143
rect 23021 133 23028 143
rect 23148 133 23155 143
rect 23164 123 23165 143
rect 23184 118 23187 143
rect 23197 123 23198 143
rect 23207 133 23214 143
rect 22978 109 23012 113
rect 23164 109 23198 113
rect 23258 109 23260 159
rect 22864 103 22906 104
rect 23270 103 23312 104
rect 22864 96 22868 103
rect 22759 62 22764 96
rect 22788 62 22793 96
rect 22831 79 22902 96
rect 23274 79 23308 96
rect 23311 79 23345 96
rect 22831 62 22906 79
rect 22864 61 22906 62
rect 23270 62 23345 79
rect 23270 61 23312 62
rect 22842 55 22928 61
rect 23248 55 23334 61
rect 23376 55 23380 233
rect 23564 183 23568 251
rect 23573 207 23583 241
rect 23593 213 23613 241
rect 23593 207 23607 213
rect 23632 207 23643 251
rect 23674 246 23750 253
rect 23783 251 23792 279
rect 23695 228 23729 246
rect 23737 228 23739 246
rect 23674 221 23750 228
rect 23737 213 23739 221
rect 23781 213 23792 251
rect 23856 241 23860 395
rect 23863 378 23868 412
rect 23892 378 23897 412
rect 23898 400 23909 412
rect 24112 395 24154 421
rect 24518 395 24560 421
rect 24775 420 24787 424
rect 24797 420 24809 424
rect 24847 420 24859 424
rect 24869 421 24881 424
rect 25039 421 25051 424
rect 24869 420 24922 421
rect 24880 412 24922 420
rect 24763 400 24774 412
rect 24044 341 24048 395
rect 24104 387 24150 395
rect 24104 383 24120 387
rect 24112 380 24120 383
rect 24146 380 24150 387
rect 24154 383 24162 395
rect 24510 383 24518 395
rect 24522 387 24556 395
rect 24522 380 24526 387
rect 24552 380 24556 387
rect 24560 383 24568 395
rect 24100 379 24166 380
rect 24506 379 24572 380
rect 24112 371 24116 379
rect 24166 365 24216 367
rect 24456 365 24506 367
rect 24206 361 24260 365
rect 24412 361 24466 365
rect 24206 356 24226 361
rect 24446 356 24466 361
rect 24216 341 24218 356
rect 24044 261 24048 329
rect 24112 305 24116 341
rect 24210 331 24218 341
rect 24226 331 24227 351
rect 24216 315 24218 331
rect 24237 322 24240 356
rect 24259 331 24260 351
rect 24269 331 24276 341
rect 24396 331 24403 341
rect 24412 331 24413 351
rect 24432 322 24435 356
rect 24445 331 24446 351
rect 24455 331 24462 341
rect 24226 315 24242 321
rect 24244 315 24260 321
rect 24412 315 24428 321
rect 24430 315 24446 321
rect 24506 315 24508 365
rect 24049 267 24085 295
rect 24049 261 24063 267
rect 23728 212 23739 213
rect 23573 183 23580 207
rect 23728 183 23738 212
rect 23819 207 23831 241
rect 23841 207 23861 241
rect 23564 103 23568 171
rect 23632 133 23636 183
rect 23632 98 23636 103
rect 23383 62 23388 96
rect 23412 62 23417 96
rect 23632 94 23670 98
rect 23632 79 23640 94
rect 23666 79 23670 94
rect 23754 94 23788 98
rect 23754 79 23758 94
rect 23784 79 23788 94
rect 23632 61 23674 79
rect 23750 61 23792 79
rect 23610 55 23696 61
rect 23728 55 23814 61
rect 23856 55 23860 207
rect 23886 183 23893 211
rect 24044 183 24048 251
rect 24053 233 24063 261
rect 24073 261 24087 267
rect 24112 261 24123 305
rect 24549 267 24560 305
rect 24587 267 24623 295
rect 24624 267 24628 395
rect 24775 378 24780 412
rect 24804 378 24809 412
rect 24810 400 24821 412
rect 24835 400 24846 412
rect 24847 395 24922 412
rect 24998 420 25051 421
rect 25061 420 25073 424
rect 25111 420 25123 424
rect 25133 420 25145 424
rect 24998 412 25040 420
rect 24998 395 25073 412
rect 25074 400 25085 412
rect 25099 400 25110 412
rect 24812 341 24816 395
rect 24847 378 24918 395
rect 24922 383 24930 395
rect 24990 383 24998 395
rect 25002 378 25036 395
rect 25039 378 25073 395
rect 24880 371 24884 378
rect 24274 262 24324 264
rect 24348 262 24398 264
rect 24073 233 24093 261
rect 24112 233 24121 261
rect 24175 253 24209 261
rect 24154 246 24209 253
rect 24175 245 24209 246
rect 24277 253 24308 261
rect 24277 245 24311 253
rect 24112 213 24116 233
rect 24308 229 24311 245
rect 24175 228 24209 229
rect 24154 221 24209 228
rect 24277 221 24311 229
rect 24324 212 24326 262
rect 24364 253 24395 261
rect 24398 253 24400 262
rect 24587 261 24599 267
rect 24364 245 24400 253
rect 24463 253 24497 261
rect 24463 246 24518 253
rect 24463 245 24497 246
rect 24395 229 24400 245
rect 24589 233 24599 261
rect 24609 233 24629 267
rect 24812 261 24816 329
rect 24880 291 24884 341
rect 24880 251 24889 279
rect 24976 264 24986 291
rect 24935 262 24986 264
rect 24976 261 24987 262
rect 24943 253 24977 261
rect 24985 253 24987 261
rect 24364 221 24400 229
rect 24463 228 24497 229
rect 24463 221 24518 228
rect 24398 212 24400 221
rect 24044 103 24048 171
rect 24112 133 24116 183
rect 24166 159 24216 161
rect 24456 159 24506 161
rect 24216 143 24218 159
rect 24226 153 24242 159
rect 24244 153 24260 159
rect 24412 153 24428 159
rect 24430 153 24446 159
rect 24237 143 24260 152
rect 24412 143 24435 152
rect 24210 133 24218 143
rect 24216 109 24218 133
rect 24226 123 24227 143
rect 24237 118 24240 143
rect 24259 123 24260 143
rect 24269 133 24276 143
rect 24396 133 24403 143
rect 24412 123 24413 143
rect 24432 118 24435 143
rect 24445 123 24446 143
rect 24455 133 24462 143
rect 24226 109 24260 113
rect 24412 109 24446 113
rect 24506 109 24508 159
rect 24112 103 24154 104
rect 24518 103 24560 104
rect 24112 96 24116 103
rect 24007 62 24012 96
rect 24036 62 24041 96
rect 24079 79 24150 96
rect 24522 79 24556 96
rect 24559 79 24593 96
rect 24079 62 24154 79
rect 24112 61 24154 62
rect 24518 62 24593 79
rect 24518 61 24560 62
rect 24090 55 24176 61
rect 24496 55 24582 61
rect 24624 55 24628 233
rect 24812 183 24816 251
rect 24821 207 24831 241
rect 24841 213 24861 241
rect 24841 207 24855 213
rect 24880 207 24891 251
rect 24922 246 24998 253
rect 25031 251 25040 279
rect 24943 228 24977 246
rect 24985 228 24987 246
rect 24922 221 24998 228
rect 24985 213 24987 221
rect 25029 213 25040 251
rect 25104 241 25108 395
rect 25111 378 25116 412
rect 25140 378 25145 412
rect 25146 400 25157 412
rect 25360 395 25402 421
rect 25766 395 25808 421
rect 26023 420 26035 424
rect 26045 420 26057 424
rect 26095 420 26107 424
rect 26117 421 26129 424
rect 26287 421 26299 424
rect 26117 420 26170 421
rect 26128 412 26170 420
rect 26011 400 26022 412
rect 25292 341 25296 395
rect 25352 387 25398 395
rect 25352 383 25368 387
rect 25360 380 25368 383
rect 25394 380 25398 387
rect 25402 383 25410 395
rect 25758 383 25766 395
rect 25770 387 25804 395
rect 25770 380 25774 387
rect 25800 380 25804 387
rect 25808 383 25816 395
rect 25348 379 25414 380
rect 25754 379 25820 380
rect 25360 371 25364 379
rect 25414 365 25464 367
rect 25704 365 25754 367
rect 25454 361 25508 365
rect 25660 361 25714 365
rect 25454 356 25474 361
rect 25694 356 25714 361
rect 25464 341 25466 356
rect 25292 261 25296 329
rect 25360 305 25364 341
rect 25458 331 25466 341
rect 25474 331 25475 351
rect 25464 315 25466 331
rect 25485 322 25488 356
rect 25507 331 25508 351
rect 25517 331 25524 341
rect 25644 331 25651 341
rect 25660 331 25661 351
rect 25680 322 25683 356
rect 25693 331 25694 351
rect 25703 331 25710 341
rect 25474 315 25490 321
rect 25492 315 25508 321
rect 25660 315 25676 321
rect 25678 315 25694 321
rect 25754 315 25756 365
rect 25297 267 25333 295
rect 25297 261 25311 267
rect 24976 212 24987 213
rect 24821 183 24828 207
rect 24976 183 24986 212
rect 25067 207 25079 241
rect 25089 207 25109 241
rect 24812 103 24816 171
rect 24880 133 24884 183
rect 24880 98 24884 103
rect 24631 62 24636 96
rect 24660 62 24665 96
rect 24880 94 24918 98
rect 24880 79 24888 94
rect 24914 79 24918 94
rect 25002 94 25036 98
rect 25002 79 25006 94
rect 25032 79 25036 94
rect 24880 61 24922 79
rect 24998 61 25040 79
rect 24858 55 24944 61
rect 24976 55 25062 61
rect 25104 55 25108 207
rect 25134 183 25141 211
rect 25292 183 25296 251
rect 25301 233 25311 261
rect 25321 261 25335 267
rect 25360 261 25371 305
rect 25797 267 25808 305
rect 25835 267 25871 295
rect 25872 267 25876 395
rect 26023 378 26028 412
rect 26052 378 26057 412
rect 26058 400 26069 412
rect 26083 400 26094 412
rect 26095 395 26170 412
rect 26246 420 26299 421
rect 26309 420 26321 424
rect 26359 420 26371 424
rect 26381 420 26393 424
rect 26246 412 26288 420
rect 26246 395 26321 412
rect 26322 400 26333 412
rect 26347 400 26358 412
rect 26060 341 26064 395
rect 26095 378 26166 395
rect 26170 383 26178 395
rect 26238 383 26246 395
rect 26250 378 26284 395
rect 26287 378 26321 395
rect 26128 371 26132 378
rect 25522 262 25572 264
rect 25596 262 25646 264
rect 25321 233 25341 261
rect 25360 233 25369 261
rect 25423 253 25457 261
rect 25402 246 25457 253
rect 25423 245 25457 246
rect 25525 253 25556 261
rect 25525 245 25559 253
rect 25360 213 25364 233
rect 25556 229 25559 245
rect 25423 228 25457 229
rect 25402 221 25457 228
rect 25525 221 25559 229
rect 25572 212 25574 262
rect 25612 253 25643 261
rect 25646 253 25648 262
rect 25835 261 25847 267
rect 25612 245 25648 253
rect 25711 253 25745 261
rect 25711 246 25766 253
rect 25711 245 25745 246
rect 25643 229 25648 245
rect 25837 233 25847 261
rect 25857 233 25877 267
rect 26060 261 26064 329
rect 26128 291 26132 341
rect 26128 251 26137 279
rect 26224 264 26234 291
rect 26183 262 26234 264
rect 26224 261 26235 262
rect 26191 253 26225 261
rect 26233 253 26235 261
rect 25612 221 25648 229
rect 25711 228 25745 229
rect 25711 221 25766 228
rect 25646 212 25648 221
rect 25292 103 25296 171
rect 25360 133 25364 183
rect 25414 159 25464 161
rect 25704 159 25754 161
rect 25464 143 25466 159
rect 25474 153 25490 159
rect 25492 153 25508 159
rect 25660 153 25676 159
rect 25678 153 25694 159
rect 25485 143 25508 152
rect 25660 143 25683 152
rect 25458 133 25466 143
rect 25464 109 25466 133
rect 25474 123 25475 143
rect 25485 118 25488 143
rect 25507 123 25508 143
rect 25517 133 25524 143
rect 25644 133 25651 143
rect 25660 123 25661 143
rect 25680 118 25683 143
rect 25693 123 25694 143
rect 25703 133 25710 143
rect 25474 109 25508 113
rect 25660 109 25694 113
rect 25754 109 25756 159
rect 25360 103 25402 104
rect 25766 103 25808 104
rect 25360 96 25364 103
rect 25255 62 25260 96
rect 25284 62 25289 96
rect 25327 79 25398 96
rect 25770 79 25804 96
rect 25807 79 25841 96
rect 25327 62 25402 79
rect 25360 61 25402 62
rect 25766 62 25841 79
rect 25766 61 25808 62
rect 25338 55 25424 61
rect 25744 55 25830 61
rect 25872 55 25876 233
rect 26060 183 26064 251
rect 26069 207 26079 241
rect 26089 213 26109 241
rect 26089 207 26103 213
rect 26128 207 26139 251
rect 26170 246 26246 253
rect 26279 251 26288 279
rect 26191 228 26225 246
rect 26233 228 26235 246
rect 26170 221 26246 228
rect 26233 213 26235 221
rect 26277 213 26288 251
rect 26352 241 26356 395
rect 26359 378 26364 412
rect 26388 378 26393 412
rect 26394 400 26405 412
rect 26608 395 26650 421
rect 27014 395 27056 421
rect 27271 420 27283 424
rect 27293 420 27305 424
rect 27343 420 27355 424
rect 27365 421 27377 424
rect 27535 421 27547 424
rect 27365 420 27418 421
rect 27376 412 27418 420
rect 27259 400 27270 412
rect 26540 341 26544 395
rect 26600 387 26646 395
rect 26600 383 26616 387
rect 26608 380 26616 383
rect 26642 380 26646 387
rect 26650 383 26658 395
rect 27006 383 27014 395
rect 27018 387 27052 395
rect 27018 380 27022 387
rect 27048 380 27052 387
rect 27056 383 27064 395
rect 26596 379 26662 380
rect 27002 379 27068 380
rect 26608 371 26612 379
rect 26662 365 26712 367
rect 26952 365 27002 367
rect 26702 361 26756 365
rect 26908 361 26962 365
rect 26702 356 26722 361
rect 26942 356 26962 361
rect 26712 341 26714 356
rect 26540 261 26544 329
rect 26608 305 26612 341
rect 26706 331 26714 341
rect 26722 331 26723 351
rect 26712 315 26714 331
rect 26733 322 26736 356
rect 26755 331 26756 351
rect 26765 331 26772 341
rect 26892 331 26899 341
rect 26908 331 26909 351
rect 26928 322 26931 356
rect 26941 331 26942 351
rect 26951 331 26958 341
rect 26722 315 26738 321
rect 26740 315 26756 321
rect 26908 315 26924 321
rect 26926 315 26942 321
rect 27002 315 27004 365
rect 26545 267 26581 295
rect 26545 261 26559 267
rect 26224 212 26235 213
rect 26069 183 26076 207
rect 26224 183 26234 212
rect 26315 207 26327 241
rect 26337 207 26357 241
rect 26060 103 26064 171
rect 26128 133 26132 183
rect 26128 98 26132 103
rect 25879 62 25884 96
rect 25908 62 25913 96
rect 26128 94 26166 98
rect 26128 79 26136 94
rect 26162 79 26166 94
rect 26250 94 26284 98
rect 26250 79 26254 94
rect 26280 79 26284 94
rect 26128 61 26170 79
rect 26246 61 26288 79
rect 26106 55 26192 61
rect 26224 55 26310 61
rect 26352 55 26356 207
rect 26382 183 26389 211
rect 26540 183 26544 251
rect 26549 233 26559 261
rect 26569 261 26583 267
rect 26608 261 26619 305
rect 27045 267 27056 305
rect 27083 267 27119 295
rect 27120 267 27124 395
rect 27271 378 27276 412
rect 27300 378 27305 412
rect 27306 400 27317 412
rect 27331 400 27342 412
rect 27343 395 27418 412
rect 27494 420 27547 421
rect 27557 420 27569 424
rect 27607 420 27619 424
rect 27629 420 27641 424
rect 27494 412 27536 420
rect 27494 395 27569 412
rect 27570 400 27581 412
rect 27595 400 27606 412
rect 27308 341 27312 395
rect 27343 378 27414 395
rect 27418 383 27426 395
rect 27486 383 27494 395
rect 27498 378 27532 395
rect 27535 378 27569 395
rect 27376 371 27380 378
rect 26770 262 26820 264
rect 26844 262 26894 264
rect 26569 233 26589 261
rect 26608 233 26617 261
rect 26671 253 26705 261
rect 26650 246 26705 253
rect 26671 245 26705 246
rect 26773 253 26804 261
rect 26773 245 26807 253
rect 26608 213 26612 233
rect 26804 229 26807 245
rect 26671 228 26705 229
rect 26650 221 26705 228
rect 26773 221 26807 229
rect 26820 212 26822 262
rect 26860 253 26891 261
rect 26894 253 26896 262
rect 27083 261 27095 267
rect 26860 245 26896 253
rect 26959 253 26993 261
rect 26959 246 27014 253
rect 26959 245 26993 246
rect 26891 229 26896 245
rect 27085 233 27095 261
rect 27105 233 27125 267
rect 27308 261 27312 329
rect 27376 291 27380 341
rect 27376 251 27385 279
rect 27472 264 27482 291
rect 27431 262 27482 264
rect 27472 261 27483 262
rect 27439 253 27473 261
rect 27481 253 27483 261
rect 26860 221 26896 229
rect 26959 228 26993 229
rect 26959 221 27014 228
rect 26894 212 26896 221
rect 26540 103 26544 171
rect 26608 133 26612 183
rect 26662 159 26712 161
rect 26952 159 27002 161
rect 26712 143 26714 159
rect 26722 153 26738 159
rect 26740 153 26756 159
rect 26908 153 26924 159
rect 26926 153 26942 159
rect 26733 143 26756 152
rect 26908 143 26931 152
rect 26706 133 26714 143
rect 26712 109 26714 133
rect 26722 123 26723 143
rect 26733 118 26736 143
rect 26755 123 26756 143
rect 26765 133 26772 143
rect 26892 133 26899 143
rect 26908 123 26909 143
rect 26928 118 26931 143
rect 26941 123 26942 143
rect 26951 133 26958 143
rect 26722 109 26756 113
rect 26908 109 26942 113
rect 27002 109 27004 159
rect 26608 103 26650 104
rect 27014 103 27056 104
rect 26608 96 26612 103
rect 26503 62 26508 96
rect 26532 62 26537 96
rect 26575 79 26646 96
rect 27018 79 27052 96
rect 27055 79 27089 96
rect 26575 62 26650 79
rect 26608 61 26650 62
rect 27014 62 27089 79
rect 27014 61 27056 62
rect 26586 55 26672 61
rect 26992 55 27078 61
rect 27120 55 27124 233
rect 27308 183 27312 251
rect 27317 207 27327 241
rect 27337 213 27357 241
rect 27337 207 27351 213
rect 27376 207 27387 251
rect 27418 246 27494 253
rect 27527 251 27536 279
rect 27439 228 27473 246
rect 27481 228 27483 246
rect 27418 221 27494 228
rect 27481 213 27483 221
rect 27525 213 27536 251
rect 27600 241 27604 395
rect 27607 378 27612 412
rect 27636 378 27641 412
rect 27642 400 27653 412
rect 27856 395 27898 421
rect 28262 395 28304 421
rect 28519 420 28531 424
rect 28541 420 28553 424
rect 28591 420 28603 424
rect 28613 421 28625 424
rect 28783 421 28795 424
rect 28613 420 28666 421
rect 28624 412 28666 420
rect 28507 400 28518 412
rect 27788 341 27792 395
rect 27848 387 27894 395
rect 27848 383 27864 387
rect 27856 380 27864 383
rect 27890 380 27894 387
rect 27898 383 27906 395
rect 28254 383 28262 395
rect 28266 387 28300 395
rect 28266 380 28270 387
rect 28296 380 28300 387
rect 28304 383 28312 395
rect 27844 379 27910 380
rect 28250 379 28316 380
rect 27856 371 27860 379
rect 27910 365 27960 367
rect 28200 365 28250 367
rect 27950 361 28004 365
rect 28156 361 28210 365
rect 27950 356 27970 361
rect 28190 356 28210 361
rect 27960 341 27962 356
rect 27788 261 27792 329
rect 27856 305 27860 341
rect 27954 331 27962 341
rect 27970 331 27971 351
rect 27960 315 27962 331
rect 27981 322 27984 356
rect 28003 331 28004 351
rect 28013 331 28020 341
rect 28140 331 28147 341
rect 28156 331 28157 351
rect 28176 322 28179 356
rect 28189 331 28190 351
rect 28199 331 28206 341
rect 27970 315 27986 321
rect 27988 315 28004 321
rect 28156 315 28172 321
rect 28174 315 28190 321
rect 28250 315 28252 365
rect 27793 267 27829 295
rect 27793 261 27807 267
rect 27472 212 27483 213
rect 27317 183 27324 207
rect 27472 183 27482 212
rect 27563 207 27575 241
rect 27585 207 27605 241
rect 27308 103 27312 171
rect 27376 133 27380 183
rect 27376 98 27380 103
rect 27127 62 27132 96
rect 27156 62 27161 96
rect 27376 94 27414 98
rect 27376 79 27384 94
rect 27410 79 27414 94
rect 27498 94 27532 98
rect 27498 79 27502 94
rect 27528 79 27532 94
rect 27376 61 27418 79
rect 27494 61 27536 79
rect 27354 55 27440 61
rect 27472 55 27558 61
rect 27600 55 27604 207
rect 27630 183 27637 211
rect 27788 183 27792 251
rect 27797 233 27807 261
rect 27817 261 27831 267
rect 27856 261 27867 305
rect 28293 267 28304 305
rect 28331 267 28367 295
rect 28368 267 28372 395
rect 28519 378 28524 412
rect 28548 378 28553 412
rect 28554 400 28565 412
rect 28579 400 28590 412
rect 28591 395 28666 412
rect 28742 420 28795 421
rect 28805 420 28817 424
rect 28855 420 28867 424
rect 28877 420 28889 424
rect 28742 412 28784 420
rect 28742 395 28817 412
rect 28818 400 28829 412
rect 28843 400 28854 412
rect 28556 341 28560 395
rect 28591 378 28662 395
rect 28666 383 28674 395
rect 28734 383 28742 395
rect 28746 378 28780 395
rect 28783 378 28817 395
rect 28624 371 28628 378
rect 28018 262 28068 264
rect 28092 262 28142 264
rect 27817 233 27837 261
rect 27856 233 27865 261
rect 27919 253 27953 261
rect 27898 246 27953 253
rect 27919 245 27953 246
rect 28021 253 28052 261
rect 28021 245 28055 253
rect 27856 213 27860 233
rect 28052 229 28055 245
rect 27919 228 27953 229
rect 27898 221 27953 228
rect 28021 221 28055 229
rect 28068 212 28070 262
rect 28108 253 28139 261
rect 28142 253 28144 262
rect 28331 261 28343 267
rect 28108 245 28144 253
rect 28207 253 28241 261
rect 28207 246 28262 253
rect 28207 245 28241 246
rect 28139 229 28144 245
rect 28333 233 28343 261
rect 28353 233 28373 267
rect 28556 261 28560 329
rect 28624 291 28628 341
rect 28624 251 28633 279
rect 28720 264 28730 291
rect 28679 262 28730 264
rect 28720 261 28731 262
rect 28687 253 28721 261
rect 28729 253 28731 261
rect 28108 221 28144 229
rect 28207 228 28241 229
rect 28207 221 28262 228
rect 28142 212 28144 221
rect 27788 103 27792 171
rect 27856 133 27860 183
rect 27910 159 27960 161
rect 28200 159 28250 161
rect 27960 143 27962 159
rect 27970 153 27986 159
rect 27988 153 28004 159
rect 28156 153 28172 159
rect 28174 153 28190 159
rect 27981 143 28004 152
rect 28156 143 28179 152
rect 27954 133 27962 143
rect 27960 109 27962 133
rect 27970 123 27971 143
rect 27981 118 27984 143
rect 28003 123 28004 143
rect 28013 133 28020 143
rect 28140 133 28147 143
rect 28156 123 28157 143
rect 28176 118 28179 143
rect 28189 123 28190 143
rect 28199 133 28206 143
rect 27970 109 28004 113
rect 28156 109 28190 113
rect 28250 109 28252 159
rect 27856 103 27898 104
rect 28262 103 28304 104
rect 27856 96 27860 103
rect 27751 62 27756 96
rect 27780 62 27785 96
rect 27823 79 27894 96
rect 28266 79 28300 96
rect 28303 79 28337 96
rect 27823 62 27898 79
rect 27856 61 27898 62
rect 28262 62 28337 79
rect 28262 61 28304 62
rect 27834 55 27920 61
rect 28240 55 28326 61
rect 28368 55 28372 233
rect 28556 183 28560 251
rect 28565 207 28575 241
rect 28585 213 28605 241
rect 28585 207 28599 213
rect 28624 207 28635 251
rect 28666 246 28742 253
rect 28775 251 28784 279
rect 28687 228 28721 246
rect 28729 228 28731 246
rect 28666 221 28742 228
rect 28729 213 28731 221
rect 28773 213 28784 251
rect 28848 241 28852 395
rect 28855 378 28860 412
rect 28884 378 28889 412
rect 28890 400 28901 412
rect 29104 395 29146 421
rect 29510 395 29552 421
rect 29767 420 29779 424
rect 29789 420 29801 424
rect 29839 420 29851 424
rect 29861 421 29873 424
rect 30031 421 30043 424
rect 29861 420 29914 421
rect 29872 412 29914 420
rect 29755 400 29766 412
rect 29036 341 29040 395
rect 29096 387 29142 395
rect 29096 383 29112 387
rect 29104 380 29112 383
rect 29138 380 29142 387
rect 29146 383 29154 395
rect 29502 383 29510 395
rect 29514 387 29548 395
rect 29514 380 29518 387
rect 29544 380 29548 387
rect 29552 383 29560 395
rect 29092 379 29158 380
rect 29498 379 29564 380
rect 29104 371 29108 379
rect 29158 365 29208 367
rect 29448 365 29498 367
rect 29198 361 29252 365
rect 29404 361 29458 365
rect 29198 356 29218 361
rect 29438 356 29458 361
rect 29208 341 29210 356
rect 29036 261 29040 329
rect 29104 305 29108 341
rect 29202 331 29210 341
rect 29218 331 29219 351
rect 29208 315 29210 331
rect 29229 322 29232 356
rect 29251 331 29252 351
rect 29261 331 29268 341
rect 29388 331 29395 341
rect 29404 331 29405 351
rect 29424 322 29427 356
rect 29437 331 29438 351
rect 29447 331 29454 341
rect 29218 315 29234 321
rect 29236 315 29252 321
rect 29404 315 29420 321
rect 29422 315 29438 321
rect 29498 315 29500 365
rect 29041 267 29077 295
rect 29041 261 29055 267
rect 28720 212 28731 213
rect 28565 183 28572 207
rect 28720 183 28730 212
rect 28811 207 28823 241
rect 28833 207 28853 241
rect 28556 103 28560 171
rect 28624 133 28628 183
rect 28624 98 28628 103
rect 28375 62 28380 96
rect 28404 62 28409 96
rect 28624 94 28662 98
rect 28624 79 28632 94
rect 28658 79 28662 94
rect 28746 94 28780 98
rect 28746 79 28750 94
rect 28776 79 28780 94
rect 28624 61 28666 79
rect 28742 61 28784 79
rect 28602 55 28688 61
rect 28720 55 28806 61
rect 28848 55 28852 207
rect 28878 183 28885 211
rect 29036 183 29040 251
rect 29045 233 29055 261
rect 29065 261 29079 267
rect 29104 261 29115 305
rect 29541 267 29552 305
rect 29579 267 29615 295
rect 29616 267 29620 395
rect 29767 378 29772 412
rect 29796 378 29801 412
rect 29802 400 29813 412
rect 29827 400 29838 412
rect 29839 395 29914 412
rect 29990 420 30043 421
rect 30053 420 30065 424
rect 30103 420 30115 424
rect 30125 420 30137 424
rect 29990 412 30032 420
rect 29990 395 30065 412
rect 30066 400 30077 412
rect 30091 400 30102 412
rect 29804 341 29808 395
rect 29839 378 29910 395
rect 29914 383 29922 395
rect 29982 383 29990 395
rect 29994 378 30028 395
rect 30031 378 30065 395
rect 29872 371 29876 378
rect 29266 262 29316 264
rect 29340 262 29390 264
rect 29065 233 29085 261
rect 29104 233 29113 261
rect 29167 253 29201 261
rect 29146 246 29201 253
rect 29167 245 29201 246
rect 29269 253 29300 261
rect 29269 245 29303 253
rect 29104 213 29108 233
rect 29300 229 29303 245
rect 29167 228 29201 229
rect 29146 221 29201 228
rect 29269 221 29303 229
rect 29316 212 29318 262
rect 29356 253 29387 261
rect 29390 253 29392 262
rect 29579 261 29591 267
rect 29356 245 29392 253
rect 29455 253 29489 261
rect 29455 246 29510 253
rect 29455 245 29489 246
rect 29387 229 29392 245
rect 29581 233 29591 261
rect 29601 233 29621 267
rect 29804 261 29808 329
rect 29872 291 29876 341
rect 29872 251 29881 279
rect 29968 264 29978 291
rect 29927 262 29978 264
rect 29968 261 29979 262
rect 29935 253 29969 261
rect 29977 253 29979 261
rect 29356 221 29392 229
rect 29455 228 29489 229
rect 29455 221 29510 228
rect 29390 212 29392 221
rect 29036 103 29040 171
rect 29104 133 29108 183
rect 29158 159 29208 161
rect 29448 159 29498 161
rect 29208 143 29210 159
rect 29218 153 29234 159
rect 29236 153 29252 159
rect 29404 153 29420 159
rect 29422 153 29438 159
rect 29229 143 29252 152
rect 29404 143 29427 152
rect 29202 133 29210 143
rect 29208 109 29210 133
rect 29218 123 29219 143
rect 29229 118 29232 143
rect 29251 123 29252 143
rect 29261 133 29268 143
rect 29388 133 29395 143
rect 29404 123 29405 143
rect 29424 118 29427 143
rect 29437 123 29438 143
rect 29447 133 29454 143
rect 29218 109 29252 113
rect 29404 109 29438 113
rect 29498 109 29500 159
rect 29104 103 29146 104
rect 29510 103 29552 104
rect 29104 96 29108 103
rect 28999 62 29004 96
rect 29028 62 29033 96
rect 29071 79 29142 96
rect 29514 79 29548 96
rect 29551 79 29585 96
rect 29071 62 29146 79
rect 29104 61 29146 62
rect 29510 62 29585 79
rect 29510 61 29552 62
rect 29082 55 29168 61
rect 29488 55 29574 61
rect 29616 55 29620 233
rect 29804 183 29808 251
rect 29813 207 29823 241
rect 29833 213 29853 241
rect 29833 207 29847 213
rect 29872 207 29883 251
rect 29914 246 29990 253
rect 30023 251 30032 279
rect 29935 228 29969 246
rect 29977 228 29979 246
rect 29914 221 29990 228
rect 29977 213 29979 221
rect 30021 213 30032 251
rect 30096 241 30100 395
rect 30103 378 30108 412
rect 30132 378 30137 412
rect 30138 400 30149 412
rect 30352 395 30394 421
rect 30758 395 30800 421
rect 31015 420 31027 424
rect 31037 420 31049 424
rect 31087 420 31099 424
rect 31109 421 31121 424
rect 31279 421 31291 424
rect 31109 420 31162 421
rect 31120 412 31162 420
rect 31003 400 31014 412
rect 30284 341 30288 395
rect 30344 387 30390 395
rect 30344 383 30360 387
rect 30352 380 30360 383
rect 30386 380 30390 387
rect 30394 383 30402 395
rect 30750 383 30758 395
rect 30762 387 30796 395
rect 30762 380 30766 387
rect 30792 380 30796 387
rect 30800 383 30808 395
rect 30340 379 30406 380
rect 30746 379 30812 380
rect 30352 371 30356 379
rect 30406 365 30456 367
rect 30696 365 30746 367
rect 30446 361 30500 365
rect 30652 361 30706 365
rect 30446 356 30466 361
rect 30686 356 30706 361
rect 30456 341 30458 356
rect 30284 261 30288 329
rect 30352 305 30356 341
rect 30450 331 30458 341
rect 30466 331 30467 351
rect 30456 315 30458 331
rect 30477 322 30480 356
rect 30499 331 30500 351
rect 30509 331 30516 341
rect 30636 331 30643 341
rect 30652 331 30653 351
rect 30672 322 30675 356
rect 30685 331 30686 351
rect 30695 331 30702 341
rect 30466 315 30482 321
rect 30484 315 30500 321
rect 30652 315 30668 321
rect 30670 315 30686 321
rect 30746 315 30748 365
rect 30289 267 30325 295
rect 30289 261 30303 267
rect 29968 212 29979 213
rect 29813 183 29820 207
rect 29968 183 29978 212
rect 30059 207 30071 241
rect 30081 207 30101 241
rect 29804 103 29808 171
rect 29872 133 29876 183
rect 29872 98 29876 103
rect 29623 62 29628 96
rect 29652 62 29657 96
rect 29872 94 29910 98
rect 29872 79 29880 94
rect 29906 79 29910 94
rect 29994 94 30028 98
rect 29994 79 29998 94
rect 30024 79 30028 94
rect 29872 61 29914 79
rect 29990 61 30032 79
rect 29850 55 29936 61
rect 29968 55 30054 61
rect 30096 55 30100 207
rect 30126 183 30133 211
rect 30284 183 30288 251
rect 30293 233 30303 261
rect 30313 261 30327 267
rect 30352 261 30363 305
rect 30789 267 30800 305
rect 30827 267 30863 295
rect 30864 267 30868 395
rect 31015 378 31020 412
rect 31044 378 31049 412
rect 31050 400 31061 412
rect 31075 400 31086 412
rect 31087 395 31162 412
rect 31238 420 31291 421
rect 31301 420 31313 424
rect 31351 420 31363 424
rect 31373 420 31385 424
rect 31238 412 31280 420
rect 31238 395 31313 412
rect 31314 400 31325 412
rect 31339 400 31350 412
rect 31052 341 31056 395
rect 31087 378 31158 395
rect 31162 383 31170 395
rect 31230 383 31238 395
rect 31242 378 31276 395
rect 31279 378 31313 395
rect 31120 371 31124 378
rect 30514 262 30564 264
rect 30588 262 30638 264
rect 30313 233 30333 261
rect 30352 233 30361 261
rect 30415 253 30449 261
rect 30394 246 30449 253
rect 30415 245 30449 246
rect 30517 253 30548 261
rect 30517 245 30551 253
rect 30352 213 30356 233
rect 30548 229 30551 245
rect 30415 228 30449 229
rect 30394 221 30449 228
rect 30517 221 30551 229
rect 30564 212 30566 262
rect 30604 253 30635 261
rect 30638 253 30640 262
rect 30827 261 30839 267
rect 30604 245 30640 253
rect 30703 253 30737 261
rect 30703 246 30758 253
rect 30703 245 30737 246
rect 30635 229 30640 245
rect 30829 233 30839 261
rect 30849 233 30869 267
rect 31052 261 31056 329
rect 31120 291 31124 341
rect 31120 251 31129 279
rect 31216 264 31226 291
rect 31175 262 31226 264
rect 31216 261 31227 262
rect 31183 253 31217 261
rect 31225 253 31227 261
rect 30604 221 30640 229
rect 30703 228 30737 229
rect 30703 221 30758 228
rect 30638 212 30640 221
rect 30284 103 30288 171
rect 30352 133 30356 183
rect 30406 159 30456 161
rect 30696 159 30746 161
rect 30456 143 30458 159
rect 30466 153 30482 159
rect 30484 153 30500 159
rect 30652 153 30668 159
rect 30670 153 30686 159
rect 30477 143 30500 152
rect 30652 143 30675 152
rect 30450 133 30458 143
rect 30456 109 30458 133
rect 30466 123 30467 143
rect 30477 118 30480 143
rect 30499 123 30500 143
rect 30509 133 30516 143
rect 30636 133 30643 143
rect 30652 123 30653 143
rect 30672 118 30675 143
rect 30685 123 30686 143
rect 30695 133 30702 143
rect 30466 109 30500 113
rect 30652 109 30686 113
rect 30746 109 30748 159
rect 30352 103 30394 104
rect 30758 103 30800 104
rect 30352 96 30356 103
rect 30247 62 30252 96
rect 30276 62 30281 96
rect 30319 79 30390 96
rect 30762 79 30796 96
rect 30799 79 30833 96
rect 30319 62 30394 79
rect 30352 61 30394 62
rect 30758 62 30833 79
rect 30758 61 30800 62
rect 30330 55 30416 61
rect 30736 55 30822 61
rect 30864 55 30868 233
rect 31052 183 31056 251
rect 31061 207 31071 241
rect 31081 213 31101 241
rect 31081 207 31095 213
rect 31120 207 31131 251
rect 31162 246 31238 253
rect 31271 251 31280 279
rect 31183 228 31217 246
rect 31225 228 31227 246
rect 31162 221 31238 228
rect 31225 213 31227 221
rect 31269 213 31280 251
rect 31344 241 31348 395
rect 31351 378 31356 412
rect 31380 378 31385 412
rect 31386 400 31397 412
rect 31600 395 31642 421
rect 32006 395 32048 421
rect 32263 420 32275 424
rect 32285 420 32297 424
rect 32335 420 32347 424
rect 32357 421 32369 424
rect 32527 421 32539 424
rect 32357 420 32410 421
rect 32368 412 32410 420
rect 32251 400 32262 412
rect 31532 341 31536 395
rect 31592 387 31638 395
rect 31592 383 31608 387
rect 31600 380 31608 383
rect 31634 380 31638 387
rect 31642 383 31650 395
rect 31998 383 32006 395
rect 32010 387 32044 395
rect 32010 380 32014 387
rect 32040 380 32044 387
rect 32048 383 32056 395
rect 31588 379 31654 380
rect 31994 379 32060 380
rect 31600 371 31604 379
rect 31654 365 31704 367
rect 31944 365 31994 367
rect 31694 361 31748 365
rect 31900 361 31954 365
rect 31694 356 31714 361
rect 31934 356 31954 361
rect 31704 341 31706 356
rect 31532 261 31536 329
rect 31600 305 31604 341
rect 31698 331 31706 341
rect 31714 331 31715 351
rect 31704 315 31706 331
rect 31725 322 31728 356
rect 31747 331 31748 351
rect 31757 331 31764 341
rect 31884 331 31891 341
rect 31900 331 31901 351
rect 31920 322 31923 356
rect 31933 331 31934 351
rect 31943 331 31950 341
rect 31714 315 31730 321
rect 31732 315 31748 321
rect 31900 315 31916 321
rect 31918 315 31934 321
rect 31994 315 31996 365
rect 31537 267 31573 295
rect 31537 261 31551 267
rect 31216 212 31227 213
rect 31061 183 31068 207
rect 31216 183 31226 212
rect 31307 207 31319 241
rect 31329 207 31349 241
rect 31052 103 31056 171
rect 31120 133 31124 183
rect 31120 98 31124 103
rect 30871 62 30876 96
rect 30900 62 30905 96
rect 31120 94 31158 98
rect 31120 79 31128 94
rect 31154 79 31158 94
rect 31242 94 31276 98
rect 31242 79 31246 94
rect 31272 79 31276 94
rect 31120 61 31162 79
rect 31238 61 31280 79
rect 31098 55 31184 61
rect 31216 55 31302 61
rect 31344 55 31348 207
rect 31374 183 31381 211
rect 31532 183 31536 251
rect 31541 233 31551 261
rect 31561 261 31575 267
rect 31600 261 31611 305
rect 32037 267 32048 305
rect 32075 267 32111 295
rect 32112 267 32116 395
rect 32263 378 32268 412
rect 32292 378 32297 412
rect 32298 400 32309 412
rect 32323 400 32334 412
rect 32335 395 32410 412
rect 32486 420 32539 421
rect 32549 420 32561 424
rect 32599 420 32611 424
rect 32621 420 32633 424
rect 32486 412 32528 420
rect 32486 395 32561 412
rect 32562 400 32573 412
rect 32587 400 32598 412
rect 32300 341 32304 395
rect 32335 378 32406 395
rect 32410 383 32418 395
rect 32478 383 32486 395
rect 32490 378 32524 395
rect 32527 378 32561 395
rect 32368 371 32372 378
rect 31762 262 31812 264
rect 31836 262 31886 264
rect 31561 233 31581 261
rect 31600 233 31609 261
rect 31663 253 31697 261
rect 31642 246 31697 253
rect 31663 245 31697 246
rect 31765 253 31796 261
rect 31765 245 31799 253
rect 31600 213 31604 233
rect 31796 229 31799 245
rect 31663 228 31697 229
rect 31642 221 31697 228
rect 31765 221 31799 229
rect 31812 212 31814 262
rect 31852 253 31883 261
rect 31886 253 31888 262
rect 32075 261 32087 267
rect 31852 245 31888 253
rect 31951 253 31985 261
rect 31951 246 32006 253
rect 31951 245 31985 246
rect 31883 229 31888 245
rect 32077 233 32087 261
rect 32097 233 32117 267
rect 32300 261 32304 329
rect 32368 291 32372 341
rect 32368 251 32377 279
rect 32464 264 32474 291
rect 32423 262 32474 264
rect 32464 261 32475 262
rect 32431 253 32465 261
rect 32473 253 32475 261
rect 31852 221 31888 229
rect 31951 228 31985 229
rect 31951 221 32006 228
rect 31886 212 31888 221
rect 31532 103 31536 171
rect 31600 133 31604 183
rect 31654 159 31704 161
rect 31944 159 31994 161
rect 31704 143 31706 159
rect 31714 153 31730 159
rect 31732 153 31748 159
rect 31900 153 31916 159
rect 31918 153 31934 159
rect 31725 143 31748 152
rect 31900 143 31923 152
rect 31698 133 31706 143
rect 31704 109 31706 133
rect 31714 123 31715 143
rect 31725 118 31728 143
rect 31747 123 31748 143
rect 31757 133 31764 143
rect 31884 133 31891 143
rect 31900 123 31901 143
rect 31920 118 31923 143
rect 31933 123 31934 143
rect 31943 133 31950 143
rect 31714 109 31748 113
rect 31900 109 31934 113
rect 31994 109 31996 159
rect 31600 103 31642 104
rect 32006 103 32048 104
rect 31600 96 31604 103
rect 31495 62 31500 96
rect 31524 62 31529 96
rect 31567 79 31638 96
rect 32010 79 32044 96
rect 32047 79 32081 96
rect 31567 62 31642 79
rect 31600 61 31642 62
rect 32006 62 32081 79
rect 32006 61 32048 62
rect 31578 55 31664 61
rect 31984 55 32070 61
rect 32112 55 32116 233
rect 32300 183 32304 251
rect 32309 207 32319 241
rect 32329 213 32349 241
rect 32329 207 32343 213
rect 32368 207 32379 251
rect 32410 246 32486 253
rect 32519 251 32528 279
rect 32431 228 32465 246
rect 32473 228 32475 246
rect 32410 221 32486 228
rect 32473 213 32475 221
rect 32517 213 32528 251
rect 32592 241 32596 395
rect 32599 378 32604 412
rect 32628 378 32633 412
rect 32634 400 32645 412
rect 32848 395 32890 421
rect 33254 395 33296 421
rect 33511 420 33523 424
rect 33533 420 33545 424
rect 33583 420 33595 424
rect 33605 421 33617 424
rect 33775 421 33787 424
rect 33605 420 33658 421
rect 33616 412 33658 420
rect 33499 400 33510 412
rect 32780 341 32784 395
rect 32840 387 32886 395
rect 32840 383 32856 387
rect 32848 380 32856 383
rect 32882 380 32886 387
rect 32890 383 32898 395
rect 33246 383 33254 395
rect 33258 387 33292 395
rect 33258 380 33262 387
rect 33288 380 33292 387
rect 33296 383 33304 395
rect 32836 379 32902 380
rect 33242 379 33308 380
rect 32848 371 32852 379
rect 32902 365 32952 367
rect 33192 365 33242 367
rect 32942 361 32996 365
rect 33148 361 33202 365
rect 32942 356 32962 361
rect 33182 356 33202 361
rect 32952 341 32954 356
rect 32780 261 32784 329
rect 32848 305 32852 341
rect 32946 331 32954 341
rect 32962 331 32963 351
rect 32952 315 32954 331
rect 32973 322 32976 356
rect 32995 331 32996 351
rect 33005 331 33012 341
rect 33132 331 33139 341
rect 33148 331 33149 351
rect 33168 322 33171 356
rect 33181 331 33182 351
rect 33191 331 33198 341
rect 32962 315 32978 321
rect 32980 315 32996 321
rect 33148 315 33164 321
rect 33166 315 33182 321
rect 33242 315 33244 365
rect 32785 267 32821 295
rect 32785 261 32799 267
rect 32464 212 32475 213
rect 32309 183 32316 207
rect 32464 183 32474 212
rect 32555 207 32567 241
rect 32577 207 32597 241
rect 32300 103 32304 171
rect 32368 133 32372 183
rect 32368 98 32372 103
rect 32119 62 32124 96
rect 32148 62 32153 96
rect 32368 94 32406 98
rect 32368 79 32376 94
rect 32402 79 32406 94
rect 32490 94 32524 98
rect 32490 79 32494 94
rect 32520 79 32524 94
rect 32368 61 32410 79
rect 32486 61 32528 79
rect 32346 55 32432 61
rect 32464 55 32550 61
rect 32592 55 32596 207
rect 32622 183 32629 211
rect 32780 183 32784 251
rect 32789 233 32799 261
rect 32809 261 32823 267
rect 32848 261 32859 305
rect 33285 267 33296 305
rect 33323 267 33359 295
rect 33360 267 33364 395
rect 33511 378 33516 412
rect 33540 378 33545 412
rect 33546 400 33557 412
rect 33571 400 33582 412
rect 33583 395 33658 412
rect 33734 420 33787 421
rect 33797 420 33809 424
rect 33847 420 33859 424
rect 33869 420 33881 424
rect 33734 412 33776 420
rect 33734 395 33809 412
rect 33810 400 33821 412
rect 33835 400 33846 412
rect 33548 341 33552 395
rect 33583 378 33654 395
rect 33658 383 33666 395
rect 33726 383 33734 395
rect 33738 378 33772 395
rect 33775 378 33809 395
rect 33616 371 33620 378
rect 33010 262 33060 264
rect 33084 262 33134 264
rect 32809 233 32829 261
rect 32848 233 32857 261
rect 32911 253 32945 261
rect 32890 246 32945 253
rect 32911 245 32945 246
rect 33013 253 33044 261
rect 33013 245 33047 253
rect 32848 213 32852 233
rect 33044 229 33047 245
rect 32911 228 32945 229
rect 32890 221 32945 228
rect 33013 221 33047 229
rect 33060 212 33062 262
rect 33100 253 33131 261
rect 33134 253 33136 262
rect 33323 261 33335 267
rect 33100 245 33136 253
rect 33199 253 33233 261
rect 33199 246 33254 253
rect 33199 245 33233 246
rect 33131 229 33136 245
rect 33325 233 33335 261
rect 33345 233 33365 267
rect 33548 261 33552 329
rect 33616 291 33620 341
rect 33616 251 33625 279
rect 33712 264 33722 291
rect 33671 262 33722 264
rect 33712 261 33723 262
rect 33679 253 33713 261
rect 33721 253 33723 261
rect 33100 221 33136 229
rect 33199 228 33233 229
rect 33199 221 33254 228
rect 33134 212 33136 221
rect 32780 103 32784 171
rect 32848 133 32852 183
rect 32902 159 32952 161
rect 33192 159 33242 161
rect 32952 143 32954 159
rect 32962 153 32978 159
rect 32980 153 32996 159
rect 33148 153 33164 159
rect 33166 153 33182 159
rect 32973 143 32996 152
rect 33148 143 33171 152
rect 32946 133 32954 143
rect 32952 109 32954 133
rect 32962 123 32963 143
rect 32973 118 32976 143
rect 32995 123 32996 143
rect 33005 133 33012 143
rect 33132 133 33139 143
rect 33148 123 33149 143
rect 33168 118 33171 143
rect 33181 123 33182 143
rect 33191 133 33198 143
rect 32962 109 32996 113
rect 33148 109 33182 113
rect 33242 109 33244 159
rect 32848 103 32890 104
rect 33254 103 33296 104
rect 32848 96 32852 103
rect 32743 62 32748 96
rect 32772 62 32777 96
rect 32815 79 32886 96
rect 33258 79 33292 96
rect 33295 79 33329 96
rect 32815 62 32890 79
rect 32848 61 32890 62
rect 33254 62 33329 79
rect 33254 61 33296 62
rect 32826 55 32912 61
rect 33232 55 33318 61
rect 33360 55 33364 233
rect 33548 183 33552 251
rect 33557 207 33567 241
rect 33577 213 33597 241
rect 33577 207 33591 213
rect 33616 207 33627 251
rect 33658 246 33734 253
rect 33767 251 33776 279
rect 33679 228 33713 246
rect 33721 228 33723 246
rect 33658 221 33734 228
rect 33721 213 33723 221
rect 33765 213 33776 251
rect 33840 241 33844 395
rect 33847 378 33852 412
rect 33876 378 33881 412
rect 33882 400 33893 412
rect 34096 395 34138 421
rect 34502 395 34544 421
rect 34759 420 34771 424
rect 34781 420 34793 424
rect 34831 420 34843 424
rect 34853 421 34865 424
rect 35023 421 35035 424
rect 34853 420 34906 421
rect 34864 412 34906 420
rect 34747 400 34758 412
rect 34028 341 34032 395
rect 34088 387 34134 395
rect 34088 383 34104 387
rect 34096 380 34104 383
rect 34130 380 34134 387
rect 34138 383 34146 395
rect 34494 383 34502 395
rect 34506 387 34540 395
rect 34506 380 34510 387
rect 34536 380 34540 387
rect 34544 383 34552 395
rect 34084 379 34150 380
rect 34490 379 34556 380
rect 34096 371 34100 379
rect 34150 365 34200 367
rect 34440 365 34490 367
rect 34190 361 34244 365
rect 34396 361 34450 365
rect 34190 356 34210 361
rect 34430 356 34450 361
rect 34200 341 34202 356
rect 34028 261 34032 329
rect 34096 305 34100 341
rect 34194 331 34202 341
rect 34210 331 34211 351
rect 34200 315 34202 331
rect 34221 322 34224 356
rect 34243 331 34244 351
rect 34253 331 34260 341
rect 34380 331 34387 341
rect 34396 331 34397 351
rect 34416 322 34419 356
rect 34429 331 34430 351
rect 34439 331 34446 341
rect 34210 315 34226 321
rect 34228 315 34244 321
rect 34396 315 34412 321
rect 34414 315 34430 321
rect 34490 315 34492 365
rect 34033 267 34069 295
rect 34033 261 34047 267
rect 33712 212 33723 213
rect 33557 183 33564 207
rect 33712 183 33722 212
rect 33803 207 33815 241
rect 33825 207 33845 241
rect 33548 103 33552 171
rect 33616 133 33620 183
rect 33616 98 33620 103
rect 33367 62 33372 96
rect 33396 62 33401 96
rect 33616 94 33654 98
rect 33616 79 33624 94
rect 33650 79 33654 94
rect 33738 94 33772 98
rect 33738 79 33742 94
rect 33768 79 33772 94
rect 33616 61 33658 79
rect 33734 61 33776 79
rect 33594 55 33680 61
rect 33712 55 33798 61
rect 33840 55 33844 207
rect 33870 183 33877 211
rect 34028 183 34032 251
rect 34037 233 34047 261
rect 34057 261 34071 267
rect 34096 261 34107 305
rect 34533 267 34544 305
rect 34571 267 34607 295
rect 34608 267 34612 395
rect 34759 378 34764 412
rect 34788 378 34793 412
rect 34794 400 34805 412
rect 34819 400 34830 412
rect 34831 395 34906 412
rect 34982 420 35035 421
rect 35045 420 35057 424
rect 35095 420 35107 424
rect 35117 420 35129 424
rect 34982 412 35024 420
rect 34982 395 35057 412
rect 35058 400 35069 412
rect 35083 400 35094 412
rect 34796 341 34800 395
rect 34831 378 34902 395
rect 34906 383 34914 395
rect 34974 383 34982 395
rect 34986 378 35020 395
rect 35023 378 35057 395
rect 34864 371 34868 378
rect 34258 262 34308 264
rect 34332 262 34382 264
rect 34057 233 34077 261
rect 34096 233 34105 261
rect 34159 253 34193 261
rect 34138 246 34193 253
rect 34159 245 34193 246
rect 34261 253 34292 261
rect 34261 245 34295 253
rect 34096 213 34100 233
rect 34292 229 34295 245
rect 34159 228 34193 229
rect 34138 221 34193 228
rect 34261 221 34295 229
rect 34308 212 34310 262
rect 34348 253 34379 261
rect 34382 253 34384 262
rect 34571 261 34583 267
rect 34348 245 34384 253
rect 34447 253 34481 261
rect 34447 246 34502 253
rect 34447 245 34481 246
rect 34379 229 34384 245
rect 34573 233 34583 261
rect 34593 233 34613 267
rect 34796 261 34800 329
rect 34864 291 34868 341
rect 34864 251 34873 279
rect 34960 264 34970 291
rect 34919 262 34970 264
rect 34960 261 34971 262
rect 34927 253 34961 261
rect 34969 253 34971 261
rect 34348 221 34384 229
rect 34447 228 34481 229
rect 34447 221 34502 228
rect 34382 212 34384 221
rect 34028 103 34032 171
rect 34096 133 34100 183
rect 34150 159 34200 161
rect 34440 159 34490 161
rect 34200 143 34202 159
rect 34210 153 34226 159
rect 34228 153 34244 159
rect 34396 153 34412 159
rect 34414 153 34430 159
rect 34221 143 34244 152
rect 34396 143 34419 152
rect 34194 133 34202 143
rect 34200 109 34202 133
rect 34210 123 34211 143
rect 34221 118 34224 143
rect 34243 123 34244 143
rect 34253 133 34260 143
rect 34380 133 34387 143
rect 34396 123 34397 143
rect 34416 118 34419 143
rect 34429 123 34430 143
rect 34439 133 34446 143
rect 34210 109 34244 113
rect 34396 109 34430 113
rect 34490 109 34492 159
rect 34096 103 34138 104
rect 34502 103 34544 104
rect 34096 96 34100 103
rect 33991 62 33996 96
rect 34020 62 34025 96
rect 34063 79 34134 96
rect 34506 79 34540 96
rect 34543 79 34577 96
rect 34063 62 34138 79
rect 34096 61 34138 62
rect 34502 62 34577 79
rect 34502 61 34544 62
rect 34074 55 34160 61
rect 34480 55 34566 61
rect 34608 55 34612 233
rect 34796 183 34800 251
rect 34805 207 34815 241
rect 34825 213 34845 241
rect 34825 207 34839 213
rect 34864 207 34875 251
rect 34906 246 34982 253
rect 35015 251 35024 279
rect 34927 228 34961 246
rect 34969 228 34971 246
rect 34906 221 34982 228
rect 34969 213 34971 221
rect 35013 213 35024 251
rect 35088 241 35092 395
rect 35095 378 35100 412
rect 35124 378 35129 412
rect 35130 400 35141 412
rect 35344 395 35386 421
rect 35750 395 35792 421
rect 36007 420 36019 424
rect 36029 420 36041 424
rect 36079 420 36091 424
rect 36101 421 36113 424
rect 36271 421 36283 424
rect 36101 420 36154 421
rect 36112 412 36154 420
rect 35995 400 36006 412
rect 35276 341 35280 395
rect 35336 387 35382 395
rect 35336 383 35352 387
rect 35344 380 35352 383
rect 35378 380 35382 387
rect 35386 383 35394 395
rect 35742 383 35750 395
rect 35754 387 35788 395
rect 35754 380 35758 387
rect 35784 380 35788 387
rect 35792 383 35800 395
rect 35332 379 35398 380
rect 35738 379 35804 380
rect 35344 371 35348 379
rect 35398 365 35448 367
rect 35688 365 35738 367
rect 35438 361 35492 365
rect 35644 361 35698 365
rect 35438 356 35458 361
rect 35678 356 35698 361
rect 35448 341 35450 356
rect 35276 261 35280 329
rect 35344 305 35348 341
rect 35442 331 35450 341
rect 35458 331 35459 351
rect 35448 315 35450 331
rect 35469 322 35472 356
rect 35491 331 35492 351
rect 35501 331 35508 341
rect 35628 331 35635 341
rect 35644 331 35645 351
rect 35664 322 35667 356
rect 35677 331 35678 351
rect 35687 331 35694 341
rect 35458 315 35474 321
rect 35476 315 35492 321
rect 35644 315 35660 321
rect 35662 315 35678 321
rect 35738 315 35740 365
rect 35281 267 35317 295
rect 35281 261 35295 267
rect 34960 212 34971 213
rect 34805 183 34812 207
rect 34960 183 34970 212
rect 35051 207 35063 241
rect 35073 207 35093 241
rect 34796 103 34800 171
rect 34864 133 34868 183
rect 34864 98 34868 103
rect 34615 62 34620 96
rect 34644 62 34649 96
rect 34864 94 34902 98
rect 34864 79 34872 94
rect 34898 79 34902 94
rect 34986 94 35020 98
rect 34986 79 34990 94
rect 35016 79 35020 94
rect 34864 61 34906 79
rect 34982 61 35024 79
rect 34842 55 34928 61
rect 34960 55 35046 61
rect 35088 55 35092 207
rect 35118 183 35125 211
rect 35276 183 35280 251
rect 35285 233 35295 261
rect 35305 261 35319 267
rect 35344 261 35355 305
rect 35781 267 35792 305
rect 35819 267 35855 295
rect 35856 267 35860 395
rect 36007 378 36012 412
rect 36036 378 36041 412
rect 36042 400 36053 412
rect 36067 400 36078 412
rect 36079 395 36154 412
rect 36230 420 36283 421
rect 36293 420 36305 424
rect 36343 420 36355 424
rect 36365 420 36377 424
rect 36230 412 36272 420
rect 36230 395 36305 412
rect 36306 400 36317 412
rect 36331 400 36342 412
rect 36044 341 36048 395
rect 36079 378 36150 395
rect 36154 383 36162 395
rect 36222 383 36230 395
rect 36234 378 36268 395
rect 36271 378 36305 395
rect 36112 371 36116 378
rect 35506 262 35556 264
rect 35580 262 35630 264
rect 35305 233 35325 261
rect 35344 233 35353 261
rect 35407 253 35441 261
rect 35386 246 35441 253
rect 35407 245 35441 246
rect 35509 253 35540 261
rect 35509 245 35543 253
rect 35344 213 35348 233
rect 35540 229 35543 245
rect 35407 228 35441 229
rect 35386 221 35441 228
rect 35509 221 35543 229
rect 35556 212 35558 262
rect 35596 253 35627 261
rect 35630 253 35632 262
rect 35819 261 35831 267
rect 35596 245 35632 253
rect 35695 253 35729 261
rect 35695 246 35750 253
rect 35695 245 35729 246
rect 35627 229 35632 245
rect 35821 233 35831 261
rect 35841 233 35861 267
rect 36044 261 36048 329
rect 36112 291 36116 341
rect 36112 251 36121 279
rect 36208 264 36218 291
rect 36167 262 36218 264
rect 36208 261 36219 262
rect 36175 253 36209 261
rect 36217 253 36219 261
rect 35596 221 35632 229
rect 35695 228 35729 229
rect 35695 221 35750 228
rect 35630 212 35632 221
rect 35276 103 35280 171
rect 35344 133 35348 183
rect 35398 159 35448 161
rect 35688 159 35738 161
rect 35448 143 35450 159
rect 35458 153 35474 159
rect 35476 153 35492 159
rect 35644 153 35660 159
rect 35662 153 35678 159
rect 35469 143 35492 152
rect 35644 143 35667 152
rect 35442 133 35450 143
rect 35448 109 35450 133
rect 35458 123 35459 143
rect 35469 118 35472 143
rect 35491 123 35492 143
rect 35501 133 35508 143
rect 35628 133 35635 143
rect 35644 123 35645 143
rect 35664 118 35667 143
rect 35677 123 35678 143
rect 35687 133 35694 143
rect 35458 109 35492 113
rect 35644 109 35678 113
rect 35738 109 35740 159
rect 35344 103 35386 104
rect 35750 103 35792 104
rect 35344 96 35348 103
rect 35239 62 35244 96
rect 35268 62 35273 96
rect 35311 79 35382 96
rect 35754 79 35788 96
rect 35791 79 35825 96
rect 35311 62 35386 79
rect 35344 61 35386 62
rect 35750 62 35825 79
rect 35750 61 35792 62
rect 35322 55 35408 61
rect 35728 55 35814 61
rect 35856 55 35860 233
rect 36044 183 36048 251
rect 36053 207 36063 241
rect 36073 213 36093 241
rect 36073 207 36087 213
rect 36112 207 36123 251
rect 36154 246 36230 253
rect 36263 251 36272 279
rect 36175 228 36209 246
rect 36217 228 36219 246
rect 36154 221 36230 228
rect 36217 213 36219 221
rect 36261 213 36272 251
rect 36336 241 36340 395
rect 36343 378 36348 412
rect 36372 378 36377 412
rect 36378 400 36389 412
rect 36592 395 36634 421
rect 36998 395 37040 421
rect 37255 420 37267 424
rect 37277 420 37289 424
rect 37327 420 37339 424
rect 37349 421 37361 424
rect 37519 421 37531 424
rect 37349 420 37402 421
rect 37360 412 37402 420
rect 37243 400 37254 412
rect 36524 341 36528 395
rect 36584 387 36630 395
rect 36584 383 36600 387
rect 36592 380 36600 383
rect 36626 380 36630 387
rect 36634 383 36642 395
rect 36990 383 36998 395
rect 37002 387 37036 395
rect 37002 380 37006 387
rect 37032 380 37036 387
rect 37040 383 37048 395
rect 36580 379 36646 380
rect 36986 379 37052 380
rect 36592 371 36596 379
rect 36646 365 36696 367
rect 36936 365 36986 367
rect 36686 361 36740 365
rect 36892 361 36946 365
rect 36686 356 36706 361
rect 36926 356 36946 361
rect 36696 341 36698 356
rect 36524 261 36528 329
rect 36592 305 36596 341
rect 36690 331 36698 341
rect 36706 331 36707 351
rect 36696 315 36698 331
rect 36717 322 36720 356
rect 36739 331 36740 351
rect 36749 331 36756 341
rect 36876 331 36883 341
rect 36892 331 36893 351
rect 36912 322 36915 356
rect 36925 331 36926 351
rect 36935 331 36942 341
rect 36706 315 36722 321
rect 36724 315 36740 321
rect 36892 315 36908 321
rect 36910 315 36926 321
rect 36986 315 36988 365
rect 36529 267 36565 295
rect 36529 261 36543 267
rect 36208 212 36219 213
rect 36053 183 36060 207
rect 36208 183 36218 212
rect 36299 207 36311 241
rect 36321 207 36341 241
rect 36044 103 36048 171
rect 36112 133 36116 183
rect 36112 98 36116 103
rect 35863 62 35868 96
rect 35892 62 35897 96
rect 36112 94 36150 98
rect 36112 79 36120 94
rect 36146 79 36150 94
rect 36234 94 36268 98
rect 36234 79 36238 94
rect 36264 79 36268 94
rect 36112 61 36154 79
rect 36230 61 36272 79
rect 36090 55 36176 61
rect 36208 55 36294 61
rect 36336 55 36340 207
rect 36366 183 36373 211
rect 36524 183 36528 251
rect 36533 233 36543 261
rect 36553 261 36567 267
rect 36592 261 36603 305
rect 37029 267 37040 305
rect 37067 267 37103 295
rect 37104 267 37108 395
rect 37255 378 37260 412
rect 37284 378 37289 412
rect 37290 400 37301 412
rect 37315 400 37326 412
rect 37327 395 37402 412
rect 37478 420 37531 421
rect 37541 420 37553 424
rect 37591 420 37603 424
rect 37613 420 37625 424
rect 37478 412 37520 420
rect 37478 395 37553 412
rect 37554 400 37565 412
rect 37579 400 37590 412
rect 37292 341 37296 395
rect 37327 378 37398 395
rect 37402 383 37410 395
rect 37470 383 37478 395
rect 37482 378 37516 395
rect 37519 378 37553 395
rect 37360 371 37364 378
rect 36754 262 36804 264
rect 36828 262 36878 264
rect 36553 233 36573 261
rect 36592 233 36601 261
rect 36655 253 36689 261
rect 36634 246 36689 253
rect 36655 245 36689 246
rect 36757 253 36788 261
rect 36757 245 36791 253
rect 36592 213 36596 233
rect 36788 229 36791 245
rect 36655 228 36689 229
rect 36634 221 36689 228
rect 36757 221 36791 229
rect 36804 212 36806 262
rect 36844 253 36875 261
rect 36878 253 36880 262
rect 37067 261 37079 267
rect 36844 245 36880 253
rect 36943 253 36977 261
rect 36943 246 36998 253
rect 36943 245 36977 246
rect 36875 229 36880 245
rect 37069 233 37079 261
rect 37089 233 37109 267
rect 37292 261 37296 329
rect 37360 291 37364 341
rect 37360 251 37369 279
rect 37456 264 37466 291
rect 37415 262 37466 264
rect 37456 261 37467 262
rect 37423 253 37457 261
rect 37465 253 37467 261
rect 36844 221 36880 229
rect 36943 228 36977 229
rect 36943 221 36998 228
rect 36878 212 36880 221
rect 36524 103 36528 171
rect 36592 133 36596 183
rect 36646 159 36696 161
rect 36936 159 36986 161
rect 36696 143 36698 159
rect 36706 153 36722 159
rect 36724 153 36740 159
rect 36892 153 36908 159
rect 36910 153 36926 159
rect 36717 143 36740 152
rect 36892 143 36915 152
rect 36690 133 36698 143
rect 36696 109 36698 133
rect 36706 123 36707 143
rect 36717 118 36720 143
rect 36739 123 36740 143
rect 36749 133 36756 143
rect 36876 133 36883 143
rect 36892 123 36893 143
rect 36912 118 36915 143
rect 36925 123 36926 143
rect 36935 133 36942 143
rect 36706 109 36740 113
rect 36892 109 36926 113
rect 36986 109 36988 159
rect 36592 103 36634 104
rect 36998 103 37040 104
rect 36592 96 36596 103
rect 36487 62 36492 96
rect 36516 62 36521 96
rect 36559 79 36630 96
rect 37002 79 37036 96
rect 37039 79 37073 96
rect 36559 62 36634 79
rect 36592 61 36634 62
rect 36998 62 37073 79
rect 36998 61 37040 62
rect 36570 55 36656 61
rect 36976 55 37062 61
rect 37104 55 37108 233
rect 37292 183 37296 251
rect 37301 207 37311 241
rect 37321 213 37341 241
rect 37321 207 37335 213
rect 37360 207 37371 251
rect 37402 246 37478 253
rect 37511 251 37520 279
rect 37423 228 37457 246
rect 37465 228 37467 246
rect 37402 221 37478 228
rect 37465 213 37467 221
rect 37509 213 37520 251
rect 37584 241 37588 395
rect 37591 378 37596 412
rect 37620 378 37625 412
rect 37626 400 37637 412
rect 37840 395 37882 421
rect 38246 395 38288 421
rect 38503 420 38515 424
rect 38525 420 38537 424
rect 38575 420 38587 424
rect 38597 421 38609 424
rect 38767 421 38779 424
rect 38597 420 38650 421
rect 38608 412 38650 420
rect 38491 400 38502 412
rect 37772 341 37776 395
rect 37832 387 37878 395
rect 37832 383 37848 387
rect 37840 380 37848 383
rect 37874 380 37878 387
rect 37882 383 37890 395
rect 38238 383 38246 395
rect 38250 387 38284 395
rect 38250 380 38254 387
rect 38280 380 38284 387
rect 38288 383 38296 395
rect 37828 379 37894 380
rect 38234 379 38300 380
rect 37840 371 37844 379
rect 37894 365 37944 367
rect 38184 365 38234 367
rect 37934 361 37988 365
rect 38140 361 38194 365
rect 37934 356 37954 361
rect 38174 356 38194 361
rect 37944 341 37946 356
rect 37772 261 37776 329
rect 37840 305 37844 341
rect 37938 331 37946 341
rect 37954 331 37955 351
rect 37944 315 37946 331
rect 37965 322 37968 356
rect 37987 331 37988 351
rect 37997 331 38004 341
rect 38124 331 38131 341
rect 38140 331 38141 351
rect 38160 322 38163 356
rect 38173 331 38174 351
rect 38183 331 38190 341
rect 37954 315 37970 321
rect 37972 315 37988 321
rect 38140 315 38156 321
rect 38158 315 38174 321
rect 38234 315 38236 365
rect 37777 267 37813 295
rect 37777 261 37791 267
rect 37456 212 37467 213
rect 37301 183 37308 207
rect 37456 183 37466 212
rect 37547 207 37559 241
rect 37569 207 37589 241
rect 37292 103 37296 171
rect 37360 133 37364 183
rect 37360 98 37364 103
rect 37111 62 37116 96
rect 37140 62 37145 96
rect 37360 94 37398 98
rect 37360 79 37368 94
rect 37394 79 37398 94
rect 37482 94 37516 98
rect 37482 79 37486 94
rect 37512 79 37516 94
rect 37360 61 37402 79
rect 37478 61 37520 79
rect 37338 55 37424 61
rect 37456 55 37542 61
rect 37584 55 37588 207
rect 37614 183 37621 211
rect 37772 183 37776 251
rect 37781 233 37791 261
rect 37801 261 37815 267
rect 37840 261 37851 305
rect 38277 267 38288 305
rect 38315 267 38351 295
rect 38352 267 38356 395
rect 38503 378 38508 412
rect 38532 378 38537 412
rect 38538 400 38549 412
rect 38563 400 38574 412
rect 38575 395 38650 412
rect 38726 420 38779 421
rect 38789 420 38801 424
rect 38839 420 38851 424
rect 38861 420 38873 424
rect 38726 412 38768 420
rect 38726 395 38801 412
rect 38802 400 38813 412
rect 38827 400 38838 412
rect 38540 341 38544 395
rect 38575 378 38646 395
rect 38650 383 38658 395
rect 38718 383 38726 395
rect 38730 378 38764 395
rect 38767 378 38801 395
rect 38608 371 38612 378
rect 38002 262 38052 264
rect 38076 262 38126 264
rect 37801 233 37821 261
rect 37840 233 37849 261
rect 37903 253 37937 261
rect 37882 246 37937 253
rect 37903 245 37937 246
rect 38005 253 38036 261
rect 38005 245 38039 253
rect 37840 213 37844 233
rect 38036 229 38039 245
rect 37903 228 37937 229
rect 37882 221 37937 228
rect 38005 221 38039 229
rect 38052 212 38054 262
rect 38092 253 38123 261
rect 38126 253 38128 262
rect 38315 261 38327 267
rect 38092 245 38128 253
rect 38191 253 38225 261
rect 38191 246 38246 253
rect 38191 245 38225 246
rect 38123 229 38128 245
rect 38317 233 38327 261
rect 38337 233 38357 267
rect 38540 261 38544 329
rect 38608 291 38612 341
rect 38608 251 38617 279
rect 38704 264 38714 291
rect 38663 262 38714 264
rect 38704 261 38715 262
rect 38671 253 38705 261
rect 38713 253 38715 261
rect 38092 221 38128 229
rect 38191 228 38225 229
rect 38191 221 38246 228
rect 38126 212 38128 221
rect 37772 103 37776 171
rect 37840 133 37844 183
rect 37894 159 37944 161
rect 38184 159 38234 161
rect 37944 143 37946 159
rect 37954 153 37970 159
rect 37972 153 37988 159
rect 38140 153 38156 159
rect 38158 153 38174 159
rect 37965 143 37988 152
rect 38140 143 38163 152
rect 37938 133 37946 143
rect 37944 109 37946 133
rect 37954 123 37955 143
rect 37965 118 37968 143
rect 37987 123 37988 143
rect 37997 133 38004 143
rect 38124 133 38131 143
rect 38140 123 38141 143
rect 38160 118 38163 143
rect 38173 123 38174 143
rect 38183 133 38190 143
rect 37954 109 37988 113
rect 38140 109 38174 113
rect 38234 109 38236 159
rect 37840 103 37882 104
rect 38246 103 38288 104
rect 37840 96 37844 103
rect 37735 62 37740 96
rect 37764 62 37769 96
rect 37807 79 37878 96
rect 38250 79 38284 96
rect 38287 79 38321 96
rect 37807 62 37882 79
rect 37840 61 37882 62
rect 38246 62 38321 79
rect 38246 61 38288 62
rect 37818 55 37904 61
rect 38224 55 38310 61
rect 38352 55 38356 233
rect 38540 183 38544 251
rect 38549 207 38559 241
rect 38569 213 38589 241
rect 38569 207 38583 213
rect 38608 207 38619 251
rect 38650 246 38726 253
rect 38759 251 38768 279
rect 38671 228 38705 246
rect 38713 228 38715 246
rect 38650 221 38726 228
rect 38713 213 38715 221
rect 38757 213 38768 251
rect 38832 241 38836 395
rect 38839 378 38844 412
rect 38868 378 38873 412
rect 38874 400 38885 412
rect 39088 395 39130 421
rect 39494 395 39536 421
rect 39751 420 39763 424
rect 39773 420 39785 424
rect 39823 420 39835 424
rect 39845 421 39857 424
rect 40015 421 40027 424
rect 39845 420 39898 421
rect 39856 412 39898 420
rect 39739 400 39750 412
rect 39020 341 39024 395
rect 39080 387 39126 395
rect 39080 383 39096 387
rect 39088 380 39096 383
rect 39122 380 39126 387
rect 39130 383 39138 395
rect 39486 383 39494 395
rect 39498 387 39532 395
rect 39498 380 39502 387
rect 39528 380 39532 387
rect 39536 383 39544 395
rect 39076 379 39142 380
rect 39482 379 39548 380
rect 39088 371 39092 379
rect 39142 365 39192 367
rect 39432 365 39482 367
rect 39182 361 39236 365
rect 39388 361 39442 365
rect 39182 356 39202 361
rect 39422 356 39442 361
rect 39192 341 39194 356
rect 39020 261 39024 329
rect 39088 305 39092 341
rect 39186 331 39194 341
rect 39202 331 39203 351
rect 39192 315 39194 331
rect 39213 322 39216 356
rect 39235 331 39236 351
rect 39245 331 39252 341
rect 39372 331 39379 341
rect 39388 331 39389 351
rect 39408 322 39411 356
rect 39421 331 39422 351
rect 39431 331 39438 341
rect 39202 315 39218 321
rect 39220 315 39236 321
rect 39388 315 39404 321
rect 39406 315 39422 321
rect 39482 315 39484 365
rect 39025 267 39061 295
rect 39025 261 39039 267
rect 38704 212 38715 213
rect 38549 183 38556 207
rect 38704 183 38714 212
rect 38795 207 38807 241
rect 38817 207 38837 241
rect 38540 103 38544 171
rect 38608 133 38612 183
rect 38608 98 38612 103
rect 38359 62 38364 96
rect 38388 62 38393 96
rect 38608 94 38646 98
rect 38608 79 38616 94
rect 38642 79 38646 94
rect 38730 94 38764 98
rect 38730 79 38734 94
rect 38760 79 38764 94
rect 38608 61 38650 79
rect 38726 61 38768 79
rect 38586 55 38672 61
rect 38704 55 38790 61
rect 38832 55 38836 207
rect 38862 183 38869 211
rect 39020 183 39024 251
rect 39029 233 39039 261
rect 39049 261 39063 267
rect 39088 261 39099 305
rect 39525 267 39536 305
rect 39563 267 39599 295
rect 39600 267 39604 395
rect 39751 378 39756 412
rect 39780 378 39785 412
rect 39786 400 39797 412
rect 39811 400 39822 412
rect 39823 395 39898 412
rect 39974 420 40027 421
rect 40037 420 40049 424
rect 40087 420 40099 424
rect 40109 420 40121 424
rect 39974 412 40016 420
rect 39974 395 40049 412
rect 40050 400 40061 412
rect 40075 400 40086 412
rect 39788 341 39792 395
rect 39823 378 39894 395
rect 39898 383 39906 395
rect 39966 383 39974 395
rect 39978 378 40012 395
rect 40015 378 40049 395
rect 39856 371 39860 378
rect 39250 262 39300 264
rect 39324 262 39374 264
rect 39049 233 39069 261
rect 39088 233 39097 261
rect 39151 253 39185 261
rect 39130 246 39185 253
rect 39151 245 39185 246
rect 39253 253 39284 261
rect 39253 245 39287 253
rect 39088 213 39092 233
rect 39284 229 39287 245
rect 39151 228 39185 229
rect 39130 221 39185 228
rect 39253 221 39287 229
rect 39300 212 39302 262
rect 39340 253 39371 261
rect 39374 253 39376 262
rect 39563 261 39575 267
rect 39340 245 39376 253
rect 39439 253 39473 261
rect 39439 246 39494 253
rect 39439 245 39473 246
rect 39371 229 39376 245
rect 39565 233 39575 261
rect 39585 233 39605 267
rect 39788 261 39792 329
rect 39856 291 39860 341
rect 39856 251 39865 279
rect 39952 264 39962 291
rect 39911 262 39962 264
rect 39952 261 39963 262
rect 39919 253 39953 261
rect 39961 253 39963 261
rect 39340 221 39376 229
rect 39439 228 39473 229
rect 39439 221 39494 228
rect 39374 212 39376 221
rect 39020 103 39024 171
rect 39088 133 39092 183
rect 39142 159 39192 161
rect 39432 159 39482 161
rect 39192 143 39194 159
rect 39202 153 39218 159
rect 39220 153 39236 159
rect 39388 153 39404 159
rect 39406 153 39422 159
rect 39213 143 39236 152
rect 39388 143 39411 152
rect 39186 133 39194 143
rect 39192 109 39194 133
rect 39202 123 39203 143
rect 39213 118 39216 143
rect 39235 123 39236 143
rect 39245 133 39252 143
rect 39372 133 39379 143
rect 39388 123 39389 143
rect 39408 118 39411 143
rect 39421 123 39422 143
rect 39431 133 39438 143
rect 39202 109 39236 113
rect 39388 109 39422 113
rect 39482 109 39484 159
rect 39088 103 39130 104
rect 39494 103 39536 104
rect 39088 96 39092 103
rect 38983 62 38988 96
rect 39012 62 39017 96
rect 39055 79 39126 96
rect 39498 79 39532 96
rect 39535 79 39569 96
rect 39055 62 39130 79
rect 39088 61 39130 62
rect 39494 62 39569 79
rect 39494 61 39536 62
rect 39066 55 39152 61
rect 39472 55 39558 61
rect 39600 55 39604 233
rect 39788 183 39792 251
rect 39797 207 39807 241
rect 39817 213 39837 241
rect 39817 207 39831 213
rect 39856 207 39867 251
rect 39898 246 39974 253
rect 40007 251 40016 279
rect 39919 228 39953 246
rect 39961 228 39963 246
rect 39898 221 39974 228
rect 39961 213 39963 221
rect 40005 213 40016 251
rect 40080 241 40084 395
rect 40087 378 40092 412
rect 40116 378 40121 412
rect 40122 400 40133 412
rect 40336 395 40378 421
rect 40742 395 40784 421
rect 40999 420 41011 424
rect 41021 420 41033 424
rect 41071 420 41083 424
rect 41093 421 41105 424
rect 41263 421 41275 424
rect 41093 420 41146 421
rect 41104 412 41146 420
rect 40987 400 40998 412
rect 40268 341 40272 395
rect 40328 387 40374 395
rect 40328 383 40344 387
rect 40336 380 40344 383
rect 40370 380 40374 387
rect 40378 383 40386 395
rect 40734 383 40742 395
rect 40746 387 40780 395
rect 40746 380 40750 387
rect 40776 380 40780 387
rect 40784 383 40792 395
rect 40324 379 40390 380
rect 40730 379 40796 380
rect 40336 371 40340 379
rect 40390 365 40440 367
rect 40680 365 40730 367
rect 40430 361 40484 365
rect 40636 361 40690 365
rect 40430 356 40450 361
rect 40670 356 40690 361
rect 40440 341 40442 356
rect 40268 261 40272 329
rect 40336 305 40340 341
rect 40434 331 40442 341
rect 40450 331 40451 351
rect 40440 315 40442 331
rect 40461 322 40464 356
rect 40483 331 40484 351
rect 40493 331 40500 341
rect 40620 331 40627 341
rect 40636 331 40637 351
rect 40656 322 40659 356
rect 40669 331 40670 351
rect 40679 331 40686 341
rect 40450 315 40466 321
rect 40468 315 40484 321
rect 40636 315 40652 321
rect 40654 315 40670 321
rect 40730 315 40732 365
rect 40273 267 40309 295
rect 40273 261 40287 267
rect 39952 212 39963 213
rect 39797 183 39804 207
rect 39952 183 39962 212
rect 40043 207 40055 241
rect 40065 207 40085 241
rect 39788 103 39792 171
rect 39856 133 39860 183
rect 39856 98 39860 103
rect 39607 62 39612 96
rect 39636 62 39641 96
rect 39856 94 39894 98
rect 39856 79 39864 94
rect 39890 79 39894 94
rect 39978 94 40012 98
rect 39978 79 39982 94
rect 40008 79 40012 94
rect 39856 61 39898 79
rect 39974 61 40016 79
rect 39834 55 39920 61
rect 39952 55 40038 61
rect 40080 55 40084 207
rect 40110 183 40117 211
rect 40268 183 40272 251
rect 40277 233 40287 261
rect 40297 261 40311 267
rect 40336 261 40347 305
rect 40773 267 40784 305
rect 40811 267 40847 295
rect 40848 267 40852 395
rect 40999 378 41004 412
rect 41028 378 41033 412
rect 41034 400 41045 412
rect 41059 400 41070 412
rect 41071 395 41146 412
rect 41222 420 41275 421
rect 41285 420 41297 424
rect 41335 420 41347 424
rect 41357 420 41369 424
rect 41222 412 41264 420
rect 41222 395 41297 412
rect 41298 400 41309 412
rect 41323 400 41334 412
rect 41036 341 41040 395
rect 41071 378 41142 395
rect 41146 383 41154 395
rect 41214 383 41222 395
rect 41226 378 41260 395
rect 41263 378 41297 395
rect 41104 371 41108 378
rect 40498 262 40548 264
rect 40572 262 40622 264
rect 40297 233 40317 261
rect 40336 233 40345 261
rect 40399 253 40433 261
rect 40378 246 40433 253
rect 40399 245 40433 246
rect 40501 253 40532 261
rect 40501 245 40535 253
rect 40336 213 40340 233
rect 40532 229 40535 245
rect 40399 228 40433 229
rect 40378 221 40433 228
rect 40501 221 40535 229
rect 40548 212 40550 262
rect 40588 253 40619 261
rect 40622 253 40624 262
rect 40811 261 40823 267
rect 40588 245 40624 253
rect 40687 253 40721 261
rect 40687 246 40742 253
rect 40687 245 40721 246
rect 40619 229 40624 245
rect 40813 233 40823 261
rect 40833 233 40853 267
rect 41036 261 41040 329
rect 41104 291 41108 341
rect 41104 251 41113 279
rect 41200 264 41210 291
rect 41159 262 41210 264
rect 41200 261 41211 262
rect 41167 253 41201 261
rect 41209 253 41211 261
rect 40588 221 40624 229
rect 40687 228 40721 229
rect 40687 221 40742 228
rect 40622 212 40624 221
rect 40268 103 40272 171
rect 40336 133 40340 183
rect 40390 159 40440 161
rect 40680 159 40730 161
rect 40440 143 40442 159
rect 40450 153 40466 159
rect 40468 153 40484 159
rect 40636 153 40652 159
rect 40654 153 40670 159
rect 40461 143 40484 152
rect 40636 143 40659 152
rect 40434 133 40442 143
rect 40440 109 40442 133
rect 40450 123 40451 143
rect 40461 118 40464 143
rect 40483 123 40484 143
rect 40493 133 40500 143
rect 40620 133 40627 143
rect 40636 123 40637 143
rect 40656 118 40659 143
rect 40669 123 40670 143
rect 40679 133 40686 143
rect 40450 109 40484 113
rect 40636 109 40670 113
rect 40730 109 40732 159
rect 40336 103 40378 104
rect 40742 103 40784 104
rect 40336 96 40340 103
rect 40231 62 40236 96
rect 40260 62 40265 96
rect 40303 79 40374 96
rect 40746 79 40780 96
rect 40783 79 40817 96
rect 40303 62 40378 79
rect 40336 61 40378 62
rect 40742 62 40817 79
rect 40742 61 40784 62
rect 40320 55 40400 61
rect 40720 55 40806 61
rect 40848 55 40852 233
rect 41036 183 41040 251
rect 41045 207 41055 241
rect 41065 213 41085 241
rect 41065 207 41079 213
rect 41104 207 41115 251
rect 41146 246 41222 253
rect 41255 251 41264 279
rect 41167 228 41201 246
rect 41209 228 41211 246
rect 41146 221 41222 228
rect 41209 213 41211 221
rect 41253 213 41264 251
rect 41328 241 41332 395
rect 41335 378 41340 412
rect 41364 378 41369 412
rect 41370 400 41381 412
rect 41584 395 41626 421
rect 41990 395 42032 421
rect 42247 420 42259 424
rect 42269 420 42281 424
rect 42319 420 42331 424
rect 42341 421 42353 424
rect 42511 421 42523 424
rect 42341 420 42394 421
rect 42352 412 42394 420
rect 42235 400 42246 412
rect 41516 341 41520 395
rect 41576 387 41622 395
rect 41576 383 41592 387
rect 41584 380 41592 383
rect 41618 380 41622 387
rect 41626 383 41634 395
rect 41982 383 41990 395
rect 41994 387 42028 395
rect 41994 380 41998 387
rect 42024 380 42028 387
rect 42032 383 42040 395
rect 41572 379 41638 380
rect 41978 379 42044 380
rect 41584 371 41588 379
rect 41638 365 41688 367
rect 41928 365 41978 367
rect 41678 361 41732 365
rect 41884 361 41938 365
rect 41678 356 41698 361
rect 41918 356 41938 361
rect 41688 341 41690 356
rect 41516 261 41520 329
rect 41584 305 41588 341
rect 41682 331 41690 341
rect 41698 331 41699 351
rect 41688 315 41690 331
rect 41709 322 41712 356
rect 41731 331 41732 351
rect 41741 331 41748 341
rect 41868 331 41875 341
rect 41884 331 41885 351
rect 41904 322 41907 356
rect 41917 331 41918 351
rect 41927 331 41934 341
rect 41698 315 41714 321
rect 41716 315 41732 321
rect 41884 315 41900 321
rect 41902 315 41918 321
rect 41978 315 41980 365
rect 41521 267 41557 295
rect 41521 261 41535 267
rect 41200 212 41211 213
rect 41045 183 41052 207
rect 41200 183 41210 212
rect 41291 207 41303 241
rect 41313 207 41333 241
rect 41036 103 41040 171
rect 41104 133 41108 183
rect 41104 98 41108 103
rect 40855 62 40860 96
rect 40884 62 40889 96
rect 41104 94 41142 98
rect 41104 79 41112 94
rect 41138 79 41142 94
rect 41226 94 41260 98
rect 41226 79 41230 94
rect 41256 79 41260 94
rect 41104 61 41146 79
rect 41222 61 41264 79
rect 41082 55 41168 61
rect 41200 55 41286 61
rect 41328 55 41332 207
rect 41358 183 41365 211
rect 41516 183 41520 251
rect 41525 233 41535 261
rect 41545 261 41559 267
rect 41584 261 41595 305
rect 42021 267 42032 305
rect 42059 267 42095 295
rect 42096 267 42100 395
rect 42247 378 42252 412
rect 42276 378 42281 412
rect 42282 400 42293 412
rect 42307 400 42318 412
rect 42319 395 42394 412
rect 42470 420 42523 421
rect 42533 420 42545 424
rect 42583 420 42595 424
rect 42605 420 42617 424
rect 42470 412 42512 420
rect 42470 395 42545 412
rect 42546 400 42557 412
rect 42571 400 42582 412
rect 42284 341 42288 395
rect 42319 378 42390 395
rect 42394 383 42402 395
rect 42462 383 42470 395
rect 42474 378 42508 395
rect 42511 378 42545 395
rect 42352 371 42356 378
rect 41746 262 41796 264
rect 41820 262 41870 264
rect 41545 233 41565 261
rect 41584 233 41593 261
rect 41647 253 41681 261
rect 41626 246 41681 253
rect 41647 245 41681 246
rect 41749 253 41780 261
rect 41749 245 41783 253
rect 41584 213 41588 233
rect 41780 229 41783 245
rect 41647 228 41681 229
rect 41626 221 41681 228
rect 41749 221 41783 229
rect 41796 212 41798 262
rect 41836 253 41867 261
rect 41870 253 41872 262
rect 42059 261 42071 267
rect 41836 245 41872 253
rect 41935 253 41969 261
rect 41935 246 41990 253
rect 41935 245 41969 246
rect 41867 229 41872 245
rect 42061 233 42071 261
rect 42081 233 42101 267
rect 42284 261 42288 329
rect 42352 291 42356 341
rect 42352 251 42361 279
rect 42448 264 42458 291
rect 42407 262 42458 264
rect 42448 261 42459 262
rect 42415 253 42449 261
rect 42457 253 42459 261
rect 41836 221 41872 229
rect 41935 228 41969 229
rect 41935 221 41990 228
rect 41870 212 41872 221
rect 41516 103 41520 171
rect 41584 133 41588 183
rect 41638 159 41688 161
rect 41928 159 41978 161
rect 41688 143 41690 159
rect 41698 153 41714 159
rect 41716 153 41732 159
rect 41884 153 41900 159
rect 41902 153 41918 159
rect 41709 143 41732 152
rect 41884 143 41907 152
rect 41682 133 41690 143
rect 41688 109 41690 133
rect 41698 123 41699 143
rect 41709 118 41712 143
rect 41731 123 41732 143
rect 41741 133 41748 143
rect 41868 133 41875 143
rect 41884 123 41885 143
rect 41904 118 41907 143
rect 41917 123 41918 143
rect 41927 133 41934 143
rect 41698 109 41732 113
rect 41884 109 41918 113
rect 41978 109 41980 159
rect 41584 103 41626 104
rect 41990 103 42032 104
rect 41584 96 41588 103
rect 41479 62 41484 96
rect 41508 62 41513 96
rect 41551 79 41622 96
rect 41994 79 42028 96
rect 42031 79 42065 96
rect 41551 62 41626 79
rect 41584 61 41626 62
rect 41990 62 42065 79
rect 41990 61 42032 62
rect 41562 55 41648 61
rect 41968 55 42054 61
rect 42096 55 42100 233
rect 42284 183 42288 251
rect 42293 207 42303 241
rect 42313 213 42333 241
rect 42313 207 42327 213
rect 42352 207 42363 251
rect 42394 246 42470 253
rect 42503 251 42512 279
rect 42415 228 42449 246
rect 42457 228 42459 246
rect 42394 221 42470 228
rect 42457 213 42459 221
rect 42501 213 42512 251
rect 42576 241 42580 395
rect 42583 378 42588 412
rect 42612 378 42617 412
rect 42618 400 42629 412
rect 42832 395 42874 421
rect 43238 395 43280 421
rect 43495 420 43507 424
rect 43517 420 43529 424
rect 43567 420 43579 424
rect 43589 421 43601 424
rect 43759 421 43771 424
rect 43589 420 43642 421
rect 43600 412 43642 420
rect 43483 400 43494 412
rect 42764 341 42768 395
rect 42824 387 42870 395
rect 42824 383 42840 387
rect 42832 380 42840 383
rect 42866 380 42870 387
rect 42874 383 42882 395
rect 43230 383 43238 395
rect 43242 387 43276 395
rect 43242 380 43246 387
rect 43272 380 43276 387
rect 43280 383 43288 395
rect 42820 379 42886 380
rect 43226 379 43292 380
rect 42832 371 42836 379
rect 42886 365 42936 367
rect 43176 365 43226 367
rect 42926 361 42980 365
rect 43132 361 43186 365
rect 42926 356 42946 361
rect 43166 356 43186 361
rect 42936 341 42938 356
rect 42764 261 42768 329
rect 42832 305 42836 341
rect 42930 331 42938 341
rect 42946 331 42947 351
rect 42936 315 42938 331
rect 42957 322 42960 356
rect 42979 331 42980 351
rect 42989 331 42996 341
rect 43116 331 43123 341
rect 43132 331 43133 351
rect 43152 322 43155 356
rect 43165 331 43166 351
rect 43175 331 43182 341
rect 42946 315 42962 321
rect 42964 315 42980 321
rect 43132 315 43148 321
rect 43150 315 43166 321
rect 43226 315 43228 365
rect 42769 267 42805 295
rect 42769 261 42783 267
rect 42448 212 42459 213
rect 42293 183 42300 207
rect 42448 183 42458 212
rect 42539 207 42551 241
rect 42561 207 42581 241
rect 42284 103 42288 171
rect 42352 133 42356 183
rect 42352 98 42356 103
rect 42103 62 42108 96
rect 42132 62 42137 96
rect 42352 94 42390 98
rect 42352 79 42360 94
rect 42386 79 42390 94
rect 42474 94 42508 98
rect 42474 79 42478 94
rect 42504 79 42508 94
rect 42352 61 42394 79
rect 42470 61 42512 79
rect 42330 55 42416 61
rect 42448 55 42534 61
rect 42576 55 42580 207
rect 42606 183 42613 211
rect 42764 183 42768 251
rect 42773 233 42783 261
rect 42793 261 42807 267
rect 42832 261 42843 305
rect 43269 267 43280 305
rect 43307 267 43343 295
rect 43344 267 43348 395
rect 43495 378 43500 412
rect 43524 378 43529 412
rect 43530 400 43541 412
rect 43555 400 43566 412
rect 43567 395 43642 412
rect 43718 420 43771 421
rect 43781 420 43793 424
rect 43831 420 43843 424
rect 43853 420 43865 424
rect 43718 412 43760 420
rect 43718 395 43793 412
rect 43794 400 43805 412
rect 43819 400 43830 412
rect 43532 341 43536 395
rect 43567 378 43638 395
rect 43642 383 43650 395
rect 43710 383 43718 395
rect 43722 378 43756 395
rect 43759 378 43793 395
rect 43600 371 43604 378
rect 42994 262 43044 264
rect 43068 262 43118 264
rect 42793 233 42813 261
rect 42832 233 42841 261
rect 42895 253 42929 261
rect 42874 246 42929 253
rect 42895 245 42929 246
rect 42997 253 43028 261
rect 42997 245 43031 253
rect 42832 213 42836 233
rect 43028 229 43031 245
rect 42895 228 42929 229
rect 42874 221 42929 228
rect 42997 221 43031 229
rect 43044 212 43046 262
rect 43084 253 43115 261
rect 43118 253 43120 262
rect 43307 261 43319 267
rect 43084 245 43120 253
rect 43183 253 43217 261
rect 43183 246 43238 253
rect 43183 245 43217 246
rect 43115 229 43120 245
rect 43309 233 43319 261
rect 43329 233 43349 267
rect 43532 261 43536 329
rect 43600 291 43604 341
rect 43600 251 43609 279
rect 43696 264 43706 291
rect 43655 262 43706 264
rect 43696 261 43707 262
rect 43663 253 43697 261
rect 43705 253 43707 261
rect 43084 221 43120 229
rect 43183 228 43217 229
rect 43183 221 43238 228
rect 43118 212 43120 221
rect 42764 103 42768 171
rect 42832 133 42836 183
rect 42886 159 42936 161
rect 43176 159 43226 161
rect 42936 143 42938 159
rect 42946 153 42962 159
rect 42964 153 42980 159
rect 43132 153 43148 159
rect 43150 153 43166 159
rect 42957 143 42980 152
rect 43132 143 43155 152
rect 42930 133 42938 143
rect 42936 109 42938 133
rect 42946 123 42947 143
rect 42957 118 42960 143
rect 42979 123 42980 143
rect 42989 133 42996 143
rect 43116 133 43123 143
rect 43132 123 43133 143
rect 43152 118 43155 143
rect 43165 123 43166 143
rect 43175 133 43182 143
rect 42946 109 42980 113
rect 43132 109 43166 113
rect 43226 109 43228 159
rect 42832 103 42874 104
rect 43238 103 43280 104
rect 42832 96 42836 103
rect 42727 62 42732 96
rect 42756 62 42761 96
rect 42799 79 42870 96
rect 43242 79 43276 96
rect 43279 79 43313 96
rect 42799 62 42874 79
rect 42832 61 42874 62
rect 43238 62 43313 79
rect 43238 61 43280 62
rect 42810 55 42896 61
rect 43216 55 43302 61
rect 43344 55 43348 233
rect 43532 183 43536 251
rect 43541 207 43551 241
rect 43561 213 43581 241
rect 43561 207 43575 213
rect 43600 207 43611 251
rect 43642 246 43718 253
rect 43751 251 43760 279
rect 43663 228 43697 246
rect 43705 228 43707 246
rect 43642 221 43718 228
rect 43705 213 43707 221
rect 43749 213 43760 251
rect 43824 241 43828 395
rect 43831 378 43836 412
rect 43860 378 43865 412
rect 43866 400 43877 412
rect 44080 395 44122 421
rect 44486 395 44528 421
rect 44743 420 44755 424
rect 44765 420 44777 424
rect 44815 420 44827 424
rect 44837 421 44849 424
rect 45007 421 45019 424
rect 44837 420 44890 421
rect 44848 412 44890 420
rect 44731 400 44742 412
rect 44012 341 44016 395
rect 44072 387 44118 395
rect 44072 383 44088 387
rect 44080 380 44088 383
rect 44114 380 44118 387
rect 44122 383 44130 395
rect 44478 383 44486 395
rect 44490 387 44524 395
rect 44490 380 44494 387
rect 44520 380 44524 387
rect 44528 383 44536 395
rect 44068 379 44134 380
rect 44474 379 44540 380
rect 44080 371 44084 379
rect 44134 365 44184 367
rect 44424 365 44474 367
rect 44174 361 44228 365
rect 44380 361 44434 365
rect 44174 356 44194 361
rect 44414 356 44434 361
rect 44184 341 44186 356
rect 44012 261 44016 329
rect 44080 305 44084 341
rect 44178 331 44186 341
rect 44194 331 44195 351
rect 44184 315 44186 331
rect 44205 322 44208 356
rect 44227 331 44228 351
rect 44237 331 44244 341
rect 44364 331 44371 341
rect 44380 331 44381 351
rect 44400 322 44403 356
rect 44413 331 44414 351
rect 44423 331 44430 341
rect 44194 315 44210 321
rect 44212 315 44228 321
rect 44380 315 44396 321
rect 44398 315 44414 321
rect 44474 315 44476 365
rect 44017 267 44053 295
rect 44017 261 44031 267
rect 43696 212 43707 213
rect 43541 183 43548 207
rect 43696 183 43706 212
rect 43787 207 43799 241
rect 43809 207 43829 241
rect 43532 103 43536 171
rect 43600 133 43604 183
rect 43600 98 43604 103
rect 43351 62 43356 96
rect 43380 62 43385 96
rect 43600 94 43638 98
rect 43600 79 43608 94
rect 43634 79 43638 94
rect 43722 94 43756 98
rect 43722 79 43726 94
rect 43752 79 43756 94
rect 43600 61 43642 79
rect 43718 61 43760 79
rect 43578 55 43664 61
rect 43696 55 43782 61
rect 43824 55 43828 207
rect 43854 183 43861 211
rect 44012 183 44016 251
rect 44021 233 44031 261
rect 44041 261 44055 267
rect 44080 261 44091 305
rect 44517 267 44528 305
rect 44555 267 44591 295
rect 44592 267 44596 395
rect 44743 378 44748 412
rect 44772 378 44777 412
rect 44778 400 44789 412
rect 44803 400 44814 412
rect 44815 395 44890 412
rect 44966 420 45019 421
rect 45029 420 45041 424
rect 45079 420 45091 424
rect 45101 420 45113 424
rect 44966 412 45008 420
rect 44966 395 45041 412
rect 45042 400 45053 412
rect 45067 400 45078 412
rect 44780 341 44784 395
rect 44815 378 44886 395
rect 44890 383 44898 395
rect 44958 383 44966 395
rect 44970 378 45004 395
rect 45007 378 45041 395
rect 44848 371 44852 378
rect 44242 262 44292 264
rect 44316 262 44366 264
rect 44041 233 44061 261
rect 44080 233 44089 261
rect 44143 253 44177 261
rect 44122 246 44177 253
rect 44143 245 44177 246
rect 44245 253 44276 261
rect 44245 245 44279 253
rect 44080 213 44084 233
rect 44276 229 44279 245
rect 44143 228 44177 229
rect 44122 221 44177 228
rect 44245 221 44279 229
rect 44292 212 44294 262
rect 44332 253 44363 261
rect 44366 253 44368 262
rect 44555 261 44567 267
rect 44332 245 44368 253
rect 44431 253 44465 261
rect 44431 246 44486 253
rect 44431 245 44465 246
rect 44363 229 44368 245
rect 44557 233 44567 261
rect 44577 233 44597 267
rect 44780 261 44784 329
rect 44848 291 44852 341
rect 44848 251 44857 279
rect 44944 264 44954 291
rect 44903 262 44954 264
rect 44944 261 44955 262
rect 44911 253 44945 261
rect 44953 253 44955 261
rect 44332 221 44368 229
rect 44431 228 44465 229
rect 44431 221 44486 228
rect 44366 212 44368 221
rect 44012 103 44016 171
rect 44080 133 44084 183
rect 44134 159 44184 161
rect 44424 159 44474 161
rect 44184 143 44186 159
rect 44194 153 44210 159
rect 44212 153 44228 159
rect 44380 153 44396 159
rect 44398 153 44414 159
rect 44205 143 44228 152
rect 44380 143 44403 152
rect 44178 133 44186 143
rect 44184 109 44186 133
rect 44194 123 44195 143
rect 44205 118 44208 143
rect 44227 123 44228 143
rect 44237 133 44244 143
rect 44364 133 44371 143
rect 44380 123 44381 143
rect 44400 118 44403 143
rect 44413 123 44414 143
rect 44423 133 44430 143
rect 44194 109 44228 113
rect 44380 109 44414 113
rect 44474 109 44476 159
rect 44080 103 44122 104
rect 44486 103 44528 104
rect 44080 96 44084 103
rect 43975 62 43980 96
rect 44004 62 44009 96
rect 44047 79 44118 96
rect 44490 79 44524 96
rect 44527 79 44561 96
rect 44047 62 44122 79
rect 44080 61 44122 62
rect 44486 62 44561 79
rect 44486 61 44528 62
rect 44058 55 44144 61
rect 44464 55 44550 61
rect 44592 55 44596 233
rect 44780 183 44784 251
rect 44789 207 44799 241
rect 44809 213 44829 241
rect 44809 207 44823 213
rect 44848 207 44859 251
rect 44890 246 44966 253
rect 44999 251 45008 279
rect 44911 228 44945 246
rect 44953 228 44955 246
rect 44890 221 44966 228
rect 44953 213 44955 221
rect 44997 213 45008 251
rect 45072 241 45076 395
rect 45079 378 45084 412
rect 45108 378 45113 412
rect 45114 400 45125 412
rect 45328 395 45370 421
rect 45734 395 45776 421
rect 45991 420 46003 424
rect 46013 420 46025 424
rect 46063 420 46075 424
rect 46085 421 46097 424
rect 46255 421 46267 424
rect 46085 420 46138 421
rect 46096 412 46138 420
rect 45979 400 45990 412
rect 45260 341 45264 395
rect 45320 387 45366 395
rect 45320 383 45336 387
rect 45328 380 45336 383
rect 45362 380 45366 387
rect 45370 383 45378 395
rect 45726 383 45734 395
rect 45738 387 45772 395
rect 45738 380 45742 387
rect 45768 380 45772 387
rect 45776 383 45784 395
rect 45316 379 45382 380
rect 45722 379 45788 380
rect 45328 371 45332 379
rect 45382 365 45432 367
rect 45672 365 45722 367
rect 45422 361 45476 365
rect 45628 361 45682 365
rect 45422 356 45442 361
rect 45662 356 45682 361
rect 45432 341 45434 356
rect 45260 261 45264 329
rect 45328 305 45332 341
rect 45426 331 45434 341
rect 45442 331 45443 351
rect 45432 315 45434 331
rect 45453 322 45456 356
rect 45475 331 45476 351
rect 45485 331 45492 341
rect 45612 331 45619 341
rect 45628 331 45629 351
rect 45648 322 45651 356
rect 45661 331 45662 351
rect 45671 331 45678 341
rect 45442 315 45458 321
rect 45460 315 45476 321
rect 45628 315 45644 321
rect 45646 315 45662 321
rect 45722 315 45724 365
rect 45265 267 45301 295
rect 45265 261 45279 267
rect 44944 212 44955 213
rect 44789 183 44796 207
rect 44944 183 44954 212
rect 45035 207 45047 241
rect 45057 207 45077 241
rect 44780 103 44784 171
rect 44848 133 44852 183
rect 44848 98 44852 103
rect 44599 62 44604 96
rect 44628 62 44633 96
rect 44848 94 44886 98
rect 44848 79 44856 94
rect 44882 79 44886 94
rect 44970 94 45004 98
rect 44970 79 44974 94
rect 45000 79 45004 94
rect 44848 61 44890 79
rect 44966 61 45008 79
rect 44826 55 44912 61
rect 44944 55 45030 61
rect 45072 55 45076 207
rect 45102 183 45109 211
rect 45260 183 45264 251
rect 45269 233 45279 261
rect 45289 261 45303 267
rect 45328 261 45339 305
rect 45765 267 45776 305
rect 45803 267 45839 295
rect 45840 267 45844 395
rect 45991 378 45996 412
rect 46020 378 46025 412
rect 46026 400 46037 412
rect 46051 400 46062 412
rect 46063 395 46138 412
rect 46214 420 46267 421
rect 46277 420 46289 424
rect 46327 420 46339 424
rect 46349 420 46361 424
rect 46214 412 46256 420
rect 46214 395 46289 412
rect 46290 400 46301 412
rect 46315 400 46326 412
rect 46028 341 46032 395
rect 46063 378 46134 395
rect 46138 383 46146 395
rect 46206 383 46214 395
rect 46218 378 46252 395
rect 46255 378 46289 395
rect 46096 371 46100 378
rect 45490 262 45540 264
rect 45564 262 45614 264
rect 45289 233 45309 261
rect 45328 233 45337 261
rect 45391 253 45425 261
rect 45370 246 45425 253
rect 45391 245 45425 246
rect 45493 253 45524 261
rect 45493 245 45527 253
rect 45328 213 45332 233
rect 45524 229 45527 245
rect 45391 228 45425 229
rect 45370 221 45425 228
rect 45493 221 45527 229
rect 45540 212 45542 262
rect 45580 253 45611 261
rect 45614 253 45616 262
rect 45803 261 45815 267
rect 45580 245 45616 253
rect 45679 253 45713 261
rect 45679 246 45734 253
rect 45679 245 45713 246
rect 45611 229 45616 245
rect 45805 233 45815 261
rect 45825 233 45845 267
rect 46028 261 46032 329
rect 46096 291 46100 341
rect 46096 251 46105 279
rect 46192 264 46202 291
rect 46151 262 46202 264
rect 46192 261 46203 262
rect 46159 253 46193 261
rect 46201 253 46203 261
rect 45580 221 45616 229
rect 45679 228 45713 229
rect 45679 221 45734 228
rect 45614 212 45616 221
rect 45260 103 45264 171
rect 45328 133 45332 183
rect 45382 159 45432 161
rect 45672 159 45722 161
rect 45432 143 45434 159
rect 45442 153 45458 159
rect 45460 153 45476 159
rect 45628 153 45644 159
rect 45646 153 45662 159
rect 45453 143 45476 152
rect 45628 143 45651 152
rect 45426 133 45434 143
rect 45432 109 45434 133
rect 45442 123 45443 143
rect 45453 118 45456 143
rect 45475 123 45476 143
rect 45485 133 45492 143
rect 45612 133 45619 143
rect 45628 123 45629 143
rect 45648 118 45651 143
rect 45661 123 45662 143
rect 45671 133 45678 143
rect 45442 109 45476 113
rect 45628 109 45662 113
rect 45722 109 45724 159
rect 45328 103 45370 104
rect 45734 103 45776 104
rect 45328 96 45332 103
rect 45223 62 45228 96
rect 45252 62 45257 96
rect 45295 79 45366 96
rect 45738 79 45772 96
rect 45775 79 45809 96
rect 45295 62 45370 79
rect 45328 61 45370 62
rect 45734 62 45809 79
rect 45734 61 45776 62
rect 45306 55 45392 61
rect 45712 55 45798 61
rect 45840 55 45844 233
rect 46028 183 46032 251
rect 46037 207 46047 241
rect 46057 213 46077 241
rect 46057 207 46071 213
rect 46096 207 46107 251
rect 46138 246 46214 253
rect 46247 251 46256 279
rect 46159 228 46193 246
rect 46201 228 46203 246
rect 46138 221 46214 228
rect 46201 213 46203 221
rect 46245 213 46256 251
rect 46320 241 46324 395
rect 46327 378 46332 412
rect 46356 378 46361 412
rect 46362 400 46373 412
rect 46576 395 46618 421
rect 46982 395 47024 421
rect 47239 420 47251 424
rect 47261 420 47273 424
rect 47311 420 47323 424
rect 47333 421 47345 424
rect 47503 421 47515 424
rect 47333 420 47386 421
rect 47344 412 47386 420
rect 47227 400 47238 412
rect 46508 341 46512 395
rect 46568 387 46614 395
rect 46568 383 46584 387
rect 46576 380 46584 383
rect 46610 380 46614 387
rect 46618 383 46626 395
rect 46974 383 46982 395
rect 46986 387 47020 395
rect 46986 380 46990 387
rect 47016 380 47020 387
rect 47024 383 47032 395
rect 46564 379 46630 380
rect 46970 379 47036 380
rect 46576 371 46580 379
rect 46630 365 46680 367
rect 46920 365 46970 367
rect 46670 361 46724 365
rect 46876 361 46930 365
rect 46670 356 46690 361
rect 46910 356 46930 361
rect 46680 341 46682 356
rect 46508 261 46512 329
rect 46576 305 46580 341
rect 46674 331 46682 341
rect 46690 331 46691 351
rect 46680 315 46682 331
rect 46701 322 46704 356
rect 46723 331 46724 351
rect 46733 331 46740 341
rect 46860 331 46867 341
rect 46876 331 46877 351
rect 46896 322 46899 356
rect 46909 331 46910 351
rect 46919 331 46926 341
rect 46690 315 46706 321
rect 46708 315 46724 321
rect 46876 315 46892 321
rect 46894 315 46910 321
rect 46970 315 46972 365
rect 46513 267 46549 295
rect 46513 261 46527 267
rect 46192 212 46203 213
rect 46037 183 46044 207
rect 46192 183 46202 212
rect 46283 207 46295 241
rect 46305 207 46325 241
rect 46028 103 46032 171
rect 46096 133 46100 183
rect 46096 98 46100 103
rect 45847 62 45852 96
rect 45876 62 45881 96
rect 46096 94 46134 98
rect 46096 79 46104 94
rect 46130 79 46134 94
rect 46218 94 46252 98
rect 46218 79 46222 94
rect 46248 79 46252 94
rect 46096 61 46138 79
rect 46214 61 46256 79
rect 46074 55 46160 61
rect 46192 55 46278 61
rect 46320 55 46324 207
rect 46350 183 46357 211
rect 46508 183 46512 251
rect 46517 233 46527 261
rect 46537 261 46551 267
rect 46576 261 46587 305
rect 47013 267 47024 305
rect 47051 267 47087 295
rect 47088 267 47092 395
rect 47239 378 47244 412
rect 47268 378 47273 412
rect 47274 400 47285 412
rect 47299 400 47310 412
rect 47311 395 47386 412
rect 47462 420 47515 421
rect 47525 420 47537 424
rect 47575 420 47587 424
rect 47597 420 47609 424
rect 47462 412 47504 420
rect 47462 395 47537 412
rect 47538 400 47549 412
rect 47563 400 47574 412
rect 47276 341 47280 395
rect 47311 378 47382 395
rect 47386 383 47394 395
rect 47454 383 47462 395
rect 47466 378 47500 395
rect 47503 378 47537 395
rect 47344 371 47348 378
rect 46738 262 46788 264
rect 46812 262 46862 264
rect 46537 233 46557 261
rect 46576 233 46585 261
rect 46639 253 46673 261
rect 46618 246 46673 253
rect 46639 245 46673 246
rect 46741 253 46772 261
rect 46741 245 46775 253
rect 46576 213 46580 233
rect 46772 229 46775 245
rect 46639 228 46673 229
rect 46618 221 46673 228
rect 46741 221 46775 229
rect 46788 212 46790 262
rect 46828 253 46859 261
rect 46862 253 46864 262
rect 47051 261 47063 267
rect 46828 245 46864 253
rect 46927 253 46961 261
rect 46927 246 46982 253
rect 46927 245 46961 246
rect 46859 229 46864 245
rect 47053 233 47063 261
rect 47073 233 47093 267
rect 47276 261 47280 329
rect 47344 291 47348 341
rect 47344 251 47353 279
rect 47440 264 47450 291
rect 47399 262 47450 264
rect 47440 261 47451 262
rect 47407 253 47441 261
rect 47449 253 47451 261
rect 46828 221 46864 229
rect 46927 228 46961 229
rect 46927 221 46982 228
rect 46862 212 46864 221
rect 46508 103 46512 171
rect 46576 133 46580 183
rect 46630 159 46680 161
rect 46920 159 46970 161
rect 46680 143 46682 159
rect 46690 153 46706 159
rect 46708 153 46724 159
rect 46876 153 46892 159
rect 46894 153 46910 159
rect 46701 143 46724 152
rect 46876 143 46899 152
rect 46674 133 46682 143
rect 46680 109 46682 133
rect 46690 123 46691 143
rect 46701 118 46704 143
rect 46723 123 46724 143
rect 46733 133 46740 143
rect 46860 133 46867 143
rect 46876 123 46877 143
rect 46896 118 46899 143
rect 46909 123 46910 143
rect 46919 133 46926 143
rect 46690 109 46724 113
rect 46876 109 46910 113
rect 46970 109 46972 159
rect 46576 103 46618 104
rect 46982 103 47024 104
rect 46576 96 46580 103
rect 46471 62 46476 96
rect 46500 62 46505 96
rect 46543 79 46614 96
rect 46986 79 47020 96
rect 47023 79 47057 96
rect 46543 62 46618 79
rect 46576 61 46618 62
rect 46982 62 47057 79
rect 46982 61 47024 62
rect 46554 55 46640 61
rect 46960 55 47046 61
rect 47088 55 47092 233
rect 47276 183 47280 251
rect 47285 207 47295 241
rect 47305 213 47325 241
rect 47305 207 47319 213
rect 47344 207 47355 251
rect 47386 246 47462 253
rect 47495 251 47504 279
rect 47407 228 47441 246
rect 47449 228 47451 246
rect 47386 221 47462 228
rect 47449 213 47451 221
rect 47493 213 47504 251
rect 47568 241 47572 395
rect 47575 378 47580 412
rect 47604 378 47609 412
rect 47610 400 47621 412
rect 47824 395 47866 421
rect 48230 395 48272 421
rect 48487 420 48499 424
rect 48509 420 48521 424
rect 48559 420 48571 424
rect 48581 421 48593 424
rect 48751 421 48763 424
rect 48581 420 48634 421
rect 48592 412 48634 420
rect 48475 400 48486 412
rect 47756 341 47760 395
rect 47816 387 47862 395
rect 47816 383 47832 387
rect 47824 380 47832 383
rect 47858 380 47862 387
rect 47866 383 47874 395
rect 48222 383 48230 395
rect 48234 387 48268 395
rect 48234 380 48238 387
rect 48264 380 48268 387
rect 48272 383 48280 395
rect 47812 379 47878 380
rect 48218 379 48284 380
rect 47824 371 47828 379
rect 47878 365 47928 367
rect 48168 365 48218 367
rect 47918 361 47972 365
rect 48124 361 48178 365
rect 47918 356 47938 361
rect 48158 356 48178 361
rect 47928 341 47930 356
rect 47756 261 47760 329
rect 47824 305 47828 341
rect 47922 331 47930 341
rect 47938 331 47939 351
rect 47928 315 47930 331
rect 47949 322 47952 356
rect 47971 331 47972 351
rect 47981 331 47988 341
rect 48108 331 48115 341
rect 48124 331 48125 351
rect 48144 322 48147 356
rect 48157 331 48158 351
rect 48167 331 48174 341
rect 47938 315 47954 321
rect 47956 315 47972 321
rect 48124 315 48140 321
rect 48142 315 48158 321
rect 48218 315 48220 365
rect 47761 267 47797 295
rect 47761 261 47775 267
rect 47440 212 47451 213
rect 47285 183 47292 207
rect 47440 183 47450 212
rect 47531 207 47543 241
rect 47553 207 47573 241
rect 47276 103 47280 171
rect 47344 133 47348 183
rect 47344 98 47348 103
rect 47095 62 47100 96
rect 47124 62 47129 96
rect 47344 94 47382 98
rect 47344 79 47352 94
rect 47378 79 47382 94
rect 47466 94 47500 98
rect 47466 79 47470 94
rect 47496 79 47500 94
rect 47344 61 47386 79
rect 47462 61 47504 79
rect 47322 55 47408 61
rect 47440 55 47526 61
rect 47568 55 47572 207
rect 47598 183 47605 211
rect 47756 183 47760 251
rect 47765 233 47775 261
rect 47785 261 47799 267
rect 47824 261 47835 305
rect 48261 267 48272 305
rect 48299 267 48335 295
rect 48336 267 48340 395
rect 48487 378 48492 412
rect 48516 378 48521 412
rect 48522 400 48533 412
rect 48547 400 48558 412
rect 48559 395 48634 412
rect 48710 420 48763 421
rect 48773 420 48785 424
rect 48823 420 48835 424
rect 48845 420 48857 424
rect 48710 412 48752 420
rect 48710 395 48785 412
rect 48786 400 48797 412
rect 48811 400 48822 412
rect 48524 341 48528 395
rect 48559 378 48630 395
rect 48634 383 48642 395
rect 48702 383 48710 395
rect 48714 378 48748 395
rect 48751 378 48785 395
rect 48592 371 48596 378
rect 47986 262 48036 264
rect 48060 262 48110 264
rect 47785 233 47805 261
rect 47824 233 47833 261
rect 47887 253 47921 261
rect 47866 246 47921 253
rect 47887 245 47921 246
rect 47989 253 48020 261
rect 47989 245 48023 253
rect 47824 213 47828 233
rect 48020 229 48023 245
rect 47887 228 47921 229
rect 47866 221 47921 228
rect 47989 221 48023 229
rect 48036 212 48038 262
rect 48076 253 48107 261
rect 48110 253 48112 262
rect 48299 261 48311 267
rect 48076 245 48112 253
rect 48175 253 48209 261
rect 48175 246 48230 253
rect 48175 245 48209 246
rect 48107 229 48112 245
rect 48301 233 48311 261
rect 48321 233 48341 267
rect 48524 261 48528 329
rect 48592 291 48596 341
rect 48592 251 48601 279
rect 48688 264 48698 291
rect 48647 262 48698 264
rect 48688 261 48699 262
rect 48655 253 48689 261
rect 48697 253 48699 261
rect 48076 221 48112 229
rect 48175 228 48209 229
rect 48175 221 48230 228
rect 48110 212 48112 221
rect 47756 103 47760 171
rect 47824 133 47828 183
rect 47878 159 47928 161
rect 48168 159 48218 161
rect 47928 143 47930 159
rect 47938 153 47954 159
rect 47956 153 47972 159
rect 48124 153 48140 159
rect 48142 153 48158 159
rect 47949 143 47972 152
rect 48124 143 48147 152
rect 47922 133 47930 143
rect 47928 109 47930 133
rect 47938 123 47939 143
rect 47949 118 47952 143
rect 47971 123 47972 143
rect 47981 133 47988 143
rect 48108 133 48115 143
rect 48124 123 48125 143
rect 48144 118 48147 143
rect 48157 123 48158 143
rect 48167 133 48174 143
rect 47938 109 47972 113
rect 48124 109 48158 113
rect 48218 109 48220 159
rect 47824 103 47866 104
rect 48230 103 48272 104
rect 47824 96 47828 103
rect 47719 62 47724 96
rect 47748 62 47753 96
rect 47791 79 47862 96
rect 48234 79 48268 96
rect 48271 79 48305 96
rect 47791 62 47866 79
rect 47824 61 47866 62
rect 48230 62 48305 79
rect 48230 61 48272 62
rect 47802 55 47888 61
rect 48208 55 48294 61
rect 48336 55 48340 233
rect 48524 183 48528 251
rect 48533 207 48543 241
rect 48553 213 48573 241
rect 48553 207 48567 213
rect 48592 207 48603 251
rect 48634 246 48710 253
rect 48743 251 48752 279
rect 48655 228 48689 246
rect 48697 228 48699 246
rect 48634 221 48710 228
rect 48697 213 48699 221
rect 48741 213 48752 251
rect 48816 241 48820 395
rect 48823 378 48828 412
rect 48852 378 48857 412
rect 48858 400 48869 412
rect 49072 395 49114 421
rect 49478 395 49520 421
rect 49735 420 49747 424
rect 49757 420 49769 424
rect 49807 420 49819 424
rect 49829 421 49841 424
rect 49999 421 50011 424
rect 49829 420 49882 421
rect 49840 412 49882 420
rect 49723 400 49734 412
rect 49004 341 49008 395
rect 49064 387 49110 395
rect 49064 383 49080 387
rect 49072 380 49080 383
rect 49106 380 49110 387
rect 49114 383 49122 395
rect 49470 383 49478 395
rect 49482 387 49516 395
rect 49482 380 49486 387
rect 49512 380 49516 387
rect 49520 383 49528 395
rect 49060 379 49126 380
rect 49466 379 49532 380
rect 49072 371 49076 379
rect 49126 365 49176 367
rect 49416 365 49466 367
rect 49166 361 49220 365
rect 49372 361 49426 365
rect 49166 356 49186 361
rect 49406 356 49426 361
rect 49176 341 49178 356
rect 49004 261 49008 329
rect 49072 305 49076 341
rect 49170 331 49178 341
rect 49186 331 49187 351
rect 49176 315 49178 331
rect 49197 322 49200 356
rect 49219 331 49220 351
rect 49229 331 49236 341
rect 49356 331 49363 341
rect 49372 331 49373 351
rect 49392 322 49395 356
rect 49405 331 49406 351
rect 49415 331 49422 341
rect 49186 315 49202 321
rect 49204 315 49220 321
rect 49372 315 49388 321
rect 49390 315 49406 321
rect 49466 315 49468 365
rect 49009 267 49045 295
rect 49009 261 49023 267
rect 48688 212 48699 213
rect 48533 183 48540 207
rect 48688 183 48698 212
rect 48779 207 48791 241
rect 48801 207 48821 241
rect 48524 103 48528 171
rect 48592 133 48596 183
rect 48592 98 48596 103
rect 48343 62 48348 96
rect 48372 62 48377 96
rect 48592 94 48630 98
rect 48592 79 48600 94
rect 48626 79 48630 94
rect 48714 94 48748 98
rect 48714 79 48718 94
rect 48744 79 48748 94
rect 48592 61 48634 79
rect 48710 61 48752 79
rect 48570 55 48656 61
rect 48688 55 48774 61
rect 48816 55 48820 207
rect 48846 183 48853 211
rect 49004 183 49008 251
rect 49013 233 49023 261
rect 49033 261 49047 267
rect 49072 261 49083 305
rect 49509 267 49520 305
rect 49547 267 49583 295
rect 49584 267 49588 395
rect 49735 378 49740 412
rect 49764 378 49769 412
rect 49770 400 49781 412
rect 49795 400 49806 412
rect 49807 395 49882 412
rect 49958 420 50011 421
rect 50021 420 50033 424
rect 50071 420 50083 424
rect 50093 420 50105 424
rect 49958 412 50000 420
rect 49958 395 50033 412
rect 50034 400 50045 412
rect 50059 400 50070 412
rect 49772 341 49776 395
rect 49807 378 49878 395
rect 49882 383 49890 395
rect 49950 383 49958 395
rect 49962 378 49996 395
rect 49999 378 50033 395
rect 49840 371 49844 378
rect 49234 262 49284 264
rect 49308 262 49358 264
rect 49033 233 49053 261
rect 49072 233 49081 261
rect 49135 253 49169 261
rect 49114 246 49169 253
rect 49135 245 49169 246
rect 49237 253 49268 261
rect 49237 245 49271 253
rect 49072 213 49076 233
rect 49268 229 49271 245
rect 49135 228 49169 229
rect 49114 221 49169 228
rect 49237 221 49271 229
rect 49284 212 49286 262
rect 49324 253 49355 261
rect 49358 253 49360 262
rect 49547 261 49559 267
rect 49324 245 49360 253
rect 49423 253 49457 261
rect 49423 246 49478 253
rect 49423 245 49457 246
rect 49355 229 49360 245
rect 49549 233 49559 261
rect 49569 233 49589 267
rect 49772 261 49776 329
rect 49840 291 49844 341
rect 49840 251 49849 279
rect 49936 264 49946 291
rect 49895 262 49946 264
rect 49936 261 49947 262
rect 49903 253 49937 261
rect 49945 253 49947 261
rect 49324 221 49360 229
rect 49423 228 49457 229
rect 49423 221 49478 228
rect 49358 212 49360 221
rect 49004 103 49008 171
rect 49072 133 49076 183
rect 49126 159 49176 161
rect 49416 159 49466 161
rect 49176 143 49178 159
rect 49186 153 49202 159
rect 49204 153 49220 159
rect 49372 153 49388 159
rect 49390 153 49406 159
rect 49197 143 49220 152
rect 49372 143 49395 152
rect 49170 133 49178 143
rect 49176 109 49178 133
rect 49186 123 49187 143
rect 49197 118 49200 143
rect 49219 123 49220 143
rect 49229 133 49236 143
rect 49356 133 49363 143
rect 49372 123 49373 143
rect 49392 118 49395 143
rect 49405 123 49406 143
rect 49415 133 49422 143
rect 49186 109 49220 113
rect 49372 109 49406 113
rect 49466 109 49468 159
rect 49072 103 49114 104
rect 49478 103 49520 104
rect 49072 96 49076 103
rect 48967 62 48972 96
rect 48996 62 49001 96
rect 49039 79 49110 96
rect 49482 79 49516 96
rect 49519 79 49553 96
rect 49039 62 49114 79
rect 49072 61 49114 62
rect 49478 62 49553 79
rect 49478 61 49520 62
rect 49050 55 49136 61
rect 49456 55 49542 61
rect 49584 55 49588 233
rect 49772 183 49776 251
rect 49781 207 49791 241
rect 49801 213 49821 241
rect 49801 207 49815 213
rect 49840 207 49851 251
rect 49882 246 49958 253
rect 49991 251 50000 279
rect 49903 228 49937 246
rect 49945 228 49947 246
rect 49882 221 49958 228
rect 49945 213 49947 221
rect 49989 213 50000 251
rect 50064 241 50068 395
rect 50071 378 50076 412
rect 50100 378 50105 412
rect 50106 400 50117 412
rect 50320 395 50362 421
rect 50726 395 50768 421
rect 50983 420 50995 424
rect 51005 420 51017 424
rect 51055 420 51067 424
rect 51077 421 51089 424
rect 51247 421 51259 424
rect 51077 420 51130 421
rect 51088 412 51130 420
rect 50971 400 50982 412
rect 50252 341 50256 395
rect 50312 387 50358 395
rect 50312 383 50328 387
rect 50320 380 50328 383
rect 50354 380 50358 387
rect 50362 383 50370 395
rect 50718 383 50726 395
rect 50730 387 50764 395
rect 50730 380 50734 387
rect 50760 380 50764 387
rect 50768 383 50776 395
rect 50308 379 50374 380
rect 50714 379 50780 380
rect 50320 371 50324 379
rect 50374 365 50424 367
rect 50664 365 50714 367
rect 50414 361 50468 365
rect 50620 361 50674 365
rect 50414 356 50434 361
rect 50654 356 50674 361
rect 50424 341 50426 356
rect 50252 261 50256 329
rect 50320 305 50324 341
rect 50418 331 50426 341
rect 50434 331 50435 351
rect 50424 315 50426 331
rect 50445 322 50448 356
rect 50467 331 50468 351
rect 50477 331 50484 341
rect 50604 331 50611 341
rect 50620 331 50621 351
rect 50640 322 50643 356
rect 50653 331 50654 351
rect 50663 331 50670 341
rect 50434 315 50450 321
rect 50452 315 50468 321
rect 50620 315 50636 321
rect 50638 315 50654 321
rect 50714 315 50716 365
rect 50257 267 50293 295
rect 50257 261 50271 267
rect 49936 212 49947 213
rect 49781 183 49788 207
rect 49936 183 49946 212
rect 50027 207 50039 241
rect 50049 207 50069 241
rect 49772 103 49776 171
rect 49840 133 49844 183
rect 49840 98 49844 103
rect 49591 62 49596 96
rect 49620 62 49625 96
rect 49840 94 49878 98
rect 49840 79 49848 94
rect 49874 79 49878 94
rect 49962 94 49996 98
rect 49962 79 49966 94
rect 49992 79 49996 94
rect 49840 61 49882 79
rect 49958 61 50000 79
rect 49818 55 49904 61
rect 49936 55 50022 61
rect 50064 55 50068 207
rect 50094 183 50101 211
rect 50252 183 50256 251
rect 50261 233 50271 261
rect 50281 261 50295 267
rect 50320 261 50331 305
rect 50757 267 50768 305
rect 50795 267 50831 295
rect 50832 267 50836 395
rect 50983 378 50988 412
rect 51012 378 51017 412
rect 51018 400 51029 412
rect 51043 400 51054 412
rect 51055 395 51130 412
rect 51206 420 51259 421
rect 51269 420 51281 424
rect 51319 420 51331 424
rect 51341 420 51353 424
rect 51206 412 51248 420
rect 51206 395 51281 412
rect 51282 400 51293 412
rect 51307 400 51318 412
rect 51020 341 51024 395
rect 51055 378 51126 395
rect 51130 383 51138 395
rect 51198 383 51206 395
rect 51210 378 51244 395
rect 51247 378 51281 395
rect 51088 371 51092 378
rect 50482 262 50532 264
rect 50556 262 50606 264
rect 50281 233 50301 261
rect 50320 233 50329 261
rect 50383 253 50417 261
rect 50362 246 50417 253
rect 50383 245 50417 246
rect 50485 253 50516 261
rect 50485 245 50519 253
rect 50320 213 50324 233
rect 50516 229 50519 245
rect 50383 228 50417 229
rect 50362 221 50417 228
rect 50485 221 50519 229
rect 50532 212 50534 262
rect 50572 253 50603 261
rect 50606 253 50608 262
rect 50795 261 50807 267
rect 50572 245 50608 253
rect 50671 253 50705 261
rect 50671 246 50726 253
rect 50671 245 50705 246
rect 50603 229 50608 245
rect 50797 233 50807 261
rect 50817 233 50837 267
rect 51020 261 51024 329
rect 51088 291 51092 341
rect 51088 251 51097 279
rect 51184 264 51194 291
rect 51143 262 51194 264
rect 51184 261 51195 262
rect 51151 253 51185 261
rect 51193 253 51195 261
rect 50572 221 50608 229
rect 50671 228 50705 229
rect 50671 221 50726 228
rect 50606 212 50608 221
rect 50252 103 50256 171
rect 50320 133 50324 183
rect 50374 159 50424 161
rect 50664 159 50714 161
rect 50424 143 50426 159
rect 50434 153 50450 159
rect 50452 153 50468 159
rect 50620 153 50636 159
rect 50638 153 50654 159
rect 50445 143 50468 152
rect 50620 143 50643 152
rect 50418 133 50426 143
rect 50424 109 50426 133
rect 50434 123 50435 143
rect 50445 118 50448 143
rect 50467 123 50468 143
rect 50477 133 50484 143
rect 50604 133 50611 143
rect 50620 123 50621 143
rect 50640 118 50643 143
rect 50653 123 50654 143
rect 50663 133 50670 143
rect 50434 109 50468 113
rect 50620 109 50654 113
rect 50714 109 50716 159
rect 50320 103 50362 104
rect 50726 103 50768 104
rect 50320 96 50324 103
rect 50215 62 50220 96
rect 50244 62 50249 96
rect 50287 79 50358 96
rect 50730 79 50764 96
rect 50767 79 50801 96
rect 50287 62 50362 79
rect 50320 61 50362 62
rect 50726 62 50801 79
rect 50726 61 50768 62
rect 50298 55 50384 61
rect 50704 55 50790 61
rect 50832 55 50836 233
rect 51020 183 51024 251
rect 51029 207 51039 241
rect 51049 213 51069 241
rect 51049 207 51063 213
rect 51088 207 51099 251
rect 51130 246 51206 253
rect 51239 251 51248 279
rect 51151 228 51185 246
rect 51193 228 51195 246
rect 51130 221 51206 228
rect 51193 213 51195 221
rect 51237 213 51248 251
rect 51312 241 51316 395
rect 51319 378 51324 412
rect 51348 378 51353 412
rect 51354 400 51365 412
rect 51568 395 51610 421
rect 51974 395 52016 421
rect 52231 420 52243 424
rect 52253 420 52265 424
rect 52303 420 52315 424
rect 52325 421 52337 424
rect 52495 421 52507 424
rect 52325 420 52378 421
rect 52336 412 52378 420
rect 52219 400 52230 412
rect 51500 341 51504 395
rect 51560 387 51606 395
rect 51560 383 51576 387
rect 51568 380 51576 383
rect 51602 380 51606 387
rect 51610 383 51618 395
rect 51966 383 51974 395
rect 51978 387 52012 395
rect 51978 380 51982 387
rect 52008 380 52012 387
rect 52016 383 52024 395
rect 51556 379 51622 380
rect 51962 379 52028 380
rect 51568 371 51572 379
rect 51622 365 51672 367
rect 51912 365 51962 367
rect 51662 361 51716 365
rect 51868 361 51922 365
rect 51662 356 51682 361
rect 51902 356 51922 361
rect 51672 341 51674 356
rect 51500 261 51504 329
rect 51568 305 51572 341
rect 51666 331 51674 341
rect 51682 331 51683 351
rect 51672 315 51674 331
rect 51693 322 51696 356
rect 51715 331 51716 351
rect 51725 331 51732 341
rect 51852 331 51859 341
rect 51868 331 51869 351
rect 51888 322 51891 356
rect 51901 331 51902 351
rect 51911 331 51918 341
rect 51682 315 51698 321
rect 51700 315 51716 321
rect 51868 315 51884 321
rect 51886 315 51902 321
rect 51962 315 51964 365
rect 51505 267 51541 295
rect 51505 261 51519 267
rect 51184 212 51195 213
rect 51029 183 51036 207
rect 51184 183 51194 212
rect 51275 207 51287 241
rect 51297 207 51317 241
rect 51020 103 51024 171
rect 51088 133 51092 183
rect 51088 98 51092 103
rect 50839 62 50844 96
rect 50868 62 50873 96
rect 51088 94 51126 98
rect 51088 79 51096 94
rect 51122 79 51126 94
rect 51210 94 51244 98
rect 51210 79 51214 94
rect 51240 79 51244 94
rect 51088 61 51130 79
rect 51206 61 51248 79
rect 51066 55 51152 61
rect 51184 55 51270 61
rect 51312 55 51316 207
rect 51342 183 51349 211
rect 51500 183 51504 251
rect 51509 233 51519 261
rect 51529 261 51543 267
rect 51568 261 51579 305
rect 52005 267 52016 305
rect 52043 267 52079 295
rect 52080 267 52084 395
rect 52231 378 52236 412
rect 52260 378 52265 412
rect 52266 400 52277 412
rect 52291 400 52302 412
rect 52303 395 52378 412
rect 52454 420 52507 421
rect 52517 420 52529 424
rect 52567 420 52579 424
rect 52589 420 52601 424
rect 52454 412 52496 420
rect 52454 395 52529 412
rect 52530 400 52541 412
rect 52555 400 52566 412
rect 52268 341 52272 395
rect 52303 378 52374 395
rect 52378 383 52386 395
rect 52446 383 52454 395
rect 52458 378 52492 395
rect 52495 378 52529 395
rect 52336 371 52340 378
rect 51730 262 51780 264
rect 51804 262 51854 264
rect 51529 233 51549 261
rect 51568 233 51577 261
rect 51631 253 51665 261
rect 51610 246 51665 253
rect 51631 245 51665 246
rect 51733 253 51764 261
rect 51733 245 51767 253
rect 51568 213 51572 233
rect 51764 229 51767 245
rect 51631 228 51665 229
rect 51610 221 51665 228
rect 51733 221 51767 229
rect 51780 212 51782 262
rect 51820 253 51851 261
rect 51854 253 51856 262
rect 52043 261 52055 267
rect 51820 245 51856 253
rect 51919 253 51953 261
rect 51919 246 51974 253
rect 51919 245 51953 246
rect 51851 229 51856 245
rect 52045 233 52055 261
rect 52065 233 52085 267
rect 52268 261 52272 329
rect 52336 291 52340 341
rect 52336 251 52345 279
rect 52432 264 52442 291
rect 52391 262 52442 264
rect 52432 261 52443 262
rect 52399 253 52433 261
rect 52441 253 52443 261
rect 51820 221 51856 229
rect 51919 228 51953 229
rect 51919 221 51974 228
rect 51854 212 51856 221
rect 51500 103 51504 171
rect 51568 133 51572 183
rect 51622 159 51672 161
rect 51912 159 51962 161
rect 51672 143 51674 159
rect 51682 153 51698 159
rect 51700 153 51716 159
rect 51868 153 51884 159
rect 51886 153 51902 159
rect 51693 143 51716 152
rect 51868 143 51891 152
rect 51666 133 51674 143
rect 51672 109 51674 133
rect 51682 123 51683 143
rect 51693 118 51696 143
rect 51715 123 51716 143
rect 51725 133 51732 143
rect 51852 133 51859 143
rect 51868 123 51869 143
rect 51888 118 51891 143
rect 51901 123 51902 143
rect 51911 133 51918 143
rect 51682 109 51716 113
rect 51868 109 51902 113
rect 51962 109 51964 159
rect 51568 103 51610 104
rect 51974 103 52016 104
rect 51568 96 51572 103
rect 51463 62 51468 96
rect 51492 62 51497 96
rect 51535 79 51606 96
rect 51978 79 52012 96
rect 52015 79 52049 96
rect 51535 62 51610 79
rect 51568 61 51610 62
rect 51974 62 52049 79
rect 51974 61 52016 62
rect 51546 55 51632 61
rect 51952 55 52038 61
rect 52080 55 52084 233
rect 52268 183 52272 251
rect 52277 207 52287 241
rect 52297 213 52317 241
rect 52297 207 52311 213
rect 52336 207 52347 251
rect 52378 246 52454 253
rect 52487 251 52496 279
rect 52399 228 52433 246
rect 52441 228 52443 246
rect 52378 221 52454 228
rect 52441 213 52443 221
rect 52485 213 52496 251
rect 52560 241 52564 395
rect 52567 378 52572 412
rect 52596 378 52601 412
rect 52602 400 52613 412
rect 52816 395 52858 421
rect 53222 395 53264 421
rect 53479 420 53491 424
rect 53501 420 53513 424
rect 53551 420 53563 424
rect 53573 421 53585 424
rect 53743 421 53755 424
rect 53573 420 53626 421
rect 53584 412 53626 420
rect 53467 400 53478 412
rect 52748 341 52752 395
rect 52808 387 52854 395
rect 52808 383 52824 387
rect 52816 380 52824 383
rect 52850 380 52854 387
rect 52858 383 52866 395
rect 53214 383 53222 395
rect 53226 387 53260 395
rect 53226 380 53230 387
rect 53256 380 53260 387
rect 53264 383 53272 395
rect 52804 379 52870 380
rect 53210 379 53276 380
rect 52816 371 52820 379
rect 52870 365 52920 367
rect 53160 365 53210 367
rect 52910 361 52964 365
rect 53116 361 53170 365
rect 52910 356 52930 361
rect 53150 356 53170 361
rect 52920 341 52922 356
rect 52748 261 52752 329
rect 52816 305 52820 341
rect 52914 331 52922 341
rect 52930 331 52931 351
rect 52920 315 52922 331
rect 52941 322 52944 356
rect 52963 331 52964 351
rect 52973 331 52980 341
rect 53100 331 53107 341
rect 53116 331 53117 351
rect 53136 322 53139 356
rect 53149 331 53150 351
rect 53159 331 53166 341
rect 52930 315 52946 321
rect 52948 315 52964 321
rect 53116 315 53132 321
rect 53134 315 53150 321
rect 53210 315 53212 365
rect 52753 267 52789 295
rect 52753 261 52767 267
rect 52432 212 52443 213
rect 52277 183 52284 207
rect 52432 183 52442 212
rect 52523 207 52535 241
rect 52545 207 52565 241
rect 52268 103 52272 171
rect 52336 133 52340 183
rect 52336 98 52340 103
rect 52087 62 52092 96
rect 52116 62 52121 96
rect 52336 94 52374 98
rect 52336 79 52344 94
rect 52370 79 52374 94
rect 52458 94 52492 98
rect 52458 79 52462 94
rect 52488 79 52492 94
rect 52336 61 52378 79
rect 52454 61 52496 79
rect 52314 55 52400 61
rect 52432 55 52518 61
rect 52560 55 52564 207
rect 52590 183 52597 211
rect 52748 183 52752 251
rect 52757 233 52767 261
rect 52777 261 52791 267
rect 52816 261 52827 305
rect 53253 267 53264 305
rect 53291 267 53327 295
rect 53328 267 53332 395
rect 53479 378 53484 412
rect 53508 378 53513 412
rect 53514 400 53525 412
rect 53539 400 53550 412
rect 53551 395 53626 412
rect 53702 420 53755 421
rect 53765 420 53777 424
rect 53815 420 53827 424
rect 53837 420 53849 424
rect 53702 412 53744 420
rect 53702 395 53777 412
rect 53778 400 53789 412
rect 53803 400 53814 412
rect 53516 341 53520 395
rect 53551 378 53622 395
rect 53626 383 53634 395
rect 53694 383 53702 395
rect 53706 378 53740 395
rect 53743 378 53777 395
rect 53584 371 53588 378
rect 52978 262 53028 264
rect 53052 262 53102 264
rect 52777 233 52797 261
rect 52816 233 52825 261
rect 52879 253 52913 261
rect 52858 246 52913 253
rect 52879 245 52913 246
rect 52981 253 53012 261
rect 52981 245 53015 253
rect 52816 213 52820 233
rect 53012 229 53015 245
rect 52879 228 52913 229
rect 52858 221 52913 228
rect 52981 221 53015 229
rect 53028 212 53030 262
rect 53068 253 53099 261
rect 53102 253 53104 262
rect 53291 261 53303 267
rect 53068 245 53104 253
rect 53167 253 53201 261
rect 53167 246 53222 253
rect 53167 245 53201 246
rect 53099 229 53104 245
rect 53293 233 53303 261
rect 53313 233 53333 267
rect 53516 261 53520 329
rect 53584 291 53588 341
rect 53584 251 53593 279
rect 53680 264 53690 291
rect 53639 262 53690 264
rect 53680 261 53691 262
rect 53647 253 53681 261
rect 53689 253 53691 261
rect 53068 221 53104 229
rect 53167 228 53201 229
rect 53167 221 53222 228
rect 53102 212 53104 221
rect 52748 103 52752 171
rect 52816 133 52820 183
rect 52870 159 52920 161
rect 53160 159 53210 161
rect 52920 143 52922 159
rect 52930 153 52946 159
rect 52948 153 52964 159
rect 53116 153 53132 159
rect 53134 153 53150 159
rect 52941 143 52964 152
rect 53116 143 53139 152
rect 52914 133 52922 143
rect 52920 109 52922 133
rect 52930 123 52931 143
rect 52941 118 52944 143
rect 52963 123 52964 143
rect 52973 133 52980 143
rect 53100 133 53107 143
rect 53116 123 53117 143
rect 53136 118 53139 143
rect 53149 123 53150 143
rect 53159 133 53166 143
rect 52930 109 52964 113
rect 53116 109 53150 113
rect 53210 109 53212 159
rect 52816 103 52858 104
rect 53222 103 53264 104
rect 52816 96 52820 103
rect 52711 62 52716 96
rect 52740 62 52745 96
rect 52783 79 52854 96
rect 53226 79 53260 96
rect 53263 79 53297 96
rect 52783 62 52858 79
rect 52816 61 52858 62
rect 53222 62 53297 79
rect 53222 61 53264 62
rect 52794 55 52880 61
rect 53200 55 53286 61
rect 53328 55 53332 233
rect 53516 183 53520 251
rect 53525 207 53535 241
rect 53545 213 53565 241
rect 53545 207 53559 213
rect 53584 207 53595 251
rect 53626 246 53702 253
rect 53735 251 53744 279
rect 53647 228 53681 246
rect 53689 228 53691 246
rect 53626 221 53702 228
rect 53689 213 53691 221
rect 53733 213 53744 251
rect 53808 241 53812 395
rect 53815 378 53820 412
rect 53844 378 53849 412
rect 53850 400 53861 412
rect 54064 395 54106 421
rect 54470 395 54512 421
rect 54727 420 54739 424
rect 54749 420 54761 424
rect 54799 420 54811 424
rect 54821 421 54833 424
rect 54991 421 55003 424
rect 54821 420 54874 421
rect 54832 412 54874 420
rect 54715 400 54726 412
rect 53996 341 54000 395
rect 54056 387 54102 395
rect 54056 383 54072 387
rect 54064 380 54072 383
rect 54098 380 54102 387
rect 54106 383 54114 395
rect 54462 383 54470 395
rect 54474 387 54508 395
rect 54474 380 54478 387
rect 54504 380 54508 387
rect 54512 383 54520 395
rect 54052 379 54118 380
rect 54458 379 54524 380
rect 54064 371 54068 379
rect 54118 365 54168 367
rect 54408 365 54458 367
rect 54158 361 54212 365
rect 54364 361 54418 365
rect 54158 356 54178 361
rect 54398 356 54418 361
rect 54168 341 54170 356
rect 53996 261 54000 329
rect 54064 305 54068 341
rect 54162 331 54170 341
rect 54178 331 54179 351
rect 54168 315 54170 331
rect 54189 322 54192 356
rect 54211 331 54212 351
rect 54221 331 54228 341
rect 54348 331 54355 341
rect 54364 331 54365 351
rect 54384 322 54387 356
rect 54397 331 54398 351
rect 54407 331 54414 341
rect 54178 315 54194 321
rect 54196 315 54212 321
rect 54364 315 54380 321
rect 54382 315 54398 321
rect 54458 315 54460 365
rect 54001 267 54037 295
rect 54001 261 54015 267
rect 53680 212 53691 213
rect 53525 183 53532 207
rect 53680 183 53690 212
rect 53771 207 53783 241
rect 53793 207 53813 241
rect 53516 103 53520 171
rect 53584 133 53588 183
rect 53584 98 53588 103
rect 53335 62 53340 96
rect 53364 62 53369 96
rect 53584 94 53622 98
rect 53584 79 53592 94
rect 53618 79 53622 94
rect 53706 94 53740 98
rect 53706 79 53710 94
rect 53736 79 53740 94
rect 53584 61 53626 79
rect 53702 61 53744 79
rect 53562 55 53648 61
rect 53680 55 53766 61
rect 53808 55 53812 207
rect 53838 183 53845 211
rect 53996 183 54000 251
rect 54005 233 54015 261
rect 54025 261 54039 267
rect 54064 261 54075 305
rect 54501 267 54512 305
rect 54539 267 54575 295
rect 54576 267 54580 395
rect 54727 378 54732 412
rect 54756 378 54761 412
rect 54762 400 54773 412
rect 54787 400 54798 412
rect 54799 395 54874 412
rect 54950 420 55003 421
rect 55013 420 55025 424
rect 55063 420 55075 424
rect 55085 420 55097 424
rect 54950 412 54992 420
rect 54950 395 55025 412
rect 55026 400 55037 412
rect 55051 400 55062 412
rect 54764 341 54768 395
rect 54799 378 54870 395
rect 54874 383 54882 395
rect 54942 383 54950 395
rect 54954 378 54988 395
rect 54991 378 55025 395
rect 54832 371 54836 378
rect 54226 262 54276 264
rect 54300 262 54350 264
rect 54025 233 54045 261
rect 54064 233 54073 261
rect 54127 253 54161 261
rect 54106 246 54161 253
rect 54127 245 54161 246
rect 54229 253 54260 261
rect 54229 245 54263 253
rect 54064 213 54068 233
rect 54260 229 54263 245
rect 54127 228 54161 229
rect 54106 221 54161 228
rect 54229 221 54263 229
rect 54276 212 54278 262
rect 54316 253 54347 261
rect 54350 253 54352 262
rect 54539 261 54551 267
rect 54316 245 54352 253
rect 54415 253 54449 261
rect 54415 246 54470 253
rect 54415 245 54449 246
rect 54347 229 54352 245
rect 54541 233 54551 261
rect 54561 233 54581 267
rect 54764 261 54768 329
rect 54832 291 54836 341
rect 54832 251 54841 279
rect 54928 264 54938 291
rect 54887 262 54938 264
rect 54928 261 54939 262
rect 54895 253 54929 261
rect 54937 253 54939 261
rect 54316 221 54352 229
rect 54415 228 54449 229
rect 54415 221 54470 228
rect 54350 212 54352 221
rect 53996 103 54000 171
rect 54064 133 54068 183
rect 54118 159 54168 161
rect 54408 159 54458 161
rect 54168 143 54170 159
rect 54178 153 54194 159
rect 54196 153 54212 159
rect 54364 153 54380 159
rect 54382 153 54398 159
rect 54189 143 54212 152
rect 54364 143 54387 152
rect 54162 133 54170 143
rect 54168 109 54170 133
rect 54178 123 54179 143
rect 54189 118 54192 143
rect 54211 123 54212 143
rect 54221 133 54228 143
rect 54348 133 54355 143
rect 54364 123 54365 143
rect 54384 118 54387 143
rect 54397 123 54398 143
rect 54407 133 54414 143
rect 54178 109 54212 113
rect 54364 109 54398 113
rect 54458 109 54460 159
rect 54064 103 54106 104
rect 54470 103 54512 104
rect 54064 96 54068 103
rect 53959 62 53964 96
rect 53988 62 53993 96
rect 54031 79 54102 96
rect 54474 79 54508 96
rect 54511 79 54545 96
rect 54031 62 54106 79
rect 54064 61 54106 62
rect 54470 62 54545 79
rect 54470 61 54512 62
rect 54042 55 54128 61
rect 54448 55 54534 61
rect 54576 55 54580 233
rect 54764 183 54768 251
rect 54773 207 54783 241
rect 54793 213 54813 241
rect 54793 207 54807 213
rect 54832 207 54843 251
rect 54874 246 54950 253
rect 54983 251 54992 279
rect 54895 228 54929 246
rect 54937 228 54939 246
rect 54874 221 54950 228
rect 54937 213 54939 221
rect 54981 213 54992 251
rect 55056 241 55060 395
rect 55063 378 55068 412
rect 55092 378 55097 412
rect 55098 400 55109 412
rect 55312 395 55354 421
rect 55718 395 55760 421
rect 55975 420 55987 424
rect 55997 420 56009 424
rect 56047 420 56059 424
rect 56069 421 56081 424
rect 56239 421 56251 424
rect 56069 420 56122 421
rect 56080 412 56122 420
rect 55963 400 55974 412
rect 55244 341 55248 395
rect 55304 387 55350 395
rect 55304 383 55320 387
rect 55312 380 55320 383
rect 55346 380 55350 387
rect 55354 383 55362 395
rect 55710 383 55718 395
rect 55722 387 55756 395
rect 55722 380 55726 387
rect 55752 380 55756 387
rect 55760 383 55768 395
rect 55300 379 55366 380
rect 55706 379 55772 380
rect 55312 371 55316 379
rect 55366 365 55416 367
rect 55656 365 55706 367
rect 55406 361 55460 365
rect 55612 361 55666 365
rect 55406 356 55426 361
rect 55646 356 55666 361
rect 55416 341 55418 356
rect 55244 261 55248 329
rect 55312 305 55316 341
rect 55410 331 55418 341
rect 55426 331 55427 351
rect 55416 315 55418 331
rect 55437 322 55440 356
rect 55459 331 55460 351
rect 55469 331 55476 341
rect 55596 331 55603 341
rect 55612 331 55613 351
rect 55632 322 55635 356
rect 55645 331 55646 351
rect 55655 331 55662 341
rect 55426 315 55442 321
rect 55444 315 55460 321
rect 55612 315 55628 321
rect 55630 315 55646 321
rect 55706 315 55708 365
rect 55249 267 55285 295
rect 55249 261 55263 267
rect 54928 212 54939 213
rect 54773 183 54780 207
rect 54928 183 54938 212
rect 55019 207 55031 241
rect 55041 207 55061 241
rect 54764 103 54768 171
rect 54832 133 54836 183
rect 54832 98 54836 103
rect 54583 62 54588 96
rect 54612 62 54617 96
rect 54832 94 54870 98
rect 54832 79 54840 94
rect 54866 79 54870 94
rect 54954 94 54988 98
rect 54954 79 54958 94
rect 54984 79 54988 94
rect 54832 61 54874 79
rect 54950 61 54992 79
rect 54810 55 54896 61
rect 54928 55 55014 61
rect 55056 55 55060 207
rect 55086 183 55093 211
rect 55244 183 55248 251
rect 55253 233 55263 261
rect 55273 261 55287 267
rect 55312 261 55323 305
rect 55749 267 55760 305
rect 55787 267 55823 295
rect 55824 267 55828 395
rect 55975 378 55980 412
rect 56004 378 56009 412
rect 56010 400 56021 412
rect 56035 400 56046 412
rect 56047 395 56122 412
rect 56198 420 56251 421
rect 56261 420 56273 424
rect 56311 420 56323 424
rect 56333 420 56345 424
rect 56198 412 56240 420
rect 56198 395 56273 412
rect 56274 400 56285 412
rect 56299 400 56310 412
rect 56012 341 56016 395
rect 56047 378 56118 395
rect 56122 383 56130 395
rect 56190 383 56198 395
rect 56202 378 56236 395
rect 56239 378 56273 395
rect 56080 371 56084 378
rect 55474 262 55524 264
rect 55548 262 55598 264
rect 55273 233 55293 261
rect 55312 233 55321 261
rect 55375 253 55409 261
rect 55354 246 55409 253
rect 55375 245 55409 246
rect 55477 253 55508 261
rect 55477 245 55511 253
rect 55312 213 55316 233
rect 55508 229 55511 245
rect 55375 228 55409 229
rect 55354 221 55409 228
rect 55477 221 55511 229
rect 55524 212 55526 262
rect 55564 253 55595 261
rect 55598 253 55600 262
rect 55787 261 55799 267
rect 55564 245 55600 253
rect 55663 253 55697 261
rect 55663 246 55718 253
rect 55663 245 55697 246
rect 55595 229 55600 245
rect 55789 233 55799 261
rect 55809 233 55829 267
rect 56012 261 56016 329
rect 56080 291 56084 341
rect 56080 251 56089 279
rect 56176 264 56186 291
rect 56135 262 56186 264
rect 56176 261 56187 262
rect 56143 253 56177 261
rect 56185 253 56187 261
rect 55564 221 55600 229
rect 55663 228 55697 229
rect 55663 221 55718 228
rect 55598 212 55600 221
rect 55244 103 55248 171
rect 55312 133 55316 183
rect 55366 159 55416 161
rect 55656 159 55706 161
rect 55416 143 55418 159
rect 55426 153 55442 159
rect 55444 153 55460 159
rect 55612 153 55628 159
rect 55630 153 55646 159
rect 55437 143 55460 152
rect 55612 143 55635 152
rect 55410 133 55418 143
rect 55416 109 55418 133
rect 55426 123 55427 143
rect 55437 118 55440 143
rect 55459 123 55460 143
rect 55469 133 55476 143
rect 55596 133 55603 143
rect 55612 123 55613 143
rect 55632 118 55635 143
rect 55645 123 55646 143
rect 55655 133 55662 143
rect 55426 109 55460 113
rect 55612 109 55646 113
rect 55706 109 55708 159
rect 55312 103 55354 104
rect 55718 103 55760 104
rect 55312 96 55316 103
rect 55207 62 55212 96
rect 55236 62 55241 96
rect 55279 79 55350 96
rect 55722 79 55756 96
rect 55759 79 55793 96
rect 55279 62 55354 79
rect 55312 61 55354 62
rect 55718 62 55793 79
rect 55718 61 55760 62
rect 55290 55 55376 61
rect 55696 55 55782 61
rect 55824 55 55828 233
rect 56012 183 56016 251
rect 56021 207 56031 241
rect 56041 213 56061 241
rect 56041 207 56055 213
rect 56080 207 56091 251
rect 56122 246 56198 253
rect 56231 251 56240 279
rect 56143 228 56177 246
rect 56185 228 56187 246
rect 56122 221 56198 228
rect 56185 213 56187 221
rect 56229 213 56240 251
rect 56304 241 56308 395
rect 56311 378 56316 412
rect 56340 378 56345 412
rect 56346 400 56357 412
rect 56560 395 56602 421
rect 56966 395 57008 421
rect 57223 420 57235 424
rect 57245 420 57257 424
rect 57295 420 57307 424
rect 57317 421 57329 424
rect 57487 421 57499 424
rect 57317 420 57370 421
rect 57328 412 57370 420
rect 57211 400 57222 412
rect 56492 341 56496 395
rect 56552 387 56598 395
rect 56552 383 56568 387
rect 56560 380 56568 383
rect 56594 380 56598 387
rect 56602 383 56610 395
rect 56958 383 56966 395
rect 56970 387 57004 395
rect 56970 380 56974 387
rect 57000 380 57004 387
rect 57008 383 57016 395
rect 56548 379 56614 380
rect 56954 379 57020 380
rect 56560 371 56564 379
rect 56614 365 56664 367
rect 56904 365 56954 367
rect 56654 361 56708 365
rect 56860 361 56914 365
rect 56654 356 56674 361
rect 56894 356 56914 361
rect 56664 341 56666 356
rect 56492 261 56496 329
rect 56560 305 56564 341
rect 56658 331 56666 341
rect 56674 331 56675 351
rect 56664 315 56666 331
rect 56685 322 56688 356
rect 56707 331 56708 351
rect 56717 331 56724 341
rect 56844 331 56851 341
rect 56860 331 56861 351
rect 56880 322 56883 356
rect 56893 331 56894 351
rect 56903 331 56910 341
rect 56674 315 56690 321
rect 56692 315 56708 321
rect 56860 315 56876 321
rect 56878 315 56894 321
rect 56954 315 56956 365
rect 56497 267 56533 295
rect 56497 261 56511 267
rect 56176 212 56187 213
rect 56021 183 56028 207
rect 56176 183 56186 212
rect 56267 207 56279 241
rect 56289 207 56309 241
rect 56012 103 56016 171
rect 56080 133 56084 183
rect 56080 98 56084 103
rect 55831 62 55836 96
rect 55860 62 55865 96
rect 56080 94 56118 98
rect 56080 79 56088 94
rect 56114 79 56118 94
rect 56202 94 56236 98
rect 56202 79 56206 94
rect 56232 79 56236 94
rect 56080 61 56122 79
rect 56198 61 56240 79
rect 56058 55 56144 61
rect 56176 55 56262 61
rect 56304 55 56308 207
rect 56334 183 56341 211
rect 56492 183 56496 251
rect 56501 233 56511 261
rect 56521 261 56535 267
rect 56560 261 56571 305
rect 56997 267 57008 305
rect 57035 267 57071 295
rect 57072 267 57076 395
rect 57223 378 57228 412
rect 57252 378 57257 412
rect 57258 400 57269 412
rect 57283 400 57294 412
rect 57295 395 57370 412
rect 57446 420 57499 421
rect 57509 420 57521 424
rect 57559 420 57571 424
rect 57581 420 57593 424
rect 57446 412 57488 420
rect 57446 395 57521 412
rect 57522 400 57533 412
rect 57547 400 57558 412
rect 57260 341 57264 395
rect 57295 378 57366 395
rect 57370 383 57378 395
rect 57438 383 57446 395
rect 57450 378 57484 395
rect 57487 378 57521 395
rect 57328 371 57332 378
rect 56722 262 56772 264
rect 56796 262 56846 264
rect 56521 233 56541 261
rect 56560 233 56569 261
rect 56623 253 56657 261
rect 56602 246 56657 253
rect 56623 245 56657 246
rect 56725 253 56756 261
rect 56725 245 56759 253
rect 56560 213 56564 233
rect 56756 229 56759 245
rect 56623 228 56657 229
rect 56602 221 56657 228
rect 56725 221 56759 229
rect 56772 212 56774 262
rect 56812 253 56843 261
rect 56846 253 56848 262
rect 57035 261 57047 267
rect 56812 245 56848 253
rect 56911 253 56945 261
rect 56911 246 56966 253
rect 56911 245 56945 246
rect 56843 229 56848 245
rect 57037 233 57047 261
rect 57057 233 57077 267
rect 57260 261 57264 329
rect 57328 291 57332 341
rect 57328 251 57337 279
rect 57424 264 57434 291
rect 57383 262 57434 264
rect 57424 261 57435 262
rect 57391 253 57425 261
rect 57433 253 57435 261
rect 56812 221 56848 229
rect 56911 228 56945 229
rect 56911 221 56966 228
rect 56846 212 56848 221
rect 56492 103 56496 171
rect 56560 133 56564 183
rect 56614 159 56664 161
rect 56904 159 56954 161
rect 56664 143 56666 159
rect 56674 153 56690 159
rect 56692 153 56708 159
rect 56860 153 56876 159
rect 56878 153 56894 159
rect 56685 143 56708 152
rect 56860 143 56883 152
rect 56658 133 56666 143
rect 56664 109 56666 133
rect 56674 123 56675 143
rect 56685 118 56688 143
rect 56707 123 56708 143
rect 56717 133 56724 143
rect 56844 133 56851 143
rect 56860 123 56861 143
rect 56880 118 56883 143
rect 56893 123 56894 143
rect 56903 133 56910 143
rect 56674 109 56708 113
rect 56860 109 56894 113
rect 56954 109 56956 159
rect 56560 103 56602 104
rect 56966 103 57008 104
rect 56560 96 56564 103
rect 56455 62 56460 96
rect 56484 62 56489 96
rect 56527 79 56598 96
rect 56970 79 57004 96
rect 57007 79 57041 96
rect 56527 62 56602 79
rect 56560 61 56602 62
rect 56966 62 57041 79
rect 56966 61 57008 62
rect 56538 55 56624 61
rect 56944 55 57030 61
rect 57072 55 57076 233
rect 57260 183 57264 251
rect 57269 207 57279 241
rect 57289 213 57309 241
rect 57289 207 57303 213
rect 57328 207 57339 251
rect 57370 246 57446 253
rect 57479 251 57488 279
rect 57391 228 57425 246
rect 57433 228 57435 246
rect 57370 221 57446 228
rect 57433 213 57435 221
rect 57477 213 57488 251
rect 57552 241 57556 395
rect 57559 378 57564 412
rect 57588 378 57593 412
rect 57594 400 57605 412
rect 57808 395 57850 421
rect 58214 395 58256 421
rect 58471 420 58483 424
rect 58493 420 58505 424
rect 58543 420 58555 424
rect 58565 421 58577 424
rect 58735 421 58747 424
rect 58565 420 58618 421
rect 58576 412 58618 420
rect 58459 400 58470 412
rect 57740 341 57744 395
rect 57800 387 57846 395
rect 57800 383 57816 387
rect 57808 380 57816 383
rect 57842 380 57846 387
rect 57850 383 57858 395
rect 58206 383 58214 395
rect 58218 387 58252 395
rect 58218 380 58222 387
rect 58248 380 58252 387
rect 58256 383 58264 395
rect 57796 379 57862 380
rect 58202 379 58268 380
rect 57808 371 57812 379
rect 57862 365 57912 367
rect 58152 365 58202 367
rect 57902 361 57956 365
rect 58108 361 58162 365
rect 57902 356 57922 361
rect 58142 356 58162 361
rect 57912 341 57914 356
rect 57740 261 57744 329
rect 57808 305 57812 341
rect 57906 331 57914 341
rect 57922 331 57923 351
rect 57912 315 57914 331
rect 57933 322 57936 356
rect 57955 331 57956 351
rect 57965 331 57972 341
rect 58092 331 58099 341
rect 58108 331 58109 351
rect 58128 322 58131 356
rect 58141 331 58142 351
rect 58151 331 58158 341
rect 57922 315 57938 321
rect 57940 315 57956 321
rect 58108 315 58124 321
rect 58126 315 58142 321
rect 58202 315 58204 365
rect 57745 267 57781 295
rect 57745 261 57759 267
rect 57424 212 57435 213
rect 57269 183 57276 207
rect 57424 183 57434 212
rect 57515 207 57527 241
rect 57537 207 57557 241
rect 57260 103 57264 171
rect 57328 133 57332 183
rect 57328 98 57332 103
rect 57079 62 57084 96
rect 57108 62 57113 96
rect 57328 94 57366 98
rect 57328 79 57336 94
rect 57362 79 57366 94
rect 57450 94 57484 98
rect 57450 79 57454 94
rect 57480 79 57484 94
rect 57328 61 57370 79
rect 57446 61 57488 79
rect 57306 55 57392 61
rect 57424 55 57510 61
rect 57552 55 57556 207
rect 57582 183 57589 211
rect 57740 183 57744 251
rect 57749 233 57759 261
rect 57769 261 57783 267
rect 57808 261 57819 305
rect 58245 267 58256 305
rect 58283 267 58319 295
rect 58320 267 58324 395
rect 58471 378 58476 412
rect 58500 378 58505 412
rect 58506 400 58517 412
rect 58531 400 58542 412
rect 58543 395 58618 412
rect 58694 420 58747 421
rect 58757 420 58769 424
rect 58807 420 58819 424
rect 58829 420 58841 424
rect 58694 412 58736 420
rect 58694 395 58769 412
rect 58770 400 58781 412
rect 58795 400 58806 412
rect 58508 341 58512 395
rect 58543 378 58614 395
rect 58618 383 58626 395
rect 58686 383 58694 395
rect 58698 378 58732 395
rect 58735 378 58769 395
rect 58576 371 58580 378
rect 57970 262 58020 264
rect 58044 262 58094 264
rect 57769 233 57789 261
rect 57808 233 57817 261
rect 57871 253 57905 261
rect 57850 246 57905 253
rect 57871 245 57905 246
rect 57973 253 58004 261
rect 57973 245 58007 253
rect 57808 213 57812 233
rect 58004 229 58007 245
rect 57871 228 57905 229
rect 57850 221 57905 228
rect 57973 221 58007 229
rect 58020 212 58022 262
rect 58060 253 58091 261
rect 58094 253 58096 262
rect 58283 261 58295 267
rect 58060 245 58096 253
rect 58159 253 58193 261
rect 58159 246 58214 253
rect 58159 245 58193 246
rect 58091 229 58096 245
rect 58285 233 58295 261
rect 58305 233 58325 267
rect 58508 261 58512 329
rect 58576 291 58580 341
rect 58576 251 58585 279
rect 58672 264 58682 291
rect 58631 262 58682 264
rect 58672 261 58683 262
rect 58639 253 58673 261
rect 58681 253 58683 261
rect 58060 221 58096 229
rect 58159 228 58193 229
rect 58159 221 58214 228
rect 58094 212 58096 221
rect 57740 103 57744 171
rect 57808 133 57812 183
rect 57862 159 57912 161
rect 58152 159 58202 161
rect 57912 143 57914 159
rect 57922 153 57938 159
rect 57940 153 57956 159
rect 58108 153 58124 159
rect 58126 153 58142 159
rect 57933 143 57956 152
rect 58108 143 58131 152
rect 57906 133 57914 143
rect 57912 109 57914 133
rect 57922 123 57923 143
rect 57933 118 57936 143
rect 57955 123 57956 143
rect 57965 133 57972 143
rect 58092 133 58099 143
rect 58108 123 58109 143
rect 58128 118 58131 143
rect 58141 123 58142 143
rect 58151 133 58158 143
rect 57922 109 57956 113
rect 58108 109 58142 113
rect 58202 109 58204 159
rect 57808 103 57850 104
rect 58214 103 58256 104
rect 57808 96 57812 103
rect 57703 62 57708 96
rect 57732 62 57737 96
rect 57775 79 57846 96
rect 58218 79 58252 96
rect 58255 79 58289 96
rect 57775 62 57850 79
rect 57808 61 57850 62
rect 58214 62 58289 79
rect 58214 61 58256 62
rect 57786 55 57872 61
rect 58192 55 58278 61
rect 58320 55 58324 233
rect 58508 183 58512 251
rect 58517 207 58527 241
rect 58537 213 58557 241
rect 58537 207 58551 213
rect 58576 207 58587 251
rect 58618 246 58694 253
rect 58727 251 58736 279
rect 58639 228 58673 246
rect 58681 228 58683 246
rect 58618 221 58694 228
rect 58681 213 58683 221
rect 58725 213 58736 251
rect 58800 241 58804 395
rect 58807 378 58812 412
rect 58836 378 58841 412
rect 58842 400 58853 412
rect 59056 395 59098 421
rect 59462 395 59504 421
rect 59719 420 59731 424
rect 59741 420 59753 424
rect 59791 420 59803 424
rect 59813 421 59825 424
rect 59983 421 59995 424
rect 59813 420 59866 421
rect 59824 412 59866 420
rect 59707 400 59718 412
rect 58988 341 58992 395
rect 59048 387 59094 395
rect 59048 383 59064 387
rect 59056 380 59064 383
rect 59090 380 59094 387
rect 59098 383 59106 395
rect 59454 383 59462 395
rect 59466 387 59500 395
rect 59466 380 59470 387
rect 59496 380 59500 387
rect 59504 383 59512 395
rect 59044 379 59110 380
rect 59450 379 59516 380
rect 59056 371 59060 379
rect 59110 365 59160 367
rect 59400 365 59450 367
rect 59150 361 59204 365
rect 59356 361 59410 365
rect 59150 356 59170 361
rect 59390 356 59410 361
rect 59160 341 59162 356
rect 58988 261 58992 329
rect 59056 305 59060 341
rect 59154 331 59162 341
rect 59170 331 59171 351
rect 59160 315 59162 331
rect 59181 322 59184 356
rect 59203 331 59204 351
rect 59213 331 59220 341
rect 59340 331 59347 341
rect 59356 331 59357 351
rect 59376 322 59379 356
rect 59389 331 59390 351
rect 59399 331 59406 341
rect 59170 315 59186 321
rect 59188 315 59204 321
rect 59356 315 59372 321
rect 59374 315 59390 321
rect 59450 315 59452 365
rect 58993 267 59029 295
rect 58993 261 59007 267
rect 58672 212 58683 213
rect 58517 183 58524 207
rect 58672 183 58682 212
rect 58763 207 58775 241
rect 58785 207 58805 241
rect 58508 103 58512 171
rect 58576 133 58580 183
rect 58576 98 58580 103
rect 58327 62 58332 96
rect 58356 62 58361 96
rect 58576 94 58614 98
rect 58576 79 58584 94
rect 58610 79 58614 94
rect 58698 94 58732 98
rect 58698 79 58702 94
rect 58728 79 58732 94
rect 58576 61 58618 79
rect 58694 61 58736 79
rect 58554 55 58640 61
rect 58672 55 58758 61
rect 58800 55 58804 207
rect 58830 183 58837 211
rect 58988 183 58992 251
rect 58997 233 59007 261
rect 59017 261 59031 267
rect 59056 261 59067 305
rect 59493 267 59504 305
rect 59531 267 59567 295
rect 59568 267 59572 395
rect 59719 378 59724 412
rect 59748 378 59753 412
rect 59754 400 59765 412
rect 59779 400 59790 412
rect 59791 395 59866 412
rect 59942 420 59995 421
rect 60005 420 60017 424
rect 60055 420 60067 424
rect 60077 420 60089 424
rect 59942 412 59984 420
rect 59942 395 60017 412
rect 60018 400 60029 412
rect 60043 400 60054 412
rect 59756 341 59760 395
rect 59791 378 59862 395
rect 59866 383 59874 395
rect 59934 383 59942 395
rect 59946 378 59980 395
rect 59983 378 60017 395
rect 59824 371 59828 378
rect 59218 262 59268 264
rect 59292 262 59342 264
rect 59017 233 59037 261
rect 59056 233 59065 261
rect 59119 253 59153 261
rect 59098 246 59153 253
rect 59119 245 59153 246
rect 59221 253 59252 261
rect 59221 245 59255 253
rect 59056 213 59060 233
rect 59252 229 59255 245
rect 59119 228 59153 229
rect 59098 221 59153 228
rect 59221 221 59255 229
rect 59268 212 59270 262
rect 59308 253 59339 261
rect 59342 253 59344 262
rect 59531 261 59543 267
rect 59308 245 59344 253
rect 59407 253 59441 261
rect 59407 246 59462 253
rect 59407 245 59441 246
rect 59339 229 59344 245
rect 59533 233 59543 261
rect 59553 233 59573 267
rect 59756 261 59760 329
rect 59824 291 59828 341
rect 59824 251 59833 279
rect 59920 264 59930 291
rect 59879 262 59930 264
rect 59920 261 59931 262
rect 59887 253 59921 261
rect 59929 253 59931 261
rect 59308 221 59344 229
rect 59407 228 59441 229
rect 59407 221 59462 228
rect 59342 212 59344 221
rect 58988 103 58992 171
rect 59056 133 59060 183
rect 59110 159 59160 161
rect 59400 159 59450 161
rect 59160 143 59162 159
rect 59170 153 59186 159
rect 59188 153 59204 159
rect 59356 153 59372 159
rect 59374 153 59390 159
rect 59181 143 59204 152
rect 59356 143 59379 152
rect 59154 133 59162 143
rect 59160 109 59162 133
rect 59170 123 59171 143
rect 59181 118 59184 143
rect 59203 123 59204 143
rect 59213 133 59220 143
rect 59340 133 59347 143
rect 59356 123 59357 143
rect 59376 118 59379 143
rect 59389 123 59390 143
rect 59399 133 59406 143
rect 59170 109 59204 113
rect 59356 109 59390 113
rect 59450 109 59452 159
rect 59056 103 59098 104
rect 59462 103 59504 104
rect 59056 96 59060 103
rect 58951 62 58956 96
rect 58980 62 58985 96
rect 59023 79 59094 96
rect 59466 79 59500 96
rect 59503 79 59537 96
rect 59023 62 59098 79
rect 59056 61 59098 62
rect 59462 62 59537 79
rect 59462 61 59504 62
rect 59034 55 59120 61
rect 59440 55 59526 61
rect 59568 55 59572 233
rect 59756 183 59760 251
rect 59765 207 59775 241
rect 59785 213 59805 241
rect 59785 207 59799 213
rect 59824 207 59835 251
rect 59866 246 59942 253
rect 59975 251 59984 279
rect 59887 228 59921 246
rect 59929 228 59931 246
rect 59866 221 59942 228
rect 59929 213 59931 221
rect 59973 213 59984 251
rect 60048 241 60052 395
rect 60055 378 60060 412
rect 60084 378 60089 412
rect 60090 400 60101 412
rect 60304 395 60346 421
rect 60710 395 60752 421
rect 60967 420 60979 424
rect 60989 420 61001 424
rect 61039 420 61051 424
rect 61061 421 61073 424
rect 61231 421 61243 424
rect 61061 420 61114 421
rect 61072 412 61114 420
rect 60955 400 60966 412
rect 60236 341 60240 395
rect 60296 387 60342 395
rect 60296 383 60312 387
rect 60304 380 60312 383
rect 60338 380 60342 387
rect 60346 383 60354 395
rect 60702 383 60710 395
rect 60714 387 60748 395
rect 60714 380 60718 387
rect 60744 380 60748 387
rect 60752 383 60760 395
rect 60292 379 60358 380
rect 60698 379 60764 380
rect 60304 371 60308 379
rect 60358 365 60408 367
rect 60648 365 60698 367
rect 60398 361 60452 365
rect 60604 361 60658 365
rect 60398 356 60418 361
rect 60638 356 60658 361
rect 60408 341 60410 356
rect 60236 261 60240 329
rect 60304 305 60308 341
rect 60402 331 60410 341
rect 60418 331 60419 351
rect 60408 315 60410 331
rect 60429 322 60432 356
rect 60451 331 60452 351
rect 60461 331 60468 341
rect 60588 331 60595 341
rect 60604 331 60605 351
rect 60624 322 60627 356
rect 60637 331 60638 351
rect 60647 331 60654 341
rect 60418 315 60434 321
rect 60436 315 60452 321
rect 60604 315 60620 321
rect 60622 315 60638 321
rect 60698 315 60700 365
rect 60241 267 60277 295
rect 60241 261 60255 267
rect 59920 212 59931 213
rect 59765 183 59772 207
rect 59920 183 59930 212
rect 60011 207 60023 241
rect 60033 207 60053 241
rect 59756 103 59760 171
rect 59824 133 59828 183
rect 59824 98 59828 103
rect 59575 62 59580 96
rect 59604 62 59609 96
rect 59824 94 59862 98
rect 59824 79 59832 94
rect 59858 79 59862 94
rect 59946 94 59980 98
rect 59946 79 59950 94
rect 59976 79 59980 94
rect 59824 61 59866 79
rect 59942 61 59984 79
rect 59802 55 59888 61
rect 59920 55 60006 61
rect 60048 55 60052 207
rect 60078 183 60085 211
rect 60236 183 60240 251
rect 60245 233 60255 261
rect 60265 261 60279 267
rect 60304 261 60315 305
rect 60741 267 60752 305
rect 60779 267 60815 295
rect 60816 267 60820 395
rect 60967 378 60972 412
rect 60996 378 61001 412
rect 61002 400 61013 412
rect 61027 400 61038 412
rect 61039 395 61114 412
rect 61190 420 61243 421
rect 61253 420 61265 424
rect 61303 420 61315 424
rect 61325 420 61337 424
rect 61190 412 61232 420
rect 61190 395 61265 412
rect 61266 400 61277 412
rect 61291 400 61302 412
rect 61004 341 61008 395
rect 61039 378 61110 395
rect 61114 383 61122 395
rect 61182 383 61190 395
rect 61194 378 61228 395
rect 61231 378 61265 395
rect 61072 371 61076 378
rect 60466 262 60516 264
rect 60540 262 60590 264
rect 60265 233 60285 261
rect 60304 233 60313 261
rect 60367 253 60401 261
rect 60346 246 60401 253
rect 60367 245 60401 246
rect 60469 253 60500 261
rect 60469 245 60503 253
rect 60304 213 60308 233
rect 60500 229 60503 245
rect 60367 228 60401 229
rect 60346 221 60401 228
rect 60469 221 60503 229
rect 60516 212 60518 262
rect 60556 253 60587 261
rect 60590 253 60592 262
rect 60779 261 60791 267
rect 60556 245 60592 253
rect 60655 253 60689 261
rect 60655 246 60710 253
rect 60655 245 60689 246
rect 60587 229 60592 245
rect 60781 233 60791 261
rect 60801 233 60821 267
rect 61004 261 61008 329
rect 61072 291 61076 341
rect 61072 251 61081 279
rect 61168 264 61178 291
rect 61127 262 61178 264
rect 61168 261 61179 262
rect 61135 253 61169 261
rect 61177 253 61179 261
rect 60556 221 60592 229
rect 60655 228 60689 229
rect 60655 221 60710 228
rect 60590 212 60592 221
rect 60236 103 60240 171
rect 60304 133 60308 183
rect 60358 159 60408 161
rect 60648 159 60698 161
rect 60408 143 60410 159
rect 60418 153 60434 159
rect 60436 153 60452 159
rect 60604 153 60620 159
rect 60622 153 60638 159
rect 60429 143 60452 152
rect 60604 143 60627 152
rect 60402 133 60410 143
rect 60408 109 60410 133
rect 60418 123 60419 143
rect 60429 118 60432 143
rect 60451 123 60452 143
rect 60461 133 60468 143
rect 60588 133 60595 143
rect 60604 123 60605 143
rect 60624 118 60627 143
rect 60637 123 60638 143
rect 60647 133 60654 143
rect 60418 109 60452 113
rect 60604 109 60638 113
rect 60698 109 60700 159
rect 60304 103 60346 104
rect 60710 103 60752 104
rect 60304 96 60308 103
rect 60199 62 60204 96
rect 60228 62 60233 96
rect 60271 79 60342 96
rect 60714 79 60748 96
rect 60751 79 60785 96
rect 60271 62 60346 79
rect 60304 61 60346 62
rect 60710 62 60785 79
rect 60710 61 60752 62
rect 60282 55 60368 61
rect 60688 55 60774 61
rect 60816 55 60820 233
rect 61004 183 61008 251
rect 61013 207 61023 241
rect 61033 213 61053 241
rect 61033 207 61047 213
rect 61072 207 61083 251
rect 61114 246 61190 253
rect 61223 251 61232 279
rect 61135 228 61169 246
rect 61177 228 61179 246
rect 61114 221 61190 228
rect 61177 213 61179 221
rect 61221 213 61232 251
rect 61296 241 61300 395
rect 61303 378 61308 412
rect 61332 378 61337 412
rect 61338 400 61349 412
rect 61552 395 61594 421
rect 61958 395 62000 421
rect 62215 420 62227 424
rect 62237 420 62249 424
rect 62287 420 62299 424
rect 62309 421 62321 424
rect 62479 421 62491 424
rect 62309 420 62362 421
rect 62320 412 62362 420
rect 62203 400 62214 412
rect 61484 341 61488 395
rect 61544 387 61590 395
rect 61544 383 61560 387
rect 61552 380 61560 383
rect 61586 380 61590 387
rect 61594 383 61602 395
rect 61950 383 61958 395
rect 61962 387 61996 395
rect 61962 380 61966 387
rect 61992 380 61996 387
rect 62000 383 62008 395
rect 61540 379 61606 380
rect 61946 379 62012 380
rect 61552 371 61556 379
rect 61606 365 61656 367
rect 61896 365 61946 367
rect 61646 361 61700 365
rect 61852 361 61906 365
rect 61646 356 61666 361
rect 61886 356 61906 361
rect 61656 341 61658 356
rect 61484 261 61488 329
rect 61552 305 61556 341
rect 61650 331 61658 341
rect 61666 331 61667 351
rect 61656 315 61658 331
rect 61677 322 61680 356
rect 61699 331 61700 351
rect 61709 331 61716 341
rect 61836 331 61843 341
rect 61852 331 61853 351
rect 61872 322 61875 356
rect 61885 331 61886 351
rect 61895 331 61902 341
rect 61666 315 61682 321
rect 61684 315 61700 321
rect 61852 315 61868 321
rect 61870 315 61886 321
rect 61946 315 61948 365
rect 61489 267 61525 295
rect 61489 261 61503 267
rect 61168 212 61179 213
rect 61013 183 61020 207
rect 61168 183 61178 212
rect 61259 207 61271 241
rect 61281 207 61301 241
rect 61004 103 61008 171
rect 61072 133 61076 183
rect 61072 98 61076 103
rect 60823 62 60828 96
rect 60852 62 60857 96
rect 61072 94 61110 98
rect 61072 79 61080 94
rect 61106 79 61110 94
rect 61194 94 61228 98
rect 61194 79 61198 94
rect 61224 79 61228 94
rect 61072 61 61114 79
rect 61190 61 61232 79
rect 61050 55 61136 61
rect 61168 55 61254 61
rect 61296 55 61300 207
rect 61326 183 61333 211
rect 61484 183 61488 251
rect 61493 233 61503 261
rect 61513 261 61527 267
rect 61552 261 61563 305
rect 61989 267 62000 305
rect 62027 267 62063 295
rect 62064 267 62068 395
rect 62215 378 62220 412
rect 62244 378 62249 412
rect 62250 400 62261 412
rect 62275 400 62286 412
rect 62287 395 62362 412
rect 62438 420 62491 421
rect 62501 420 62513 424
rect 62551 420 62563 424
rect 62573 420 62585 424
rect 62438 412 62480 420
rect 62438 395 62513 412
rect 62514 400 62525 412
rect 62539 400 62550 412
rect 62252 341 62256 395
rect 62287 378 62358 395
rect 62362 383 62370 395
rect 62430 383 62438 395
rect 62442 378 62476 395
rect 62479 378 62513 395
rect 62320 371 62324 378
rect 61714 262 61764 264
rect 61788 262 61838 264
rect 61513 233 61533 261
rect 61552 233 61561 261
rect 61615 253 61649 261
rect 61594 246 61649 253
rect 61615 245 61649 246
rect 61717 253 61748 261
rect 61717 245 61751 253
rect 61552 213 61556 233
rect 61748 229 61751 245
rect 61615 228 61649 229
rect 61594 221 61649 228
rect 61717 221 61751 229
rect 61764 212 61766 262
rect 61804 253 61835 261
rect 61838 253 61840 262
rect 62027 261 62039 267
rect 61804 245 61840 253
rect 61903 253 61937 261
rect 61903 246 61958 253
rect 61903 245 61937 246
rect 61835 229 61840 245
rect 62029 233 62039 261
rect 62049 233 62069 267
rect 62252 261 62256 329
rect 62320 291 62324 341
rect 62320 251 62329 279
rect 62416 264 62426 291
rect 62375 262 62426 264
rect 62416 261 62427 262
rect 62383 253 62417 261
rect 62425 253 62427 261
rect 61804 221 61840 229
rect 61903 228 61937 229
rect 61903 221 61958 228
rect 61838 212 61840 221
rect 61484 103 61488 171
rect 61552 133 61556 183
rect 61606 159 61656 161
rect 61896 159 61946 161
rect 61656 143 61658 159
rect 61666 153 61682 159
rect 61684 153 61700 159
rect 61852 153 61868 159
rect 61870 153 61886 159
rect 61677 143 61700 152
rect 61852 143 61875 152
rect 61650 133 61658 143
rect 61656 109 61658 133
rect 61666 123 61667 143
rect 61677 118 61680 143
rect 61699 123 61700 143
rect 61709 133 61716 143
rect 61836 133 61843 143
rect 61852 123 61853 143
rect 61872 118 61875 143
rect 61885 123 61886 143
rect 61895 133 61902 143
rect 61666 109 61700 113
rect 61852 109 61886 113
rect 61946 109 61948 159
rect 61552 103 61594 104
rect 61958 103 62000 104
rect 61552 96 61556 103
rect 61447 62 61452 96
rect 61476 62 61481 96
rect 61519 79 61590 96
rect 61962 79 61996 96
rect 61999 79 62033 96
rect 61519 62 61594 79
rect 61552 61 61594 62
rect 61958 62 62033 79
rect 61958 61 62000 62
rect 61530 55 61616 61
rect 61936 55 62022 61
rect 62064 55 62068 233
rect 62252 183 62256 251
rect 62261 207 62271 241
rect 62281 213 62301 241
rect 62281 207 62295 213
rect 62320 207 62331 251
rect 62362 246 62438 253
rect 62471 251 62480 279
rect 62383 228 62417 246
rect 62425 228 62427 246
rect 62362 221 62438 228
rect 62425 213 62427 221
rect 62469 213 62480 251
rect 62544 241 62548 395
rect 62551 378 62556 412
rect 62580 378 62585 412
rect 62586 400 62597 412
rect 62800 395 62842 421
rect 63206 395 63248 421
rect 63463 420 63475 424
rect 63485 420 63497 424
rect 63535 420 63547 424
rect 63557 421 63569 424
rect 63727 421 63739 424
rect 63557 420 63610 421
rect 63568 412 63610 420
rect 63451 400 63462 412
rect 62732 341 62736 395
rect 62792 387 62838 395
rect 62792 383 62808 387
rect 62800 380 62808 383
rect 62834 380 62838 387
rect 62842 383 62850 395
rect 63198 383 63206 395
rect 63210 387 63244 395
rect 63210 380 63214 387
rect 63240 380 63244 387
rect 63248 383 63256 395
rect 62788 379 62854 380
rect 63194 379 63260 380
rect 62800 371 62804 379
rect 62854 365 62904 367
rect 63144 365 63194 367
rect 62894 361 62948 365
rect 63100 361 63154 365
rect 62894 356 62914 361
rect 63134 356 63154 361
rect 62904 341 62906 356
rect 62732 261 62736 329
rect 62800 305 62804 341
rect 62898 331 62906 341
rect 62914 331 62915 351
rect 62904 315 62906 331
rect 62925 322 62928 356
rect 62947 331 62948 351
rect 62957 331 62964 341
rect 63084 331 63091 341
rect 63100 331 63101 351
rect 63120 322 63123 356
rect 63133 331 63134 351
rect 63143 331 63150 341
rect 62914 315 62930 321
rect 62932 315 62948 321
rect 63100 315 63116 321
rect 63118 315 63134 321
rect 63194 315 63196 365
rect 62737 267 62773 295
rect 62737 261 62751 267
rect 62416 212 62427 213
rect 62261 183 62268 207
rect 62416 183 62426 212
rect 62507 207 62519 241
rect 62529 207 62549 241
rect 62252 103 62256 171
rect 62320 133 62324 183
rect 62320 98 62324 103
rect 62071 62 62076 96
rect 62100 62 62105 96
rect 62320 94 62358 98
rect 62320 79 62328 94
rect 62354 79 62358 94
rect 62442 94 62476 98
rect 62442 79 62446 94
rect 62472 79 62476 94
rect 62320 61 62362 79
rect 62438 61 62480 79
rect 62298 55 62384 61
rect 62416 55 62502 61
rect 62544 55 62548 207
rect 62574 183 62581 211
rect 62732 183 62736 251
rect 62741 233 62751 261
rect 62761 261 62775 267
rect 62800 261 62811 305
rect 63237 267 63248 305
rect 63275 267 63311 295
rect 63312 267 63316 395
rect 63463 378 63468 412
rect 63492 378 63497 412
rect 63498 400 63509 412
rect 63523 400 63534 412
rect 63535 395 63610 412
rect 63686 420 63739 421
rect 63749 420 63761 424
rect 63799 420 63811 424
rect 63821 420 63833 424
rect 63686 412 63728 420
rect 63686 395 63761 412
rect 63762 400 63773 412
rect 63787 400 63798 412
rect 63500 341 63504 395
rect 63535 378 63606 395
rect 63610 383 63618 395
rect 63678 383 63686 395
rect 63690 378 63724 395
rect 63727 378 63761 395
rect 63568 371 63572 378
rect 62962 262 63012 264
rect 63036 262 63086 264
rect 62761 233 62781 261
rect 62800 233 62809 261
rect 62863 253 62897 261
rect 62842 246 62897 253
rect 62863 245 62897 246
rect 62965 253 62996 261
rect 62965 245 62999 253
rect 62800 213 62804 233
rect 62996 229 62999 245
rect 62863 228 62897 229
rect 62842 221 62897 228
rect 62965 221 62999 229
rect 63012 212 63014 262
rect 63052 253 63083 261
rect 63086 253 63088 262
rect 63275 261 63287 267
rect 63052 245 63088 253
rect 63151 253 63185 261
rect 63151 246 63206 253
rect 63151 245 63185 246
rect 63083 229 63088 245
rect 63277 233 63287 261
rect 63297 233 63317 267
rect 63500 261 63504 329
rect 63568 291 63572 341
rect 63568 251 63577 279
rect 63664 264 63674 291
rect 63623 262 63674 264
rect 63664 261 63675 262
rect 63631 253 63665 261
rect 63673 253 63675 261
rect 63052 221 63088 229
rect 63151 228 63185 229
rect 63151 221 63206 228
rect 63086 212 63088 221
rect 62732 103 62736 171
rect 62800 133 62804 183
rect 62854 159 62904 161
rect 63144 159 63194 161
rect 62904 143 62906 159
rect 62914 153 62930 159
rect 62932 153 62948 159
rect 63100 153 63116 159
rect 63118 153 63134 159
rect 62925 143 62948 152
rect 63100 143 63123 152
rect 62898 133 62906 143
rect 62904 109 62906 133
rect 62914 123 62915 143
rect 62925 118 62928 143
rect 62947 123 62948 143
rect 62957 133 62964 143
rect 63084 133 63091 143
rect 63100 123 63101 143
rect 63120 118 63123 143
rect 63133 123 63134 143
rect 63143 133 63150 143
rect 62914 109 62948 113
rect 63100 109 63134 113
rect 63194 109 63196 159
rect 62800 103 62842 104
rect 63206 103 63248 104
rect 62800 96 62804 103
rect 62695 62 62700 96
rect 62724 62 62729 96
rect 62767 79 62838 96
rect 63210 79 63244 96
rect 63247 79 63281 96
rect 62767 62 62842 79
rect 62800 61 62842 62
rect 63206 62 63281 79
rect 63206 61 63248 62
rect 62778 55 62864 61
rect 63184 55 63270 61
rect 63312 55 63316 233
rect 63500 183 63504 251
rect 63509 207 63519 241
rect 63529 213 63549 241
rect 63529 207 63543 213
rect 63568 207 63579 251
rect 63610 246 63686 253
rect 63719 251 63728 279
rect 63631 228 63665 246
rect 63673 228 63675 246
rect 63610 221 63686 228
rect 63673 213 63675 221
rect 63717 213 63728 251
rect 63792 241 63796 395
rect 63799 378 63804 412
rect 63828 378 63833 412
rect 63834 400 63845 412
rect 64048 395 64090 421
rect 64454 395 64496 421
rect 64711 420 64723 424
rect 64733 420 64745 424
rect 64783 420 64795 424
rect 64805 421 64817 424
rect 64975 421 64987 424
rect 64805 420 64858 421
rect 64816 412 64858 420
rect 64699 400 64710 412
rect 63980 341 63984 395
rect 64040 387 64086 395
rect 64040 383 64056 387
rect 64048 380 64056 383
rect 64082 380 64086 387
rect 64090 383 64098 395
rect 64446 383 64454 395
rect 64458 387 64492 395
rect 64458 380 64462 387
rect 64488 380 64492 387
rect 64496 383 64504 395
rect 64036 379 64102 380
rect 64442 379 64508 380
rect 64048 371 64052 379
rect 64102 365 64152 367
rect 64392 365 64442 367
rect 64142 361 64196 365
rect 64348 361 64402 365
rect 64142 356 64162 361
rect 64382 356 64402 361
rect 64152 341 64154 356
rect 63980 261 63984 329
rect 64048 305 64052 341
rect 64146 331 64154 341
rect 64162 331 64163 351
rect 64152 315 64154 331
rect 64173 322 64176 356
rect 64195 331 64196 351
rect 64205 331 64212 341
rect 64332 331 64339 341
rect 64348 331 64349 351
rect 64368 322 64371 356
rect 64381 331 64382 351
rect 64391 331 64398 341
rect 64162 315 64178 321
rect 64180 315 64196 321
rect 64348 315 64364 321
rect 64366 315 64382 321
rect 64442 315 64444 365
rect 63985 267 64021 295
rect 63985 261 63999 267
rect 63664 212 63675 213
rect 63509 183 63516 207
rect 63664 183 63674 212
rect 63755 207 63767 241
rect 63777 207 63797 241
rect 63500 103 63504 171
rect 63568 133 63572 183
rect 63568 98 63572 103
rect 63319 62 63324 96
rect 63348 62 63353 96
rect 63568 94 63606 98
rect 63568 79 63576 94
rect 63602 79 63606 94
rect 63690 94 63724 98
rect 63690 79 63694 94
rect 63720 79 63724 94
rect 63568 61 63610 79
rect 63686 61 63728 79
rect 63546 55 63632 61
rect 63664 55 63750 61
rect 63792 55 63796 207
rect 63822 183 63829 211
rect 63980 183 63984 251
rect 63989 233 63999 261
rect 64009 261 64023 267
rect 64048 261 64059 305
rect 64485 267 64496 305
rect 64523 267 64559 295
rect 64560 267 64564 395
rect 64711 378 64716 412
rect 64740 378 64745 412
rect 64746 400 64757 412
rect 64771 400 64782 412
rect 64783 395 64858 412
rect 64934 420 64987 421
rect 64997 420 65009 424
rect 65047 420 65059 424
rect 65069 420 65081 424
rect 64934 412 64976 420
rect 64934 395 65009 412
rect 65010 400 65021 412
rect 65035 400 65046 412
rect 64748 341 64752 395
rect 64783 378 64854 395
rect 64858 383 64866 395
rect 64926 383 64934 395
rect 64938 378 64972 395
rect 64975 378 65009 395
rect 64816 371 64820 378
rect 64210 262 64260 264
rect 64284 262 64334 264
rect 64009 233 64029 261
rect 64048 233 64057 261
rect 64111 253 64145 261
rect 64090 246 64145 253
rect 64111 245 64145 246
rect 64213 253 64244 261
rect 64213 245 64247 253
rect 64048 213 64052 233
rect 64244 229 64247 245
rect 64111 228 64145 229
rect 64090 221 64145 228
rect 64213 221 64247 229
rect 64260 212 64262 262
rect 64300 253 64331 261
rect 64334 253 64336 262
rect 64523 261 64535 267
rect 64300 245 64336 253
rect 64399 253 64433 261
rect 64399 246 64454 253
rect 64399 245 64433 246
rect 64331 229 64336 245
rect 64525 233 64535 261
rect 64545 233 64565 267
rect 64748 261 64752 329
rect 64816 291 64820 341
rect 64816 251 64825 279
rect 64912 264 64922 291
rect 64871 262 64922 264
rect 64912 261 64923 262
rect 64879 253 64913 261
rect 64921 253 64923 261
rect 64300 221 64336 229
rect 64399 228 64433 229
rect 64399 221 64454 228
rect 64334 212 64336 221
rect 63980 103 63984 171
rect 64048 133 64052 183
rect 64102 159 64152 161
rect 64392 159 64442 161
rect 64152 143 64154 159
rect 64162 153 64178 159
rect 64180 153 64196 159
rect 64348 153 64364 159
rect 64366 153 64382 159
rect 64173 143 64196 152
rect 64348 143 64371 152
rect 64146 133 64154 143
rect 64152 109 64154 133
rect 64162 123 64163 143
rect 64173 118 64176 143
rect 64195 123 64196 143
rect 64205 133 64212 143
rect 64332 133 64339 143
rect 64348 123 64349 143
rect 64368 118 64371 143
rect 64381 123 64382 143
rect 64391 133 64398 143
rect 64162 109 64196 113
rect 64348 109 64382 113
rect 64442 109 64444 159
rect 64048 103 64090 104
rect 64454 103 64496 104
rect 64048 96 64052 103
rect 63943 62 63948 96
rect 63972 62 63977 96
rect 64015 79 64086 96
rect 64458 79 64492 96
rect 64495 79 64529 96
rect 64015 62 64090 79
rect 64048 61 64090 62
rect 64454 62 64529 79
rect 64454 61 64496 62
rect 64026 55 64112 61
rect 64432 55 64518 61
rect 64560 55 64564 233
rect 64748 183 64752 251
rect 64757 207 64767 241
rect 64777 213 64797 241
rect 64777 207 64791 213
rect 64816 207 64827 251
rect 64858 246 64934 253
rect 64967 251 64976 279
rect 64879 228 64913 246
rect 64921 228 64923 246
rect 64858 221 64934 228
rect 64921 213 64923 221
rect 64965 213 64976 251
rect 65040 241 65044 395
rect 65047 378 65052 412
rect 65076 378 65081 412
rect 65082 400 65093 412
rect 65296 395 65338 421
rect 65702 395 65744 421
rect 65959 420 65971 424
rect 65981 420 65993 424
rect 66031 420 66043 424
rect 66053 421 66065 424
rect 66223 421 66235 424
rect 66053 420 66106 421
rect 66064 412 66106 420
rect 65947 400 65958 412
rect 65228 341 65232 395
rect 65288 387 65334 395
rect 65288 383 65304 387
rect 65296 380 65304 383
rect 65330 380 65334 387
rect 65338 383 65346 395
rect 65694 383 65702 395
rect 65706 387 65740 395
rect 65706 380 65710 387
rect 65736 380 65740 387
rect 65744 383 65752 395
rect 65284 379 65350 380
rect 65690 379 65756 380
rect 65296 371 65300 379
rect 65350 365 65400 367
rect 65640 365 65690 367
rect 65390 361 65444 365
rect 65596 361 65650 365
rect 65390 356 65410 361
rect 65630 356 65650 361
rect 65400 341 65402 356
rect 65228 261 65232 329
rect 65296 305 65300 341
rect 65394 331 65402 341
rect 65410 331 65411 351
rect 65400 315 65402 331
rect 65421 322 65424 356
rect 65443 331 65444 351
rect 65453 331 65460 341
rect 65580 331 65587 341
rect 65596 331 65597 351
rect 65616 322 65619 356
rect 65629 331 65630 351
rect 65639 331 65646 341
rect 65410 315 65426 321
rect 65428 315 65444 321
rect 65596 315 65612 321
rect 65614 315 65630 321
rect 65690 315 65692 365
rect 65233 267 65269 295
rect 65233 261 65247 267
rect 64912 212 64923 213
rect 64757 183 64764 207
rect 64912 183 64922 212
rect 65003 207 65015 241
rect 65025 207 65045 241
rect 64748 103 64752 171
rect 64816 133 64820 183
rect 64816 98 64820 103
rect 64567 62 64572 96
rect 64596 62 64601 96
rect 64816 94 64854 98
rect 64816 79 64824 94
rect 64850 79 64854 94
rect 64938 94 64972 98
rect 64938 79 64942 94
rect 64968 79 64972 94
rect 64816 61 64858 79
rect 64934 61 64976 79
rect 64794 55 64880 61
rect 64912 55 64998 61
rect 65040 55 65044 207
rect 65070 183 65077 211
rect 65228 183 65232 251
rect 65237 233 65247 261
rect 65257 261 65271 267
rect 65296 261 65307 305
rect 65733 267 65744 305
rect 65771 267 65807 295
rect 65808 267 65812 395
rect 65959 378 65964 412
rect 65988 378 65993 412
rect 65994 400 66005 412
rect 66019 400 66030 412
rect 66031 395 66106 412
rect 66182 420 66235 421
rect 66245 420 66257 424
rect 66295 420 66307 424
rect 66317 420 66329 424
rect 66182 412 66224 420
rect 66182 395 66257 412
rect 66258 400 66269 412
rect 66283 400 66294 412
rect 65996 341 66000 395
rect 66031 378 66102 395
rect 66106 383 66114 395
rect 66174 383 66182 395
rect 66186 378 66220 395
rect 66223 378 66257 395
rect 66064 371 66068 378
rect 65458 262 65508 264
rect 65532 262 65582 264
rect 65257 233 65277 261
rect 65296 233 65305 261
rect 65359 253 65393 261
rect 65338 246 65393 253
rect 65359 245 65393 246
rect 65461 253 65492 261
rect 65461 245 65495 253
rect 65296 213 65300 233
rect 65492 229 65495 245
rect 65359 228 65393 229
rect 65338 221 65393 228
rect 65461 221 65495 229
rect 65508 212 65510 262
rect 65548 253 65579 261
rect 65582 253 65584 262
rect 65771 261 65783 267
rect 65548 245 65584 253
rect 65647 253 65681 261
rect 65647 246 65702 253
rect 65647 245 65681 246
rect 65579 229 65584 245
rect 65773 233 65783 261
rect 65793 233 65813 267
rect 65996 261 66000 329
rect 66064 291 66068 341
rect 66064 251 66073 279
rect 66160 264 66170 291
rect 66119 262 66170 264
rect 66160 261 66171 262
rect 66127 253 66161 261
rect 66169 253 66171 261
rect 65548 221 65584 229
rect 65647 228 65681 229
rect 65647 221 65702 228
rect 65582 212 65584 221
rect 65228 103 65232 171
rect 65296 133 65300 183
rect 65350 159 65400 161
rect 65640 159 65690 161
rect 65400 143 65402 159
rect 65410 153 65426 159
rect 65428 153 65444 159
rect 65596 153 65612 159
rect 65614 153 65630 159
rect 65421 143 65444 152
rect 65596 143 65619 152
rect 65394 133 65402 143
rect 65400 109 65402 133
rect 65410 123 65411 143
rect 65421 118 65424 143
rect 65443 123 65444 143
rect 65453 133 65460 143
rect 65580 133 65587 143
rect 65596 123 65597 143
rect 65616 118 65619 143
rect 65629 123 65630 143
rect 65639 133 65646 143
rect 65410 109 65444 113
rect 65596 109 65630 113
rect 65690 109 65692 159
rect 65296 103 65338 104
rect 65702 103 65744 104
rect 65296 96 65300 103
rect 65191 62 65196 96
rect 65220 62 65225 96
rect 65263 79 65334 96
rect 65706 79 65740 96
rect 65743 79 65777 96
rect 65263 62 65338 79
rect 65296 61 65338 62
rect 65702 62 65777 79
rect 65702 61 65744 62
rect 65274 55 65360 61
rect 65680 55 65766 61
rect 65808 55 65812 233
rect 65996 183 66000 251
rect 66005 207 66015 241
rect 66025 213 66045 241
rect 66025 207 66039 213
rect 66064 207 66075 251
rect 66106 246 66182 253
rect 66215 251 66224 279
rect 66127 228 66161 246
rect 66169 228 66171 246
rect 66106 221 66182 228
rect 66169 213 66171 221
rect 66213 213 66224 251
rect 66288 241 66292 395
rect 66295 378 66300 412
rect 66324 378 66329 412
rect 66330 400 66341 412
rect 66544 395 66586 421
rect 66950 395 66992 421
rect 67207 420 67219 424
rect 67229 420 67241 424
rect 67279 420 67291 424
rect 67301 421 67313 424
rect 67471 421 67483 424
rect 67301 420 67354 421
rect 67312 412 67354 420
rect 67195 400 67206 412
rect 66476 341 66480 395
rect 66536 387 66582 395
rect 66536 383 66552 387
rect 66544 380 66552 383
rect 66578 380 66582 387
rect 66586 383 66594 395
rect 66942 383 66950 395
rect 66954 387 66988 395
rect 66954 380 66958 387
rect 66984 380 66988 387
rect 66992 383 67000 395
rect 66532 379 66598 380
rect 66938 379 67004 380
rect 66544 371 66548 379
rect 66598 365 66648 367
rect 66888 365 66938 367
rect 66638 361 66692 365
rect 66844 361 66898 365
rect 66638 356 66658 361
rect 66878 356 66898 361
rect 66648 341 66650 356
rect 66476 261 66480 329
rect 66544 305 66548 341
rect 66642 331 66650 341
rect 66658 331 66659 351
rect 66648 315 66650 331
rect 66669 322 66672 356
rect 66691 331 66692 351
rect 66701 331 66708 341
rect 66828 331 66835 341
rect 66844 331 66845 351
rect 66864 322 66867 356
rect 66877 331 66878 351
rect 66887 331 66894 341
rect 66658 315 66674 321
rect 66676 315 66692 321
rect 66844 315 66860 321
rect 66862 315 66878 321
rect 66938 315 66940 365
rect 66481 267 66517 295
rect 66481 261 66495 267
rect 66160 212 66171 213
rect 66005 183 66012 207
rect 66160 183 66170 212
rect 66251 207 66263 241
rect 66273 207 66293 241
rect 65996 103 66000 171
rect 66064 133 66068 183
rect 66064 98 66068 103
rect 65815 62 65820 96
rect 65844 62 65849 96
rect 66064 94 66102 98
rect 66064 79 66072 94
rect 66098 79 66102 94
rect 66186 94 66220 98
rect 66186 79 66190 94
rect 66216 79 66220 94
rect 66064 61 66106 79
rect 66182 61 66224 79
rect 66042 55 66128 61
rect 66160 55 66246 61
rect 66288 55 66292 207
rect 66318 183 66325 211
rect 66476 183 66480 251
rect 66485 233 66495 261
rect 66505 261 66519 267
rect 66544 261 66555 305
rect 66981 267 66992 305
rect 67019 267 67055 295
rect 67056 267 67060 395
rect 67207 378 67212 412
rect 67236 378 67241 412
rect 67242 400 67253 412
rect 67267 400 67278 412
rect 67279 395 67354 412
rect 67430 420 67483 421
rect 67493 420 67505 424
rect 67543 420 67555 424
rect 67565 420 67577 424
rect 67430 412 67472 420
rect 67430 395 67505 412
rect 67506 400 67517 412
rect 67531 400 67542 412
rect 67244 341 67248 395
rect 67279 378 67350 395
rect 67354 383 67362 395
rect 67422 383 67430 395
rect 67434 378 67468 395
rect 67471 378 67505 395
rect 67312 371 67316 378
rect 66706 262 66756 264
rect 66780 262 66830 264
rect 66505 233 66525 261
rect 66544 233 66553 261
rect 66607 253 66641 261
rect 66586 246 66641 253
rect 66607 245 66641 246
rect 66709 253 66740 261
rect 66709 245 66743 253
rect 66544 213 66548 233
rect 66740 229 66743 245
rect 66607 228 66641 229
rect 66586 221 66641 228
rect 66709 221 66743 229
rect 66756 212 66758 262
rect 66796 253 66827 261
rect 66830 253 66832 262
rect 67019 261 67031 267
rect 66796 245 66832 253
rect 66895 253 66929 261
rect 66895 246 66950 253
rect 66895 245 66929 246
rect 66827 229 66832 245
rect 67021 233 67031 261
rect 67041 233 67061 267
rect 67244 261 67248 329
rect 67312 291 67316 341
rect 67312 251 67321 279
rect 67408 264 67418 291
rect 67367 262 67418 264
rect 67408 261 67419 262
rect 67375 253 67409 261
rect 67417 253 67419 261
rect 66796 221 66832 229
rect 66895 228 66929 229
rect 66895 221 66950 228
rect 66830 212 66832 221
rect 66476 103 66480 171
rect 66544 133 66548 183
rect 66598 159 66648 161
rect 66888 159 66938 161
rect 66648 143 66650 159
rect 66658 153 66674 159
rect 66676 153 66692 159
rect 66844 153 66860 159
rect 66862 153 66878 159
rect 66669 143 66692 152
rect 66844 143 66867 152
rect 66642 133 66650 143
rect 66648 109 66650 133
rect 66658 123 66659 143
rect 66669 118 66672 143
rect 66691 123 66692 143
rect 66701 133 66708 143
rect 66828 133 66835 143
rect 66844 123 66845 143
rect 66864 118 66867 143
rect 66877 123 66878 143
rect 66887 133 66894 143
rect 66658 109 66692 113
rect 66844 109 66878 113
rect 66938 109 66940 159
rect 66544 103 66586 104
rect 66950 103 66992 104
rect 66544 96 66548 103
rect 66439 62 66444 96
rect 66468 62 66473 96
rect 66511 79 66582 96
rect 66954 79 66988 96
rect 66991 79 67025 96
rect 66511 62 66586 79
rect 66544 61 66586 62
rect 66950 62 67025 79
rect 66950 61 66992 62
rect 66522 55 66608 61
rect 66928 55 67014 61
rect 67056 55 67060 233
rect 67244 183 67248 251
rect 67253 207 67263 241
rect 67273 213 67293 241
rect 67273 207 67287 213
rect 67312 207 67323 251
rect 67354 246 67430 253
rect 67463 251 67472 279
rect 67375 228 67409 246
rect 67417 228 67419 246
rect 67354 221 67430 228
rect 67417 213 67419 221
rect 67461 213 67472 251
rect 67536 241 67540 395
rect 67543 378 67548 412
rect 67572 378 67577 412
rect 67578 400 67589 412
rect 67792 395 67834 421
rect 68198 395 68240 421
rect 68455 420 68467 424
rect 68477 420 68489 424
rect 68527 420 68539 424
rect 68549 421 68561 424
rect 68719 421 68731 424
rect 68549 420 68602 421
rect 68560 412 68602 420
rect 68443 400 68454 412
rect 67724 341 67728 395
rect 67784 387 67830 395
rect 67784 383 67800 387
rect 67792 380 67800 383
rect 67826 380 67830 387
rect 67834 383 67842 395
rect 68190 383 68198 395
rect 68202 387 68236 395
rect 68202 380 68206 387
rect 68232 380 68236 387
rect 68240 383 68248 395
rect 67780 379 67846 380
rect 68186 379 68252 380
rect 67792 371 67796 379
rect 67846 365 67896 367
rect 68136 365 68186 367
rect 67886 361 67940 365
rect 68092 361 68146 365
rect 67886 356 67906 361
rect 68126 356 68146 361
rect 67896 341 67898 356
rect 67724 261 67728 329
rect 67792 305 67796 341
rect 67890 331 67898 341
rect 67906 331 67907 351
rect 67896 315 67898 331
rect 67917 322 67920 356
rect 67939 331 67940 351
rect 67949 331 67956 341
rect 68076 331 68083 341
rect 68092 331 68093 351
rect 68112 322 68115 356
rect 68125 331 68126 351
rect 68135 331 68142 341
rect 67906 315 67922 321
rect 67924 315 67940 321
rect 68092 315 68108 321
rect 68110 315 68126 321
rect 68186 315 68188 365
rect 67729 267 67765 295
rect 67729 261 67743 267
rect 67408 212 67419 213
rect 67253 183 67260 207
rect 67408 183 67418 212
rect 67499 207 67511 241
rect 67521 207 67541 241
rect 67244 103 67248 171
rect 67312 133 67316 183
rect 67312 98 67316 103
rect 67063 62 67068 96
rect 67092 62 67097 96
rect 67312 94 67350 98
rect 67312 79 67320 94
rect 67346 79 67350 94
rect 67434 94 67468 98
rect 67434 79 67438 94
rect 67464 79 67468 94
rect 67312 61 67354 79
rect 67430 61 67472 79
rect 67290 55 67376 61
rect 67408 55 67494 61
rect 67536 55 67540 207
rect 67566 183 67573 211
rect 67724 183 67728 251
rect 67733 233 67743 261
rect 67753 261 67767 267
rect 67792 261 67803 305
rect 68229 267 68240 305
rect 68267 267 68303 295
rect 68304 267 68308 395
rect 68455 378 68460 412
rect 68484 378 68489 412
rect 68490 400 68501 412
rect 68515 400 68526 412
rect 68527 395 68602 412
rect 68678 420 68731 421
rect 68741 420 68753 424
rect 68791 420 68803 424
rect 68813 420 68825 424
rect 68678 412 68720 420
rect 68678 395 68753 412
rect 68754 400 68765 412
rect 68779 400 68790 412
rect 68492 341 68496 395
rect 68527 378 68598 395
rect 68602 383 68610 395
rect 68670 383 68678 395
rect 68682 378 68716 395
rect 68719 378 68753 395
rect 68560 371 68564 378
rect 67954 262 68004 264
rect 68028 262 68078 264
rect 67753 233 67773 261
rect 67792 233 67801 261
rect 67855 253 67889 261
rect 67834 246 67889 253
rect 67855 245 67889 246
rect 67957 253 67988 261
rect 67957 245 67991 253
rect 67792 213 67796 233
rect 67988 229 67991 245
rect 67855 228 67889 229
rect 67834 221 67889 228
rect 67957 221 67991 229
rect 68004 212 68006 262
rect 68044 253 68075 261
rect 68078 253 68080 262
rect 68267 261 68279 267
rect 68044 245 68080 253
rect 68143 253 68177 261
rect 68143 246 68198 253
rect 68143 245 68177 246
rect 68075 229 68080 245
rect 68269 233 68279 261
rect 68289 233 68309 267
rect 68492 261 68496 329
rect 68560 291 68564 341
rect 68560 251 68569 279
rect 68656 264 68666 291
rect 68615 262 68666 264
rect 68656 261 68667 262
rect 68623 253 68657 261
rect 68665 253 68667 261
rect 68044 221 68080 229
rect 68143 228 68177 229
rect 68143 221 68198 228
rect 68078 212 68080 221
rect 67724 103 67728 171
rect 67792 133 67796 183
rect 67846 159 67896 161
rect 68136 159 68186 161
rect 67896 143 67898 159
rect 67906 153 67922 159
rect 67924 153 67940 159
rect 68092 153 68108 159
rect 68110 153 68126 159
rect 67917 143 67940 152
rect 68092 143 68115 152
rect 67890 133 67898 143
rect 67896 109 67898 133
rect 67906 123 67907 143
rect 67917 118 67920 143
rect 67939 123 67940 143
rect 67949 133 67956 143
rect 68076 133 68083 143
rect 68092 123 68093 143
rect 68112 118 68115 143
rect 68125 123 68126 143
rect 68135 133 68142 143
rect 67906 109 67940 113
rect 68092 109 68126 113
rect 68186 109 68188 159
rect 67792 103 67834 104
rect 68198 103 68240 104
rect 67792 96 67796 103
rect 67687 62 67692 96
rect 67716 62 67721 96
rect 67759 79 67830 96
rect 68202 79 68236 96
rect 68239 79 68273 96
rect 67759 62 67834 79
rect 67792 61 67834 62
rect 68198 62 68273 79
rect 68198 61 68240 62
rect 67770 55 67856 61
rect 68176 55 68262 61
rect 68304 55 68308 233
rect 68492 183 68496 251
rect 68501 207 68511 241
rect 68521 213 68541 241
rect 68521 207 68535 213
rect 68560 207 68571 251
rect 68602 246 68678 253
rect 68711 251 68720 279
rect 68623 228 68657 246
rect 68665 228 68667 246
rect 68602 221 68678 228
rect 68665 213 68667 221
rect 68709 213 68720 251
rect 68784 241 68788 395
rect 68791 378 68796 412
rect 68820 378 68825 412
rect 68826 400 68837 412
rect 69040 395 69082 421
rect 69446 395 69488 421
rect 69703 420 69715 424
rect 69725 420 69737 424
rect 69775 420 69787 424
rect 69797 421 69809 424
rect 69967 421 69979 424
rect 69797 420 69850 421
rect 69808 412 69850 420
rect 69691 400 69702 412
rect 68972 341 68976 395
rect 69032 387 69078 395
rect 69032 383 69048 387
rect 69040 380 69048 383
rect 69074 380 69078 387
rect 69082 383 69090 395
rect 69438 383 69446 395
rect 69450 387 69484 395
rect 69450 380 69454 387
rect 69480 380 69484 387
rect 69488 383 69496 395
rect 69028 379 69094 380
rect 69434 379 69500 380
rect 69040 371 69044 379
rect 69094 365 69144 367
rect 69384 365 69434 367
rect 69134 361 69188 365
rect 69340 361 69394 365
rect 69134 356 69154 361
rect 69374 356 69394 361
rect 69144 341 69146 356
rect 68972 261 68976 329
rect 69040 305 69044 341
rect 69138 331 69146 341
rect 69154 331 69155 351
rect 69144 315 69146 331
rect 69165 322 69168 356
rect 69187 331 69188 351
rect 69197 331 69204 341
rect 69324 331 69331 341
rect 69340 331 69341 351
rect 69360 322 69363 356
rect 69373 331 69374 351
rect 69383 331 69390 341
rect 69154 315 69170 321
rect 69172 315 69188 321
rect 69340 315 69356 321
rect 69358 315 69374 321
rect 69434 315 69436 365
rect 68977 267 69013 295
rect 68977 261 68991 267
rect 68656 212 68667 213
rect 68501 183 68508 207
rect 68656 183 68666 212
rect 68747 207 68759 241
rect 68769 207 68789 241
rect 68492 103 68496 171
rect 68560 133 68564 183
rect 68560 98 68564 103
rect 68311 62 68316 96
rect 68340 62 68345 96
rect 68560 94 68598 98
rect 68560 79 68568 94
rect 68594 79 68598 94
rect 68682 94 68716 98
rect 68682 79 68686 94
rect 68712 79 68716 94
rect 68560 61 68602 79
rect 68678 61 68720 79
rect 68538 55 68624 61
rect 68656 55 68742 61
rect 68784 55 68788 207
rect 68814 183 68821 211
rect 68972 183 68976 251
rect 68981 233 68991 261
rect 69001 261 69015 267
rect 69040 261 69051 305
rect 69477 267 69488 305
rect 69515 267 69551 295
rect 69552 267 69556 395
rect 69703 378 69708 412
rect 69732 378 69737 412
rect 69738 400 69749 412
rect 69763 400 69774 412
rect 69775 395 69850 412
rect 69926 420 69979 421
rect 69989 420 70001 424
rect 70039 420 70051 424
rect 70061 420 70073 424
rect 69926 412 69968 420
rect 69926 395 70001 412
rect 70002 400 70013 412
rect 70027 400 70038 412
rect 69740 341 69744 395
rect 69775 378 69846 395
rect 69850 383 69858 395
rect 69918 383 69926 395
rect 69930 378 69964 395
rect 69967 378 70001 395
rect 69808 371 69812 378
rect 69202 262 69252 264
rect 69276 262 69326 264
rect 69001 233 69021 261
rect 69040 233 69049 261
rect 69103 253 69137 261
rect 69082 246 69137 253
rect 69103 245 69137 246
rect 69205 253 69236 261
rect 69205 245 69239 253
rect 69040 213 69044 233
rect 69236 229 69239 245
rect 69103 228 69137 229
rect 69082 221 69137 228
rect 69205 221 69239 229
rect 69252 212 69254 262
rect 69292 253 69323 261
rect 69326 253 69328 262
rect 69515 261 69527 267
rect 69292 245 69328 253
rect 69391 253 69425 261
rect 69391 246 69446 253
rect 69391 245 69425 246
rect 69323 229 69328 245
rect 69517 233 69527 261
rect 69537 233 69557 267
rect 69740 261 69744 329
rect 69808 291 69812 341
rect 69808 251 69817 279
rect 69904 264 69914 291
rect 69863 262 69914 264
rect 69904 261 69915 262
rect 69871 253 69905 261
rect 69913 253 69915 261
rect 69292 221 69328 229
rect 69391 228 69425 229
rect 69391 221 69446 228
rect 69326 212 69328 221
rect 68972 103 68976 171
rect 69040 133 69044 183
rect 69094 159 69144 161
rect 69384 159 69434 161
rect 69144 143 69146 159
rect 69154 153 69170 159
rect 69172 153 69188 159
rect 69340 153 69356 159
rect 69358 153 69374 159
rect 69165 143 69188 152
rect 69340 143 69363 152
rect 69138 133 69146 143
rect 69144 109 69146 133
rect 69154 123 69155 143
rect 69165 118 69168 143
rect 69187 123 69188 143
rect 69197 133 69204 143
rect 69324 133 69331 143
rect 69340 123 69341 143
rect 69360 118 69363 143
rect 69373 123 69374 143
rect 69383 133 69390 143
rect 69154 109 69188 113
rect 69340 109 69374 113
rect 69434 109 69436 159
rect 69040 103 69082 104
rect 69446 103 69488 104
rect 69040 96 69044 103
rect 68935 62 68940 96
rect 68964 62 68969 96
rect 69007 79 69078 96
rect 69450 79 69484 96
rect 69487 79 69521 96
rect 69007 62 69082 79
rect 69040 61 69082 62
rect 69446 62 69521 79
rect 69446 61 69488 62
rect 69018 55 69104 61
rect 69424 55 69510 61
rect 69552 55 69556 233
rect 69740 183 69744 251
rect 69749 207 69759 241
rect 69769 213 69789 241
rect 69769 207 69783 213
rect 69808 207 69819 251
rect 69850 246 69926 253
rect 69959 251 69968 279
rect 69871 228 69905 246
rect 69913 228 69915 246
rect 69850 221 69926 228
rect 69913 213 69915 221
rect 69957 213 69968 251
rect 70032 241 70036 395
rect 70039 378 70044 412
rect 70068 378 70073 412
rect 70074 400 70085 412
rect 70288 395 70330 421
rect 70694 395 70736 421
rect 70951 420 70963 424
rect 70973 420 70985 424
rect 71023 420 71035 424
rect 71045 421 71057 424
rect 71215 421 71227 424
rect 71045 420 71098 421
rect 71056 412 71098 420
rect 70939 400 70950 412
rect 70220 341 70224 395
rect 70280 387 70326 395
rect 70280 383 70296 387
rect 70288 380 70296 383
rect 70322 380 70326 387
rect 70330 383 70338 395
rect 70686 383 70694 395
rect 70698 387 70732 395
rect 70698 380 70702 387
rect 70728 380 70732 387
rect 70736 383 70744 395
rect 70276 379 70342 380
rect 70682 379 70748 380
rect 70288 371 70292 379
rect 70342 365 70392 367
rect 70632 365 70682 367
rect 70382 361 70436 365
rect 70588 361 70642 365
rect 70382 356 70402 361
rect 70622 356 70642 361
rect 70392 341 70394 356
rect 70220 261 70224 329
rect 70288 305 70292 341
rect 70386 331 70394 341
rect 70402 331 70403 351
rect 70392 315 70394 331
rect 70413 322 70416 356
rect 70435 331 70436 351
rect 70445 331 70452 341
rect 70572 331 70579 341
rect 70588 331 70589 351
rect 70608 322 70611 356
rect 70621 331 70622 351
rect 70631 331 70638 341
rect 70402 315 70418 321
rect 70420 315 70436 321
rect 70588 315 70604 321
rect 70606 315 70622 321
rect 70682 315 70684 365
rect 70225 267 70261 295
rect 70225 261 70239 267
rect 69904 212 69915 213
rect 69749 183 69756 207
rect 69904 183 69914 212
rect 69995 207 70007 241
rect 70017 207 70037 241
rect 69740 103 69744 171
rect 69808 133 69812 183
rect 69808 98 69812 103
rect 69559 62 69564 96
rect 69588 62 69593 96
rect 69808 94 69846 98
rect 69808 79 69816 94
rect 69842 79 69846 94
rect 69930 94 69964 98
rect 69930 79 69934 94
rect 69960 79 69964 94
rect 69808 61 69850 79
rect 69926 61 69968 79
rect 69786 55 69872 61
rect 69904 55 69990 61
rect 70032 55 70036 207
rect 70062 183 70069 211
rect 70220 183 70224 251
rect 70229 233 70239 261
rect 70249 261 70263 267
rect 70288 261 70299 305
rect 70725 267 70736 305
rect 70763 267 70799 295
rect 70800 267 70804 395
rect 70951 378 70956 412
rect 70980 378 70985 412
rect 70986 400 70997 412
rect 71011 400 71022 412
rect 71023 395 71098 412
rect 71174 420 71227 421
rect 71237 420 71249 424
rect 71287 420 71299 424
rect 71309 420 71321 424
rect 71174 412 71216 420
rect 71174 395 71249 412
rect 71250 400 71261 412
rect 71275 400 71286 412
rect 70988 341 70992 395
rect 71023 378 71094 395
rect 71098 383 71106 395
rect 71166 383 71174 395
rect 71178 378 71212 395
rect 71215 378 71249 395
rect 71056 371 71060 378
rect 70450 262 70500 264
rect 70524 262 70574 264
rect 70249 233 70269 261
rect 70288 233 70297 261
rect 70351 253 70385 261
rect 70330 246 70385 253
rect 70351 245 70385 246
rect 70453 253 70484 261
rect 70453 245 70487 253
rect 70288 213 70292 233
rect 70484 229 70487 245
rect 70351 228 70385 229
rect 70330 221 70385 228
rect 70453 221 70487 229
rect 70500 212 70502 262
rect 70540 253 70571 261
rect 70574 253 70576 262
rect 70763 261 70775 267
rect 70540 245 70576 253
rect 70639 253 70673 261
rect 70639 246 70694 253
rect 70639 245 70673 246
rect 70571 229 70576 245
rect 70765 233 70775 261
rect 70785 233 70805 267
rect 70988 261 70992 329
rect 71056 291 71060 341
rect 71056 251 71065 279
rect 71152 264 71162 291
rect 71111 262 71162 264
rect 71152 261 71163 262
rect 71119 253 71153 261
rect 71161 253 71163 261
rect 70540 221 70576 229
rect 70639 228 70673 229
rect 70639 221 70694 228
rect 70574 212 70576 221
rect 70220 103 70224 171
rect 70288 133 70292 183
rect 70342 159 70392 161
rect 70632 159 70682 161
rect 70392 143 70394 159
rect 70402 153 70418 159
rect 70420 153 70436 159
rect 70588 153 70604 159
rect 70606 153 70622 159
rect 70413 143 70436 152
rect 70588 143 70611 152
rect 70386 133 70394 143
rect 70392 109 70394 133
rect 70402 123 70403 143
rect 70413 118 70416 143
rect 70435 123 70436 143
rect 70445 133 70452 143
rect 70572 133 70579 143
rect 70588 123 70589 143
rect 70608 118 70611 143
rect 70621 123 70622 143
rect 70631 133 70638 143
rect 70402 109 70436 113
rect 70588 109 70622 113
rect 70682 109 70684 159
rect 70288 103 70330 104
rect 70694 103 70736 104
rect 70288 96 70292 103
rect 70183 62 70188 96
rect 70212 62 70217 96
rect 70255 79 70326 96
rect 70698 79 70732 96
rect 70735 79 70769 96
rect 70255 62 70330 79
rect 70288 61 70330 62
rect 70694 62 70769 79
rect 70694 61 70736 62
rect 70266 55 70352 61
rect 70672 55 70758 61
rect 70800 55 70804 233
rect 70988 183 70992 251
rect 70997 207 71007 241
rect 71017 213 71037 241
rect 71017 207 71031 213
rect 71056 207 71067 251
rect 71098 246 71174 253
rect 71207 251 71216 279
rect 71119 228 71153 246
rect 71161 228 71163 246
rect 71098 221 71174 228
rect 71161 213 71163 221
rect 71205 213 71216 251
rect 71280 241 71284 395
rect 71287 378 71292 412
rect 71316 378 71321 412
rect 71322 400 71333 412
rect 71536 395 71578 421
rect 71942 395 71984 421
rect 72199 420 72211 424
rect 72221 420 72233 424
rect 72271 420 72283 424
rect 72293 421 72305 424
rect 72463 421 72475 424
rect 72293 420 72346 421
rect 72304 412 72346 420
rect 72187 400 72198 412
rect 71468 341 71472 395
rect 71528 387 71574 395
rect 71528 383 71544 387
rect 71536 380 71544 383
rect 71570 380 71574 387
rect 71578 383 71586 395
rect 71934 383 71942 395
rect 71946 387 71980 395
rect 71946 380 71950 387
rect 71976 380 71980 387
rect 71984 383 71992 395
rect 71524 379 71590 380
rect 71930 379 71996 380
rect 71536 371 71540 379
rect 71590 365 71640 367
rect 71880 365 71930 367
rect 71630 361 71684 365
rect 71836 361 71890 365
rect 71630 356 71650 361
rect 71870 356 71890 361
rect 71640 341 71642 356
rect 71468 261 71472 329
rect 71536 305 71540 341
rect 71634 331 71642 341
rect 71650 331 71651 351
rect 71640 315 71642 331
rect 71661 322 71664 356
rect 71683 331 71684 351
rect 71693 331 71700 341
rect 71820 331 71827 341
rect 71836 331 71837 351
rect 71856 322 71859 356
rect 71869 331 71870 351
rect 71879 331 71886 341
rect 71650 315 71666 321
rect 71668 315 71684 321
rect 71836 315 71852 321
rect 71854 315 71870 321
rect 71930 315 71932 365
rect 71473 267 71509 295
rect 71473 261 71487 267
rect 71152 212 71163 213
rect 70997 183 71004 207
rect 71152 183 71162 212
rect 71243 207 71255 241
rect 71265 207 71285 241
rect 70988 103 70992 171
rect 71056 133 71060 183
rect 71056 98 71060 103
rect 70807 62 70812 96
rect 70836 62 70841 96
rect 71056 94 71094 98
rect 71056 79 71064 94
rect 71090 79 71094 94
rect 71178 94 71212 98
rect 71178 79 71182 94
rect 71208 79 71212 94
rect 71056 61 71098 79
rect 71174 61 71216 79
rect 71034 55 71120 61
rect 71152 55 71238 61
rect 71280 55 71284 207
rect 71310 183 71317 211
rect 71468 183 71472 251
rect 71477 233 71487 261
rect 71497 261 71511 267
rect 71536 261 71547 305
rect 71973 267 71984 305
rect 72011 267 72047 295
rect 72048 267 72052 395
rect 72199 378 72204 412
rect 72228 378 72233 412
rect 72234 400 72245 412
rect 72259 400 72270 412
rect 72271 395 72346 412
rect 72422 420 72475 421
rect 72485 420 72497 424
rect 72535 420 72547 424
rect 72557 420 72569 424
rect 72422 412 72464 420
rect 72422 395 72497 412
rect 72498 400 72509 412
rect 72523 400 72534 412
rect 72236 341 72240 395
rect 72271 378 72342 395
rect 72346 383 72354 395
rect 72414 383 72422 395
rect 72426 378 72460 395
rect 72463 378 72497 395
rect 72304 371 72308 378
rect 71698 262 71748 264
rect 71772 262 71822 264
rect 71497 233 71517 261
rect 71536 233 71545 261
rect 71599 253 71633 261
rect 71578 246 71633 253
rect 71599 245 71633 246
rect 71701 253 71732 261
rect 71701 245 71735 253
rect 71536 213 71540 233
rect 71732 229 71735 245
rect 71599 228 71633 229
rect 71578 221 71633 228
rect 71701 221 71735 229
rect 71748 212 71750 262
rect 71788 253 71819 261
rect 71822 253 71824 262
rect 72011 261 72023 267
rect 71788 245 71824 253
rect 71887 253 71921 261
rect 71887 246 71942 253
rect 71887 245 71921 246
rect 71819 229 71824 245
rect 72013 233 72023 261
rect 72033 233 72053 267
rect 72236 261 72240 329
rect 72304 291 72308 341
rect 72304 251 72313 279
rect 72400 264 72410 291
rect 72359 262 72410 264
rect 72400 261 72411 262
rect 72367 253 72401 261
rect 72409 253 72411 261
rect 71788 221 71824 229
rect 71887 228 71921 229
rect 71887 221 71942 228
rect 71822 212 71824 221
rect 71468 103 71472 171
rect 71536 133 71540 183
rect 71590 159 71640 161
rect 71880 159 71930 161
rect 71640 143 71642 159
rect 71650 153 71666 159
rect 71668 153 71684 159
rect 71836 153 71852 159
rect 71854 153 71870 159
rect 71661 143 71684 152
rect 71836 143 71859 152
rect 71634 133 71642 143
rect 71640 109 71642 133
rect 71650 123 71651 143
rect 71661 118 71664 143
rect 71683 123 71684 143
rect 71693 133 71700 143
rect 71820 133 71827 143
rect 71836 123 71837 143
rect 71856 118 71859 143
rect 71869 123 71870 143
rect 71879 133 71886 143
rect 71650 109 71684 113
rect 71836 109 71870 113
rect 71930 109 71932 159
rect 71536 103 71578 104
rect 71942 103 71984 104
rect 71536 96 71540 103
rect 71431 62 71436 96
rect 71460 62 71465 96
rect 71503 79 71574 96
rect 71946 79 71980 96
rect 71983 79 72017 96
rect 71503 62 71578 79
rect 71536 61 71578 62
rect 71942 62 72017 79
rect 71942 61 71984 62
rect 71514 55 71600 61
rect 71920 55 72006 61
rect 72048 55 72052 233
rect 72236 183 72240 251
rect 72245 207 72255 241
rect 72265 213 72285 241
rect 72265 207 72279 213
rect 72304 207 72315 251
rect 72346 246 72422 253
rect 72455 251 72464 279
rect 72367 228 72401 246
rect 72409 228 72411 246
rect 72346 221 72422 228
rect 72409 213 72411 221
rect 72453 213 72464 251
rect 72528 241 72532 395
rect 72535 378 72540 412
rect 72564 378 72569 412
rect 72570 400 72581 412
rect 72784 395 72826 421
rect 73190 395 73232 421
rect 73447 420 73459 424
rect 73469 420 73481 424
rect 73519 420 73531 424
rect 73541 421 73553 424
rect 73711 421 73723 424
rect 73541 420 73594 421
rect 73552 412 73594 420
rect 73435 400 73446 412
rect 72716 341 72720 395
rect 72776 387 72822 395
rect 72776 383 72792 387
rect 72784 380 72792 383
rect 72818 380 72822 387
rect 72826 383 72834 395
rect 73182 383 73190 395
rect 73194 387 73228 395
rect 73194 380 73198 387
rect 73224 380 73228 387
rect 73232 383 73240 395
rect 72772 379 72838 380
rect 73178 379 73244 380
rect 72784 371 72788 379
rect 72838 365 72888 367
rect 73128 365 73178 367
rect 72878 361 72932 365
rect 73084 361 73138 365
rect 72878 356 72898 361
rect 73118 356 73138 361
rect 72888 341 72890 356
rect 72716 261 72720 329
rect 72784 305 72788 341
rect 72882 331 72890 341
rect 72898 331 72899 351
rect 72888 315 72890 331
rect 72909 322 72912 356
rect 72931 331 72932 351
rect 72941 331 72948 341
rect 73068 331 73075 341
rect 73084 331 73085 351
rect 73104 322 73107 356
rect 73117 331 73118 351
rect 73127 331 73134 341
rect 72898 315 72914 321
rect 72916 315 72932 321
rect 73084 315 73100 321
rect 73102 315 73118 321
rect 73178 315 73180 365
rect 72721 267 72757 295
rect 72721 261 72735 267
rect 72400 212 72411 213
rect 72245 183 72252 207
rect 72400 183 72410 212
rect 72491 207 72503 241
rect 72513 207 72533 241
rect 72236 103 72240 171
rect 72304 133 72308 183
rect 72304 98 72308 103
rect 72055 62 72060 96
rect 72084 62 72089 96
rect 72304 94 72342 98
rect 72304 79 72312 94
rect 72338 79 72342 94
rect 72426 94 72460 98
rect 72426 79 72430 94
rect 72456 79 72460 94
rect 72304 61 72346 79
rect 72422 61 72464 79
rect 72282 55 72368 61
rect 72400 55 72486 61
rect 72528 55 72532 207
rect 72558 183 72565 211
rect 72716 183 72720 251
rect 72725 233 72735 261
rect 72745 261 72759 267
rect 72784 261 72795 305
rect 73221 267 73232 305
rect 73259 267 73295 295
rect 73296 267 73300 395
rect 73447 378 73452 412
rect 73476 378 73481 412
rect 73482 400 73493 412
rect 73507 400 73518 412
rect 73519 395 73594 412
rect 73670 420 73723 421
rect 73733 420 73745 424
rect 73783 420 73795 424
rect 73805 420 73817 424
rect 73670 412 73712 420
rect 73670 395 73745 412
rect 73746 400 73757 412
rect 73771 400 73782 412
rect 73484 341 73488 395
rect 73519 378 73590 395
rect 73594 383 73602 395
rect 73662 383 73670 395
rect 73674 378 73708 395
rect 73711 378 73745 395
rect 73552 371 73556 378
rect 72946 262 72996 264
rect 73020 262 73070 264
rect 72745 233 72765 261
rect 72784 233 72793 261
rect 72847 253 72881 261
rect 72826 246 72881 253
rect 72847 245 72881 246
rect 72949 253 72980 261
rect 72949 245 72983 253
rect 72784 213 72788 233
rect 72980 229 72983 245
rect 72847 228 72881 229
rect 72826 221 72881 228
rect 72949 221 72983 229
rect 72996 212 72998 262
rect 73036 253 73067 261
rect 73070 253 73072 262
rect 73259 261 73271 267
rect 73036 245 73072 253
rect 73135 253 73169 261
rect 73135 246 73190 253
rect 73135 245 73169 246
rect 73067 229 73072 245
rect 73261 233 73271 261
rect 73281 233 73301 267
rect 73484 261 73488 329
rect 73552 291 73556 341
rect 73552 251 73561 279
rect 73648 264 73658 291
rect 73607 262 73658 264
rect 73648 261 73659 262
rect 73615 253 73649 261
rect 73657 253 73659 261
rect 73036 221 73072 229
rect 73135 228 73169 229
rect 73135 221 73190 228
rect 73070 212 73072 221
rect 72716 103 72720 171
rect 72784 133 72788 183
rect 72838 159 72888 161
rect 73128 159 73178 161
rect 72888 143 72890 159
rect 72898 153 72914 159
rect 72916 153 72932 159
rect 73084 153 73100 159
rect 73102 153 73118 159
rect 72909 143 72932 152
rect 73084 143 73107 152
rect 72882 133 72890 143
rect 72888 109 72890 133
rect 72898 123 72899 143
rect 72909 118 72912 143
rect 72931 123 72932 143
rect 72941 133 72948 143
rect 73068 133 73075 143
rect 73084 123 73085 143
rect 73104 118 73107 143
rect 73117 123 73118 143
rect 73127 133 73134 143
rect 72898 109 72932 113
rect 73084 109 73118 113
rect 73178 109 73180 159
rect 72784 103 72826 104
rect 73190 103 73232 104
rect 72784 96 72788 103
rect 72679 62 72684 96
rect 72708 62 72713 96
rect 72751 79 72822 96
rect 73194 79 73228 96
rect 73231 79 73265 96
rect 72751 62 72826 79
rect 72784 61 72826 62
rect 73190 62 73265 79
rect 73190 61 73232 62
rect 72762 55 72848 61
rect 73168 55 73254 61
rect 73296 55 73300 233
rect 73484 183 73488 251
rect 73493 207 73503 241
rect 73513 213 73533 241
rect 73513 207 73527 213
rect 73552 207 73563 251
rect 73594 246 73670 253
rect 73703 251 73712 279
rect 73615 228 73649 246
rect 73657 228 73659 246
rect 73594 221 73670 228
rect 73657 213 73659 221
rect 73701 213 73712 251
rect 73776 241 73780 395
rect 73783 378 73788 412
rect 73812 378 73817 412
rect 73818 400 73829 412
rect 74032 395 74074 421
rect 74438 395 74480 421
rect 74695 420 74707 424
rect 74717 420 74729 424
rect 74767 420 74779 424
rect 74789 421 74801 424
rect 74959 421 74971 424
rect 74789 420 74842 421
rect 74800 412 74842 420
rect 74683 400 74694 412
rect 73964 341 73968 395
rect 74024 387 74070 395
rect 74024 383 74040 387
rect 74032 380 74040 383
rect 74066 380 74070 387
rect 74074 383 74082 395
rect 74430 383 74438 395
rect 74442 387 74476 395
rect 74442 380 74446 387
rect 74472 380 74476 387
rect 74480 383 74488 395
rect 74020 379 74086 380
rect 74426 379 74492 380
rect 74032 371 74036 379
rect 74086 365 74136 367
rect 74376 365 74426 367
rect 74126 361 74180 365
rect 74332 361 74386 365
rect 74126 356 74146 361
rect 74366 356 74386 361
rect 74136 341 74138 356
rect 73964 261 73968 329
rect 74032 305 74036 341
rect 74130 331 74138 341
rect 74146 331 74147 351
rect 74136 315 74138 331
rect 74157 322 74160 356
rect 74179 331 74180 351
rect 74189 331 74196 341
rect 74316 331 74323 341
rect 74332 331 74333 351
rect 74352 322 74355 356
rect 74365 331 74366 351
rect 74375 331 74382 341
rect 74146 315 74162 321
rect 74164 315 74180 321
rect 74332 315 74348 321
rect 74350 315 74366 321
rect 74426 315 74428 365
rect 73969 267 74005 295
rect 73969 261 73983 267
rect 73648 212 73659 213
rect 73493 183 73500 207
rect 73648 183 73658 212
rect 73739 207 73751 241
rect 73761 207 73781 241
rect 73484 103 73488 171
rect 73552 133 73556 183
rect 73552 98 73556 103
rect 73303 62 73308 96
rect 73332 62 73337 96
rect 73552 94 73590 98
rect 73552 79 73560 94
rect 73586 79 73590 94
rect 73674 94 73708 98
rect 73674 79 73678 94
rect 73704 79 73708 94
rect 73552 61 73594 79
rect 73670 61 73712 79
rect 73530 55 73616 61
rect 73648 55 73734 61
rect 73776 55 73780 207
rect 73806 183 73813 211
rect 73964 183 73968 251
rect 73973 233 73983 261
rect 73993 261 74007 267
rect 74032 261 74043 305
rect 74469 267 74480 305
rect 74507 267 74543 295
rect 74544 267 74548 395
rect 74695 378 74700 412
rect 74724 378 74729 412
rect 74730 400 74741 412
rect 74755 400 74766 412
rect 74767 395 74842 412
rect 74918 420 74971 421
rect 74981 420 74993 424
rect 75031 420 75043 424
rect 75053 420 75065 424
rect 74918 412 74960 420
rect 74918 395 74993 412
rect 74994 400 75005 412
rect 75019 400 75030 412
rect 74732 341 74736 395
rect 74767 378 74838 395
rect 74842 383 74850 395
rect 74910 383 74918 395
rect 74922 378 74956 395
rect 74959 378 74993 395
rect 74800 371 74804 378
rect 74194 262 74244 264
rect 74268 262 74318 264
rect 73993 233 74013 261
rect 74032 233 74041 261
rect 74095 253 74129 261
rect 74074 246 74129 253
rect 74095 245 74129 246
rect 74197 253 74228 261
rect 74197 245 74231 253
rect 74032 213 74036 233
rect 74228 229 74231 245
rect 74095 228 74129 229
rect 74074 221 74129 228
rect 74197 221 74231 229
rect 74244 212 74246 262
rect 74284 253 74315 261
rect 74318 253 74320 262
rect 74507 261 74519 267
rect 74284 245 74320 253
rect 74383 253 74417 261
rect 74383 246 74438 253
rect 74383 245 74417 246
rect 74315 229 74320 245
rect 74509 233 74519 261
rect 74529 233 74549 267
rect 74732 261 74736 329
rect 74800 291 74804 341
rect 74800 251 74809 279
rect 74896 264 74906 291
rect 74855 262 74906 264
rect 74896 261 74907 262
rect 74863 253 74897 261
rect 74905 253 74907 261
rect 74284 221 74320 229
rect 74383 228 74417 229
rect 74383 221 74438 228
rect 74318 212 74320 221
rect 73964 103 73968 171
rect 74032 133 74036 183
rect 74086 159 74136 161
rect 74376 159 74426 161
rect 74136 143 74138 159
rect 74146 153 74162 159
rect 74164 153 74180 159
rect 74332 153 74348 159
rect 74350 153 74366 159
rect 74157 143 74180 152
rect 74332 143 74355 152
rect 74130 133 74138 143
rect 74136 109 74138 133
rect 74146 123 74147 143
rect 74157 118 74160 143
rect 74179 123 74180 143
rect 74189 133 74196 143
rect 74316 133 74323 143
rect 74332 123 74333 143
rect 74352 118 74355 143
rect 74365 123 74366 143
rect 74375 133 74382 143
rect 74146 109 74180 113
rect 74332 109 74366 113
rect 74426 109 74428 159
rect 74032 103 74074 104
rect 74438 103 74480 104
rect 74032 96 74036 103
rect 73927 62 73932 96
rect 73956 62 73961 96
rect 73999 79 74070 96
rect 74442 79 74476 96
rect 74479 79 74513 96
rect 73999 62 74074 79
rect 74032 61 74074 62
rect 74438 62 74513 79
rect 74438 61 74480 62
rect 74010 55 74096 61
rect 74416 55 74502 61
rect 74544 55 74548 233
rect 74732 183 74736 251
rect 74741 207 74751 241
rect 74761 213 74781 241
rect 74761 207 74775 213
rect 74800 207 74811 251
rect 74842 246 74918 253
rect 74951 251 74960 279
rect 74863 228 74897 246
rect 74905 228 74907 246
rect 74842 221 74918 228
rect 74905 213 74907 221
rect 74949 213 74960 251
rect 75024 241 75028 395
rect 75031 378 75036 412
rect 75060 378 75065 412
rect 75066 400 75077 412
rect 75280 395 75322 421
rect 75686 395 75728 421
rect 75943 420 75955 424
rect 75965 420 75977 424
rect 76015 420 76027 424
rect 76037 421 76049 424
rect 76207 421 76219 424
rect 76037 420 76090 421
rect 76048 412 76090 420
rect 75931 400 75942 412
rect 75212 341 75216 395
rect 75272 387 75318 395
rect 75272 383 75288 387
rect 75280 380 75288 383
rect 75314 380 75318 387
rect 75322 383 75330 395
rect 75678 383 75686 395
rect 75690 387 75724 395
rect 75690 380 75694 387
rect 75720 380 75724 387
rect 75728 383 75736 395
rect 75268 379 75334 380
rect 75674 379 75740 380
rect 75280 371 75284 379
rect 75334 365 75384 367
rect 75624 365 75674 367
rect 75374 361 75428 365
rect 75580 361 75634 365
rect 75374 356 75394 361
rect 75614 356 75634 361
rect 75384 341 75386 356
rect 75212 261 75216 329
rect 75280 305 75284 341
rect 75378 331 75386 341
rect 75394 331 75395 351
rect 75384 315 75386 331
rect 75405 322 75408 356
rect 75427 331 75428 351
rect 75437 331 75444 341
rect 75564 331 75571 341
rect 75580 331 75581 351
rect 75600 322 75603 356
rect 75613 331 75614 351
rect 75623 331 75630 341
rect 75394 315 75410 321
rect 75412 315 75428 321
rect 75580 315 75596 321
rect 75598 315 75614 321
rect 75674 315 75676 365
rect 75217 267 75253 295
rect 75217 261 75231 267
rect 74896 212 74907 213
rect 74741 183 74748 207
rect 74896 183 74906 212
rect 74987 207 74999 241
rect 75009 207 75029 241
rect 74732 103 74736 171
rect 74800 133 74804 183
rect 74800 98 74804 103
rect 74551 62 74556 96
rect 74580 62 74585 96
rect 74800 94 74838 98
rect 74800 79 74808 94
rect 74834 79 74838 94
rect 74922 94 74956 98
rect 74922 79 74926 94
rect 74952 79 74956 94
rect 74800 61 74842 79
rect 74918 61 74960 79
rect 74778 55 74864 61
rect 74896 55 74982 61
rect 75024 55 75028 207
rect 75054 183 75061 211
rect 75212 183 75216 251
rect 75221 233 75231 261
rect 75241 261 75255 267
rect 75280 261 75291 305
rect 75717 267 75728 305
rect 75755 267 75791 295
rect 75792 267 75796 395
rect 75943 378 75948 412
rect 75972 378 75977 412
rect 75978 400 75989 412
rect 76003 400 76014 412
rect 76015 395 76090 412
rect 76166 420 76219 421
rect 76229 420 76241 424
rect 76279 420 76291 424
rect 76301 420 76313 424
rect 76166 412 76208 420
rect 76166 395 76241 412
rect 76242 400 76253 412
rect 76267 400 76278 412
rect 75980 341 75984 395
rect 76015 378 76086 395
rect 76090 383 76098 395
rect 76158 383 76166 395
rect 76170 378 76204 395
rect 76207 378 76241 395
rect 76048 371 76052 378
rect 75442 262 75492 264
rect 75516 262 75566 264
rect 75241 233 75261 261
rect 75280 233 75289 261
rect 75343 253 75377 261
rect 75322 246 75377 253
rect 75343 245 75377 246
rect 75445 253 75476 261
rect 75445 245 75479 253
rect 75280 213 75284 233
rect 75476 229 75479 245
rect 75343 228 75377 229
rect 75322 221 75377 228
rect 75445 221 75479 229
rect 75492 212 75494 262
rect 75532 253 75563 261
rect 75566 253 75568 262
rect 75755 261 75767 267
rect 75532 245 75568 253
rect 75631 253 75665 261
rect 75631 246 75686 253
rect 75631 245 75665 246
rect 75563 229 75568 245
rect 75757 233 75767 261
rect 75777 233 75797 267
rect 75980 261 75984 329
rect 76048 291 76052 341
rect 76048 251 76057 279
rect 76144 264 76154 291
rect 76103 262 76154 264
rect 76144 261 76155 262
rect 76111 253 76145 261
rect 76153 253 76155 261
rect 75532 221 75568 229
rect 75631 228 75665 229
rect 75631 221 75686 228
rect 75566 212 75568 221
rect 75212 103 75216 171
rect 75280 133 75284 183
rect 75334 159 75384 161
rect 75624 159 75674 161
rect 75384 143 75386 159
rect 75394 153 75410 159
rect 75412 153 75428 159
rect 75580 153 75596 159
rect 75598 153 75614 159
rect 75405 143 75428 152
rect 75580 143 75603 152
rect 75378 133 75386 143
rect 75384 109 75386 133
rect 75394 123 75395 143
rect 75405 118 75408 143
rect 75427 123 75428 143
rect 75437 133 75444 143
rect 75564 133 75571 143
rect 75580 123 75581 143
rect 75600 118 75603 143
rect 75613 123 75614 143
rect 75623 133 75630 143
rect 75394 109 75428 113
rect 75580 109 75614 113
rect 75674 109 75676 159
rect 75280 103 75322 104
rect 75686 103 75728 104
rect 75280 96 75284 103
rect 75175 62 75180 96
rect 75204 62 75209 96
rect 75247 79 75318 96
rect 75690 79 75724 96
rect 75727 79 75761 96
rect 75247 62 75322 79
rect 75280 61 75322 62
rect 75686 62 75761 79
rect 75686 61 75728 62
rect 75258 55 75344 61
rect 75664 55 75750 61
rect 75792 55 75796 233
rect 75980 183 75984 251
rect 75989 207 75999 241
rect 76009 213 76029 241
rect 76009 207 76023 213
rect 76048 207 76059 251
rect 76090 246 76166 253
rect 76199 251 76208 279
rect 76111 228 76145 246
rect 76153 228 76155 246
rect 76090 221 76166 228
rect 76153 213 76155 221
rect 76197 213 76208 251
rect 76272 241 76276 395
rect 76279 378 76284 412
rect 76308 378 76313 412
rect 76314 400 76325 412
rect 76528 395 76570 421
rect 76934 395 76976 421
rect 77191 420 77203 424
rect 77213 420 77225 424
rect 77263 420 77275 424
rect 77285 421 77297 424
rect 77455 421 77467 424
rect 77285 420 77338 421
rect 77296 412 77338 420
rect 77179 400 77190 412
rect 76460 341 76464 395
rect 76520 387 76566 395
rect 76520 383 76536 387
rect 76528 380 76536 383
rect 76562 380 76566 387
rect 76570 383 76578 395
rect 76926 383 76934 395
rect 76938 387 76972 395
rect 76938 380 76942 387
rect 76968 380 76972 387
rect 76976 383 76984 395
rect 76516 379 76582 380
rect 76922 379 76988 380
rect 76528 371 76532 379
rect 76582 365 76632 367
rect 76872 365 76922 367
rect 76622 361 76676 365
rect 76828 361 76882 365
rect 76622 356 76642 361
rect 76862 356 76882 361
rect 76632 341 76634 356
rect 76460 261 76464 329
rect 76528 305 76532 341
rect 76626 331 76634 341
rect 76642 331 76643 351
rect 76632 315 76634 331
rect 76653 322 76656 356
rect 76675 331 76676 351
rect 76685 331 76692 341
rect 76812 331 76819 341
rect 76828 331 76829 351
rect 76848 322 76851 356
rect 76861 331 76862 351
rect 76871 331 76878 341
rect 76642 315 76658 321
rect 76660 315 76676 321
rect 76828 315 76844 321
rect 76846 315 76862 321
rect 76922 315 76924 365
rect 76465 267 76501 295
rect 76465 261 76479 267
rect 76144 212 76155 213
rect 75989 183 75996 207
rect 76144 183 76154 212
rect 76235 207 76247 241
rect 76257 207 76277 241
rect 75980 103 75984 171
rect 76048 133 76052 183
rect 76048 98 76052 103
rect 75799 62 75804 96
rect 75828 62 75833 96
rect 76048 94 76086 98
rect 76048 79 76056 94
rect 76082 79 76086 94
rect 76170 94 76204 98
rect 76170 79 76174 94
rect 76200 79 76204 94
rect 76048 61 76090 79
rect 76166 61 76208 79
rect 76026 55 76112 61
rect 76144 55 76230 61
rect 76272 55 76276 207
rect 76302 183 76309 211
rect 76460 183 76464 251
rect 76469 233 76479 261
rect 76489 261 76503 267
rect 76528 261 76539 305
rect 76965 267 76976 305
rect 77003 267 77039 295
rect 77040 267 77044 395
rect 77191 378 77196 412
rect 77220 378 77225 412
rect 77226 400 77237 412
rect 77251 400 77262 412
rect 77263 395 77338 412
rect 77414 420 77467 421
rect 77477 420 77489 424
rect 77527 420 77539 424
rect 77549 420 77561 424
rect 77414 412 77456 420
rect 77414 395 77489 412
rect 77490 400 77501 412
rect 77515 400 77526 412
rect 77228 341 77232 395
rect 77263 378 77334 395
rect 77338 383 77346 395
rect 77406 383 77414 395
rect 77418 378 77452 395
rect 77455 378 77489 395
rect 77296 371 77300 378
rect 76690 262 76740 264
rect 76764 262 76814 264
rect 76489 233 76509 261
rect 76528 233 76537 261
rect 76591 253 76625 261
rect 76570 246 76625 253
rect 76591 245 76625 246
rect 76693 253 76724 261
rect 76693 245 76727 253
rect 76528 213 76532 233
rect 76724 229 76727 245
rect 76591 228 76625 229
rect 76570 221 76625 228
rect 76693 221 76727 229
rect 76740 212 76742 262
rect 76780 253 76811 261
rect 76814 253 76816 262
rect 77003 261 77015 267
rect 76780 245 76816 253
rect 76879 253 76913 261
rect 76879 246 76934 253
rect 76879 245 76913 246
rect 76811 229 76816 245
rect 77005 233 77015 261
rect 77025 233 77045 267
rect 77228 261 77232 329
rect 77296 291 77300 341
rect 77296 251 77305 279
rect 77392 264 77402 291
rect 77351 262 77402 264
rect 77392 261 77403 262
rect 77359 253 77393 261
rect 77401 253 77403 261
rect 76780 221 76816 229
rect 76879 228 76913 229
rect 76879 221 76934 228
rect 76814 212 76816 221
rect 76460 103 76464 171
rect 76528 133 76532 183
rect 76582 159 76632 161
rect 76872 159 76922 161
rect 76632 143 76634 159
rect 76642 153 76658 159
rect 76660 153 76676 159
rect 76828 153 76844 159
rect 76846 153 76862 159
rect 76653 143 76676 152
rect 76828 143 76851 152
rect 76626 133 76634 143
rect 76632 109 76634 133
rect 76642 123 76643 143
rect 76653 118 76656 143
rect 76675 123 76676 143
rect 76685 133 76692 143
rect 76812 133 76819 143
rect 76828 123 76829 143
rect 76848 118 76851 143
rect 76861 123 76862 143
rect 76871 133 76878 143
rect 76642 109 76676 113
rect 76828 109 76862 113
rect 76922 109 76924 159
rect 76528 103 76570 104
rect 76934 103 76976 104
rect 76528 96 76532 103
rect 76423 62 76428 96
rect 76452 62 76457 96
rect 76495 79 76566 96
rect 76938 79 76972 96
rect 76975 79 77009 96
rect 76495 62 76570 79
rect 76528 61 76570 62
rect 76934 62 77009 79
rect 76934 61 76976 62
rect 76506 55 76592 61
rect 76912 55 76998 61
rect 77040 55 77044 233
rect 77228 183 77232 251
rect 77237 207 77247 241
rect 77257 213 77277 241
rect 77257 207 77271 213
rect 77296 207 77307 251
rect 77338 246 77414 253
rect 77447 251 77456 279
rect 77359 228 77393 246
rect 77401 228 77403 246
rect 77338 221 77414 228
rect 77401 213 77403 221
rect 77445 213 77456 251
rect 77520 241 77524 395
rect 77527 378 77532 412
rect 77556 378 77561 412
rect 77562 400 77573 412
rect 77776 395 77818 421
rect 78182 395 78224 421
rect 78439 420 78451 424
rect 78461 420 78473 424
rect 78511 420 78523 424
rect 78533 421 78545 424
rect 78703 421 78715 424
rect 78533 420 78586 421
rect 78544 412 78586 420
rect 78427 400 78438 412
rect 77708 341 77712 395
rect 77768 387 77814 395
rect 77768 383 77784 387
rect 77776 380 77784 383
rect 77810 380 77814 387
rect 77818 383 77826 395
rect 78174 383 78182 395
rect 78186 387 78220 395
rect 78186 380 78190 387
rect 78216 380 78220 387
rect 78224 383 78232 395
rect 77764 379 77830 380
rect 78170 379 78236 380
rect 77776 371 77780 379
rect 77830 365 77880 367
rect 78120 365 78170 367
rect 77870 361 77924 365
rect 78076 361 78130 365
rect 77870 356 77890 361
rect 78110 356 78130 361
rect 77880 341 77882 356
rect 77708 261 77712 329
rect 77776 305 77780 341
rect 77874 331 77882 341
rect 77890 331 77891 351
rect 77880 315 77882 331
rect 77901 322 77904 356
rect 77923 331 77924 351
rect 77933 331 77940 341
rect 78060 331 78067 341
rect 78076 331 78077 351
rect 78096 322 78099 356
rect 78109 331 78110 351
rect 78119 331 78126 341
rect 77890 315 77906 321
rect 77908 315 77924 321
rect 78076 315 78092 321
rect 78094 315 78110 321
rect 78170 315 78172 365
rect 77713 267 77749 295
rect 77713 261 77727 267
rect 77392 212 77403 213
rect 77237 183 77244 207
rect 77392 183 77402 212
rect 77483 207 77495 241
rect 77505 207 77525 241
rect 77228 103 77232 171
rect 77296 133 77300 183
rect 77296 98 77300 103
rect 77047 62 77052 96
rect 77076 62 77081 96
rect 77296 94 77334 98
rect 77296 79 77304 94
rect 77330 79 77334 94
rect 77418 94 77452 98
rect 77418 79 77422 94
rect 77448 79 77452 94
rect 77296 61 77338 79
rect 77414 61 77456 79
rect 77274 55 77360 61
rect 77392 55 77478 61
rect 77520 55 77524 207
rect 77550 183 77557 211
rect 77708 183 77712 251
rect 77717 233 77727 261
rect 77737 261 77751 267
rect 77776 261 77787 305
rect 78213 267 78224 305
rect 78251 267 78287 295
rect 78288 267 78292 395
rect 78439 378 78444 412
rect 78468 378 78473 412
rect 78474 400 78485 412
rect 78499 400 78510 412
rect 78511 395 78586 412
rect 78662 420 78715 421
rect 78725 420 78737 424
rect 78775 420 78787 424
rect 78797 420 78809 424
rect 78662 412 78704 420
rect 78662 395 78737 412
rect 78738 400 78749 412
rect 78763 400 78774 412
rect 78476 341 78480 395
rect 78511 378 78582 395
rect 78586 383 78594 395
rect 78654 383 78662 395
rect 78666 378 78700 395
rect 78703 378 78737 395
rect 78544 371 78548 378
rect 77938 262 77988 264
rect 78012 262 78062 264
rect 77737 233 77757 261
rect 77776 233 77785 261
rect 77839 253 77873 261
rect 77818 246 77873 253
rect 77839 245 77873 246
rect 77941 253 77972 261
rect 77941 245 77975 253
rect 77776 213 77780 233
rect 77972 229 77975 245
rect 77839 228 77873 229
rect 77818 221 77873 228
rect 77941 221 77975 229
rect 77988 212 77990 262
rect 78028 253 78059 261
rect 78062 253 78064 262
rect 78251 261 78263 267
rect 78028 245 78064 253
rect 78127 253 78161 261
rect 78127 246 78182 253
rect 78127 245 78161 246
rect 78059 229 78064 245
rect 78253 233 78263 261
rect 78273 233 78293 267
rect 78476 261 78480 329
rect 78544 291 78548 341
rect 78544 251 78553 279
rect 78640 264 78650 291
rect 78599 262 78650 264
rect 78640 261 78651 262
rect 78607 253 78641 261
rect 78649 253 78651 261
rect 78028 221 78064 229
rect 78127 228 78161 229
rect 78127 221 78182 228
rect 78062 212 78064 221
rect 77708 103 77712 171
rect 77776 133 77780 183
rect 77830 159 77880 161
rect 78120 159 78170 161
rect 77880 143 77882 159
rect 77890 153 77906 159
rect 77908 153 77924 159
rect 78076 153 78092 159
rect 78094 153 78110 159
rect 77901 143 77924 152
rect 78076 143 78099 152
rect 77874 133 77882 143
rect 77880 109 77882 133
rect 77890 123 77891 143
rect 77901 118 77904 143
rect 77923 123 77924 143
rect 77933 133 77940 143
rect 78060 133 78067 143
rect 78076 123 78077 143
rect 78096 118 78099 143
rect 78109 123 78110 143
rect 78119 133 78126 143
rect 77890 109 77924 113
rect 78076 109 78110 113
rect 78170 109 78172 159
rect 77776 103 77818 104
rect 78182 103 78224 104
rect 77776 96 77780 103
rect 77671 62 77676 96
rect 77700 62 77705 96
rect 77743 79 77814 96
rect 78186 79 78220 96
rect 78223 79 78257 96
rect 77743 62 77818 79
rect 77776 61 77818 62
rect 78182 62 78257 79
rect 78182 61 78224 62
rect 77754 55 77840 61
rect 78160 55 78246 61
rect 78288 55 78292 233
rect 78476 183 78480 251
rect 78485 207 78495 241
rect 78505 213 78525 241
rect 78505 207 78519 213
rect 78544 207 78555 251
rect 78586 246 78662 253
rect 78695 251 78704 279
rect 78607 228 78641 246
rect 78649 228 78651 246
rect 78586 221 78662 228
rect 78649 213 78651 221
rect 78693 213 78704 251
rect 78768 241 78772 395
rect 78775 378 78780 412
rect 78804 378 78809 412
rect 78810 400 78821 412
rect 79024 395 79066 421
rect 79430 395 79472 421
rect 79687 420 79699 424
rect 79709 420 79721 424
rect 79759 420 79771 424
rect 79781 421 79793 424
rect 79781 420 79834 421
rect 79792 412 79834 420
rect 79675 400 79686 412
rect 78956 341 78960 395
rect 79016 387 79062 395
rect 79016 383 79032 387
rect 79024 380 79032 383
rect 79058 380 79062 387
rect 79066 383 79074 395
rect 79422 383 79430 395
rect 79434 387 79468 395
rect 79434 380 79438 387
rect 79464 380 79468 387
rect 79472 383 79480 395
rect 79012 379 79078 380
rect 79418 379 79484 380
rect 79024 371 79028 379
rect 79078 365 79128 367
rect 79368 365 79418 367
rect 79118 361 79172 365
rect 79324 361 79378 365
rect 79118 356 79138 361
rect 79358 356 79378 361
rect 79128 341 79130 356
rect 78956 261 78960 329
rect 79024 305 79028 341
rect 79122 331 79130 341
rect 79138 331 79139 351
rect 79128 315 79130 331
rect 79149 322 79152 356
rect 79171 331 79172 351
rect 79181 331 79188 341
rect 79308 331 79315 341
rect 79324 331 79325 351
rect 79344 322 79347 356
rect 79357 331 79358 351
rect 79367 331 79374 341
rect 79138 315 79154 321
rect 79156 315 79172 321
rect 79324 315 79340 321
rect 79342 315 79358 321
rect 79418 315 79420 365
rect 78961 267 78997 295
rect 78961 261 78975 267
rect 78640 212 78651 213
rect 78485 183 78492 207
rect 78640 183 78650 212
rect 78731 207 78743 241
rect 78753 207 78773 241
rect 78476 103 78480 171
rect 78544 133 78548 183
rect 78544 98 78548 103
rect 78295 62 78300 96
rect 78324 62 78329 96
rect 78544 94 78582 98
rect 78544 79 78552 94
rect 78578 79 78582 94
rect 78666 94 78700 98
rect 78666 79 78670 94
rect 78696 79 78700 94
rect 78544 61 78586 79
rect 78662 61 78704 79
rect 78522 55 78608 61
rect 78640 55 78726 61
rect 78768 55 78772 207
rect 78798 183 78805 211
rect 78956 183 78960 251
rect 78965 233 78975 261
rect 78985 261 78999 267
rect 79024 261 79035 305
rect 79461 267 79472 305
rect 79499 267 79535 295
rect 79536 267 79540 395
rect 79687 378 79692 412
rect 79716 378 79721 412
rect 79722 400 79733 412
rect 79747 400 79758 412
rect 79759 395 79834 412
rect 79724 341 79728 395
rect 79759 378 79830 395
rect 79834 383 79842 395
rect 79792 371 79796 378
rect 79186 262 79236 264
rect 79260 262 79310 264
rect 78985 233 79005 261
rect 79024 233 79033 261
rect 79087 253 79121 261
rect 79066 246 79121 253
rect 79087 245 79121 246
rect 79189 253 79220 261
rect 79189 245 79223 253
rect 79024 213 79028 233
rect 79220 229 79223 245
rect 79087 228 79121 229
rect 79066 221 79121 228
rect 79189 221 79223 229
rect 79236 212 79238 262
rect 79276 253 79307 261
rect 79310 253 79312 262
rect 79499 261 79511 267
rect 79276 245 79312 253
rect 79375 253 79409 261
rect 79375 246 79430 253
rect 79375 245 79409 246
rect 79307 229 79312 245
rect 79501 233 79511 261
rect 79521 233 79541 267
rect 79724 261 79728 329
rect 79792 291 79796 341
rect 79792 251 79801 279
rect 79860 264 79872 265
rect 79847 262 79897 264
rect 79860 261 79872 262
rect 79855 253 79880 261
rect 79276 221 79312 229
rect 79375 228 79409 229
rect 79375 221 79430 228
rect 79310 212 79312 221
rect 78956 103 78960 171
rect 79024 133 79028 183
rect 79078 159 79128 161
rect 79368 159 79418 161
rect 79128 143 79130 159
rect 79138 153 79154 159
rect 79156 153 79172 159
rect 79324 153 79340 159
rect 79342 153 79358 159
rect 79149 143 79172 152
rect 79324 143 79347 152
rect 79122 133 79130 143
rect 79128 109 79130 133
rect 79138 123 79139 143
rect 79149 118 79152 143
rect 79171 123 79172 143
rect 79181 133 79188 143
rect 79308 133 79315 143
rect 79324 123 79325 143
rect 79344 118 79347 143
rect 79357 123 79358 143
rect 79367 133 79374 143
rect 79138 109 79172 113
rect 79324 109 79358 113
rect 79418 109 79420 159
rect 79024 103 79066 104
rect 79430 103 79472 104
rect 79024 96 79028 103
rect 78919 62 78924 96
rect 78948 62 78953 96
rect 78991 79 79062 96
rect 79434 79 79468 96
rect 79471 79 79505 96
rect 78991 62 79066 79
rect 79024 61 79066 62
rect 79430 62 79505 79
rect 79430 61 79472 62
rect 79002 55 79088 61
rect 79408 55 79494 61
rect 79536 55 79540 233
rect 79724 183 79728 251
rect 79733 207 79743 241
rect 79753 213 79773 241
rect 79753 207 79767 213
rect 79792 207 79803 251
rect 79834 246 79889 253
rect 79855 245 79889 246
rect 79864 229 79889 245
rect 79855 228 79889 229
rect 79834 221 79889 228
rect 79860 213 79880 221
rect 79860 209 79872 213
rect 79897 212 79899 262
rect 79733 183 79740 207
rect 79724 103 79728 171
rect 79792 133 79796 183
rect 79792 98 79796 103
rect 79543 62 79548 96
rect 79572 62 79577 96
rect 79792 94 79830 98
rect 79792 79 79800 94
rect 79826 79 79830 94
rect 79792 61 79834 79
rect 79770 55 79856 61
rect 38 39 80 55
rect 400 39 442 55
rect 806 39 848 55
rect 1168 39 1210 55
rect 1286 39 1328 55
rect 1648 39 1690 55
rect 2054 39 2096 55
rect 2416 39 2458 55
rect 2534 39 2576 55
rect 2896 39 2938 55
rect 3302 39 3344 55
rect 3664 39 3706 55
rect 3782 39 3824 55
rect 4144 39 4186 55
rect 4550 39 4592 55
rect 4912 39 4954 55
rect 5030 39 5072 55
rect 5392 39 5434 55
rect 5798 39 5840 55
rect 6160 39 6202 55
rect 6278 39 6320 55
rect 6640 39 6682 55
rect 7046 39 7088 55
rect 7408 39 7450 55
rect 7526 39 7568 55
rect 7888 39 7930 55
rect 8294 39 8336 55
rect 8656 39 8698 55
rect 8774 39 8816 55
rect 9136 39 9178 55
rect 9542 39 9584 55
rect 9904 39 9946 55
rect 10022 39 10064 55
rect 10384 39 10426 55
rect 10790 39 10832 55
rect 11152 39 11194 55
rect 11270 39 11312 55
rect 11632 39 11674 55
rect 12038 39 12080 55
rect 12400 39 12442 55
rect 12518 39 12560 55
rect 12880 39 12922 55
rect 13286 39 13328 55
rect 13648 39 13690 55
rect 13766 39 13808 55
rect 14128 39 14170 55
rect 14534 39 14576 55
rect 14896 39 14938 55
rect 15014 39 15056 55
rect 15376 39 15418 55
rect 15782 39 15824 55
rect 16144 39 16186 55
rect 16262 39 16304 55
rect 16624 39 16666 55
rect 17030 39 17072 55
rect 17392 39 17434 55
rect 17510 39 17552 55
rect 17872 39 17914 55
rect 18278 39 18320 55
rect 18640 39 18682 55
rect 18758 39 18800 55
rect 19120 39 19162 55
rect 19526 39 19568 55
rect 19888 39 19930 55
rect 20006 39 20048 55
rect 20368 39 20410 55
rect 20774 39 20816 55
rect 21136 39 21178 55
rect 21254 39 21296 55
rect 21616 39 21658 55
rect 22022 39 22064 55
rect 22384 39 22426 55
rect 22502 39 22544 55
rect 22864 39 22906 55
rect 23270 39 23312 55
rect 23632 39 23674 55
rect 23750 39 23792 55
rect 24112 39 24154 55
rect 24518 39 24560 55
rect 24880 39 24922 55
rect 24998 39 25040 55
rect 25360 39 25402 55
rect 25766 39 25808 55
rect 26128 39 26170 55
rect 26246 39 26288 55
rect 26608 39 26650 55
rect 27014 39 27056 55
rect 27376 39 27418 55
rect 27494 39 27536 55
rect 27856 39 27898 55
rect 28262 39 28304 55
rect 28624 39 28666 55
rect 28742 39 28784 55
rect 29104 39 29146 55
rect 29510 39 29552 55
rect 29872 39 29914 55
rect 29990 39 30032 55
rect 30352 39 30394 55
rect 30758 39 30800 55
rect 31120 39 31162 55
rect 31238 39 31280 55
rect 31600 39 31642 55
rect 32006 39 32048 55
rect 32368 39 32410 55
rect 32486 39 32528 55
rect 32848 39 32890 55
rect 33254 39 33296 55
rect 33616 39 33658 55
rect 33734 39 33776 55
rect 34096 39 34138 55
rect 34502 39 34544 55
rect 34864 39 34906 55
rect 34982 39 35024 55
rect 35344 39 35386 55
rect 35750 39 35792 55
rect 36112 39 36154 55
rect 36230 39 36272 55
rect 36592 39 36634 55
rect 36998 39 37040 55
rect 37360 39 37402 55
rect 37478 39 37520 55
rect 37840 39 37882 55
rect 38246 39 38288 55
rect 38608 39 38650 55
rect 38726 39 38768 55
rect 39088 39 39130 55
rect 39494 39 39536 55
rect 39856 39 39898 55
rect 39974 39 40016 55
rect 40336 39 40378 55
rect 40742 39 40784 55
rect 41104 39 41146 55
rect 41222 39 41264 55
rect 41584 39 41626 55
rect 41990 39 42032 55
rect 42352 39 42394 55
rect 42470 39 42512 55
rect 42832 39 42874 55
rect 43238 39 43280 55
rect 43600 39 43642 55
rect 43718 39 43760 55
rect 44080 39 44122 55
rect 44486 39 44528 55
rect 44848 39 44890 55
rect 44966 39 45008 55
rect 45328 39 45370 55
rect 45734 39 45776 55
rect 46096 39 46138 55
rect 46214 39 46256 55
rect 46576 39 46618 55
rect 46982 39 47024 55
rect 47344 39 47386 55
rect 47462 39 47504 55
rect 47824 39 47866 55
rect 48230 39 48272 55
rect 48592 39 48634 55
rect 48710 39 48752 55
rect 49072 39 49114 55
rect 49478 39 49520 55
rect 49840 39 49882 55
rect 49958 39 50000 55
rect 50320 39 50362 55
rect 50726 39 50768 55
rect 51088 39 51130 55
rect 51206 39 51248 55
rect 51568 39 51610 55
rect 51974 39 52016 55
rect 52336 39 52378 55
rect 52454 39 52496 55
rect 52816 39 52858 55
rect 53222 39 53264 55
rect 53584 39 53626 55
rect 53702 39 53744 55
rect 54064 39 54106 55
rect 54470 39 54512 55
rect 54832 39 54874 55
rect 54950 39 54992 55
rect 55312 39 55354 55
rect 55718 39 55760 55
rect 56080 39 56122 55
rect 56198 39 56240 55
rect 56560 39 56602 55
rect 56966 39 57008 55
rect 57328 39 57370 55
rect 57446 39 57488 55
rect 57808 39 57850 55
rect 58214 39 58256 55
rect 58576 39 58618 55
rect 58694 39 58736 55
rect 59056 39 59098 55
rect 59462 39 59504 55
rect 59824 39 59866 55
rect 59942 39 59984 55
rect 60304 39 60346 55
rect 60710 39 60752 55
rect 61072 39 61114 55
rect 61190 39 61232 55
rect 61552 39 61594 55
rect 61958 39 62000 55
rect 62320 39 62362 55
rect 62438 39 62480 55
rect 62800 39 62842 55
rect 63206 39 63248 55
rect 63568 39 63610 55
rect 63686 39 63728 55
rect 64048 39 64090 55
rect 64454 39 64496 55
rect 64816 39 64858 55
rect 64934 39 64976 55
rect 65296 39 65338 55
rect 65702 39 65744 55
rect 66064 39 66106 55
rect 66182 39 66224 55
rect 66544 39 66586 55
rect 66950 39 66992 55
rect 67312 39 67354 55
rect 67430 39 67472 55
rect 67792 39 67834 55
rect 68198 39 68240 55
rect 68560 39 68602 55
rect 68678 39 68720 55
rect 69040 39 69082 55
rect 69446 39 69488 55
rect 69808 39 69850 55
rect 69926 39 69968 55
rect 70288 39 70330 55
rect 70694 39 70736 55
rect 71056 39 71098 55
rect 71174 39 71216 55
rect 71536 39 71578 55
rect 71942 39 71984 55
rect 72304 39 72346 55
rect 72422 39 72464 55
rect 72784 39 72826 55
rect 73190 39 73232 55
rect 73552 39 73594 55
rect 73670 39 73712 55
rect 74032 39 74074 55
rect 74438 39 74480 55
rect 74800 39 74842 55
rect 74918 39 74960 55
rect 75280 39 75322 55
rect 75686 39 75728 55
rect 76048 39 76090 55
rect 76166 39 76208 55
rect 76528 39 76570 55
rect 76934 39 76976 55
rect 77296 39 77338 55
rect 77414 39 77456 55
rect 77776 39 77818 55
rect 78182 39 78224 55
rect 78544 39 78586 55
rect 78662 39 78704 55
rect 79024 39 79066 55
rect 79430 39 79472 55
rect 79792 39 79834 55
rect -25 25 25 27
rect 42 25 76 39
rect 404 25 438 39
rect 455 25 505 27
rect 557 25 607 27
rect 641 25 691 27
rect 743 25 793 27
rect 810 25 844 39
rect 1172 25 1206 39
rect 1223 25 1273 27
rect 1290 25 1324 39
rect 1652 25 1686 39
rect 1703 25 1753 27
rect 1805 25 1855 27
rect 1889 25 1939 27
rect 1991 25 2041 27
rect 2058 25 2092 39
rect 2420 25 2454 39
rect 2471 25 2521 27
rect 2538 25 2572 39
rect 2900 25 2934 39
rect 2951 25 3001 27
rect 3053 25 3103 27
rect 3137 25 3187 27
rect 3239 25 3289 27
rect 3306 25 3340 39
rect 3668 25 3702 39
rect 3719 25 3769 27
rect 3786 25 3820 39
rect 4148 25 4182 39
rect 4199 25 4249 27
rect 4301 25 4351 27
rect 4385 25 4435 27
rect 4487 25 4537 27
rect 4554 25 4588 39
rect 4916 25 4950 39
rect 4967 25 5017 27
rect 5034 25 5068 39
rect 5396 25 5430 39
rect 5447 25 5497 27
rect 5549 25 5599 27
rect 5633 25 5683 27
rect 5735 25 5785 27
rect 5802 25 5836 39
rect 6164 25 6198 39
rect 6215 25 6265 27
rect 6282 25 6316 39
rect 6644 25 6678 39
rect 6695 25 6745 27
rect 6797 25 6847 27
rect 6881 25 6931 27
rect 6983 25 7033 27
rect 7050 25 7084 39
rect 7412 25 7446 39
rect 7463 25 7513 27
rect 7530 25 7564 39
rect 7892 25 7926 39
rect 7943 25 7993 27
rect 8045 25 8095 27
rect 8129 25 8179 27
rect 8231 25 8281 27
rect 8298 25 8332 39
rect 8660 25 8694 39
rect 8711 25 8761 27
rect 8778 25 8812 39
rect 9140 25 9174 39
rect 9191 25 9241 27
rect 9293 25 9343 27
rect 9377 25 9427 27
rect 9479 25 9529 27
rect 9546 25 9580 39
rect 9908 25 9942 39
rect 9959 25 10009 27
rect 10026 25 10060 39
rect 10388 25 10422 39
rect 10439 25 10489 27
rect 10541 25 10591 27
rect 10625 25 10675 27
rect 10727 25 10777 27
rect 10794 25 10828 39
rect 11156 25 11190 39
rect 11207 25 11257 27
rect 11274 25 11308 39
rect 11636 25 11670 39
rect 11687 25 11737 27
rect 11789 25 11839 27
rect 11873 25 11923 27
rect 11975 25 12025 27
rect 12042 25 12076 39
rect 12404 25 12438 39
rect 12455 25 12505 27
rect 12522 25 12556 39
rect 12884 25 12918 39
rect 12935 25 12985 27
rect 13037 25 13087 27
rect 13121 25 13171 27
rect 13223 25 13273 27
rect 13290 25 13324 39
rect 13652 25 13686 39
rect 13703 25 13753 27
rect 13770 25 13804 39
rect 14132 25 14166 39
rect 14183 25 14233 27
rect 14285 25 14335 27
rect 14369 25 14419 27
rect 14471 25 14521 27
rect 14538 25 14572 39
rect 14900 25 14934 39
rect 14951 25 15001 27
rect 15018 25 15052 39
rect 15380 25 15414 39
rect 15431 25 15481 27
rect 15533 25 15583 27
rect 15617 25 15667 27
rect 15719 25 15769 27
rect 15786 25 15820 39
rect 16148 25 16182 39
rect 16199 25 16249 27
rect 16266 25 16300 39
rect 16628 25 16662 39
rect 16679 25 16729 27
rect 16781 25 16831 27
rect 16865 25 16915 27
rect 16967 25 17017 27
rect 17034 25 17068 39
rect 17396 25 17430 39
rect 17447 25 17497 27
rect 17514 25 17548 39
rect 17876 25 17910 39
rect 17927 25 17977 27
rect 18029 25 18079 27
rect 18113 25 18163 27
rect 18215 25 18265 27
rect 18282 25 18316 39
rect 18644 25 18678 39
rect 18695 25 18745 27
rect 18762 25 18796 39
rect 19124 25 19158 39
rect 19175 25 19225 27
rect 19277 25 19327 27
rect 19361 25 19411 27
rect 19463 25 19513 27
rect 19530 25 19564 39
rect 19892 25 19926 39
rect 19943 25 19993 27
rect 20010 25 20044 39
rect 20372 25 20406 39
rect 20423 25 20473 27
rect 20525 25 20575 27
rect 20609 25 20659 27
rect 20711 25 20761 27
rect 20778 25 20812 39
rect 21140 25 21174 39
rect 21191 25 21241 27
rect 21258 25 21292 39
rect 21620 25 21654 39
rect 21671 25 21721 27
rect 21773 25 21823 27
rect 21857 25 21907 27
rect 21959 25 22009 27
rect 22026 25 22060 39
rect 22388 25 22422 39
rect 22439 25 22489 27
rect 22506 25 22540 39
rect 22868 25 22902 39
rect 22919 25 22969 27
rect 23021 25 23071 27
rect 23105 25 23155 27
rect 23207 25 23257 27
rect 23274 25 23308 39
rect 23636 25 23670 39
rect 23687 25 23737 27
rect 23754 25 23788 39
rect 24116 25 24150 39
rect 24167 25 24217 27
rect 24269 25 24319 27
rect 24353 25 24403 27
rect 24455 25 24505 27
rect 24522 25 24556 39
rect 24884 25 24918 39
rect 24935 25 24985 27
rect 25002 25 25036 39
rect 25364 25 25398 39
rect 25415 25 25465 27
rect 25517 25 25567 27
rect 25601 25 25651 27
rect 25703 25 25753 27
rect 25770 25 25804 39
rect 26132 25 26166 39
rect 26183 25 26233 27
rect 26250 25 26284 39
rect 26612 25 26646 39
rect 26663 25 26713 27
rect 26765 25 26815 27
rect 26849 25 26899 27
rect 26951 25 27001 27
rect 27018 25 27052 39
rect 27380 25 27414 39
rect 27431 25 27481 27
rect 27498 25 27532 39
rect 27860 25 27894 39
rect 27911 25 27961 27
rect 28013 25 28063 27
rect 28097 25 28147 27
rect 28199 25 28249 27
rect 28266 25 28300 39
rect 28628 25 28662 39
rect 28679 25 28729 27
rect 28746 25 28780 39
rect 29108 25 29142 39
rect 29159 25 29209 27
rect 29261 25 29311 27
rect 29345 25 29395 27
rect 29447 25 29497 27
rect 29514 25 29548 39
rect 29876 25 29910 39
rect 29927 25 29977 27
rect 29994 25 30028 39
rect 30356 25 30390 39
rect 30407 25 30457 27
rect 30509 25 30559 27
rect 30593 25 30643 27
rect 30695 25 30745 27
rect 30762 25 30796 39
rect 31124 25 31158 39
rect 31175 25 31225 27
rect 31242 25 31276 39
rect 31604 25 31638 39
rect 31655 25 31705 27
rect 31757 25 31807 27
rect 31841 25 31891 27
rect 31943 25 31993 27
rect 32010 25 32044 39
rect 32372 25 32406 39
rect 32423 25 32473 27
rect 32490 25 32524 39
rect 32852 25 32886 39
rect 32903 25 32953 27
rect 33005 25 33055 27
rect 33089 25 33139 27
rect 33191 25 33241 27
rect 33258 25 33292 39
rect 33620 25 33654 39
rect 33671 25 33721 27
rect 33738 25 33772 39
rect 34100 25 34134 39
rect 34151 25 34201 27
rect 34253 25 34303 27
rect 34337 25 34387 27
rect 34439 25 34489 27
rect 34506 25 34540 39
rect 34868 25 34902 39
rect 34919 25 34969 27
rect 34986 25 35020 39
rect 35348 25 35382 39
rect 35399 25 35449 27
rect 35501 25 35551 27
rect 35585 25 35635 27
rect 35687 25 35737 27
rect 35754 25 35788 39
rect 36116 25 36150 39
rect 36167 25 36217 27
rect 36234 25 36268 39
rect 36596 25 36630 39
rect 36647 25 36697 27
rect 36749 25 36799 27
rect 36833 25 36883 27
rect 36935 25 36985 27
rect 37002 25 37036 39
rect 37364 25 37398 39
rect 37415 25 37465 27
rect 37482 25 37516 39
rect 37844 25 37878 39
rect 37895 25 37945 27
rect 37997 25 38047 27
rect 38081 25 38131 27
rect 38183 25 38233 27
rect 38250 25 38284 39
rect 38612 25 38646 39
rect 38663 25 38713 27
rect 38730 25 38764 39
rect 39092 25 39126 39
rect 39143 25 39193 27
rect 39245 25 39295 27
rect 39329 25 39379 27
rect 39431 25 39481 27
rect 39498 25 39532 39
rect 39860 25 39894 39
rect 39911 25 39961 27
rect 39978 25 40012 39
rect 40340 25 40374 39
rect 40391 25 40441 27
rect 40493 25 40543 27
rect 40577 25 40627 27
rect 40679 25 40729 27
rect 40746 25 40780 39
rect 41108 25 41142 39
rect 41159 25 41209 27
rect 41226 25 41260 39
rect 41588 25 41622 39
rect 41639 25 41689 27
rect 41741 25 41791 27
rect 41825 25 41875 27
rect 41927 25 41977 27
rect 41994 25 42028 39
rect 42356 25 42390 39
rect 42407 25 42457 27
rect 42474 25 42508 39
rect 42836 25 42870 39
rect 42887 25 42937 27
rect 42989 25 43039 27
rect 43073 25 43123 27
rect 43175 25 43225 27
rect 43242 25 43276 39
rect 43604 25 43638 39
rect 43655 25 43705 27
rect 43722 25 43756 39
rect 44084 25 44118 39
rect 44135 25 44185 27
rect 44237 25 44287 27
rect 44321 25 44371 27
rect 44423 25 44473 27
rect 44490 25 44524 39
rect 44852 25 44886 39
rect 44903 25 44953 27
rect 44970 25 45004 39
rect 45332 25 45366 39
rect 45383 25 45433 27
rect 45485 25 45535 27
rect 45569 25 45619 27
rect 45671 25 45721 27
rect 45738 25 45772 39
rect 46100 25 46134 39
rect 46151 25 46201 27
rect 46218 25 46252 39
rect 46580 25 46614 39
rect 46631 25 46681 27
rect 46733 25 46783 27
rect 46817 25 46867 27
rect 46919 25 46969 27
rect 46986 25 47020 39
rect 47348 25 47382 39
rect 47399 25 47449 27
rect 47466 25 47500 39
rect 47828 25 47862 39
rect 47879 25 47929 27
rect 47981 25 48031 27
rect 48065 25 48115 27
rect 48167 25 48217 27
rect 48234 25 48268 39
rect 48596 25 48630 39
rect 48647 25 48697 27
rect 48714 25 48748 39
rect 49076 25 49110 39
rect 49127 25 49177 27
rect 49229 25 49279 27
rect 49313 25 49363 27
rect 49415 25 49465 27
rect 49482 25 49516 39
rect 49844 25 49878 39
rect 49895 25 49945 27
rect 49962 25 49996 39
rect 50324 25 50358 39
rect 50375 25 50425 27
rect 50477 25 50527 27
rect 50561 25 50611 27
rect 50663 25 50713 27
rect 50730 25 50764 39
rect 51092 25 51126 39
rect 51143 25 51193 27
rect 51210 25 51244 39
rect 51572 25 51606 39
rect 51623 25 51673 27
rect 51725 25 51775 27
rect 51809 25 51859 27
rect 51911 25 51961 27
rect 51978 25 52012 39
rect 52340 25 52374 39
rect 52391 25 52441 27
rect 52458 25 52492 39
rect 52820 25 52854 39
rect 52871 25 52921 27
rect 52973 25 53023 27
rect 53057 25 53107 27
rect 53159 25 53209 27
rect 53226 25 53260 39
rect 53588 25 53622 39
rect 53639 25 53689 27
rect 53706 25 53740 39
rect 54068 25 54102 39
rect 54119 25 54169 27
rect 54221 25 54271 27
rect 54305 25 54355 27
rect 54407 25 54457 27
rect 54474 25 54508 39
rect 54836 25 54870 39
rect 54887 25 54937 27
rect 54954 25 54988 39
rect 55316 25 55350 39
rect 55367 25 55417 27
rect 55469 25 55519 27
rect 55553 25 55603 27
rect 55655 25 55705 27
rect 55722 25 55756 39
rect 56084 25 56118 39
rect 56135 25 56185 27
rect 56202 25 56236 39
rect 56564 25 56598 39
rect 56615 25 56665 27
rect 56717 25 56767 27
rect 56801 25 56851 27
rect 56903 25 56953 27
rect 56970 25 57004 39
rect 57332 25 57366 39
rect 57383 25 57433 27
rect 57450 25 57484 39
rect 57812 25 57846 39
rect 57863 25 57913 27
rect 57965 25 58015 27
rect 58049 25 58099 27
rect 58151 25 58201 27
rect 58218 25 58252 39
rect 58580 25 58614 39
rect 58631 25 58681 27
rect 58698 25 58732 39
rect 59060 25 59094 39
rect 59111 25 59161 27
rect 59213 25 59263 27
rect 59297 25 59347 27
rect 59399 25 59449 27
rect 59466 25 59500 39
rect 59828 25 59862 39
rect 59879 25 59929 27
rect 59946 25 59980 39
rect 60308 25 60342 39
rect 60359 25 60409 27
rect 60461 25 60511 27
rect 60545 25 60595 27
rect 60647 25 60697 27
rect 60714 25 60748 39
rect 61076 25 61110 39
rect 61127 25 61177 27
rect 61194 25 61228 39
rect 61556 25 61590 39
rect 61607 25 61657 27
rect 61709 25 61759 27
rect 61793 25 61843 27
rect 61895 25 61945 27
rect 61962 25 61996 39
rect 62324 25 62358 39
rect 62375 25 62425 27
rect 62442 25 62476 39
rect 62804 25 62838 39
rect 62855 25 62905 27
rect 62957 25 63007 27
rect 63041 25 63091 27
rect 63143 25 63193 27
rect 63210 25 63244 39
rect 63572 25 63606 39
rect 63623 25 63673 27
rect 63690 25 63724 39
rect 64052 25 64086 39
rect 64103 25 64153 27
rect 64205 25 64255 27
rect 64289 25 64339 27
rect 64391 25 64441 27
rect 64458 25 64492 39
rect 64820 25 64854 39
rect 64871 25 64921 27
rect 64938 25 64972 39
rect 65300 25 65334 39
rect 65351 25 65401 27
rect 65453 25 65503 27
rect 65537 25 65587 27
rect 65639 25 65689 27
rect 65706 25 65740 39
rect 66068 25 66102 39
rect 66119 25 66169 27
rect 66186 25 66220 39
rect 66548 25 66582 39
rect 66599 25 66649 27
rect 66701 25 66751 27
rect 66785 25 66835 27
rect 66887 25 66937 27
rect 66954 25 66988 39
rect 67316 25 67350 39
rect 67367 25 67417 27
rect 67434 25 67468 39
rect 67796 25 67830 39
rect 67847 25 67897 27
rect 67949 25 67999 27
rect 68033 25 68083 27
rect 68135 25 68185 27
rect 68202 25 68236 39
rect 68564 25 68598 39
rect 68615 25 68665 27
rect 68682 25 68716 39
rect 69044 25 69078 39
rect 69095 25 69145 27
rect 69197 25 69247 27
rect 69281 25 69331 27
rect 69383 25 69433 27
rect 69450 25 69484 39
rect 69812 25 69846 39
rect 69863 25 69913 27
rect 69930 25 69964 39
rect 70292 25 70326 39
rect 70343 25 70393 27
rect 70445 25 70495 27
rect 70529 25 70579 27
rect 70631 25 70681 27
rect 70698 25 70732 39
rect 71060 25 71094 39
rect 71111 25 71161 27
rect 71178 25 71212 39
rect 71540 25 71574 39
rect 71591 25 71641 27
rect 71693 25 71743 27
rect 71777 25 71827 27
rect 71879 25 71929 27
rect 71946 25 71980 39
rect 72308 25 72342 39
rect 72359 25 72409 27
rect 72426 25 72460 39
rect 72788 25 72822 39
rect 72839 25 72889 27
rect 72941 25 72991 27
rect 73025 25 73075 27
rect 73127 25 73177 27
rect 73194 25 73228 39
rect 73556 25 73590 39
rect 73607 25 73657 27
rect 73674 25 73708 39
rect 74036 25 74070 39
rect 74087 25 74137 27
rect 74189 25 74239 27
rect 74273 25 74323 27
rect 74375 25 74425 27
rect 74442 25 74476 39
rect 74804 25 74838 39
rect 74855 25 74905 27
rect 74922 25 74956 39
rect 75284 25 75318 39
rect 75335 25 75385 27
rect 75437 25 75487 27
rect 75521 25 75571 27
rect 75623 25 75673 27
rect 75690 25 75724 39
rect 76052 25 76086 39
rect 76103 25 76153 27
rect 76170 25 76204 39
rect 76532 25 76566 39
rect 76583 25 76633 27
rect 76685 25 76735 27
rect 76769 25 76819 27
rect 76871 25 76921 27
rect 76938 25 76972 39
rect 77300 25 77334 39
rect 77351 25 77401 27
rect 77418 25 77452 39
rect 77780 25 77814 39
rect 77831 25 77881 27
rect 77933 25 77983 27
rect 78017 25 78067 27
rect 78119 25 78169 27
rect 78186 25 78220 39
rect 78548 25 78582 39
rect 78599 25 78649 27
rect 78666 25 78700 39
rect 79028 25 79062 39
rect 79079 25 79129 27
rect 79181 25 79231 27
rect 79265 25 79315 27
rect 79367 25 79417 27
rect 79434 25 79468 39
rect 79796 25 79830 39
rect 79847 25 79897 27
rect 16 17 102 25
rect 378 17 464 25
rect 8 -17 17 17
rect 18 15 51 17
rect 80 15 100 17
rect 18 -17 100 15
rect 380 15 404 17
rect 429 15 438 17
rect 442 15 462 17
rect 16 -25 102 -17
rect 42 -41 76 -25
rect 16 -61 38 -55
rect 80 -61 102 -55
rect 144 -79 148 0
rect 332 -55 336 0
rect 380 -17 462 15
rect 463 -17 472 17
rect 480 -17 497 17
rect 378 -25 464 -17
rect 505 -25 507 25
rect 514 -17 548 17
rect 565 -17 582 17
rect 607 -25 609 25
rect 666 -17 683 17
rect 691 -25 693 25
rect 784 17 870 25
rect 1146 17 1232 25
rect 1264 17 1350 25
rect 1626 17 1712 25
rect 700 -17 734 17
rect 751 -17 768 17
rect 776 -17 785 17
rect 786 15 819 17
rect 848 15 868 17
rect 786 -17 868 15
rect 1148 15 1172 17
rect 1197 15 1206 17
rect 1210 15 1230 17
rect 784 -25 870 -17
rect 404 -41 438 -25
rect 810 -41 844 -25
rect 378 -61 404 -55
rect 442 -61 464 -55
rect 784 -61 806 -55
rect 848 -61 870 -55
rect 400 -79 404 -61
rect 912 -79 916 0
rect 1100 -55 1104 0
rect 1148 -17 1230 15
rect 1231 -17 1240 17
rect 1256 -17 1265 17
rect 1266 15 1299 17
rect 1328 15 1348 17
rect 1266 -17 1348 15
rect 1628 15 1652 17
rect 1677 15 1686 17
rect 1690 15 1710 17
rect 1146 -25 1232 -17
rect 1264 -25 1350 -17
rect 1172 -41 1206 -25
rect 1290 -41 1324 -25
rect 1146 -61 1172 -55
rect 1210 -61 1232 -55
rect 1264 -61 1286 -55
rect 1328 -61 1350 -55
rect 1168 -79 1172 -61
rect 1392 -79 1396 0
rect 1580 -55 1584 0
rect 1628 -17 1710 15
rect 1711 -17 1720 17
rect 1728 -17 1745 17
rect 1626 -25 1712 -17
rect 1753 -25 1755 25
rect 1762 -17 1796 17
rect 1813 -17 1830 17
rect 1855 -25 1857 25
rect 1914 -17 1931 17
rect 1939 -25 1941 25
rect 2032 17 2118 25
rect 2394 17 2480 25
rect 2512 17 2598 25
rect 2874 17 2960 25
rect 1948 -17 1982 17
rect 1999 -17 2016 17
rect 2024 -17 2033 17
rect 2034 15 2067 17
rect 2096 15 2116 17
rect 2034 -17 2116 15
rect 2396 15 2420 17
rect 2445 15 2454 17
rect 2458 15 2478 17
rect 2032 -25 2118 -17
rect 1652 -41 1686 -25
rect 2058 -41 2092 -25
rect 1626 -61 1652 -55
rect 1690 -61 1712 -55
rect 2032 -61 2054 -55
rect 2096 -61 2118 -55
rect 1648 -79 1652 -61
rect 2160 -79 2164 0
rect 2348 -55 2352 0
rect 2396 -17 2478 15
rect 2479 -17 2488 17
rect 2504 -17 2513 17
rect 2514 15 2547 17
rect 2576 15 2596 17
rect 2514 -17 2596 15
rect 2876 15 2900 17
rect 2925 15 2934 17
rect 2938 15 2958 17
rect 2394 -25 2480 -17
rect 2512 -25 2598 -17
rect 2420 -41 2454 -25
rect 2538 -41 2572 -25
rect 2394 -61 2420 -55
rect 2458 -61 2480 -55
rect 2512 -61 2534 -55
rect 2576 -61 2598 -55
rect 2416 -79 2420 -61
rect 2640 -79 2644 0
rect 2828 -55 2832 0
rect 2876 -17 2958 15
rect 2959 -17 2968 17
rect 2976 -17 2993 17
rect 2874 -25 2960 -17
rect 3001 -25 3003 25
rect 3010 -17 3044 17
rect 3061 -17 3078 17
rect 3103 -25 3105 25
rect 3162 -17 3179 17
rect 3187 -25 3189 25
rect 3280 17 3366 25
rect 3642 17 3728 25
rect 3760 17 3846 25
rect 4122 17 4208 25
rect 3196 -17 3230 17
rect 3247 -17 3264 17
rect 3272 -17 3281 17
rect 3282 15 3315 17
rect 3344 15 3364 17
rect 3282 -17 3364 15
rect 3644 15 3668 17
rect 3693 15 3702 17
rect 3706 15 3726 17
rect 3280 -25 3366 -17
rect 2900 -41 2934 -25
rect 3306 -41 3340 -25
rect 2874 -61 2900 -55
rect 2938 -61 2960 -55
rect 3280 -61 3302 -55
rect 3344 -61 3366 -55
rect 2896 -79 2900 -61
rect 3408 -79 3412 0
rect 3596 -55 3600 0
rect 3644 -17 3726 15
rect 3727 -17 3736 17
rect 3752 -17 3761 17
rect 3762 15 3795 17
rect 3824 15 3844 17
rect 3762 -17 3844 15
rect 4124 15 4148 17
rect 4173 15 4182 17
rect 4186 15 4206 17
rect 3642 -25 3728 -17
rect 3760 -25 3846 -17
rect 3668 -41 3702 -25
rect 3786 -41 3820 -25
rect 3642 -61 3668 -55
rect 3706 -61 3728 -55
rect 3760 -61 3782 -55
rect 3824 -61 3846 -55
rect 3664 -79 3668 -61
rect 3888 -79 3892 0
rect 4076 -55 4080 0
rect 4124 -17 4206 15
rect 4207 -17 4216 17
rect 4224 -17 4241 17
rect 4122 -25 4208 -17
rect 4249 -25 4251 25
rect 4258 -17 4292 17
rect 4309 -17 4326 17
rect 4351 -25 4353 25
rect 4410 -17 4427 17
rect 4435 -25 4437 25
rect 4528 17 4614 25
rect 4890 17 4976 25
rect 5008 17 5094 25
rect 5370 17 5456 25
rect 4444 -17 4478 17
rect 4495 -17 4512 17
rect 4520 -17 4529 17
rect 4530 15 4563 17
rect 4592 15 4612 17
rect 4530 -17 4612 15
rect 4892 15 4916 17
rect 4941 15 4950 17
rect 4954 15 4974 17
rect 4528 -25 4614 -17
rect 4148 -41 4182 -25
rect 4554 -41 4588 -25
rect 4122 -61 4148 -55
rect 4186 -61 4208 -55
rect 4528 -61 4550 -55
rect 4592 -61 4614 -55
rect 4144 -79 4148 -61
rect 4656 -79 4660 0
rect 4844 -55 4848 0
rect 4892 -17 4974 15
rect 4975 -17 4984 17
rect 5000 -17 5009 17
rect 5010 15 5043 17
rect 5072 15 5092 17
rect 5010 -17 5092 15
rect 5372 15 5396 17
rect 5421 15 5430 17
rect 5434 15 5454 17
rect 4890 -25 4976 -17
rect 5008 -25 5094 -17
rect 4916 -41 4950 -25
rect 5034 -41 5068 -25
rect 4890 -61 4916 -55
rect 4954 -61 4976 -55
rect 5008 -61 5030 -55
rect 5072 -61 5094 -55
rect 4912 -79 4916 -61
rect 5136 -79 5140 0
rect 5324 -55 5328 0
rect 5372 -17 5454 15
rect 5455 -17 5464 17
rect 5472 -17 5489 17
rect 5370 -25 5456 -17
rect 5497 -25 5499 25
rect 5506 -17 5540 17
rect 5557 -17 5574 17
rect 5599 -25 5601 25
rect 5658 -17 5675 17
rect 5683 -25 5685 25
rect 5776 17 5862 25
rect 6138 17 6224 25
rect 6256 17 6342 25
rect 6618 17 6704 25
rect 5692 -17 5726 17
rect 5743 -17 5760 17
rect 5768 -17 5777 17
rect 5778 15 5811 17
rect 5840 15 5860 17
rect 5778 -17 5860 15
rect 6140 15 6164 17
rect 6189 15 6198 17
rect 6202 15 6222 17
rect 5776 -25 5862 -17
rect 5396 -41 5430 -25
rect 5802 -41 5836 -25
rect 5370 -61 5396 -55
rect 5434 -61 5456 -55
rect 5776 -61 5798 -55
rect 5840 -61 5862 -55
rect 5392 -79 5396 -61
rect 5904 -79 5908 0
rect 6092 -55 6096 0
rect 6140 -17 6222 15
rect 6223 -17 6232 17
rect 6248 -17 6257 17
rect 6258 15 6291 17
rect 6320 15 6340 17
rect 6258 -17 6340 15
rect 6620 15 6644 17
rect 6669 15 6678 17
rect 6682 15 6702 17
rect 6138 -25 6224 -17
rect 6256 -25 6342 -17
rect 6164 -41 6198 -25
rect 6282 -41 6316 -25
rect 6138 -61 6164 -55
rect 6202 -61 6224 -55
rect 6256 -61 6278 -55
rect 6320 -61 6342 -55
rect 6160 -79 6164 -61
rect 6384 -79 6388 0
rect 6572 -55 6576 0
rect 6620 -17 6702 15
rect 6703 -17 6712 17
rect 6720 -17 6737 17
rect 6618 -25 6704 -17
rect 6745 -25 6747 25
rect 6754 -17 6788 17
rect 6805 -17 6822 17
rect 6847 -25 6849 25
rect 6906 -17 6923 17
rect 6931 -25 6933 25
rect 7024 17 7110 25
rect 7386 17 7472 25
rect 7504 17 7590 25
rect 7866 17 7952 25
rect 6940 -17 6974 17
rect 6991 -17 7008 17
rect 7016 -17 7025 17
rect 7026 15 7059 17
rect 7088 15 7108 17
rect 7026 -17 7108 15
rect 7388 15 7412 17
rect 7437 15 7446 17
rect 7450 15 7470 17
rect 7024 -25 7110 -17
rect 6644 -41 6678 -25
rect 7050 -41 7084 -25
rect 6618 -61 6644 -55
rect 6682 -61 6704 -55
rect 7024 -61 7046 -55
rect 7088 -61 7110 -55
rect 6640 -79 6644 -61
rect 7152 -79 7156 0
rect 7340 -55 7344 0
rect 7388 -17 7470 15
rect 7471 -17 7480 17
rect 7496 -17 7505 17
rect 7506 15 7539 17
rect 7568 15 7588 17
rect 7506 -17 7588 15
rect 7868 15 7892 17
rect 7917 15 7926 17
rect 7930 15 7950 17
rect 7386 -25 7472 -17
rect 7504 -25 7590 -17
rect 7412 -41 7446 -25
rect 7530 -41 7564 -25
rect 7386 -61 7412 -55
rect 7450 -61 7472 -55
rect 7504 -61 7526 -55
rect 7568 -61 7590 -55
rect 7408 -79 7412 -61
rect 7632 -79 7636 0
rect 7820 -55 7824 0
rect 7868 -17 7950 15
rect 7951 -17 7960 17
rect 7968 -17 7985 17
rect 7866 -25 7952 -17
rect 7993 -25 7995 25
rect 8002 -17 8036 17
rect 8053 -17 8070 17
rect 8095 -25 8097 25
rect 8154 -17 8171 17
rect 8179 -25 8181 25
rect 8272 17 8358 25
rect 8634 17 8720 25
rect 8752 17 8838 25
rect 9114 17 9200 25
rect 8188 -17 8222 17
rect 8239 -17 8256 17
rect 8264 -17 8273 17
rect 8274 15 8307 17
rect 8336 15 8356 17
rect 8274 -17 8356 15
rect 8636 15 8660 17
rect 8685 15 8694 17
rect 8698 15 8718 17
rect 8272 -25 8358 -17
rect 7892 -41 7926 -25
rect 8298 -41 8332 -25
rect 7866 -61 7892 -55
rect 7930 -61 7952 -55
rect 8272 -61 8294 -55
rect 8336 -61 8358 -55
rect 7888 -79 7892 -61
rect 8400 -79 8404 0
rect 8588 -55 8592 0
rect 8636 -17 8718 15
rect 8719 -17 8728 17
rect 8744 -17 8753 17
rect 8754 15 8787 17
rect 8816 15 8836 17
rect 8754 -17 8836 15
rect 9116 15 9140 17
rect 9165 15 9174 17
rect 9178 15 9198 17
rect 8634 -25 8720 -17
rect 8752 -25 8838 -17
rect 8660 -41 8694 -25
rect 8778 -41 8812 -25
rect 8634 -61 8660 -55
rect 8698 -61 8720 -55
rect 8752 -61 8774 -55
rect 8816 -61 8838 -55
rect 8656 -79 8660 -61
rect 8880 -79 8884 0
rect 9068 -55 9072 0
rect 9116 -17 9198 15
rect 9199 -17 9208 17
rect 9216 -17 9233 17
rect 9114 -25 9200 -17
rect 9241 -25 9243 25
rect 9250 -17 9284 17
rect 9301 -17 9318 17
rect 9343 -25 9345 25
rect 9402 -17 9419 17
rect 9427 -25 9429 25
rect 9520 17 9606 25
rect 9882 17 9968 25
rect 10000 17 10086 25
rect 10362 17 10448 25
rect 9436 -17 9470 17
rect 9487 -17 9504 17
rect 9512 -17 9521 17
rect 9522 15 9555 17
rect 9584 15 9604 17
rect 9522 -17 9604 15
rect 9884 15 9908 17
rect 9933 15 9942 17
rect 9946 15 9966 17
rect 9520 -25 9606 -17
rect 9140 -41 9174 -25
rect 9546 -41 9580 -25
rect 9114 -61 9140 -55
rect 9178 -61 9200 -55
rect 9520 -61 9542 -55
rect 9584 -61 9606 -55
rect 9136 -79 9140 -61
rect 9648 -79 9652 0
rect 9836 -55 9840 0
rect 9884 -17 9966 15
rect 9967 -17 9976 17
rect 9992 -17 10001 17
rect 10002 15 10035 17
rect 10064 15 10084 17
rect 10002 -17 10084 15
rect 10364 15 10388 17
rect 10413 15 10422 17
rect 10426 15 10446 17
rect 9882 -25 9968 -17
rect 10000 -25 10086 -17
rect 9908 -41 9942 -25
rect 10026 -41 10060 -25
rect 9882 -61 9908 -55
rect 9946 -61 9968 -55
rect 10000 -61 10022 -55
rect 10064 -61 10086 -55
rect 9904 -79 9908 -61
rect 10128 -79 10132 0
rect 10316 -55 10320 0
rect 10364 -17 10446 15
rect 10447 -17 10456 17
rect 10464 -17 10481 17
rect 10362 -25 10448 -17
rect 10489 -25 10491 25
rect 10498 -17 10532 17
rect 10549 -17 10566 17
rect 10591 -25 10593 25
rect 10650 -17 10667 17
rect 10675 -25 10677 25
rect 10768 17 10854 25
rect 11130 17 11216 25
rect 11248 17 11334 25
rect 11610 17 11696 25
rect 10684 -17 10718 17
rect 10735 -17 10752 17
rect 10760 -17 10769 17
rect 10770 15 10803 17
rect 10832 15 10852 17
rect 10770 -17 10852 15
rect 11132 15 11156 17
rect 11181 15 11190 17
rect 11194 15 11214 17
rect 10768 -25 10854 -17
rect 10388 -41 10422 -25
rect 10794 -41 10828 -25
rect 10362 -61 10388 -55
rect 10426 -61 10448 -55
rect 10768 -61 10790 -55
rect 10832 -61 10854 -55
rect 10384 -79 10388 -61
rect 10896 -79 10900 0
rect 11084 -55 11088 0
rect 11132 -17 11214 15
rect 11215 -17 11224 17
rect 11240 -17 11249 17
rect 11250 15 11283 17
rect 11312 15 11332 17
rect 11250 -17 11332 15
rect 11612 15 11636 17
rect 11661 15 11670 17
rect 11674 15 11694 17
rect 11130 -25 11216 -17
rect 11248 -25 11334 -17
rect 11156 -41 11190 -25
rect 11274 -41 11308 -25
rect 11130 -61 11156 -55
rect 11194 -61 11216 -55
rect 11248 -61 11270 -55
rect 11312 -61 11334 -55
rect 11152 -79 11156 -61
rect 11376 -79 11380 0
rect 11564 -55 11568 0
rect 11612 -17 11694 15
rect 11695 -17 11704 17
rect 11712 -17 11729 17
rect 11610 -25 11696 -17
rect 11737 -25 11739 25
rect 11746 -17 11780 17
rect 11797 -17 11814 17
rect 11839 -25 11841 25
rect 11898 -17 11915 17
rect 11923 -25 11925 25
rect 12016 17 12102 25
rect 12378 17 12464 25
rect 12496 17 12582 25
rect 12858 17 12944 25
rect 11932 -17 11966 17
rect 11983 -17 12000 17
rect 12008 -17 12017 17
rect 12018 15 12051 17
rect 12080 15 12100 17
rect 12018 -17 12100 15
rect 12380 15 12404 17
rect 12429 15 12438 17
rect 12442 15 12462 17
rect 12016 -25 12102 -17
rect 11636 -41 11670 -25
rect 12042 -41 12076 -25
rect 11610 -61 11636 -55
rect 11674 -61 11696 -55
rect 12016 -61 12038 -55
rect 12080 -61 12102 -55
rect 11632 -79 11636 -61
rect 12144 -79 12148 0
rect 12332 -55 12336 0
rect 12380 -17 12462 15
rect 12463 -17 12472 17
rect 12488 -17 12497 17
rect 12498 15 12531 17
rect 12560 15 12580 17
rect 12498 -17 12580 15
rect 12860 15 12884 17
rect 12909 15 12918 17
rect 12922 15 12942 17
rect 12378 -25 12464 -17
rect 12496 -25 12582 -17
rect 12404 -41 12438 -25
rect 12522 -41 12556 -25
rect 12378 -61 12404 -55
rect 12442 -61 12464 -55
rect 12496 -61 12518 -55
rect 12560 -61 12582 -55
rect 12400 -79 12404 -61
rect 12624 -79 12628 0
rect 12812 -55 12816 0
rect 12860 -17 12942 15
rect 12943 -17 12952 17
rect 12960 -17 12977 17
rect 12858 -25 12944 -17
rect 12985 -25 12987 25
rect 12994 -17 13028 17
rect 13045 -17 13062 17
rect 13087 -25 13089 25
rect 13146 -17 13163 17
rect 13171 -25 13173 25
rect 13264 17 13350 25
rect 13626 17 13712 25
rect 13744 17 13830 25
rect 14106 17 14192 25
rect 13180 -17 13214 17
rect 13231 -17 13248 17
rect 13256 -17 13265 17
rect 13266 15 13299 17
rect 13328 15 13348 17
rect 13266 -17 13348 15
rect 13628 15 13652 17
rect 13677 15 13686 17
rect 13690 15 13710 17
rect 13264 -25 13350 -17
rect 12884 -41 12918 -25
rect 13290 -41 13324 -25
rect 12858 -61 12884 -55
rect 12922 -61 12944 -55
rect 13264 -61 13286 -55
rect 13328 -61 13350 -55
rect 12880 -79 12884 -61
rect 13392 -79 13396 0
rect 13580 -55 13584 0
rect 13628 -17 13710 15
rect 13711 -17 13720 17
rect 13736 -17 13745 17
rect 13746 15 13779 17
rect 13808 15 13828 17
rect 13746 -17 13828 15
rect 14108 15 14132 17
rect 14157 15 14166 17
rect 14170 15 14190 17
rect 13626 -25 13712 -17
rect 13744 -25 13830 -17
rect 13652 -41 13686 -25
rect 13770 -41 13804 -25
rect 13626 -61 13652 -55
rect 13690 -61 13712 -55
rect 13744 -61 13766 -55
rect 13808 -61 13830 -55
rect 13648 -79 13652 -61
rect 13872 -79 13876 0
rect 14060 -55 14064 0
rect 14108 -17 14190 15
rect 14191 -17 14200 17
rect 14208 -17 14225 17
rect 14106 -25 14192 -17
rect 14233 -25 14235 25
rect 14242 -17 14276 17
rect 14293 -17 14310 17
rect 14335 -25 14337 25
rect 14394 -17 14411 17
rect 14419 -25 14421 25
rect 14512 17 14598 25
rect 14874 17 14960 25
rect 14992 17 15078 25
rect 15354 17 15440 25
rect 14428 -17 14462 17
rect 14479 -17 14496 17
rect 14504 -17 14513 17
rect 14514 15 14547 17
rect 14576 15 14596 17
rect 14514 -17 14596 15
rect 14876 15 14900 17
rect 14925 15 14934 17
rect 14938 15 14958 17
rect 14512 -25 14598 -17
rect 14132 -41 14166 -25
rect 14538 -41 14572 -25
rect 14106 -61 14132 -55
rect 14170 -61 14192 -55
rect 14512 -61 14534 -55
rect 14576 -61 14598 -55
rect 14128 -79 14132 -61
rect 14640 -79 14644 0
rect 14828 -55 14832 0
rect 14876 -17 14958 15
rect 14959 -17 14968 17
rect 14984 -17 14993 17
rect 14994 15 15027 17
rect 15056 15 15076 17
rect 14994 -17 15076 15
rect 15356 15 15380 17
rect 15405 15 15414 17
rect 15418 15 15438 17
rect 14874 -25 14960 -17
rect 14992 -25 15078 -17
rect 14900 -41 14934 -25
rect 15018 -41 15052 -25
rect 14874 -61 14900 -55
rect 14938 -61 14960 -55
rect 14992 -61 15014 -55
rect 15056 -61 15078 -55
rect 14896 -79 14900 -61
rect 15120 -79 15124 0
rect 15308 -55 15312 0
rect 15356 -17 15438 15
rect 15439 -17 15448 17
rect 15456 -17 15473 17
rect 15354 -25 15440 -17
rect 15481 -25 15483 25
rect 15490 -17 15524 17
rect 15541 -17 15558 17
rect 15583 -25 15585 25
rect 15642 -17 15659 17
rect 15667 -25 15669 25
rect 15760 17 15846 25
rect 16122 17 16208 25
rect 16240 17 16326 25
rect 16602 17 16688 25
rect 15676 -17 15710 17
rect 15727 -17 15744 17
rect 15752 -17 15761 17
rect 15762 15 15795 17
rect 15824 15 15844 17
rect 15762 -17 15844 15
rect 16124 15 16148 17
rect 16173 15 16182 17
rect 16186 15 16206 17
rect 15760 -25 15846 -17
rect 15380 -41 15414 -25
rect 15786 -41 15820 -25
rect 15354 -61 15380 -55
rect 15418 -61 15440 -55
rect 15760 -61 15782 -55
rect 15824 -61 15846 -55
rect 15376 -79 15380 -61
rect 15888 -79 15892 0
rect 16076 -55 16080 0
rect 16124 -17 16206 15
rect 16207 -17 16216 17
rect 16232 -17 16241 17
rect 16242 15 16275 17
rect 16304 15 16324 17
rect 16242 -17 16324 15
rect 16604 15 16628 17
rect 16653 15 16662 17
rect 16666 15 16686 17
rect 16122 -25 16208 -17
rect 16240 -25 16326 -17
rect 16148 -41 16182 -25
rect 16266 -41 16300 -25
rect 16122 -61 16148 -55
rect 16186 -61 16208 -55
rect 16240 -61 16262 -55
rect 16304 -61 16326 -55
rect 16144 -79 16148 -61
rect 16368 -79 16372 0
rect 16556 -55 16560 0
rect 16604 -17 16686 15
rect 16687 -17 16696 17
rect 16704 -17 16721 17
rect 16602 -25 16688 -17
rect 16729 -25 16731 25
rect 16738 -17 16772 17
rect 16789 -17 16806 17
rect 16831 -25 16833 25
rect 16890 -17 16907 17
rect 16915 -25 16917 25
rect 17008 17 17094 25
rect 17370 17 17456 25
rect 17488 17 17574 25
rect 17850 17 17936 25
rect 16924 -17 16958 17
rect 16975 -17 16992 17
rect 17000 -17 17009 17
rect 17010 15 17043 17
rect 17072 15 17092 17
rect 17010 -17 17092 15
rect 17372 15 17396 17
rect 17421 15 17430 17
rect 17434 15 17454 17
rect 17008 -25 17094 -17
rect 16628 -41 16662 -25
rect 17034 -41 17068 -25
rect 16602 -61 16628 -55
rect 16666 -61 16688 -55
rect 17008 -61 17030 -55
rect 17072 -61 17094 -55
rect 16624 -79 16628 -61
rect 17136 -79 17140 0
rect 17324 -55 17328 0
rect 17372 -17 17454 15
rect 17455 -17 17464 17
rect 17480 -17 17489 17
rect 17490 15 17523 17
rect 17552 15 17572 17
rect 17490 -17 17572 15
rect 17852 15 17876 17
rect 17901 15 17910 17
rect 17914 15 17934 17
rect 17370 -25 17456 -17
rect 17488 -25 17574 -17
rect 17396 -41 17430 -25
rect 17514 -41 17548 -25
rect 17370 -61 17396 -55
rect 17434 -61 17456 -55
rect 17488 -61 17510 -55
rect 17552 -61 17574 -55
rect 17392 -79 17396 -61
rect 17616 -79 17620 0
rect 17804 -55 17808 0
rect 17852 -17 17934 15
rect 17935 -17 17944 17
rect 17952 -17 17969 17
rect 17850 -25 17936 -17
rect 17977 -25 17979 25
rect 17986 -17 18020 17
rect 18037 -17 18054 17
rect 18079 -25 18081 25
rect 18138 -17 18155 17
rect 18163 -25 18165 25
rect 18256 17 18342 25
rect 18618 17 18704 25
rect 18736 17 18822 25
rect 19098 17 19184 25
rect 18172 -17 18206 17
rect 18223 -17 18240 17
rect 18248 -17 18257 17
rect 18258 15 18291 17
rect 18320 15 18340 17
rect 18258 -17 18340 15
rect 18620 15 18644 17
rect 18669 15 18678 17
rect 18682 15 18702 17
rect 18256 -25 18342 -17
rect 17876 -41 17910 -25
rect 18282 -41 18316 -25
rect 17850 -61 17876 -55
rect 17914 -61 17936 -55
rect 18256 -61 18278 -55
rect 18320 -61 18342 -55
rect 17872 -79 17876 -61
rect 18384 -79 18388 0
rect 18572 -55 18576 0
rect 18620 -17 18702 15
rect 18703 -17 18712 17
rect 18728 -17 18737 17
rect 18738 15 18771 17
rect 18800 15 18820 17
rect 18738 -17 18820 15
rect 19100 15 19124 17
rect 19149 15 19158 17
rect 19162 15 19182 17
rect 18618 -25 18704 -17
rect 18736 -25 18822 -17
rect 18644 -41 18678 -25
rect 18762 -41 18796 -25
rect 18618 -61 18644 -55
rect 18682 -61 18704 -55
rect 18736 -61 18758 -55
rect 18800 -61 18822 -55
rect 18640 -79 18644 -61
rect 18864 -79 18868 0
rect 19052 -55 19056 0
rect 19100 -17 19182 15
rect 19183 -17 19192 17
rect 19200 -17 19217 17
rect 19098 -25 19184 -17
rect 19225 -25 19227 25
rect 19234 -17 19268 17
rect 19285 -17 19302 17
rect 19327 -25 19329 25
rect 19386 -17 19403 17
rect 19411 -25 19413 25
rect 19504 17 19590 25
rect 19866 17 19952 25
rect 19984 17 20070 25
rect 20346 17 20432 25
rect 19420 -17 19454 17
rect 19471 -17 19488 17
rect 19496 -17 19505 17
rect 19506 15 19539 17
rect 19568 15 19588 17
rect 19506 -17 19588 15
rect 19868 15 19892 17
rect 19917 15 19926 17
rect 19930 15 19950 17
rect 19504 -25 19590 -17
rect 19124 -41 19158 -25
rect 19530 -41 19564 -25
rect 19098 -61 19124 -55
rect 19162 -61 19184 -55
rect 19504 -61 19526 -55
rect 19568 -61 19590 -55
rect 19120 -79 19124 -61
rect 19632 -79 19636 0
rect 19820 -55 19824 0
rect 19868 -17 19950 15
rect 19951 -17 19960 17
rect 19976 -17 19985 17
rect 19986 15 20019 17
rect 20048 15 20068 17
rect 19986 -17 20068 15
rect 20348 15 20372 17
rect 20397 15 20406 17
rect 20410 15 20430 17
rect 19866 -25 19952 -17
rect 19984 -25 20070 -17
rect 19892 -41 19926 -25
rect 20010 -41 20044 -25
rect 19866 -61 19892 -55
rect 19930 -61 19952 -55
rect 19984 -61 20006 -55
rect 20048 -61 20070 -55
rect 19888 -79 19892 -61
rect 20112 -79 20116 0
rect 20300 -55 20304 0
rect 20348 -17 20430 15
rect 20431 -17 20440 17
rect 20448 -17 20465 17
rect 20346 -25 20432 -17
rect 20473 -25 20475 25
rect 20482 -17 20516 17
rect 20533 -17 20550 17
rect 20575 -25 20577 25
rect 20634 -17 20651 17
rect 20659 -25 20661 25
rect 20752 17 20838 25
rect 21114 17 21200 25
rect 21232 17 21318 25
rect 21594 17 21680 25
rect 20668 -17 20702 17
rect 20719 -17 20736 17
rect 20744 -17 20753 17
rect 20754 15 20787 17
rect 20816 15 20836 17
rect 20754 -17 20836 15
rect 21116 15 21140 17
rect 21165 15 21174 17
rect 21178 15 21198 17
rect 20752 -25 20838 -17
rect 20372 -41 20406 -25
rect 20778 -41 20812 -25
rect 20346 -61 20372 -55
rect 20410 -61 20432 -55
rect 20752 -61 20774 -55
rect 20816 -61 20838 -55
rect 20368 -79 20372 -61
rect 20880 -79 20884 0
rect 21068 -55 21072 0
rect 21116 -17 21198 15
rect 21199 -17 21208 17
rect 21224 -17 21233 17
rect 21234 15 21267 17
rect 21296 15 21316 17
rect 21234 -17 21316 15
rect 21596 15 21620 17
rect 21645 15 21654 17
rect 21658 15 21678 17
rect 21114 -25 21200 -17
rect 21232 -25 21318 -17
rect 21140 -41 21174 -25
rect 21258 -41 21292 -25
rect 21114 -61 21140 -55
rect 21178 -61 21200 -55
rect 21232 -61 21254 -55
rect 21296 -61 21318 -55
rect 21136 -79 21140 -61
rect 21360 -79 21364 0
rect 21548 -55 21552 0
rect 21596 -17 21678 15
rect 21679 -17 21688 17
rect 21696 -17 21713 17
rect 21594 -25 21680 -17
rect 21721 -25 21723 25
rect 21730 -17 21764 17
rect 21781 -17 21798 17
rect 21823 -25 21825 25
rect 21882 -17 21899 17
rect 21907 -25 21909 25
rect 22000 17 22086 25
rect 22362 17 22448 25
rect 22480 17 22566 25
rect 22842 17 22928 25
rect 21916 -17 21950 17
rect 21967 -17 21984 17
rect 21992 -17 22001 17
rect 22002 15 22035 17
rect 22064 15 22084 17
rect 22002 -17 22084 15
rect 22364 15 22388 17
rect 22413 15 22422 17
rect 22426 15 22446 17
rect 22000 -25 22086 -17
rect 21620 -41 21654 -25
rect 22026 -41 22060 -25
rect 21594 -61 21620 -55
rect 21658 -61 21680 -55
rect 22000 -61 22022 -55
rect 22064 -61 22086 -55
rect 21616 -79 21620 -61
rect 22128 -79 22132 0
rect 22316 -55 22320 0
rect 22364 -17 22446 15
rect 22447 -17 22456 17
rect 22472 -17 22481 17
rect 22482 15 22515 17
rect 22544 15 22564 17
rect 22482 -17 22564 15
rect 22844 15 22868 17
rect 22893 15 22902 17
rect 22906 15 22926 17
rect 22362 -25 22448 -17
rect 22480 -25 22566 -17
rect 22388 -41 22422 -25
rect 22506 -41 22540 -25
rect 22362 -61 22388 -55
rect 22426 -61 22448 -55
rect 22480 -61 22502 -55
rect 22544 -61 22566 -55
rect 22384 -79 22388 -61
rect 22608 -79 22612 0
rect 22796 -55 22800 0
rect 22844 -17 22926 15
rect 22927 -17 22936 17
rect 22944 -17 22961 17
rect 22842 -25 22928 -17
rect 22969 -25 22971 25
rect 22978 -17 23012 17
rect 23029 -17 23046 17
rect 23071 -25 23073 25
rect 23130 -17 23147 17
rect 23155 -25 23157 25
rect 23248 17 23334 25
rect 23610 17 23696 25
rect 23728 17 23814 25
rect 24090 17 24176 25
rect 23164 -17 23198 17
rect 23215 -17 23232 17
rect 23240 -17 23249 17
rect 23250 15 23283 17
rect 23312 15 23332 17
rect 23250 -17 23332 15
rect 23612 15 23636 17
rect 23661 15 23670 17
rect 23674 15 23694 17
rect 23248 -25 23334 -17
rect 22868 -41 22902 -25
rect 23274 -41 23308 -25
rect 22842 -61 22868 -55
rect 22906 -61 22928 -55
rect 23248 -61 23270 -55
rect 23312 -61 23334 -55
rect 22864 -79 22868 -61
rect 23376 -79 23380 0
rect 23564 -55 23568 0
rect 23612 -17 23694 15
rect 23695 -17 23704 17
rect 23720 -17 23729 17
rect 23730 15 23763 17
rect 23792 15 23812 17
rect 23730 -17 23812 15
rect 24092 15 24116 17
rect 24141 15 24150 17
rect 24154 15 24174 17
rect 23610 -25 23696 -17
rect 23728 -25 23814 -17
rect 23636 -41 23670 -25
rect 23754 -41 23788 -25
rect 23610 -61 23636 -55
rect 23674 -61 23696 -55
rect 23728 -61 23750 -55
rect 23792 -61 23814 -55
rect 23632 -79 23636 -61
rect 23856 -79 23860 0
rect 24044 -55 24048 0
rect 24092 -17 24174 15
rect 24175 -17 24184 17
rect 24192 -17 24209 17
rect 24090 -25 24176 -17
rect 24217 -25 24219 25
rect 24226 -17 24260 17
rect 24277 -17 24294 17
rect 24319 -25 24321 25
rect 24378 -17 24395 17
rect 24403 -25 24405 25
rect 24496 17 24582 25
rect 24858 17 24944 25
rect 24976 17 25062 25
rect 25338 17 25424 25
rect 24412 -17 24446 17
rect 24463 -17 24480 17
rect 24488 -17 24497 17
rect 24498 15 24531 17
rect 24560 15 24580 17
rect 24498 -17 24580 15
rect 24860 15 24884 17
rect 24909 15 24918 17
rect 24922 15 24942 17
rect 24496 -25 24582 -17
rect 24116 -41 24150 -25
rect 24522 -41 24556 -25
rect 24090 -61 24116 -55
rect 24154 -61 24176 -55
rect 24496 -61 24518 -55
rect 24560 -61 24582 -55
rect 24112 -79 24116 -61
rect 24624 -79 24628 0
rect 24812 -55 24816 0
rect 24860 -17 24942 15
rect 24943 -17 24952 17
rect 24968 -17 24977 17
rect 24978 15 25011 17
rect 25040 15 25060 17
rect 24978 -17 25060 15
rect 25340 15 25364 17
rect 25389 15 25398 17
rect 25402 15 25422 17
rect 24858 -25 24944 -17
rect 24976 -25 25062 -17
rect 24884 -41 24918 -25
rect 25002 -41 25036 -25
rect 24858 -61 24884 -55
rect 24922 -61 24944 -55
rect 24976 -61 24998 -55
rect 25040 -61 25062 -55
rect 24880 -79 24884 -61
rect 25104 -79 25108 0
rect 25292 -55 25296 0
rect 25340 -17 25422 15
rect 25423 -17 25432 17
rect 25440 -17 25457 17
rect 25338 -25 25424 -17
rect 25465 -25 25467 25
rect 25474 -17 25508 17
rect 25525 -17 25542 17
rect 25567 -25 25569 25
rect 25626 -17 25643 17
rect 25651 -25 25653 25
rect 25744 17 25830 25
rect 26106 17 26192 25
rect 26224 17 26310 25
rect 26586 17 26672 25
rect 25660 -17 25694 17
rect 25711 -17 25728 17
rect 25736 -17 25745 17
rect 25746 15 25779 17
rect 25808 15 25828 17
rect 25746 -17 25828 15
rect 26108 15 26132 17
rect 26157 15 26166 17
rect 26170 15 26190 17
rect 25744 -25 25830 -17
rect 25364 -41 25398 -25
rect 25770 -41 25804 -25
rect 25338 -61 25364 -55
rect 25402 -61 25424 -55
rect 25744 -61 25766 -55
rect 25808 -61 25830 -55
rect 25360 -79 25364 -61
rect 25872 -79 25876 0
rect 26060 -55 26064 0
rect 26108 -17 26190 15
rect 26191 -17 26200 17
rect 26216 -17 26225 17
rect 26226 15 26259 17
rect 26288 15 26308 17
rect 26226 -17 26308 15
rect 26588 15 26612 17
rect 26637 15 26646 17
rect 26650 15 26670 17
rect 26106 -25 26192 -17
rect 26224 -25 26310 -17
rect 26132 -41 26166 -25
rect 26250 -41 26284 -25
rect 26106 -61 26132 -55
rect 26170 -61 26192 -55
rect 26224 -61 26246 -55
rect 26288 -61 26310 -55
rect 26128 -79 26132 -61
rect 26352 -79 26356 0
rect 26540 -55 26544 0
rect 26588 -17 26670 15
rect 26671 -17 26680 17
rect 26688 -17 26705 17
rect 26586 -25 26672 -17
rect 26713 -25 26715 25
rect 26722 -17 26756 17
rect 26773 -17 26790 17
rect 26815 -25 26817 25
rect 26874 -17 26891 17
rect 26899 -25 26901 25
rect 26992 17 27078 25
rect 27354 17 27440 25
rect 27472 17 27558 25
rect 27834 17 27920 25
rect 26908 -17 26942 17
rect 26959 -17 26976 17
rect 26984 -17 26993 17
rect 26994 15 27027 17
rect 27056 15 27076 17
rect 26994 -17 27076 15
rect 27356 15 27380 17
rect 27405 15 27414 17
rect 27418 15 27438 17
rect 26992 -25 27078 -17
rect 26612 -41 26646 -25
rect 27018 -41 27052 -25
rect 26586 -61 26612 -55
rect 26650 -61 26672 -55
rect 26992 -61 27014 -55
rect 27056 -61 27078 -55
rect 26608 -79 26612 -61
rect 27120 -79 27124 0
rect 27308 -55 27312 0
rect 27356 -17 27438 15
rect 27439 -17 27448 17
rect 27464 -17 27473 17
rect 27474 15 27507 17
rect 27536 15 27556 17
rect 27474 -17 27556 15
rect 27836 15 27860 17
rect 27885 15 27894 17
rect 27898 15 27918 17
rect 27354 -25 27440 -17
rect 27472 -25 27558 -17
rect 27380 -41 27414 -25
rect 27498 -41 27532 -25
rect 27354 -61 27380 -55
rect 27418 -61 27440 -55
rect 27472 -61 27494 -55
rect 27536 -61 27558 -55
rect 27376 -79 27380 -61
rect 27600 -79 27604 0
rect 27788 -55 27792 0
rect 27836 -17 27918 15
rect 27919 -17 27928 17
rect 27936 -17 27953 17
rect 27834 -25 27920 -17
rect 27961 -25 27963 25
rect 27970 -17 28004 17
rect 28021 -17 28038 17
rect 28063 -25 28065 25
rect 28122 -17 28139 17
rect 28147 -25 28149 25
rect 28240 17 28326 25
rect 28602 17 28688 25
rect 28720 17 28806 25
rect 29082 17 29168 25
rect 28156 -17 28190 17
rect 28207 -17 28224 17
rect 28232 -17 28241 17
rect 28242 15 28275 17
rect 28304 15 28324 17
rect 28242 -17 28324 15
rect 28604 15 28628 17
rect 28653 15 28662 17
rect 28666 15 28686 17
rect 28240 -25 28326 -17
rect 27860 -41 27894 -25
rect 28266 -41 28300 -25
rect 27834 -61 27860 -55
rect 27898 -61 27920 -55
rect 28240 -61 28262 -55
rect 28304 -61 28326 -55
rect 27856 -79 27860 -61
rect 28368 -79 28372 0
rect 28556 -55 28560 0
rect 28604 -17 28686 15
rect 28687 -17 28696 17
rect 28712 -17 28721 17
rect 28722 15 28755 17
rect 28784 15 28804 17
rect 28722 -17 28804 15
rect 29084 15 29108 17
rect 29133 15 29142 17
rect 29146 15 29166 17
rect 28602 -25 28688 -17
rect 28720 -25 28806 -17
rect 28628 -41 28662 -25
rect 28746 -41 28780 -25
rect 28602 -61 28628 -55
rect 28666 -61 28688 -55
rect 28720 -61 28742 -55
rect 28784 -61 28806 -55
rect 28624 -79 28628 -61
rect 28848 -79 28852 0
rect 29036 -55 29040 0
rect 29084 -17 29166 15
rect 29167 -17 29176 17
rect 29184 -17 29201 17
rect 29082 -25 29168 -17
rect 29209 -25 29211 25
rect 29218 -17 29252 17
rect 29269 -17 29286 17
rect 29311 -25 29313 25
rect 29370 -17 29387 17
rect 29395 -25 29397 25
rect 29488 17 29574 25
rect 29850 17 29936 25
rect 29968 17 30054 25
rect 30330 17 30416 25
rect 29404 -17 29438 17
rect 29455 -17 29472 17
rect 29480 -17 29489 17
rect 29490 15 29523 17
rect 29552 15 29572 17
rect 29490 -17 29572 15
rect 29852 15 29876 17
rect 29901 15 29910 17
rect 29914 15 29934 17
rect 29488 -25 29574 -17
rect 29108 -41 29142 -25
rect 29514 -41 29548 -25
rect 29082 -61 29108 -55
rect 29146 -61 29168 -55
rect 29488 -61 29510 -55
rect 29552 -61 29574 -55
rect 29104 -79 29108 -61
rect 29616 -79 29620 0
rect 29804 -55 29808 0
rect 29852 -17 29934 15
rect 29935 -17 29944 17
rect 29960 -17 29969 17
rect 29970 15 30003 17
rect 30032 15 30052 17
rect 29970 -17 30052 15
rect 30332 15 30356 17
rect 30381 15 30390 17
rect 30394 15 30414 17
rect 29850 -25 29936 -17
rect 29968 -25 30054 -17
rect 29876 -41 29910 -25
rect 29994 -41 30028 -25
rect 29850 -61 29876 -55
rect 29914 -61 29936 -55
rect 29968 -61 29990 -55
rect 30032 -61 30054 -55
rect 29872 -79 29876 -61
rect 30096 -79 30100 0
rect 30284 -55 30288 0
rect 30332 -17 30414 15
rect 30415 -17 30424 17
rect 30432 -17 30449 17
rect 30330 -25 30416 -17
rect 30457 -25 30459 25
rect 30466 -17 30500 17
rect 30517 -17 30534 17
rect 30559 -25 30561 25
rect 30618 -17 30635 17
rect 30643 -25 30645 25
rect 30736 17 30822 25
rect 31098 17 31184 25
rect 31216 17 31302 25
rect 31578 17 31664 25
rect 30652 -17 30686 17
rect 30703 -17 30720 17
rect 30728 -17 30737 17
rect 30738 15 30771 17
rect 30800 15 30820 17
rect 30738 -17 30820 15
rect 31100 15 31124 17
rect 31149 15 31158 17
rect 31162 15 31182 17
rect 30736 -25 30822 -17
rect 30356 -41 30390 -25
rect 30762 -41 30796 -25
rect 30330 -61 30356 -55
rect 30394 -61 30416 -55
rect 30736 -61 30758 -55
rect 30800 -61 30822 -55
rect 30352 -79 30356 -61
rect 30864 -79 30868 0
rect 31052 -55 31056 0
rect 31100 -17 31182 15
rect 31183 -17 31192 17
rect 31208 -17 31217 17
rect 31218 15 31251 17
rect 31280 15 31300 17
rect 31218 -17 31300 15
rect 31580 15 31604 17
rect 31629 15 31638 17
rect 31642 15 31662 17
rect 31098 -25 31184 -17
rect 31216 -25 31302 -17
rect 31124 -41 31158 -25
rect 31242 -41 31276 -25
rect 31098 -61 31124 -55
rect 31162 -61 31184 -55
rect 31216 -61 31238 -55
rect 31280 -61 31302 -55
rect 31120 -79 31124 -61
rect 31344 -79 31348 0
rect 31532 -55 31536 0
rect 31580 -17 31662 15
rect 31663 -17 31672 17
rect 31680 -17 31697 17
rect 31578 -25 31664 -17
rect 31705 -25 31707 25
rect 31714 -17 31748 17
rect 31765 -17 31782 17
rect 31807 -25 31809 25
rect 31866 -17 31883 17
rect 31891 -25 31893 25
rect 31984 17 32070 25
rect 32346 17 32432 25
rect 32464 17 32550 25
rect 32826 17 32912 25
rect 31900 -17 31934 17
rect 31951 -17 31968 17
rect 31976 -17 31985 17
rect 31986 15 32019 17
rect 32048 15 32068 17
rect 31986 -17 32068 15
rect 32348 15 32372 17
rect 32397 15 32406 17
rect 32410 15 32430 17
rect 31984 -25 32070 -17
rect 31604 -41 31638 -25
rect 32010 -41 32044 -25
rect 31578 -61 31604 -55
rect 31642 -61 31664 -55
rect 31984 -61 32006 -55
rect 32048 -61 32070 -55
rect 31600 -79 31604 -61
rect 32112 -79 32116 0
rect 32300 -55 32304 0
rect 32348 -17 32430 15
rect 32431 -17 32440 17
rect 32456 -17 32465 17
rect 32466 15 32499 17
rect 32528 15 32548 17
rect 32466 -17 32548 15
rect 32828 15 32852 17
rect 32877 15 32886 17
rect 32890 15 32910 17
rect 32346 -25 32432 -17
rect 32464 -25 32550 -17
rect 32372 -41 32406 -25
rect 32490 -41 32524 -25
rect 32346 -61 32372 -55
rect 32410 -61 32432 -55
rect 32464 -61 32486 -55
rect 32528 -61 32550 -55
rect 32368 -79 32372 -61
rect 32592 -79 32596 0
rect 32780 -55 32784 0
rect 32828 -17 32910 15
rect 32911 -17 32920 17
rect 32928 -17 32945 17
rect 32826 -25 32912 -17
rect 32953 -25 32955 25
rect 32962 -17 32996 17
rect 33013 -17 33030 17
rect 33055 -25 33057 25
rect 33114 -17 33131 17
rect 33139 -25 33141 25
rect 33232 17 33318 25
rect 33594 17 33680 25
rect 33712 17 33798 25
rect 34074 17 34160 25
rect 33148 -17 33182 17
rect 33199 -17 33216 17
rect 33224 -17 33233 17
rect 33234 15 33267 17
rect 33296 15 33316 17
rect 33234 -17 33316 15
rect 33596 15 33620 17
rect 33645 15 33654 17
rect 33658 15 33678 17
rect 33232 -25 33318 -17
rect 32852 -41 32886 -25
rect 33258 -41 33292 -25
rect 32826 -61 32852 -55
rect 32890 -61 32912 -55
rect 33232 -61 33254 -55
rect 33296 -61 33318 -55
rect 32848 -79 32852 -61
rect 33360 -79 33364 0
rect 33548 -55 33552 0
rect 33596 -17 33678 15
rect 33679 -17 33688 17
rect 33704 -17 33713 17
rect 33714 15 33747 17
rect 33776 15 33796 17
rect 33714 -17 33796 15
rect 34076 15 34100 17
rect 34125 15 34134 17
rect 34138 15 34158 17
rect 33594 -25 33680 -17
rect 33712 -25 33798 -17
rect 33620 -41 33654 -25
rect 33738 -41 33772 -25
rect 33594 -61 33620 -55
rect 33658 -61 33680 -55
rect 33712 -61 33734 -55
rect 33776 -61 33798 -55
rect 33616 -79 33620 -61
rect 33840 -79 33844 0
rect 34028 -55 34032 0
rect 34076 -17 34158 15
rect 34159 -17 34168 17
rect 34176 -17 34193 17
rect 34074 -25 34160 -17
rect 34201 -25 34203 25
rect 34210 -17 34244 17
rect 34261 -17 34278 17
rect 34303 -25 34305 25
rect 34362 -17 34379 17
rect 34387 -25 34389 25
rect 34480 17 34566 25
rect 34842 17 34928 25
rect 34960 17 35046 25
rect 35322 17 35408 25
rect 34396 -17 34430 17
rect 34447 -17 34464 17
rect 34472 -17 34481 17
rect 34482 15 34515 17
rect 34544 15 34564 17
rect 34482 -17 34564 15
rect 34844 15 34868 17
rect 34893 15 34902 17
rect 34906 15 34926 17
rect 34480 -25 34566 -17
rect 34100 -41 34134 -25
rect 34506 -41 34540 -25
rect 34074 -61 34100 -55
rect 34138 -61 34160 -55
rect 34480 -61 34502 -55
rect 34544 -61 34566 -55
rect 34096 -79 34100 -61
rect 34608 -79 34612 0
rect 34796 -55 34800 0
rect 34844 -17 34926 15
rect 34927 -17 34936 17
rect 34952 -17 34961 17
rect 34962 15 34995 17
rect 35024 15 35044 17
rect 34962 -17 35044 15
rect 35324 15 35348 17
rect 35373 15 35382 17
rect 35386 15 35406 17
rect 34842 -25 34928 -17
rect 34960 -25 35046 -17
rect 34868 -41 34902 -25
rect 34986 -41 35020 -25
rect 34842 -61 34868 -55
rect 34906 -61 34928 -55
rect 34960 -61 34982 -55
rect 35024 -61 35046 -55
rect 34864 -79 34868 -61
rect 35088 -79 35092 0
rect 35276 -55 35280 0
rect 35324 -17 35406 15
rect 35407 -17 35416 17
rect 35424 -17 35441 17
rect 35322 -25 35408 -17
rect 35449 -25 35451 25
rect 35458 -17 35492 17
rect 35509 -17 35526 17
rect 35551 -25 35553 25
rect 35610 -17 35627 17
rect 35635 -25 35637 25
rect 35728 17 35814 25
rect 36090 17 36176 25
rect 36208 17 36294 25
rect 36570 17 36656 25
rect 35644 -17 35678 17
rect 35695 -17 35712 17
rect 35720 -17 35729 17
rect 35730 15 35763 17
rect 35792 15 35812 17
rect 35730 -17 35812 15
rect 36092 15 36116 17
rect 36141 15 36150 17
rect 36154 15 36174 17
rect 35728 -25 35814 -17
rect 35348 -41 35382 -25
rect 35754 -41 35788 -25
rect 35322 -61 35348 -55
rect 35386 -61 35408 -55
rect 35728 -61 35750 -55
rect 35792 -61 35814 -55
rect 35344 -79 35348 -61
rect 35856 -79 35860 0
rect 36044 -55 36048 0
rect 36092 -17 36174 15
rect 36175 -17 36184 17
rect 36200 -17 36209 17
rect 36210 15 36243 17
rect 36272 15 36292 17
rect 36210 -17 36292 15
rect 36572 15 36596 17
rect 36621 15 36630 17
rect 36634 15 36654 17
rect 36090 -25 36176 -17
rect 36208 -25 36294 -17
rect 36116 -41 36150 -25
rect 36234 -41 36268 -25
rect 36090 -61 36116 -55
rect 36154 -61 36176 -55
rect 36208 -61 36230 -55
rect 36272 -61 36294 -55
rect 36112 -79 36116 -61
rect 36336 -79 36340 0
rect 36524 -55 36528 0
rect 36572 -17 36654 15
rect 36655 -17 36664 17
rect 36672 -17 36689 17
rect 36570 -25 36656 -17
rect 36697 -25 36699 25
rect 36706 -17 36740 17
rect 36757 -17 36774 17
rect 36799 -25 36801 25
rect 36858 -17 36875 17
rect 36883 -25 36885 25
rect 36976 17 37062 25
rect 37338 17 37424 25
rect 37456 17 37542 25
rect 37818 17 37904 25
rect 36892 -17 36926 17
rect 36943 -17 36960 17
rect 36968 -17 36977 17
rect 36978 15 37011 17
rect 37040 15 37060 17
rect 36978 -17 37060 15
rect 37340 15 37364 17
rect 37389 15 37398 17
rect 37402 15 37422 17
rect 36976 -25 37062 -17
rect 36596 -41 36630 -25
rect 37002 -41 37036 -25
rect 36570 -61 36596 -55
rect 36634 -61 36656 -55
rect 36976 -61 36998 -55
rect 37040 -61 37062 -55
rect 36592 -79 36596 -61
rect 37104 -79 37108 0
rect 37292 -55 37296 0
rect 37340 -17 37422 15
rect 37423 -17 37432 17
rect 37448 -17 37457 17
rect 37458 15 37491 17
rect 37520 15 37540 17
rect 37458 -17 37540 15
rect 37820 15 37844 17
rect 37869 15 37878 17
rect 37882 15 37902 17
rect 37338 -25 37424 -17
rect 37456 -25 37542 -17
rect 37364 -41 37398 -25
rect 37482 -41 37516 -25
rect 37338 -61 37364 -55
rect 37402 -61 37424 -55
rect 37456 -61 37478 -55
rect 37520 -61 37542 -55
rect 37360 -79 37364 -61
rect 37584 -79 37588 0
rect 37772 -55 37776 0
rect 37820 -17 37902 15
rect 37903 -17 37912 17
rect 37920 -17 37937 17
rect 37818 -25 37904 -17
rect 37945 -25 37947 25
rect 37954 -17 37988 17
rect 38005 -17 38022 17
rect 38047 -25 38049 25
rect 38106 -17 38123 17
rect 38131 -25 38133 25
rect 38224 17 38310 25
rect 38586 17 38672 25
rect 38704 17 38790 25
rect 39066 17 39152 25
rect 38140 -17 38174 17
rect 38191 -17 38208 17
rect 38216 -17 38225 17
rect 38226 15 38259 17
rect 38288 15 38308 17
rect 38226 -17 38308 15
rect 38588 15 38612 17
rect 38637 15 38646 17
rect 38650 15 38670 17
rect 38224 -25 38310 -17
rect 37844 -41 37878 -25
rect 38250 -41 38284 -25
rect 37818 -61 37844 -55
rect 37882 -61 37904 -55
rect 38224 -61 38246 -55
rect 38288 -61 38310 -55
rect 37840 -79 37844 -61
rect 38352 -79 38356 0
rect 38540 -55 38544 0
rect 38588 -17 38670 15
rect 38671 -17 38680 17
rect 38696 -17 38705 17
rect 38706 15 38739 17
rect 38768 15 38788 17
rect 38706 -17 38788 15
rect 39068 15 39092 17
rect 39117 15 39126 17
rect 39130 15 39150 17
rect 38586 -25 38672 -17
rect 38704 -25 38790 -17
rect 38612 -41 38646 -25
rect 38730 -41 38764 -25
rect 38586 -61 38612 -55
rect 38650 -61 38672 -55
rect 38704 -61 38726 -55
rect 38768 -61 38790 -55
rect 38608 -79 38612 -61
rect 38832 -79 38836 0
rect 39020 -55 39024 0
rect 39068 -17 39150 15
rect 39151 -17 39160 17
rect 39168 -17 39185 17
rect 39066 -25 39152 -17
rect 39193 -25 39195 25
rect 39202 -17 39236 17
rect 39253 -17 39270 17
rect 39295 -25 39297 25
rect 39354 -17 39371 17
rect 39379 -25 39381 25
rect 39472 17 39558 25
rect 39834 17 39920 25
rect 39952 17 40038 25
rect 40314 17 40400 25
rect 39388 -17 39422 17
rect 39439 -17 39456 17
rect 39464 -17 39473 17
rect 39474 15 39507 17
rect 39536 15 39556 17
rect 39474 -17 39556 15
rect 39836 15 39860 17
rect 39885 15 39894 17
rect 39898 15 39918 17
rect 39472 -25 39558 -17
rect 39092 -41 39126 -25
rect 39498 -41 39532 -25
rect 39066 -61 39092 -55
rect 39130 -61 39152 -55
rect 39472 -61 39494 -55
rect 39536 -61 39558 -55
rect 39088 -79 39092 -61
rect 39600 -79 39604 0
rect 39788 -55 39792 0
rect 39836 -17 39918 15
rect 39919 -17 39928 17
rect 39944 -17 39953 17
rect 39954 15 39987 17
rect 40016 15 40036 17
rect 39954 -17 40036 15
rect 40316 15 40340 17
rect 40365 15 40374 17
rect 40378 15 40398 17
rect 39834 -25 39920 -17
rect 39952 -25 40038 -17
rect 39860 -41 39894 -25
rect 39978 -41 40012 -25
rect 39834 -61 39860 -55
rect 39898 -61 39920 -55
rect 39952 -61 39974 -55
rect 40016 -61 40038 -55
rect 39856 -79 39860 -61
rect 40080 -79 40084 0
rect 40268 -55 40272 0
rect 40316 -17 40398 15
rect 40399 -17 40408 17
rect 40416 -17 40433 17
rect 40314 -25 40400 -17
rect 40441 -25 40443 25
rect 40450 -17 40484 17
rect 40501 -17 40518 17
rect 40543 -25 40545 25
rect 40602 -17 40619 17
rect 40627 -25 40629 25
rect 40720 17 40806 25
rect 41082 17 41168 25
rect 41200 17 41286 25
rect 41562 17 41648 25
rect 40636 -17 40670 17
rect 40687 -17 40704 17
rect 40712 -17 40721 17
rect 40722 15 40755 17
rect 40784 15 40804 17
rect 40722 -17 40804 15
rect 41084 15 41108 17
rect 41133 15 41142 17
rect 41146 15 41166 17
rect 40720 -25 40806 -17
rect 40340 -41 40374 -25
rect 40746 -41 40780 -25
rect 40320 -61 40340 -55
rect 40378 -61 40400 -55
rect 40720 -61 40742 -55
rect 40784 -61 40806 -55
rect 40336 -79 40340 -61
rect 40848 -79 40852 0
rect 41036 -55 41040 0
rect 41084 -17 41166 15
rect 41167 -17 41176 17
rect 41192 -17 41201 17
rect 41202 15 41235 17
rect 41264 15 41284 17
rect 41202 -17 41284 15
rect 41564 15 41588 17
rect 41613 15 41622 17
rect 41626 15 41646 17
rect 41082 -25 41168 -17
rect 41200 -25 41286 -17
rect 41108 -41 41142 -25
rect 41226 -41 41260 -25
rect 41082 -61 41108 -55
rect 41146 -61 41168 -55
rect 41200 -61 41222 -55
rect 41264 -61 41286 -55
rect 41104 -79 41108 -61
rect 41328 -79 41332 0
rect 41516 -55 41520 0
rect 41564 -17 41646 15
rect 41647 -17 41656 17
rect 41664 -17 41681 17
rect 41562 -25 41648 -17
rect 41689 -25 41691 25
rect 41698 -17 41732 17
rect 41749 -17 41766 17
rect 41791 -25 41793 25
rect 41850 -17 41867 17
rect 41875 -25 41877 25
rect 41968 17 42054 25
rect 42330 17 42416 25
rect 42448 17 42534 25
rect 42810 17 42896 25
rect 41884 -17 41918 17
rect 41935 -17 41952 17
rect 41960 -17 41969 17
rect 41970 15 42003 17
rect 42032 15 42052 17
rect 41970 -17 42052 15
rect 42332 15 42356 17
rect 42381 15 42390 17
rect 42394 15 42414 17
rect 41968 -25 42054 -17
rect 41588 -41 41622 -25
rect 41994 -41 42028 -25
rect 41562 -61 41588 -55
rect 41626 -61 41648 -55
rect 41968 -61 41990 -55
rect 42032 -61 42054 -55
rect 41584 -79 41588 -61
rect 42096 -79 42100 0
rect 42284 -55 42288 0
rect 42332 -17 42414 15
rect 42415 -17 42424 17
rect 42440 -17 42449 17
rect 42450 15 42483 17
rect 42512 15 42532 17
rect 42450 -17 42532 15
rect 42812 15 42836 17
rect 42861 15 42870 17
rect 42874 15 42894 17
rect 42330 -25 42416 -17
rect 42448 -25 42534 -17
rect 42356 -41 42390 -25
rect 42474 -41 42508 -25
rect 42330 -61 42356 -55
rect 42394 -61 42416 -55
rect 42448 -61 42470 -55
rect 42512 -61 42534 -55
rect 42352 -79 42356 -61
rect 42576 -79 42580 0
rect 42764 -55 42768 0
rect 42812 -17 42894 15
rect 42895 -17 42904 17
rect 42912 -17 42929 17
rect 42810 -25 42896 -17
rect 42937 -25 42939 25
rect 42946 -17 42980 17
rect 42997 -17 43014 17
rect 43039 -25 43041 25
rect 43098 -17 43115 17
rect 43123 -25 43125 25
rect 43216 17 43302 25
rect 43578 17 43664 25
rect 43696 17 43782 25
rect 44058 17 44144 25
rect 43132 -17 43166 17
rect 43183 -17 43200 17
rect 43208 -17 43217 17
rect 43218 15 43251 17
rect 43280 15 43300 17
rect 43218 -17 43300 15
rect 43580 15 43604 17
rect 43629 15 43638 17
rect 43642 15 43662 17
rect 43216 -25 43302 -17
rect 42836 -41 42870 -25
rect 43242 -41 43276 -25
rect 42810 -61 42836 -55
rect 42874 -61 42896 -55
rect 43216 -61 43238 -55
rect 43280 -61 43302 -55
rect 42832 -79 42836 -61
rect 43344 -79 43348 0
rect 43532 -55 43536 0
rect 43580 -17 43662 15
rect 43663 -17 43672 17
rect 43688 -17 43697 17
rect 43698 15 43731 17
rect 43760 15 43780 17
rect 43698 -17 43780 15
rect 44060 15 44084 17
rect 44109 15 44118 17
rect 44122 15 44142 17
rect 43578 -25 43664 -17
rect 43696 -25 43782 -17
rect 43604 -41 43638 -25
rect 43722 -41 43756 -25
rect 43578 -61 43604 -55
rect 43642 -61 43664 -55
rect 43696 -61 43718 -55
rect 43760 -61 43782 -55
rect 43600 -79 43604 -61
rect 43824 -79 43828 0
rect 44012 -55 44016 0
rect 44060 -17 44142 15
rect 44143 -17 44152 17
rect 44160 -17 44177 17
rect 44058 -25 44144 -17
rect 44185 -25 44187 25
rect 44194 -17 44228 17
rect 44245 -17 44262 17
rect 44287 -25 44289 25
rect 44346 -17 44363 17
rect 44371 -25 44373 25
rect 44464 17 44550 25
rect 44826 17 44912 25
rect 44944 17 45030 25
rect 45306 17 45392 25
rect 44380 -17 44414 17
rect 44431 -17 44448 17
rect 44456 -17 44465 17
rect 44466 15 44499 17
rect 44528 15 44548 17
rect 44466 -17 44548 15
rect 44828 15 44852 17
rect 44877 15 44886 17
rect 44890 15 44910 17
rect 44464 -25 44550 -17
rect 44084 -41 44118 -25
rect 44490 -41 44524 -25
rect 44058 -61 44084 -55
rect 44122 -61 44144 -55
rect 44464 -61 44486 -55
rect 44528 -61 44550 -55
rect 44080 -79 44084 -61
rect 44592 -79 44596 0
rect 44780 -55 44784 0
rect 44828 -17 44910 15
rect 44911 -17 44920 17
rect 44936 -17 44945 17
rect 44946 15 44979 17
rect 45008 15 45028 17
rect 44946 -17 45028 15
rect 45308 15 45332 17
rect 45357 15 45366 17
rect 45370 15 45390 17
rect 44826 -25 44912 -17
rect 44944 -25 45030 -17
rect 44852 -41 44886 -25
rect 44970 -41 45004 -25
rect 44826 -61 44852 -55
rect 44890 -61 44912 -55
rect 44944 -61 44966 -55
rect 45008 -61 45030 -55
rect 44848 -79 44852 -61
rect 45072 -79 45076 0
rect 45260 -55 45264 0
rect 45308 -17 45390 15
rect 45391 -17 45400 17
rect 45408 -17 45425 17
rect 45306 -25 45392 -17
rect 45433 -25 45435 25
rect 45442 -17 45476 17
rect 45493 -17 45510 17
rect 45535 -25 45537 25
rect 45594 -17 45611 17
rect 45619 -25 45621 25
rect 45712 17 45798 25
rect 46074 17 46160 25
rect 46192 17 46278 25
rect 46554 17 46640 25
rect 45628 -17 45662 17
rect 45679 -17 45696 17
rect 45704 -17 45713 17
rect 45714 15 45747 17
rect 45776 15 45796 17
rect 45714 -17 45796 15
rect 46076 15 46100 17
rect 46125 15 46134 17
rect 46138 15 46158 17
rect 45712 -25 45798 -17
rect 45332 -41 45366 -25
rect 45738 -41 45772 -25
rect 45306 -61 45332 -55
rect 45370 -61 45392 -55
rect 45712 -61 45734 -55
rect 45776 -61 45798 -55
rect 45328 -79 45332 -61
rect 45840 -79 45844 0
rect 46028 -55 46032 0
rect 46076 -17 46158 15
rect 46159 -17 46168 17
rect 46184 -17 46193 17
rect 46194 15 46227 17
rect 46256 15 46276 17
rect 46194 -17 46276 15
rect 46556 15 46580 17
rect 46605 15 46614 17
rect 46618 15 46638 17
rect 46074 -25 46160 -17
rect 46192 -25 46278 -17
rect 46100 -41 46134 -25
rect 46218 -41 46252 -25
rect 46074 -61 46100 -55
rect 46138 -61 46160 -55
rect 46192 -61 46214 -55
rect 46256 -61 46278 -55
rect 46096 -79 46100 -61
rect 46320 -79 46324 0
rect 46508 -55 46512 0
rect 46556 -17 46638 15
rect 46639 -17 46648 17
rect 46656 -17 46673 17
rect 46554 -25 46640 -17
rect 46681 -25 46683 25
rect 46690 -17 46724 17
rect 46741 -17 46758 17
rect 46783 -25 46785 25
rect 46842 -17 46859 17
rect 46867 -25 46869 25
rect 46960 17 47046 25
rect 47322 17 47408 25
rect 47440 17 47526 25
rect 47802 17 47888 25
rect 46876 -17 46910 17
rect 46927 -17 46944 17
rect 46952 -17 46961 17
rect 46962 15 46995 17
rect 47024 15 47044 17
rect 46962 -17 47044 15
rect 47324 15 47348 17
rect 47373 15 47382 17
rect 47386 15 47406 17
rect 46960 -25 47046 -17
rect 46580 -41 46614 -25
rect 46986 -41 47020 -25
rect 46554 -61 46580 -55
rect 46618 -61 46640 -55
rect 46960 -61 46982 -55
rect 47024 -61 47046 -55
rect 46576 -79 46580 -61
rect 47088 -79 47092 0
rect 47276 -55 47280 0
rect 47324 -17 47406 15
rect 47407 -17 47416 17
rect 47432 -17 47441 17
rect 47442 15 47475 17
rect 47504 15 47524 17
rect 47442 -17 47524 15
rect 47804 15 47828 17
rect 47853 15 47862 17
rect 47866 15 47886 17
rect 47322 -25 47408 -17
rect 47440 -25 47526 -17
rect 47348 -41 47382 -25
rect 47466 -41 47500 -25
rect 47322 -61 47348 -55
rect 47386 -61 47408 -55
rect 47440 -61 47462 -55
rect 47504 -61 47526 -55
rect 47344 -79 47348 -61
rect 47568 -79 47572 0
rect 47756 -55 47760 0
rect 47804 -17 47886 15
rect 47887 -17 47896 17
rect 47904 -17 47921 17
rect 47802 -25 47888 -17
rect 47929 -25 47931 25
rect 47938 -17 47972 17
rect 47989 -17 48006 17
rect 48031 -25 48033 25
rect 48090 -17 48107 17
rect 48115 -25 48117 25
rect 48208 17 48294 25
rect 48570 17 48656 25
rect 48688 17 48774 25
rect 49050 17 49136 25
rect 48124 -17 48158 17
rect 48175 -17 48192 17
rect 48200 -17 48209 17
rect 48210 15 48243 17
rect 48272 15 48292 17
rect 48210 -17 48292 15
rect 48572 15 48596 17
rect 48621 15 48630 17
rect 48634 15 48654 17
rect 48208 -25 48294 -17
rect 47828 -41 47862 -25
rect 48234 -41 48268 -25
rect 47802 -61 47828 -55
rect 47866 -61 47888 -55
rect 48208 -61 48230 -55
rect 48272 -61 48294 -55
rect 47824 -79 47828 -61
rect 48336 -79 48340 0
rect 48524 -55 48528 0
rect 48572 -17 48654 15
rect 48655 -17 48664 17
rect 48680 -17 48689 17
rect 48690 15 48723 17
rect 48752 15 48772 17
rect 48690 -17 48772 15
rect 49052 15 49076 17
rect 49101 15 49110 17
rect 49114 15 49134 17
rect 48570 -25 48656 -17
rect 48688 -25 48774 -17
rect 48596 -41 48630 -25
rect 48714 -41 48748 -25
rect 48570 -61 48596 -55
rect 48634 -61 48656 -55
rect 48688 -61 48710 -55
rect 48752 -61 48774 -55
rect 48592 -79 48596 -61
rect 48816 -79 48820 0
rect 49004 -55 49008 0
rect 49052 -17 49134 15
rect 49135 -17 49144 17
rect 49152 -17 49169 17
rect 49050 -25 49136 -17
rect 49177 -25 49179 25
rect 49186 -17 49220 17
rect 49237 -17 49254 17
rect 49279 -25 49281 25
rect 49338 -17 49355 17
rect 49363 -25 49365 25
rect 49456 17 49542 25
rect 49818 17 49904 25
rect 49936 17 50022 25
rect 50298 17 50384 25
rect 49372 -17 49406 17
rect 49423 -17 49440 17
rect 49448 -17 49457 17
rect 49458 15 49491 17
rect 49520 15 49540 17
rect 49458 -17 49540 15
rect 49820 15 49844 17
rect 49869 15 49878 17
rect 49882 15 49902 17
rect 49456 -25 49542 -17
rect 49076 -41 49110 -25
rect 49482 -41 49516 -25
rect 49050 -61 49076 -55
rect 49114 -61 49136 -55
rect 49456 -61 49478 -55
rect 49520 -61 49542 -55
rect 49072 -79 49076 -61
rect 49584 -79 49588 0
rect 49772 -55 49776 0
rect 49820 -17 49902 15
rect 49903 -17 49912 17
rect 49928 -17 49937 17
rect 49938 15 49971 17
rect 50000 15 50020 17
rect 49938 -17 50020 15
rect 50300 15 50324 17
rect 50349 15 50358 17
rect 50362 15 50382 17
rect 49818 -25 49904 -17
rect 49936 -25 50022 -17
rect 49844 -41 49878 -25
rect 49962 -41 49996 -25
rect 49818 -61 49844 -55
rect 49882 -61 49904 -55
rect 49936 -61 49958 -55
rect 50000 -61 50022 -55
rect 49840 -79 49844 -61
rect 50064 -79 50068 0
rect 50252 -55 50256 0
rect 50300 -17 50382 15
rect 50383 -17 50392 17
rect 50400 -17 50417 17
rect 50298 -25 50384 -17
rect 50425 -25 50427 25
rect 50434 -17 50468 17
rect 50485 -17 50502 17
rect 50527 -25 50529 25
rect 50586 -17 50603 17
rect 50611 -25 50613 25
rect 50704 17 50790 25
rect 51066 17 51152 25
rect 51184 17 51270 25
rect 51546 17 51632 25
rect 50620 -17 50654 17
rect 50671 -17 50688 17
rect 50696 -17 50705 17
rect 50706 15 50739 17
rect 50768 15 50788 17
rect 50706 -17 50788 15
rect 51068 15 51092 17
rect 51117 15 51126 17
rect 51130 15 51150 17
rect 50704 -25 50790 -17
rect 50324 -41 50358 -25
rect 50730 -41 50764 -25
rect 50298 -61 50324 -55
rect 50362 -61 50384 -55
rect 50704 -61 50726 -55
rect 50768 -61 50790 -55
rect 50320 -79 50324 -61
rect 50832 -79 50836 0
rect 51020 -55 51024 0
rect 51068 -17 51150 15
rect 51151 -17 51160 17
rect 51176 -17 51185 17
rect 51186 15 51219 17
rect 51248 15 51268 17
rect 51186 -17 51268 15
rect 51548 15 51572 17
rect 51597 15 51606 17
rect 51610 15 51630 17
rect 51066 -25 51152 -17
rect 51184 -25 51270 -17
rect 51092 -41 51126 -25
rect 51210 -41 51244 -25
rect 51066 -61 51092 -55
rect 51130 -61 51152 -55
rect 51184 -61 51206 -55
rect 51248 -61 51270 -55
rect 51088 -79 51092 -61
rect 51312 -79 51316 0
rect 51500 -55 51504 0
rect 51548 -17 51630 15
rect 51631 -17 51640 17
rect 51648 -17 51665 17
rect 51546 -25 51632 -17
rect 51673 -25 51675 25
rect 51682 -17 51716 17
rect 51733 -17 51750 17
rect 51775 -25 51777 25
rect 51834 -17 51851 17
rect 51859 -25 51861 25
rect 51952 17 52038 25
rect 52314 17 52400 25
rect 52432 17 52518 25
rect 52794 17 52880 25
rect 51868 -17 51902 17
rect 51919 -17 51936 17
rect 51944 -17 51953 17
rect 51954 15 51987 17
rect 52016 15 52036 17
rect 51954 -17 52036 15
rect 52316 15 52340 17
rect 52365 15 52374 17
rect 52378 15 52398 17
rect 51952 -25 52038 -17
rect 51572 -41 51606 -25
rect 51978 -41 52012 -25
rect 51546 -61 51572 -55
rect 51610 -61 51632 -55
rect 51952 -61 51974 -55
rect 52016 -61 52038 -55
rect 51568 -79 51572 -61
rect 52080 -79 52084 0
rect 52268 -55 52272 0
rect 52316 -17 52398 15
rect 52399 -17 52408 17
rect 52424 -17 52433 17
rect 52434 15 52467 17
rect 52496 15 52516 17
rect 52434 -17 52516 15
rect 52796 15 52820 17
rect 52845 15 52854 17
rect 52858 15 52878 17
rect 52314 -25 52400 -17
rect 52432 -25 52518 -17
rect 52340 -41 52374 -25
rect 52458 -41 52492 -25
rect 52314 -61 52340 -55
rect 52378 -61 52400 -55
rect 52432 -61 52454 -55
rect 52496 -61 52518 -55
rect 52336 -79 52340 -61
rect 52560 -79 52564 0
rect 52748 -55 52752 0
rect 52796 -17 52878 15
rect 52879 -17 52888 17
rect 52896 -17 52913 17
rect 52794 -25 52880 -17
rect 52921 -25 52923 25
rect 52930 -17 52964 17
rect 52981 -17 52998 17
rect 53023 -25 53025 25
rect 53082 -17 53099 17
rect 53107 -25 53109 25
rect 53200 17 53286 25
rect 53562 17 53648 25
rect 53680 17 53766 25
rect 54042 17 54128 25
rect 53116 -17 53150 17
rect 53167 -17 53184 17
rect 53192 -17 53201 17
rect 53202 15 53235 17
rect 53264 15 53284 17
rect 53202 -17 53284 15
rect 53564 15 53588 17
rect 53613 15 53622 17
rect 53626 15 53646 17
rect 53200 -25 53286 -17
rect 52820 -41 52854 -25
rect 53226 -41 53260 -25
rect 52794 -61 52820 -55
rect 52858 -61 52880 -55
rect 53200 -61 53222 -55
rect 53264 -61 53286 -55
rect 52816 -79 52820 -61
rect 53328 -79 53332 0
rect 53516 -55 53520 0
rect 53564 -17 53646 15
rect 53647 -17 53656 17
rect 53672 -17 53681 17
rect 53682 15 53715 17
rect 53744 15 53764 17
rect 53682 -17 53764 15
rect 54044 15 54068 17
rect 54093 15 54102 17
rect 54106 15 54126 17
rect 53562 -25 53648 -17
rect 53680 -25 53766 -17
rect 53588 -41 53622 -25
rect 53706 -41 53740 -25
rect 53562 -61 53588 -55
rect 53626 -61 53648 -55
rect 53680 -61 53702 -55
rect 53744 -61 53766 -55
rect 53584 -79 53588 -61
rect 53808 -79 53812 0
rect 53996 -55 54000 0
rect 54044 -17 54126 15
rect 54127 -17 54136 17
rect 54144 -17 54161 17
rect 54042 -25 54128 -17
rect 54169 -25 54171 25
rect 54178 -17 54212 17
rect 54229 -17 54246 17
rect 54271 -25 54273 25
rect 54330 -17 54347 17
rect 54355 -25 54357 25
rect 54448 17 54534 25
rect 54810 17 54896 25
rect 54928 17 55014 25
rect 55290 17 55376 25
rect 54364 -17 54398 17
rect 54415 -17 54432 17
rect 54440 -17 54449 17
rect 54450 15 54483 17
rect 54512 15 54532 17
rect 54450 -17 54532 15
rect 54812 15 54836 17
rect 54861 15 54870 17
rect 54874 15 54894 17
rect 54448 -25 54534 -17
rect 54068 -41 54102 -25
rect 54474 -41 54508 -25
rect 54042 -61 54068 -55
rect 54106 -61 54128 -55
rect 54448 -61 54470 -55
rect 54512 -61 54534 -55
rect 54064 -79 54068 -61
rect 54576 -79 54580 0
rect 54764 -55 54768 0
rect 54812 -17 54894 15
rect 54895 -17 54904 17
rect 54920 -17 54929 17
rect 54930 15 54963 17
rect 54992 15 55012 17
rect 54930 -17 55012 15
rect 55292 15 55316 17
rect 55341 15 55350 17
rect 55354 15 55374 17
rect 54810 -25 54896 -17
rect 54928 -25 55014 -17
rect 54836 -41 54870 -25
rect 54954 -41 54988 -25
rect 54810 -61 54836 -55
rect 54874 -61 54896 -55
rect 54928 -61 54950 -55
rect 54992 -61 55014 -55
rect 54832 -79 54836 -61
rect 55056 -79 55060 0
rect 55244 -55 55248 0
rect 55292 -17 55374 15
rect 55375 -17 55384 17
rect 55392 -17 55409 17
rect 55290 -25 55376 -17
rect 55417 -25 55419 25
rect 55426 -17 55460 17
rect 55477 -17 55494 17
rect 55519 -25 55521 25
rect 55578 -17 55595 17
rect 55603 -25 55605 25
rect 55696 17 55782 25
rect 56058 17 56144 25
rect 56176 17 56262 25
rect 56538 17 56624 25
rect 55612 -17 55646 17
rect 55663 -17 55680 17
rect 55688 -17 55697 17
rect 55698 15 55731 17
rect 55760 15 55780 17
rect 55698 -17 55780 15
rect 56060 15 56084 17
rect 56109 15 56118 17
rect 56122 15 56142 17
rect 55696 -25 55782 -17
rect 55316 -41 55350 -25
rect 55722 -41 55756 -25
rect 55290 -61 55316 -55
rect 55354 -61 55376 -55
rect 55696 -61 55718 -55
rect 55760 -61 55782 -55
rect 55312 -79 55316 -61
rect 55824 -79 55828 0
rect 56012 -55 56016 0
rect 56060 -17 56142 15
rect 56143 -17 56152 17
rect 56168 -17 56177 17
rect 56178 15 56211 17
rect 56240 15 56260 17
rect 56178 -17 56260 15
rect 56540 15 56564 17
rect 56589 15 56598 17
rect 56602 15 56622 17
rect 56058 -25 56144 -17
rect 56176 -25 56262 -17
rect 56084 -41 56118 -25
rect 56202 -41 56236 -25
rect 56058 -61 56084 -55
rect 56122 -61 56144 -55
rect 56176 -61 56198 -55
rect 56240 -61 56262 -55
rect 56080 -79 56084 -61
rect 56304 -79 56308 0
rect 56492 -55 56496 0
rect 56540 -17 56622 15
rect 56623 -17 56632 17
rect 56640 -17 56657 17
rect 56538 -25 56624 -17
rect 56665 -25 56667 25
rect 56674 -17 56708 17
rect 56725 -17 56742 17
rect 56767 -25 56769 25
rect 56826 -17 56843 17
rect 56851 -25 56853 25
rect 56944 17 57030 25
rect 57306 17 57392 25
rect 57424 17 57510 25
rect 57786 17 57872 25
rect 56860 -17 56894 17
rect 56911 -17 56928 17
rect 56936 -17 56945 17
rect 56946 15 56979 17
rect 57008 15 57028 17
rect 56946 -17 57028 15
rect 57308 15 57332 17
rect 57357 15 57366 17
rect 57370 15 57390 17
rect 56944 -25 57030 -17
rect 56564 -41 56598 -25
rect 56970 -41 57004 -25
rect 56538 -61 56564 -55
rect 56602 -61 56624 -55
rect 56944 -61 56966 -55
rect 57008 -61 57030 -55
rect 56560 -79 56564 -61
rect 57072 -79 57076 0
rect 57260 -55 57264 0
rect 57308 -17 57390 15
rect 57391 -17 57400 17
rect 57416 -17 57425 17
rect 57426 15 57459 17
rect 57488 15 57508 17
rect 57426 -17 57508 15
rect 57788 15 57812 17
rect 57837 15 57846 17
rect 57850 15 57870 17
rect 57306 -25 57392 -17
rect 57424 -25 57510 -17
rect 57332 -41 57366 -25
rect 57450 -41 57484 -25
rect 57306 -61 57332 -55
rect 57370 -61 57392 -55
rect 57424 -61 57446 -55
rect 57488 -61 57510 -55
rect 57328 -79 57332 -61
rect 57552 -79 57556 0
rect 57740 -55 57744 0
rect 57788 -17 57870 15
rect 57871 -17 57880 17
rect 57888 -17 57905 17
rect 57786 -25 57872 -17
rect 57913 -25 57915 25
rect 57922 -17 57956 17
rect 57973 -17 57990 17
rect 58015 -25 58017 25
rect 58074 -17 58091 17
rect 58099 -25 58101 25
rect 58192 17 58278 25
rect 58554 17 58640 25
rect 58672 17 58758 25
rect 59034 17 59120 25
rect 58108 -17 58142 17
rect 58159 -17 58176 17
rect 58184 -17 58193 17
rect 58194 15 58227 17
rect 58256 15 58276 17
rect 58194 -17 58276 15
rect 58556 15 58580 17
rect 58605 15 58614 17
rect 58618 15 58638 17
rect 58192 -25 58278 -17
rect 57812 -41 57846 -25
rect 58218 -41 58252 -25
rect 57786 -61 57812 -55
rect 57850 -61 57872 -55
rect 58192 -61 58214 -55
rect 58256 -61 58278 -55
rect 57808 -79 57812 -61
rect 58320 -79 58324 0
rect 58508 -55 58512 0
rect 58556 -17 58638 15
rect 58639 -17 58648 17
rect 58664 -17 58673 17
rect 58674 15 58707 17
rect 58736 15 58756 17
rect 58674 -17 58756 15
rect 59036 15 59060 17
rect 59085 15 59094 17
rect 59098 15 59118 17
rect 58554 -25 58640 -17
rect 58672 -25 58758 -17
rect 58580 -41 58614 -25
rect 58698 -41 58732 -25
rect 58554 -61 58580 -55
rect 58618 -61 58640 -55
rect 58672 -61 58694 -55
rect 58736 -61 58758 -55
rect 58576 -79 58580 -61
rect 58800 -79 58804 0
rect 58988 -55 58992 0
rect 59036 -17 59118 15
rect 59119 -17 59128 17
rect 59136 -17 59153 17
rect 59034 -25 59120 -17
rect 59161 -25 59163 25
rect 59170 -17 59204 17
rect 59221 -17 59238 17
rect 59263 -25 59265 25
rect 59322 -17 59339 17
rect 59347 -25 59349 25
rect 59440 17 59526 25
rect 59802 17 59888 25
rect 59920 17 60006 25
rect 60282 17 60368 25
rect 59356 -17 59390 17
rect 59407 -17 59424 17
rect 59432 -17 59441 17
rect 59442 15 59475 17
rect 59504 15 59524 17
rect 59442 -17 59524 15
rect 59804 15 59828 17
rect 59853 15 59862 17
rect 59866 15 59886 17
rect 59440 -25 59526 -17
rect 59060 -41 59094 -25
rect 59466 -41 59500 -25
rect 59034 -61 59060 -55
rect 59098 -61 59120 -55
rect 59440 -61 59462 -55
rect 59504 -61 59526 -55
rect 59056 -79 59060 -61
rect 59568 -79 59572 0
rect 59756 -55 59760 0
rect 59804 -17 59886 15
rect 59887 -17 59896 17
rect 59912 -17 59921 17
rect 59922 15 59955 17
rect 59984 15 60004 17
rect 59922 -17 60004 15
rect 60284 15 60308 17
rect 60333 15 60342 17
rect 60346 15 60366 17
rect 59802 -25 59888 -17
rect 59920 -25 60006 -17
rect 59828 -41 59862 -25
rect 59946 -41 59980 -25
rect 59802 -61 59828 -55
rect 59866 -61 59888 -55
rect 59920 -61 59942 -55
rect 59984 -61 60006 -55
rect 59824 -79 59828 -61
rect 60048 -79 60052 0
rect 60236 -55 60240 0
rect 60284 -17 60366 15
rect 60367 -17 60376 17
rect 60384 -17 60401 17
rect 60282 -25 60368 -17
rect 60409 -25 60411 25
rect 60418 -17 60452 17
rect 60469 -17 60486 17
rect 60511 -25 60513 25
rect 60570 -17 60587 17
rect 60595 -25 60597 25
rect 60688 17 60774 25
rect 61050 17 61136 25
rect 61168 17 61254 25
rect 61530 17 61616 25
rect 60604 -17 60638 17
rect 60655 -17 60672 17
rect 60680 -17 60689 17
rect 60690 15 60723 17
rect 60752 15 60772 17
rect 60690 -17 60772 15
rect 61052 15 61076 17
rect 61101 15 61110 17
rect 61114 15 61134 17
rect 60688 -25 60774 -17
rect 60308 -41 60342 -25
rect 60714 -41 60748 -25
rect 60282 -61 60308 -55
rect 60346 -61 60368 -55
rect 60688 -61 60710 -55
rect 60752 -61 60774 -55
rect 60304 -79 60308 -61
rect 60816 -79 60820 0
rect 61004 -55 61008 0
rect 61052 -17 61134 15
rect 61135 -17 61144 17
rect 61160 -17 61169 17
rect 61170 15 61203 17
rect 61232 15 61252 17
rect 61170 -17 61252 15
rect 61532 15 61556 17
rect 61581 15 61590 17
rect 61594 15 61614 17
rect 61050 -25 61136 -17
rect 61168 -25 61254 -17
rect 61076 -41 61110 -25
rect 61194 -41 61228 -25
rect 61050 -61 61076 -55
rect 61114 -61 61136 -55
rect 61168 -61 61190 -55
rect 61232 -61 61254 -55
rect 61072 -79 61076 -61
rect 61296 -79 61300 0
rect 61484 -55 61488 0
rect 61532 -17 61614 15
rect 61615 -17 61624 17
rect 61632 -17 61649 17
rect 61530 -25 61616 -17
rect 61657 -25 61659 25
rect 61666 -17 61700 17
rect 61717 -17 61734 17
rect 61759 -25 61761 25
rect 61818 -17 61835 17
rect 61843 -25 61845 25
rect 61936 17 62022 25
rect 62298 17 62384 25
rect 62416 17 62502 25
rect 62778 17 62864 25
rect 61852 -17 61886 17
rect 61903 -17 61920 17
rect 61928 -17 61937 17
rect 61938 15 61971 17
rect 62000 15 62020 17
rect 61938 -17 62020 15
rect 62300 15 62324 17
rect 62349 15 62358 17
rect 62362 15 62382 17
rect 61936 -25 62022 -17
rect 61556 -41 61590 -25
rect 61962 -41 61996 -25
rect 61530 -61 61556 -55
rect 61594 -61 61616 -55
rect 61936 -61 61958 -55
rect 62000 -61 62022 -55
rect 61552 -79 61556 -61
rect 62064 -79 62068 0
rect 62252 -55 62256 0
rect 62300 -17 62382 15
rect 62383 -17 62392 17
rect 62408 -17 62417 17
rect 62418 15 62451 17
rect 62480 15 62500 17
rect 62418 -17 62500 15
rect 62780 15 62804 17
rect 62829 15 62838 17
rect 62842 15 62862 17
rect 62298 -25 62384 -17
rect 62416 -25 62502 -17
rect 62324 -41 62358 -25
rect 62442 -41 62476 -25
rect 62298 -61 62324 -55
rect 62362 -61 62384 -55
rect 62416 -61 62438 -55
rect 62480 -61 62502 -55
rect 62320 -79 62324 -61
rect 62544 -79 62548 0
rect 62732 -55 62736 0
rect 62780 -17 62862 15
rect 62863 -17 62872 17
rect 62880 -17 62897 17
rect 62778 -25 62864 -17
rect 62905 -25 62907 25
rect 62914 -17 62948 17
rect 62965 -17 62982 17
rect 63007 -25 63009 25
rect 63066 -17 63083 17
rect 63091 -25 63093 25
rect 63184 17 63270 25
rect 63546 17 63632 25
rect 63664 17 63750 25
rect 64026 17 64112 25
rect 63100 -17 63134 17
rect 63151 -17 63168 17
rect 63176 -17 63185 17
rect 63186 15 63219 17
rect 63248 15 63268 17
rect 63186 -17 63268 15
rect 63548 15 63572 17
rect 63597 15 63606 17
rect 63610 15 63630 17
rect 63184 -25 63270 -17
rect 62804 -41 62838 -25
rect 63210 -41 63244 -25
rect 62778 -61 62804 -55
rect 62842 -61 62864 -55
rect 63184 -61 63206 -55
rect 63248 -61 63270 -55
rect 62800 -79 62804 -61
rect 63312 -79 63316 0
rect 63500 -55 63504 0
rect 63548 -17 63630 15
rect 63631 -17 63640 17
rect 63656 -17 63665 17
rect 63666 15 63699 17
rect 63728 15 63748 17
rect 63666 -17 63748 15
rect 64028 15 64052 17
rect 64077 15 64086 17
rect 64090 15 64110 17
rect 63546 -25 63632 -17
rect 63664 -25 63750 -17
rect 63572 -41 63606 -25
rect 63690 -41 63724 -25
rect 63546 -61 63572 -55
rect 63610 -61 63632 -55
rect 63664 -61 63686 -55
rect 63728 -61 63750 -55
rect 63568 -79 63572 -61
rect 63792 -79 63796 0
rect 63980 -55 63984 0
rect 64028 -17 64110 15
rect 64111 -17 64120 17
rect 64128 -17 64145 17
rect 64026 -25 64112 -17
rect 64153 -25 64155 25
rect 64162 -17 64196 17
rect 64213 -17 64230 17
rect 64255 -25 64257 25
rect 64314 -17 64331 17
rect 64339 -25 64341 25
rect 64432 17 64518 25
rect 64794 17 64880 25
rect 64912 17 64998 25
rect 65274 17 65360 25
rect 64348 -17 64382 17
rect 64399 -17 64416 17
rect 64424 -17 64433 17
rect 64434 15 64467 17
rect 64496 15 64516 17
rect 64434 -17 64516 15
rect 64796 15 64820 17
rect 64845 15 64854 17
rect 64858 15 64878 17
rect 64432 -25 64518 -17
rect 64052 -41 64086 -25
rect 64458 -41 64492 -25
rect 64026 -61 64052 -55
rect 64090 -61 64112 -55
rect 64432 -61 64454 -55
rect 64496 -61 64518 -55
rect 64048 -79 64052 -61
rect 64560 -79 64564 0
rect 64748 -55 64752 0
rect 64796 -17 64878 15
rect 64879 -17 64888 17
rect 64904 -17 64913 17
rect 64914 15 64947 17
rect 64976 15 64996 17
rect 64914 -17 64996 15
rect 65276 15 65300 17
rect 65325 15 65334 17
rect 65338 15 65358 17
rect 64794 -25 64880 -17
rect 64912 -25 64998 -17
rect 64820 -41 64854 -25
rect 64938 -41 64972 -25
rect 64794 -61 64820 -55
rect 64858 -61 64880 -55
rect 64912 -61 64934 -55
rect 64976 -61 64998 -55
rect 64816 -79 64820 -61
rect 65040 -79 65044 0
rect 65228 -55 65232 0
rect 65276 -17 65358 15
rect 65359 -17 65368 17
rect 65376 -17 65393 17
rect 65274 -25 65360 -17
rect 65401 -25 65403 25
rect 65410 -17 65444 17
rect 65461 -17 65478 17
rect 65503 -25 65505 25
rect 65562 -17 65579 17
rect 65587 -25 65589 25
rect 65680 17 65766 25
rect 66042 17 66128 25
rect 66160 17 66246 25
rect 66522 17 66608 25
rect 65596 -17 65630 17
rect 65647 -17 65664 17
rect 65672 -17 65681 17
rect 65682 15 65715 17
rect 65744 15 65764 17
rect 65682 -17 65764 15
rect 66044 15 66068 17
rect 66093 15 66102 17
rect 66106 15 66126 17
rect 65680 -25 65766 -17
rect 65300 -41 65334 -25
rect 65706 -41 65740 -25
rect 65274 -61 65300 -55
rect 65338 -61 65360 -55
rect 65680 -61 65702 -55
rect 65744 -61 65766 -55
rect 65296 -79 65300 -61
rect 65808 -79 65812 0
rect 65996 -55 66000 0
rect 66044 -17 66126 15
rect 66127 -17 66136 17
rect 66152 -17 66161 17
rect 66162 15 66195 17
rect 66224 15 66244 17
rect 66162 -17 66244 15
rect 66524 15 66548 17
rect 66573 15 66582 17
rect 66586 15 66606 17
rect 66042 -25 66128 -17
rect 66160 -25 66246 -17
rect 66068 -41 66102 -25
rect 66186 -41 66220 -25
rect 66042 -61 66068 -55
rect 66106 -61 66128 -55
rect 66160 -61 66182 -55
rect 66224 -61 66246 -55
rect 66064 -79 66068 -61
rect 66288 -79 66292 0
rect 66476 -55 66480 0
rect 66524 -17 66606 15
rect 66607 -17 66616 17
rect 66624 -17 66641 17
rect 66522 -25 66608 -17
rect 66649 -25 66651 25
rect 66658 -17 66692 17
rect 66709 -17 66726 17
rect 66751 -25 66753 25
rect 66810 -17 66827 17
rect 66835 -25 66837 25
rect 66928 17 67014 25
rect 67290 17 67376 25
rect 67408 17 67494 25
rect 67770 17 67856 25
rect 66844 -17 66878 17
rect 66895 -17 66912 17
rect 66920 -17 66929 17
rect 66930 15 66963 17
rect 66992 15 67012 17
rect 66930 -17 67012 15
rect 67292 15 67316 17
rect 67341 15 67350 17
rect 67354 15 67374 17
rect 66928 -25 67014 -17
rect 66548 -41 66582 -25
rect 66954 -41 66988 -25
rect 66522 -61 66548 -55
rect 66586 -61 66608 -55
rect 66928 -61 66950 -55
rect 66992 -61 67014 -55
rect 66544 -79 66548 -61
rect 67056 -79 67060 0
rect 67244 -55 67248 0
rect 67292 -17 67374 15
rect 67375 -17 67384 17
rect 67400 -17 67409 17
rect 67410 15 67443 17
rect 67472 15 67492 17
rect 67410 -17 67492 15
rect 67772 15 67796 17
rect 67821 15 67830 17
rect 67834 15 67854 17
rect 67290 -25 67376 -17
rect 67408 -25 67494 -17
rect 67316 -41 67350 -25
rect 67434 -41 67468 -25
rect 67290 -61 67316 -55
rect 67354 -61 67376 -55
rect 67408 -61 67430 -55
rect 67472 -61 67494 -55
rect 67312 -79 67316 -61
rect 67536 -79 67540 0
rect 67724 -55 67728 0
rect 67772 -17 67854 15
rect 67855 -17 67864 17
rect 67872 -17 67889 17
rect 67770 -25 67856 -17
rect 67897 -25 67899 25
rect 67906 -17 67940 17
rect 67957 -17 67974 17
rect 67999 -25 68001 25
rect 68058 -17 68075 17
rect 68083 -25 68085 25
rect 68176 17 68262 25
rect 68538 17 68624 25
rect 68656 17 68742 25
rect 69018 17 69104 25
rect 68092 -17 68126 17
rect 68143 -17 68160 17
rect 68168 -17 68177 17
rect 68178 15 68211 17
rect 68240 15 68260 17
rect 68178 -17 68260 15
rect 68540 15 68564 17
rect 68589 15 68598 17
rect 68602 15 68622 17
rect 68176 -25 68262 -17
rect 67796 -41 67830 -25
rect 68202 -41 68236 -25
rect 67770 -61 67796 -55
rect 67834 -61 67856 -55
rect 68176 -61 68198 -55
rect 68240 -61 68262 -55
rect 67792 -79 67796 -61
rect 68304 -79 68308 0
rect 68492 -55 68496 0
rect 68540 -17 68622 15
rect 68623 -17 68632 17
rect 68648 -17 68657 17
rect 68658 15 68691 17
rect 68720 15 68740 17
rect 68658 -17 68740 15
rect 69020 15 69044 17
rect 69069 15 69078 17
rect 69082 15 69102 17
rect 68538 -25 68624 -17
rect 68656 -25 68742 -17
rect 68564 -41 68598 -25
rect 68682 -41 68716 -25
rect 68538 -61 68564 -55
rect 68602 -61 68624 -55
rect 68656 -61 68678 -55
rect 68720 -61 68742 -55
rect 68560 -79 68564 -61
rect 68784 -79 68788 0
rect 68972 -55 68976 0
rect 69020 -17 69102 15
rect 69103 -17 69112 17
rect 69120 -17 69137 17
rect 69018 -25 69104 -17
rect 69145 -25 69147 25
rect 69154 -17 69188 17
rect 69205 -17 69222 17
rect 69247 -25 69249 25
rect 69306 -17 69323 17
rect 69331 -25 69333 25
rect 69424 17 69510 25
rect 69786 17 69872 25
rect 69904 17 69990 25
rect 70266 17 70352 25
rect 69340 -17 69374 17
rect 69391 -17 69408 17
rect 69416 -17 69425 17
rect 69426 15 69459 17
rect 69488 15 69508 17
rect 69426 -17 69508 15
rect 69788 15 69812 17
rect 69837 15 69846 17
rect 69850 15 69870 17
rect 69424 -25 69510 -17
rect 69044 -41 69078 -25
rect 69450 -41 69484 -25
rect 69018 -61 69044 -55
rect 69082 -61 69104 -55
rect 69424 -61 69446 -55
rect 69488 -61 69510 -55
rect 69040 -79 69044 -61
rect 69552 -79 69556 0
rect 69740 -55 69744 0
rect 69788 -17 69870 15
rect 69871 -17 69880 17
rect 69896 -17 69905 17
rect 69906 15 69939 17
rect 69968 15 69988 17
rect 69906 -17 69988 15
rect 70268 15 70292 17
rect 70317 15 70326 17
rect 70330 15 70350 17
rect 69786 -25 69872 -17
rect 69904 -25 69990 -17
rect 69812 -41 69846 -25
rect 69930 -41 69964 -25
rect 69786 -61 69812 -55
rect 69850 -61 69872 -55
rect 69904 -61 69926 -55
rect 69968 -61 69990 -55
rect 69808 -79 69812 -61
rect 70032 -79 70036 0
rect 70220 -55 70224 0
rect 70268 -17 70350 15
rect 70351 -17 70360 17
rect 70368 -17 70385 17
rect 70266 -25 70352 -17
rect 70393 -25 70395 25
rect 70402 -17 70436 17
rect 70453 -17 70470 17
rect 70495 -25 70497 25
rect 70554 -17 70571 17
rect 70579 -25 70581 25
rect 70672 17 70758 25
rect 71034 17 71120 25
rect 71152 17 71238 25
rect 71514 17 71600 25
rect 70588 -17 70622 17
rect 70639 -17 70656 17
rect 70664 -17 70673 17
rect 70674 15 70707 17
rect 70736 15 70756 17
rect 70674 -17 70756 15
rect 71036 15 71060 17
rect 71085 15 71094 17
rect 71098 15 71118 17
rect 70672 -25 70758 -17
rect 70292 -41 70326 -25
rect 70698 -41 70732 -25
rect 70266 -61 70292 -55
rect 70330 -61 70352 -55
rect 70672 -61 70694 -55
rect 70736 -61 70758 -55
rect 70288 -79 70292 -61
rect 70800 -79 70804 0
rect 70988 -55 70992 0
rect 71036 -17 71118 15
rect 71119 -17 71128 17
rect 71144 -17 71153 17
rect 71154 15 71187 17
rect 71216 15 71236 17
rect 71154 -17 71236 15
rect 71516 15 71540 17
rect 71565 15 71574 17
rect 71578 15 71598 17
rect 71034 -25 71120 -17
rect 71152 -25 71238 -17
rect 71060 -41 71094 -25
rect 71178 -41 71212 -25
rect 71034 -61 71060 -55
rect 71098 -61 71120 -55
rect 71152 -61 71174 -55
rect 71216 -61 71238 -55
rect 71056 -79 71060 -61
rect 71280 -79 71284 0
rect 71468 -55 71472 0
rect 71516 -17 71598 15
rect 71599 -17 71608 17
rect 71616 -17 71633 17
rect 71514 -25 71600 -17
rect 71641 -25 71643 25
rect 71650 -17 71684 17
rect 71701 -17 71718 17
rect 71743 -25 71745 25
rect 71802 -17 71819 17
rect 71827 -25 71829 25
rect 71920 17 72006 25
rect 72282 17 72368 25
rect 72400 17 72486 25
rect 72762 17 72848 25
rect 71836 -17 71870 17
rect 71887 -17 71904 17
rect 71912 -17 71921 17
rect 71922 15 71955 17
rect 71984 15 72004 17
rect 71922 -17 72004 15
rect 72284 15 72308 17
rect 72333 15 72342 17
rect 72346 15 72366 17
rect 71920 -25 72006 -17
rect 71540 -41 71574 -25
rect 71946 -41 71980 -25
rect 71514 -61 71540 -55
rect 71578 -61 71600 -55
rect 71920 -61 71942 -55
rect 71984 -61 72006 -55
rect 71536 -79 71540 -61
rect 72048 -79 72052 0
rect 72236 -55 72240 0
rect 72284 -17 72366 15
rect 72367 -17 72376 17
rect 72392 -17 72401 17
rect 72402 15 72435 17
rect 72464 15 72484 17
rect 72402 -17 72484 15
rect 72764 15 72788 17
rect 72813 15 72822 17
rect 72826 15 72846 17
rect 72282 -25 72368 -17
rect 72400 -25 72486 -17
rect 72308 -41 72342 -25
rect 72426 -41 72460 -25
rect 72282 -61 72308 -55
rect 72346 -61 72368 -55
rect 72400 -61 72422 -55
rect 72464 -61 72486 -55
rect 72304 -79 72308 -61
rect 72528 -79 72532 0
rect 72716 -55 72720 0
rect 72764 -17 72846 15
rect 72847 -17 72856 17
rect 72864 -17 72881 17
rect 72762 -25 72848 -17
rect 72889 -25 72891 25
rect 72898 -17 72932 17
rect 72949 -17 72966 17
rect 72991 -25 72993 25
rect 73050 -17 73067 17
rect 73075 -25 73077 25
rect 73168 17 73254 25
rect 73530 17 73616 25
rect 73648 17 73734 25
rect 74010 17 74096 25
rect 73084 -17 73118 17
rect 73135 -17 73152 17
rect 73160 -17 73169 17
rect 73170 15 73203 17
rect 73232 15 73252 17
rect 73170 -17 73252 15
rect 73532 15 73556 17
rect 73581 15 73590 17
rect 73594 15 73614 17
rect 73168 -25 73254 -17
rect 72788 -41 72822 -25
rect 73194 -41 73228 -25
rect 72762 -61 72788 -55
rect 72826 -61 72848 -55
rect 73168 -61 73190 -55
rect 73232 -61 73254 -55
rect 72784 -79 72788 -61
rect 73296 -79 73300 0
rect 73484 -55 73488 0
rect 73532 -17 73614 15
rect 73615 -17 73624 17
rect 73640 -17 73649 17
rect 73650 15 73683 17
rect 73712 15 73732 17
rect 73650 -17 73732 15
rect 74012 15 74036 17
rect 74061 15 74070 17
rect 74074 15 74094 17
rect 73530 -25 73616 -17
rect 73648 -25 73734 -17
rect 73556 -41 73590 -25
rect 73674 -41 73708 -25
rect 73530 -61 73556 -55
rect 73594 -61 73616 -55
rect 73648 -61 73670 -55
rect 73712 -61 73734 -55
rect 73552 -79 73556 -61
rect 73776 -79 73780 0
rect 73964 -55 73968 0
rect 74012 -17 74094 15
rect 74095 -17 74104 17
rect 74112 -17 74129 17
rect 74010 -25 74096 -17
rect 74137 -25 74139 25
rect 74146 -17 74180 17
rect 74197 -17 74214 17
rect 74239 -25 74241 25
rect 74298 -17 74315 17
rect 74323 -25 74325 25
rect 74416 17 74502 25
rect 74778 17 74864 25
rect 74896 17 74982 25
rect 75258 17 75344 25
rect 74332 -17 74366 17
rect 74383 -17 74400 17
rect 74408 -17 74417 17
rect 74418 15 74451 17
rect 74480 15 74500 17
rect 74418 -17 74500 15
rect 74780 15 74804 17
rect 74829 15 74838 17
rect 74842 15 74862 17
rect 74416 -25 74502 -17
rect 74036 -41 74070 -25
rect 74442 -41 74476 -25
rect 74010 -61 74036 -55
rect 74074 -61 74096 -55
rect 74416 -61 74438 -55
rect 74480 -61 74502 -55
rect 74032 -79 74036 -61
rect 74544 -79 74548 0
rect 74732 -55 74736 0
rect 74780 -17 74862 15
rect 74863 -17 74872 17
rect 74888 -17 74897 17
rect 74898 15 74931 17
rect 74960 15 74980 17
rect 74898 -17 74980 15
rect 75260 15 75284 17
rect 75309 15 75318 17
rect 75322 15 75342 17
rect 74778 -25 74864 -17
rect 74896 -25 74982 -17
rect 74804 -41 74838 -25
rect 74922 -41 74956 -25
rect 74778 -61 74804 -55
rect 74842 -61 74864 -55
rect 74896 -61 74918 -55
rect 74960 -61 74982 -55
rect 74800 -79 74804 -61
rect 75024 -79 75028 0
rect 75212 -55 75216 0
rect 75260 -17 75342 15
rect 75343 -17 75352 17
rect 75360 -17 75377 17
rect 75258 -25 75344 -17
rect 75385 -25 75387 25
rect 75394 -17 75428 17
rect 75445 -17 75462 17
rect 75487 -25 75489 25
rect 75546 -17 75563 17
rect 75571 -25 75573 25
rect 75664 17 75750 25
rect 76026 17 76112 25
rect 76144 17 76230 25
rect 76506 17 76592 25
rect 75580 -17 75614 17
rect 75631 -17 75648 17
rect 75656 -17 75665 17
rect 75666 15 75699 17
rect 75728 15 75748 17
rect 75666 -17 75748 15
rect 76028 15 76052 17
rect 76077 15 76086 17
rect 76090 15 76110 17
rect 75664 -25 75750 -17
rect 75284 -41 75318 -25
rect 75690 -41 75724 -25
rect 75258 -61 75284 -55
rect 75322 -61 75344 -55
rect 75664 -61 75686 -55
rect 75728 -61 75750 -55
rect 75280 -79 75284 -61
rect 75792 -79 75796 0
rect 75980 -55 75984 0
rect 76028 -17 76110 15
rect 76111 -17 76120 17
rect 76136 -17 76145 17
rect 76146 15 76179 17
rect 76208 15 76228 17
rect 76146 -17 76228 15
rect 76508 15 76532 17
rect 76557 15 76566 17
rect 76570 15 76590 17
rect 76026 -25 76112 -17
rect 76144 -25 76230 -17
rect 76052 -41 76086 -25
rect 76170 -41 76204 -25
rect 76026 -61 76052 -55
rect 76090 -61 76112 -55
rect 76144 -61 76166 -55
rect 76208 -61 76230 -55
rect 76048 -79 76052 -61
rect 76272 -79 76276 0
rect 76460 -55 76464 0
rect 76508 -17 76590 15
rect 76591 -17 76600 17
rect 76608 -17 76625 17
rect 76506 -25 76592 -17
rect 76633 -25 76635 25
rect 76642 -17 76676 17
rect 76693 -17 76710 17
rect 76735 -25 76737 25
rect 76794 -17 76811 17
rect 76819 -25 76821 25
rect 76912 17 76998 25
rect 77274 17 77360 25
rect 77392 17 77478 25
rect 77754 17 77840 25
rect 76828 -17 76862 17
rect 76879 -17 76896 17
rect 76904 -17 76913 17
rect 76914 15 76947 17
rect 76976 15 76996 17
rect 76914 -17 76996 15
rect 77276 15 77300 17
rect 77325 15 77334 17
rect 77338 15 77358 17
rect 76912 -25 76998 -17
rect 76532 -41 76566 -25
rect 76938 -41 76972 -25
rect 76506 -61 76532 -55
rect 76570 -61 76592 -55
rect 76912 -61 76934 -55
rect 76976 -61 76998 -55
rect 76528 -79 76532 -61
rect 77040 -79 77044 0
rect 77228 -55 77232 0
rect 77276 -17 77358 15
rect 77359 -17 77368 17
rect 77384 -17 77393 17
rect 77394 15 77427 17
rect 77456 15 77476 17
rect 77394 -17 77476 15
rect 77756 15 77780 17
rect 77805 15 77814 17
rect 77818 15 77838 17
rect 77274 -25 77360 -17
rect 77392 -25 77478 -17
rect 77300 -41 77334 -25
rect 77418 -41 77452 -25
rect 77274 -61 77300 -55
rect 77338 -61 77360 -55
rect 77392 -61 77414 -55
rect 77456 -61 77478 -55
rect 77296 -79 77300 -61
rect 77520 -79 77524 0
rect 77708 -55 77712 0
rect 77756 -17 77838 15
rect 77839 -17 77848 17
rect 77856 -17 77873 17
rect 77754 -25 77840 -17
rect 77881 -25 77883 25
rect 77890 -17 77924 17
rect 77941 -17 77958 17
rect 77983 -25 77985 25
rect 78042 -17 78059 17
rect 78067 -25 78069 25
rect 78160 17 78246 25
rect 78522 17 78608 25
rect 78640 17 78726 25
rect 79002 17 79088 25
rect 78076 -17 78110 17
rect 78127 -17 78144 17
rect 78152 -17 78161 17
rect 78162 15 78195 17
rect 78224 15 78244 17
rect 78162 -17 78244 15
rect 78524 15 78548 17
rect 78573 15 78582 17
rect 78586 15 78606 17
rect 78160 -25 78246 -17
rect 77780 -41 77814 -25
rect 78186 -41 78220 -25
rect 77754 -61 77780 -55
rect 77818 -61 77840 -55
rect 78160 -61 78182 -55
rect 78224 -61 78246 -55
rect 77776 -79 77780 -61
rect 78288 -79 78292 0
rect 78476 -55 78480 0
rect 78524 -17 78606 15
rect 78607 -17 78616 17
rect 78632 -17 78641 17
rect 78642 15 78675 17
rect 78704 15 78724 17
rect 78642 -17 78724 15
rect 79004 15 79028 17
rect 79053 15 79062 17
rect 79066 15 79086 17
rect 78522 -25 78608 -17
rect 78640 -25 78726 -17
rect 78548 -41 78582 -25
rect 78666 -41 78700 -25
rect 78522 -61 78548 -55
rect 78586 -61 78608 -55
rect 78640 -61 78662 -55
rect 78704 -61 78726 -55
rect 78544 -79 78548 -61
rect 78768 -79 78772 0
rect 78956 -55 78960 0
rect 79004 -17 79086 15
rect 79087 -17 79096 17
rect 79104 -17 79121 17
rect 79002 -25 79088 -17
rect 79129 -25 79131 25
rect 79138 -17 79172 17
rect 79189 -17 79206 17
rect 79231 -25 79233 25
rect 79290 -17 79307 17
rect 79315 -25 79317 25
rect 79408 17 79494 25
rect 79770 17 79856 25
rect 79324 -17 79358 17
rect 79375 -17 79392 17
rect 79400 -17 79409 17
rect 79410 15 79443 17
rect 79472 15 79492 17
rect 79410 -17 79492 15
rect 79772 15 79796 17
rect 79821 15 79830 17
rect 79834 15 79854 17
rect 79408 -25 79494 -17
rect 79028 -41 79062 -25
rect 79434 -41 79468 -25
rect 79002 -61 79028 -55
rect 79066 -61 79088 -55
rect 79408 -61 79430 -55
rect 79472 -61 79494 -55
rect 79024 -79 79028 -61
rect 79536 -79 79540 0
rect 79724 -55 79728 0
rect 79772 -17 79854 15
rect 79855 -17 79864 17
rect 79770 -25 79856 -17
rect 79897 -25 79899 25
rect 79796 -41 79830 -25
rect 79770 -61 79796 -55
rect 79834 -61 79856 -55
rect 79792 -79 79796 -61
rect 38 -105 80 -79
rect 400 -105 442 -79
rect 806 -105 848 -79
rect 1168 -105 1210 -79
rect 1286 -105 1328 -79
rect 1648 -105 1690 -79
rect 2054 -105 2096 -79
rect 2416 -105 2458 -79
rect 2534 -105 2576 -79
rect 2896 -105 2938 -79
rect 3302 -105 3344 -79
rect 3664 -105 3706 -79
rect 3782 -105 3824 -79
rect 4144 -105 4186 -79
rect 4550 -105 4592 -79
rect 4912 -105 4954 -79
rect 5030 -105 5072 -79
rect 5392 -105 5434 -79
rect 5798 -105 5840 -79
rect 6160 -105 6202 -79
rect 6278 -105 6320 -79
rect 6640 -105 6682 -79
rect 7046 -105 7088 -79
rect 7408 -105 7450 -79
rect 7526 -105 7568 -79
rect 7888 -105 7930 -79
rect 8294 -105 8336 -79
rect 8656 -105 8698 -79
rect 8774 -105 8816 -79
rect 9136 -105 9178 -79
rect 9542 -105 9584 -79
rect 9904 -105 9946 -79
rect 10022 -105 10064 -79
rect 10384 -105 10426 -79
rect 10790 -105 10832 -79
rect 11152 -105 11194 -79
rect 11270 -105 11312 -79
rect 11632 -105 11674 -79
rect 12038 -105 12080 -79
rect 12400 -105 12442 -79
rect 12518 -105 12560 -79
rect 12880 -105 12922 -79
rect 13286 -105 13328 -79
rect 13648 -105 13690 -79
rect 13766 -105 13808 -79
rect 14128 -105 14170 -79
rect 14534 -105 14576 -79
rect 14896 -105 14938 -79
rect 15014 -105 15056 -79
rect 15376 -105 15418 -79
rect 15782 -105 15824 -79
rect 16144 -105 16186 -79
rect 16262 -105 16304 -79
rect 16624 -105 16666 -79
rect 17030 -105 17072 -79
rect 17392 -105 17434 -79
rect 17510 -105 17552 -79
rect 17872 -105 17914 -79
rect 18278 -105 18320 -79
rect 18640 -105 18682 -79
rect 18758 -105 18800 -79
rect 19120 -105 19162 -79
rect 19526 -105 19568 -79
rect 19888 -105 19930 -79
rect 20006 -105 20048 -79
rect 20368 -105 20410 -79
rect 20774 -105 20816 -79
rect 21136 -105 21178 -79
rect 21254 -105 21296 -79
rect 21616 -105 21658 -79
rect 22022 -105 22064 -79
rect 22384 -105 22426 -79
rect 22502 -105 22544 -79
rect 22864 -105 22906 -79
rect 23270 -105 23312 -79
rect 23632 -105 23674 -79
rect 23750 -105 23792 -79
rect 24112 -105 24154 -79
rect 24518 -105 24560 -79
rect 24880 -105 24922 -79
rect 24998 -105 25040 -79
rect 25360 -105 25402 -79
rect 25766 -105 25808 -79
rect 26128 -105 26170 -79
rect 26246 -105 26288 -79
rect 26608 -105 26650 -79
rect 27014 -105 27056 -79
rect 27376 -105 27418 -79
rect 27494 -105 27536 -79
rect 27856 -105 27898 -79
rect 28262 -105 28304 -79
rect 28624 -105 28666 -79
rect 28742 -105 28784 -79
rect 29104 -105 29146 -79
rect 29510 -105 29552 -79
rect 29872 -105 29914 -79
rect 29990 -105 30032 -79
rect 30352 -105 30394 -79
rect 30758 -105 30800 -79
rect 31120 -105 31162 -79
rect 31238 -105 31280 -79
rect 31600 -105 31642 -79
rect 32006 -105 32048 -79
rect 32368 -105 32410 -79
rect 32486 -105 32528 -79
rect 32848 -105 32890 -79
rect 33254 -105 33296 -79
rect 33616 -105 33658 -79
rect 33734 -105 33776 -79
rect 34096 -105 34138 -79
rect 34502 -105 34544 -79
rect 34864 -105 34906 -79
rect 34982 -105 35024 -79
rect 35344 -105 35386 -79
rect 35750 -105 35792 -79
rect 36112 -105 36154 -79
rect 36230 -105 36272 -79
rect 36592 -105 36634 -79
rect 36998 -105 37040 -79
rect 37360 -105 37402 -79
rect 37478 -105 37520 -79
rect 37840 -105 37882 -79
rect 38246 -105 38288 -79
rect 38608 -105 38650 -79
rect 38726 -105 38768 -79
rect 39088 -105 39130 -79
rect 39494 -105 39536 -79
rect 39856 -105 39898 -79
rect 39974 -105 40016 -79
rect 40336 -105 40378 -79
rect 40742 -105 40784 -79
rect 41104 -105 41146 -79
rect 41222 -105 41264 -79
rect 41584 -105 41626 -79
rect 41990 -105 42032 -79
rect 42352 -105 42394 -79
rect 42470 -105 42512 -79
rect 42832 -105 42874 -79
rect 43238 -105 43280 -79
rect 43600 -105 43642 -79
rect 43718 -105 43760 -79
rect 44080 -105 44122 -79
rect 44486 -105 44528 -79
rect 44848 -105 44890 -79
rect 44966 -105 45008 -79
rect 45328 -105 45370 -79
rect 45734 -105 45776 -79
rect 46096 -105 46138 -79
rect 46214 -105 46256 -79
rect 46576 -105 46618 -79
rect 46982 -105 47024 -79
rect 47344 -105 47386 -79
rect 47462 -105 47504 -79
rect 47824 -105 47866 -79
rect 48230 -105 48272 -79
rect 48592 -105 48634 -79
rect 48710 -105 48752 -79
rect 49072 -105 49114 -79
rect 49478 -105 49520 -79
rect 49840 -105 49882 -79
rect 49958 -105 50000 -79
rect 50320 -105 50362 -79
rect 50726 -105 50768 -79
rect 51088 -105 51130 -79
rect 51206 -105 51248 -79
rect 51568 -105 51610 -79
rect 51974 -105 52016 -79
rect 52336 -105 52378 -79
rect 52454 -105 52496 -79
rect 52816 -105 52858 -79
rect 53222 -105 53264 -79
rect 53584 -105 53626 -79
rect 53702 -105 53744 -79
rect 54064 -105 54106 -79
rect 54470 -105 54512 -79
rect 54832 -105 54874 -79
rect 54950 -105 54992 -79
rect 55312 -105 55354 -79
rect 55718 -105 55760 -79
rect 56080 -105 56122 -79
rect 56198 -105 56240 -79
rect 56560 -105 56602 -79
rect 56966 -105 57008 -79
rect 57328 -105 57370 -79
rect 57446 -105 57488 -79
rect 57808 -105 57850 -79
rect 58214 -105 58256 -79
rect 58576 -105 58618 -79
rect 58694 -105 58736 -79
rect 59056 -105 59098 -79
rect 59462 -105 59504 -79
rect 59824 -105 59866 -79
rect 59942 -105 59984 -79
rect 60304 -105 60346 -79
rect 60710 -105 60752 -79
rect 61072 -105 61114 -79
rect 61190 -105 61232 -79
rect 61552 -105 61594 -79
rect 61958 -105 62000 -79
rect 62320 -105 62362 -79
rect 62438 -105 62480 -79
rect 62800 -105 62842 -79
rect 63206 -105 63248 -79
rect 63568 -105 63610 -79
rect 63686 -105 63728 -79
rect 64048 -105 64090 -79
rect 64454 -105 64496 -79
rect 64816 -105 64858 -79
rect 64934 -105 64976 -79
rect 65296 -105 65338 -79
rect 65702 -105 65744 -79
rect 66064 -105 66106 -79
rect 66182 -105 66224 -79
rect 66544 -105 66586 -79
rect 66950 -105 66992 -79
rect 67312 -105 67354 -79
rect 67430 -105 67472 -79
rect 67792 -105 67834 -79
rect 68198 -105 68240 -79
rect 68560 -105 68602 -79
rect 68678 -105 68720 -79
rect 69040 -105 69082 -79
rect 69446 -105 69488 -79
rect 69808 -105 69850 -79
rect 69926 -105 69968 -79
rect 70288 -105 70330 -79
rect 70694 -105 70736 -79
rect 71056 -105 71098 -79
rect 71174 -105 71216 -79
rect 71536 -105 71578 -79
rect 71942 -105 71984 -79
rect 72304 -105 72346 -79
rect 72422 -105 72464 -79
rect 72784 -105 72826 -79
rect 73190 -105 73232 -79
rect 73552 -105 73594 -79
rect 73670 -105 73712 -79
rect 74032 -105 74074 -79
rect 74438 -105 74480 -79
rect 74800 -105 74842 -79
rect 74918 -105 74960 -79
rect 75280 -105 75322 -79
rect 75686 -105 75728 -79
rect 76048 -105 76090 -79
rect 76166 -105 76208 -79
rect 76528 -105 76570 -79
rect 76934 -105 76976 -79
rect 77296 -105 77338 -79
rect 77414 -105 77456 -79
rect 77776 -105 77818 -79
rect 78182 -105 78224 -79
rect 78544 -105 78586 -79
rect 78662 -105 78704 -79
rect 79024 -105 79066 -79
rect 79430 -105 79472 -79
rect 79792 -105 79834 -79
<< metal1 >>
rect 78 0 114 395
rect 150 0 186 395
rect 222 79 258 420
rect 294 0 330 395
rect 366 0 402 395
rect 846 0 882 395
rect 918 0 954 395
rect 990 79 1026 420
rect 1062 0 1098 395
rect 1134 0 1170 395
rect 1326 0 1362 395
rect 1398 0 1434 395
rect 1470 79 1506 420
rect 1542 0 1578 395
rect 1614 0 1650 395
rect 2094 0 2130 395
rect 2166 0 2202 395
rect 2238 79 2274 420
rect 2310 0 2346 395
rect 2382 0 2418 395
rect 2574 0 2610 395
rect 2646 0 2682 395
rect 2718 79 2754 420
rect 2790 0 2826 395
rect 2862 0 2898 395
rect 3342 0 3378 395
rect 3414 0 3450 395
rect 3486 79 3522 420
rect 3558 0 3594 395
rect 3630 0 3666 395
rect 3822 0 3858 395
rect 3894 0 3930 395
rect 3966 79 4002 420
rect 4038 0 4074 395
rect 4110 0 4146 395
rect 4590 0 4626 395
rect 4662 0 4698 395
rect 4734 79 4770 420
rect 4806 0 4842 395
rect 4878 0 4914 395
rect 5070 0 5106 395
rect 5142 0 5178 395
rect 5214 79 5250 420
rect 5286 0 5322 395
rect 5358 0 5394 395
rect 5838 0 5874 395
rect 5910 0 5946 395
rect 5982 79 6018 420
rect 6054 0 6090 395
rect 6126 0 6162 395
rect 6318 0 6354 395
rect 6390 0 6426 395
rect 6462 79 6498 420
rect 6534 0 6570 395
rect 6606 0 6642 395
rect 7086 0 7122 395
rect 7158 0 7194 395
rect 7230 79 7266 420
rect 7302 0 7338 395
rect 7374 0 7410 395
rect 7566 0 7602 395
rect 7638 0 7674 395
rect 7710 79 7746 420
rect 7782 0 7818 395
rect 7854 0 7890 395
rect 8334 0 8370 395
rect 8406 0 8442 395
rect 8478 79 8514 420
rect 8550 0 8586 395
rect 8622 0 8658 395
rect 8814 0 8850 395
rect 8886 0 8922 395
rect 8958 79 8994 420
rect 9030 0 9066 395
rect 9102 0 9138 395
rect 9582 0 9618 395
rect 9654 0 9690 395
rect 9726 79 9762 420
rect 9798 0 9834 395
rect 9870 0 9906 395
rect 10062 0 10098 395
rect 10134 0 10170 395
rect 10206 79 10242 420
rect 10278 0 10314 395
rect 10350 0 10386 395
rect 10830 0 10866 395
rect 10902 0 10938 395
rect 10974 79 11010 420
rect 11046 0 11082 395
rect 11118 0 11154 395
rect 11310 0 11346 395
rect 11382 0 11418 395
rect 11454 79 11490 420
rect 11526 0 11562 395
rect 11598 0 11634 395
rect 12078 0 12114 395
rect 12150 0 12186 395
rect 12222 79 12258 420
rect 12294 0 12330 395
rect 12366 0 12402 395
rect 12558 0 12594 395
rect 12630 0 12666 395
rect 12702 79 12738 420
rect 12774 0 12810 395
rect 12846 0 12882 395
rect 13326 0 13362 395
rect 13398 0 13434 395
rect 13470 79 13506 420
rect 13542 0 13578 395
rect 13614 0 13650 395
rect 13806 0 13842 395
rect 13878 0 13914 395
rect 13950 79 13986 420
rect 14022 0 14058 395
rect 14094 0 14130 395
rect 14574 0 14610 395
rect 14646 0 14682 395
rect 14718 79 14754 420
rect 14790 0 14826 395
rect 14862 0 14898 395
rect 15054 0 15090 395
rect 15126 0 15162 395
rect 15198 79 15234 420
rect 15270 0 15306 395
rect 15342 0 15378 395
rect 15822 0 15858 395
rect 15894 0 15930 395
rect 15966 79 16002 420
rect 16038 0 16074 395
rect 16110 0 16146 395
rect 16302 0 16338 395
rect 16374 0 16410 395
rect 16446 79 16482 420
rect 16518 0 16554 395
rect 16590 0 16626 395
rect 17070 0 17106 395
rect 17142 0 17178 395
rect 17214 79 17250 420
rect 17286 0 17322 395
rect 17358 0 17394 395
rect 17550 0 17586 395
rect 17622 0 17658 395
rect 17694 79 17730 420
rect 17766 0 17802 395
rect 17838 0 17874 395
rect 18318 0 18354 395
rect 18390 0 18426 395
rect 18462 79 18498 420
rect 18534 0 18570 395
rect 18606 0 18642 395
rect 18798 0 18834 395
rect 18870 0 18906 395
rect 18942 79 18978 420
rect 19014 0 19050 395
rect 19086 0 19122 395
rect 19566 0 19602 395
rect 19638 0 19674 395
rect 19710 79 19746 420
rect 19782 0 19818 395
rect 19854 0 19890 395
rect 20046 0 20082 395
rect 20118 0 20154 395
rect 20190 79 20226 420
rect 20262 0 20298 395
rect 20334 0 20370 395
rect 20814 0 20850 395
rect 20886 0 20922 395
rect 20958 79 20994 420
rect 21030 0 21066 395
rect 21102 0 21138 395
rect 21294 0 21330 395
rect 21366 0 21402 395
rect 21438 79 21474 420
rect 21510 0 21546 395
rect 21582 0 21618 395
rect 22062 0 22098 395
rect 22134 0 22170 395
rect 22206 79 22242 420
rect 22278 0 22314 395
rect 22350 0 22386 395
rect 22542 0 22578 395
rect 22614 0 22650 395
rect 22686 79 22722 420
rect 22758 0 22794 395
rect 22830 0 22866 395
rect 23310 0 23346 395
rect 23382 0 23418 395
rect 23454 79 23490 420
rect 23526 0 23562 395
rect 23598 0 23634 395
rect 23790 0 23826 395
rect 23862 0 23898 395
rect 23934 79 23970 420
rect 24006 0 24042 395
rect 24078 0 24114 395
rect 24558 0 24594 395
rect 24630 0 24666 395
rect 24702 79 24738 420
rect 24774 0 24810 395
rect 24846 0 24882 395
rect 25038 0 25074 395
rect 25110 0 25146 395
rect 25182 79 25218 420
rect 25254 0 25290 395
rect 25326 0 25362 395
rect 25806 0 25842 395
rect 25878 0 25914 395
rect 25950 79 25986 420
rect 26022 0 26058 395
rect 26094 0 26130 395
rect 26286 0 26322 395
rect 26358 0 26394 395
rect 26430 79 26466 420
rect 26502 0 26538 395
rect 26574 0 26610 395
rect 27054 0 27090 395
rect 27126 0 27162 395
rect 27198 79 27234 420
rect 27270 0 27306 395
rect 27342 0 27378 395
rect 27534 0 27570 395
rect 27606 0 27642 395
rect 27678 79 27714 420
rect 27750 0 27786 395
rect 27822 0 27858 395
rect 28302 0 28338 395
rect 28374 0 28410 395
rect 28446 79 28482 420
rect 28518 0 28554 395
rect 28590 0 28626 395
rect 28782 0 28818 395
rect 28854 0 28890 395
rect 28926 79 28962 420
rect 28998 0 29034 395
rect 29070 0 29106 395
rect 29550 0 29586 395
rect 29622 0 29658 395
rect 29694 79 29730 420
rect 29766 0 29802 395
rect 29838 0 29874 395
rect 30030 0 30066 395
rect 30102 0 30138 395
rect 30174 79 30210 420
rect 30246 0 30282 395
rect 30318 0 30354 395
rect 30798 0 30834 395
rect 30870 0 30906 395
rect 30942 79 30978 420
rect 31014 0 31050 395
rect 31086 0 31122 395
rect 31278 0 31314 395
rect 31350 0 31386 395
rect 31422 79 31458 420
rect 31494 0 31530 395
rect 31566 0 31602 395
rect 32046 0 32082 395
rect 32118 0 32154 395
rect 32190 79 32226 420
rect 32262 0 32298 395
rect 32334 0 32370 395
rect 32526 0 32562 395
rect 32598 0 32634 395
rect 32670 79 32706 420
rect 32742 0 32778 395
rect 32814 0 32850 395
rect 33294 0 33330 395
rect 33366 0 33402 395
rect 33438 79 33474 420
rect 33510 0 33546 395
rect 33582 0 33618 395
rect 33774 0 33810 395
rect 33846 0 33882 395
rect 33918 79 33954 420
rect 33990 0 34026 395
rect 34062 0 34098 395
rect 34542 0 34578 395
rect 34614 0 34650 395
rect 34686 79 34722 420
rect 34758 0 34794 395
rect 34830 0 34866 395
rect 35022 0 35058 395
rect 35094 0 35130 395
rect 35166 79 35202 420
rect 35238 0 35274 395
rect 35310 0 35346 395
rect 35790 0 35826 395
rect 35862 0 35898 395
rect 35934 79 35970 420
rect 36006 0 36042 395
rect 36078 0 36114 395
rect 36270 0 36306 395
rect 36342 0 36378 395
rect 36414 79 36450 420
rect 36486 0 36522 395
rect 36558 0 36594 395
rect 37038 0 37074 395
rect 37110 0 37146 395
rect 37182 79 37218 420
rect 37254 0 37290 395
rect 37326 0 37362 395
rect 37518 0 37554 395
rect 37590 0 37626 395
rect 37662 79 37698 420
rect 37734 0 37770 395
rect 37806 0 37842 395
rect 38286 0 38322 395
rect 38358 0 38394 395
rect 38430 79 38466 420
rect 38502 0 38538 395
rect 38574 0 38610 395
rect 38766 0 38802 395
rect 38838 0 38874 395
rect 38910 79 38946 420
rect 38982 0 39018 395
rect 39054 0 39090 395
rect 39534 0 39570 395
rect 39606 0 39642 395
rect 39678 79 39714 420
rect 39750 0 39786 395
rect 39822 0 39858 395
rect 40014 0 40050 395
rect 40086 0 40122 395
rect 40158 79 40194 420
rect 40230 0 40266 395
rect 40302 0 40338 395
rect 40782 0 40818 395
rect 40854 0 40890 395
rect 40926 79 40962 420
rect 40998 0 41034 395
rect 41070 0 41106 395
rect 41262 0 41298 395
rect 41334 0 41370 395
rect 41406 79 41442 420
rect 41478 0 41514 395
rect 41550 0 41586 395
rect 42030 0 42066 395
rect 42102 0 42138 395
rect 42174 79 42210 420
rect 42246 0 42282 395
rect 42318 0 42354 395
rect 42510 0 42546 395
rect 42582 0 42618 395
rect 42654 79 42690 420
rect 42726 0 42762 395
rect 42798 0 42834 395
rect 43278 0 43314 395
rect 43350 0 43386 395
rect 43422 79 43458 420
rect 43494 0 43530 395
rect 43566 0 43602 395
rect 43758 0 43794 395
rect 43830 0 43866 395
rect 43902 79 43938 420
rect 43974 0 44010 395
rect 44046 0 44082 395
rect 44526 0 44562 395
rect 44598 0 44634 395
rect 44670 79 44706 420
rect 44742 0 44778 395
rect 44814 0 44850 395
rect 45006 0 45042 395
rect 45078 0 45114 395
rect 45150 79 45186 420
rect 45222 0 45258 395
rect 45294 0 45330 395
rect 45774 0 45810 395
rect 45846 0 45882 395
rect 45918 79 45954 420
rect 45990 0 46026 395
rect 46062 0 46098 395
rect 46254 0 46290 395
rect 46326 0 46362 395
rect 46398 79 46434 420
rect 46470 0 46506 395
rect 46542 0 46578 395
rect 47022 0 47058 395
rect 47094 0 47130 395
rect 47166 79 47202 420
rect 47238 0 47274 395
rect 47310 0 47346 395
rect 47502 0 47538 395
rect 47574 0 47610 395
rect 47646 79 47682 420
rect 47718 0 47754 395
rect 47790 0 47826 395
rect 48270 0 48306 395
rect 48342 0 48378 395
rect 48414 79 48450 420
rect 48486 0 48522 395
rect 48558 0 48594 395
rect 48750 0 48786 395
rect 48822 0 48858 395
rect 48894 79 48930 420
rect 48966 0 49002 395
rect 49038 0 49074 395
rect 49518 0 49554 395
rect 49590 0 49626 395
rect 49662 79 49698 420
rect 49734 0 49770 395
rect 49806 0 49842 395
rect 49998 0 50034 395
rect 50070 0 50106 395
rect 50142 79 50178 420
rect 50214 0 50250 395
rect 50286 0 50322 395
rect 50766 0 50802 395
rect 50838 0 50874 395
rect 50910 79 50946 420
rect 50982 0 51018 395
rect 51054 0 51090 395
rect 51246 0 51282 395
rect 51318 0 51354 395
rect 51390 79 51426 420
rect 51462 0 51498 395
rect 51534 0 51570 395
rect 52014 0 52050 395
rect 52086 0 52122 395
rect 52158 79 52194 420
rect 52230 0 52266 395
rect 52302 0 52338 395
rect 52494 0 52530 395
rect 52566 0 52602 395
rect 52638 79 52674 420
rect 52710 0 52746 395
rect 52782 0 52818 395
rect 53262 0 53298 395
rect 53334 0 53370 395
rect 53406 79 53442 420
rect 53478 0 53514 395
rect 53550 0 53586 395
rect 53742 0 53778 395
rect 53814 0 53850 395
rect 53886 79 53922 420
rect 53958 0 53994 395
rect 54030 0 54066 395
rect 54510 0 54546 395
rect 54582 0 54618 395
rect 54654 79 54690 420
rect 54726 0 54762 395
rect 54798 0 54834 395
rect 54990 0 55026 395
rect 55062 0 55098 395
rect 55134 79 55170 420
rect 55206 0 55242 395
rect 55278 0 55314 395
rect 55758 0 55794 395
rect 55830 0 55866 395
rect 55902 79 55938 420
rect 55974 0 56010 395
rect 56046 0 56082 395
rect 56238 0 56274 395
rect 56310 0 56346 395
rect 56382 79 56418 420
rect 56454 0 56490 395
rect 56526 0 56562 395
rect 57006 0 57042 395
rect 57078 0 57114 395
rect 57150 79 57186 420
rect 57222 0 57258 395
rect 57294 0 57330 395
rect 57486 0 57522 395
rect 57558 0 57594 395
rect 57630 79 57666 420
rect 57702 0 57738 395
rect 57774 0 57810 395
rect 58254 0 58290 395
rect 58326 0 58362 395
rect 58398 79 58434 420
rect 58470 0 58506 395
rect 58542 0 58578 395
rect 58734 0 58770 395
rect 58806 0 58842 395
rect 58878 79 58914 420
rect 58950 0 58986 395
rect 59022 0 59058 395
rect 59502 0 59538 395
rect 59574 0 59610 395
rect 59646 79 59682 420
rect 59718 0 59754 395
rect 59790 0 59826 395
rect 59982 0 60018 395
rect 60054 0 60090 395
rect 60126 79 60162 420
rect 60198 0 60234 395
rect 60270 0 60306 395
rect 60750 0 60786 395
rect 60822 0 60858 395
rect 60894 79 60930 420
rect 60966 0 61002 395
rect 61038 0 61074 395
rect 61230 0 61266 395
rect 61302 0 61338 395
rect 61374 79 61410 420
rect 61446 0 61482 395
rect 61518 0 61554 395
rect 61998 0 62034 395
rect 62070 0 62106 395
rect 62142 79 62178 420
rect 62214 0 62250 395
rect 62286 0 62322 395
rect 62478 0 62514 395
rect 62550 0 62586 395
rect 62622 79 62658 420
rect 62694 0 62730 395
rect 62766 0 62802 395
rect 63246 0 63282 395
rect 63318 0 63354 395
rect 63390 79 63426 420
rect 63462 0 63498 395
rect 63534 0 63570 395
rect 63726 0 63762 395
rect 63798 0 63834 395
rect 63870 79 63906 420
rect 63942 0 63978 395
rect 64014 0 64050 395
rect 64494 0 64530 395
rect 64566 0 64602 395
rect 64638 79 64674 420
rect 64710 0 64746 395
rect 64782 0 64818 395
rect 64974 0 65010 395
rect 65046 0 65082 395
rect 65118 79 65154 420
rect 65190 0 65226 395
rect 65262 0 65298 395
rect 65742 0 65778 395
rect 65814 0 65850 395
rect 65886 79 65922 420
rect 65958 0 65994 395
rect 66030 0 66066 395
rect 66222 0 66258 395
rect 66294 0 66330 395
rect 66366 79 66402 420
rect 66438 0 66474 395
rect 66510 0 66546 395
rect 66990 0 67026 395
rect 67062 0 67098 395
rect 67134 79 67170 420
rect 67206 0 67242 395
rect 67278 0 67314 395
rect 67470 0 67506 395
rect 67542 0 67578 395
rect 67614 79 67650 420
rect 67686 0 67722 395
rect 67758 0 67794 395
rect 68238 0 68274 395
rect 68310 0 68346 395
rect 68382 79 68418 420
rect 68454 0 68490 395
rect 68526 0 68562 395
rect 68718 0 68754 395
rect 68790 0 68826 395
rect 68862 79 68898 420
rect 68934 0 68970 395
rect 69006 0 69042 395
rect 69486 0 69522 395
rect 69558 0 69594 395
rect 69630 79 69666 420
rect 69702 0 69738 395
rect 69774 0 69810 395
rect 69966 0 70002 395
rect 70038 0 70074 395
rect 70110 79 70146 420
rect 70182 0 70218 395
rect 70254 0 70290 395
rect 70734 0 70770 395
rect 70806 0 70842 395
rect 70878 79 70914 420
rect 70950 0 70986 395
rect 71022 0 71058 395
rect 71214 0 71250 395
rect 71286 0 71322 395
rect 71358 79 71394 420
rect 71430 0 71466 395
rect 71502 0 71538 395
rect 71982 0 72018 395
rect 72054 0 72090 395
rect 72126 79 72162 420
rect 72198 0 72234 395
rect 72270 0 72306 395
rect 72462 0 72498 395
rect 72534 0 72570 395
rect 72606 79 72642 420
rect 72678 0 72714 395
rect 72750 0 72786 395
rect 73230 0 73266 395
rect 73302 0 73338 395
rect 73374 79 73410 420
rect 73446 0 73482 395
rect 73518 0 73554 395
rect 73710 0 73746 395
rect 73782 0 73818 395
rect 73854 79 73890 420
rect 73926 0 73962 395
rect 73998 0 74034 395
rect 74478 0 74514 395
rect 74550 0 74586 395
rect 74622 79 74658 420
rect 74694 0 74730 395
rect 74766 0 74802 395
rect 74958 0 74994 395
rect 75030 0 75066 395
rect 75102 79 75138 420
rect 75174 0 75210 395
rect 75246 0 75282 395
rect 75726 0 75762 395
rect 75798 0 75834 395
rect 75870 79 75906 420
rect 75942 0 75978 395
rect 76014 0 76050 395
rect 76206 0 76242 395
rect 76278 0 76314 395
rect 76350 79 76386 420
rect 76422 0 76458 395
rect 76494 0 76530 395
rect 76974 0 77010 395
rect 77046 0 77082 395
rect 77118 79 77154 420
rect 77190 0 77226 395
rect 77262 0 77298 395
rect 77454 0 77490 395
rect 77526 0 77562 395
rect 77598 79 77634 420
rect 77670 0 77706 395
rect 77742 0 77778 395
rect 78222 0 78258 395
rect 78294 0 78330 395
rect 78366 79 78402 420
rect 78438 0 78474 395
rect 78510 0 78546 395
rect 78702 0 78738 395
rect 78774 0 78810 395
rect 78846 79 78882 420
rect 78918 0 78954 395
rect 78990 0 79026 395
rect 79470 0 79506 395
rect 79542 0 79578 395
rect 79614 79 79650 420
rect 79686 0 79722 395
rect 79758 0 79794 395
<< metal2 >>
rect 0 323 79872 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 5178 199 5286 275
rect 5946 199 6054 275
rect 6426 199 6534 275
rect 7194 199 7302 275
rect 7674 199 7782 275
rect 8442 199 8550 275
rect 8922 199 9030 275
rect 9690 199 9798 275
rect 10170 199 10278 275
rect 10938 199 11046 275
rect 11418 199 11526 275
rect 12186 199 12294 275
rect 12666 199 12774 275
rect 13434 199 13542 275
rect 13914 199 14022 275
rect 14682 199 14790 275
rect 15162 199 15270 275
rect 15930 199 16038 275
rect 16410 199 16518 275
rect 17178 199 17286 275
rect 17658 199 17766 275
rect 18426 199 18534 275
rect 18906 199 19014 275
rect 19674 199 19782 275
rect 20154 199 20262 275
rect 20922 199 21030 275
rect 21402 199 21510 275
rect 22170 199 22278 275
rect 22650 199 22758 275
rect 23418 199 23526 275
rect 23898 199 24006 275
rect 24666 199 24774 275
rect 25146 199 25254 275
rect 25914 199 26022 275
rect 26394 199 26502 275
rect 27162 199 27270 275
rect 27642 199 27750 275
rect 28410 199 28518 275
rect 28890 199 28998 275
rect 29658 199 29766 275
rect 30138 199 30246 275
rect 30906 199 31014 275
rect 31386 199 31494 275
rect 32154 199 32262 275
rect 32634 199 32742 275
rect 33402 199 33510 275
rect 33882 199 33990 275
rect 34650 199 34758 275
rect 35130 199 35238 275
rect 35898 199 36006 275
rect 36378 199 36486 275
rect 37146 199 37254 275
rect 37626 199 37734 275
rect 38394 199 38502 275
rect 38874 199 38982 275
rect 39642 199 39750 275
rect 40122 199 40230 275
rect 40890 199 40998 275
rect 41370 199 41478 275
rect 42138 199 42246 275
rect 42618 199 42726 275
rect 43386 199 43494 275
rect 43866 199 43974 275
rect 44634 199 44742 275
rect 45114 199 45222 275
rect 45882 199 45990 275
rect 46362 199 46470 275
rect 47130 199 47238 275
rect 47610 199 47718 275
rect 48378 199 48486 275
rect 48858 199 48966 275
rect 49626 199 49734 275
rect 50106 199 50214 275
rect 50874 199 50982 275
rect 51354 199 51462 275
rect 52122 199 52230 275
rect 52602 199 52710 275
rect 53370 199 53478 275
rect 53850 199 53958 275
rect 54618 199 54726 275
rect 55098 199 55206 275
rect 55866 199 55974 275
rect 56346 199 56454 275
rect 57114 199 57222 275
rect 57594 199 57702 275
rect 58362 199 58470 275
rect 58842 199 58950 275
rect 59610 199 59718 275
rect 60090 199 60198 275
rect 60858 199 60966 275
rect 61338 199 61446 275
rect 62106 199 62214 275
rect 62586 199 62694 275
rect 63354 199 63462 275
rect 63834 199 63942 275
rect 64602 199 64710 275
rect 65082 199 65190 275
rect 65850 199 65958 275
rect 66330 199 66438 275
rect 67098 199 67206 275
rect 67578 199 67686 275
rect 68346 199 68454 275
rect 68826 199 68934 275
rect 69594 199 69702 275
rect 70074 199 70182 275
rect 70842 199 70950 275
rect 71322 199 71430 275
rect 72090 199 72198 275
rect 72570 199 72678 275
rect 73338 199 73446 275
rect 73818 199 73926 275
rect 74586 199 74694 275
rect 75066 199 75174 275
rect 75834 199 75942 275
rect 76314 199 76422 275
rect 77082 199 77190 275
rect 77562 199 77670 275
rect 78330 199 78438 275
rect 78810 199 78918 275
rect 79578 199 79686 275
rect 0 103 79872 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
rect 5178 -55 5286 55
rect 5946 -55 6054 55
rect 6426 -55 6534 55
rect 7194 -55 7302 55
rect 7674 -55 7782 55
rect 8442 -55 8550 55
rect 8922 -55 9030 55
rect 9690 -55 9798 55
rect 10170 -55 10278 55
rect 10938 -55 11046 55
rect 11418 -55 11526 55
rect 12186 -55 12294 55
rect 12666 -55 12774 55
rect 13434 -55 13542 55
rect 13914 -55 14022 55
rect 14682 -55 14790 55
rect 15162 -55 15270 55
rect 15930 -55 16038 55
rect 16410 -55 16518 55
rect 17178 -55 17286 55
rect 17658 -55 17766 55
rect 18426 -55 18534 55
rect 18906 -55 19014 55
rect 19674 -55 19782 55
rect 20154 -55 20262 55
rect 20922 -55 21030 55
rect 21402 -55 21510 55
rect 22170 -55 22278 55
rect 22650 -55 22758 55
rect 23418 -55 23526 55
rect 23898 -55 24006 55
rect 24666 -55 24774 55
rect 25146 -55 25254 55
rect 25914 -55 26022 55
rect 26394 -55 26502 55
rect 27162 -55 27270 55
rect 27642 -55 27750 55
rect 28410 -55 28518 55
rect 28890 -55 28998 55
rect 29658 -55 29766 55
rect 30138 -55 30246 55
rect 30906 -55 31014 55
rect 31386 -55 31494 55
rect 32154 -55 32262 55
rect 32634 -55 32742 55
rect 33402 -55 33510 55
rect 33882 -55 33990 55
rect 34650 -55 34758 55
rect 35130 -55 35238 55
rect 35898 -55 36006 55
rect 36378 -55 36486 55
rect 37146 -55 37254 55
rect 37626 -55 37734 55
rect 38394 -55 38502 55
rect 38874 -55 38982 55
rect 39642 -55 39750 55
rect 40122 -55 40230 55
rect 40890 -55 40998 55
rect 41370 -55 41478 55
rect 42138 -55 42246 55
rect 42618 -55 42726 55
rect 43386 -55 43494 55
rect 43866 -55 43974 55
rect 44634 -55 44742 55
rect 45114 -55 45222 55
rect 45882 -55 45990 55
rect 46362 -55 46470 55
rect 47130 -55 47238 55
rect 47610 -55 47718 55
rect 48378 -55 48486 55
rect 48858 -55 48966 55
rect 49626 -55 49734 55
rect 50106 -55 50214 55
rect 50874 -55 50982 55
rect 51354 -55 51462 55
rect 52122 -55 52230 55
rect 52602 -55 52710 55
rect 53370 -55 53478 55
rect 53850 -55 53958 55
rect 54618 -55 54726 55
rect 55098 -55 55206 55
rect 55866 -55 55974 55
rect 56346 -55 56454 55
rect 57114 -55 57222 55
rect 57594 -55 57702 55
rect 58362 -55 58470 55
rect 58842 -55 58950 55
rect 59610 -55 59718 55
rect 60090 -55 60198 55
rect 60858 -55 60966 55
rect 61338 -55 61446 55
rect 62106 -55 62214 55
rect 62586 -55 62694 55
rect 63354 -55 63462 55
rect 63834 -55 63942 55
rect 64602 -55 64710 55
rect 65082 -55 65190 55
rect 65850 -55 65958 55
rect 66330 -55 66438 55
rect 67098 -55 67206 55
rect 67578 -55 67686 55
rect 68346 -55 68454 55
rect 68826 -55 68934 55
rect 69594 -55 69702 55
rect 70074 -55 70182 55
rect 70842 -55 70950 55
rect 71322 -55 71430 55
rect 72090 -55 72198 55
rect 72570 -55 72678 55
rect 73338 -55 73446 55
rect 73818 -55 73926 55
rect 74586 -55 74694 55
rect 75066 -55 75174 55
rect 75834 -55 75942 55
rect 76314 -55 76422 55
rect 77082 -55 77190 55
rect 77562 -55 77670 55
rect 78330 -55 78438 55
rect 78810 -55 78918 55
rect 79578 -55 79686 55
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_127
timestamp 1624494425
transform 1 0 0 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_126
timestamp 1624494425
transform -1 0 1248 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_125
timestamp 1624494425
transform 1 0 1248 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_124
timestamp 1624494425
transform -1 0 2496 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_123
timestamp 1624494425
transform 1 0 2496 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_122
timestamp 1624494425
transform -1 0 3744 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_121
timestamp 1624494425
transform 1 0 3744 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_120
timestamp 1624494425
transform -1 0 4992 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_119
timestamp 1624494425
transform 1 0 4992 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_118
timestamp 1624494425
transform -1 0 6240 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_117
timestamp 1624494425
transform 1 0 6240 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_116
timestamp 1624494425
transform -1 0 7488 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_115
timestamp 1624494425
transform 1 0 7488 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_114
timestamp 1624494425
transform -1 0 8736 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_113
timestamp 1624494425
transform 1 0 8736 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_112
timestamp 1624494425
transform -1 0 9984 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_111
timestamp 1624494425
transform 1 0 9984 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_110
timestamp 1624494425
transform -1 0 11232 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_109
timestamp 1624494425
transform 1 0 11232 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_108
timestamp 1624494425
transform -1 0 12480 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_107
timestamp 1624494425
transform 1 0 12480 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_106
timestamp 1624494425
transform -1 0 13728 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_105
timestamp 1624494425
transform 1 0 13728 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_104
timestamp 1624494425
transform -1 0 14976 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_103
timestamp 1624494425
transform 1 0 14976 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_102
timestamp 1624494425
transform -1 0 16224 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_101
timestamp 1624494425
transform 1 0 16224 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_100
timestamp 1624494425
transform -1 0 17472 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_99
timestamp 1624494425
transform 1 0 17472 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_98
timestamp 1624494425
transform -1 0 18720 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_97
timestamp 1624494425
transform 1 0 18720 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_96
timestamp 1624494425
transform -1 0 19968 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_95
timestamp 1624494425
transform 1 0 19968 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_94
timestamp 1624494425
transform -1 0 21216 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_93
timestamp 1624494425
transform 1 0 21216 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_92
timestamp 1624494425
transform -1 0 22464 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_91
timestamp 1624494425
transform 1 0 22464 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_90
timestamp 1624494425
transform -1 0 23712 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_89
timestamp 1624494425
transform 1 0 23712 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_88
timestamp 1624494425
transform -1 0 24960 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_87
timestamp 1624494425
transform 1 0 24960 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_86
timestamp 1624494425
transform -1 0 26208 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_85
timestamp 1624494425
transform 1 0 26208 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_84
timestamp 1624494425
transform -1 0 27456 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_83
timestamp 1624494425
transform 1 0 27456 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_82
timestamp 1624494425
transform -1 0 28704 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_81
timestamp 1624494425
transform 1 0 28704 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_80
timestamp 1624494425
transform -1 0 29952 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_79
timestamp 1624494425
transform 1 0 29952 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_78
timestamp 1624494425
transform -1 0 31200 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_77
timestamp 1624494425
transform 1 0 31200 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_76
timestamp 1624494425
transform -1 0 32448 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_75
timestamp 1624494425
transform 1 0 32448 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_74
timestamp 1624494425
transform -1 0 33696 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_73
timestamp 1624494425
transform 1 0 33696 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_72
timestamp 1624494425
transform -1 0 34944 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_71
timestamp 1624494425
transform 1 0 34944 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_70
timestamp 1624494425
transform -1 0 36192 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_69
timestamp 1624494425
transform 1 0 36192 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_68
timestamp 1624494425
transform -1 0 37440 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_67
timestamp 1624494425
transform 1 0 37440 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_66
timestamp 1624494425
transform -1 0 38688 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_65
timestamp 1624494425
transform 1 0 38688 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_64
timestamp 1624494425
transform -1 0 39936 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_63
timestamp 1624494425
transform 1 0 39936 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_62
timestamp 1624494425
transform -1 0 41184 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_61
timestamp 1624494425
transform 1 0 41184 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_60
timestamp 1624494425
transform -1 0 42432 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_59
timestamp 1624494425
transform 1 0 42432 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_58
timestamp 1624494425
transform -1 0 43680 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_57
timestamp 1624494425
transform 1 0 43680 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_56
timestamp 1624494425
transform -1 0 44928 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_55
timestamp 1624494425
transform 1 0 44928 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_54
timestamp 1624494425
transform -1 0 46176 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_53
timestamp 1624494425
transform 1 0 46176 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_52
timestamp 1624494425
transform -1 0 47424 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_51
timestamp 1624494425
transform 1 0 47424 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_50
timestamp 1624494425
transform -1 0 48672 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_49
timestamp 1624494425
transform 1 0 48672 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_48
timestamp 1624494425
transform -1 0 49920 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_47
timestamp 1624494425
transform 1 0 49920 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_46
timestamp 1624494425
transform -1 0 51168 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_45
timestamp 1624494425
transform 1 0 51168 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_44
timestamp 1624494425
transform -1 0 52416 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_43
timestamp 1624494425
transform 1 0 52416 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_42
timestamp 1624494425
transform -1 0 53664 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_41
timestamp 1624494425
transform 1 0 53664 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_40
timestamp 1624494425
transform -1 0 54912 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_39
timestamp 1624494425
transform 1 0 54912 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_38
timestamp 1624494425
transform -1 0 56160 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_37
timestamp 1624494425
transform 1 0 56160 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_36
timestamp 1624494425
transform -1 0 57408 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_35
timestamp 1624494425
transform 1 0 57408 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_34
timestamp 1624494425
transform -1 0 58656 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_33
timestamp 1624494425
transform 1 0 58656 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_32
timestamp 1624494425
transform -1 0 59904 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_31
timestamp 1624494425
transform 1 0 59904 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_30
timestamp 1624494425
transform -1 0 61152 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_29
timestamp 1624494425
transform 1 0 61152 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_28
timestamp 1624494425
transform -1 0 62400 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_27
timestamp 1624494425
transform 1 0 62400 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_26
timestamp 1624494425
transform -1 0 63648 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_25
timestamp 1624494425
transform 1 0 63648 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_24
timestamp 1624494425
transform -1 0 64896 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_23
timestamp 1624494425
transform 1 0 64896 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_22
timestamp 1624494425
transform -1 0 66144 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_21
timestamp 1624494425
transform 1 0 66144 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_20
timestamp 1624494425
transform -1 0 67392 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_19
timestamp 1624494425
transform 1 0 67392 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_18
timestamp 1624494425
transform -1 0 68640 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_17
timestamp 1624494425
transform 1 0 68640 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_16
timestamp 1624494425
transform -1 0 69888 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_15
timestamp 1624494425
transform 1 0 69888 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_14
timestamp 1624494425
transform -1 0 71136 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_13
timestamp 1624494425
transform 1 0 71136 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_12
timestamp 1624494425
transform -1 0 72384 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_11
timestamp 1624494425
transform 1 0 72384 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_10
timestamp 1624494425
transform -1 0 73632 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_9
timestamp 1624494425
transform 1 0 73632 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_8
timestamp 1624494425
transform -1 0 74880 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_7
timestamp 1624494425
transform 1 0 74880 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_6
timestamp 1624494425
transform -1 0 76128 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_5
timestamp 1624494425
transform 1 0 76128 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_4
timestamp 1624494425
transform -1 0 77376 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_3
timestamp 1624494425
transform 1 0 77376 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_2
timestamp 1624494425
transform -1 0 78624 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_1
timestamp 1624494425
transform 1 0 78624 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1624494425
transform -1 0 79872 0 1 0
box -42 -105 650 424
<< labels >>
rlabel metal1 s 78 0 114 395 4 bl_0_0
rlabel metal1 s 150 0 186 395 4 br_0_0
rlabel metal1 s 294 0 330 395 4 bl_1_0
rlabel metal1 s 366 0 402 395 4 br_1_0
rlabel metal1 s 1134 0 1170 395 4 bl_0_1
rlabel metal1 s 1062 0 1098 395 4 br_0_1
rlabel metal1 s 918 0 954 395 4 bl_1_1
rlabel metal1 s 846 0 882 395 4 br_1_1
rlabel metal1 s 1326 0 1362 395 4 bl_0_2
rlabel metal1 s 1398 0 1434 395 4 br_0_2
rlabel metal1 s 1542 0 1578 395 4 bl_1_2
rlabel metal1 s 1614 0 1650 395 4 br_1_2
rlabel metal1 s 2382 0 2418 395 4 bl_0_3
rlabel metal1 s 2310 0 2346 395 4 br_0_3
rlabel metal1 s 2166 0 2202 395 4 bl_1_3
rlabel metal1 s 2094 0 2130 395 4 br_1_3
rlabel metal1 s 2574 0 2610 395 4 bl_0_4
rlabel metal1 s 2646 0 2682 395 4 br_0_4
rlabel metal1 s 2790 0 2826 395 4 bl_1_4
rlabel metal1 s 2862 0 2898 395 4 br_1_4
rlabel metal1 s 3630 0 3666 395 4 bl_0_5
rlabel metal1 s 3558 0 3594 395 4 br_0_5
rlabel metal1 s 3414 0 3450 395 4 bl_1_5
rlabel metal1 s 3342 0 3378 395 4 br_1_5
rlabel metal1 s 3822 0 3858 395 4 bl_0_6
rlabel metal1 s 3894 0 3930 395 4 br_0_6
rlabel metal1 s 4038 0 4074 395 4 bl_1_6
rlabel metal1 s 4110 0 4146 395 4 br_1_6
rlabel metal1 s 4878 0 4914 395 4 bl_0_7
rlabel metal1 s 4806 0 4842 395 4 br_0_7
rlabel metal1 s 4662 0 4698 395 4 bl_1_7
rlabel metal1 s 4590 0 4626 395 4 br_1_7
rlabel metal1 s 5070 0 5106 395 4 bl_0_8
rlabel metal1 s 5142 0 5178 395 4 br_0_8
rlabel metal1 s 5286 0 5322 395 4 bl_1_8
rlabel metal1 s 5358 0 5394 395 4 br_1_8
rlabel metal1 s 6126 0 6162 395 4 bl_0_9
rlabel metal1 s 6054 0 6090 395 4 br_0_9
rlabel metal1 s 5910 0 5946 395 4 bl_1_9
rlabel metal1 s 5838 0 5874 395 4 br_1_9
rlabel metal1 s 6318 0 6354 395 4 bl_0_10
rlabel metal1 s 6390 0 6426 395 4 br_0_10
rlabel metal1 s 6534 0 6570 395 4 bl_1_10
rlabel metal1 s 6606 0 6642 395 4 br_1_10
rlabel metal1 s 7374 0 7410 395 4 bl_0_11
rlabel metal1 s 7302 0 7338 395 4 br_0_11
rlabel metal1 s 7158 0 7194 395 4 bl_1_11
rlabel metal1 s 7086 0 7122 395 4 br_1_11
rlabel metal1 s 7566 0 7602 395 4 bl_0_12
rlabel metal1 s 7638 0 7674 395 4 br_0_12
rlabel metal1 s 7782 0 7818 395 4 bl_1_12
rlabel metal1 s 7854 0 7890 395 4 br_1_12
rlabel metal1 s 8622 0 8658 395 4 bl_0_13
rlabel metal1 s 8550 0 8586 395 4 br_0_13
rlabel metal1 s 8406 0 8442 395 4 bl_1_13
rlabel metal1 s 8334 0 8370 395 4 br_1_13
rlabel metal1 s 8814 0 8850 395 4 bl_0_14
rlabel metal1 s 8886 0 8922 395 4 br_0_14
rlabel metal1 s 9030 0 9066 395 4 bl_1_14
rlabel metal1 s 9102 0 9138 395 4 br_1_14
rlabel metal1 s 9870 0 9906 395 4 bl_0_15
rlabel metal1 s 9798 0 9834 395 4 br_0_15
rlabel metal1 s 9654 0 9690 395 4 bl_1_15
rlabel metal1 s 9582 0 9618 395 4 br_1_15
rlabel metal1 s 10062 0 10098 395 4 bl_0_16
rlabel metal1 s 10134 0 10170 395 4 br_0_16
rlabel metal1 s 10278 0 10314 395 4 bl_1_16
rlabel metal1 s 10350 0 10386 395 4 br_1_16
rlabel metal1 s 11118 0 11154 395 4 bl_0_17
rlabel metal1 s 11046 0 11082 395 4 br_0_17
rlabel metal1 s 10902 0 10938 395 4 bl_1_17
rlabel metal1 s 10830 0 10866 395 4 br_1_17
rlabel metal1 s 11310 0 11346 395 4 bl_0_18
rlabel metal1 s 11382 0 11418 395 4 br_0_18
rlabel metal1 s 11526 0 11562 395 4 bl_1_18
rlabel metal1 s 11598 0 11634 395 4 br_1_18
rlabel metal1 s 12366 0 12402 395 4 bl_0_19
rlabel metal1 s 12294 0 12330 395 4 br_0_19
rlabel metal1 s 12150 0 12186 395 4 bl_1_19
rlabel metal1 s 12078 0 12114 395 4 br_1_19
rlabel metal1 s 12558 0 12594 395 4 bl_0_20
rlabel metal1 s 12630 0 12666 395 4 br_0_20
rlabel metal1 s 12774 0 12810 395 4 bl_1_20
rlabel metal1 s 12846 0 12882 395 4 br_1_20
rlabel metal1 s 13614 0 13650 395 4 bl_0_21
rlabel metal1 s 13542 0 13578 395 4 br_0_21
rlabel metal1 s 13398 0 13434 395 4 bl_1_21
rlabel metal1 s 13326 0 13362 395 4 br_1_21
rlabel metal1 s 13806 0 13842 395 4 bl_0_22
rlabel metal1 s 13878 0 13914 395 4 br_0_22
rlabel metal1 s 14022 0 14058 395 4 bl_1_22
rlabel metal1 s 14094 0 14130 395 4 br_1_22
rlabel metal1 s 14862 0 14898 395 4 bl_0_23
rlabel metal1 s 14790 0 14826 395 4 br_0_23
rlabel metal1 s 14646 0 14682 395 4 bl_1_23
rlabel metal1 s 14574 0 14610 395 4 br_1_23
rlabel metal1 s 15054 0 15090 395 4 bl_0_24
rlabel metal1 s 15126 0 15162 395 4 br_0_24
rlabel metal1 s 15270 0 15306 395 4 bl_1_24
rlabel metal1 s 15342 0 15378 395 4 br_1_24
rlabel metal1 s 16110 0 16146 395 4 bl_0_25
rlabel metal1 s 16038 0 16074 395 4 br_0_25
rlabel metal1 s 15894 0 15930 395 4 bl_1_25
rlabel metal1 s 15822 0 15858 395 4 br_1_25
rlabel metal1 s 16302 0 16338 395 4 bl_0_26
rlabel metal1 s 16374 0 16410 395 4 br_0_26
rlabel metal1 s 16518 0 16554 395 4 bl_1_26
rlabel metal1 s 16590 0 16626 395 4 br_1_26
rlabel metal1 s 17358 0 17394 395 4 bl_0_27
rlabel metal1 s 17286 0 17322 395 4 br_0_27
rlabel metal1 s 17142 0 17178 395 4 bl_1_27
rlabel metal1 s 17070 0 17106 395 4 br_1_27
rlabel metal1 s 17550 0 17586 395 4 bl_0_28
rlabel metal1 s 17622 0 17658 395 4 br_0_28
rlabel metal1 s 17766 0 17802 395 4 bl_1_28
rlabel metal1 s 17838 0 17874 395 4 br_1_28
rlabel metal1 s 18606 0 18642 395 4 bl_0_29
rlabel metal1 s 18534 0 18570 395 4 br_0_29
rlabel metal1 s 18390 0 18426 395 4 bl_1_29
rlabel metal1 s 18318 0 18354 395 4 br_1_29
rlabel metal1 s 18798 0 18834 395 4 bl_0_30
rlabel metal1 s 18870 0 18906 395 4 br_0_30
rlabel metal1 s 19014 0 19050 395 4 bl_1_30
rlabel metal1 s 19086 0 19122 395 4 br_1_30
rlabel metal1 s 19854 0 19890 395 4 bl_0_31
rlabel metal1 s 19782 0 19818 395 4 br_0_31
rlabel metal1 s 19638 0 19674 395 4 bl_1_31
rlabel metal1 s 19566 0 19602 395 4 br_1_31
rlabel metal1 s 20046 0 20082 395 4 bl_0_32
rlabel metal1 s 20118 0 20154 395 4 br_0_32
rlabel metal1 s 20262 0 20298 395 4 bl_1_32
rlabel metal1 s 20334 0 20370 395 4 br_1_32
rlabel metal1 s 21102 0 21138 395 4 bl_0_33
rlabel metal1 s 21030 0 21066 395 4 br_0_33
rlabel metal1 s 20886 0 20922 395 4 bl_1_33
rlabel metal1 s 20814 0 20850 395 4 br_1_33
rlabel metal1 s 21294 0 21330 395 4 bl_0_34
rlabel metal1 s 21366 0 21402 395 4 br_0_34
rlabel metal1 s 21510 0 21546 395 4 bl_1_34
rlabel metal1 s 21582 0 21618 395 4 br_1_34
rlabel metal1 s 22350 0 22386 395 4 bl_0_35
rlabel metal1 s 22278 0 22314 395 4 br_0_35
rlabel metal1 s 22134 0 22170 395 4 bl_1_35
rlabel metal1 s 22062 0 22098 395 4 br_1_35
rlabel metal1 s 22542 0 22578 395 4 bl_0_36
rlabel metal1 s 22614 0 22650 395 4 br_0_36
rlabel metal1 s 22758 0 22794 395 4 bl_1_36
rlabel metal1 s 22830 0 22866 395 4 br_1_36
rlabel metal1 s 23598 0 23634 395 4 bl_0_37
rlabel metal1 s 23526 0 23562 395 4 br_0_37
rlabel metal1 s 23382 0 23418 395 4 bl_1_37
rlabel metal1 s 23310 0 23346 395 4 br_1_37
rlabel metal1 s 23790 0 23826 395 4 bl_0_38
rlabel metal1 s 23862 0 23898 395 4 br_0_38
rlabel metal1 s 24006 0 24042 395 4 bl_1_38
rlabel metal1 s 24078 0 24114 395 4 br_1_38
rlabel metal1 s 24846 0 24882 395 4 bl_0_39
rlabel metal1 s 24774 0 24810 395 4 br_0_39
rlabel metal1 s 24630 0 24666 395 4 bl_1_39
rlabel metal1 s 24558 0 24594 395 4 br_1_39
rlabel metal1 s 25038 0 25074 395 4 bl_0_40
rlabel metal1 s 25110 0 25146 395 4 br_0_40
rlabel metal1 s 25254 0 25290 395 4 bl_1_40
rlabel metal1 s 25326 0 25362 395 4 br_1_40
rlabel metal1 s 26094 0 26130 395 4 bl_0_41
rlabel metal1 s 26022 0 26058 395 4 br_0_41
rlabel metal1 s 25878 0 25914 395 4 bl_1_41
rlabel metal1 s 25806 0 25842 395 4 br_1_41
rlabel metal1 s 26286 0 26322 395 4 bl_0_42
rlabel metal1 s 26358 0 26394 395 4 br_0_42
rlabel metal1 s 26502 0 26538 395 4 bl_1_42
rlabel metal1 s 26574 0 26610 395 4 br_1_42
rlabel metal1 s 27342 0 27378 395 4 bl_0_43
rlabel metal1 s 27270 0 27306 395 4 br_0_43
rlabel metal1 s 27126 0 27162 395 4 bl_1_43
rlabel metal1 s 27054 0 27090 395 4 br_1_43
rlabel metal1 s 27534 0 27570 395 4 bl_0_44
rlabel metal1 s 27606 0 27642 395 4 br_0_44
rlabel metal1 s 27750 0 27786 395 4 bl_1_44
rlabel metal1 s 27822 0 27858 395 4 br_1_44
rlabel metal1 s 28590 0 28626 395 4 bl_0_45
rlabel metal1 s 28518 0 28554 395 4 br_0_45
rlabel metal1 s 28374 0 28410 395 4 bl_1_45
rlabel metal1 s 28302 0 28338 395 4 br_1_45
rlabel metal1 s 28782 0 28818 395 4 bl_0_46
rlabel metal1 s 28854 0 28890 395 4 br_0_46
rlabel metal1 s 28998 0 29034 395 4 bl_1_46
rlabel metal1 s 29070 0 29106 395 4 br_1_46
rlabel metal1 s 29838 0 29874 395 4 bl_0_47
rlabel metal1 s 29766 0 29802 395 4 br_0_47
rlabel metal1 s 29622 0 29658 395 4 bl_1_47
rlabel metal1 s 29550 0 29586 395 4 br_1_47
rlabel metal1 s 30030 0 30066 395 4 bl_0_48
rlabel metal1 s 30102 0 30138 395 4 br_0_48
rlabel metal1 s 30246 0 30282 395 4 bl_1_48
rlabel metal1 s 30318 0 30354 395 4 br_1_48
rlabel metal1 s 31086 0 31122 395 4 bl_0_49
rlabel metal1 s 31014 0 31050 395 4 br_0_49
rlabel metal1 s 30870 0 30906 395 4 bl_1_49
rlabel metal1 s 30798 0 30834 395 4 br_1_49
rlabel metal1 s 31278 0 31314 395 4 bl_0_50
rlabel metal1 s 31350 0 31386 395 4 br_0_50
rlabel metal1 s 31494 0 31530 395 4 bl_1_50
rlabel metal1 s 31566 0 31602 395 4 br_1_50
rlabel metal1 s 32334 0 32370 395 4 bl_0_51
rlabel metal1 s 32262 0 32298 395 4 br_0_51
rlabel metal1 s 32118 0 32154 395 4 bl_1_51
rlabel metal1 s 32046 0 32082 395 4 br_1_51
rlabel metal1 s 32526 0 32562 395 4 bl_0_52
rlabel metal1 s 32598 0 32634 395 4 br_0_52
rlabel metal1 s 32742 0 32778 395 4 bl_1_52
rlabel metal1 s 32814 0 32850 395 4 br_1_52
rlabel metal1 s 33582 0 33618 395 4 bl_0_53
rlabel metal1 s 33510 0 33546 395 4 br_0_53
rlabel metal1 s 33366 0 33402 395 4 bl_1_53
rlabel metal1 s 33294 0 33330 395 4 br_1_53
rlabel metal1 s 33774 0 33810 395 4 bl_0_54
rlabel metal1 s 33846 0 33882 395 4 br_0_54
rlabel metal1 s 33990 0 34026 395 4 bl_1_54
rlabel metal1 s 34062 0 34098 395 4 br_1_54
rlabel metal1 s 34830 0 34866 395 4 bl_0_55
rlabel metal1 s 34758 0 34794 395 4 br_0_55
rlabel metal1 s 34614 0 34650 395 4 bl_1_55
rlabel metal1 s 34542 0 34578 395 4 br_1_55
rlabel metal1 s 35022 0 35058 395 4 bl_0_56
rlabel metal1 s 35094 0 35130 395 4 br_0_56
rlabel metal1 s 35238 0 35274 395 4 bl_1_56
rlabel metal1 s 35310 0 35346 395 4 br_1_56
rlabel metal1 s 36078 0 36114 395 4 bl_0_57
rlabel metal1 s 36006 0 36042 395 4 br_0_57
rlabel metal1 s 35862 0 35898 395 4 bl_1_57
rlabel metal1 s 35790 0 35826 395 4 br_1_57
rlabel metal1 s 36270 0 36306 395 4 bl_0_58
rlabel metal1 s 36342 0 36378 395 4 br_0_58
rlabel metal1 s 36486 0 36522 395 4 bl_1_58
rlabel metal1 s 36558 0 36594 395 4 br_1_58
rlabel metal1 s 37326 0 37362 395 4 bl_0_59
rlabel metal1 s 37254 0 37290 395 4 br_0_59
rlabel metal1 s 37110 0 37146 395 4 bl_1_59
rlabel metal1 s 37038 0 37074 395 4 br_1_59
rlabel metal1 s 37518 0 37554 395 4 bl_0_60
rlabel metal1 s 37590 0 37626 395 4 br_0_60
rlabel metal1 s 37734 0 37770 395 4 bl_1_60
rlabel metal1 s 37806 0 37842 395 4 br_1_60
rlabel metal1 s 38574 0 38610 395 4 bl_0_61
rlabel metal1 s 38502 0 38538 395 4 br_0_61
rlabel metal1 s 38358 0 38394 395 4 bl_1_61
rlabel metal1 s 38286 0 38322 395 4 br_1_61
rlabel metal1 s 38766 0 38802 395 4 bl_0_62
rlabel metal1 s 38838 0 38874 395 4 br_0_62
rlabel metal1 s 38982 0 39018 395 4 bl_1_62
rlabel metal1 s 39054 0 39090 395 4 br_1_62
rlabel metal1 s 39822 0 39858 395 4 bl_0_63
rlabel metal1 s 39750 0 39786 395 4 br_0_63
rlabel metal1 s 39606 0 39642 395 4 bl_1_63
rlabel metal1 s 39534 0 39570 395 4 br_1_63
rlabel metal1 s 40014 0 40050 395 4 bl_0_64
rlabel metal1 s 40086 0 40122 395 4 br_0_64
rlabel metal1 s 40230 0 40266 395 4 bl_1_64
rlabel metal1 s 40302 0 40338 395 4 br_1_64
rlabel metal1 s 41070 0 41106 395 4 bl_0_65
rlabel metal1 s 40998 0 41034 395 4 br_0_65
rlabel metal1 s 40854 0 40890 395 4 bl_1_65
rlabel metal1 s 40782 0 40818 395 4 br_1_65
rlabel metal1 s 41262 0 41298 395 4 bl_0_66
rlabel metal1 s 41334 0 41370 395 4 br_0_66
rlabel metal1 s 41478 0 41514 395 4 bl_1_66
rlabel metal1 s 41550 0 41586 395 4 br_1_66
rlabel metal1 s 42318 0 42354 395 4 bl_0_67
rlabel metal1 s 42246 0 42282 395 4 br_0_67
rlabel metal1 s 42102 0 42138 395 4 bl_1_67
rlabel metal1 s 42030 0 42066 395 4 br_1_67
rlabel metal1 s 42510 0 42546 395 4 bl_0_68
rlabel metal1 s 42582 0 42618 395 4 br_0_68
rlabel metal1 s 42726 0 42762 395 4 bl_1_68
rlabel metal1 s 42798 0 42834 395 4 br_1_68
rlabel metal1 s 43566 0 43602 395 4 bl_0_69
rlabel metal1 s 43494 0 43530 395 4 br_0_69
rlabel metal1 s 43350 0 43386 395 4 bl_1_69
rlabel metal1 s 43278 0 43314 395 4 br_1_69
rlabel metal1 s 43758 0 43794 395 4 bl_0_70
rlabel metal1 s 43830 0 43866 395 4 br_0_70
rlabel metal1 s 43974 0 44010 395 4 bl_1_70
rlabel metal1 s 44046 0 44082 395 4 br_1_70
rlabel metal1 s 44814 0 44850 395 4 bl_0_71
rlabel metal1 s 44742 0 44778 395 4 br_0_71
rlabel metal1 s 44598 0 44634 395 4 bl_1_71
rlabel metal1 s 44526 0 44562 395 4 br_1_71
rlabel metal1 s 45006 0 45042 395 4 bl_0_72
rlabel metal1 s 45078 0 45114 395 4 br_0_72
rlabel metal1 s 45222 0 45258 395 4 bl_1_72
rlabel metal1 s 45294 0 45330 395 4 br_1_72
rlabel metal1 s 46062 0 46098 395 4 bl_0_73
rlabel metal1 s 45990 0 46026 395 4 br_0_73
rlabel metal1 s 45846 0 45882 395 4 bl_1_73
rlabel metal1 s 45774 0 45810 395 4 br_1_73
rlabel metal1 s 46254 0 46290 395 4 bl_0_74
rlabel metal1 s 46326 0 46362 395 4 br_0_74
rlabel metal1 s 46470 0 46506 395 4 bl_1_74
rlabel metal1 s 46542 0 46578 395 4 br_1_74
rlabel metal1 s 47310 0 47346 395 4 bl_0_75
rlabel metal1 s 47238 0 47274 395 4 br_0_75
rlabel metal1 s 47094 0 47130 395 4 bl_1_75
rlabel metal1 s 47022 0 47058 395 4 br_1_75
rlabel metal1 s 47502 0 47538 395 4 bl_0_76
rlabel metal1 s 47574 0 47610 395 4 br_0_76
rlabel metal1 s 47718 0 47754 395 4 bl_1_76
rlabel metal1 s 47790 0 47826 395 4 br_1_76
rlabel metal1 s 48558 0 48594 395 4 bl_0_77
rlabel metal1 s 48486 0 48522 395 4 br_0_77
rlabel metal1 s 48342 0 48378 395 4 bl_1_77
rlabel metal1 s 48270 0 48306 395 4 br_1_77
rlabel metal1 s 48750 0 48786 395 4 bl_0_78
rlabel metal1 s 48822 0 48858 395 4 br_0_78
rlabel metal1 s 48966 0 49002 395 4 bl_1_78
rlabel metal1 s 49038 0 49074 395 4 br_1_78
rlabel metal1 s 49806 0 49842 395 4 bl_0_79
rlabel metal1 s 49734 0 49770 395 4 br_0_79
rlabel metal1 s 49590 0 49626 395 4 bl_1_79
rlabel metal1 s 49518 0 49554 395 4 br_1_79
rlabel metal1 s 49998 0 50034 395 4 bl_0_80
rlabel metal1 s 50070 0 50106 395 4 br_0_80
rlabel metal1 s 50214 0 50250 395 4 bl_1_80
rlabel metal1 s 50286 0 50322 395 4 br_1_80
rlabel metal1 s 51054 0 51090 395 4 bl_0_81
rlabel metal1 s 50982 0 51018 395 4 br_0_81
rlabel metal1 s 50838 0 50874 395 4 bl_1_81
rlabel metal1 s 50766 0 50802 395 4 br_1_81
rlabel metal1 s 51246 0 51282 395 4 bl_0_82
rlabel metal1 s 51318 0 51354 395 4 br_0_82
rlabel metal1 s 51462 0 51498 395 4 bl_1_82
rlabel metal1 s 51534 0 51570 395 4 br_1_82
rlabel metal1 s 52302 0 52338 395 4 bl_0_83
rlabel metal1 s 52230 0 52266 395 4 br_0_83
rlabel metal1 s 52086 0 52122 395 4 bl_1_83
rlabel metal1 s 52014 0 52050 395 4 br_1_83
rlabel metal1 s 52494 0 52530 395 4 bl_0_84
rlabel metal1 s 52566 0 52602 395 4 br_0_84
rlabel metal1 s 52710 0 52746 395 4 bl_1_84
rlabel metal1 s 52782 0 52818 395 4 br_1_84
rlabel metal1 s 53550 0 53586 395 4 bl_0_85
rlabel metal1 s 53478 0 53514 395 4 br_0_85
rlabel metal1 s 53334 0 53370 395 4 bl_1_85
rlabel metal1 s 53262 0 53298 395 4 br_1_85
rlabel metal1 s 53742 0 53778 395 4 bl_0_86
rlabel metal1 s 53814 0 53850 395 4 br_0_86
rlabel metal1 s 53958 0 53994 395 4 bl_1_86
rlabel metal1 s 54030 0 54066 395 4 br_1_86
rlabel metal1 s 54798 0 54834 395 4 bl_0_87
rlabel metal1 s 54726 0 54762 395 4 br_0_87
rlabel metal1 s 54582 0 54618 395 4 bl_1_87
rlabel metal1 s 54510 0 54546 395 4 br_1_87
rlabel metal1 s 54990 0 55026 395 4 bl_0_88
rlabel metal1 s 55062 0 55098 395 4 br_0_88
rlabel metal1 s 55206 0 55242 395 4 bl_1_88
rlabel metal1 s 55278 0 55314 395 4 br_1_88
rlabel metal1 s 56046 0 56082 395 4 bl_0_89
rlabel metal1 s 55974 0 56010 395 4 br_0_89
rlabel metal1 s 55830 0 55866 395 4 bl_1_89
rlabel metal1 s 55758 0 55794 395 4 br_1_89
rlabel metal1 s 56238 0 56274 395 4 bl_0_90
rlabel metal1 s 56310 0 56346 395 4 br_0_90
rlabel metal1 s 56454 0 56490 395 4 bl_1_90
rlabel metal1 s 56526 0 56562 395 4 br_1_90
rlabel metal1 s 57294 0 57330 395 4 bl_0_91
rlabel metal1 s 57222 0 57258 395 4 br_0_91
rlabel metal1 s 57078 0 57114 395 4 bl_1_91
rlabel metal1 s 57006 0 57042 395 4 br_1_91
rlabel metal1 s 57486 0 57522 395 4 bl_0_92
rlabel metal1 s 57558 0 57594 395 4 br_0_92
rlabel metal1 s 57702 0 57738 395 4 bl_1_92
rlabel metal1 s 57774 0 57810 395 4 br_1_92
rlabel metal1 s 58542 0 58578 395 4 bl_0_93
rlabel metal1 s 58470 0 58506 395 4 br_0_93
rlabel metal1 s 58326 0 58362 395 4 bl_1_93
rlabel metal1 s 58254 0 58290 395 4 br_1_93
rlabel metal1 s 58734 0 58770 395 4 bl_0_94
rlabel metal1 s 58806 0 58842 395 4 br_0_94
rlabel metal1 s 58950 0 58986 395 4 bl_1_94
rlabel metal1 s 59022 0 59058 395 4 br_1_94
rlabel metal1 s 59790 0 59826 395 4 bl_0_95
rlabel metal1 s 59718 0 59754 395 4 br_0_95
rlabel metal1 s 59574 0 59610 395 4 bl_1_95
rlabel metal1 s 59502 0 59538 395 4 br_1_95
rlabel metal1 s 59982 0 60018 395 4 bl_0_96
rlabel metal1 s 60054 0 60090 395 4 br_0_96
rlabel metal1 s 60198 0 60234 395 4 bl_1_96
rlabel metal1 s 60270 0 60306 395 4 br_1_96
rlabel metal1 s 61038 0 61074 395 4 bl_0_97
rlabel metal1 s 60966 0 61002 395 4 br_0_97
rlabel metal1 s 60822 0 60858 395 4 bl_1_97
rlabel metal1 s 60750 0 60786 395 4 br_1_97
rlabel metal1 s 61230 0 61266 395 4 bl_0_98
rlabel metal1 s 61302 0 61338 395 4 br_0_98
rlabel metal1 s 61446 0 61482 395 4 bl_1_98
rlabel metal1 s 61518 0 61554 395 4 br_1_98
rlabel metal1 s 62286 0 62322 395 4 bl_0_99
rlabel metal1 s 62214 0 62250 395 4 br_0_99
rlabel metal1 s 62070 0 62106 395 4 bl_1_99
rlabel metal1 s 61998 0 62034 395 4 br_1_99
rlabel metal1 s 62478 0 62514 395 4 bl_0_100
rlabel metal1 s 62550 0 62586 395 4 br_0_100
rlabel metal1 s 62694 0 62730 395 4 bl_1_100
rlabel metal1 s 62766 0 62802 395 4 br_1_100
rlabel metal1 s 63534 0 63570 395 4 bl_0_101
rlabel metal1 s 63462 0 63498 395 4 br_0_101
rlabel metal1 s 63318 0 63354 395 4 bl_1_101
rlabel metal1 s 63246 0 63282 395 4 br_1_101
rlabel metal1 s 63726 0 63762 395 4 bl_0_102
rlabel metal1 s 63798 0 63834 395 4 br_0_102
rlabel metal1 s 63942 0 63978 395 4 bl_1_102
rlabel metal1 s 64014 0 64050 395 4 br_1_102
rlabel metal1 s 64782 0 64818 395 4 bl_0_103
rlabel metal1 s 64710 0 64746 395 4 br_0_103
rlabel metal1 s 64566 0 64602 395 4 bl_1_103
rlabel metal1 s 64494 0 64530 395 4 br_1_103
rlabel metal1 s 64974 0 65010 395 4 bl_0_104
rlabel metal1 s 65046 0 65082 395 4 br_0_104
rlabel metal1 s 65190 0 65226 395 4 bl_1_104
rlabel metal1 s 65262 0 65298 395 4 br_1_104
rlabel metal1 s 66030 0 66066 395 4 bl_0_105
rlabel metal1 s 65958 0 65994 395 4 br_0_105
rlabel metal1 s 65814 0 65850 395 4 bl_1_105
rlabel metal1 s 65742 0 65778 395 4 br_1_105
rlabel metal1 s 66222 0 66258 395 4 bl_0_106
rlabel metal1 s 66294 0 66330 395 4 br_0_106
rlabel metal1 s 66438 0 66474 395 4 bl_1_106
rlabel metal1 s 66510 0 66546 395 4 br_1_106
rlabel metal1 s 67278 0 67314 395 4 bl_0_107
rlabel metal1 s 67206 0 67242 395 4 br_0_107
rlabel metal1 s 67062 0 67098 395 4 bl_1_107
rlabel metal1 s 66990 0 67026 395 4 br_1_107
rlabel metal1 s 67470 0 67506 395 4 bl_0_108
rlabel metal1 s 67542 0 67578 395 4 br_0_108
rlabel metal1 s 67686 0 67722 395 4 bl_1_108
rlabel metal1 s 67758 0 67794 395 4 br_1_108
rlabel metal1 s 68526 0 68562 395 4 bl_0_109
rlabel metal1 s 68454 0 68490 395 4 br_0_109
rlabel metal1 s 68310 0 68346 395 4 bl_1_109
rlabel metal1 s 68238 0 68274 395 4 br_1_109
rlabel metal1 s 68718 0 68754 395 4 bl_0_110
rlabel metal1 s 68790 0 68826 395 4 br_0_110
rlabel metal1 s 68934 0 68970 395 4 bl_1_110
rlabel metal1 s 69006 0 69042 395 4 br_1_110
rlabel metal1 s 69774 0 69810 395 4 bl_0_111
rlabel metal1 s 69702 0 69738 395 4 br_0_111
rlabel metal1 s 69558 0 69594 395 4 bl_1_111
rlabel metal1 s 69486 0 69522 395 4 br_1_111
rlabel metal1 s 69966 0 70002 395 4 bl_0_112
rlabel metal1 s 70038 0 70074 395 4 br_0_112
rlabel metal1 s 70182 0 70218 395 4 bl_1_112
rlabel metal1 s 70254 0 70290 395 4 br_1_112
rlabel metal1 s 71022 0 71058 395 4 bl_0_113
rlabel metal1 s 70950 0 70986 395 4 br_0_113
rlabel metal1 s 70806 0 70842 395 4 bl_1_113
rlabel metal1 s 70734 0 70770 395 4 br_1_113
rlabel metal1 s 71214 0 71250 395 4 bl_0_114
rlabel metal1 s 71286 0 71322 395 4 br_0_114
rlabel metal1 s 71430 0 71466 395 4 bl_1_114
rlabel metal1 s 71502 0 71538 395 4 br_1_114
rlabel metal1 s 72270 0 72306 395 4 bl_0_115
rlabel metal1 s 72198 0 72234 395 4 br_0_115
rlabel metal1 s 72054 0 72090 395 4 bl_1_115
rlabel metal1 s 71982 0 72018 395 4 br_1_115
rlabel metal1 s 72462 0 72498 395 4 bl_0_116
rlabel metal1 s 72534 0 72570 395 4 br_0_116
rlabel metal1 s 72678 0 72714 395 4 bl_1_116
rlabel metal1 s 72750 0 72786 395 4 br_1_116
rlabel metal1 s 73518 0 73554 395 4 bl_0_117
rlabel metal1 s 73446 0 73482 395 4 br_0_117
rlabel metal1 s 73302 0 73338 395 4 bl_1_117
rlabel metal1 s 73230 0 73266 395 4 br_1_117
rlabel metal1 s 73710 0 73746 395 4 bl_0_118
rlabel metal1 s 73782 0 73818 395 4 br_0_118
rlabel metal1 s 73926 0 73962 395 4 bl_1_118
rlabel metal1 s 73998 0 74034 395 4 br_1_118
rlabel metal1 s 74766 0 74802 395 4 bl_0_119
rlabel metal1 s 74694 0 74730 395 4 br_0_119
rlabel metal1 s 74550 0 74586 395 4 bl_1_119
rlabel metal1 s 74478 0 74514 395 4 br_1_119
rlabel metal1 s 74958 0 74994 395 4 bl_0_120
rlabel metal1 s 75030 0 75066 395 4 br_0_120
rlabel metal1 s 75174 0 75210 395 4 bl_1_120
rlabel metal1 s 75246 0 75282 395 4 br_1_120
rlabel metal1 s 76014 0 76050 395 4 bl_0_121
rlabel metal1 s 75942 0 75978 395 4 br_0_121
rlabel metal1 s 75798 0 75834 395 4 bl_1_121
rlabel metal1 s 75726 0 75762 395 4 br_1_121
rlabel metal1 s 76206 0 76242 395 4 bl_0_122
rlabel metal1 s 76278 0 76314 395 4 br_0_122
rlabel metal1 s 76422 0 76458 395 4 bl_1_122
rlabel metal1 s 76494 0 76530 395 4 br_1_122
rlabel metal1 s 77262 0 77298 395 4 bl_0_123
rlabel metal1 s 77190 0 77226 395 4 br_0_123
rlabel metal1 s 77046 0 77082 395 4 bl_1_123
rlabel metal1 s 76974 0 77010 395 4 br_1_123
rlabel metal1 s 77454 0 77490 395 4 bl_0_124
rlabel metal1 s 77526 0 77562 395 4 br_0_124
rlabel metal1 s 77670 0 77706 395 4 bl_1_124
rlabel metal1 s 77742 0 77778 395 4 br_1_124
rlabel metal1 s 78510 0 78546 395 4 bl_0_125
rlabel metal1 s 78438 0 78474 395 4 br_0_125
rlabel metal1 s 78294 0 78330 395 4 bl_1_125
rlabel metal1 s 78222 0 78258 395 4 br_1_125
rlabel metal1 s 78702 0 78738 395 4 bl_0_126
rlabel metal1 s 78774 0 78810 395 4 br_0_126
rlabel metal1 s 78918 0 78954 395 4 bl_1_126
rlabel metal1 s 78990 0 79026 395 4 br_1_126
rlabel metal1 s 79758 0 79794 395 4 bl_0_127
rlabel metal1 s 79686 0 79722 395 4 br_0_127
rlabel metal1 s 79542 0 79578 395 4 bl_1_127
rlabel metal1 s 79470 0 79506 395 4 br_1_127
rlabel metal2 s 0 323 79872 371 4 wl_0_0
rlabel metal2 s 0 103 79872 151 4 wl_1_0
rlabel metal1 s 10206 79 10242 420 4 vdd
rlabel metal1 s 53406 79 53442 420 4 vdd
rlabel metal1 s 38910 79 38946 420 4 vdd
rlabel metal1 s 12222 79 12258 420 4 vdd
rlabel metal1 s 12702 79 12738 420 4 vdd
rlabel metal1 s 21438 79 21474 420 4 vdd
rlabel metal1 s 66366 79 66402 420 4 vdd
rlabel metal1 s 25950 79 25986 420 4 vdd
rlabel metal1 s 30174 79 30210 420 4 vdd
rlabel metal1 s 55134 79 55170 420 4 vdd
rlabel metal1 s 42174 79 42210 420 4 vdd
rlabel metal1 s 3966 79 4002 420 4 vdd
rlabel metal1 s 75870 79 75906 420 4 vdd
rlabel metal1 s 22686 79 22722 420 4 vdd
rlabel metal1 s 14718 79 14754 420 4 vdd
rlabel metal1 s 58878 79 58914 420 4 vdd
rlabel metal1 s 41406 79 41442 420 4 vdd
rlabel metal1 s 25182 79 25218 420 4 vdd
rlabel metal1 s 8958 79 8994 420 4 vdd
rlabel metal1 s 70878 79 70914 420 4 vdd
rlabel metal1 s 24702 79 24738 420 4 vdd
rlabel metal1 s 47166 79 47202 420 4 vdd
rlabel metal1 s 3486 79 3522 420 4 vdd
rlabel metal1 s 48894 79 48930 420 4 vdd
rlabel metal1 s 49662 79 49698 420 4 vdd
rlabel metal1 s 53886 79 53922 420 4 vdd
rlabel metal1 s 29694 79 29730 420 4 vdd
rlabel metal1 s 78846 79 78882 420 4 vdd
rlabel metal1 s 13470 79 13506 420 4 vdd
rlabel metal1 s 38430 79 38466 420 4 vdd
rlabel metal1 s 72126 79 72162 420 4 vdd
rlabel metal1 s 75102 79 75138 420 4 vdd
rlabel metal1 s 73854 79 73890 420 4 vdd
rlabel metal1 s 77118 79 77154 420 4 vdd
rlabel metal1 s 39678 79 39714 420 4 vdd
rlabel metal1 s 26430 79 26466 420 4 vdd
rlabel metal1 s 64638 79 64674 420 4 vdd
rlabel metal1 s 60126 79 60162 420 4 vdd
rlabel metal1 s 65886 79 65922 420 4 vdd
rlabel metal1 s 52638 79 52674 420 4 vdd
rlabel metal1 s 48414 79 48450 420 4 vdd
rlabel metal1 s 47646 79 47682 420 4 vdd
rlabel metal1 s 42654 79 42690 420 4 vdd
rlabel metal1 s 35934 79 35970 420 4 vdd
rlabel metal1 s 37182 79 37218 420 4 vdd
rlabel metal1 s 63390 79 63426 420 4 vdd
rlabel metal1 s 4734 79 4770 420 4 vdd
rlabel metal1 s 28446 79 28482 420 4 vdd
rlabel metal1 s 60894 79 60930 420 4 vdd
rlabel metal1 s 72606 79 72642 420 4 vdd
rlabel metal1 s 43902 79 43938 420 4 vdd
rlabel metal1 s 67614 79 67650 420 4 vdd
rlabel metal1 s 17694 79 17730 420 4 vdd
rlabel metal1 s 28926 79 28962 420 4 vdd
rlabel metal1 s 27678 79 27714 420 4 vdd
rlabel metal1 s 18462 79 18498 420 4 vdd
rlabel metal1 s 30942 79 30978 420 4 vdd
rlabel metal1 s 68862 79 68898 420 4 vdd
rlabel metal1 s 68382 79 68418 420 4 vdd
rlabel metal1 s 40926 79 40962 420 4 vdd
rlabel metal1 s 74622 79 74658 420 4 vdd
rlabel metal1 s 32670 79 32706 420 4 vdd
rlabel metal1 s 33918 79 33954 420 4 vdd
rlabel metal1 s 23934 79 23970 420 4 vdd
rlabel metal1 s 8478 79 8514 420 4 vdd
rlabel metal1 s 20190 79 20226 420 4 vdd
rlabel metal1 s 37662 79 37698 420 4 vdd
rlabel metal1 s 35166 79 35202 420 4 vdd
rlabel metal1 s 76350 79 76386 420 4 vdd
rlabel metal1 s 11454 79 11490 420 4 vdd
rlabel metal1 s 15198 79 15234 420 4 vdd
rlabel metal1 s 1470 79 1506 420 4 vdd
rlabel metal1 s 46398 79 46434 420 4 vdd
rlabel metal1 s 79614 79 79650 420 4 vdd
rlabel metal1 s 50142 79 50178 420 4 vdd
rlabel metal1 s 57630 79 57666 420 4 vdd
rlabel metal1 s 59646 79 59682 420 4 vdd
rlabel metal1 s 18942 79 18978 420 4 vdd
rlabel metal1 s 54654 79 54690 420 4 vdd
rlabel metal1 s 70110 79 70146 420 4 vdd
rlabel metal1 s 77598 79 77634 420 4 vdd
rlabel metal1 s 56382 79 56418 420 4 vdd
rlabel metal1 s 27198 79 27234 420 4 vdd
rlabel metal1 s 51390 79 51426 420 4 vdd
rlabel metal1 s 45918 79 45954 420 4 vdd
rlabel metal1 s 31422 79 31458 420 4 vdd
rlabel metal1 s 990 79 1026 420 4 vdd
rlabel metal1 s 22206 79 22242 420 4 vdd
rlabel metal1 s 67134 79 67170 420 4 vdd
rlabel metal1 s 73374 79 73410 420 4 vdd
rlabel metal1 s 7710 79 7746 420 4 vdd
rlabel metal1 s 62142 79 62178 420 4 vdd
rlabel metal1 s 78366 79 78402 420 4 vdd
rlabel metal1 s 61374 79 61410 420 4 vdd
rlabel metal1 s 9726 79 9762 420 4 vdd
rlabel metal1 s 5982 79 6018 420 4 vdd
rlabel metal1 s 33438 79 33474 420 4 vdd
rlabel metal1 s 43422 79 43458 420 4 vdd
rlabel metal1 s 55902 79 55938 420 4 vdd
rlabel metal1 s 65118 79 65154 420 4 vdd
rlabel metal1 s 19710 79 19746 420 4 vdd
rlabel metal1 s 50910 79 50946 420 4 vdd
rlabel metal1 s 23454 79 23490 420 4 vdd
rlabel metal1 s 58398 79 58434 420 4 vdd
rlabel metal1 s 36414 79 36450 420 4 vdd
rlabel metal1 s 69630 79 69666 420 4 vdd
rlabel metal1 s 2238 79 2274 420 4 vdd
rlabel metal1 s 62622 79 62658 420 4 vdd
rlabel metal1 s 10974 79 11010 420 4 vdd
rlabel metal1 s 2718 79 2754 420 4 vdd
rlabel metal1 s 57150 79 57186 420 4 vdd
rlabel metal1 s 44670 79 44706 420 4 vdd
rlabel metal1 s 52158 79 52194 420 4 vdd
rlabel metal1 s 6462 79 6498 420 4 vdd
rlabel metal1 s 32190 79 32226 420 4 vdd
rlabel metal1 s 34686 79 34722 420 4 vdd
rlabel metal1 s 17214 79 17250 420 4 vdd
rlabel metal1 s 222 79 258 420 4 vdd
rlabel metal1 s 15966 79 16002 420 4 vdd
rlabel metal1 s 20958 79 20994 420 4 vdd
rlabel metal1 s 7230 79 7266 420 4 vdd
rlabel metal1 s 40158 79 40194 420 4 vdd
rlabel metal1 s 63870 79 63906 420 4 vdd
rlabel metal1 s 5214 79 5250 420 4 vdd
rlabel metal1 s 16446 79 16482 420 4 vdd
rlabel metal1 s 13950 79 13986 420 4 vdd
rlabel metal1 s 45150 79 45186 420 4 vdd
rlabel metal1 s 71358 79 71394 420 4 vdd
rlabel metal2 s 2202 199 2310 275 4 gnd
rlabel metal2 s 35898 -55 36006 55 4 gnd
rlabel metal2 s 24666 -55 24774 55 4 gnd
rlabel metal2 s 33882 199 33990 275 4 gnd
rlabel metal2 s 70842 199 70950 275 4 gnd
rlabel metal2 s 58362 -55 58470 55 4 gnd
rlabel metal2 s 52602 199 52710 275 4 gnd
rlabel metal2 s 68826 199 68934 275 4 gnd
rlabel metal2 s 47130 199 47238 275 4 gnd
rlabel metal2 s 38394 -55 38502 55 4 gnd
rlabel metal2 s 38874 199 38982 275 4 gnd
rlabel metal2 s 43386 -55 43494 55 4 gnd
rlabel metal2 s 76314 -55 76422 55 4 gnd
rlabel metal2 s 6426 199 6534 275 4 gnd
rlabel metal2 s 37146 -55 37254 55 4 gnd
rlabel metal2 s 67578 199 67686 275 4 gnd
rlabel metal2 s 12666 199 12774 275 4 gnd
rlabel metal2 s 41370 -55 41478 55 4 gnd
rlabel metal2 s 45882 -55 45990 55 4 gnd
rlabel metal2 s 35130 -55 35238 55 4 gnd
rlabel metal2 s 36378 199 36486 275 4 gnd
rlabel metal2 s 73338 -55 73446 55 4 gnd
rlabel metal2 s 77562 -55 77670 55 4 gnd
rlabel metal2 s 1434 199 1542 275 4 gnd
rlabel metal2 s 6426 -55 6534 55 4 gnd
rlabel metal2 s 9690 -55 9798 55 4 gnd
rlabel metal2 s 18906 199 19014 275 4 gnd
rlabel metal2 s 44634 199 44742 275 4 gnd
rlabel metal2 s 49626 199 49734 275 4 gnd
rlabel metal2 s 14682 199 14790 275 4 gnd
rlabel metal2 s 58842 199 58950 275 4 gnd
rlabel metal2 s 17658 199 17766 275 4 gnd
rlabel metal2 s 25146 199 25254 275 4 gnd
rlabel metal2 s 78330 -55 78438 55 4 gnd
rlabel metal2 s 60090 -55 60198 55 4 gnd
rlabel metal2 s 65850 199 65958 275 4 gnd
rlabel metal2 s 5178 -55 5286 55 4 gnd
rlabel metal2 s 51354 199 51462 275 4 gnd
rlabel metal2 s 28410 -55 28518 55 4 gnd
rlabel metal2 s 52602 -55 52710 55 4 gnd
rlabel metal2 s 15162 -55 15270 55 4 gnd
rlabel metal2 s 7194 199 7302 275 4 gnd
rlabel metal2 s 8922 199 9030 275 4 gnd
rlabel metal2 s 17658 -55 17766 55 4 gnd
rlabel metal2 s 21402 -55 21510 55 4 gnd
rlabel metal2 s 58842 -55 58950 55 4 gnd
rlabel metal2 s 18426 199 18534 275 4 gnd
rlabel metal2 s 63834 199 63942 275 4 gnd
rlabel metal2 s 8442 199 8550 275 4 gnd
rlabel metal2 s 52122 199 52230 275 4 gnd
rlabel metal2 s 59610 -55 59718 55 4 gnd
rlabel metal2 s 2682 -55 2790 55 4 gnd
rlabel metal2 s 13434 -55 13542 55 4 gnd
rlabel metal2 s 28410 199 28518 275 4 gnd
rlabel metal2 s 48378 -55 48486 55 4 gnd
rlabel metal2 s 53370 199 53478 275 4 gnd
rlabel metal2 s 10170 -55 10278 55 4 gnd
rlabel metal2 s 14682 -55 14790 55 4 gnd
rlabel metal2 s 75066 199 75174 275 4 gnd
rlabel metal2 s 13914 199 14022 275 4 gnd
rlabel metal2 s 186 199 294 275 4 gnd
rlabel metal2 s 5946 199 6054 275 4 gnd
rlabel metal2 s 53850 199 53958 275 4 gnd
rlabel metal2 s 47130 -55 47238 55 4 gnd
rlabel metal2 s 78810 199 78918 275 4 gnd
rlabel metal2 s 186 -55 294 55 4 gnd
rlabel metal2 s 20922 -55 21030 55 4 gnd
rlabel metal2 s 8442 -55 8550 55 4 gnd
rlabel metal2 s 22170 199 22278 275 4 gnd
rlabel metal2 s 39642 199 39750 275 4 gnd
rlabel metal2 s 46362 -55 46470 55 4 gnd
rlabel metal2 s 54618 -55 54726 55 4 gnd
rlabel metal2 s 34650 199 34758 275 4 gnd
rlabel metal2 s 61338 199 61446 275 4 gnd
rlabel metal2 s 59610 199 59718 275 4 gnd
rlabel metal2 s 49626 -55 49734 55 4 gnd
rlabel metal2 s 7674 199 7782 275 4 gnd
rlabel metal2 s 65082 199 65190 275 4 gnd
rlabel metal2 s 15162 199 15270 275 4 gnd
rlabel metal2 s 40890 199 40998 275 4 gnd
rlabel metal2 s 44634 -55 44742 55 4 gnd
rlabel metal2 s 45114 -55 45222 55 4 gnd
rlabel metal2 s 68826 -55 68934 55 4 gnd
rlabel metal2 s 63354 -55 63462 55 4 gnd
rlabel metal2 s 71322 -55 71430 55 4 gnd
rlabel metal2 s 10938 -55 11046 55 4 gnd
rlabel metal2 s 56346 199 56454 275 4 gnd
rlabel metal2 s 79578 -55 79686 55 4 gnd
rlabel metal2 s 37626 199 37734 275 4 gnd
rlabel metal2 s 34650 -55 34758 55 4 gnd
rlabel metal2 s 63834 -55 63942 55 4 gnd
rlabel metal2 s 57114 199 57222 275 4 gnd
rlabel metal2 s 32154 -55 32262 55 4 gnd
rlabel metal2 s 50106 -55 50214 55 4 gnd
rlabel metal2 s 3450 -55 3558 55 4 gnd
rlabel metal2 s 61338 -55 61446 55 4 gnd
rlabel metal2 s 35130 199 35238 275 4 gnd
rlabel metal2 s 42618 199 42726 275 4 gnd
rlabel metal2 s 69594 -55 69702 55 4 gnd
rlabel metal2 s 27642 199 27750 275 4 gnd
rlabel metal2 s 15930 199 16038 275 4 gnd
rlabel metal2 s 55098 199 55206 275 4 gnd
rlabel metal2 s 56346 -55 56454 55 4 gnd
rlabel metal2 s 19674 -55 19782 55 4 gnd
rlabel metal2 s 37626 -55 37734 55 4 gnd
rlabel metal2 s 55866 199 55974 275 4 gnd
rlabel metal2 s 16410 199 16518 275 4 gnd
rlabel metal2 s 17178 199 17286 275 4 gnd
rlabel metal2 s 71322 199 71430 275 4 gnd
rlabel metal2 s 74586 -55 74694 55 4 gnd
rlabel metal2 s 30138 199 30246 275 4 gnd
rlabel metal2 s 23898 199 24006 275 4 gnd
rlabel metal2 s 20922 199 21030 275 4 gnd
rlabel metal2 s 1434 -55 1542 55 4 gnd
rlabel metal2 s 954 -55 1062 55 4 gnd
rlabel metal2 s 32634 199 32742 275 4 gnd
rlabel metal2 s 12186 199 12294 275 4 gnd
rlabel metal2 s 52122 -55 52230 55 4 gnd
rlabel metal2 s 79578 199 79686 275 4 gnd
rlabel metal2 s 13434 199 13542 275 4 gnd
rlabel metal2 s 78810 -55 78918 55 4 gnd
rlabel metal2 s 66330 -55 66438 55 4 gnd
rlabel metal2 s 57594 -55 57702 55 4 gnd
rlabel metal2 s 51354 -55 51462 55 4 gnd
rlabel metal2 s 3930 199 4038 275 4 gnd
rlabel metal2 s 30906 -55 31014 55 4 gnd
rlabel metal2 s 50874 199 50982 275 4 gnd
rlabel metal2 s 77562 199 77670 275 4 gnd
rlabel metal2 s 48858 199 48966 275 4 gnd
rlabel metal2 s 37146 199 37254 275 4 gnd
rlabel metal2 s 57114 -55 57222 55 4 gnd
rlabel metal2 s 66330 199 66438 275 4 gnd
rlabel metal2 s 8922 -55 9030 55 4 gnd
rlabel metal2 s 12666 -55 12774 55 4 gnd
rlabel metal2 s 13914 -55 14022 55 4 gnd
rlabel metal2 s 23418 -55 23526 55 4 gnd
rlabel metal2 s 45114 199 45222 275 4 gnd
rlabel metal2 s 3930 -55 4038 55 4 gnd
rlabel metal2 s 11418 199 11526 275 4 gnd
rlabel metal2 s 7194 -55 7302 55 4 gnd
rlabel metal2 s 31386 199 31494 275 4 gnd
rlabel metal2 s 42618 -55 42726 55 4 gnd
rlabel metal2 s 65850 -55 65958 55 4 gnd
rlabel metal2 s 39642 -55 39750 55 4 gnd
rlabel metal2 s 18906 -55 19014 55 4 gnd
rlabel metal2 s 27162 -55 27270 55 4 gnd
rlabel metal2 s 67098 -55 67206 55 4 gnd
rlabel metal2 s 63354 199 63462 275 4 gnd
rlabel metal2 s 33402 -55 33510 55 4 gnd
rlabel metal2 s 70074 199 70182 275 4 gnd
rlabel metal2 s 68346 -55 68454 55 4 gnd
rlabel metal2 s 31386 -55 31494 55 4 gnd
rlabel metal2 s 30138 -55 30246 55 4 gnd
rlabel metal2 s 21402 199 21510 275 4 gnd
rlabel metal2 s 25914 199 26022 275 4 gnd
rlabel metal2 s 75066 -55 75174 55 4 gnd
rlabel metal2 s 15930 -55 16038 55 4 gnd
rlabel metal2 s 43386 199 43494 275 4 gnd
rlabel metal2 s 33882 -55 33990 55 4 gnd
rlabel metal2 s 42138 199 42246 275 4 gnd
rlabel metal2 s 10938 199 11046 275 4 gnd
rlabel metal2 s 40122 -55 40230 55 4 gnd
rlabel metal2 s 29658 199 29766 275 4 gnd
rlabel metal2 s 10170 199 10278 275 4 gnd
rlabel metal2 s 69594 199 69702 275 4 gnd
rlabel metal2 s 27642 -55 27750 55 4 gnd
rlabel metal2 s 2682 199 2790 275 4 gnd
rlabel metal2 s 41370 199 41478 275 4 gnd
rlabel metal2 s 40890 -55 40998 55 4 gnd
rlabel metal2 s 43866 199 43974 275 4 gnd
rlabel metal2 s 46362 199 46470 275 4 gnd
rlabel metal2 s 55866 -55 55974 55 4 gnd
rlabel metal2 s 60858 199 60966 275 4 gnd
rlabel metal2 s 4698 -55 4806 55 4 gnd
rlabel metal2 s 25914 -55 26022 55 4 gnd
rlabel metal2 s 48378 199 48486 275 4 gnd
rlabel metal2 s 53370 -55 53478 55 4 gnd
rlabel metal2 s 22170 -55 22278 55 4 gnd
rlabel metal2 s 32634 -55 32742 55 4 gnd
rlabel metal2 s 40122 199 40230 275 4 gnd
rlabel metal2 s 62586 -55 62694 55 4 gnd
rlabel metal2 s 64602 -55 64710 55 4 gnd
rlabel metal2 s 76314 199 76422 275 4 gnd
rlabel metal2 s 19674 199 19782 275 4 gnd
rlabel metal2 s 18426 -55 18534 55 4 gnd
rlabel metal2 s 20154 -55 20262 55 4 gnd
rlabel metal2 s 68346 199 68454 275 4 gnd
rlabel metal2 s 72570 -55 72678 55 4 gnd
rlabel metal2 s 57594 199 57702 275 4 gnd
rlabel metal2 s 5946 -55 6054 55 4 gnd
rlabel metal2 s 25146 -55 25254 55 4 gnd
rlabel metal2 s 73818 -55 73926 55 4 gnd
rlabel metal2 s 62106 -55 62214 55 4 gnd
rlabel metal2 s 54618 199 54726 275 4 gnd
rlabel metal2 s 38394 199 38502 275 4 gnd
rlabel metal2 s 7674 -55 7782 55 4 gnd
rlabel metal2 s 20154 199 20262 275 4 gnd
rlabel metal2 s 70842 -55 70950 55 4 gnd
rlabel metal2 s 47610 -55 47718 55 4 gnd
rlabel metal2 s 72090 -55 72198 55 4 gnd
rlabel metal2 s 78330 199 78438 275 4 gnd
rlabel metal2 s 33402 199 33510 275 4 gnd
rlabel metal2 s 77082 -55 77190 55 4 gnd
rlabel metal2 s 62106 199 62214 275 4 gnd
rlabel metal2 s 9690 199 9798 275 4 gnd
rlabel metal2 s 62586 199 62694 275 4 gnd
rlabel metal2 s 954 199 1062 275 4 gnd
rlabel metal2 s 3450 199 3558 275 4 gnd
rlabel metal2 s 2202 -55 2310 55 4 gnd
rlabel metal2 s 12186 -55 12294 55 4 gnd
rlabel metal2 s 70074 -55 70182 55 4 gnd
rlabel metal2 s 77082 199 77190 275 4 gnd
rlabel metal2 s 22650 199 22758 275 4 gnd
rlabel metal2 s 73338 199 73446 275 4 gnd
rlabel metal2 s 72090 199 72198 275 4 gnd
rlabel metal2 s 5178 199 5286 275 4 gnd
rlabel metal2 s 16410 -55 16518 55 4 gnd
rlabel metal2 s 50106 199 50214 275 4 gnd
rlabel metal2 s 53850 -55 53958 55 4 gnd
rlabel metal2 s 75834 -55 75942 55 4 gnd
rlabel metal2 s 32154 199 32262 275 4 gnd
rlabel metal2 s 55098 -55 55206 55 4 gnd
rlabel metal2 s 47610 199 47718 275 4 gnd
rlabel metal2 s 23898 -55 24006 55 4 gnd
rlabel metal2 s 28890 199 28998 275 4 gnd
rlabel metal2 s 11418 -55 11526 55 4 gnd
rlabel metal2 s 28890 -55 28998 55 4 gnd
rlabel metal2 s 27162 199 27270 275 4 gnd
rlabel metal2 s 42138 -55 42246 55 4 gnd
rlabel metal2 s 17178 -55 17286 55 4 gnd
rlabel metal2 s 74586 199 74694 275 4 gnd
rlabel metal2 s 43866 -55 43974 55 4 gnd
rlabel metal2 s 30906 199 31014 275 4 gnd
rlabel metal2 s 72570 199 72678 275 4 gnd
rlabel metal2 s 67098 199 67206 275 4 gnd
rlabel metal2 s 4698 199 4806 275 4 gnd
rlabel metal2 s 36378 -55 36486 55 4 gnd
rlabel metal2 s 24666 199 24774 275 4 gnd
rlabel metal2 s 65082 -55 65190 55 4 gnd
rlabel metal2 s 60090 199 60198 275 4 gnd
rlabel metal2 s 67578 -55 67686 55 4 gnd
rlabel metal2 s 35898 199 36006 275 4 gnd
rlabel metal2 s 50874 -55 50982 55 4 gnd
rlabel metal2 s 64602 199 64710 275 4 gnd
rlabel metal2 s 22650 -55 22758 55 4 gnd
rlabel metal2 s 29658 -55 29766 55 4 gnd
rlabel metal2 s 60858 -55 60966 55 4 gnd
rlabel metal2 s 73818 199 73926 275 4 gnd
rlabel metal2 s 26394 -55 26502 55 4 gnd
rlabel metal2 s 58362 199 58470 275 4 gnd
rlabel metal2 s 75834 199 75942 275 4 gnd
rlabel metal2 s 38874 -55 38982 55 4 gnd
rlabel metal2 s 45882 199 45990 275 4 gnd
rlabel metal2 s 48858 -55 48966 55 4 gnd
rlabel metal2 s 23418 199 23526 275 4 gnd
rlabel metal2 s 26394 199 26502 275 4 gnd
<< properties >>
string FIXED_BBOX 0 0 79872 395
<< end >>
