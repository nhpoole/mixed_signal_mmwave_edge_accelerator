magic
tech sky130A
magscale 1 2
timestamp 1621486730
<< pwell >>
rect -2741 -310 2741 310
<< nmos >>
rect -2545 -100 -1745 100
rect -1687 -100 -887 100
rect -829 -100 -29 100
rect 29 -100 829 100
rect 887 -100 1687 100
rect 1745 -100 2545 100
<< ndiff >>
rect -2603 88 -2545 100
rect -2603 -88 -2591 88
rect -2557 -88 -2545 88
rect -2603 -100 -2545 -88
rect -1745 88 -1687 100
rect -1745 -88 -1733 88
rect -1699 -88 -1687 88
rect -1745 -100 -1687 -88
rect -887 88 -829 100
rect -887 -88 -875 88
rect -841 -88 -829 88
rect -887 -100 -829 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 829 88 887 100
rect 829 -88 841 88
rect 875 -88 887 88
rect 829 -100 887 -88
rect 1687 88 1745 100
rect 1687 -88 1699 88
rect 1733 -88 1745 88
rect 1687 -100 1745 -88
rect 2545 88 2603 100
rect 2545 -88 2557 88
rect 2591 -88 2603 88
rect 2545 -100 2603 -88
<< ndiffc >>
rect -2591 -88 -2557 88
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect 2557 -88 2591 88
<< psubdiff >>
rect -2705 240 -2609 274
rect 2609 240 2705 274
rect -2705 178 -2671 240
rect 2671 178 2705 240
rect -2705 -240 -2671 -178
rect 2671 -240 2705 -178
rect -2705 -274 -2609 -240
rect 2609 -274 2705 -240
<< psubdiffcont >>
rect -2609 240 2609 274
rect -2705 -178 -2671 178
rect 2671 -178 2705 178
rect -2609 -274 2609 -240
<< poly >>
rect -2391 172 -1899 188
rect -2391 155 -2375 172
rect -2545 138 -2375 155
rect -1915 155 -1899 172
rect -1533 172 -1041 188
rect -1533 155 -1517 172
rect -1915 138 -1745 155
rect -2545 100 -1745 138
rect -1687 138 -1517 155
rect -1057 155 -1041 172
rect -675 172 -183 188
rect -675 155 -659 172
rect -1057 138 -887 155
rect -1687 100 -887 138
rect -829 138 -659 155
rect -199 155 -183 172
rect 183 172 675 188
rect 183 155 199 172
rect -199 138 -29 155
rect -829 100 -29 138
rect 29 138 199 155
rect 659 155 675 172
rect 1041 172 1533 188
rect 1041 155 1057 172
rect 659 138 829 155
rect 29 100 829 138
rect 887 138 1057 155
rect 1517 155 1533 172
rect 1899 172 2391 188
rect 1899 155 1915 172
rect 1517 138 1687 155
rect 887 100 1687 138
rect 1745 138 1915 155
rect 2375 155 2391 172
rect 2375 138 2545 155
rect 1745 100 2545 138
rect -2545 -138 -1745 -100
rect -2545 -155 -2375 -138
rect -2391 -172 -2375 -155
rect -1915 -155 -1745 -138
rect -1687 -138 -887 -100
rect -1687 -155 -1517 -138
rect -1915 -172 -1899 -155
rect -2391 -188 -1899 -172
rect -1533 -172 -1517 -155
rect -1057 -155 -887 -138
rect -829 -138 -29 -100
rect -829 -155 -659 -138
rect -1057 -172 -1041 -155
rect -1533 -188 -1041 -172
rect -675 -172 -659 -155
rect -199 -155 -29 -138
rect 29 -138 829 -100
rect 29 -155 199 -138
rect -199 -172 -183 -155
rect -675 -188 -183 -172
rect 183 -172 199 -155
rect 659 -155 829 -138
rect 887 -138 1687 -100
rect 887 -155 1057 -138
rect 659 -172 675 -155
rect 183 -188 675 -172
rect 1041 -172 1057 -155
rect 1517 -155 1687 -138
rect 1745 -138 2545 -100
rect 1745 -155 1915 -138
rect 1517 -172 1533 -155
rect 1041 -188 1533 -172
rect 1899 -172 1915 -155
rect 2375 -155 2545 -138
rect 2375 -172 2391 -155
rect 1899 -188 2391 -172
<< polycont >>
rect -2375 138 -1915 172
rect -1517 138 -1057 172
rect -659 138 -199 172
rect 199 138 659 172
rect 1057 138 1517 172
rect 1915 138 2375 172
rect -2375 -172 -1915 -138
rect -1517 -172 -1057 -138
rect -659 -172 -199 -138
rect 199 -172 659 -138
rect 1057 -172 1517 -138
rect 1915 -172 2375 -138
<< locali >>
rect -2705 240 -2609 274
rect 2609 240 2705 274
rect -2705 178 -2671 240
rect 2671 178 2705 240
rect -2391 138 -2375 172
rect -1915 138 -1899 172
rect -1533 138 -1517 172
rect -1057 138 -1041 172
rect -675 138 -659 172
rect -199 138 -183 172
rect 183 138 199 172
rect 659 138 675 172
rect 1041 138 1057 172
rect 1517 138 1533 172
rect 1899 138 1915 172
rect 2375 138 2391 172
rect -2591 88 -2557 104
rect -2591 -104 -2557 -88
rect -1733 88 -1699 104
rect -1733 -104 -1699 -88
rect -875 88 -841 104
rect -875 -104 -841 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 841 88 875 104
rect 841 -104 875 -88
rect 1699 88 1733 104
rect 1699 -104 1733 -88
rect 2557 88 2591 104
rect 2557 -104 2591 -88
rect -2391 -172 -2375 -138
rect -1915 -172 -1899 -138
rect -1533 -172 -1517 -138
rect -1057 -172 -1041 -138
rect -675 -172 -659 -138
rect -199 -172 -183 -138
rect 183 -172 199 -138
rect 659 -172 675 -138
rect 1041 -172 1057 -138
rect 1517 -172 1533 -138
rect 1899 -172 1915 -138
rect 2375 -172 2391 -138
rect -2705 -240 -2671 -178
rect 2671 -240 2705 -178
rect -2705 -274 -2609 -240
rect 2609 -274 2705 -240
<< viali >>
rect -2337 138 -1953 172
rect -1479 138 -1095 172
rect -621 138 -237 172
rect 237 138 621 172
rect 1095 138 1479 172
rect 1953 138 2337 172
rect -2591 -88 -2557 88
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect 2557 -88 2591 88
rect -2337 -172 -1953 -138
rect -1479 -172 -1095 -138
rect -621 -172 -237 -138
rect 237 -172 621 -138
rect 1095 -172 1479 -138
rect 1953 -172 2337 -138
<< metal1 >>
rect -2349 172 -1941 178
rect -2349 138 -2337 172
rect -1953 138 -1941 172
rect -2349 132 -1941 138
rect -1491 172 -1083 178
rect -1491 138 -1479 172
rect -1095 138 -1083 172
rect -1491 132 -1083 138
rect -633 172 -225 178
rect -633 138 -621 172
rect -237 138 -225 172
rect -633 132 -225 138
rect 225 172 633 178
rect 225 138 237 172
rect 621 138 633 172
rect 225 132 633 138
rect 1083 172 1491 178
rect 1083 138 1095 172
rect 1479 138 1491 172
rect 1083 132 1491 138
rect 1941 172 2349 178
rect 1941 138 1953 172
rect 2337 138 2349 172
rect 1941 132 2349 138
rect -2597 88 -2551 100
rect -2597 -88 -2591 88
rect -2557 -88 -2551 88
rect -2597 -100 -2551 -88
rect -1739 88 -1693 100
rect -1739 -88 -1733 88
rect -1699 -88 -1693 88
rect -1739 -100 -1693 -88
rect -881 88 -835 100
rect -881 -88 -875 88
rect -841 -88 -835 88
rect -881 -100 -835 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 835 88 881 100
rect 835 -88 841 88
rect 875 -88 881 88
rect 835 -100 881 -88
rect 1693 88 1739 100
rect 1693 -88 1699 88
rect 1733 -88 1739 88
rect 1693 -100 1739 -88
rect 2551 88 2597 100
rect 2551 -88 2557 88
rect 2591 -88 2597 88
rect 2551 -100 2597 -88
rect -2349 -138 -1941 -132
rect -2349 -172 -2337 -138
rect -1953 -172 -1941 -138
rect -2349 -178 -1941 -172
rect -1491 -138 -1083 -132
rect -1491 -172 -1479 -138
rect -1095 -172 -1083 -138
rect -1491 -178 -1083 -172
rect -633 -138 -225 -132
rect -633 -172 -621 -138
rect -237 -172 -225 -138
rect -633 -178 -225 -172
rect 225 -138 633 -132
rect 225 -172 237 -138
rect 621 -172 633 -138
rect 225 -178 633 -172
rect 1083 -138 1491 -132
rect 1083 -172 1095 -138
rect 1479 -172 1491 -138
rect 1083 -178 1491 -172
rect 1941 -138 2349 -132
rect 1941 -172 1953 -138
rect 2337 -172 2349 -138
rect 1941 -178 2349 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2688 -257 2688 257
string parameters w 1 l 4 m 1 nf 6 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
