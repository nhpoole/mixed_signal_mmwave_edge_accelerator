magic
tech sky130A
magscale 1 2
timestamp 1621819980
<< metal3 >>
rect -350 972 349 1000
rect -350 428 265 972
rect 329 428 349 972
rect -350 400 349 428
rect -350 272 349 300
rect -350 -272 265 272
rect 329 -272 349 272
rect -350 -300 349 -272
rect -350 -428 349 -400
rect -350 -972 265 -428
rect 329 -972 349 -428
rect -350 -1000 349 -972
<< via3 >>
rect 265 428 329 972
rect 265 -272 329 272
rect 265 -972 329 -428
<< mimcap >>
rect -250 860 150 900
rect -250 540 -210 860
rect 110 540 150 860
rect -250 500 150 540
rect -250 160 150 200
rect -250 -160 -210 160
rect 110 -160 150 160
rect -250 -200 150 -160
rect -250 -540 150 -500
rect -250 -860 -210 -540
rect 110 -860 150 -540
rect -250 -900 150 -860
<< mimcapcontact >>
rect -210 540 110 860
rect -210 -160 110 160
rect -210 -860 110 -540
<< metal4 >>
rect -102 861 2 1050
rect 218 988 322 1050
rect 218 972 345 988
rect -211 860 111 861
rect -211 540 -210 860
rect 110 540 111 860
rect -211 539 111 540
rect -102 161 2 539
rect 218 428 265 972
rect 329 428 345 972
rect 218 412 345 428
rect 218 288 322 412
rect 218 272 345 288
rect -211 160 111 161
rect -211 -160 -210 160
rect 110 -160 111 160
rect -211 -161 111 -160
rect -102 -539 2 -161
rect 218 -272 265 272
rect 329 -272 345 272
rect 218 -288 345 -272
rect 218 -412 322 -288
rect 218 -428 345 -412
rect -211 -540 111 -539
rect -211 -860 -210 -540
rect 110 -860 111 -540
rect -211 -861 111 -860
rect -102 -1050 2 -861
rect 218 -972 265 -428
rect 329 -972 345 -428
rect 218 -988 345 -972
rect 218 -1050 322 -988
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -350 400 250 1000
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
