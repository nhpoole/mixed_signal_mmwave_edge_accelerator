magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -732 -654 732 654
<< metal3 >>
rect -102 16 102 24
rect -102 -16 -96 16
rect -64 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 64 16
rect 96 -16 102 16
rect -102 -24 102 -16
<< via3 >>
rect -96 -16 -64 16
rect -56 -16 -24 16
rect -16 -16 16 16
rect 24 -16 56 16
rect 64 -16 96 16
<< metal4 >>
rect -102 16 102 24
rect -102 -16 -96 16
rect -64 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 64 16
rect 96 -16 102 16
rect -102 -24 102 -16
<< end >>
