magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -798 -654 798 654
<< metal3 >>
rect -168 16 168 24
rect -168 -16 -156 16
rect -124 -16 -116 16
rect -84 -16 -76 16
rect -44 -16 -36 16
rect -4 -16 4 16
rect 36 -16 44 16
rect 76 -16 84 16
rect 116 -16 124 16
rect 156 -16 168 16
rect -168 -24 168 -16
<< via3 >>
rect -156 -16 -124 16
rect -116 -16 -84 16
rect -76 -16 -44 16
rect -36 -16 -4 16
rect 4 -16 36 16
rect 44 -16 76 16
rect 84 -16 116 16
rect 124 -16 156 16
<< metal4 >>
rect -168 16 168 24
rect -168 -16 -156 16
rect -124 -16 -116 16
rect -84 -16 -76 16
rect -44 -16 -36 16
rect -4 -16 4 16
rect 36 -16 44 16
rect 76 -16 84 16
rect 116 -16 124 16
rect 156 -16 168 16
rect -168 -24 168 -16
<< end >>
