magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 28 -17 62 17
<< locali >>
rect 17 211 111 323
rect 488 299 540 493
rect 506 165 540 299
rect 482 51 540 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 401 76 493
rect 110 435 153 527
rect 187 435 264 493
rect 17 357 179 401
rect 145 265 179 357
rect 145 199 196 265
rect 230 255 264 435
rect 303 349 348 486
rect 382 383 454 527
rect 303 315 448 349
rect 414 265 448 315
rect 230 215 380 255
rect 145 177 179 199
rect 19 143 179 177
rect 19 51 76 143
rect 230 109 264 215
rect 414 199 472 265
rect 414 181 448 199
rect 110 17 153 109
rect 187 51 264 109
rect 303 147 448 181
rect 303 51 348 147
rect 382 17 448 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 17 211 111 323 6 A
port 1 nsew signal input
rlabel locali s 506 165 540 299 6 X
port 2 nsew signal output
rlabel locali s 488 299 540 493 6 X
port 2 nsew signal output
rlabel locali s 482 51 540 165 6 X
port 2 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 28 -17 62 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
