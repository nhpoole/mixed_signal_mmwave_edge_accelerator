magic
tech sky130A
magscale 1 2
timestamp 1622534145
<< error_p >>
rect -35 20161084 35 20161228
rect -35 20080116 35 20080260
rect -35 19999148 35 19999292
rect -35 19918180 35 19918324
rect -35 19837212 35 19837356
rect -35 19756244 35 19756388
rect -35 19675276 35 19675420
rect -35 19594308 35 19594452
rect -35 19513340 35 19513484
rect -35 19432372 35 19432516
rect -35 19351404 35 19351548
rect -35 19270436 35 19270580
rect -35 19189468 35 19189612
rect -35 19108500 35 19108644
rect -35 19027532 35 19027676
rect -35 18946564 35 18946708
rect -35 18865596 35 18865740
rect -35 18784628 35 18784772
rect -35 18703660 35 18703804
rect -35 18622692 35 18622836
rect -35 18541724 35 18541868
rect -35 18460756 35 18460900
rect -35 18379788 35 18379932
rect -35 18298820 35 18298964
rect -35 18217852 35 18217996
rect -35 18136884 35 18137028
rect -35 18055916 35 18056060
rect -35 17974948 35 17975092
rect -35 17893980 35 17894124
rect -35 17813012 35 17813156
rect -35 17732044 35 17732188
rect -35 17651076 35 17651220
rect -35 17570108 35 17570252
rect -35 17489140 35 17489284
rect -35 17408172 35 17408316
rect -35 17327204 35 17327348
rect -35 17246236 35 17246380
rect -35 17165268 35 17165412
rect -35 17084300 35 17084444
rect -35 17003332 35 17003476
rect -35 16922364 35 16922508
rect -35 16841396 35 16841540
rect -35 16760428 35 16760572
rect -35 16679460 35 16679604
rect -35 16598492 35 16598636
rect -35 16517524 35 16517668
rect -35 16436556 35 16436700
rect -35 16355588 35 16355732
rect -35 16274620 35 16274764
rect -35 16193652 35 16193796
rect -35 16112684 35 16112828
rect -35 16031716 35 16031860
rect -35 15950748 35 15950892
rect -35 15869780 35 15869924
rect -35 15788812 35 15788956
rect -35 15707844 35 15707988
rect -35 15626876 35 15627020
rect -35 15545908 35 15546052
rect -35 15464940 35 15465084
rect -35 15383972 35 15384116
rect -35 15303004 35 15303148
rect -35 15222036 35 15222180
rect -35 15141068 35 15141212
rect -35 15060100 35 15060244
rect -35 14979132 35 14979276
rect -35 14898164 35 14898308
rect -35 14817196 35 14817340
rect -35 14736228 35 14736372
rect -35 14655260 35 14655404
rect -35 14574292 35 14574436
rect -35 14493324 35 14493468
rect -35 14412356 35 14412500
rect -35 14331388 35 14331532
rect -35 14250420 35 14250564
rect -35 14169452 35 14169596
rect -35 14088484 35 14088628
rect -35 14007516 35 14007660
rect -35 13926548 35 13926692
rect -35 13845580 35 13845724
rect -35 13764612 35 13764756
rect -35 13683644 35 13683788
rect -35 13602676 35 13602820
rect -35 13521708 35 13521852
rect -35 13440740 35 13440884
rect -35 13359772 35 13359916
rect -35 13278804 35 13278948
rect -35 13197836 35 13197980
rect -35 13116868 35 13117012
rect -35 13035900 35 13036044
rect -35 12954932 35 12955076
rect -35 12873964 35 12874108
rect -35 12792996 35 12793140
rect -35 12712028 35 12712172
rect -35 12631060 35 12631204
rect -35 12550092 35 12550236
rect -35 12469124 35 12469268
rect -35 12388156 35 12388300
rect -35 12307188 35 12307332
rect -35 12226220 35 12226364
rect -35 12145252 35 12145396
rect -35 12064284 35 12064428
rect -35 11983316 35 11983460
rect -35 11902348 35 11902492
rect -35 11821380 35 11821524
rect -35 11740412 35 11740556
rect -35 11659444 35 11659588
rect -35 11578476 35 11578620
rect -35 11497508 35 11497652
rect -35 11416540 35 11416684
rect -35 11335572 35 11335716
rect -35 11254604 35 11254748
rect -35 11173636 35 11173780
rect -35 11092668 35 11092812
rect -35 11011700 35 11011844
rect -35 10930732 35 10930876
rect -35 10849764 35 10849908
rect -35 10768796 35 10768940
rect -35 10687828 35 10687972
rect -35 10606860 35 10607004
rect -35 10525892 35 10526036
rect -35 10444924 35 10445068
rect -35 10363956 35 10364100
rect -35 10282988 35 10283132
rect -35 10202020 35 10202164
rect -35 10121052 35 10121196
rect -35 10040084 35 10040228
rect -35 9959116 35 9959260
rect -35 9878148 35 9878292
rect -35 9797180 35 9797324
rect -35 9716212 35 9716356
rect -35 9635244 35 9635388
rect -35 9554276 35 9554420
rect -35 9473308 35 9473452
rect -35 9392340 35 9392484
rect -35 9311372 35 9311516
rect -35 9230404 35 9230548
rect -35 9149436 35 9149580
rect -35 9068468 35 9068612
rect -35 8987500 35 8987644
rect -35 8906532 35 8906676
rect -35 8825564 35 8825708
rect -35 8744596 35 8744740
rect -35 8663628 35 8663772
rect -35 8582660 35 8582804
rect -35 8501692 35 8501836
rect -35 8420724 35 8420868
rect -35 8339756 35 8339900
rect -35 8258788 35 8258932
rect -35 8177820 35 8177964
rect -35 8096852 35 8096996
rect -35 8015884 35 8016028
rect -35 7934916 35 7935060
rect -35 7853948 35 7854092
rect -35 7772980 35 7773124
rect -35 7692012 35 7692156
rect -35 7611044 35 7611188
rect -35 7530076 35 7530220
rect -35 7449108 35 7449252
rect -35 7368140 35 7368284
rect -35 7287172 35 7287316
rect -35 7206204 35 7206348
rect -35 7125236 35 7125380
rect -35 7044268 35 7044412
rect -35 6963300 35 6963444
rect -35 6882332 35 6882476
rect -35 6801364 35 6801508
rect -35 6720396 35 6720540
rect -35 6639428 35 6639572
rect -35 6558460 35 6558604
rect -35 6477492 35 6477636
rect -35 6396524 35 6396668
rect -35 6315556 35 6315700
rect -35 6234588 35 6234732
rect -35 6153620 35 6153764
rect -35 6072652 35 6072796
rect -35 5991684 35 5991828
rect -35 5910716 35 5910860
rect -35 5829748 35 5829892
rect -35 5748780 35 5748924
rect -35 5667812 35 5667956
rect -35 5586844 35 5586988
rect -35 5505876 35 5506020
rect -35 5424908 35 5425052
rect -35 5343940 35 5344084
rect -35 5262972 35 5263116
rect -35 5182004 35 5182148
rect -35 5101036 35 5101180
rect -35 5020068 35 5020212
rect -35 4939100 35 4939244
rect -35 4858132 35 4858276
rect -35 4777164 35 4777308
rect -35 4696196 35 4696340
rect -35 4615228 35 4615372
rect -35 4534260 35 4534404
rect -35 4453292 35 4453436
rect -35 4372324 35 4372468
rect -35 4291356 35 4291500
rect -35 4210388 35 4210532
rect -35 4129420 35 4129564
rect -35 4048452 35 4048596
rect -35 3967484 35 3967628
rect -35 3886516 35 3886660
rect -35 3805548 35 3805692
rect -35 3724580 35 3724724
rect -35 3643612 35 3643756
rect -35 3562644 35 3562788
rect -35 3481676 35 3481820
rect -35 3400708 35 3400852
rect -35 3319740 35 3319884
rect -35 3238772 35 3238916
rect -35 3157804 35 3157948
rect -35 3076836 35 3076980
rect -35 2995868 35 2996012
rect -35 2914900 35 2915044
rect -35 2833932 35 2834076
rect -35 2752964 35 2753108
rect -35 2671996 35 2672140
rect -35 2591028 35 2591172
rect -35 2510060 35 2510204
rect -35 2429092 35 2429236
rect -35 2348124 35 2348268
rect -35 2267156 35 2267300
rect -35 2186188 35 2186332
rect -35 2105220 35 2105364
rect -35 2024252 35 2024396
rect -35 1943284 35 1943428
rect -35 1862316 35 1862460
rect -35 1781348 35 1781492
rect -35 1700380 35 1700524
rect -35 1619412 35 1619556
rect -35 1538444 35 1538588
rect -35 1457476 35 1457620
rect -35 1376508 35 1376652
rect -35 1295540 35 1295684
rect -35 1214572 35 1214716
rect -35 1133604 35 1133748
rect -35 1052636 35 1052780
rect -35 971668 35 971812
rect -35 890700 35 890844
rect -35 809732 35 809876
rect -35 728764 35 728908
rect -35 647796 35 647940
rect -35 566828 35 566972
rect -35 485860 35 486004
rect -35 404892 35 405036
rect -35 323924 35 324068
rect -35 242956 35 243100
rect -35 161988 35 162132
rect -35 81020 35 81164
rect -35 52 35 196
rect -35 -80916 35 -80772
rect -35 -161884 35 -161740
rect -35 -242852 35 -242708
rect -35 -323820 35 -323676
rect -35 -404788 35 -404644
rect -35 -485756 35 -485612
rect -35 -566724 35 -566580
rect -35 -647692 35 -647548
rect -35 -728660 35 -728516
rect -35 -809628 35 -809484
rect -35 -890596 35 -890452
rect -35 -971564 35 -971420
rect -35 -1052532 35 -1052388
rect -35 -1133500 35 -1133356
rect -35 -1214468 35 -1214324
rect -35 -1295436 35 -1295292
rect -35 -1376404 35 -1376260
rect -35 -1457372 35 -1457228
rect -35 -1538340 35 -1538196
rect -35 -1619308 35 -1619164
rect -35 -1700276 35 -1700132
rect -35 -1781244 35 -1781100
rect -35 -1862212 35 -1862068
rect -35 -1943180 35 -1943036
rect -35 -2024148 35 -2024004
rect -35 -2105116 35 -2104972
rect -35 -2186084 35 -2185940
rect -35 -2267052 35 -2266908
rect -35 -2348020 35 -2347876
rect -35 -2428988 35 -2428844
rect -35 -2509956 35 -2509812
rect -35 -2590924 35 -2590780
rect -35 -2671892 35 -2671748
rect -35 -2752860 35 -2752716
rect -35 -2833828 35 -2833684
rect -35 -2914796 35 -2914652
rect -35 -2995764 35 -2995620
rect -35 -3076732 35 -3076588
rect -35 -3157700 35 -3157556
rect -35 -3238668 35 -3238524
rect -35 -3319636 35 -3319492
rect -35 -3400604 35 -3400460
rect -35 -3481572 35 -3481428
rect -35 -3562540 35 -3562396
rect -35 -3643508 35 -3643364
rect -35 -3724476 35 -3724332
rect -35 -3805444 35 -3805300
rect -35 -3886412 35 -3886268
rect -35 -3967380 35 -3967236
rect -35 -4048348 35 -4048204
rect -35 -4129316 35 -4129172
rect -35 -4210284 35 -4210140
rect -35 -4291252 35 -4291108
rect -35 -4372220 35 -4372076
rect -35 -4453188 35 -4453044
rect -35 -4534156 35 -4534012
rect -35 -4615124 35 -4614980
rect -35 -4696092 35 -4695948
rect -35 -4777060 35 -4776916
rect -35 -4858028 35 -4857884
rect -35 -4938996 35 -4938852
rect -35 -5019964 35 -5019820
rect -35 -5100932 35 -5100788
rect -35 -5181900 35 -5181756
rect -35 -5262868 35 -5262724
rect -35 -5343836 35 -5343692
rect -35 -5424804 35 -5424660
rect -35 -5505772 35 -5505628
rect -35 -5586740 35 -5586596
rect -35 -5667708 35 -5667564
rect -35 -5748676 35 -5748532
rect -35 -5829644 35 -5829500
rect -35 -5910612 35 -5910468
rect -35 -5991580 35 -5991436
rect -35 -6072548 35 -6072404
rect -35 -6153516 35 -6153372
rect -35 -6234484 35 -6234340
rect -35 -6315452 35 -6315308
rect -35 -6396420 35 -6396276
rect -35 -6477388 35 -6477244
rect -35 -6558356 35 -6558212
rect -35 -6639324 35 -6639180
rect -35 -6720292 35 -6720148
rect -35 -6801260 35 -6801116
rect -35 -6882228 35 -6882084
rect -35 -6963196 35 -6963052
rect -35 -7044164 35 -7044020
rect -35 -7125132 35 -7124988
rect -35 -7206100 35 -7205956
rect -35 -7287068 35 -7286924
rect -35 -7368036 35 -7367892
rect -35 -7449004 35 -7448860
rect -35 -7529972 35 -7529828
rect -35 -7610940 35 -7610796
rect -35 -7691908 35 -7691764
rect -35 -7772876 35 -7772732
rect -35 -7853844 35 -7853700
rect -35 -7934812 35 -7934668
rect -35 -8015780 35 -8015636
rect -35 -8096748 35 -8096604
rect -35 -8177716 35 -8177572
rect -35 -8258684 35 -8258540
rect -35 -8339652 35 -8339508
rect -35 -8420620 35 -8420476
rect -35 -8501588 35 -8501444
rect -35 -8582556 35 -8582412
rect -35 -8663524 35 -8663380
rect -35 -8744492 35 -8744348
rect -35 -8825460 35 -8825316
rect -35 -8906428 35 -8906284
rect -35 -8987396 35 -8987252
rect -35 -9068364 35 -9068220
rect -35 -9149332 35 -9149188
rect -35 -9230300 35 -9230156
rect -35 -9311268 35 -9311124
rect -35 -9392236 35 -9392092
rect -35 -9473204 35 -9473060
rect -35 -9554172 35 -9554028
rect -35 -9635140 35 -9634996
rect -35 -9716108 35 -9715964
rect -35 -9797076 35 -9796932
rect -35 -9878044 35 -9877900
rect -35 -9959012 35 -9958868
rect -35 -10039980 35 -10039836
rect -35 -10120948 35 -10120804
rect -35 -10201916 35 -10201772
rect -35 -10282884 35 -10282740
rect -35 -10363852 35 -10363708
rect -35 -10444820 35 -10444676
rect -35 -10525788 35 -10525644
rect -35 -10606756 35 -10606612
rect -35 -10687724 35 -10687580
rect -35 -10768692 35 -10768548
rect -35 -10849660 35 -10849516
rect -35 -10930628 35 -10930484
rect -35 -11011596 35 -11011452
rect -35 -11092564 35 -11092420
rect -35 -11173532 35 -11173388
rect -35 -11254500 35 -11254356
rect -35 -11335468 35 -11335324
rect -35 -11416436 35 -11416292
rect -35 -11497404 35 -11497260
rect -35 -11578372 35 -11578228
rect -35 -11659340 35 -11659196
rect -35 -11740308 35 -11740164
rect -35 -11821276 35 -11821132
rect -35 -11902244 35 -11902100
rect -35 -11983212 35 -11983068
rect -35 -12064180 35 -12064036
rect -35 -12145148 35 -12145004
rect -35 -12226116 35 -12225972
rect -35 -12307084 35 -12306940
rect -35 -12388052 35 -12387908
rect -35 -12469020 35 -12468876
rect -35 -12549988 35 -12549844
rect -35 -12630956 35 -12630812
rect -35 -12711924 35 -12711780
rect -35 -12792892 35 -12792748
rect -35 -12873860 35 -12873716
rect -35 -12954828 35 -12954684
rect -35 -13035796 35 -13035652
rect -35 -13116764 35 -13116620
rect -35 -13197732 35 -13197588
rect -35 -13278700 35 -13278556
rect -35 -13359668 35 -13359524
rect -35 -13440636 35 -13440492
rect -35 -13521604 35 -13521460
rect -35 -13602572 35 -13602428
rect -35 -13683540 35 -13683396
rect -35 -13764508 35 -13764364
rect -35 -13845476 35 -13845332
rect -35 -13926444 35 -13926300
rect -35 -14007412 35 -14007268
rect -35 -14088380 35 -14088236
rect -35 -14169348 35 -14169204
rect -35 -14250316 35 -14250172
rect -35 -14331284 35 -14331140
rect -35 -14412252 35 -14412108
rect -35 -14493220 35 -14493076
rect -35 -14574188 35 -14574044
rect -35 -14655156 35 -14655012
rect -35 -14736124 35 -14735980
rect -35 -14817092 35 -14816948
rect -35 -14898060 35 -14897916
rect -35 -14979028 35 -14978884
rect -35 -15059996 35 -15059852
rect -35 -15140964 35 -15140820
rect -35 -15221932 35 -15221788
rect -35 -15302900 35 -15302756
rect -35 -15383868 35 -15383724
rect -35 -15464836 35 -15464692
rect -35 -15545804 35 -15545660
rect -35 -15626772 35 -15626628
rect -35 -15707740 35 -15707596
rect -35 -15788708 35 -15788564
rect -35 -15869676 35 -15869532
rect -35 -15950644 35 -15950500
rect -35 -16031612 35 -16031468
rect -35 -16112580 35 -16112436
rect -35 -16193548 35 -16193404
rect -35 -16274516 35 -16274372
rect -35 -16355484 35 -16355340
rect -35 -16436452 35 -16436308
rect -35 -16517420 35 -16517276
rect -35 -16598388 35 -16598244
rect -35 -16679356 35 -16679212
rect -35 -16760324 35 -16760180
rect -35 -16841292 35 -16841148
rect -35 -16922260 35 -16922116
rect -35 -17003228 35 -17003084
rect -35 -17084196 35 -17084052
rect -35 -17165164 35 -17165020
rect -35 -17246132 35 -17245988
rect -35 -17327100 35 -17326956
rect -35 -17408068 35 -17407924
rect -35 -17489036 35 -17488892
rect -35 -17570004 35 -17569860
rect -35 -17650972 35 -17650828
rect -35 -17731940 35 -17731796
rect -35 -17812908 35 -17812764
rect -35 -17893876 35 -17893732
rect -35 -17974844 35 -17974700
rect -35 -18055812 35 -18055668
rect -35 -18136780 35 -18136636
rect -35 -18217748 35 -18217604
rect -35 -18298716 35 -18298572
rect -35 -18379684 35 -18379540
rect -35 -18460652 35 -18460508
rect -35 -18541620 35 -18541476
rect -35 -18622588 35 -18622444
rect -35 -18703556 35 -18703412
rect -35 -18784524 35 -18784380
rect -35 -18865492 35 -18865348
rect -35 -18946460 35 -18946316
rect -35 -19027428 35 -19027284
rect -35 -19108396 35 -19108252
rect -35 -19189364 35 -19189220
rect -35 -19270332 35 -19270188
rect -35 -19351300 35 -19351156
rect -35 -19432268 35 -19432124
rect -35 -19513236 35 -19513092
rect -35 -19594204 35 -19594060
rect -35 -19675172 35 -19675028
rect -35 -19756140 35 -19755996
rect -35 -19837108 35 -19836964
rect -35 -19918076 35 -19917932
rect -35 -19999044 35 -19998900
rect -35 -20080012 35 -20079868
rect -35 -20160980 35 -20160836
<< pwell >>
rect -201 -20242114 201 20242114
<< psubdiff >>
rect -165 20242044 -69 20242078
rect 69 20242044 165 20242078
rect -165 20241982 -131 20242044
rect 131 20241982 165 20242044
rect -165 -20242044 -131 -20241982
rect 131 -20242044 165 -20241982
rect -165 -20242078 -69 -20242044
rect 69 -20242078 165 -20242044
<< psubdiffcont >>
rect -69 20242044 69 20242078
rect -165 -20241982 -131 20241982
rect 131 -20241982 165 20241982
rect -69 -20242078 69 -20242044
<< xpolycontact >>
rect -35 20241516 35 20241948
rect -35 20161084 35 20161516
rect -35 20160548 35 20160980
rect -35 20080116 35 20080548
rect -35 20079580 35 20080012
rect -35 19999148 35 19999580
rect -35 19998612 35 19999044
rect -35 19918180 35 19918612
rect -35 19917644 35 19918076
rect -35 19837212 35 19837644
rect -35 19836676 35 19837108
rect -35 19756244 35 19756676
rect -35 19755708 35 19756140
rect -35 19675276 35 19675708
rect -35 19674740 35 19675172
rect -35 19594308 35 19594740
rect -35 19593772 35 19594204
rect -35 19513340 35 19513772
rect -35 19512804 35 19513236
rect -35 19432372 35 19432804
rect -35 19431836 35 19432268
rect -35 19351404 35 19351836
rect -35 19350868 35 19351300
rect -35 19270436 35 19270868
rect -35 19269900 35 19270332
rect -35 19189468 35 19189900
rect -35 19188932 35 19189364
rect -35 19108500 35 19108932
rect -35 19107964 35 19108396
rect -35 19027532 35 19027964
rect -35 19026996 35 19027428
rect -35 18946564 35 18946996
rect -35 18946028 35 18946460
rect -35 18865596 35 18866028
rect -35 18865060 35 18865492
rect -35 18784628 35 18785060
rect -35 18784092 35 18784524
rect -35 18703660 35 18704092
rect -35 18703124 35 18703556
rect -35 18622692 35 18623124
rect -35 18622156 35 18622588
rect -35 18541724 35 18542156
rect -35 18541188 35 18541620
rect -35 18460756 35 18461188
rect -35 18460220 35 18460652
rect -35 18379788 35 18380220
rect -35 18379252 35 18379684
rect -35 18298820 35 18299252
rect -35 18298284 35 18298716
rect -35 18217852 35 18218284
rect -35 18217316 35 18217748
rect -35 18136884 35 18137316
rect -35 18136348 35 18136780
rect -35 18055916 35 18056348
rect -35 18055380 35 18055812
rect -35 17974948 35 17975380
rect -35 17974412 35 17974844
rect -35 17893980 35 17894412
rect -35 17893444 35 17893876
rect -35 17813012 35 17813444
rect -35 17812476 35 17812908
rect -35 17732044 35 17732476
rect -35 17731508 35 17731940
rect -35 17651076 35 17651508
rect -35 17650540 35 17650972
rect -35 17570108 35 17570540
rect -35 17569572 35 17570004
rect -35 17489140 35 17489572
rect -35 17488604 35 17489036
rect -35 17408172 35 17408604
rect -35 17407636 35 17408068
rect -35 17327204 35 17327636
rect -35 17326668 35 17327100
rect -35 17246236 35 17246668
rect -35 17245700 35 17246132
rect -35 17165268 35 17165700
rect -35 17164732 35 17165164
rect -35 17084300 35 17084732
rect -35 17083764 35 17084196
rect -35 17003332 35 17003764
rect -35 17002796 35 17003228
rect -35 16922364 35 16922796
rect -35 16921828 35 16922260
rect -35 16841396 35 16841828
rect -35 16840860 35 16841292
rect -35 16760428 35 16760860
rect -35 16759892 35 16760324
rect -35 16679460 35 16679892
rect -35 16678924 35 16679356
rect -35 16598492 35 16598924
rect -35 16597956 35 16598388
rect -35 16517524 35 16517956
rect -35 16516988 35 16517420
rect -35 16436556 35 16436988
rect -35 16436020 35 16436452
rect -35 16355588 35 16356020
rect -35 16355052 35 16355484
rect -35 16274620 35 16275052
rect -35 16274084 35 16274516
rect -35 16193652 35 16194084
rect -35 16193116 35 16193548
rect -35 16112684 35 16113116
rect -35 16112148 35 16112580
rect -35 16031716 35 16032148
rect -35 16031180 35 16031612
rect -35 15950748 35 15951180
rect -35 15950212 35 15950644
rect -35 15869780 35 15870212
rect -35 15869244 35 15869676
rect -35 15788812 35 15789244
rect -35 15788276 35 15788708
rect -35 15707844 35 15708276
rect -35 15707308 35 15707740
rect -35 15626876 35 15627308
rect -35 15626340 35 15626772
rect -35 15545908 35 15546340
rect -35 15545372 35 15545804
rect -35 15464940 35 15465372
rect -35 15464404 35 15464836
rect -35 15383972 35 15384404
rect -35 15383436 35 15383868
rect -35 15303004 35 15303436
rect -35 15302468 35 15302900
rect -35 15222036 35 15222468
rect -35 15221500 35 15221932
rect -35 15141068 35 15141500
rect -35 15140532 35 15140964
rect -35 15060100 35 15060532
rect -35 15059564 35 15059996
rect -35 14979132 35 14979564
rect -35 14978596 35 14979028
rect -35 14898164 35 14898596
rect -35 14897628 35 14898060
rect -35 14817196 35 14817628
rect -35 14816660 35 14817092
rect -35 14736228 35 14736660
rect -35 14735692 35 14736124
rect -35 14655260 35 14655692
rect -35 14654724 35 14655156
rect -35 14574292 35 14574724
rect -35 14573756 35 14574188
rect -35 14493324 35 14493756
rect -35 14492788 35 14493220
rect -35 14412356 35 14412788
rect -35 14411820 35 14412252
rect -35 14331388 35 14331820
rect -35 14330852 35 14331284
rect -35 14250420 35 14250852
rect -35 14249884 35 14250316
rect -35 14169452 35 14169884
rect -35 14168916 35 14169348
rect -35 14088484 35 14088916
rect -35 14087948 35 14088380
rect -35 14007516 35 14007948
rect -35 14006980 35 14007412
rect -35 13926548 35 13926980
rect -35 13926012 35 13926444
rect -35 13845580 35 13846012
rect -35 13845044 35 13845476
rect -35 13764612 35 13765044
rect -35 13764076 35 13764508
rect -35 13683644 35 13684076
rect -35 13683108 35 13683540
rect -35 13602676 35 13603108
rect -35 13602140 35 13602572
rect -35 13521708 35 13522140
rect -35 13521172 35 13521604
rect -35 13440740 35 13441172
rect -35 13440204 35 13440636
rect -35 13359772 35 13360204
rect -35 13359236 35 13359668
rect -35 13278804 35 13279236
rect -35 13278268 35 13278700
rect -35 13197836 35 13198268
rect -35 13197300 35 13197732
rect -35 13116868 35 13117300
rect -35 13116332 35 13116764
rect -35 13035900 35 13036332
rect -35 13035364 35 13035796
rect -35 12954932 35 12955364
rect -35 12954396 35 12954828
rect -35 12873964 35 12874396
rect -35 12873428 35 12873860
rect -35 12792996 35 12793428
rect -35 12792460 35 12792892
rect -35 12712028 35 12712460
rect -35 12711492 35 12711924
rect -35 12631060 35 12631492
rect -35 12630524 35 12630956
rect -35 12550092 35 12550524
rect -35 12549556 35 12549988
rect -35 12469124 35 12469556
rect -35 12468588 35 12469020
rect -35 12388156 35 12388588
rect -35 12387620 35 12388052
rect -35 12307188 35 12307620
rect -35 12306652 35 12307084
rect -35 12226220 35 12226652
rect -35 12225684 35 12226116
rect -35 12145252 35 12145684
rect -35 12144716 35 12145148
rect -35 12064284 35 12064716
rect -35 12063748 35 12064180
rect -35 11983316 35 11983748
rect -35 11982780 35 11983212
rect -35 11902348 35 11902780
rect -35 11901812 35 11902244
rect -35 11821380 35 11821812
rect -35 11820844 35 11821276
rect -35 11740412 35 11740844
rect -35 11739876 35 11740308
rect -35 11659444 35 11659876
rect -35 11658908 35 11659340
rect -35 11578476 35 11578908
rect -35 11577940 35 11578372
rect -35 11497508 35 11497940
rect -35 11496972 35 11497404
rect -35 11416540 35 11416972
rect -35 11416004 35 11416436
rect -35 11335572 35 11336004
rect -35 11335036 35 11335468
rect -35 11254604 35 11255036
rect -35 11254068 35 11254500
rect -35 11173636 35 11174068
rect -35 11173100 35 11173532
rect -35 11092668 35 11093100
rect -35 11092132 35 11092564
rect -35 11011700 35 11012132
rect -35 11011164 35 11011596
rect -35 10930732 35 10931164
rect -35 10930196 35 10930628
rect -35 10849764 35 10850196
rect -35 10849228 35 10849660
rect -35 10768796 35 10769228
rect -35 10768260 35 10768692
rect -35 10687828 35 10688260
rect -35 10687292 35 10687724
rect -35 10606860 35 10607292
rect -35 10606324 35 10606756
rect -35 10525892 35 10526324
rect -35 10525356 35 10525788
rect -35 10444924 35 10445356
rect -35 10444388 35 10444820
rect -35 10363956 35 10364388
rect -35 10363420 35 10363852
rect -35 10282988 35 10283420
rect -35 10282452 35 10282884
rect -35 10202020 35 10202452
rect -35 10201484 35 10201916
rect -35 10121052 35 10121484
rect -35 10120516 35 10120948
rect -35 10040084 35 10040516
rect -35 10039548 35 10039980
rect -35 9959116 35 9959548
rect -35 9958580 35 9959012
rect -35 9878148 35 9878580
rect -35 9877612 35 9878044
rect -35 9797180 35 9797612
rect -35 9796644 35 9797076
rect -35 9716212 35 9716644
rect -35 9715676 35 9716108
rect -35 9635244 35 9635676
rect -35 9634708 35 9635140
rect -35 9554276 35 9554708
rect -35 9553740 35 9554172
rect -35 9473308 35 9473740
rect -35 9472772 35 9473204
rect -35 9392340 35 9392772
rect -35 9391804 35 9392236
rect -35 9311372 35 9311804
rect -35 9310836 35 9311268
rect -35 9230404 35 9230836
rect -35 9229868 35 9230300
rect -35 9149436 35 9149868
rect -35 9148900 35 9149332
rect -35 9068468 35 9068900
rect -35 9067932 35 9068364
rect -35 8987500 35 8987932
rect -35 8986964 35 8987396
rect -35 8906532 35 8906964
rect -35 8905996 35 8906428
rect -35 8825564 35 8825996
rect -35 8825028 35 8825460
rect -35 8744596 35 8745028
rect -35 8744060 35 8744492
rect -35 8663628 35 8664060
rect -35 8663092 35 8663524
rect -35 8582660 35 8583092
rect -35 8582124 35 8582556
rect -35 8501692 35 8502124
rect -35 8501156 35 8501588
rect -35 8420724 35 8421156
rect -35 8420188 35 8420620
rect -35 8339756 35 8340188
rect -35 8339220 35 8339652
rect -35 8258788 35 8259220
rect -35 8258252 35 8258684
rect -35 8177820 35 8178252
rect -35 8177284 35 8177716
rect -35 8096852 35 8097284
rect -35 8096316 35 8096748
rect -35 8015884 35 8016316
rect -35 8015348 35 8015780
rect -35 7934916 35 7935348
rect -35 7934380 35 7934812
rect -35 7853948 35 7854380
rect -35 7853412 35 7853844
rect -35 7772980 35 7773412
rect -35 7772444 35 7772876
rect -35 7692012 35 7692444
rect -35 7691476 35 7691908
rect -35 7611044 35 7611476
rect -35 7610508 35 7610940
rect -35 7530076 35 7530508
rect -35 7529540 35 7529972
rect -35 7449108 35 7449540
rect -35 7448572 35 7449004
rect -35 7368140 35 7368572
rect -35 7367604 35 7368036
rect -35 7287172 35 7287604
rect -35 7286636 35 7287068
rect -35 7206204 35 7206636
rect -35 7205668 35 7206100
rect -35 7125236 35 7125668
rect -35 7124700 35 7125132
rect -35 7044268 35 7044700
rect -35 7043732 35 7044164
rect -35 6963300 35 6963732
rect -35 6962764 35 6963196
rect -35 6882332 35 6882764
rect -35 6881796 35 6882228
rect -35 6801364 35 6801796
rect -35 6800828 35 6801260
rect -35 6720396 35 6720828
rect -35 6719860 35 6720292
rect -35 6639428 35 6639860
rect -35 6638892 35 6639324
rect -35 6558460 35 6558892
rect -35 6557924 35 6558356
rect -35 6477492 35 6477924
rect -35 6476956 35 6477388
rect -35 6396524 35 6396956
rect -35 6395988 35 6396420
rect -35 6315556 35 6315988
rect -35 6315020 35 6315452
rect -35 6234588 35 6235020
rect -35 6234052 35 6234484
rect -35 6153620 35 6154052
rect -35 6153084 35 6153516
rect -35 6072652 35 6073084
rect -35 6072116 35 6072548
rect -35 5991684 35 5992116
rect -35 5991148 35 5991580
rect -35 5910716 35 5911148
rect -35 5910180 35 5910612
rect -35 5829748 35 5830180
rect -35 5829212 35 5829644
rect -35 5748780 35 5749212
rect -35 5748244 35 5748676
rect -35 5667812 35 5668244
rect -35 5667276 35 5667708
rect -35 5586844 35 5587276
rect -35 5586308 35 5586740
rect -35 5505876 35 5506308
rect -35 5505340 35 5505772
rect -35 5424908 35 5425340
rect -35 5424372 35 5424804
rect -35 5343940 35 5344372
rect -35 5343404 35 5343836
rect -35 5262972 35 5263404
rect -35 5262436 35 5262868
rect -35 5182004 35 5182436
rect -35 5181468 35 5181900
rect -35 5101036 35 5101468
rect -35 5100500 35 5100932
rect -35 5020068 35 5020500
rect -35 5019532 35 5019964
rect -35 4939100 35 4939532
rect -35 4938564 35 4938996
rect -35 4858132 35 4858564
rect -35 4857596 35 4858028
rect -35 4777164 35 4777596
rect -35 4776628 35 4777060
rect -35 4696196 35 4696628
rect -35 4695660 35 4696092
rect -35 4615228 35 4615660
rect -35 4614692 35 4615124
rect -35 4534260 35 4534692
rect -35 4533724 35 4534156
rect -35 4453292 35 4453724
rect -35 4452756 35 4453188
rect -35 4372324 35 4372756
rect -35 4371788 35 4372220
rect -35 4291356 35 4291788
rect -35 4290820 35 4291252
rect -35 4210388 35 4210820
rect -35 4209852 35 4210284
rect -35 4129420 35 4129852
rect -35 4128884 35 4129316
rect -35 4048452 35 4048884
rect -35 4047916 35 4048348
rect -35 3967484 35 3967916
rect -35 3966948 35 3967380
rect -35 3886516 35 3886948
rect -35 3885980 35 3886412
rect -35 3805548 35 3805980
rect -35 3805012 35 3805444
rect -35 3724580 35 3725012
rect -35 3724044 35 3724476
rect -35 3643612 35 3644044
rect -35 3643076 35 3643508
rect -35 3562644 35 3563076
rect -35 3562108 35 3562540
rect -35 3481676 35 3482108
rect -35 3481140 35 3481572
rect -35 3400708 35 3401140
rect -35 3400172 35 3400604
rect -35 3319740 35 3320172
rect -35 3319204 35 3319636
rect -35 3238772 35 3239204
rect -35 3238236 35 3238668
rect -35 3157804 35 3158236
rect -35 3157268 35 3157700
rect -35 3076836 35 3077268
rect -35 3076300 35 3076732
rect -35 2995868 35 2996300
rect -35 2995332 35 2995764
rect -35 2914900 35 2915332
rect -35 2914364 35 2914796
rect -35 2833932 35 2834364
rect -35 2833396 35 2833828
rect -35 2752964 35 2753396
rect -35 2752428 35 2752860
rect -35 2671996 35 2672428
rect -35 2671460 35 2671892
rect -35 2591028 35 2591460
rect -35 2590492 35 2590924
rect -35 2510060 35 2510492
rect -35 2509524 35 2509956
rect -35 2429092 35 2429524
rect -35 2428556 35 2428988
rect -35 2348124 35 2348556
rect -35 2347588 35 2348020
rect -35 2267156 35 2267588
rect -35 2266620 35 2267052
rect -35 2186188 35 2186620
rect -35 2185652 35 2186084
rect -35 2105220 35 2105652
rect -35 2104684 35 2105116
rect -35 2024252 35 2024684
rect -35 2023716 35 2024148
rect -35 1943284 35 1943716
rect -35 1942748 35 1943180
rect -35 1862316 35 1862748
rect -35 1861780 35 1862212
rect -35 1781348 35 1781780
rect -35 1780812 35 1781244
rect -35 1700380 35 1700812
rect -35 1699844 35 1700276
rect -35 1619412 35 1619844
rect -35 1618876 35 1619308
rect -35 1538444 35 1538876
rect -35 1537908 35 1538340
rect -35 1457476 35 1457908
rect -35 1456940 35 1457372
rect -35 1376508 35 1376940
rect -35 1375972 35 1376404
rect -35 1295540 35 1295972
rect -35 1295004 35 1295436
rect -35 1214572 35 1215004
rect -35 1214036 35 1214468
rect -35 1133604 35 1134036
rect -35 1133068 35 1133500
rect -35 1052636 35 1053068
rect -35 1052100 35 1052532
rect -35 971668 35 972100
rect -35 971132 35 971564
rect -35 890700 35 891132
rect -35 890164 35 890596
rect -35 809732 35 810164
rect -35 809196 35 809628
rect -35 728764 35 729196
rect -35 728228 35 728660
rect -35 647796 35 648228
rect -35 647260 35 647692
rect -35 566828 35 567260
rect -35 566292 35 566724
rect -35 485860 35 486292
rect -35 485324 35 485756
rect -35 404892 35 405324
rect -35 404356 35 404788
rect -35 323924 35 324356
rect -35 323388 35 323820
rect -35 242956 35 243388
rect -35 242420 35 242852
rect -35 161988 35 162420
rect -35 161452 35 161884
rect -35 81020 35 81452
rect -35 80484 35 80916
rect -35 52 35 484
rect -35 -484 35 -52
rect -35 -80916 35 -80484
rect -35 -81452 35 -81020
rect -35 -161884 35 -161452
rect -35 -162420 35 -161988
rect -35 -242852 35 -242420
rect -35 -243388 35 -242956
rect -35 -323820 35 -323388
rect -35 -324356 35 -323924
rect -35 -404788 35 -404356
rect -35 -405324 35 -404892
rect -35 -485756 35 -485324
rect -35 -486292 35 -485860
rect -35 -566724 35 -566292
rect -35 -567260 35 -566828
rect -35 -647692 35 -647260
rect -35 -648228 35 -647796
rect -35 -728660 35 -728228
rect -35 -729196 35 -728764
rect -35 -809628 35 -809196
rect -35 -810164 35 -809732
rect -35 -890596 35 -890164
rect -35 -891132 35 -890700
rect -35 -971564 35 -971132
rect -35 -972100 35 -971668
rect -35 -1052532 35 -1052100
rect -35 -1053068 35 -1052636
rect -35 -1133500 35 -1133068
rect -35 -1134036 35 -1133604
rect -35 -1214468 35 -1214036
rect -35 -1215004 35 -1214572
rect -35 -1295436 35 -1295004
rect -35 -1295972 35 -1295540
rect -35 -1376404 35 -1375972
rect -35 -1376940 35 -1376508
rect -35 -1457372 35 -1456940
rect -35 -1457908 35 -1457476
rect -35 -1538340 35 -1537908
rect -35 -1538876 35 -1538444
rect -35 -1619308 35 -1618876
rect -35 -1619844 35 -1619412
rect -35 -1700276 35 -1699844
rect -35 -1700812 35 -1700380
rect -35 -1781244 35 -1780812
rect -35 -1781780 35 -1781348
rect -35 -1862212 35 -1861780
rect -35 -1862748 35 -1862316
rect -35 -1943180 35 -1942748
rect -35 -1943716 35 -1943284
rect -35 -2024148 35 -2023716
rect -35 -2024684 35 -2024252
rect -35 -2105116 35 -2104684
rect -35 -2105652 35 -2105220
rect -35 -2186084 35 -2185652
rect -35 -2186620 35 -2186188
rect -35 -2267052 35 -2266620
rect -35 -2267588 35 -2267156
rect -35 -2348020 35 -2347588
rect -35 -2348556 35 -2348124
rect -35 -2428988 35 -2428556
rect -35 -2429524 35 -2429092
rect -35 -2509956 35 -2509524
rect -35 -2510492 35 -2510060
rect -35 -2590924 35 -2590492
rect -35 -2591460 35 -2591028
rect -35 -2671892 35 -2671460
rect -35 -2672428 35 -2671996
rect -35 -2752860 35 -2752428
rect -35 -2753396 35 -2752964
rect -35 -2833828 35 -2833396
rect -35 -2834364 35 -2833932
rect -35 -2914796 35 -2914364
rect -35 -2915332 35 -2914900
rect -35 -2995764 35 -2995332
rect -35 -2996300 35 -2995868
rect -35 -3076732 35 -3076300
rect -35 -3077268 35 -3076836
rect -35 -3157700 35 -3157268
rect -35 -3158236 35 -3157804
rect -35 -3238668 35 -3238236
rect -35 -3239204 35 -3238772
rect -35 -3319636 35 -3319204
rect -35 -3320172 35 -3319740
rect -35 -3400604 35 -3400172
rect -35 -3401140 35 -3400708
rect -35 -3481572 35 -3481140
rect -35 -3482108 35 -3481676
rect -35 -3562540 35 -3562108
rect -35 -3563076 35 -3562644
rect -35 -3643508 35 -3643076
rect -35 -3644044 35 -3643612
rect -35 -3724476 35 -3724044
rect -35 -3725012 35 -3724580
rect -35 -3805444 35 -3805012
rect -35 -3805980 35 -3805548
rect -35 -3886412 35 -3885980
rect -35 -3886948 35 -3886516
rect -35 -3967380 35 -3966948
rect -35 -3967916 35 -3967484
rect -35 -4048348 35 -4047916
rect -35 -4048884 35 -4048452
rect -35 -4129316 35 -4128884
rect -35 -4129852 35 -4129420
rect -35 -4210284 35 -4209852
rect -35 -4210820 35 -4210388
rect -35 -4291252 35 -4290820
rect -35 -4291788 35 -4291356
rect -35 -4372220 35 -4371788
rect -35 -4372756 35 -4372324
rect -35 -4453188 35 -4452756
rect -35 -4453724 35 -4453292
rect -35 -4534156 35 -4533724
rect -35 -4534692 35 -4534260
rect -35 -4615124 35 -4614692
rect -35 -4615660 35 -4615228
rect -35 -4696092 35 -4695660
rect -35 -4696628 35 -4696196
rect -35 -4777060 35 -4776628
rect -35 -4777596 35 -4777164
rect -35 -4858028 35 -4857596
rect -35 -4858564 35 -4858132
rect -35 -4938996 35 -4938564
rect -35 -4939532 35 -4939100
rect -35 -5019964 35 -5019532
rect -35 -5020500 35 -5020068
rect -35 -5100932 35 -5100500
rect -35 -5101468 35 -5101036
rect -35 -5181900 35 -5181468
rect -35 -5182436 35 -5182004
rect -35 -5262868 35 -5262436
rect -35 -5263404 35 -5262972
rect -35 -5343836 35 -5343404
rect -35 -5344372 35 -5343940
rect -35 -5424804 35 -5424372
rect -35 -5425340 35 -5424908
rect -35 -5505772 35 -5505340
rect -35 -5506308 35 -5505876
rect -35 -5586740 35 -5586308
rect -35 -5587276 35 -5586844
rect -35 -5667708 35 -5667276
rect -35 -5668244 35 -5667812
rect -35 -5748676 35 -5748244
rect -35 -5749212 35 -5748780
rect -35 -5829644 35 -5829212
rect -35 -5830180 35 -5829748
rect -35 -5910612 35 -5910180
rect -35 -5911148 35 -5910716
rect -35 -5991580 35 -5991148
rect -35 -5992116 35 -5991684
rect -35 -6072548 35 -6072116
rect -35 -6073084 35 -6072652
rect -35 -6153516 35 -6153084
rect -35 -6154052 35 -6153620
rect -35 -6234484 35 -6234052
rect -35 -6235020 35 -6234588
rect -35 -6315452 35 -6315020
rect -35 -6315988 35 -6315556
rect -35 -6396420 35 -6395988
rect -35 -6396956 35 -6396524
rect -35 -6477388 35 -6476956
rect -35 -6477924 35 -6477492
rect -35 -6558356 35 -6557924
rect -35 -6558892 35 -6558460
rect -35 -6639324 35 -6638892
rect -35 -6639860 35 -6639428
rect -35 -6720292 35 -6719860
rect -35 -6720828 35 -6720396
rect -35 -6801260 35 -6800828
rect -35 -6801796 35 -6801364
rect -35 -6882228 35 -6881796
rect -35 -6882764 35 -6882332
rect -35 -6963196 35 -6962764
rect -35 -6963732 35 -6963300
rect -35 -7044164 35 -7043732
rect -35 -7044700 35 -7044268
rect -35 -7125132 35 -7124700
rect -35 -7125668 35 -7125236
rect -35 -7206100 35 -7205668
rect -35 -7206636 35 -7206204
rect -35 -7287068 35 -7286636
rect -35 -7287604 35 -7287172
rect -35 -7368036 35 -7367604
rect -35 -7368572 35 -7368140
rect -35 -7449004 35 -7448572
rect -35 -7449540 35 -7449108
rect -35 -7529972 35 -7529540
rect -35 -7530508 35 -7530076
rect -35 -7610940 35 -7610508
rect -35 -7611476 35 -7611044
rect -35 -7691908 35 -7691476
rect -35 -7692444 35 -7692012
rect -35 -7772876 35 -7772444
rect -35 -7773412 35 -7772980
rect -35 -7853844 35 -7853412
rect -35 -7854380 35 -7853948
rect -35 -7934812 35 -7934380
rect -35 -7935348 35 -7934916
rect -35 -8015780 35 -8015348
rect -35 -8016316 35 -8015884
rect -35 -8096748 35 -8096316
rect -35 -8097284 35 -8096852
rect -35 -8177716 35 -8177284
rect -35 -8178252 35 -8177820
rect -35 -8258684 35 -8258252
rect -35 -8259220 35 -8258788
rect -35 -8339652 35 -8339220
rect -35 -8340188 35 -8339756
rect -35 -8420620 35 -8420188
rect -35 -8421156 35 -8420724
rect -35 -8501588 35 -8501156
rect -35 -8502124 35 -8501692
rect -35 -8582556 35 -8582124
rect -35 -8583092 35 -8582660
rect -35 -8663524 35 -8663092
rect -35 -8664060 35 -8663628
rect -35 -8744492 35 -8744060
rect -35 -8745028 35 -8744596
rect -35 -8825460 35 -8825028
rect -35 -8825996 35 -8825564
rect -35 -8906428 35 -8905996
rect -35 -8906964 35 -8906532
rect -35 -8987396 35 -8986964
rect -35 -8987932 35 -8987500
rect -35 -9068364 35 -9067932
rect -35 -9068900 35 -9068468
rect -35 -9149332 35 -9148900
rect -35 -9149868 35 -9149436
rect -35 -9230300 35 -9229868
rect -35 -9230836 35 -9230404
rect -35 -9311268 35 -9310836
rect -35 -9311804 35 -9311372
rect -35 -9392236 35 -9391804
rect -35 -9392772 35 -9392340
rect -35 -9473204 35 -9472772
rect -35 -9473740 35 -9473308
rect -35 -9554172 35 -9553740
rect -35 -9554708 35 -9554276
rect -35 -9635140 35 -9634708
rect -35 -9635676 35 -9635244
rect -35 -9716108 35 -9715676
rect -35 -9716644 35 -9716212
rect -35 -9797076 35 -9796644
rect -35 -9797612 35 -9797180
rect -35 -9878044 35 -9877612
rect -35 -9878580 35 -9878148
rect -35 -9959012 35 -9958580
rect -35 -9959548 35 -9959116
rect -35 -10039980 35 -10039548
rect -35 -10040516 35 -10040084
rect -35 -10120948 35 -10120516
rect -35 -10121484 35 -10121052
rect -35 -10201916 35 -10201484
rect -35 -10202452 35 -10202020
rect -35 -10282884 35 -10282452
rect -35 -10283420 35 -10282988
rect -35 -10363852 35 -10363420
rect -35 -10364388 35 -10363956
rect -35 -10444820 35 -10444388
rect -35 -10445356 35 -10444924
rect -35 -10525788 35 -10525356
rect -35 -10526324 35 -10525892
rect -35 -10606756 35 -10606324
rect -35 -10607292 35 -10606860
rect -35 -10687724 35 -10687292
rect -35 -10688260 35 -10687828
rect -35 -10768692 35 -10768260
rect -35 -10769228 35 -10768796
rect -35 -10849660 35 -10849228
rect -35 -10850196 35 -10849764
rect -35 -10930628 35 -10930196
rect -35 -10931164 35 -10930732
rect -35 -11011596 35 -11011164
rect -35 -11012132 35 -11011700
rect -35 -11092564 35 -11092132
rect -35 -11093100 35 -11092668
rect -35 -11173532 35 -11173100
rect -35 -11174068 35 -11173636
rect -35 -11254500 35 -11254068
rect -35 -11255036 35 -11254604
rect -35 -11335468 35 -11335036
rect -35 -11336004 35 -11335572
rect -35 -11416436 35 -11416004
rect -35 -11416972 35 -11416540
rect -35 -11497404 35 -11496972
rect -35 -11497940 35 -11497508
rect -35 -11578372 35 -11577940
rect -35 -11578908 35 -11578476
rect -35 -11659340 35 -11658908
rect -35 -11659876 35 -11659444
rect -35 -11740308 35 -11739876
rect -35 -11740844 35 -11740412
rect -35 -11821276 35 -11820844
rect -35 -11821812 35 -11821380
rect -35 -11902244 35 -11901812
rect -35 -11902780 35 -11902348
rect -35 -11983212 35 -11982780
rect -35 -11983748 35 -11983316
rect -35 -12064180 35 -12063748
rect -35 -12064716 35 -12064284
rect -35 -12145148 35 -12144716
rect -35 -12145684 35 -12145252
rect -35 -12226116 35 -12225684
rect -35 -12226652 35 -12226220
rect -35 -12307084 35 -12306652
rect -35 -12307620 35 -12307188
rect -35 -12388052 35 -12387620
rect -35 -12388588 35 -12388156
rect -35 -12469020 35 -12468588
rect -35 -12469556 35 -12469124
rect -35 -12549988 35 -12549556
rect -35 -12550524 35 -12550092
rect -35 -12630956 35 -12630524
rect -35 -12631492 35 -12631060
rect -35 -12711924 35 -12711492
rect -35 -12712460 35 -12712028
rect -35 -12792892 35 -12792460
rect -35 -12793428 35 -12792996
rect -35 -12873860 35 -12873428
rect -35 -12874396 35 -12873964
rect -35 -12954828 35 -12954396
rect -35 -12955364 35 -12954932
rect -35 -13035796 35 -13035364
rect -35 -13036332 35 -13035900
rect -35 -13116764 35 -13116332
rect -35 -13117300 35 -13116868
rect -35 -13197732 35 -13197300
rect -35 -13198268 35 -13197836
rect -35 -13278700 35 -13278268
rect -35 -13279236 35 -13278804
rect -35 -13359668 35 -13359236
rect -35 -13360204 35 -13359772
rect -35 -13440636 35 -13440204
rect -35 -13441172 35 -13440740
rect -35 -13521604 35 -13521172
rect -35 -13522140 35 -13521708
rect -35 -13602572 35 -13602140
rect -35 -13603108 35 -13602676
rect -35 -13683540 35 -13683108
rect -35 -13684076 35 -13683644
rect -35 -13764508 35 -13764076
rect -35 -13765044 35 -13764612
rect -35 -13845476 35 -13845044
rect -35 -13846012 35 -13845580
rect -35 -13926444 35 -13926012
rect -35 -13926980 35 -13926548
rect -35 -14007412 35 -14006980
rect -35 -14007948 35 -14007516
rect -35 -14088380 35 -14087948
rect -35 -14088916 35 -14088484
rect -35 -14169348 35 -14168916
rect -35 -14169884 35 -14169452
rect -35 -14250316 35 -14249884
rect -35 -14250852 35 -14250420
rect -35 -14331284 35 -14330852
rect -35 -14331820 35 -14331388
rect -35 -14412252 35 -14411820
rect -35 -14412788 35 -14412356
rect -35 -14493220 35 -14492788
rect -35 -14493756 35 -14493324
rect -35 -14574188 35 -14573756
rect -35 -14574724 35 -14574292
rect -35 -14655156 35 -14654724
rect -35 -14655692 35 -14655260
rect -35 -14736124 35 -14735692
rect -35 -14736660 35 -14736228
rect -35 -14817092 35 -14816660
rect -35 -14817628 35 -14817196
rect -35 -14898060 35 -14897628
rect -35 -14898596 35 -14898164
rect -35 -14979028 35 -14978596
rect -35 -14979564 35 -14979132
rect -35 -15059996 35 -15059564
rect -35 -15060532 35 -15060100
rect -35 -15140964 35 -15140532
rect -35 -15141500 35 -15141068
rect -35 -15221932 35 -15221500
rect -35 -15222468 35 -15222036
rect -35 -15302900 35 -15302468
rect -35 -15303436 35 -15303004
rect -35 -15383868 35 -15383436
rect -35 -15384404 35 -15383972
rect -35 -15464836 35 -15464404
rect -35 -15465372 35 -15464940
rect -35 -15545804 35 -15545372
rect -35 -15546340 35 -15545908
rect -35 -15626772 35 -15626340
rect -35 -15627308 35 -15626876
rect -35 -15707740 35 -15707308
rect -35 -15708276 35 -15707844
rect -35 -15788708 35 -15788276
rect -35 -15789244 35 -15788812
rect -35 -15869676 35 -15869244
rect -35 -15870212 35 -15869780
rect -35 -15950644 35 -15950212
rect -35 -15951180 35 -15950748
rect -35 -16031612 35 -16031180
rect -35 -16032148 35 -16031716
rect -35 -16112580 35 -16112148
rect -35 -16113116 35 -16112684
rect -35 -16193548 35 -16193116
rect -35 -16194084 35 -16193652
rect -35 -16274516 35 -16274084
rect -35 -16275052 35 -16274620
rect -35 -16355484 35 -16355052
rect -35 -16356020 35 -16355588
rect -35 -16436452 35 -16436020
rect -35 -16436988 35 -16436556
rect -35 -16517420 35 -16516988
rect -35 -16517956 35 -16517524
rect -35 -16598388 35 -16597956
rect -35 -16598924 35 -16598492
rect -35 -16679356 35 -16678924
rect -35 -16679892 35 -16679460
rect -35 -16760324 35 -16759892
rect -35 -16760860 35 -16760428
rect -35 -16841292 35 -16840860
rect -35 -16841828 35 -16841396
rect -35 -16922260 35 -16921828
rect -35 -16922796 35 -16922364
rect -35 -17003228 35 -17002796
rect -35 -17003764 35 -17003332
rect -35 -17084196 35 -17083764
rect -35 -17084732 35 -17084300
rect -35 -17165164 35 -17164732
rect -35 -17165700 35 -17165268
rect -35 -17246132 35 -17245700
rect -35 -17246668 35 -17246236
rect -35 -17327100 35 -17326668
rect -35 -17327636 35 -17327204
rect -35 -17408068 35 -17407636
rect -35 -17408604 35 -17408172
rect -35 -17489036 35 -17488604
rect -35 -17489572 35 -17489140
rect -35 -17570004 35 -17569572
rect -35 -17570540 35 -17570108
rect -35 -17650972 35 -17650540
rect -35 -17651508 35 -17651076
rect -35 -17731940 35 -17731508
rect -35 -17732476 35 -17732044
rect -35 -17812908 35 -17812476
rect -35 -17813444 35 -17813012
rect -35 -17893876 35 -17893444
rect -35 -17894412 35 -17893980
rect -35 -17974844 35 -17974412
rect -35 -17975380 35 -17974948
rect -35 -18055812 35 -18055380
rect -35 -18056348 35 -18055916
rect -35 -18136780 35 -18136348
rect -35 -18137316 35 -18136884
rect -35 -18217748 35 -18217316
rect -35 -18218284 35 -18217852
rect -35 -18298716 35 -18298284
rect -35 -18299252 35 -18298820
rect -35 -18379684 35 -18379252
rect -35 -18380220 35 -18379788
rect -35 -18460652 35 -18460220
rect -35 -18461188 35 -18460756
rect -35 -18541620 35 -18541188
rect -35 -18542156 35 -18541724
rect -35 -18622588 35 -18622156
rect -35 -18623124 35 -18622692
rect -35 -18703556 35 -18703124
rect -35 -18704092 35 -18703660
rect -35 -18784524 35 -18784092
rect -35 -18785060 35 -18784628
rect -35 -18865492 35 -18865060
rect -35 -18866028 35 -18865596
rect -35 -18946460 35 -18946028
rect -35 -18946996 35 -18946564
rect -35 -19027428 35 -19026996
rect -35 -19027964 35 -19027532
rect -35 -19108396 35 -19107964
rect -35 -19108932 35 -19108500
rect -35 -19189364 35 -19188932
rect -35 -19189900 35 -19189468
rect -35 -19270332 35 -19269900
rect -35 -19270868 35 -19270436
rect -35 -19351300 35 -19350868
rect -35 -19351836 35 -19351404
rect -35 -19432268 35 -19431836
rect -35 -19432804 35 -19432372
rect -35 -19513236 35 -19512804
rect -35 -19513772 35 -19513340
rect -35 -19594204 35 -19593772
rect -35 -19594740 35 -19594308
rect -35 -19675172 35 -19674740
rect -35 -19675708 35 -19675276
rect -35 -19756140 35 -19755708
rect -35 -19756676 35 -19756244
rect -35 -19837108 35 -19836676
rect -35 -19837644 35 -19837212
rect -35 -19918076 35 -19917644
rect -35 -19918612 35 -19918180
rect -35 -19999044 35 -19998612
rect -35 -19999580 35 -19999148
rect -35 -20080012 35 -20079580
rect -35 -20080548 35 -20080116
rect -35 -20160980 35 -20160548
rect -35 -20161516 35 -20161084
rect -35 -20241948 35 -20241516
<< xpolyres >>
rect -35 20161516 35 20241516
rect -35 20080548 35 20160548
rect -35 19999580 35 20079580
rect -35 19918612 35 19998612
rect -35 19837644 35 19917644
rect -35 19756676 35 19836676
rect -35 19675708 35 19755708
rect -35 19594740 35 19674740
rect -35 19513772 35 19593772
rect -35 19432804 35 19512804
rect -35 19351836 35 19431836
rect -35 19270868 35 19350868
rect -35 19189900 35 19269900
rect -35 19108932 35 19188932
rect -35 19027964 35 19107964
rect -35 18946996 35 19026996
rect -35 18866028 35 18946028
rect -35 18785060 35 18865060
rect -35 18704092 35 18784092
rect -35 18623124 35 18703124
rect -35 18542156 35 18622156
rect -35 18461188 35 18541188
rect -35 18380220 35 18460220
rect -35 18299252 35 18379252
rect -35 18218284 35 18298284
rect -35 18137316 35 18217316
rect -35 18056348 35 18136348
rect -35 17975380 35 18055380
rect -35 17894412 35 17974412
rect -35 17813444 35 17893444
rect -35 17732476 35 17812476
rect -35 17651508 35 17731508
rect -35 17570540 35 17650540
rect -35 17489572 35 17569572
rect -35 17408604 35 17488604
rect -35 17327636 35 17407636
rect -35 17246668 35 17326668
rect -35 17165700 35 17245700
rect -35 17084732 35 17164732
rect -35 17003764 35 17083764
rect -35 16922796 35 17002796
rect -35 16841828 35 16921828
rect -35 16760860 35 16840860
rect -35 16679892 35 16759892
rect -35 16598924 35 16678924
rect -35 16517956 35 16597956
rect -35 16436988 35 16516988
rect -35 16356020 35 16436020
rect -35 16275052 35 16355052
rect -35 16194084 35 16274084
rect -35 16113116 35 16193116
rect -35 16032148 35 16112148
rect -35 15951180 35 16031180
rect -35 15870212 35 15950212
rect -35 15789244 35 15869244
rect -35 15708276 35 15788276
rect -35 15627308 35 15707308
rect -35 15546340 35 15626340
rect -35 15465372 35 15545372
rect -35 15384404 35 15464404
rect -35 15303436 35 15383436
rect -35 15222468 35 15302468
rect -35 15141500 35 15221500
rect -35 15060532 35 15140532
rect -35 14979564 35 15059564
rect -35 14898596 35 14978596
rect -35 14817628 35 14897628
rect -35 14736660 35 14816660
rect -35 14655692 35 14735692
rect -35 14574724 35 14654724
rect -35 14493756 35 14573756
rect -35 14412788 35 14492788
rect -35 14331820 35 14411820
rect -35 14250852 35 14330852
rect -35 14169884 35 14249884
rect -35 14088916 35 14168916
rect -35 14007948 35 14087948
rect -35 13926980 35 14006980
rect -35 13846012 35 13926012
rect -35 13765044 35 13845044
rect -35 13684076 35 13764076
rect -35 13603108 35 13683108
rect -35 13522140 35 13602140
rect -35 13441172 35 13521172
rect -35 13360204 35 13440204
rect -35 13279236 35 13359236
rect -35 13198268 35 13278268
rect -35 13117300 35 13197300
rect -35 13036332 35 13116332
rect -35 12955364 35 13035364
rect -35 12874396 35 12954396
rect -35 12793428 35 12873428
rect -35 12712460 35 12792460
rect -35 12631492 35 12711492
rect -35 12550524 35 12630524
rect -35 12469556 35 12549556
rect -35 12388588 35 12468588
rect -35 12307620 35 12387620
rect -35 12226652 35 12306652
rect -35 12145684 35 12225684
rect -35 12064716 35 12144716
rect -35 11983748 35 12063748
rect -35 11902780 35 11982780
rect -35 11821812 35 11901812
rect -35 11740844 35 11820844
rect -35 11659876 35 11739876
rect -35 11578908 35 11658908
rect -35 11497940 35 11577940
rect -35 11416972 35 11496972
rect -35 11336004 35 11416004
rect -35 11255036 35 11335036
rect -35 11174068 35 11254068
rect -35 11093100 35 11173100
rect -35 11012132 35 11092132
rect -35 10931164 35 11011164
rect -35 10850196 35 10930196
rect -35 10769228 35 10849228
rect -35 10688260 35 10768260
rect -35 10607292 35 10687292
rect -35 10526324 35 10606324
rect -35 10445356 35 10525356
rect -35 10364388 35 10444388
rect -35 10283420 35 10363420
rect -35 10202452 35 10282452
rect -35 10121484 35 10201484
rect -35 10040516 35 10120516
rect -35 9959548 35 10039548
rect -35 9878580 35 9958580
rect -35 9797612 35 9877612
rect -35 9716644 35 9796644
rect -35 9635676 35 9715676
rect -35 9554708 35 9634708
rect -35 9473740 35 9553740
rect -35 9392772 35 9472772
rect -35 9311804 35 9391804
rect -35 9230836 35 9310836
rect -35 9149868 35 9229868
rect -35 9068900 35 9148900
rect -35 8987932 35 9067932
rect -35 8906964 35 8986964
rect -35 8825996 35 8905996
rect -35 8745028 35 8825028
rect -35 8664060 35 8744060
rect -35 8583092 35 8663092
rect -35 8502124 35 8582124
rect -35 8421156 35 8501156
rect -35 8340188 35 8420188
rect -35 8259220 35 8339220
rect -35 8178252 35 8258252
rect -35 8097284 35 8177284
rect -35 8016316 35 8096316
rect -35 7935348 35 8015348
rect -35 7854380 35 7934380
rect -35 7773412 35 7853412
rect -35 7692444 35 7772444
rect -35 7611476 35 7691476
rect -35 7530508 35 7610508
rect -35 7449540 35 7529540
rect -35 7368572 35 7448572
rect -35 7287604 35 7367604
rect -35 7206636 35 7286636
rect -35 7125668 35 7205668
rect -35 7044700 35 7124700
rect -35 6963732 35 7043732
rect -35 6882764 35 6962764
rect -35 6801796 35 6881796
rect -35 6720828 35 6800828
rect -35 6639860 35 6719860
rect -35 6558892 35 6638892
rect -35 6477924 35 6557924
rect -35 6396956 35 6476956
rect -35 6315988 35 6395988
rect -35 6235020 35 6315020
rect -35 6154052 35 6234052
rect -35 6073084 35 6153084
rect -35 5992116 35 6072116
rect -35 5911148 35 5991148
rect -35 5830180 35 5910180
rect -35 5749212 35 5829212
rect -35 5668244 35 5748244
rect -35 5587276 35 5667276
rect -35 5506308 35 5586308
rect -35 5425340 35 5505340
rect -35 5344372 35 5424372
rect -35 5263404 35 5343404
rect -35 5182436 35 5262436
rect -35 5101468 35 5181468
rect -35 5020500 35 5100500
rect -35 4939532 35 5019532
rect -35 4858564 35 4938564
rect -35 4777596 35 4857596
rect -35 4696628 35 4776628
rect -35 4615660 35 4695660
rect -35 4534692 35 4614692
rect -35 4453724 35 4533724
rect -35 4372756 35 4452756
rect -35 4291788 35 4371788
rect -35 4210820 35 4290820
rect -35 4129852 35 4209852
rect -35 4048884 35 4128884
rect -35 3967916 35 4047916
rect -35 3886948 35 3966948
rect -35 3805980 35 3885980
rect -35 3725012 35 3805012
rect -35 3644044 35 3724044
rect -35 3563076 35 3643076
rect -35 3482108 35 3562108
rect -35 3401140 35 3481140
rect -35 3320172 35 3400172
rect -35 3239204 35 3319204
rect -35 3158236 35 3238236
rect -35 3077268 35 3157268
rect -35 2996300 35 3076300
rect -35 2915332 35 2995332
rect -35 2834364 35 2914364
rect -35 2753396 35 2833396
rect -35 2672428 35 2752428
rect -35 2591460 35 2671460
rect -35 2510492 35 2590492
rect -35 2429524 35 2509524
rect -35 2348556 35 2428556
rect -35 2267588 35 2347588
rect -35 2186620 35 2266620
rect -35 2105652 35 2185652
rect -35 2024684 35 2104684
rect -35 1943716 35 2023716
rect -35 1862748 35 1942748
rect -35 1781780 35 1861780
rect -35 1700812 35 1780812
rect -35 1619844 35 1699844
rect -35 1538876 35 1618876
rect -35 1457908 35 1537908
rect -35 1376940 35 1456940
rect -35 1295972 35 1375972
rect -35 1215004 35 1295004
rect -35 1134036 35 1214036
rect -35 1053068 35 1133068
rect -35 972100 35 1052100
rect -35 891132 35 971132
rect -35 810164 35 890164
rect -35 729196 35 809196
rect -35 648228 35 728228
rect -35 567260 35 647260
rect -35 486292 35 566292
rect -35 405324 35 485324
rect -35 324356 35 404356
rect -35 243388 35 323388
rect -35 162420 35 242420
rect -35 81452 35 161452
rect -35 484 35 80484
rect -35 -80484 35 -484
rect -35 -161452 35 -81452
rect -35 -242420 35 -162420
rect -35 -323388 35 -243388
rect -35 -404356 35 -324356
rect -35 -485324 35 -405324
rect -35 -566292 35 -486292
rect -35 -647260 35 -567260
rect -35 -728228 35 -648228
rect -35 -809196 35 -729196
rect -35 -890164 35 -810164
rect -35 -971132 35 -891132
rect -35 -1052100 35 -972100
rect -35 -1133068 35 -1053068
rect -35 -1214036 35 -1134036
rect -35 -1295004 35 -1215004
rect -35 -1375972 35 -1295972
rect -35 -1456940 35 -1376940
rect -35 -1537908 35 -1457908
rect -35 -1618876 35 -1538876
rect -35 -1699844 35 -1619844
rect -35 -1780812 35 -1700812
rect -35 -1861780 35 -1781780
rect -35 -1942748 35 -1862748
rect -35 -2023716 35 -1943716
rect -35 -2104684 35 -2024684
rect -35 -2185652 35 -2105652
rect -35 -2266620 35 -2186620
rect -35 -2347588 35 -2267588
rect -35 -2428556 35 -2348556
rect -35 -2509524 35 -2429524
rect -35 -2590492 35 -2510492
rect -35 -2671460 35 -2591460
rect -35 -2752428 35 -2672428
rect -35 -2833396 35 -2753396
rect -35 -2914364 35 -2834364
rect -35 -2995332 35 -2915332
rect -35 -3076300 35 -2996300
rect -35 -3157268 35 -3077268
rect -35 -3238236 35 -3158236
rect -35 -3319204 35 -3239204
rect -35 -3400172 35 -3320172
rect -35 -3481140 35 -3401140
rect -35 -3562108 35 -3482108
rect -35 -3643076 35 -3563076
rect -35 -3724044 35 -3644044
rect -35 -3805012 35 -3725012
rect -35 -3885980 35 -3805980
rect -35 -3966948 35 -3886948
rect -35 -4047916 35 -3967916
rect -35 -4128884 35 -4048884
rect -35 -4209852 35 -4129852
rect -35 -4290820 35 -4210820
rect -35 -4371788 35 -4291788
rect -35 -4452756 35 -4372756
rect -35 -4533724 35 -4453724
rect -35 -4614692 35 -4534692
rect -35 -4695660 35 -4615660
rect -35 -4776628 35 -4696628
rect -35 -4857596 35 -4777596
rect -35 -4938564 35 -4858564
rect -35 -5019532 35 -4939532
rect -35 -5100500 35 -5020500
rect -35 -5181468 35 -5101468
rect -35 -5262436 35 -5182436
rect -35 -5343404 35 -5263404
rect -35 -5424372 35 -5344372
rect -35 -5505340 35 -5425340
rect -35 -5586308 35 -5506308
rect -35 -5667276 35 -5587276
rect -35 -5748244 35 -5668244
rect -35 -5829212 35 -5749212
rect -35 -5910180 35 -5830180
rect -35 -5991148 35 -5911148
rect -35 -6072116 35 -5992116
rect -35 -6153084 35 -6073084
rect -35 -6234052 35 -6154052
rect -35 -6315020 35 -6235020
rect -35 -6395988 35 -6315988
rect -35 -6476956 35 -6396956
rect -35 -6557924 35 -6477924
rect -35 -6638892 35 -6558892
rect -35 -6719860 35 -6639860
rect -35 -6800828 35 -6720828
rect -35 -6881796 35 -6801796
rect -35 -6962764 35 -6882764
rect -35 -7043732 35 -6963732
rect -35 -7124700 35 -7044700
rect -35 -7205668 35 -7125668
rect -35 -7286636 35 -7206636
rect -35 -7367604 35 -7287604
rect -35 -7448572 35 -7368572
rect -35 -7529540 35 -7449540
rect -35 -7610508 35 -7530508
rect -35 -7691476 35 -7611476
rect -35 -7772444 35 -7692444
rect -35 -7853412 35 -7773412
rect -35 -7934380 35 -7854380
rect -35 -8015348 35 -7935348
rect -35 -8096316 35 -8016316
rect -35 -8177284 35 -8097284
rect -35 -8258252 35 -8178252
rect -35 -8339220 35 -8259220
rect -35 -8420188 35 -8340188
rect -35 -8501156 35 -8421156
rect -35 -8582124 35 -8502124
rect -35 -8663092 35 -8583092
rect -35 -8744060 35 -8664060
rect -35 -8825028 35 -8745028
rect -35 -8905996 35 -8825996
rect -35 -8986964 35 -8906964
rect -35 -9067932 35 -8987932
rect -35 -9148900 35 -9068900
rect -35 -9229868 35 -9149868
rect -35 -9310836 35 -9230836
rect -35 -9391804 35 -9311804
rect -35 -9472772 35 -9392772
rect -35 -9553740 35 -9473740
rect -35 -9634708 35 -9554708
rect -35 -9715676 35 -9635676
rect -35 -9796644 35 -9716644
rect -35 -9877612 35 -9797612
rect -35 -9958580 35 -9878580
rect -35 -10039548 35 -9959548
rect -35 -10120516 35 -10040516
rect -35 -10201484 35 -10121484
rect -35 -10282452 35 -10202452
rect -35 -10363420 35 -10283420
rect -35 -10444388 35 -10364388
rect -35 -10525356 35 -10445356
rect -35 -10606324 35 -10526324
rect -35 -10687292 35 -10607292
rect -35 -10768260 35 -10688260
rect -35 -10849228 35 -10769228
rect -35 -10930196 35 -10850196
rect -35 -11011164 35 -10931164
rect -35 -11092132 35 -11012132
rect -35 -11173100 35 -11093100
rect -35 -11254068 35 -11174068
rect -35 -11335036 35 -11255036
rect -35 -11416004 35 -11336004
rect -35 -11496972 35 -11416972
rect -35 -11577940 35 -11497940
rect -35 -11658908 35 -11578908
rect -35 -11739876 35 -11659876
rect -35 -11820844 35 -11740844
rect -35 -11901812 35 -11821812
rect -35 -11982780 35 -11902780
rect -35 -12063748 35 -11983748
rect -35 -12144716 35 -12064716
rect -35 -12225684 35 -12145684
rect -35 -12306652 35 -12226652
rect -35 -12387620 35 -12307620
rect -35 -12468588 35 -12388588
rect -35 -12549556 35 -12469556
rect -35 -12630524 35 -12550524
rect -35 -12711492 35 -12631492
rect -35 -12792460 35 -12712460
rect -35 -12873428 35 -12793428
rect -35 -12954396 35 -12874396
rect -35 -13035364 35 -12955364
rect -35 -13116332 35 -13036332
rect -35 -13197300 35 -13117300
rect -35 -13278268 35 -13198268
rect -35 -13359236 35 -13279236
rect -35 -13440204 35 -13360204
rect -35 -13521172 35 -13441172
rect -35 -13602140 35 -13522140
rect -35 -13683108 35 -13603108
rect -35 -13764076 35 -13684076
rect -35 -13845044 35 -13765044
rect -35 -13926012 35 -13846012
rect -35 -14006980 35 -13926980
rect -35 -14087948 35 -14007948
rect -35 -14168916 35 -14088916
rect -35 -14249884 35 -14169884
rect -35 -14330852 35 -14250852
rect -35 -14411820 35 -14331820
rect -35 -14492788 35 -14412788
rect -35 -14573756 35 -14493756
rect -35 -14654724 35 -14574724
rect -35 -14735692 35 -14655692
rect -35 -14816660 35 -14736660
rect -35 -14897628 35 -14817628
rect -35 -14978596 35 -14898596
rect -35 -15059564 35 -14979564
rect -35 -15140532 35 -15060532
rect -35 -15221500 35 -15141500
rect -35 -15302468 35 -15222468
rect -35 -15383436 35 -15303436
rect -35 -15464404 35 -15384404
rect -35 -15545372 35 -15465372
rect -35 -15626340 35 -15546340
rect -35 -15707308 35 -15627308
rect -35 -15788276 35 -15708276
rect -35 -15869244 35 -15789244
rect -35 -15950212 35 -15870212
rect -35 -16031180 35 -15951180
rect -35 -16112148 35 -16032148
rect -35 -16193116 35 -16113116
rect -35 -16274084 35 -16194084
rect -35 -16355052 35 -16275052
rect -35 -16436020 35 -16356020
rect -35 -16516988 35 -16436988
rect -35 -16597956 35 -16517956
rect -35 -16678924 35 -16598924
rect -35 -16759892 35 -16679892
rect -35 -16840860 35 -16760860
rect -35 -16921828 35 -16841828
rect -35 -17002796 35 -16922796
rect -35 -17083764 35 -17003764
rect -35 -17164732 35 -17084732
rect -35 -17245700 35 -17165700
rect -35 -17326668 35 -17246668
rect -35 -17407636 35 -17327636
rect -35 -17488604 35 -17408604
rect -35 -17569572 35 -17489572
rect -35 -17650540 35 -17570540
rect -35 -17731508 35 -17651508
rect -35 -17812476 35 -17732476
rect -35 -17893444 35 -17813444
rect -35 -17974412 35 -17894412
rect -35 -18055380 35 -17975380
rect -35 -18136348 35 -18056348
rect -35 -18217316 35 -18137316
rect -35 -18298284 35 -18218284
rect -35 -18379252 35 -18299252
rect -35 -18460220 35 -18380220
rect -35 -18541188 35 -18461188
rect -35 -18622156 35 -18542156
rect -35 -18703124 35 -18623124
rect -35 -18784092 35 -18704092
rect -35 -18865060 35 -18785060
rect -35 -18946028 35 -18866028
rect -35 -19026996 35 -18946996
rect -35 -19107964 35 -19027964
rect -35 -19188932 35 -19108932
rect -35 -19269900 35 -19189900
rect -35 -19350868 35 -19270868
rect -35 -19431836 35 -19351836
rect -35 -19512804 35 -19432804
rect -35 -19593772 35 -19513772
rect -35 -19674740 35 -19594740
rect -35 -19755708 35 -19675708
rect -35 -19836676 35 -19756676
rect -35 -19917644 35 -19837644
rect -35 -19998612 35 -19918612
rect -35 -20079580 35 -19999580
rect -35 -20160548 35 -20080548
rect -35 -20241516 35 -20161516
<< locali >>
rect -165 20242044 -69 20242078
rect 69 20242044 165 20242078
rect -165 20241982 -131 20242044
rect 131 20241982 165 20242044
rect -165 -20242044 -131 -20241982
rect 131 -20242044 165 -20241982
rect -165 -20242078 -69 -20242044
rect 69 -20242078 165 -20242044
<< viali >>
rect -19 20241533 19 20241930
rect -19 20161102 19 20161499
rect -19 20160565 19 20160962
rect -19 20080134 19 20080531
rect -19 20079597 19 20079994
rect -19 19999166 19 19999563
rect -19 19998629 19 19999026
rect -19 19918198 19 19918595
rect -19 19917661 19 19918058
rect -19 19837230 19 19837627
rect -19 19836693 19 19837090
rect -19 19756262 19 19756659
rect -19 19755725 19 19756122
rect -19 19675294 19 19675691
rect -19 19674757 19 19675154
rect -19 19594326 19 19594723
rect -19 19593789 19 19594186
rect -19 19513358 19 19513755
rect -19 19512821 19 19513218
rect -19 19432390 19 19432787
rect -19 19431853 19 19432250
rect -19 19351422 19 19351819
rect -19 19350885 19 19351282
rect -19 19270454 19 19270851
rect -19 19269917 19 19270314
rect -19 19189486 19 19189883
rect -19 19188949 19 19189346
rect -19 19108518 19 19108915
rect -19 19107981 19 19108378
rect -19 19027550 19 19027947
rect -19 19027013 19 19027410
rect -19 18946582 19 18946979
rect -19 18946045 19 18946442
rect -19 18865614 19 18866011
rect -19 18865077 19 18865474
rect -19 18784646 19 18785043
rect -19 18784109 19 18784506
rect -19 18703678 19 18704075
rect -19 18703141 19 18703538
rect -19 18622710 19 18623107
rect -19 18622173 19 18622570
rect -19 18541742 19 18542139
rect -19 18541205 19 18541602
rect -19 18460774 19 18461171
rect -19 18460237 19 18460634
rect -19 18379806 19 18380203
rect -19 18379269 19 18379666
rect -19 18298838 19 18299235
rect -19 18298301 19 18298698
rect -19 18217870 19 18218267
rect -19 18217333 19 18217730
rect -19 18136902 19 18137299
rect -19 18136365 19 18136762
rect -19 18055934 19 18056331
rect -19 18055397 19 18055794
rect -19 17974966 19 17975363
rect -19 17974429 19 17974826
rect -19 17893998 19 17894395
rect -19 17893461 19 17893858
rect -19 17813030 19 17813427
rect -19 17812493 19 17812890
rect -19 17732062 19 17732459
rect -19 17731525 19 17731922
rect -19 17651094 19 17651491
rect -19 17650557 19 17650954
rect -19 17570126 19 17570523
rect -19 17569589 19 17569986
rect -19 17489158 19 17489555
rect -19 17488621 19 17489018
rect -19 17408190 19 17408587
rect -19 17407653 19 17408050
rect -19 17327222 19 17327619
rect -19 17326685 19 17327082
rect -19 17246254 19 17246651
rect -19 17245717 19 17246114
rect -19 17165286 19 17165683
rect -19 17164749 19 17165146
rect -19 17084318 19 17084715
rect -19 17083781 19 17084178
rect -19 17003350 19 17003747
rect -19 17002813 19 17003210
rect -19 16922382 19 16922779
rect -19 16921845 19 16922242
rect -19 16841414 19 16841811
rect -19 16840877 19 16841274
rect -19 16760446 19 16760843
rect -19 16759909 19 16760306
rect -19 16679478 19 16679875
rect -19 16678941 19 16679338
rect -19 16598510 19 16598907
rect -19 16597973 19 16598370
rect -19 16517542 19 16517939
rect -19 16517005 19 16517402
rect -19 16436574 19 16436971
rect -19 16436037 19 16436434
rect -19 16355606 19 16356003
rect -19 16355069 19 16355466
rect -19 16274638 19 16275035
rect -19 16274101 19 16274498
rect -19 16193670 19 16194067
rect -19 16193133 19 16193530
rect -19 16112702 19 16113099
rect -19 16112165 19 16112562
rect -19 16031734 19 16032131
rect -19 16031197 19 16031594
rect -19 15950766 19 15951163
rect -19 15950229 19 15950626
rect -19 15869798 19 15870195
rect -19 15869261 19 15869658
rect -19 15788830 19 15789227
rect -19 15788293 19 15788690
rect -19 15707862 19 15708259
rect -19 15707325 19 15707722
rect -19 15626894 19 15627291
rect -19 15626357 19 15626754
rect -19 15545926 19 15546323
rect -19 15545389 19 15545786
rect -19 15464958 19 15465355
rect -19 15464421 19 15464818
rect -19 15383990 19 15384387
rect -19 15383453 19 15383850
rect -19 15303022 19 15303419
rect -19 15302485 19 15302882
rect -19 15222054 19 15222451
rect -19 15221517 19 15221914
rect -19 15141086 19 15141483
rect -19 15140549 19 15140946
rect -19 15060118 19 15060515
rect -19 15059581 19 15059978
rect -19 14979150 19 14979547
rect -19 14978613 19 14979010
rect -19 14898182 19 14898579
rect -19 14897645 19 14898042
rect -19 14817214 19 14817611
rect -19 14816677 19 14817074
rect -19 14736246 19 14736643
rect -19 14735709 19 14736106
rect -19 14655278 19 14655675
rect -19 14654741 19 14655138
rect -19 14574310 19 14574707
rect -19 14573773 19 14574170
rect -19 14493342 19 14493739
rect -19 14492805 19 14493202
rect -19 14412374 19 14412771
rect -19 14411837 19 14412234
rect -19 14331406 19 14331803
rect -19 14330869 19 14331266
rect -19 14250438 19 14250835
rect -19 14249901 19 14250298
rect -19 14169470 19 14169867
rect -19 14168933 19 14169330
rect -19 14088502 19 14088899
rect -19 14087965 19 14088362
rect -19 14007534 19 14007931
rect -19 14006997 19 14007394
rect -19 13926566 19 13926963
rect -19 13926029 19 13926426
rect -19 13845598 19 13845995
rect -19 13845061 19 13845458
rect -19 13764630 19 13765027
rect -19 13764093 19 13764490
rect -19 13683662 19 13684059
rect -19 13683125 19 13683522
rect -19 13602694 19 13603091
rect -19 13602157 19 13602554
rect -19 13521726 19 13522123
rect -19 13521189 19 13521586
rect -19 13440758 19 13441155
rect -19 13440221 19 13440618
rect -19 13359790 19 13360187
rect -19 13359253 19 13359650
rect -19 13278822 19 13279219
rect -19 13278285 19 13278682
rect -19 13197854 19 13198251
rect -19 13197317 19 13197714
rect -19 13116886 19 13117283
rect -19 13116349 19 13116746
rect -19 13035918 19 13036315
rect -19 13035381 19 13035778
rect -19 12954950 19 12955347
rect -19 12954413 19 12954810
rect -19 12873982 19 12874379
rect -19 12873445 19 12873842
rect -19 12793014 19 12793411
rect -19 12792477 19 12792874
rect -19 12712046 19 12712443
rect -19 12711509 19 12711906
rect -19 12631078 19 12631475
rect -19 12630541 19 12630938
rect -19 12550110 19 12550507
rect -19 12549573 19 12549970
rect -19 12469142 19 12469539
rect -19 12468605 19 12469002
rect -19 12388174 19 12388571
rect -19 12387637 19 12388034
rect -19 12307206 19 12307603
rect -19 12306669 19 12307066
rect -19 12226238 19 12226635
rect -19 12225701 19 12226098
rect -19 12145270 19 12145667
rect -19 12144733 19 12145130
rect -19 12064302 19 12064699
rect -19 12063765 19 12064162
rect -19 11983334 19 11983731
rect -19 11982797 19 11983194
rect -19 11902366 19 11902763
rect -19 11901829 19 11902226
rect -19 11821398 19 11821795
rect -19 11820861 19 11821258
rect -19 11740430 19 11740827
rect -19 11739893 19 11740290
rect -19 11659462 19 11659859
rect -19 11658925 19 11659322
rect -19 11578494 19 11578891
rect -19 11577957 19 11578354
rect -19 11497526 19 11497923
rect -19 11496989 19 11497386
rect -19 11416558 19 11416955
rect -19 11416021 19 11416418
rect -19 11335590 19 11335987
rect -19 11335053 19 11335450
rect -19 11254622 19 11255019
rect -19 11254085 19 11254482
rect -19 11173654 19 11174051
rect -19 11173117 19 11173514
rect -19 11092686 19 11093083
rect -19 11092149 19 11092546
rect -19 11011718 19 11012115
rect -19 11011181 19 11011578
rect -19 10930750 19 10931147
rect -19 10930213 19 10930610
rect -19 10849782 19 10850179
rect -19 10849245 19 10849642
rect -19 10768814 19 10769211
rect -19 10768277 19 10768674
rect -19 10687846 19 10688243
rect -19 10687309 19 10687706
rect -19 10606878 19 10607275
rect -19 10606341 19 10606738
rect -19 10525910 19 10526307
rect -19 10525373 19 10525770
rect -19 10444942 19 10445339
rect -19 10444405 19 10444802
rect -19 10363974 19 10364371
rect -19 10363437 19 10363834
rect -19 10283006 19 10283403
rect -19 10282469 19 10282866
rect -19 10202038 19 10202435
rect -19 10201501 19 10201898
rect -19 10121070 19 10121467
rect -19 10120533 19 10120930
rect -19 10040102 19 10040499
rect -19 10039565 19 10039962
rect -19 9959134 19 9959531
rect -19 9958597 19 9958994
rect -19 9878166 19 9878563
rect -19 9877629 19 9878026
rect -19 9797198 19 9797595
rect -19 9796661 19 9797058
rect -19 9716230 19 9716627
rect -19 9715693 19 9716090
rect -19 9635262 19 9635659
rect -19 9634725 19 9635122
rect -19 9554294 19 9554691
rect -19 9553757 19 9554154
rect -19 9473326 19 9473723
rect -19 9472789 19 9473186
rect -19 9392358 19 9392755
rect -19 9391821 19 9392218
rect -19 9311390 19 9311787
rect -19 9310853 19 9311250
rect -19 9230422 19 9230819
rect -19 9229885 19 9230282
rect -19 9149454 19 9149851
rect -19 9148917 19 9149314
rect -19 9068486 19 9068883
rect -19 9067949 19 9068346
rect -19 8987518 19 8987915
rect -19 8986981 19 8987378
rect -19 8906550 19 8906947
rect -19 8906013 19 8906410
rect -19 8825582 19 8825979
rect -19 8825045 19 8825442
rect -19 8744614 19 8745011
rect -19 8744077 19 8744474
rect -19 8663646 19 8664043
rect -19 8663109 19 8663506
rect -19 8582678 19 8583075
rect -19 8582141 19 8582538
rect -19 8501710 19 8502107
rect -19 8501173 19 8501570
rect -19 8420742 19 8421139
rect -19 8420205 19 8420602
rect -19 8339774 19 8340171
rect -19 8339237 19 8339634
rect -19 8258806 19 8259203
rect -19 8258269 19 8258666
rect -19 8177838 19 8178235
rect -19 8177301 19 8177698
rect -19 8096870 19 8097267
rect -19 8096333 19 8096730
rect -19 8015902 19 8016299
rect -19 8015365 19 8015762
rect -19 7934934 19 7935331
rect -19 7934397 19 7934794
rect -19 7853966 19 7854363
rect -19 7853429 19 7853826
rect -19 7772998 19 7773395
rect -19 7772461 19 7772858
rect -19 7692030 19 7692427
rect -19 7691493 19 7691890
rect -19 7611062 19 7611459
rect -19 7610525 19 7610922
rect -19 7530094 19 7530491
rect -19 7529557 19 7529954
rect -19 7449126 19 7449523
rect -19 7448589 19 7448986
rect -19 7368158 19 7368555
rect -19 7367621 19 7368018
rect -19 7287190 19 7287587
rect -19 7286653 19 7287050
rect -19 7206222 19 7206619
rect -19 7205685 19 7206082
rect -19 7125254 19 7125651
rect -19 7124717 19 7125114
rect -19 7044286 19 7044683
rect -19 7043749 19 7044146
rect -19 6963318 19 6963715
rect -19 6962781 19 6963178
rect -19 6882350 19 6882747
rect -19 6881813 19 6882210
rect -19 6801382 19 6801779
rect -19 6800845 19 6801242
rect -19 6720414 19 6720811
rect -19 6719877 19 6720274
rect -19 6639446 19 6639843
rect -19 6638909 19 6639306
rect -19 6558478 19 6558875
rect -19 6557941 19 6558338
rect -19 6477510 19 6477907
rect -19 6476973 19 6477370
rect -19 6396542 19 6396939
rect -19 6396005 19 6396402
rect -19 6315574 19 6315971
rect -19 6315037 19 6315434
rect -19 6234606 19 6235003
rect -19 6234069 19 6234466
rect -19 6153638 19 6154035
rect -19 6153101 19 6153498
rect -19 6072670 19 6073067
rect -19 6072133 19 6072530
rect -19 5991702 19 5992099
rect -19 5991165 19 5991562
rect -19 5910734 19 5911131
rect -19 5910197 19 5910594
rect -19 5829766 19 5830163
rect -19 5829229 19 5829626
rect -19 5748798 19 5749195
rect -19 5748261 19 5748658
rect -19 5667830 19 5668227
rect -19 5667293 19 5667690
rect -19 5586862 19 5587259
rect -19 5586325 19 5586722
rect -19 5505894 19 5506291
rect -19 5505357 19 5505754
rect -19 5424926 19 5425323
rect -19 5424389 19 5424786
rect -19 5343958 19 5344355
rect -19 5343421 19 5343818
rect -19 5262990 19 5263387
rect -19 5262453 19 5262850
rect -19 5182022 19 5182419
rect -19 5181485 19 5181882
rect -19 5101054 19 5101451
rect -19 5100517 19 5100914
rect -19 5020086 19 5020483
rect -19 5019549 19 5019946
rect -19 4939118 19 4939515
rect -19 4938581 19 4938978
rect -19 4858150 19 4858547
rect -19 4857613 19 4858010
rect -19 4777182 19 4777579
rect -19 4776645 19 4777042
rect -19 4696214 19 4696611
rect -19 4695677 19 4696074
rect -19 4615246 19 4615643
rect -19 4614709 19 4615106
rect -19 4534278 19 4534675
rect -19 4533741 19 4534138
rect -19 4453310 19 4453707
rect -19 4452773 19 4453170
rect -19 4372342 19 4372739
rect -19 4371805 19 4372202
rect -19 4291374 19 4291771
rect -19 4290837 19 4291234
rect -19 4210406 19 4210803
rect -19 4209869 19 4210266
rect -19 4129438 19 4129835
rect -19 4128901 19 4129298
rect -19 4048470 19 4048867
rect -19 4047933 19 4048330
rect -19 3967502 19 3967899
rect -19 3966965 19 3967362
rect -19 3886534 19 3886931
rect -19 3885997 19 3886394
rect -19 3805566 19 3805963
rect -19 3805029 19 3805426
rect -19 3724598 19 3724995
rect -19 3724061 19 3724458
rect -19 3643630 19 3644027
rect -19 3643093 19 3643490
rect -19 3562662 19 3563059
rect -19 3562125 19 3562522
rect -19 3481694 19 3482091
rect -19 3481157 19 3481554
rect -19 3400726 19 3401123
rect -19 3400189 19 3400586
rect -19 3319758 19 3320155
rect -19 3319221 19 3319618
rect -19 3238790 19 3239187
rect -19 3238253 19 3238650
rect -19 3157822 19 3158219
rect -19 3157285 19 3157682
rect -19 3076854 19 3077251
rect -19 3076317 19 3076714
rect -19 2995886 19 2996283
rect -19 2995349 19 2995746
rect -19 2914918 19 2915315
rect -19 2914381 19 2914778
rect -19 2833950 19 2834347
rect -19 2833413 19 2833810
rect -19 2752982 19 2753379
rect -19 2752445 19 2752842
rect -19 2672014 19 2672411
rect -19 2671477 19 2671874
rect -19 2591046 19 2591443
rect -19 2590509 19 2590906
rect -19 2510078 19 2510475
rect -19 2509541 19 2509938
rect -19 2429110 19 2429507
rect -19 2428573 19 2428970
rect -19 2348142 19 2348539
rect -19 2347605 19 2348002
rect -19 2267174 19 2267571
rect -19 2266637 19 2267034
rect -19 2186206 19 2186603
rect -19 2185669 19 2186066
rect -19 2105238 19 2105635
rect -19 2104701 19 2105098
rect -19 2024270 19 2024667
rect -19 2023733 19 2024130
rect -19 1943302 19 1943699
rect -19 1942765 19 1943162
rect -19 1862334 19 1862731
rect -19 1861797 19 1862194
rect -19 1781366 19 1781763
rect -19 1780829 19 1781226
rect -19 1700398 19 1700795
rect -19 1699861 19 1700258
rect -19 1619430 19 1619827
rect -19 1618893 19 1619290
rect -19 1538462 19 1538859
rect -19 1537925 19 1538322
rect -19 1457494 19 1457891
rect -19 1456957 19 1457354
rect -19 1376526 19 1376923
rect -19 1375989 19 1376386
rect -19 1295558 19 1295955
rect -19 1295021 19 1295418
rect -19 1214590 19 1214987
rect -19 1214053 19 1214450
rect -19 1133622 19 1134019
rect -19 1133085 19 1133482
rect -19 1052654 19 1053051
rect -19 1052117 19 1052514
rect -19 971686 19 972083
rect -19 971149 19 971546
rect -19 890718 19 891115
rect -19 890181 19 890578
rect -19 809750 19 810147
rect -19 809213 19 809610
rect -19 728782 19 729179
rect -19 728245 19 728642
rect -19 647814 19 648211
rect -19 647277 19 647674
rect -19 566846 19 567243
rect -19 566309 19 566706
rect -19 485878 19 486275
rect -19 485341 19 485738
rect -19 404910 19 405307
rect -19 404373 19 404770
rect -19 323942 19 324339
rect -19 323405 19 323802
rect -19 242974 19 243371
rect -19 242437 19 242834
rect -19 162006 19 162403
rect -19 161469 19 161866
rect -19 81038 19 81435
rect -19 80501 19 80898
rect -19 70 19 467
rect -19 -467 19 -70
rect -19 -80898 19 -80501
rect -19 -81435 19 -81038
rect -19 -161866 19 -161469
rect -19 -162403 19 -162006
rect -19 -242834 19 -242437
rect -19 -243371 19 -242974
rect -19 -323802 19 -323405
rect -19 -324339 19 -323942
rect -19 -404770 19 -404373
rect -19 -405307 19 -404910
rect -19 -485738 19 -485341
rect -19 -486275 19 -485878
rect -19 -566706 19 -566309
rect -19 -567243 19 -566846
rect -19 -647674 19 -647277
rect -19 -648211 19 -647814
rect -19 -728642 19 -728245
rect -19 -729179 19 -728782
rect -19 -809610 19 -809213
rect -19 -810147 19 -809750
rect -19 -890578 19 -890181
rect -19 -891115 19 -890718
rect -19 -971546 19 -971149
rect -19 -972083 19 -971686
rect -19 -1052514 19 -1052117
rect -19 -1053051 19 -1052654
rect -19 -1133482 19 -1133085
rect -19 -1134019 19 -1133622
rect -19 -1214450 19 -1214053
rect -19 -1214987 19 -1214590
rect -19 -1295418 19 -1295021
rect -19 -1295955 19 -1295558
rect -19 -1376386 19 -1375989
rect -19 -1376923 19 -1376526
rect -19 -1457354 19 -1456957
rect -19 -1457891 19 -1457494
rect -19 -1538322 19 -1537925
rect -19 -1538859 19 -1538462
rect -19 -1619290 19 -1618893
rect -19 -1619827 19 -1619430
rect -19 -1700258 19 -1699861
rect -19 -1700795 19 -1700398
rect -19 -1781226 19 -1780829
rect -19 -1781763 19 -1781366
rect -19 -1862194 19 -1861797
rect -19 -1862731 19 -1862334
rect -19 -1943162 19 -1942765
rect -19 -1943699 19 -1943302
rect -19 -2024130 19 -2023733
rect -19 -2024667 19 -2024270
rect -19 -2105098 19 -2104701
rect -19 -2105635 19 -2105238
rect -19 -2186066 19 -2185669
rect -19 -2186603 19 -2186206
rect -19 -2267034 19 -2266637
rect -19 -2267571 19 -2267174
rect -19 -2348002 19 -2347605
rect -19 -2348539 19 -2348142
rect -19 -2428970 19 -2428573
rect -19 -2429507 19 -2429110
rect -19 -2509938 19 -2509541
rect -19 -2510475 19 -2510078
rect -19 -2590906 19 -2590509
rect -19 -2591443 19 -2591046
rect -19 -2671874 19 -2671477
rect -19 -2672411 19 -2672014
rect -19 -2752842 19 -2752445
rect -19 -2753379 19 -2752982
rect -19 -2833810 19 -2833413
rect -19 -2834347 19 -2833950
rect -19 -2914778 19 -2914381
rect -19 -2915315 19 -2914918
rect -19 -2995746 19 -2995349
rect -19 -2996283 19 -2995886
rect -19 -3076714 19 -3076317
rect -19 -3077251 19 -3076854
rect -19 -3157682 19 -3157285
rect -19 -3158219 19 -3157822
rect -19 -3238650 19 -3238253
rect -19 -3239187 19 -3238790
rect -19 -3319618 19 -3319221
rect -19 -3320155 19 -3319758
rect -19 -3400586 19 -3400189
rect -19 -3401123 19 -3400726
rect -19 -3481554 19 -3481157
rect -19 -3482091 19 -3481694
rect -19 -3562522 19 -3562125
rect -19 -3563059 19 -3562662
rect -19 -3643490 19 -3643093
rect -19 -3644027 19 -3643630
rect -19 -3724458 19 -3724061
rect -19 -3724995 19 -3724598
rect -19 -3805426 19 -3805029
rect -19 -3805963 19 -3805566
rect -19 -3886394 19 -3885997
rect -19 -3886931 19 -3886534
rect -19 -3967362 19 -3966965
rect -19 -3967899 19 -3967502
rect -19 -4048330 19 -4047933
rect -19 -4048867 19 -4048470
rect -19 -4129298 19 -4128901
rect -19 -4129835 19 -4129438
rect -19 -4210266 19 -4209869
rect -19 -4210803 19 -4210406
rect -19 -4291234 19 -4290837
rect -19 -4291771 19 -4291374
rect -19 -4372202 19 -4371805
rect -19 -4372739 19 -4372342
rect -19 -4453170 19 -4452773
rect -19 -4453707 19 -4453310
rect -19 -4534138 19 -4533741
rect -19 -4534675 19 -4534278
rect -19 -4615106 19 -4614709
rect -19 -4615643 19 -4615246
rect -19 -4696074 19 -4695677
rect -19 -4696611 19 -4696214
rect -19 -4777042 19 -4776645
rect -19 -4777579 19 -4777182
rect -19 -4858010 19 -4857613
rect -19 -4858547 19 -4858150
rect -19 -4938978 19 -4938581
rect -19 -4939515 19 -4939118
rect -19 -5019946 19 -5019549
rect -19 -5020483 19 -5020086
rect -19 -5100914 19 -5100517
rect -19 -5101451 19 -5101054
rect -19 -5181882 19 -5181485
rect -19 -5182419 19 -5182022
rect -19 -5262850 19 -5262453
rect -19 -5263387 19 -5262990
rect -19 -5343818 19 -5343421
rect -19 -5344355 19 -5343958
rect -19 -5424786 19 -5424389
rect -19 -5425323 19 -5424926
rect -19 -5505754 19 -5505357
rect -19 -5506291 19 -5505894
rect -19 -5586722 19 -5586325
rect -19 -5587259 19 -5586862
rect -19 -5667690 19 -5667293
rect -19 -5668227 19 -5667830
rect -19 -5748658 19 -5748261
rect -19 -5749195 19 -5748798
rect -19 -5829626 19 -5829229
rect -19 -5830163 19 -5829766
rect -19 -5910594 19 -5910197
rect -19 -5911131 19 -5910734
rect -19 -5991562 19 -5991165
rect -19 -5992099 19 -5991702
rect -19 -6072530 19 -6072133
rect -19 -6073067 19 -6072670
rect -19 -6153498 19 -6153101
rect -19 -6154035 19 -6153638
rect -19 -6234466 19 -6234069
rect -19 -6235003 19 -6234606
rect -19 -6315434 19 -6315037
rect -19 -6315971 19 -6315574
rect -19 -6396402 19 -6396005
rect -19 -6396939 19 -6396542
rect -19 -6477370 19 -6476973
rect -19 -6477907 19 -6477510
rect -19 -6558338 19 -6557941
rect -19 -6558875 19 -6558478
rect -19 -6639306 19 -6638909
rect -19 -6639843 19 -6639446
rect -19 -6720274 19 -6719877
rect -19 -6720811 19 -6720414
rect -19 -6801242 19 -6800845
rect -19 -6801779 19 -6801382
rect -19 -6882210 19 -6881813
rect -19 -6882747 19 -6882350
rect -19 -6963178 19 -6962781
rect -19 -6963715 19 -6963318
rect -19 -7044146 19 -7043749
rect -19 -7044683 19 -7044286
rect -19 -7125114 19 -7124717
rect -19 -7125651 19 -7125254
rect -19 -7206082 19 -7205685
rect -19 -7206619 19 -7206222
rect -19 -7287050 19 -7286653
rect -19 -7287587 19 -7287190
rect -19 -7368018 19 -7367621
rect -19 -7368555 19 -7368158
rect -19 -7448986 19 -7448589
rect -19 -7449523 19 -7449126
rect -19 -7529954 19 -7529557
rect -19 -7530491 19 -7530094
rect -19 -7610922 19 -7610525
rect -19 -7611459 19 -7611062
rect -19 -7691890 19 -7691493
rect -19 -7692427 19 -7692030
rect -19 -7772858 19 -7772461
rect -19 -7773395 19 -7772998
rect -19 -7853826 19 -7853429
rect -19 -7854363 19 -7853966
rect -19 -7934794 19 -7934397
rect -19 -7935331 19 -7934934
rect -19 -8015762 19 -8015365
rect -19 -8016299 19 -8015902
rect -19 -8096730 19 -8096333
rect -19 -8097267 19 -8096870
rect -19 -8177698 19 -8177301
rect -19 -8178235 19 -8177838
rect -19 -8258666 19 -8258269
rect -19 -8259203 19 -8258806
rect -19 -8339634 19 -8339237
rect -19 -8340171 19 -8339774
rect -19 -8420602 19 -8420205
rect -19 -8421139 19 -8420742
rect -19 -8501570 19 -8501173
rect -19 -8502107 19 -8501710
rect -19 -8582538 19 -8582141
rect -19 -8583075 19 -8582678
rect -19 -8663506 19 -8663109
rect -19 -8664043 19 -8663646
rect -19 -8744474 19 -8744077
rect -19 -8745011 19 -8744614
rect -19 -8825442 19 -8825045
rect -19 -8825979 19 -8825582
rect -19 -8906410 19 -8906013
rect -19 -8906947 19 -8906550
rect -19 -8987378 19 -8986981
rect -19 -8987915 19 -8987518
rect -19 -9068346 19 -9067949
rect -19 -9068883 19 -9068486
rect -19 -9149314 19 -9148917
rect -19 -9149851 19 -9149454
rect -19 -9230282 19 -9229885
rect -19 -9230819 19 -9230422
rect -19 -9311250 19 -9310853
rect -19 -9311787 19 -9311390
rect -19 -9392218 19 -9391821
rect -19 -9392755 19 -9392358
rect -19 -9473186 19 -9472789
rect -19 -9473723 19 -9473326
rect -19 -9554154 19 -9553757
rect -19 -9554691 19 -9554294
rect -19 -9635122 19 -9634725
rect -19 -9635659 19 -9635262
rect -19 -9716090 19 -9715693
rect -19 -9716627 19 -9716230
rect -19 -9797058 19 -9796661
rect -19 -9797595 19 -9797198
rect -19 -9878026 19 -9877629
rect -19 -9878563 19 -9878166
rect -19 -9958994 19 -9958597
rect -19 -9959531 19 -9959134
rect -19 -10039962 19 -10039565
rect -19 -10040499 19 -10040102
rect -19 -10120930 19 -10120533
rect -19 -10121467 19 -10121070
rect -19 -10201898 19 -10201501
rect -19 -10202435 19 -10202038
rect -19 -10282866 19 -10282469
rect -19 -10283403 19 -10283006
rect -19 -10363834 19 -10363437
rect -19 -10364371 19 -10363974
rect -19 -10444802 19 -10444405
rect -19 -10445339 19 -10444942
rect -19 -10525770 19 -10525373
rect -19 -10526307 19 -10525910
rect -19 -10606738 19 -10606341
rect -19 -10607275 19 -10606878
rect -19 -10687706 19 -10687309
rect -19 -10688243 19 -10687846
rect -19 -10768674 19 -10768277
rect -19 -10769211 19 -10768814
rect -19 -10849642 19 -10849245
rect -19 -10850179 19 -10849782
rect -19 -10930610 19 -10930213
rect -19 -10931147 19 -10930750
rect -19 -11011578 19 -11011181
rect -19 -11012115 19 -11011718
rect -19 -11092546 19 -11092149
rect -19 -11093083 19 -11092686
rect -19 -11173514 19 -11173117
rect -19 -11174051 19 -11173654
rect -19 -11254482 19 -11254085
rect -19 -11255019 19 -11254622
rect -19 -11335450 19 -11335053
rect -19 -11335987 19 -11335590
rect -19 -11416418 19 -11416021
rect -19 -11416955 19 -11416558
rect -19 -11497386 19 -11496989
rect -19 -11497923 19 -11497526
rect -19 -11578354 19 -11577957
rect -19 -11578891 19 -11578494
rect -19 -11659322 19 -11658925
rect -19 -11659859 19 -11659462
rect -19 -11740290 19 -11739893
rect -19 -11740827 19 -11740430
rect -19 -11821258 19 -11820861
rect -19 -11821795 19 -11821398
rect -19 -11902226 19 -11901829
rect -19 -11902763 19 -11902366
rect -19 -11983194 19 -11982797
rect -19 -11983731 19 -11983334
rect -19 -12064162 19 -12063765
rect -19 -12064699 19 -12064302
rect -19 -12145130 19 -12144733
rect -19 -12145667 19 -12145270
rect -19 -12226098 19 -12225701
rect -19 -12226635 19 -12226238
rect -19 -12307066 19 -12306669
rect -19 -12307603 19 -12307206
rect -19 -12388034 19 -12387637
rect -19 -12388571 19 -12388174
rect -19 -12469002 19 -12468605
rect -19 -12469539 19 -12469142
rect -19 -12549970 19 -12549573
rect -19 -12550507 19 -12550110
rect -19 -12630938 19 -12630541
rect -19 -12631475 19 -12631078
rect -19 -12711906 19 -12711509
rect -19 -12712443 19 -12712046
rect -19 -12792874 19 -12792477
rect -19 -12793411 19 -12793014
rect -19 -12873842 19 -12873445
rect -19 -12874379 19 -12873982
rect -19 -12954810 19 -12954413
rect -19 -12955347 19 -12954950
rect -19 -13035778 19 -13035381
rect -19 -13036315 19 -13035918
rect -19 -13116746 19 -13116349
rect -19 -13117283 19 -13116886
rect -19 -13197714 19 -13197317
rect -19 -13198251 19 -13197854
rect -19 -13278682 19 -13278285
rect -19 -13279219 19 -13278822
rect -19 -13359650 19 -13359253
rect -19 -13360187 19 -13359790
rect -19 -13440618 19 -13440221
rect -19 -13441155 19 -13440758
rect -19 -13521586 19 -13521189
rect -19 -13522123 19 -13521726
rect -19 -13602554 19 -13602157
rect -19 -13603091 19 -13602694
rect -19 -13683522 19 -13683125
rect -19 -13684059 19 -13683662
rect -19 -13764490 19 -13764093
rect -19 -13765027 19 -13764630
rect -19 -13845458 19 -13845061
rect -19 -13845995 19 -13845598
rect -19 -13926426 19 -13926029
rect -19 -13926963 19 -13926566
rect -19 -14007394 19 -14006997
rect -19 -14007931 19 -14007534
rect -19 -14088362 19 -14087965
rect -19 -14088899 19 -14088502
rect -19 -14169330 19 -14168933
rect -19 -14169867 19 -14169470
rect -19 -14250298 19 -14249901
rect -19 -14250835 19 -14250438
rect -19 -14331266 19 -14330869
rect -19 -14331803 19 -14331406
rect -19 -14412234 19 -14411837
rect -19 -14412771 19 -14412374
rect -19 -14493202 19 -14492805
rect -19 -14493739 19 -14493342
rect -19 -14574170 19 -14573773
rect -19 -14574707 19 -14574310
rect -19 -14655138 19 -14654741
rect -19 -14655675 19 -14655278
rect -19 -14736106 19 -14735709
rect -19 -14736643 19 -14736246
rect -19 -14817074 19 -14816677
rect -19 -14817611 19 -14817214
rect -19 -14898042 19 -14897645
rect -19 -14898579 19 -14898182
rect -19 -14979010 19 -14978613
rect -19 -14979547 19 -14979150
rect -19 -15059978 19 -15059581
rect -19 -15060515 19 -15060118
rect -19 -15140946 19 -15140549
rect -19 -15141483 19 -15141086
rect -19 -15221914 19 -15221517
rect -19 -15222451 19 -15222054
rect -19 -15302882 19 -15302485
rect -19 -15303419 19 -15303022
rect -19 -15383850 19 -15383453
rect -19 -15384387 19 -15383990
rect -19 -15464818 19 -15464421
rect -19 -15465355 19 -15464958
rect -19 -15545786 19 -15545389
rect -19 -15546323 19 -15545926
rect -19 -15626754 19 -15626357
rect -19 -15627291 19 -15626894
rect -19 -15707722 19 -15707325
rect -19 -15708259 19 -15707862
rect -19 -15788690 19 -15788293
rect -19 -15789227 19 -15788830
rect -19 -15869658 19 -15869261
rect -19 -15870195 19 -15869798
rect -19 -15950626 19 -15950229
rect -19 -15951163 19 -15950766
rect -19 -16031594 19 -16031197
rect -19 -16032131 19 -16031734
rect -19 -16112562 19 -16112165
rect -19 -16113099 19 -16112702
rect -19 -16193530 19 -16193133
rect -19 -16194067 19 -16193670
rect -19 -16274498 19 -16274101
rect -19 -16275035 19 -16274638
rect -19 -16355466 19 -16355069
rect -19 -16356003 19 -16355606
rect -19 -16436434 19 -16436037
rect -19 -16436971 19 -16436574
rect -19 -16517402 19 -16517005
rect -19 -16517939 19 -16517542
rect -19 -16598370 19 -16597973
rect -19 -16598907 19 -16598510
rect -19 -16679338 19 -16678941
rect -19 -16679875 19 -16679478
rect -19 -16760306 19 -16759909
rect -19 -16760843 19 -16760446
rect -19 -16841274 19 -16840877
rect -19 -16841811 19 -16841414
rect -19 -16922242 19 -16921845
rect -19 -16922779 19 -16922382
rect -19 -17003210 19 -17002813
rect -19 -17003747 19 -17003350
rect -19 -17084178 19 -17083781
rect -19 -17084715 19 -17084318
rect -19 -17165146 19 -17164749
rect -19 -17165683 19 -17165286
rect -19 -17246114 19 -17245717
rect -19 -17246651 19 -17246254
rect -19 -17327082 19 -17326685
rect -19 -17327619 19 -17327222
rect -19 -17408050 19 -17407653
rect -19 -17408587 19 -17408190
rect -19 -17489018 19 -17488621
rect -19 -17489555 19 -17489158
rect -19 -17569986 19 -17569589
rect -19 -17570523 19 -17570126
rect -19 -17650954 19 -17650557
rect -19 -17651491 19 -17651094
rect -19 -17731922 19 -17731525
rect -19 -17732459 19 -17732062
rect -19 -17812890 19 -17812493
rect -19 -17813427 19 -17813030
rect -19 -17893858 19 -17893461
rect -19 -17894395 19 -17893998
rect -19 -17974826 19 -17974429
rect -19 -17975363 19 -17974966
rect -19 -18055794 19 -18055397
rect -19 -18056331 19 -18055934
rect -19 -18136762 19 -18136365
rect -19 -18137299 19 -18136902
rect -19 -18217730 19 -18217333
rect -19 -18218267 19 -18217870
rect -19 -18298698 19 -18298301
rect -19 -18299235 19 -18298838
rect -19 -18379666 19 -18379269
rect -19 -18380203 19 -18379806
rect -19 -18460634 19 -18460237
rect -19 -18461171 19 -18460774
rect -19 -18541602 19 -18541205
rect -19 -18542139 19 -18541742
rect -19 -18622570 19 -18622173
rect -19 -18623107 19 -18622710
rect -19 -18703538 19 -18703141
rect -19 -18704075 19 -18703678
rect -19 -18784506 19 -18784109
rect -19 -18785043 19 -18784646
rect -19 -18865474 19 -18865077
rect -19 -18866011 19 -18865614
rect -19 -18946442 19 -18946045
rect -19 -18946979 19 -18946582
rect -19 -19027410 19 -19027013
rect -19 -19027947 19 -19027550
rect -19 -19108378 19 -19107981
rect -19 -19108915 19 -19108518
rect -19 -19189346 19 -19188949
rect -19 -19189883 19 -19189486
rect -19 -19270314 19 -19269917
rect -19 -19270851 19 -19270454
rect -19 -19351282 19 -19350885
rect -19 -19351819 19 -19351422
rect -19 -19432250 19 -19431853
rect -19 -19432787 19 -19432390
rect -19 -19513218 19 -19512821
rect -19 -19513755 19 -19513358
rect -19 -19594186 19 -19593789
rect -19 -19594723 19 -19594326
rect -19 -19675154 19 -19674757
rect -19 -19675691 19 -19675294
rect -19 -19756122 19 -19755725
rect -19 -19756659 19 -19756262
rect -19 -19837090 19 -19836693
rect -19 -19837627 19 -19837230
rect -19 -19918058 19 -19917661
rect -19 -19918595 19 -19918198
rect -19 -19999026 19 -19998629
rect -19 -19999563 19 -19999166
rect -19 -20079994 19 -20079597
rect -19 -20080531 19 -20080134
rect -19 -20160962 19 -20160565
rect -19 -20161499 19 -20161102
rect -19 -20241930 19 -20241533
<< metal1 >>
rect -25 20241930 25 20241942
rect -25 20241533 -19 20241930
rect 19 20241533 25 20241930
rect -25 20241521 25 20241533
rect -25 20161499 25 20161511
rect -25 20161102 -19 20161499
rect 19 20161102 25 20161499
rect -25 20161090 25 20161102
rect -25 20160962 25 20160974
rect -25 20160565 -19 20160962
rect 19 20160565 25 20160962
rect -25 20160553 25 20160565
rect -25 20080531 25 20080543
rect -25 20080134 -19 20080531
rect 19 20080134 25 20080531
rect -25 20080122 25 20080134
rect -25 20079994 25 20080006
rect -25 20079597 -19 20079994
rect 19 20079597 25 20079994
rect -25 20079585 25 20079597
rect -25 19999563 25 19999575
rect -25 19999166 -19 19999563
rect 19 19999166 25 19999563
rect -25 19999154 25 19999166
rect -25 19999026 25 19999038
rect -25 19998629 -19 19999026
rect 19 19998629 25 19999026
rect -25 19998617 25 19998629
rect -25 19918595 25 19918607
rect -25 19918198 -19 19918595
rect 19 19918198 25 19918595
rect -25 19918186 25 19918198
rect -25 19918058 25 19918070
rect -25 19917661 -19 19918058
rect 19 19917661 25 19918058
rect -25 19917649 25 19917661
rect -25 19837627 25 19837639
rect -25 19837230 -19 19837627
rect 19 19837230 25 19837627
rect -25 19837218 25 19837230
rect -25 19837090 25 19837102
rect -25 19836693 -19 19837090
rect 19 19836693 25 19837090
rect -25 19836681 25 19836693
rect -25 19756659 25 19756671
rect -25 19756262 -19 19756659
rect 19 19756262 25 19756659
rect -25 19756250 25 19756262
rect -25 19756122 25 19756134
rect -25 19755725 -19 19756122
rect 19 19755725 25 19756122
rect -25 19755713 25 19755725
rect -25 19675691 25 19675703
rect -25 19675294 -19 19675691
rect 19 19675294 25 19675691
rect -25 19675282 25 19675294
rect -25 19675154 25 19675166
rect -25 19674757 -19 19675154
rect 19 19674757 25 19675154
rect -25 19674745 25 19674757
rect -25 19594723 25 19594735
rect -25 19594326 -19 19594723
rect 19 19594326 25 19594723
rect -25 19594314 25 19594326
rect -25 19594186 25 19594198
rect -25 19593789 -19 19594186
rect 19 19593789 25 19594186
rect -25 19593777 25 19593789
rect -25 19513755 25 19513767
rect -25 19513358 -19 19513755
rect 19 19513358 25 19513755
rect -25 19513346 25 19513358
rect -25 19513218 25 19513230
rect -25 19512821 -19 19513218
rect 19 19512821 25 19513218
rect -25 19512809 25 19512821
rect -25 19432787 25 19432799
rect -25 19432390 -19 19432787
rect 19 19432390 25 19432787
rect -25 19432378 25 19432390
rect -25 19432250 25 19432262
rect -25 19431853 -19 19432250
rect 19 19431853 25 19432250
rect -25 19431841 25 19431853
rect -25 19351819 25 19351831
rect -25 19351422 -19 19351819
rect 19 19351422 25 19351819
rect -25 19351410 25 19351422
rect -25 19351282 25 19351294
rect -25 19350885 -19 19351282
rect 19 19350885 25 19351282
rect -25 19350873 25 19350885
rect -25 19270851 25 19270863
rect -25 19270454 -19 19270851
rect 19 19270454 25 19270851
rect -25 19270442 25 19270454
rect -25 19270314 25 19270326
rect -25 19269917 -19 19270314
rect 19 19269917 25 19270314
rect -25 19269905 25 19269917
rect -25 19189883 25 19189895
rect -25 19189486 -19 19189883
rect 19 19189486 25 19189883
rect -25 19189474 25 19189486
rect -25 19189346 25 19189358
rect -25 19188949 -19 19189346
rect 19 19188949 25 19189346
rect -25 19188937 25 19188949
rect -25 19108915 25 19108927
rect -25 19108518 -19 19108915
rect 19 19108518 25 19108915
rect -25 19108506 25 19108518
rect -25 19108378 25 19108390
rect -25 19107981 -19 19108378
rect 19 19107981 25 19108378
rect -25 19107969 25 19107981
rect -25 19027947 25 19027959
rect -25 19027550 -19 19027947
rect 19 19027550 25 19027947
rect -25 19027538 25 19027550
rect -25 19027410 25 19027422
rect -25 19027013 -19 19027410
rect 19 19027013 25 19027410
rect -25 19027001 25 19027013
rect -25 18946979 25 18946991
rect -25 18946582 -19 18946979
rect 19 18946582 25 18946979
rect -25 18946570 25 18946582
rect -25 18946442 25 18946454
rect -25 18946045 -19 18946442
rect 19 18946045 25 18946442
rect -25 18946033 25 18946045
rect -25 18866011 25 18866023
rect -25 18865614 -19 18866011
rect 19 18865614 25 18866011
rect -25 18865602 25 18865614
rect -25 18865474 25 18865486
rect -25 18865077 -19 18865474
rect 19 18865077 25 18865474
rect -25 18865065 25 18865077
rect -25 18785043 25 18785055
rect -25 18784646 -19 18785043
rect 19 18784646 25 18785043
rect -25 18784634 25 18784646
rect -25 18784506 25 18784518
rect -25 18784109 -19 18784506
rect 19 18784109 25 18784506
rect -25 18784097 25 18784109
rect -25 18704075 25 18704087
rect -25 18703678 -19 18704075
rect 19 18703678 25 18704075
rect -25 18703666 25 18703678
rect -25 18703538 25 18703550
rect -25 18703141 -19 18703538
rect 19 18703141 25 18703538
rect -25 18703129 25 18703141
rect -25 18623107 25 18623119
rect -25 18622710 -19 18623107
rect 19 18622710 25 18623107
rect -25 18622698 25 18622710
rect -25 18622570 25 18622582
rect -25 18622173 -19 18622570
rect 19 18622173 25 18622570
rect -25 18622161 25 18622173
rect -25 18542139 25 18542151
rect -25 18541742 -19 18542139
rect 19 18541742 25 18542139
rect -25 18541730 25 18541742
rect -25 18541602 25 18541614
rect -25 18541205 -19 18541602
rect 19 18541205 25 18541602
rect -25 18541193 25 18541205
rect -25 18461171 25 18461183
rect -25 18460774 -19 18461171
rect 19 18460774 25 18461171
rect -25 18460762 25 18460774
rect -25 18460634 25 18460646
rect -25 18460237 -19 18460634
rect 19 18460237 25 18460634
rect -25 18460225 25 18460237
rect -25 18380203 25 18380215
rect -25 18379806 -19 18380203
rect 19 18379806 25 18380203
rect -25 18379794 25 18379806
rect -25 18379666 25 18379678
rect -25 18379269 -19 18379666
rect 19 18379269 25 18379666
rect -25 18379257 25 18379269
rect -25 18299235 25 18299247
rect -25 18298838 -19 18299235
rect 19 18298838 25 18299235
rect -25 18298826 25 18298838
rect -25 18298698 25 18298710
rect -25 18298301 -19 18298698
rect 19 18298301 25 18298698
rect -25 18298289 25 18298301
rect -25 18218267 25 18218279
rect -25 18217870 -19 18218267
rect 19 18217870 25 18218267
rect -25 18217858 25 18217870
rect -25 18217730 25 18217742
rect -25 18217333 -19 18217730
rect 19 18217333 25 18217730
rect -25 18217321 25 18217333
rect -25 18137299 25 18137311
rect -25 18136902 -19 18137299
rect 19 18136902 25 18137299
rect -25 18136890 25 18136902
rect -25 18136762 25 18136774
rect -25 18136365 -19 18136762
rect 19 18136365 25 18136762
rect -25 18136353 25 18136365
rect -25 18056331 25 18056343
rect -25 18055934 -19 18056331
rect 19 18055934 25 18056331
rect -25 18055922 25 18055934
rect -25 18055794 25 18055806
rect -25 18055397 -19 18055794
rect 19 18055397 25 18055794
rect -25 18055385 25 18055397
rect -25 17975363 25 17975375
rect -25 17974966 -19 17975363
rect 19 17974966 25 17975363
rect -25 17974954 25 17974966
rect -25 17974826 25 17974838
rect -25 17974429 -19 17974826
rect 19 17974429 25 17974826
rect -25 17974417 25 17974429
rect -25 17894395 25 17894407
rect -25 17893998 -19 17894395
rect 19 17893998 25 17894395
rect -25 17893986 25 17893998
rect -25 17893858 25 17893870
rect -25 17893461 -19 17893858
rect 19 17893461 25 17893858
rect -25 17893449 25 17893461
rect -25 17813427 25 17813439
rect -25 17813030 -19 17813427
rect 19 17813030 25 17813427
rect -25 17813018 25 17813030
rect -25 17812890 25 17812902
rect -25 17812493 -19 17812890
rect 19 17812493 25 17812890
rect -25 17812481 25 17812493
rect -25 17732459 25 17732471
rect -25 17732062 -19 17732459
rect 19 17732062 25 17732459
rect -25 17732050 25 17732062
rect -25 17731922 25 17731934
rect -25 17731525 -19 17731922
rect 19 17731525 25 17731922
rect -25 17731513 25 17731525
rect -25 17651491 25 17651503
rect -25 17651094 -19 17651491
rect 19 17651094 25 17651491
rect -25 17651082 25 17651094
rect -25 17650954 25 17650966
rect -25 17650557 -19 17650954
rect 19 17650557 25 17650954
rect -25 17650545 25 17650557
rect -25 17570523 25 17570535
rect -25 17570126 -19 17570523
rect 19 17570126 25 17570523
rect -25 17570114 25 17570126
rect -25 17569986 25 17569998
rect -25 17569589 -19 17569986
rect 19 17569589 25 17569986
rect -25 17569577 25 17569589
rect -25 17489555 25 17489567
rect -25 17489158 -19 17489555
rect 19 17489158 25 17489555
rect -25 17489146 25 17489158
rect -25 17489018 25 17489030
rect -25 17488621 -19 17489018
rect 19 17488621 25 17489018
rect -25 17488609 25 17488621
rect -25 17408587 25 17408599
rect -25 17408190 -19 17408587
rect 19 17408190 25 17408587
rect -25 17408178 25 17408190
rect -25 17408050 25 17408062
rect -25 17407653 -19 17408050
rect 19 17407653 25 17408050
rect -25 17407641 25 17407653
rect -25 17327619 25 17327631
rect -25 17327222 -19 17327619
rect 19 17327222 25 17327619
rect -25 17327210 25 17327222
rect -25 17327082 25 17327094
rect -25 17326685 -19 17327082
rect 19 17326685 25 17327082
rect -25 17326673 25 17326685
rect -25 17246651 25 17246663
rect -25 17246254 -19 17246651
rect 19 17246254 25 17246651
rect -25 17246242 25 17246254
rect -25 17246114 25 17246126
rect -25 17245717 -19 17246114
rect 19 17245717 25 17246114
rect -25 17245705 25 17245717
rect -25 17165683 25 17165695
rect -25 17165286 -19 17165683
rect 19 17165286 25 17165683
rect -25 17165274 25 17165286
rect -25 17165146 25 17165158
rect -25 17164749 -19 17165146
rect 19 17164749 25 17165146
rect -25 17164737 25 17164749
rect -25 17084715 25 17084727
rect -25 17084318 -19 17084715
rect 19 17084318 25 17084715
rect -25 17084306 25 17084318
rect -25 17084178 25 17084190
rect -25 17083781 -19 17084178
rect 19 17083781 25 17084178
rect -25 17083769 25 17083781
rect -25 17003747 25 17003759
rect -25 17003350 -19 17003747
rect 19 17003350 25 17003747
rect -25 17003338 25 17003350
rect -25 17003210 25 17003222
rect -25 17002813 -19 17003210
rect 19 17002813 25 17003210
rect -25 17002801 25 17002813
rect -25 16922779 25 16922791
rect -25 16922382 -19 16922779
rect 19 16922382 25 16922779
rect -25 16922370 25 16922382
rect -25 16922242 25 16922254
rect -25 16921845 -19 16922242
rect 19 16921845 25 16922242
rect -25 16921833 25 16921845
rect -25 16841811 25 16841823
rect -25 16841414 -19 16841811
rect 19 16841414 25 16841811
rect -25 16841402 25 16841414
rect -25 16841274 25 16841286
rect -25 16840877 -19 16841274
rect 19 16840877 25 16841274
rect -25 16840865 25 16840877
rect -25 16760843 25 16760855
rect -25 16760446 -19 16760843
rect 19 16760446 25 16760843
rect -25 16760434 25 16760446
rect -25 16760306 25 16760318
rect -25 16759909 -19 16760306
rect 19 16759909 25 16760306
rect -25 16759897 25 16759909
rect -25 16679875 25 16679887
rect -25 16679478 -19 16679875
rect 19 16679478 25 16679875
rect -25 16679466 25 16679478
rect -25 16679338 25 16679350
rect -25 16678941 -19 16679338
rect 19 16678941 25 16679338
rect -25 16678929 25 16678941
rect -25 16598907 25 16598919
rect -25 16598510 -19 16598907
rect 19 16598510 25 16598907
rect -25 16598498 25 16598510
rect -25 16598370 25 16598382
rect -25 16597973 -19 16598370
rect 19 16597973 25 16598370
rect -25 16597961 25 16597973
rect -25 16517939 25 16517951
rect -25 16517542 -19 16517939
rect 19 16517542 25 16517939
rect -25 16517530 25 16517542
rect -25 16517402 25 16517414
rect -25 16517005 -19 16517402
rect 19 16517005 25 16517402
rect -25 16516993 25 16517005
rect -25 16436971 25 16436983
rect -25 16436574 -19 16436971
rect 19 16436574 25 16436971
rect -25 16436562 25 16436574
rect -25 16436434 25 16436446
rect -25 16436037 -19 16436434
rect 19 16436037 25 16436434
rect -25 16436025 25 16436037
rect -25 16356003 25 16356015
rect -25 16355606 -19 16356003
rect 19 16355606 25 16356003
rect -25 16355594 25 16355606
rect -25 16355466 25 16355478
rect -25 16355069 -19 16355466
rect 19 16355069 25 16355466
rect -25 16355057 25 16355069
rect -25 16275035 25 16275047
rect -25 16274638 -19 16275035
rect 19 16274638 25 16275035
rect -25 16274626 25 16274638
rect -25 16274498 25 16274510
rect -25 16274101 -19 16274498
rect 19 16274101 25 16274498
rect -25 16274089 25 16274101
rect -25 16194067 25 16194079
rect -25 16193670 -19 16194067
rect 19 16193670 25 16194067
rect -25 16193658 25 16193670
rect -25 16193530 25 16193542
rect -25 16193133 -19 16193530
rect 19 16193133 25 16193530
rect -25 16193121 25 16193133
rect -25 16113099 25 16113111
rect -25 16112702 -19 16113099
rect 19 16112702 25 16113099
rect -25 16112690 25 16112702
rect -25 16112562 25 16112574
rect -25 16112165 -19 16112562
rect 19 16112165 25 16112562
rect -25 16112153 25 16112165
rect -25 16032131 25 16032143
rect -25 16031734 -19 16032131
rect 19 16031734 25 16032131
rect -25 16031722 25 16031734
rect -25 16031594 25 16031606
rect -25 16031197 -19 16031594
rect 19 16031197 25 16031594
rect -25 16031185 25 16031197
rect -25 15951163 25 15951175
rect -25 15950766 -19 15951163
rect 19 15950766 25 15951163
rect -25 15950754 25 15950766
rect -25 15950626 25 15950638
rect -25 15950229 -19 15950626
rect 19 15950229 25 15950626
rect -25 15950217 25 15950229
rect -25 15870195 25 15870207
rect -25 15869798 -19 15870195
rect 19 15869798 25 15870195
rect -25 15869786 25 15869798
rect -25 15869658 25 15869670
rect -25 15869261 -19 15869658
rect 19 15869261 25 15869658
rect -25 15869249 25 15869261
rect -25 15789227 25 15789239
rect -25 15788830 -19 15789227
rect 19 15788830 25 15789227
rect -25 15788818 25 15788830
rect -25 15788690 25 15788702
rect -25 15788293 -19 15788690
rect 19 15788293 25 15788690
rect -25 15788281 25 15788293
rect -25 15708259 25 15708271
rect -25 15707862 -19 15708259
rect 19 15707862 25 15708259
rect -25 15707850 25 15707862
rect -25 15707722 25 15707734
rect -25 15707325 -19 15707722
rect 19 15707325 25 15707722
rect -25 15707313 25 15707325
rect -25 15627291 25 15627303
rect -25 15626894 -19 15627291
rect 19 15626894 25 15627291
rect -25 15626882 25 15626894
rect -25 15626754 25 15626766
rect -25 15626357 -19 15626754
rect 19 15626357 25 15626754
rect -25 15626345 25 15626357
rect -25 15546323 25 15546335
rect -25 15545926 -19 15546323
rect 19 15545926 25 15546323
rect -25 15545914 25 15545926
rect -25 15545786 25 15545798
rect -25 15545389 -19 15545786
rect 19 15545389 25 15545786
rect -25 15545377 25 15545389
rect -25 15465355 25 15465367
rect -25 15464958 -19 15465355
rect 19 15464958 25 15465355
rect -25 15464946 25 15464958
rect -25 15464818 25 15464830
rect -25 15464421 -19 15464818
rect 19 15464421 25 15464818
rect -25 15464409 25 15464421
rect -25 15384387 25 15384399
rect -25 15383990 -19 15384387
rect 19 15383990 25 15384387
rect -25 15383978 25 15383990
rect -25 15383850 25 15383862
rect -25 15383453 -19 15383850
rect 19 15383453 25 15383850
rect -25 15383441 25 15383453
rect -25 15303419 25 15303431
rect -25 15303022 -19 15303419
rect 19 15303022 25 15303419
rect -25 15303010 25 15303022
rect -25 15302882 25 15302894
rect -25 15302485 -19 15302882
rect 19 15302485 25 15302882
rect -25 15302473 25 15302485
rect -25 15222451 25 15222463
rect -25 15222054 -19 15222451
rect 19 15222054 25 15222451
rect -25 15222042 25 15222054
rect -25 15221914 25 15221926
rect -25 15221517 -19 15221914
rect 19 15221517 25 15221914
rect -25 15221505 25 15221517
rect -25 15141483 25 15141495
rect -25 15141086 -19 15141483
rect 19 15141086 25 15141483
rect -25 15141074 25 15141086
rect -25 15140946 25 15140958
rect -25 15140549 -19 15140946
rect 19 15140549 25 15140946
rect -25 15140537 25 15140549
rect -25 15060515 25 15060527
rect -25 15060118 -19 15060515
rect 19 15060118 25 15060515
rect -25 15060106 25 15060118
rect -25 15059978 25 15059990
rect -25 15059581 -19 15059978
rect 19 15059581 25 15059978
rect -25 15059569 25 15059581
rect -25 14979547 25 14979559
rect -25 14979150 -19 14979547
rect 19 14979150 25 14979547
rect -25 14979138 25 14979150
rect -25 14979010 25 14979022
rect -25 14978613 -19 14979010
rect 19 14978613 25 14979010
rect -25 14978601 25 14978613
rect -25 14898579 25 14898591
rect -25 14898182 -19 14898579
rect 19 14898182 25 14898579
rect -25 14898170 25 14898182
rect -25 14898042 25 14898054
rect -25 14897645 -19 14898042
rect 19 14897645 25 14898042
rect -25 14897633 25 14897645
rect -25 14817611 25 14817623
rect -25 14817214 -19 14817611
rect 19 14817214 25 14817611
rect -25 14817202 25 14817214
rect -25 14817074 25 14817086
rect -25 14816677 -19 14817074
rect 19 14816677 25 14817074
rect -25 14816665 25 14816677
rect -25 14736643 25 14736655
rect -25 14736246 -19 14736643
rect 19 14736246 25 14736643
rect -25 14736234 25 14736246
rect -25 14736106 25 14736118
rect -25 14735709 -19 14736106
rect 19 14735709 25 14736106
rect -25 14735697 25 14735709
rect -25 14655675 25 14655687
rect -25 14655278 -19 14655675
rect 19 14655278 25 14655675
rect -25 14655266 25 14655278
rect -25 14655138 25 14655150
rect -25 14654741 -19 14655138
rect 19 14654741 25 14655138
rect -25 14654729 25 14654741
rect -25 14574707 25 14574719
rect -25 14574310 -19 14574707
rect 19 14574310 25 14574707
rect -25 14574298 25 14574310
rect -25 14574170 25 14574182
rect -25 14573773 -19 14574170
rect 19 14573773 25 14574170
rect -25 14573761 25 14573773
rect -25 14493739 25 14493751
rect -25 14493342 -19 14493739
rect 19 14493342 25 14493739
rect -25 14493330 25 14493342
rect -25 14493202 25 14493214
rect -25 14492805 -19 14493202
rect 19 14492805 25 14493202
rect -25 14492793 25 14492805
rect -25 14412771 25 14412783
rect -25 14412374 -19 14412771
rect 19 14412374 25 14412771
rect -25 14412362 25 14412374
rect -25 14412234 25 14412246
rect -25 14411837 -19 14412234
rect 19 14411837 25 14412234
rect -25 14411825 25 14411837
rect -25 14331803 25 14331815
rect -25 14331406 -19 14331803
rect 19 14331406 25 14331803
rect -25 14331394 25 14331406
rect -25 14331266 25 14331278
rect -25 14330869 -19 14331266
rect 19 14330869 25 14331266
rect -25 14330857 25 14330869
rect -25 14250835 25 14250847
rect -25 14250438 -19 14250835
rect 19 14250438 25 14250835
rect -25 14250426 25 14250438
rect -25 14250298 25 14250310
rect -25 14249901 -19 14250298
rect 19 14249901 25 14250298
rect -25 14249889 25 14249901
rect -25 14169867 25 14169879
rect -25 14169470 -19 14169867
rect 19 14169470 25 14169867
rect -25 14169458 25 14169470
rect -25 14169330 25 14169342
rect -25 14168933 -19 14169330
rect 19 14168933 25 14169330
rect -25 14168921 25 14168933
rect -25 14088899 25 14088911
rect -25 14088502 -19 14088899
rect 19 14088502 25 14088899
rect -25 14088490 25 14088502
rect -25 14088362 25 14088374
rect -25 14087965 -19 14088362
rect 19 14087965 25 14088362
rect -25 14087953 25 14087965
rect -25 14007931 25 14007943
rect -25 14007534 -19 14007931
rect 19 14007534 25 14007931
rect -25 14007522 25 14007534
rect -25 14007394 25 14007406
rect -25 14006997 -19 14007394
rect 19 14006997 25 14007394
rect -25 14006985 25 14006997
rect -25 13926963 25 13926975
rect -25 13926566 -19 13926963
rect 19 13926566 25 13926963
rect -25 13926554 25 13926566
rect -25 13926426 25 13926438
rect -25 13926029 -19 13926426
rect 19 13926029 25 13926426
rect -25 13926017 25 13926029
rect -25 13845995 25 13846007
rect -25 13845598 -19 13845995
rect 19 13845598 25 13845995
rect -25 13845586 25 13845598
rect -25 13845458 25 13845470
rect -25 13845061 -19 13845458
rect 19 13845061 25 13845458
rect -25 13845049 25 13845061
rect -25 13765027 25 13765039
rect -25 13764630 -19 13765027
rect 19 13764630 25 13765027
rect -25 13764618 25 13764630
rect -25 13764490 25 13764502
rect -25 13764093 -19 13764490
rect 19 13764093 25 13764490
rect -25 13764081 25 13764093
rect -25 13684059 25 13684071
rect -25 13683662 -19 13684059
rect 19 13683662 25 13684059
rect -25 13683650 25 13683662
rect -25 13683522 25 13683534
rect -25 13683125 -19 13683522
rect 19 13683125 25 13683522
rect -25 13683113 25 13683125
rect -25 13603091 25 13603103
rect -25 13602694 -19 13603091
rect 19 13602694 25 13603091
rect -25 13602682 25 13602694
rect -25 13602554 25 13602566
rect -25 13602157 -19 13602554
rect 19 13602157 25 13602554
rect -25 13602145 25 13602157
rect -25 13522123 25 13522135
rect -25 13521726 -19 13522123
rect 19 13521726 25 13522123
rect -25 13521714 25 13521726
rect -25 13521586 25 13521598
rect -25 13521189 -19 13521586
rect 19 13521189 25 13521586
rect -25 13521177 25 13521189
rect -25 13441155 25 13441167
rect -25 13440758 -19 13441155
rect 19 13440758 25 13441155
rect -25 13440746 25 13440758
rect -25 13440618 25 13440630
rect -25 13440221 -19 13440618
rect 19 13440221 25 13440618
rect -25 13440209 25 13440221
rect -25 13360187 25 13360199
rect -25 13359790 -19 13360187
rect 19 13359790 25 13360187
rect -25 13359778 25 13359790
rect -25 13359650 25 13359662
rect -25 13359253 -19 13359650
rect 19 13359253 25 13359650
rect -25 13359241 25 13359253
rect -25 13279219 25 13279231
rect -25 13278822 -19 13279219
rect 19 13278822 25 13279219
rect -25 13278810 25 13278822
rect -25 13278682 25 13278694
rect -25 13278285 -19 13278682
rect 19 13278285 25 13278682
rect -25 13278273 25 13278285
rect -25 13198251 25 13198263
rect -25 13197854 -19 13198251
rect 19 13197854 25 13198251
rect -25 13197842 25 13197854
rect -25 13197714 25 13197726
rect -25 13197317 -19 13197714
rect 19 13197317 25 13197714
rect -25 13197305 25 13197317
rect -25 13117283 25 13117295
rect -25 13116886 -19 13117283
rect 19 13116886 25 13117283
rect -25 13116874 25 13116886
rect -25 13116746 25 13116758
rect -25 13116349 -19 13116746
rect 19 13116349 25 13116746
rect -25 13116337 25 13116349
rect -25 13036315 25 13036327
rect -25 13035918 -19 13036315
rect 19 13035918 25 13036315
rect -25 13035906 25 13035918
rect -25 13035778 25 13035790
rect -25 13035381 -19 13035778
rect 19 13035381 25 13035778
rect -25 13035369 25 13035381
rect -25 12955347 25 12955359
rect -25 12954950 -19 12955347
rect 19 12954950 25 12955347
rect -25 12954938 25 12954950
rect -25 12954810 25 12954822
rect -25 12954413 -19 12954810
rect 19 12954413 25 12954810
rect -25 12954401 25 12954413
rect -25 12874379 25 12874391
rect -25 12873982 -19 12874379
rect 19 12873982 25 12874379
rect -25 12873970 25 12873982
rect -25 12873842 25 12873854
rect -25 12873445 -19 12873842
rect 19 12873445 25 12873842
rect -25 12873433 25 12873445
rect -25 12793411 25 12793423
rect -25 12793014 -19 12793411
rect 19 12793014 25 12793411
rect -25 12793002 25 12793014
rect -25 12792874 25 12792886
rect -25 12792477 -19 12792874
rect 19 12792477 25 12792874
rect -25 12792465 25 12792477
rect -25 12712443 25 12712455
rect -25 12712046 -19 12712443
rect 19 12712046 25 12712443
rect -25 12712034 25 12712046
rect -25 12711906 25 12711918
rect -25 12711509 -19 12711906
rect 19 12711509 25 12711906
rect -25 12711497 25 12711509
rect -25 12631475 25 12631487
rect -25 12631078 -19 12631475
rect 19 12631078 25 12631475
rect -25 12631066 25 12631078
rect -25 12630938 25 12630950
rect -25 12630541 -19 12630938
rect 19 12630541 25 12630938
rect -25 12630529 25 12630541
rect -25 12550507 25 12550519
rect -25 12550110 -19 12550507
rect 19 12550110 25 12550507
rect -25 12550098 25 12550110
rect -25 12549970 25 12549982
rect -25 12549573 -19 12549970
rect 19 12549573 25 12549970
rect -25 12549561 25 12549573
rect -25 12469539 25 12469551
rect -25 12469142 -19 12469539
rect 19 12469142 25 12469539
rect -25 12469130 25 12469142
rect -25 12469002 25 12469014
rect -25 12468605 -19 12469002
rect 19 12468605 25 12469002
rect -25 12468593 25 12468605
rect -25 12388571 25 12388583
rect -25 12388174 -19 12388571
rect 19 12388174 25 12388571
rect -25 12388162 25 12388174
rect -25 12388034 25 12388046
rect -25 12387637 -19 12388034
rect 19 12387637 25 12388034
rect -25 12387625 25 12387637
rect -25 12307603 25 12307615
rect -25 12307206 -19 12307603
rect 19 12307206 25 12307603
rect -25 12307194 25 12307206
rect -25 12307066 25 12307078
rect -25 12306669 -19 12307066
rect 19 12306669 25 12307066
rect -25 12306657 25 12306669
rect -25 12226635 25 12226647
rect -25 12226238 -19 12226635
rect 19 12226238 25 12226635
rect -25 12226226 25 12226238
rect -25 12226098 25 12226110
rect -25 12225701 -19 12226098
rect 19 12225701 25 12226098
rect -25 12225689 25 12225701
rect -25 12145667 25 12145679
rect -25 12145270 -19 12145667
rect 19 12145270 25 12145667
rect -25 12145258 25 12145270
rect -25 12145130 25 12145142
rect -25 12144733 -19 12145130
rect 19 12144733 25 12145130
rect -25 12144721 25 12144733
rect -25 12064699 25 12064711
rect -25 12064302 -19 12064699
rect 19 12064302 25 12064699
rect -25 12064290 25 12064302
rect -25 12064162 25 12064174
rect -25 12063765 -19 12064162
rect 19 12063765 25 12064162
rect -25 12063753 25 12063765
rect -25 11983731 25 11983743
rect -25 11983334 -19 11983731
rect 19 11983334 25 11983731
rect -25 11983322 25 11983334
rect -25 11983194 25 11983206
rect -25 11982797 -19 11983194
rect 19 11982797 25 11983194
rect -25 11982785 25 11982797
rect -25 11902763 25 11902775
rect -25 11902366 -19 11902763
rect 19 11902366 25 11902763
rect -25 11902354 25 11902366
rect -25 11902226 25 11902238
rect -25 11901829 -19 11902226
rect 19 11901829 25 11902226
rect -25 11901817 25 11901829
rect -25 11821795 25 11821807
rect -25 11821398 -19 11821795
rect 19 11821398 25 11821795
rect -25 11821386 25 11821398
rect -25 11821258 25 11821270
rect -25 11820861 -19 11821258
rect 19 11820861 25 11821258
rect -25 11820849 25 11820861
rect -25 11740827 25 11740839
rect -25 11740430 -19 11740827
rect 19 11740430 25 11740827
rect -25 11740418 25 11740430
rect -25 11740290 25 11740302
rect -25 11739893 -19 11740290
rect 19 11739893 25 11740290
rect -25 11739881 25 11739893
rect -25 11659859 25 11659871
rect -25 11659462 -19 11659859
rect 19 11659462 25 11659859
rect -25 11659450 25 11659462
rect -25 11659322 25 11659334
rect -25 11658925 -19 11659322
rect 19 11658925 25 11659322
rect -25 11658913 25 11658925
rect -25 11578891 25 11578903
rect -25 11578494 -19 11578891
rect 19 11578494 25 11578891
rect -25 11578482 25 11578494
rect -25 11578354 25 11578366
rect -25 11577957 -19 11578354
rect 19 11577957 25 11578354
rect -25 11577945 25 11577957
rect -25 11497923 25 11497935
rect -25 11497526 -19 11497923
rect 19 11497526 25 11497923
rect -25 11497514 25 11497526
rect -25 11497386 25 11497398
rect -25 11496989 -19 11497386
rect 19 11496989 25 11497386
rect -25 11496977 25 11496989
rect -25 11416955 25 11416967
rect -25 11416558 -19 11416955
rect 19 11416558 25 11416955
rect -25 11416546 25 11416558
rect -25 11416418 25 11416430
rect -25 11416021 -19 11416418
rect 19 11416021 25 11416418
rect -25 11416009 25 11416021
rect -25 11335987 25 11335999
rect -25 11335590 -19 11335987
rect 19 11335590 25 11335987
rect -25 11335578 25 11335590
rect -25 11335450 25 11335462
rect -25 11335053 -19 11335450
rect 19 11335053 25 11335450
rect -25 11335041 25 11335053
rect -25 11255019 25 11255031
rect -25 11254622 -19 11255019
rect 19 11254622 25 11255019
rect -25 11254610 25 11254622
rect -25 11254482 25 11254494
rect -25 11254085 -19 11254482
rect 19 11254085 25 11254482
rect -25 11254073 25 11254085
rect -25 11174051 25 11174063
rect -25 11173654 -19 11174051
rect 19 11173654 25 11174051
rect -25 11173642 25 11173654
rect -25 11173514 25 11173526
rect -25 11173117 -19 11173514
rect 19 11173117 25 11173514
rect -25 11173105 25 11173117
rect -25 11093083 25 11093095
rect -25 11092686 -19 11093083
rect 19 11092686 25 11093083
rect -25 11092674 25 11092686
rect -25 11092546 25 11092558
rect -25 11092149 -19 11092546
rect 19 11092149 25 11092546
rect -25 11092137 25 11092149
rect -25 11012115 25 11012127
rect -25 11011718 -19 11012115
rect 19 11011718 25 11012115
rect -25 11011706 25 11011718
rect -25 11011578 25 11011590
rect -25 11011181 -19 11011578
rect 19 11011181 25 11011578
rect -25 11011169 25 11011181
rect -25 10931147 25 10931159
rect -25 10930750 -19 10931147
rect 19 10930750 25 10931147
rect -25 10930738 25 10930750
rect -25 10930610 25 10930622
rect -25 10930213 -19 10930610
rect 19 10930213 25 10930610
rect -25 10930201 25 10930213
rect -25 10850179 25 10850191
rect -25 10849782 -19 10850179
rect 19 10849782 25 10850179
rect -25 10849770 25 10849782
rect -25 10849642 25 10849654
rect -25 10849245 -19 10849642
rect 19 10849245 25 10849642
rect -25 10849233 25 10849245
rect -25 10769211 25 10769223
rect -25 10768814 -19 10769211
rect 19 10768814 25 10769211
rect -25 10768802 25 10768814
rect -25 10768674 25 10768686
rect -25 10768277 -19 10768674
rect 19 10768277 25 10768674
rect -25 10768265 25 10768277
rect -25 10688243 25 10688255
rect -25 10687846 -19 10688243
rect 19 10687846 25 10688243
rect -25 10687834 25 10687846
rect -25 10687706 25 10687718
rect -25 10687309 -19 10687706
rect 19 10687309 25 10687706
rect -25 10687297 25 10687309
rect -25 10607275 25 10607287
rect -25 10606878 -19 10607275
rect 19 10606878 25 10607275
rect -25 10606866 25 10606878
rect -25 10606738 25 10606750
rect -25 10606341 -19 10606738
rect 19 10606341 25 10606738
rect -25 10606329 25 10606341
rect -25 10526307 25 10526319
rect -25 10525910 -19 10526307
rect 19 10525910 25 10526307
rect -25 10525898 25 10525910
rect -25 10525770 25 10525782
rect -25 10525373 -19 10525770
rect 19 10525373 25 10525770
rect -25 10525361 25 10525373
rect -25 10445339 25 10445351
rect -25 10444942 -19 10445339
rect 19 10444942 25 10445339
rect -25 10444930 25 10444942
rect -25 10444802 25 10444814
rect -25 10444405 -19 10444802
rect 19 10444405 25 10444802
rect -25 10444393 25 10444405
rect -25 10364371 25 10364383
rect -25 10363974 -19 10364371
rect 19 10363974 25 10364371
rect -25 10363962 25 10363974
rect -25 10363834 25 10363846
rect -25 10363437 -19 10363834
rect 19 10363437 25 10363834
rect -25 10363425 25 10363437
rect -25 10283403 25 10283415
rect -25 10283006 -19 10283403
rect 19 10283006 25 10283403
rect -25 10282994 25 10283006
rect -25 10282866 25 10282878
rect -25 10282469 -19 10282866
rect 19 10282469 25 10282866
rect -25 10282457 25 10282469
rect -25 10202435 25 10202447
rect -25 10202038 -19 10202435
rect 19 10202038 25 10202435
rect -25 10202026 25 10202038
rect -25 10201898 25 10201910
rect -25 10201501 -19 10201898
rect 19 10201501 25 10201898
rect -25 10201489 25 10201501
rect -25 10121467 25 10121479
rect -25 10121070 -19 10121467
rect 19 10121070 25 10121467
rect -25 10121058 25 10121070
rect -25 10120930 25 10120942
rect -25 10120533 -19 10120930
rect 19 10120533 25 10120930
rect -25 10120521 25 10120533
rect -25 10040499 25 10040511
rect -25 10040102 -19 10040499
rect 19 10040102 25 10040499
rect -25 10040090 25 10040102
rect -25 10039962 25 10039974
rect -25 10039565 -19 10039962
rect 19 10039565 25 10039962
rect -25 10039553 25 10039565
rect -25 9959531 25 9959543
rect -25 9959134 -19 9959531
rect 19 9959134 25 9959531
rect -25 9959122 25 9959134
rect -25 9958994 25 9959006
rect -25 9958597 -19 9958994
rect 19 9958597 25 9958994
rect -25 9958585 25 9958597
rect -25 9878563 25 9878575
rect -25 9878166 -19 9878563
rect 19 9878166 25 9878563
rect -25 9878154 25 9878166
rect -25 9878026 25 9878038
rect -25 9877629 -19 9878026
rect 19 9877629 25 9878026
rect -25 9877617 25 9877629
rect -25 9797595 25 9797607
rect -25 9797198 -19 9797595
rect 19 9797198 25 9797595
rect -25 9797186 25 9797198
rect -25 9797058 25 9797070
rect -25 9796661 -19 9797058
rect 19 9796661 25 9797058
rect -25 9796649 25 9796661
rect -25 9716627 25 9716639
rect -25 9716230 -19 9716627
rect 19 9716230 25 9716627
rect -25 9716218 25 9716230
rect -25 9716090 25 9716102
rect -25 9715693 -19 9716090
rect 19 9715693 25 9716090
rect -25 9715681 25 9715693
rect -25 9635659 25 9635671
rect -25 9635262 -19 9635659
rect 19 9635262 25 9635659
rect -25 9635250 25 9635262
rect -25 9635122 25 9635134
rect -25 9634725 -19 9635122
rect 19 9634725 25 9635122
rect -25 9634713 25 9634725
rect -25 9554691 25 9554703
rect -25 9554294 -19 9554691
rect 19 9554294 25 9554691
rect -25 9554282 25 9554294
rect -25 9554154 25 9554166
rect -25 9553757 -19 9554154
rect 19 9553757 25 9554154
rect -25 9553745 25 9553757
rect -25 9473723 25 9473735
rect -25 9473326 -19 9473723
rect 19 9473326 25 9473723
rect -25 9473314 25 9473326
rect -25 9473186 25 9473198
rect -25 9472789 -19 9473186
rect 19 9472789 25 9473186
rect -25 9472777 25 9472789
rect -25 9392755 25 9392767
rect -25 9392358 -19 9392755
rect 19 9392358 25 9392755
rect -25 9392346 25 9392358
rect -25 9392218 25 9392230
rect -25 9391821 -19 9392218
rect 19 9391821 25 9392218
rect -25 9391809 25 9391821
rect -25 9311787 25 9311799
rect -25 9311390 -19 9311787
rect 19 9311390 25 9311787
rect -25 9311378 25 9311390
rect -25 9311250 25 9311262
rect -25 9310853 -19 9311250
rect 19 9310853 25 9311250
rect -25 9310841 25 9310853
rect -25 9230819 25 9230831
rect -25 9230422 -19 9230819
rect 19 9230422 25 9230819
rect -25 9230410 25 9230422
rect -25 9230282 25 9230294
rect -25 9229885 -19 9230282
rect 19 9229885 25 9230282
rect -25 9229873 25 9229885
rect -25 9149851 25 9149863
rect -25 9149454 -19 9149851
rect 19 9149454 25 9149851
rect -25 9149442 25 9149454
rect -25 9149314 25 9149326
rect -25 9148917 -19 9149314
rect 19 9148917 25 9149314
rect -25 9148905 25 9148917
rect -25 9068883 25 9068895
rect -25 9068486 -19 9068883
rect 19 9068486 25 9068883
rect -25 9068474 25 9068486
rect -25 9068346 25 9068358
rect -25 9067949 -19 9068346
rect 19 9067949 25 9068346
rect -25 9067937 25 9067949
rect -25 8987915 25 8987927
rect -25 8987518 -19 8987915
rect 19 8987518 25 8987915
rect -25 8987506 25 8987518
rect -25 8987378 25 8987390
rect -25 8986981 -19 8987378
rect 19 8986981 25 8987378
rect -25 8986969 25 8986981
rect -25 8906947 25 8906959
rect -25 8906550 -19 8906947
rect 19 8906550 25 8906947
rect -25 8906538 25 8906550
rect -25 8906410 25 8906422
rect -25 8906013 -19 8906410
rect 19 8906013 25 8906410
rect -25 8906001 25 8906013
rect -25 8825979 25 8825991
rect -25 8825582 -19 8825979
rect 19 8825582 25 8825979
rect -25 8825570 25 8825582
rect -25 8825442 25 8825454
rect -25 8825045 -19 8825442
rect 19 8825045 25 8825442
rect -25 8825033 25 8825045
rect -25 8745011 25 8745023
rect -25 8744614 -19 8745011
rect 19 8744614 25 8745011
rect -25 8744602 25 8744614
rect -25 8744474 25 8744486
rect -25 8744077 -19 8744474
rect 19 8744077 25 8744474
rect -25 8744065 25 8744077
rect -25 8664043 25 8664055
rect -25 8663646 -19 8664043
rect 19 8663646 25 8664043
rect -25 8663634 25 8663646
rect -25 8663506 25 8663518
rect -25 8663109 -19 8663506
rect 19 8663109 25 8663506
rect -25 8663097 25 8663109
rect -25 8583075 25 8583087
rect -25 8582678 -19 8583075
rect 19 8582678 25 8583075
rect -25 8582666 25 8582678
rect -25 8582538 25 8582550
rect -25 8582141 -19 8582538
rect 19 8582141 25 8582538
rect -25 8582129 25 8582141
rect -25 8502107 25 8502119
rect -25 8501710 -19 8502107
rect 19 8501710 25 8502107
rect -25 8501698 25 8501710
rect -25 8501570 25 8501582
rect -25 8501173 -19 8501570
rect 19 8501173 25 8501570
rect -25 8501161 25 8501173
rect -25 8421139 25 8421151
rect -25 8420742 -19 8421139
rect 19 8420742 25 8421139
rect -25 8420730 25 8420742
rect -25 8420602 25 8420614
rect -25 8420205 -19 8420602
rect 19 8420205 25 8420602
rect -25 8420193 25 8420205
rect -25 8340171 25 8340183
rect -25 8339774 -19 8340171
rect 19 8339774 25 8340171
rect -25 8339762 25 8339774
rect -25 8339634 25 8339646
rect -25 8339237 -19 8339634
rect 19 8339237 25 8339634
rect -25 8339225 25 8339237
rect -25 8259203 25 8259215
rect -25 8258806 -19 8259203
rect 19 8258806 25 8259203
rect -25 8258794 25 8258806
rect -25 8258666 25 8258678
rect -25 8258269 -19 8258666
rect 19 8258269 25 8258666
rect -25 8258257 25 8258269
rect -25 8178235 25 8178247
rect -25 8177838 -19 8178235
rect 19 8177838 25 8178235
rect -25 8177826 25 8177838
rect -25 8177698 25 8177710
rect -25 8177301 -19 8177698
rect 19 8177301 25 8177698
rect -25 8177289 25 8177301
rect -25 8097267 25 8097279
rect -25 8096870 -19 8097267
rect 19 8096870 25 8097267
rect -25 8096858 25 8096870
rect -25 8096730 25 8096742
rect -25 8096333 -19 8096730
rect 19 8096333 25 8096730
rect -25 8096321 25 8096333
rect -25 8016299 25 8016311
rect -25 8015902 -19 8016299
rect 19 8015902 25 8016299
rect -25 8015890 25 8015902
rect -25 8015762 25 8015774
rect -25 8015365 -19 8015762
rect 19 8015365 25 8015762
rect -25 8015353 25 8015365
rect -25 7935331 25 7935343
rect -25 7934934 -19 7935331
rect 19 7934934 25 7935331
rect -25 7934922 25 7934934
rect -25 7934794 25 7934806
rect -25 7934397 -19 7934794
rect 19 7934397 25 7934794
rect -25 7934385 25 7934397
rect -25 7854363 25 7854375
rect -25 7853966 -19 7854363
rect 19 7853966 25 7854363
rect -25 7853954 25 7853966
rect -25 7853826 25 7853838
rect -25 7853429 -19 7853826
rect 19 7853429 25 7853826
rect -25 7853417 25 7853429
rect -25 7773395 25 7773407
rect -25 7772998 -19 7773395
rect 19 7772998 25 7773395
rect -25 7772986 25 7772998
rect -25 7772858 25 7772870
rect -25 7772461 -19 7772858
rect 19 7772461 25 7772858
rect -25 7772449 25 7772461
rect -25 7692427 25 7692439
rect -25 7692030 -19 7692427
rect 19 7692030 25 7692427
rect -25 7692018 25 7692030
rect -25 7691890 25 7691902
rect -25 7691493 -19 7691890
rect 19 7691493 25 7691890
rect -25 7691481 25 7691493
rect -25 7611459 25 7611471
rect -25 7611062 -19 7611459
rect 19 7611062 25 7611459
rect -25 7611050 25 7611062
rect -25 7610922 25 7610934
rect -25 7610525 -19 7610922
rect 19 7610525 25 7610922
rect -25 7610513 25 7610525
rect -25 7530491 25 7530503
rect -25 7530094 -19 7530491
rect 19 7530094 25 7530491
rect -25 7530082 25 7530094
rect -25 7529954 25 7529966
rect -25 7529557 -19 7529954
rect 19 7529557 25 7529954
rect -25 7529545 25 7529557
rect -25 7449523 25 7449535
rect -25 7449126 -19 7449523
rect 19 7449126 25 7449523
rect -25 7449114 25 7449126
rect -25 7448986 25 7448998
rect -25 7448589 -19 7448986
rect 19 7448589 25 7448986
rect -25 7448577 25 7448589
rect -25 7368555 25 7368567
rect -25 7368158 -19 7368555
rect 19 7368158 25 7368555
rect -25 7368146 25 7368158
rect -25 7368018 25 7368030
rect -25 7367621 -19 7368018
rect 19 7367621 25 7368018
rect -25 7367609 25 7367621
rect -25 7287587 25 7287599
rect -25 7287190 -19 7287587
rect 19 7287190 25 7287587
rect -25 7287178 25 7287190
rect -25 7287050 25 7287062
rect -25 7286653 -19 7287050
rect 19 7286653 25 7287050
rect -25 7286641 25 7286653
rect -25 7206619 25 7206631
rect -25 7206222 -19 7206619
rect 19 7206222 25 7206619
rect -25 7206210 25 7206222
rect -25 7206082 25 7206094
rect -25 7205685 -19 7206082
rect 19 7205685 25 7206082
rect -25 7205673 25 7205685
rect -25 7125651 25 7125663
rect -25 7125254 -19 7125651
rect 19 7125254 25 7125651
rect -25 7125242 25 7125254
rect -25 7125114 25 7125126
rect -25 7124717 -19 7125114
rect 19 7124717 25 7125114
rect -25 7124705 25 7124717
rect -25 7044683 25 7044695
rect -25 7044286 -19 7044683
rect 19 7044286 25 7044683
rect -25 7044274 25 7044286
rect -25 7044146 25 7044158
rect -25 7043749 -19 7044146
rect 19 7043749 25 7044146
rect -25 7043737 25 7043749
rect -25 6963715 25 6963727
rect -25 6963318 -19 6963715
rect 19 6963318 25 6963715
rect -25 6963306 25 6963318
rect -25 6963178 25 6963190
rect -25 6962781 -19 6963178
rect 19 6962781 25 6963178
rect -25 6962769 25 6962781
rect -25 6882747 25 6882759
rect -25 6882350 -19 6882747
rect 19 6882350 25 6882747
rect -25 6882338 25 6882350
rect -25 6882210 25 6882222
rect -25 6881813 -19 6882210
rect 19 6881813 25 6882210
rect -25 6881801 25 6881813
rect -25 6801779 25 6801791
rect -25 6801382 -19 6801779
rect 19 6801382 25 6801779
rect -25 6801370 25 6801382
rect -25 6801242 25 6801254
rect -25 6800845 -19 6801242
rect 19 6800845 25 6801242
rect -25 6800833 25 6800845
rect -25 6720811 25 6720823
rect -25 6720414 -19 6720811
rect 19 6720414 25 6720811
rect -25 6720402 25 6720414
rect -25 6720274 25 6720286
rect -25 6719877 -19 6720274
rect 19 6719877 25 6720274
rect -25 6719865 25 6719877
rect -25 6639843 25 6639855
rect -25 6639446 -19 6639843
rect 19 6639446 25 6639843
rect -25 6639434 25 6639446
rect -25 6639306 25 6639318
rect -25 6638909 -19 6639306
rect 19 6638909 25 6639306
rect -25 6638897 25 6638909
rect -25 6558875 25 6558887
rect -25 6558478 -19 6558875
rect 19 6558478 25 6558875
rect -25 6558466 25 6558478
rect -25 6558338 25 6558350
rect -25 6557941 -19 6558338
rect 19 6557941 25 6558338
rect -25 6557929 25 6557941
rect -25 6477907 25 6477919
rect -25 6477510 -19 6477907
rect 19 6477510 25 6477907
rect -25 6477498 25 6477510
rect -25 6477370 25 6477382
rect -25 6476973 -19 6477370
rect 19 6476973 25 6477370
rect -25 6476961 25 6476973
rect -25 6396939 25 6396951
rect -25 6396542 -19 6396939
rect 19 6396542 25 6396939
rect -25 6396530 25 6396542
rect -25 6396402 25 6396414
rect -25 6396005 -19 6396402
rect 19 6396005 25 6396402
rect -25 6395993 25 6396005
rect -25 6315971 25 6315983
rect -25 6315574 -19 6315971
rect 19 6315574 25 6315971
rect -25 6315562 25 6315574
rect -25 6315434 25 6315446
rect -25 6315037 -19 6315434
rect 19 6315037 25 6315434
rect -25 6315025 25 6315037
rect -25 6235003 25 6235015
rect -25 6234606 -19 6235003
rect 19 6234606 25 6235003
rect -25 6234594 25 6234606
rect -25 6234466 25 6234478
rect -25 6234069 -19 6234466
rect 19 6234069 25 6234466
rect -25 6234057 25 6234069
rect -25 6154035 25 6154047
rect -25 6153638 -19 6154035
rect 19 6153638 25 6154035
rect -25 6153626 25 6153638
rect -25 6153498 25 6153510
rect -25 6153101 -19 6153498
rect 19 6153101 25 6153498
rect -25 6153089 25 6153101
rect -25 6073067 25 6073079
rect -25 6072670 -19 6073067
rect 19 6072670 25 6073067
rect -25 6072658 25 6072670
rect -25 6072530 25 6072542
rect -25 6072133 -19 6072530
rect 19 6072133 25 6072530
rect -25 6072121 25 6072133
rect -25 5992099 25 5992111
rect -25 5991702 -19 5992099
rect 19 5991702 25 5992099
rect -25 5991690 25 5991702
rect -25 5991562 25 5991574
rect -25 5991165 -19 5991562
rect 19 5991165 25 5991562
rect -25 5991153 25 5991165
rect -25 5911131 25 5911143
rect -25 5910734 -19 5911131
rect 19 5910734 25 5911131
rect -25 5910722 25 5910734
rect -25 5910594 25 5910606
rect -25 5910197 -19 5910594
rect 19 5910197 25 5910594
rect -25 5910185 25 5910197
rect -25 5830163 25 5830175
rect -25 5829766 -19 5830163
rect 19 5829766 25 5830163
rect -25 5829754 25 5829766
rect -25 5829626 25 5829638
rect -25 5829229 -19 5829626
rect 19 5829229 25 5829626
rect -25 5829217 25 5829229
rect -25 5749195 25 5749207
rect -25 5748798 -19 5749195
rect 19 5748798 25 5749195
rect -25 5748786 25 5748798
rect -25 5748658 25 5748670
rect -25 5748261 -19 5748658
rect 19 5748261 25 5748658
rect -25 5748249 25 5748261
rect -25 5668227 25 5668239
rect -25 5667830 -19 5668227
rect 19 5667830 25 5668227
rect -25 5667818 25 5667830
rect -25 5667690 25 5667702
rect -25 5667293 -19 5667690
rect 19 5667293 25 5667690
rect -25 5667281 25 5667293
rect -25 5587259 25 5587271
rect -25 5586862 -19 5587259
rect 19 5586862 25 5587259
rect -25 5586850 25 5586862
rect -25 5586722 25 5586734
rect -25 5586325 -19 5586722
rect 19 5586325 25 5586722
rect -25 5586313 25 5586325
rect -25 5506291 25 5506303
rect -25 5505894 -19 5506291
rect 19 5505894 25 5506291
rect -25 5505882 25 5505894
rect -25 5505754 25 5505766
rect -25 5505357 -19 5505754
rect 19 5505357 25 5505754
rect -25 5505345 25 5505357
rect -25 5425323 25 5425335
rect -25 5424926 -19 5425323
rect 19 5424926 25 5425323
rect -25 5424914 25 5424926
rect -25 5424786 25 5424798
rect -25 5424389 -19 5424786
rect 19 5424389 25 5424786
rect -25 5424377 25 5424389
rect -25 5344355 25 5344367
rect -25 5343958 -19 5344355
rect 19 5343958 25 5344355
rect -25 5343946 25 5343958
rect -25 5343818 25 5343830
rect -25 5343421 -19 5343818
rect 19 5343421 25 5343818
rect -25 5343409 25 5343421
rect -25 5263387 25 5263399
rect -25 5262990 -19 5263387
rect 19 5262990 25 5263387
rect -25 5262978 25 5262990
rect -25 5262850 25 5262862
rect -25 5262453 -19 5262850
rect 19 5262453 25 5262850
rect -25 5262441 25 5262453
rect -25 5182419 25 5182431
rect -25 5182022 -19 5182419
rect 19 5182022 25 5182419
rect -25 5182010 25 5182022
rect -25 5181882 25 5181894
rect -25 5181485 -19 5181882
rect 19 5181485 25 5181882
rect -25 5181473 25 5181485
rect -25 5101451 25 5101463
rect -25 5101054 -19 5101451
rect 19 5101054 25 5101451
rect -25 5101042 25 5101054
rect -25 5100914 25 5100926
rect -25 5100517 -19 5100914
rect 19 5100517 25 5100914
rect -25 5100505 25 5100517
rect -25 5020483 25 5020495
rect -25 5020086 -19 5020483
rect 19 5020086 25 5020483
rect -25 5020074 25 5020086
rect -25 5019946 25 5019958
rect -25 5019549 -19 5019946
rect 19 5019549 25 5019946
rect -25 5019537 25 5019549
rect -25 4939515 25 4939527
rect -25 4939118 -19 4939515
rect 19 4939118 25 4939515
rect -25 4939106 25 4939118
rect -25 4938978 25 4938990
rect -25 4938581 -19 4938978
rect 19 4938581 25 4938978
rect -25 4938569 25 4938581
rect -25 4858547 25 4858559
rect -25 4858150 -19 4858547
rect 19 4858150 25 4858547
rect -25 4858138 25 4858150
rect -25 4858010 25 4858022
rect -25 4857613 -19 4858010
rect 19 4857613 25 4858010
rect -25 4857601 25 4857613
rect -25 4777579 25 4777591
rect -25 4777182 -19 4777579
rect 19 4777182 25 4777579
rect -25 4777170 25 4777182
rect -25 4777042 25 4777054
rect -25 4776645 -19 4777042
rect 19 4776645 25 4777042
rect -25 4776633 25 4776645
rect -25 4696611 25 4696623
rect -25 4696214 -19 4696611
rect 19 4696214 25 4696611
rect -25 4696202 25 4696214
rect -25 4696074 25 4696086
rect -25 4695677 -19 4696074
rect 19 4695677 25 4696074
rect -25 4695665 25 4695677
rect -25 4615643 25 4615655
rect -25 4615246 -19 4615643
rect 19 4615246 25 4615643
rect -25 4615234 25 4615246
rect -25 4615106 25 4615118
rect -25 4614709 -19 4615106
rect 19 4614709 25 4615106
rect -25 4614697 25 4614709
rect -25 4534675 25 4534687
rect -25 4534278 -19 4534675
rect 19 4534278 25 4534675
rect -25 4534266 25 4534278
rect -25 4534138 25 4534150
rect -25 4533741 -19 4534138
rect 19 4533741 25 4534138
rect -25 4533729 25 4533741
rect -25 4453707 25 4453719
rect -25 4453310 -19 4453707
rect 19 4453310 25 4453707
rect -25 4453298 25 4453310
rect -25 4453170 25 4453182
rect -25 4452773 -19 4453170
rect 19 4452773 25 4453170
rect -25 4452761 25 4452773
rect -25 4372739 25 4372751
rect -25 4372342 -19 4372739
rect 19 4372342 25 4372739
rect -25 4372330 25 4372342
rect -25 4372202 25 4372214
rect -25 4371805 -19 4372202
rect 19 4371805 25 4372202
rect -25 4371793 25 4371805
rect -25 4291771 25 4291783
rect -25 4291374 -19 4291771
rect 19 4291374 25 4291771
rect -25 4291362 25 4291374
rect -25 4291234 25 4291246
rect -25 4290837 -19 4291234
rect 19 4290837 25 4291234
rect -25 4290825 25 4290837
rect -25 4210803 25 4210815
rect -25 4210406 -19 4210803
rect 19 4210406 25 4210803
rect -25 4210394 25 4210406
rect -25 4210266 25 4210278
rect -25 4209869 -19 4210266
rect 19 4209869 25 4210266
rect -25 4209857 25 4209869
rect -25 4129835 25 4129847
rect -25 4129438 -19 4129835
rect 19 4129438 25 4129835
rect -25 4129426 25 4129438
rect -25 4129298 25 4129310
rect -25 4128901 -19 4129298
rect 19 4128901 25 4129298
rect -25 4128889 25 4128901
rect -25 4048867 25 4048879
rect -25 4048470 -19 4048867
rect 19 4048470 25 4048867
rect -25 4048458 25 4048470
rect -25 4048330 25 4048342
rect -25 4047933 -19 4048330
rect 19 4047933 25 4048330
rect -25 4047921 25 4047933
rect -25 3967899 25 3967911
rect -25 3967502 -19 3967899
rect 19 3967502 25 3967899
rect -25 3967490 25 3967502
rect -25 3967362 25 3967374
rect -25 3966965 -19 3967362
rect 19 3966965 25 3967362
rect -25 3966953 25 3966965
rect -25 3886931 25 3886943
rect -25 3886534 -19 3886931
rect 19 3886534 25 3886931
rect -25 3886522 25 3886534
rect -25 3886394 25 3886406
rect -25 3885997 -19 3886394
rect 19 3885997 25 3886394
rect -25 3885985 25 3885997
rect -25 3805963 25 3805975
rect -25 3805566 -19 3805963
rect 19 3805566 25 3805963
rect -25 3805554 25 3805566
rect -25 3805426 25 3805438
rect -25 3805029 -19 3805426
rect 19 3805029 25 3805426
rect -25 3805017 25 3805029
rect -25 3724995 25 3725007
rect -25 3724598 -19 3724995
rect 19 3724598 25 3724995
rect -25 3724586 25 3724598
rect -25 3724458 25 3724470
rect -25 3724061 -19 3724458
rect 19 3724061 25 3724458
rect -25 3724049 25 3724061
rect -25 3644027 25 3644039
rect -25 3643630 -19 3644027
rect 19 3643630 25 3644027
rect -25 3643618 25 3643630
rect -25 3643490 25 3643502
rect -25 3643093 -19 3643490
rect 19 3643093 25 3643490
rect -25 3643081 25 3643093
rect -25 3563059 25 3563071
rect -25 3562662 -19 3563059
rect 19 3562662 25 3563059
rect -25 3562650 25 3562662
rect -25 3562522 25 3562534
rect -25 3562125 -19 3562522
rect 19 3562125 25 3562522
rect -25 3562113 25 3562125
rect -25 3482091 25 3482103
rect -25 3481694 -19 3482091
rect 19 3481694 25 3482091
rect -25 3481682 25 3481694
rect -25 3481554 25 3481566
rect -25 3481157 -19 3481554
rect 19 3481157 25 3481554
rect -25 3481145 25 3481157
rect -25 3401123 25 3401135
rect -25 3400726 -19 3401123
rect 19 3400726 25 3401123
rect -25 3400714 25 3400726
rect -25 3400586 25 3400598
rect -25 3400189 -19 3400586
rect 19 3400189 25 3400586
rect -25 3400177 25 3400189
rect -25 3320155 25 3320167
rect -25 3319758 -19 3320155
rect 19 3319758 25 3320155
rect -25 3319746 25 3319758
rect -25 3319618 25 3319630
rect -25 3319221 -19 3319618
rect 19 3319221 25 3319618
rect -25 3319209 25 3319221
rect -25 3239187 25 3239199
rect -25 3238790 -19 3239187
rect 19 3238790 25 3239187
rect -25 3238778 25 3238790
rect -25 3238650 25 3238662
rect -25 3238253 -19 3238650
rect 19 3238253 25 3238650
rect -25 3238241 25 3238253
rect -25 3158219 25 3158231
rect -25 3157822 -19 3158219
rect 19 3157822 25 3158219
rect -25 3157810 25 3157822
rect -25 3157682 25 3157694
rect -25 3157285 -19 3157682
rect 19 3157285 25 3157682
rect -25 3157273 25 3157285
rect -25 3077251 25 3077263
rect -25 3076854 -19 3077251
rect 19 3076854 25 3077251
rect -25 3076842 25 3076854
rect -25 3076714 25 3076726
rect -25 3076317 -19 3076714
rect 19 3076317 25 3076714
rect -25 3076305 25 3076317
rect -25 2996283 25 2996295
rect -25 2995886 -19 2996283
rect 19 2995886 25 2996283
rect -25 2995874 25 2995886
rect -25 2995746 25 2995758
rect -25 2995349 -19 2995746
rect 19 2995349 25 2995746
rect -25 2995337 25 2995349
rect -25 2915315 25 2915327
rect -25 2914918 -19 2915315
rect 19 2914918 25 2915315
rect -25 2914906 25 2914918
rect -25 2914778 25 2914790
rect -25 2914381 -19 2914778
rect 19 2914381 25 2914778
rect -25 2914369 25 2914381
rect -25 2834347 25 2834359
rect -25 2833950 -19 2834347
rect 19 2833950 25 2834347
rect -25 2833938 25 2833950
rect -25 2833810 25 2833822
rect -25 2833413 -19 2833810
rect 19 2833413 25 2833810
rect -25 2833401 25 2833413
rect -25 2753379 25 2753391
rect -25 2752982 -19 2753379
rect 19 2752982 25 2753379
rect -25 2752970 25 2752982
rect -25 2752842 25 2752854
rect -25 2752445 -19 2752842
rect 19 2752445 25 2752842
rect -25 2752433 25 2752445
rect -25 2672411 25 2672423
rect -25 2672014 -19 2672411
rect 19 2672014 25 2672411
rect -25 2672002 25 2672014
rect -25 2671874 25 2671886
rect -25 2671477 -19 2671874
rect 19 2671477 25 2671874
rect -25 2671465 25 2671477
rect -25 2591443 25 2591455
rect -25 2591046 -19 2591443
rect 19 2591046 25 2591443
rect -25 2591034 25 2591046
rect -25 2590906 25 2590918
rect -25 2590509 -19 2590906
rect 19 2590509 25 2590906
rect -25 2590497 25 2590509
rect -25 2510475 25 2510487
rect -25 2510078 -19 2510475
rect 19 2510078 25 2510475
rect -25 2510066 25 2510078
rect -25 2509938 25 2509950
rect -25 2509541 -19 2509938
rect 19 2509541 25 2509938
rect -25 2509529 25 2509541
rect -25 2429507 25 2429519
rect -25 2429110 -19 2429507
rect 19 2429110 25 2429507
rect -25 2429098 25 2429110
rect -25 2428970 25 2428982
rect -25 2428573 -19 2428970
rect 19 2428573 25 2428970
rect -25 2428561 25 2428573
rect -25 2348539 25 2348551
rect -25 2348142 -19 2348539
rect 19 2348142 25 2348539
rect -25 2348130 25 2348142
rect -25 2348002 25 2348014
rect -25 2347605 -19 2348002
rect 19 2347605 25 2348002
rect -25 2347593 25 2347605
rect -25 2267571 25 2267583
rect -25 2267174 -19 2267571
rect 19 2267174 25 2267571
rect -25 2267162 25 2267174
rect -25 2267034 25 2267046
rect -25 2266637 -19 2267034
rect 19 2266637 25 2267034
rect -25 2266625 25 2266637
rect -25 2186603 25 2186615
rect -25 2186206 -19 2186603
rect 19 2186206 25 2186603
rect -25 2186194 25 2186206
rect -25 2186066 25 2186078
rect -25 2185669 -19 2186066
rect 19 2185669 25 2186066
rect -25 2185657 25 2185669
rect -25 2105635 25 2105647
rect -25 2105238 -19 2105635
rect 19 2105238 25 2105635
rect -25 2105226 25 2105238
rect -25 2105098 25 2105110
rect -25 2104701 -19 2105098
rect 19 2104701 25 2105098
rect -25 2104689 25 2104701
rect -25 2024667 25 2024679
rect -25 2024270 -19 2024667
rect 19 2024270 25 2024667
rect -25 2024258 25 2024270
rect -25 2024130 25 2024142
rect -25 2023733 -19 2024130
rect 19 2023733 25 2024130
rect -25 2023721 25 2023733
rect -25 1943699 25 1943711
rect -25 1943302 -19 1943699
rect 19 1943302 25 1943699
rect -25 1943290 25 1943302
rect -25 1943162 25 1943174
rect -25 1942765 -19 1943162
rect 19 1942765 25 1943162
rect -25 1942753 25 1942765
rect -25 1862731 25 1862743
rect -25 1862334 -19 1862731
rect 19 1862334 25 1862731
rect -25 1862322 25 1862334
rect -25 1862194 25 1862206
rect -25 1861797 -19 1862194
rect 19 1861797 25 1862194
rect -25 1861785 25 1861797
rect -25 1781763 25 1781775
rect -25 1781366 -19 1781763
rect 19 1781366 25 1781763
rect -25 1781354 25 1781366
rect -25 1781226 25 1781238
rect -25 1780829 -19 1781226
rect 19 1780829 25 1781226
rect -25 1780817 25 1780829
rect -25 1700795 25 1700807
rect -25 1700398 -19 1700795
rect 19 1700398 25 1700795
rect -25 1700386 25 1700398
rect -25 1700258 25 1700270
rect -25 1699861 -19 1700258
rect 19 1699861 25 1700258
rect -25 1699849 25 1699861
rect -25 1619827 25 1619839
rect -25 1619430 -19 1619827
rect 19 1619430 25 1619827
rect -25 1619418 25 1619430
rect -25 1619290 25 1619302
rect -25 1618893 -19 1619290
rect 19 1618893 25 1619290
rect -25 1618881 25 1618893
rect -25 1538859 25 1538871
rect -25 1538462 -19 1538859
rect 19 1538462 25 1538859
rect -25 1538450 25 1538462
rect -25 1538322 25 1538334
rect -25 1537925 -19 1538322
rect 19 1537925 25 1538322
rect -25 1537913 25 1537925
rect -25 1457891 25 1457903
rect -25 1457494 -19 1457891
rect 19 1457494 25 1457891
rect -25 1457482 25 1457494
rect -25 1457354 25 1457366
rect -25 1456957 -19 1457354
rect 19 1456957 25 1457354
rect -25 1456945 25 1456957
rect -25 1376923 25 1376935
rect -25 1376526 -19 1376923
rect 19 1376526 25 1376923
rect -25 1376514 25 1376526
rect -25 1376386 25 1376398
rect -25 1375989 -19 1376386
rect 19 1375989 25 1376386
rect -25 1375977 25 1375989
rect -25 1295955 25 1295967
rect -25 1295558 -19 1295955
rect 19 1295558 25 1295955
rect -25 1295546 25 1295558
rect -25 1295418 25 1295430
rect -25 1295021 -19 1295418
rect 19 1295021 25 1295418
rect -25 1295009 25 1295021
rect -25 1214987 25 1214999
rect -25 1214590 -19 1214987
rect 19 1214590 25 1214987
rect -25 1214578 25 1214590
rect -25 1214450 25 1214462
rect -25 1214053 -19 1214450
rect 19 1214053 25 1214450
rect -25 1214041 25 1214053
rect -25 1134019 25 1134031
rect -25 1133622 -19 1134019
rect 19 1133622 25 1134019
rect -25 1133610 25 1133622
rect -25 1133482 25 1133494
rect -25 1133085 -19 1133482
rect 19 1133085 25 1133482
rect -25 1133073 25 1133085
rect -25 1053051 25 1053063
rect -25 1052654 -19 1053051
rect 19 1052654 25 1053051
rect -25 1052642 25 1052654
rect -25 1052514 25 1052526
rect -25 1052117 -19 1052514
rect 19 1052117 25 1052514
rect -25 1052105 25 1052117
rect -25 972083 25 972095
rect -25 971686 -19 972083
rect 19 971686 25 972083
rect -25 971674 25 971686
rect -25 971546 25 971558
rect -25 971149 -19 971546
rect 19 971149 25 971546
rect -25 971137 25 971149
rect -25 891115 25 891127
rect -25 890718 -19 891115
rect 19 890718 25 891115
rect -25 890706 25 890718
rect -25 890578 25 890590
rect -25 890181 -19 890578
rect 19 890181 25 890578
rect -25 890169 25 890181
rect -25 810147 25 810159
rect -25 809750 -19 810147
rect 19 809750 25 810147
rect -25 809738 25 809750
rect -25 809610 25 809622
rect -25 809213 -19 809610
rect 19 809213 25 809610
rect -25 809201 25 809213
rect -25 729179 25 729191
rect -25 728782 -19 729179
rect 19 728782 25 729179
rect -25 728770 25 728782
rect -25 728642 25 728654
rect -25 728245 -19 728642
rect 19 728245 25 728642
rect -25 728233 25 728245
rect -25 648211 25 648223
rect -25 647814 -19 648211
rect 19 647814 25 648211
rect -25 647802 25 647814
rect -25 647674 25 647686
rect -25 647277 -19 647674
rect 19 647277 25 647674
rect -25 647265 25 647277
rect -25 567243 25 567255
rect -25 566846 -19 567243
rect 19 566846 25 567243
rect -25 566834 25 566846
rect -25 566706 25 566718
rect -25 566309 -19 566706
rect 19 566309 25 566706
rect -25 566297 25 566309
rect -25 486275 25 486287
rect -25 485878 -19 486275
rect 19 485878 25 486275
rect -25 485866 25 485878
rect -25 485738 25 485750
rect -25 485341 -19 485738
rect 19 485341 25 485738
rect -25 485329 25 485341
rect -25 405307 25 405319
rect -25 404910 -19 405307
rect 19 404910 25 405307
rect -25 404898 25 404910
rect -25 404770 25 404782
rect -25 404373 -19 404770
rect 19 404373 25 404770
rect -25 404361 25 404373
rect -25 324339 25 324351
rect -25 323942 -19 324339
rect 19 323942 25 324339
rect -25 323930 25 323942
rect -25 323802 25 323814
rect -25 323405 -19 323802
rect 19 323405 25 323802
rect -25 323393 25 323405
rect -25 243371 25 243383
rect -25 242974 -19 243371
rect 19 242974 25 243371
rect -25 242962 25 242974
rect -25 242834 25 242846
rect -25 242437 -19 242834
rect 19 242437 25 242834
rect -25 242425 25 242437
rect -25 162403 25 162415
rect -25 162006 -19 162403
rect 19 162006 25 162403
rect -25 161994 25 162006
rect -25 161866 25 161878
rect -25 161469 -19 161866
rect 19 161469 25 161866
rect -25 161457 25 161469
rect -25 81435 25 81447
rect -25 81038 -19 81435
rect 19 81038 25 81435
rect -25 81026 25 81038
rect -25 80898 25 80910
rect -25 80501 -19 80898
rect 19 80501 25 80898
rect -25 80489 25 80501
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect -25 -80501 25 -80489
rect -25 -80898 -19 -80501
rect 19 -80898 25 -80501
rect -25 -80910 25 -80898
rect -25 -81038 25 -81026
rect -25 -81435 -19 -81038
rect 19 -81435 25 -81038
rect -25 -81447 25 -81435
rect -25 -161469 25 -161457
rect -25 -161866 -19 -161469
rect 19 -161866 25 -161469
rect -25 -161878 25 -161866
rect -25 -162006 25 -161994
rect -25 -162403 -19 -162006
rect 19 -162403 25 -162006
rect -25 -162415 25 -162403
rect -25 -242437 25 -242425
rect -25 -242834 -19 -242437
rect 19 -242834 25 -242437
rect -25 -242846 25 -242834
rect -25 -242974 25 -242962
rect -25 -243371 -19 -242974
rect 19 -243371 25 -242974
rect -25 -243383 25 -243371
rect -25 -323405 25 -323393
rect -25 -323802 -19 -323405
rect 19 -323802 25 -323405
rect -25 -323814 25 -323802
rect -25 -323942 25 -323930
rect -25 -324339 -19 -323942
rect 19 -324339 25 -323942
rect -25 -324351 25 -324339
rect -25 -404373 25 -404361
rect -25 -404770 -19 -404373
rect 19 -404770 25 -404373
rect -25 -404782 25 -404770
rect -25 -404910 25 -404898
rect -25 -405307 -19 -404910
rect 19 -405307 25 -404910
rect -25 -405319 25 -405307
rect -25 -485341 25 -485329
rect -25 -485738 -19 -485341
rect 19 -485738 25 -485341
rect -25 -485750 25 -485738
rect -25 -485878 25 -485866
rect -25 -486275 -19 -485878
rect 19 -486275 25 -485878
rect -25 -486287 25 -486275
rect -25 -566309 25 -566297
rect -25 -566706 -19 -566309
rect 19 -566706 25 -566309
rect -25 -566718 25 -566706
rect -25 -566846 25 -566834
rect -25 -567243 -19 -566846
rect 19 -567243 25 -566846
rect -25 -567255 25 -567243
rect -25 -647277 25 -647265
rect -25 -647674 -19 -647277
rect 19 -647674 25 -647277
rect -25 -647686 25 -647674
rect -25 -647814 25 -647802
rect -25 -648211 -19 -647814
rect 19 -648211 25 -647814
rect -25 -648223 25 -648211
rect -25 -728245 25 -728233
rect -25 -728642 -19 -728245
rect 19 -728642 25 -728245
rect -25 -728654 25 -728642
rect -25 -728782 25 -728770
rect -25 -729179 -19 -728782
rect 19 -729179 25 -728782
rect -25 -729191 25 -729179
rect -25 -809213 25 -809201
rect -25 -809610 -19 -809213
rect 19 -809610 25 -809213
rect -25 -809622 25 -809610
rect -25 -809750 25 -809738
rect -25 -810147 -19 -809750
rect 19 -810147 25 -809750
rect -25 -810159 25 -810147
rect -25 -890181 25 -890169
rect -25 -890578 -19 -890181
rect 19 -890578 25 -890181
rect -25 -890590 25 -890578
rect -25 -890718 25 -890706
rect -25 -891115 -19 -890718
rect 19 -891115 25 -890718
rect -25 -891127 25 -891115
rect -25 -971149 25 -971137
rect -25 -971546 -19 -971149
rect 19 -971546 25 -971149
rect -25 -971558 25 -971546
rect -25 -971686 25 -971674
rect -25 -972083 -19 -971686
rect 19 -972083 25 -971686
rect -25 -972095 25 -972083
rect -25 -1052117 25 -1052105
rect -25 -1052514 -19 -1052117
rect 19 -1052514 25 -1052117
rect -25 -1052526 25 -1052514
rect -25 -1052654 25 -1052642
rect -25 -1053051 -19 -1052654
rect 19 -1053051 25 -1052654
rect -25 -1053063 25 -1053051
rect -25 -1133085 25 -1133073
rect -25 -1133482 -19 -1133085
rect 19 -1133482 25 -1133085
rect -25 -1133494 25 -1133482
rect -25 -1133622 25 -1133610
rect -25 -1134019 -19 -1133622
rect 19 -1134019 25 -1133622
rect -25 -1134031 25 -1134019
rect -25 -1214053 25 -1214041
rect -25 -1214450 -19 -1214053
rect 19 -1214450 25 -1214053
rect -25 -1214462 25 -1214450
rect -25 -1214590 25 -1214578
rect -25 -1214987 -19 -1214590
rect 19 -1214987 25 -1214590
rect -25 -1214999 25 -1214987
rect -25 -1295021 25 -1295009
rect -25 -1295418 -19 -1295021
rect 19 -1295418 25 -1295021
rect -25 -1295430 25 -1295418
rect -25 -1295558 25 -1295546
rect -25 -1295955 -19 -1295558
rect 19 -1295955 25 -1295558
rect -25 -1295967 25 -1295955
rect -25 -1375989 25 -1375977
rect -25 -1376386 -19 -1375989
rect 19 -1376386 25 -1375989
rect -25 -1376398 25 -1376386
rect -25 -1376526 25 -1376514
rect -25 -1376923 -19 -1376526
rect 19 -1376923 25 -1376526
rect -25 -1376935 25 -1376923
rect -25 -1456957 25 -1456945
rect -25 -1457354 -19 -1456957
rect 19 -1457354 25 -1456957
rect -25 -1457366 25 -1457354
rect -25 -1457494 25 -1457482
rect -25 -1457891 -19 -1457494
rect 19 -1457891 25 -1457494
rect -25 -1457903 25 -1457891
rect -25 -1537925 25 -1537913
rect -25 -1538322 -19 -1537925
rect 19 -1538322 25 -1537925
rect -25 -1538334 25 -1538322
rect -25 -1538462 25 -1538450
rect -25 -1538859 -19 -1538462
rect 19 -1538859 25 -1538462
rect -25 -1538871 25 -1538859
rect -25 -1618893 25 -1618881
rect -25 -1619290 -19 -1618893
rect 19 -1619290 25 -1618893
rect -25 -1619302 25 -1619290
rect -25 -1619430 25 -1619418
rect -25 -1619827 -19 -1619430
rect 19 -1619827 25 -1619430
rect -25 -1619839 25 -1619827
rect -25 -1699861 25 -1699849
rect -25 -1700258 -19 -1699861
rect 19 -1700258 25 -1699861
rect -25 -1700270 25 -1700258
rect -25 -1700398 25 -1700386
rect -25 -1700795 -19 -1700398
rect 19 -1700795 25 -1700398
rect -25 -1700807 25 -1700795
rect -25 -1780829 25 -1780817
rect -25 -1781226 -19 -1780829
rect 19 -1781226 25 -1780829
rect -25 -1781238 25 -1781226
rect -25 -1781366 25 -1781354
rect -25 -1781763 -19 -1781366
rect 19 -1781763 25 -1781366
rect -25 -1781775 25 -1781763
rect -25 -1861797 25 -1861785
rect -25 -1862194 -19 -1861797
rect 19 -1862194 25 -1861797
rect -25 -1862206 25 -1862194
rect -25 -1862334 25 -1862322
rect -25 -1862731 -19 -1862334
rect 19 -1862731 25 -1862334
rect -25 -1862743 25 -1862731
rect -25 -1942765 25 -1942753
rect -25 -1943162 -19 -1942765
rect 19 -1943162 25 -1942765
rect -25 -1943174 25 -1943162
rect -25 -1943302 25 -1943290
rect -25 -1943699 -19 -1943302
rect 19 -1943699 25 -1943302
rect -25 -1943711 25 -1943699
rect -25 -2023733 25 -2023721
rect -25 -2024130 -19 -2023733
rect 19 -2024130 25 -2023733
rect -25 -2024142 25 -2024130
rect -25 -2024270 25 -2024258
rect -25 -2024667 -19 -2024270
rect 19 -2024667 25 -2024270
rect -25 -2024679 25 -2024667
rect -25 -2104701 25 -2104689
rect -25 -2105098 -19 -2104701
rect 19 -2105098 25 -2104701
rect -25 -2105110 25 -2105098
rect -25 -2105238 25 -2105226
rect -25 -2105635 -19 -2105238
rect 19 -2105635 25 -2105238
rect -25 -2105647 25 -2105635
rect -25 -2185669 25 -2185657
rect -25 -2186066 -19 -2185669
rect 19 -2186066 25 -2185669
rect -25 -2186078 25 -2186066
rect -25 -2186206 25 -2186194
rect -25 -2186603 -19 -2186206
rect 19 -2186603 25 -2186206
rect -25 -2186615 25 -2186603
rect -25 -2266637 25 -2266625
rect -25 -2267034 -19 -2266637
rect 19 -2267034 25 -2266637
rect -25 -2267046 25 -2267034
rect -25 -2267174 25 -2267162
rect -25 -2267571 -19 -2267174
rect 19 -2267571 25 -2267174
rect -25 -2267583 25 -2267571
rect -25 -2347605 25 -2347593
rect -25 -2348002 -19 -2347605
rect 19 -2348002 25 -2347605
rect -25 -2348014 25 -2348002
rect -25 -2348142 25 -2348130
rect -25 -2348539 -19 -2348142
rect 19 -2348539 25 -2348142
rect -25 -2348551 25 -2348539
rect -25 -2428573 25 -2428561
rect -25 -2428970 -19 -2428573
rect 19 -2428970 25 -2428573
rect -25 -2428982 25 -2428970
rect -25 -2429110 25 -2429098
rect -25 -2429507 -19 -2429110
rect 19 -2429507 25 -2429110
rect -25 -2429519 25 -2429507
rect -25 -2509541 25 -2509529
rect -25 -2509938 -19 -2509541
rect 19 -2509938 25 -2509541
rect -25 -2509950 25 -2509938
rect -25 -2510078 25 -2510066
rect -25 -2510475 -19 -2510078
rect 19 -2510475 25 -2510078
rect -25 -2510487 25 -2510475
rect -25 -2590509 25 -2590497
rect -25 -2590906 -19 -2590509
rect 19 -2590906 25 -2590509
rect -25 -2590918 25 -2590906
rect -25 -2591046 25 -2591034
rect -25 -2591443 -19 -2591046
rect 19 -2591443 25 -2591046
rect -25 -2591455 25 -2591443
rect -25 -2671477 25 -2671465
rect -25 -2671874 -19 -2671477
rect 19 -2671874 25 -2671477
rect -25 -2671886 25 -2671874
rect -25 -2672014 25 -2672002
rect -25 -2672411 -19 -2672014
rect 19 -2672411 25 -2672014
rect -25 -2672423 25 -2672411
rect -25 -2752445 25 -2752433
rect -25 -2752842 -19 -2752445
rect 19 -2752842 25 -2752445
rect -25 -2752854 25 -2752842
rect -25 -2752982 25 -2752970
rect -25 -2753379 -19 -2752982
rect 19 -2753379 25 -2752982
rect -25 -2753391 25 -2753379
rect -25 -2833413 25 -2833401
rect -25 -2833810 -19 -2833413
rect 19 -2833810 25 -2833413
rect -25 -2833822 25 -2833810
rect -25 -2833950 25 -2833938
rect -25 -2834347 -19 -2833950
rect 19 -2834347 25 -2833950
rect -25 -2834359 25 -2834347
rect -25 -2914381 25 -2914369
rect -25 -2914778 -19 -2914381
rect 19 -2914778 25 -2914381
rect -25 -2914790 25 -2914778
rect -25 -2914918 25 -2914906
rect -25 -2915315 -19 -2914918
rect 19 -2915315 25 -2914918
rect -25 -2915327 25 -2915315
rect -25 -2995349 25 -2995337
rect -25 -2995746 -19 -2995349
rect 19 -2995746 25 -2995349
rect -25 -2995758 25 -2995746
rect -25 -2995886 25 -2995874
rect -25 -2996283 -19 -2995886
rect 19 -2996283 25 -2995886
rect -25 -2996295 25 -2996283
rect -25 -3076317 25 -3076305
rect -25 -3076714 -19 -3076317
rect 19 -3076714 25 -3076317
rect -25 -3076726 25 -3076714
rect -25 -3076854 25 -3076842
rect -25 -3077251 -19 -3076854
rect 19 -3077251 25 -3076854
rect -25 -3077263 25 -3077251
rect -25 -3157285 25 -3157273
rect -25 -3157682 -19 -3157285
rect 19 -3157682 25 -3157285
rect -25 -3157694 25 -3157682
rect -25 -3157822 25 -3157810
rect -25 -3158219 -19 -3157822
rect 19 -3158219 25 -3157822
rect -25 -3158231 25 -3158219
rect -25 -3238253 25 -3238241
rect -25 -3238650 -19 -3238253
rect 19 -3238650 25 -3238253
rect -25 -3238662 25 -3238650
rect -25 -3238790 25 -3238778
rect -25 -3239187 -19 -3238790
rect 19 -3239187 25 -3238790
rect -25 -3239199 25 -3239187
rect -25 -3319221 25 -3319209
rect -25 -3319618 -19 -3319221
rect 19 -3319618 25 -3319221
rect -25 -3319630 25 -3319618
rect -25 -3319758 25 -3319746
rect -25 -3320155 -19 -3319758
rect 19 -3320155 25 -3319758
rect -25 -3320167 25 -3320155
rect -25 -3400189 25 -3400177
rect -25 -3400586 -19 -3400189
rect 19 -3400586 25 -3400189
rect -25 -3400598 25 -3400586
rect -25 -3400726 25 -3400714
rect -25 -3401123 -19 -3400726
rect 19 -3401123 25 -3400726
rect -25 -3401135 25 -3401123
rect -25 -3481157 25 -3481145
rect -25 -3481554 -19 -3481157
rect 19 -3481554 25 -3481157
rect -25 -3481566 25 -3481554
rect -25 -3481694 25 -3481682
rect -25 -3482091 -19 -3481694
rect 19 -3482091 25 -3481694
rect -25 -3482103 25 -3482091
rect -25 -3562125 25 -3562113
rect -25 -3562522 -19 -3562125
rect 19 -3562522 25 -3562125
rect -25 -3562534 25 -3562522
rect -25 -3562662 25 -3562650
rect -25 -3563059 -19 -3562662
rect 19 -3563059 25 -3562662
rect -25 -3563071 25 -3563059
rect -25 -3643093 25 -3643081
rect -25 -3643490 -19 -3643093
rect 19 -3643490 25 -3643093
rect -25 -3643502 25 -3643490
rect -25 -3643630 25 -3643618
rect -25 -3644027 -19 -3643630
rect 19 -3644027 25 -3643630
rect -25 -3644039 25 -3644027
rect -25 -3724061 25 -3724049
rect -25 -3724458 -19 -3724061
rect 19 -3724458 25 -3724061
rect -25 -3724470 25 -3724458
rect -25 -3724598 25 -3724586
rect -25 -3724995 -19 -3724598
rect 19 -3724995 25 -3724598
rect -25 -3725007 25 -3724995
rect -25 -3805029 25 -3805017
rect -25 -3805426 -19 -3805029
rect 19 -3805426 25 -3805029
rect -25 -3805438 25 -3805426
rect -25 -3805566 25 -3805554
rect -25 -3805963 -19 -3805566
rect 19 -3805963 25 -3805566
rect -25 -3805975 25 -3805963
rect -25 -3885997 25 -3885985
rect -25 -3886394 -19 -3885997
rect 19 -3886394 25 -3885997
rect -25 -3886406 25 -3886394
rect -25 -3886534 25 -3886522
rect -25 -3886931 -19 -3886534
rect 19 -3886931 25 -3886534
rect -25 -3886943 25 -3886931
rect -25 -3966965 25 -3966953
rect -25 -3967362 -19 -3966965
rect 19 -3967362 25 -3966965
rect -25 -3967374 25 -3967362
rect -25 -3967502 25 -3967490
rect -25 -3967899 -19 -3967502
rect 19 -3967899 25 -3967502
rect -25 -3967911 25 -3967899
rect -25 -4047933 25 -4047921
rect -25 -4048330 -19 -4047933
rect 19 -4048330 25 -4047933
rect -25 -4048342 25 -4048330
rect -25 -4048470 25 -4048458
rect -25 -4048867 -19 -4048470
rect 19 -4048867 25 -4048470
rect -25 -4048879 25 -4048867
rect -25 -4128901 25 -4128889
rect -25 -4129298 -19 -4128901
rect 19 -4129298 25 -4128901
rect -25 -4129310 25 -4129298
rect -25 -4129438 25 -4129426
rect -25 -4129835 -19 -4129438
rect 19 -4129835 25 -4129438
rect -25 -4129847 25 -4129835
rect -25 -4209869 25 -4209857
rect -25 -4210266 -19 -4209869
rect 19 -4210266 25 -4209869
rect -25 -4210278 25 -4210266
rect -25 -4210406 25 -4210394
rect -25 -4210803 -19 -4210406
rect 19 -4210803 25 -4210406
rect -25 -4210815 25 -4210803
rect -25 -4290837 25 -4290825
rect -25 -4291234 -19 -4290837
rect 19 -4291234 25 -4290837
rect -25 -4291246 25 -4291234
rect -25 -4291374 25 -4291362
rect -25 -4291771 -19 -4291374
rect 19 -4291771 25 -4291374
rect -25 -4291783 25 -4291771
rect -25 -4371805 25 -4371793
rect -25 -4372202 -19 -4371805
rect 19 -4372202 25 -4371805
rect -25 -4372214 25 -4372202
rect -25 -4372342 25 -4372330
rect -25 -4372739 -19 -4372342
rect 19 -4372739 25 -4372342
rect -25 -4372751 25 -4372739
rect -25 -4452773 25 -4452761
rect -25 -4453170 -19 -4452773
rect 19 -4453170 25 -4452773
rect -25 -4453182 25 -4453170
rect -25 -4453310 25 -4453298
rect -25 -4453707 -19 -4453310
rect 19 -4453707 25 -4453310
rect -25 -4453719 25 -4453707
rect -25 -4533741 25 -4533729
rect -25 -4534138 -19 -4533741
rect 19 -4534138 25 -4533741
rect -25 -4534150 25 -4534138
rect -25 -4534278 25 -4534266
rect -25 -4534675 -19 -4534278
rect 19 -4534675 25 -4534278
rect -25 -4534687 25 -4534675
rect -25 -4614709 25 -4614697
rect -25 -4615106 -19 -4614709
rect 19 -4615106 25 -4614709
rect -25 -4615118 25 -4615106
rect -25 -4615246 25 -4615234
rect -25 -4615643 -19 -4615246
rect 19 -4615643 25 -4615246
rect -25 -4615655 25 -4615643
rect -25 -4695677 25 -4695665
rect -25 -4696074 -19 -4695677
rect 19 -4696074 25 -4695677
rect -25 -4696086 25 -4696074
rect -25 -4696214 25 -4696202
rect -25 -4696611 -19 -4696214
rect 19 -4696611 25 -4696214
rect -25 -4696623 25 -4696611
rect -25 -4776645 25 -4776633
rect -25 -4777042 -19 -4776645
rect 19 -4777042 25 -4776645
rect -25 -4777054 25 -4777042
rect -25 -4777182 25 -4777170
rect -25 -4777579 -19 -4777182
rect 19 -4777579 25 -4777182
rect -25 -4777591 25 -4777579
rect -25 -4857613 25 -4857601
rect -25 -4858010 -19 -4857613
rect 19 -4858010 25 -4857613
rect -25 -4858022 25 -4858010
rect -25 -4858150 25 -4858138
rect -25 -4858547 -19 -4858150
rect 19 -4858547 25 -4858150
rect -25 -4858559 25 -4858547
rect -25 -4938581 25 -4938569
rect -25 -4938978 -19 -4938581
rect 19 -4938978 25 -4938581
rect -25 -4938990 25 -4938978
rect -25 -4939118 25 -4939106
rect -25 -4939515 -19 -4939118
rect 19 -4939515 25 -4939118
rect -25 -4939527 25 -4939515
rect -25 -5019549 25 -5019537
rect -25 -5019946 -19 -5019549
rect 19 -5019946 25 -5019549
rect -25 -5019958 25 -5019946
rect -25 -5020086 25 -5020074
rect -25 -5020483 -19 -5020086
rect 19 -5020483 25 -5020086
rect -25 -5020495 25 -5020483
rect -25 -5100517 25 -5100505
rect -25 -5100914 -19 -5100517
rect 19 -5100914 25 -5100517
rect -25 -5100926 25 -5100914
rect -25 -5101054 25 -5101042
rect -25 -5101451 -19 -5101054
rect 19 -5101451 25 -5101054
rect -25 -5101463 25 -5101451
rect -25 -5181485 25 -5181473
rect -25 -5181882 -19 -5181485
rect 19 -5181882 25 -5181485
rect -25 -5181894 25 -5181882
rect -25 -5182022 25 -5182010
rect -25 -5182419 -19 -5182022
rect 19 -5182419 25 -5182022
rect -25 -5182431 25 -5182419
rect -25 -5262453 25 -5262441
rect -25 -5262850 -19 -5262453
rect 19 -5262850 25 -5262453
rect -25 -5262862 25 -5262850
rect -25 -5262990 25 -5262978
rect -25 -5263387 -19 -5262990
rect 19 -5263387 25 -5262990
rect -25 -5263399 25 -5263387
rect -25 -5343421 25 -5343409
rect -25 -5343818 -19 -5343421
rect 19 -5343818 25 -5343421
rect -25 -5343830 25 -5343818
rect -25 -5343958 25 -5343946
rect -25 -5344355 -19 -5343958
rect 19 -5344355 25 -5343958
rect -25 -5344367 25 -5344355
rect -25 -5424389 25 -5424377
rect -25 -5424786 -19 -5424389
rect 19 -5424786 25 -5424389
rect -25 -5424798 25 -5424786
rect -25 -5424926 25 -5424914
rect -25 -5425323 -19 -5424926
rect 19 -5425323 25 -5424926
rect -25 -5425335 25 -5425323
rect -25 -5505357 25 -5505345
rect -25 -5505754 -19 -5505357
rect 19 -5505754 25 -5505357
rect -25 -5505766 25 -5505754
rect -25 -5505894 25 -5505882
rect -25 -5506291 -19 -5505894
rect 19 -5506291 25 -5505894
rect -25 -5506303 25 -5506291
rect -25 -5586325 25 -5586313
rect -25 -5586722 -19 -5586325
rect 19 -5586722 25 -5586325
rect -25 -5586734 25 -5586722
rect -25 -5586862 25 -5586850
rect -25 -5587259 -19 -5586862
rect 19 -5587259 25 -5586862
rect -25 -5587271 25 -5587259
rect -25 -5667293 25 -5667281
rect -25 -5667690 -19 -5667293
rect 19 -5667690 25 -5667293
rect -25 -5667702 25 -5667690
rect -25 -5667830 25 -5667818
rect -25 -5668227 -19 -5667830
rect 19 -5668227 25 -5667830
rect -25 -5668239 25 -5668227
rect -25 -5748261 25 -5748249
rect -25 -5748658 -19 -5748261
rect 19 -5748658 25 -5748261
rect -25 -5748670 25 -5748658
rect -25 -5748798 25 -5748786
rect -25 -5749195 -19 -5748798
rect 19 -5749195 25 -5748798
rect -25 -5749207 25 -5749195
rect -25 -5829229 25 -5829217
rect -25 -5829626 -19 -5829229
rect 19 -5829626 25 -5829229
rect -25 -5829638 25 -5829626
rect -25 -5829766 25 -5829754
rect -25 -5830163 -19 -5829766
rect 19 -5830163 25 -5829766
rect -25 -5830175 25 -5830163
rect -25 -5910197 25 -5910185
rect -25 -5910594 -19 -5910197
rect 19 -5910594 25 -5910197
rect -25 -5910606 25 -5910594
rect -25 -5910734 25 -5910722
rect -25 -5911131 -19 -5910734
rect 19 -5911131 25 -5910734
rect -25 -5911143 25 -5911131
rect -25 -5991165 25 -5991153
rect -25 -5991562 -19 -5991165
rect 19 -5991562 25 -5991165
rect -25 -5991574 25 -5991562
rect -25 -5991702 25 -5991690
rect -25 -5992099 -19 -5991702
rect 19 -5992099 25 -5991702
rect -25 -5992111 25 -5992099
rect -25 -6072133 25 -6072121
rect -25 -6072530 -19 -6072133
rect 19 -6072530 25 -6072133
rect -25 -6072542 25 -6072530
rect -25 -6072670 25 -6072658
rect -25 -6073067 -19 -6072670
rect 19 -6073067 25 -6072670
rect -25 -6073079 25 -6073067
rect -25 -6153101 25 -6153089
rect -25 -6153498 -19 -6153101
rect 19 -6153498 25 -6153101
rect -25 -6153510 25 -6153498
rect -25 -6153638 25 -6153626
rect -25 -6154035 -19 -6153638
rect 19 -6154035 25 -6153638
rect -25 -6154047 25 -6154035
rect -25 -6234069 25 -6234057
rect -25 -6234466 -19 -6234069
rect 19 -6234466 25 -6234069
rect -25 -6234478 25 -6234466
rect -25 -6234606 25 -6234594
rect -25 -6235003 -19 -6234606
rect 19 -6235003 25 -6234606
rect -25 -6235015 25 -6235003
rect -25 -6315037 25 -6315025
rect -25 -6315434 -19 -6315037
rect 19 -6315434 25 -6315037
rect -25 -6315446 25 -6315434
rect -25 -6315574 25 -6315562
rect -25 -6315971 -19 -6315574
rect 19 -6315971 25 -6315574
rect -25 -6315983 25 -6315971
rect -25 -6396005 25 -6395993
rect -25 -6396402 -19 -6396005
rect 19 -6396402 25 -6396005
rect -25 -6396414 25 -6396402
rect -25 -6396542 25 -6396530
rect -25 -6396939 -19 -6396542
rect 19 -6396939 25 -6396542
rect -25 -6396951 25 -6396939
rect -25 -6476973 25 -6476961
rect -25 -6477370 -19 -6476973
rect 19 -6477370 25 -6476973
rect -25 -6477382 25 -6477370
rect -25 -6477510 25 -6477498
rect -25 -6477907 -19 -6477510
rect 19 -6477907 25 -6477510
rect -25 -6477919 25 -6477907
rect -25 -6557941 25 -6557929
rect -25 -6558338 -19 -6557941
rect 19 -6558338 25 -6557941
rect -25 -6558350 25 -6558338
rect -25 -6558478 25 -6558466
rect -25 -6558875 -19 -6558478
rect 19 -6558875 25 -6558478
rect -25 -6558887 25 -6558875
rect -25 -6638909 25 -6638897
rect -25 -6639306 -19 -6638909
rect 19 -6639306 25 -6638909
rect -25 -6639318 25 -6639306
rect -25 -6639446 25 -6639434
rect -25 -6639843 -19 -6639446
rect 19 -6639843 25 -6639446
rect -25 -6639855 25 -6639843
rect -25 -6719877 25 -6719865
rect -25 -6720274 -19 -6719877
rect 19 -6720274 25 -6719877
rect -25 -6720286 25 -6720274
rect -25 -6720414 25 -6720402
rect -25 -6720811 -19 -6720414
rect 19 -6720811 25 -6720414
rect -25 -6720823 25 -6720811
rect -25 -6800845 25 -6800833
rect -25 -6801242 -19 -6800845
rect 19 -6801242 25 -6800845
rect -25 -6801254 25 -6801242
rect -25 -6801382 25 -6801370
rect -25 -6801779 -19 -6801382
rect 19 -6801779 25 -6801382
rect -25 -6801791 25 -6801779
rect -25 -6881813 25 -6881801
rect -25 -6882210 -19 -6881813
rect 19 -6882210 25 -6881813
rect -25 -6882222 25 -6882210
rect -25 -6882350 25 -6882338
rect -25 -6882747 -19 -6882350
rect 19 -6882747 25 -6882350
rect -25 -6882759 25 -6882747
rect -25 -6962781 25 -6962769
rect -25 -6963178 -19 -6962781
rect 19 -6963178 25 -6962781
rect -25 -6963190 25 -6963178
rect -25 -6963318 25 -6963306
rect -25 -6963715 -19 -6963318
rect 19 -6963715 25 -6963318
rect -25 -6963727 25 -6963715
rect -25 -7043749 25 -7043737
rect -25 -7044146 -19 -7043749
rect 19 -7044146 25 -7043749
rect -25 -7044158 25 -7044146
rect -25 -7044286 25 -7044274
rect -25 -7044683 -19 -7044286
rect 19 -7044683 25 -7044286
rect -25 -7044695 25 -7044683
rect -25 -7124717 25 -7124705
rect -25 -7125114 -19 -7124717
rect 19 -7125114 25 -7124717
rect -25 -7125126 25 -7125114
rect -25 -7125254 25 -7125242
rect -25 -7125651 -19 -7125254
rect 19 -7125651 25 -7125254
rect -25 -7125663 25 -7125651
rect -25 -7205685 25 -7205673
rect -25 -7206082 -19 -7205685
rect 19 -7206082 25 -7205685
rect -25 -7206094 25 -7206082
rect -25 -7206222 25 -7206210
rect -25 -7206619 -19 -7206222
rect 19 -7206619 25 -7206222
rect -25 -7206631 25 -7206619
rect -25 -7286653 25 -7286641
rect -25 -7287050 -19 -7286653
rect 19 -7287050 25 -7286653
rect -25 -7287062 25 -7287050
rect -25 -7287190 25 -7287178
rect -25 -7287587 -19 -7287190
rect 19 -7287587 25 -7287190
rect -25 -7287599 25 -7287587
rect -25 -7367621 25 -7367609
rect -25 -7368018 -19 -7367621
rect 19 -7368018 25 -7367621
rect -25 -7368030 25 -7368018
rect -25 -7368158 25 -7368146
rect -25 -7368555 -19 -7368158
rect 19 -7368555 25 -7368158
rect -25 -7368567 25 -7368555
rect -25 -7448589 25 -7448577
rect -25 -7448986 -19 -7448589
rect 19 -7448986 25 -7448589
rect -25 -7448998 25 -7448986
rect -25 -7449126 25 -7449114
rect -25 -7449523 -19 -7449126
rect 19 -7449523 25 -7449126
rect -25 -7449535 25 -7449523
rect -25 -7529557 25 -7529545
rect -25 -7529954 -19 -7529557
rect 19 -7529954 25 -7529557
rect -25 -7529966 25 -7529954
rect -25 -7530094 25 -7530082
rect -25 -7530491 -19 -7530094
rect 19 -7530491 25 -7530094
rect -25 -7530503 25 -7530491
rect -25 -7610525 25 -7610513
rect -25 -7610922 -19 -7610525
rect 19 -7610922 25 -7610525
rect -25 -7610934 25 -7610922
rect -25 -7611062 25 -7611050
rect -25 -7611459 -19 -7611062
rect 19 -7611459 25 -7611062
rect -25 -7611471 25 -7611459
rect -25 -7691493 25 -7691481
rect -25 -7691890 -19 -7691493
rect 19 -7691890 25 -7691493
rect -25 -7691902 25 -7691890
rect -25 -7692030 25 -7692018
rect -25 -7692427 -19 -7692030
rect 19 -7692427 25 -7692030
rect -25 -7692439 25 -7692427
rect -25 -7772461 25 -7772449
rect -25 -7772858 -19 -7772461
rect 19 -7772858 25 -7772461
rect -25 -7772870 25 -7772858
rect -25 -7772998 25 -7772986
rect -25 -7773395 -19 -7772998
rect 19 -7773395 25 -7772998
rect -25 -7773407 25 -7773395
rect -25 -7853429 25 -7853417
rect -25 -7853826 -19 -7853429
rect 19 -7853826 25 -7853429
rect -25 -7853838 25 -7853826
rect -25 -7853966 25 -7853954
rect -25 -7854363 -19 -7853966
rect 19 -7854363 25 -7853966
rect -25 -7854375 25 -7854363
rect -25 -7934397 25 -7934385
rect -25 -7934794 -19 -7934397
rect 19 -7934794 25 -7934397
rect -25 -7934806 25 -7934794
rect -25 -7934934 25 -7934922
rect -25 -7935331 -19 -7934934
rect 19 -7935331 25 -7934934
rect -25 -7935343 25 -7935331
rect -25 -8015365 25 -8015353
rect -25 -8015762 -19 -8015365
rect 19 -8015762 25 -8015365
rect -25 -8015774 25 -8015762
rect -25 -8015902 25 -8015890
rect -25 -8016299 -19 -8015902
rect 19 -8016299 25 -8015902
rect -25 -8016311 25 -8016299
rect -25 -8096333 25 -8096321
rect -25 -8096730 -19 -8096333
rect 19 -8096730 25 -8096333
rect -25 -8096742 25 -8096730
rect -25 -8096870 25 -8096858
rect -25 -8097267 -19 -8096870
rect 19 -8097267 25 -8096870
rect -25 -8097279 25 -8097267
rect -25 -8177301 25 -8177289
rect -25 -8177698 -19 -8177301
rect 19 -8177698 25 -8177301
rect -25 -8177710 25 -8177698
rect -25 -8177838 25 -8177826
rect -25 -8178235 -19 -8177838
rect 19 -8178235 25 -8177838
rect -25 -8178247 25 -8178235
rect -25 -8258269 25 -8258257
rect -25 -8258666 -19 -8258269
rect 19 -8258666 25 -8258269
rect -25 -8258678 25 -8258666
rect -25 -8258806 25 -8258794
rect -25 -8259203 -19 -8258806
rect 19 -8259203 25 -8258806
rect -25 -8259215 25 -8259203
rect -25 -8339237 25 -8339225
rect -25 -8339634 -19 -8339237
rect 19 -8339634 25 -8339237
rect -25 -8339646 25 -8339634
rect -25 -8339774 25 -8339762
rect -25 -8340171 -19 -8339774
rect 19 -8340171 25 -8339774
rect -25 -8340183 25 -8340171
rect -25 -8420205 25 -8420193
rect -25 -8420602 -19 -8420205
rect 19 -8420602 25 -8420205
rect -25 -8420614 25 -8420602
rect -25 -8420742 25 -8420730
rect -25 -8421139 -19 -8420742
rect 19 -8421139 25 -8420742
rect -25 -8421151 25 -8421139
rect -25 -8501173 25 -8501161
rect -25 -8501570 -19 -8501173
rect 19 -8501570 25 -8501173
rect -25 -8501582 25 -8501570
rect -25 -8501710 25 -8501698
rect -25 -8502107 -19 -8501710
rect 19 -8502107 25 -8501710
rect -25 -8502119 25 -8502107
rect -25 -8582141 25 -8582129
rect -25 -8582538 -19 -8582141
rect 19 -8582538 25 -8582141
rect -25 -8582550 25 -8582538
rect -25 -8582678 25 -8582666
rect -25 -8583075 -19 -8582678
rect 19 -8583075 25 -8582678
rect -25 -8583087 25 -8583075
rect -25 -8663109 25 -8663097
rect -25 -8663506 -19 -8663109
rect 19 -8663506 25 -8663109
rect -25 -8663518 25 -8663506
rect -25 -8663646 25 -8663634
rect -25 -8664043 -19 -8663646
rect 19 -8664043 25 -8663646
rect -25 -8664055 25 -8664043
rect -25 -8744077 25 -8744065
rect -25 -8744474 -19 -8744077
rect 19 -8744474 25 -8744077
rect -25 -8744486 25 -8744474
rect -25 -8744614 25 -8744602
rect -25 -8745011 -19 -8744614
rect 19 -8745011 25 -8744614
rect -25 -8745023 25 -8745011
rect -25 -8825045 25 -8825033
rect -25 -8825442 -19 -8825045
rect 19 -8825442 25 -8825045
rect -25 -8825454 25 -8825442
rect -25 -8825582 25 -8825570
rect -25 -8825979 -19 -8825582
rect 19 -8825979 25 -8825582
rect -25 -8825991 25 -8825979
rect -25 -8906013 25 -8906001
rect -25 -8906410 -19 -8906013
rect 19 -8906410 25 -8906013
rect -25 -8906422 25 -8906410
rect -25 -8906550 25 -8906538
rect -25 -8906947 -19 -8906550
rect 19 -8906947 25 -8906550
rect -25 -8906959 25 -8906947
rect -25 -8986981 25 -8986969
rect -25 -8987378 -19 -8986981
rect 19 -8987378 25 -8986981
rect -25 -8987390 25 -8987378
rect -25 -8987518 25 -8987506
rect -25 -8987915 -19 -8987518
rect 19 -8987915 25 -8987518
rect -25 -8987927 25 -8987915
rect -25 -9067949 25 -9067937
rect -25 -9068346 -19 -9067949
rect 19 -9068346 25 -9067949
rect -25 -9068358 25 -9068346
rect -25 -9068486 25 -9068474
rect -25 -9068883 -19 -9068486
rect 19 -9068883 25 -9068486
rect -25 -9068895 25 -9068883
rect -25 -9148917 25 -9148905
rect -25 -9149314 -19 -9148917
rect 19 -9149314 25 -9148917
rect -25 -9149326 25 -9149314
rect -25 -9149454 25 -9149442
rect -25 -9149851 -19 -9149454
rect 19 -9149851 25 -9149454
rect -25 -9149863 25 -9149851
rect -25 -9229885 25 -9229873
rect -25 -9230282 -19 -9229885
rect 19 -9230282 25 -9229885
rect -25 -9230294 25 -9230282
rect -25 -9230422 25 -9230410
rect -25 -9230819 -19 -9230422
rect 19 -9230819 25 -9230422
rect -25 -9230831 25 -9230819
rect -25 -9310853 25 -9310841
rect -25 -9311250 -19 -9310853
rect 19 -9311250 25 -9310853
rect -25 -9311262 25 -9311250
rect -25 -9311390 25 -9311378
rect -25 -9311787 -19 -9311390
rect 19 -9311787 25 -9311390
rect -25 -9311799 25 -9311787
rect -25 -9391821 25 -9391809
rect -25 -9392218 -19 -9391821
rect 19 -9392218 25 -9391821
rect -25 -9392230 25 -9392218
rect -25 -9392358 25 -9392346
rect -25 -9392755 -19 -9392358
rect 19 -9392755 25 -9392358
rect -25 -9392767 25 -9392755
rect -25 -9472789 25 -9472777
rect -25 -9473186 -19 -9472789
rect 19 -9473186 25 -9472789
rect -25 -9473198 25 -9473186
rect -25 -9473326 25 -9473314
rect -25 -9473723 -19 -9473326
rect 19 -9473723 25 -9473326
rect -25 -9473735 25 -9473723
rect -25 -9553757 25 -9553745
rect -25 -9554154 -19 -9553757
rect 19 -9554154 25 -9553757
rect -25 -9554166 25 -9554154
rect -25 -9554294 25 -9554282
rect -25 -9554691 -19 -9554294
rect 19 -9554691 25 -9554294
rect -25 -9554703 25 -9554691
rect -25 -9634725 25 -9634713
rect -25 -9635122 -19 -9634725
rect 19 -9635122 25 -9634725
rect -25 -9635134 25 -9635122
rect -25 -9635262 25 -9635250
rect -25 -9635659 -19 -9635262
rect 19 -9635659 25 -9635262
rect -25 -9635671 25 -9635659
rect -25 -9715693 25 -9715681
rect -25 -9716090 -19 -9715693
rect 19 -9716090 25 -9715693
rect -25 -9716102 25 -9716090
rect -25 -9716230 25 -9716218
rect -25 -9716627 -19 -9716230
rect 19 -9716627 25 -9716230
rect -25 -9716639 25 -9716627
rect -25 -9796661 25 -9796649
rect -25 -9797058 -19 -9796661
rect 19 -9797058 25 -9796661
rect -25 -9797070 25 -9797058
rect -25 -9797198 25 -9797186
rect -25 -9797595 -19 -9797198
rect 19 -9797595 25 -9797198
rect -25 -9797607 25 -9797595
rect -25 -9877629 25 -9877617
rect -25 -9878026 -19 -9877629
rect 19 -9878026 25 -9877629
rect -25 -9878038 25 -9878026
rect -25 -9878166 25 -9878154
rect -25 -9878563 -19 -9878166
rect 19 -9878563 25 -9878166
rect -25 -9878575 25 -9878563
rect -25 -9958597 25 -9958585
rect -25 -9958994 -19 -9958597
rect 19 -9958994 25 -9958597
rect -25 -9959006 25 -9958994
rect -25 -9959134 25 -9959122
rect -25 -9959531 -19 -9959134
rect 19 -9959531 25 -9959134
rect -25 -9959543 25 -9959531
rect -25 -10039565 25 -10039553
rect -25 -10039962 -19 -10039565
rect 19 -10039962 25 -10039565
rect -25 -10039974 25 -10039962
rect -25 -10040102 25 -10040090
rect -25 -10040499 -19 -10040102
rect 19 -10040499 25 -10040102
rect -25 -10040511 25 -10040499
rect -25 -10120533 25 -10120521
rect -25 -10120930 -19 -10120533
rect 19 -10120930 25 -10120533
rect -25 -10120942 25 -10120930
rect -25 -10121070 25 -10121058
rect -25 -10121467 -19 -10121070
rect 19 -10121467 25 -10121070
rect -25 -10121479 25 -10121467
rect -25 -10201501 25 -10201489
rect -25 -10201898 -19 -10201501
rect 19 -10201898 25 -10201501
rect -25 -10201910 25 -10201898
rect -25 -10202038 25 -10202026
rect -25 -10202435 -19 -10202038
rect 19 -10202435 25 -10202038
rect -25 -10202447 25 -10202435
rect -25 -10282469 25 -10282457
rect -25 -10282866 -19 -10282469
rect 19 -10282866 25 -10282469
rect -25 -10282878 25 -10282866
rect -25 -10283006 25 -10282994
rect -25 -10283403 -19 -10283006
rect 19 -10283403 25 -10283006
rect -25 -10283415 25 -10283403
rect -25 -10363437 25 -10363425
rect -25 -10363834 -19 -10363437
rect 19 -10363834 25 -10363437
rect -25 -10363846 25 -10363834
rect -25 -10363974 25 -10363962
rect -25 -10364371 -19 -10363974
rect 19 -10364371 25 -10363974
rect -25 -10364383 25 -10364371
rect -25 -10444405 25 -10444393
rect -25 -10444802 -19 -10444405
rect 19 -10444802 25 -10444405
rect -25 -10444814 25 -10444802
rect -25 -10444942 25 -10444930
rect -25 -10445339 -19 -10444942
rect 19 -10445339 25 -10444942
rect -25 -10445351 25 -10445339
rect -25 -10525373 25 -10525361
rect -25 -10525770 -19 -10525373
rect 19 -10525770 25 -10525373
rect -25 -10525782 25 -10525770
rect -25 -10525910 25 -10525898
rect -25 -10526307 -19 -10525910
rect 19 -10526307 25 -10525910
rect -25 -10526319 25 -10526307
rect -25 -10606341 25 -10606329
rect -25 -10606738 -19 -10606341
rect 19 -10606738 25 -10606341
rect -25 -10606750 25 -10606738
rect -25 -10606878 25 -10606866
rect -25 -10607275 -19 -10606878
rect 19 -10607275 25 -10606878
rect -25 -10607287 25 -10607275
rect -25 -10687309 25 -10687297
rect -25 -10687706 -19 -10687309
rect 19 -10687706 25 -10687309
rect -25 -10687718 25 -10687706
rect -25 -10687846 25 -10687834
rect -25 -10688243 -19 -10687846
rect 19 -10688243 25 -10687846
rect -25 -10688255 25 -10688243
rect -25 -10768277 25 -10768265
rect -25 -10768674 -19 -10768277
rect 19 -10768674 25 -10768277
rect -25 -10768686 25 -10768674
rect -25 -10768814 25 -10768802
rect -25 -10769211 -19 -10768814
rect 19 -10769211 25 -10768814
rect -25 -10769223 25 -10769211
rect -25 -10849245 25 -10849233
rect -25 -10849642 -19 -10849245
rect 19 -10849642 25 -10849245
rect -25 -10849654 25 -10849642
rect -25 -10849782 25 -10849770
rect -25 -10850179 -19 -10849782
rect 19 -10850179 25 -10849782
rect -25 -10850191 25 -10850179
rect -25 -10930213 25 -10930201
rect -25 -10930610 -19 -10930213
rect 19 -10930610 25 -10930213
rect -25 -10930622 25 -10930610
rect -25 -10930750 25 -10930738
rect -25 -10931147 -19 -10930750
rect 19 -10931147 25 -10930750
rect -25 -10931159 25 -10931147
rect -25 -11011181 25 -11011169
rect -25 -11011578 -19 -11011181
rect 19 -11011578 25 -11011181
rect -25 -11011590 25 -11011578
rect -25 -11011718 25 -11011706
rect -25 -11012115 -19 -11011718
rect 19 -11012115 25 -11011718
rect -25 -11012127 25 -11012115
rect -25 -11092149 25 -11092137
rect -25 -11092546 -19 -11092149
rect 19 -11092546 25 -11092149
rect -25 -11092558 25 -11092546
rect -25 -11092686 25 -11092674
rect -25 -11093083 -19 -11092686
rect 19 -11093083 25 -11092686
rect -25 -11093095 25 -11093083
rect -25 -11173117 25 -11173105
rect -25 -11173514 -19 -11173117
rect 19 -11173514 25 -11173117
rect -25 -11173526 25 -11173514
rect -25 -11173654 25 -11173642
rect -25 -11174051 -19 -11173654
rect 19 -11174051 25 -11173654
rect -25 -11174063 25 -11174051
rect -25 -11254085 25 -11254073
rect -25 -11254482 -19 -11254085
rect 19 -11254482 25 -11254085
rect -25 -11254494 25 -11254482
rect -25 -11254622 25 -11254610
rect -25 -11255019 -19 -11254622
rect 19 -11255019 25 -11254622
rect -25 -11255031 25 -11255019
rect -25 -11335053 25 -11335041
rect -25 -11335450 -19 -11335053
rect 19 -11335450 25 -11335053
rect -25 -11335462 25 -11335450
rect -25 -11335590 25 -11335578
rect -25 -11335987 -19 -11335590
rect 19 -11335987 25 -11335590
rect -25 -11335999 25 -11335987
rect -25 -11416021 25 -11416009
rect -25 -11416418 -19 -11416021
rect 19 -11416418 25 -11416021
rect -25 -11416430 25 -11416418
rect -25 -11416558 25 -11416546
rect -25 -11416955 -19 -11416558
rect 19 -11416955 25 -11416558
rect -25 -11416967 25 -11416955
rect -25 -11496989 25 -11496977
rect -25 -11497386 -19 -11496989
rect 19 -11497386 25 -11496989
rect -25 -11497398 25 -11497386
rect -25 -11497526 25 -11497514
rect -25 -11497923 -19 -11497526
rect 19 -11497923 25 -11497526
rect -25 -11497935 25 -11497923
rect -25 -11577957 25 -11577945
rect -25 -11578354 -19 -11577957
rect 19 -11578354 25 -11577957
rect -25 -11578366 25 -11578354
rect -25 -11578494 25 -11578482
rect -25 -11578891 -19 -11578494
rect 19 -11578891 25 -11578494
rect -25 -11578903 25 -11578891
rect -25 -11658925 25 -11658913
rect -25 -11659322 -19 -11658925
rect 19 -11659322 25 -11658925
rect -25 -11659334 25 -11659322
rect -25 -11659462 25 -11659450
rect -25 -11659859 -19 -11659462
rect 19 -11659859 25 -11659462
rect -25 -11659871 25 -11659859
rect -25 -11739893 25 -11739881
rect -25 -11740290 -19 -11739893
rect 19 -11740290 25 -11739893
rect -25 -11740302 25 -11740290
rect -25 -11740430 25 -11740418
rect -25 -11740827 -19 -11740430
rect 19 -11740827 25 -11740430
rect -25 -11740839 25 -11740827
rect -25 -11820861 25 -11820849
rect -25 -11821258 -19 -11820861
rect 19 -11821258 25 -11820861
rect -25 -11821270 25 -11821258
rect -25 -11821398 25 -11821386
rect -25 -11821795 -19 -11821398
rect 19 -11821795 25 -11821398
rect -25 -11821807 25 -11821795
rect -25 -11901829 25 -11901817
rect -25 -11902226 -19 -11901829
rect 19 -11902226 25 -11901829
rect -25 -11902238 25 -11902226
rect -25 -11902366 25 -11902354
rect -25 -11902763 -19 -11902366
rect 19 -11902763 25 -11902366
rect -25 -11902775 25 -11902763
rect -25 -11982797 25 -11982785
rect -25 -11983194 -19 -11982797
rect 19 -11983194 25 -11982797
rect -25 -11983206 25 -11983194
rect -25 -11983334 25 -11983322
rect -25 -11983731 -19 -11983334
rect 19 -11983731 25 -11983334
rect -25 -11983743 25 -11983731
rect -25 -12063765 25 -12063753
rect -25 -12064162 -19 -12063765
rect 19 -12064162 25 -12063765
rect -25 -12064174 25 -12064162
rect -25 -12064302 25 -12064290
rect -25 -12064699 -19 -12064302
rect 19 -12064699 25 -12064302
rect -25 -12064711 25 -12064699
rect -25 -12144733 25 -12144721
rect -25 -12145130 -19 -12144733
rect 19 -12145130 25 -12144733
rect -25 -12145142 25 -12145130
rect -25 -12145270 25 -12145258
rect -25 -12145667 -19 -12145270
rect 19 -12145667 25 -12145270
rect -25 -12145679 25 -12145667
rect -25 -12225701 25 -12225689
rect -25 -12226098 -19 -12225701
rect 19 -12226098 25 -12225701
rect -25 -12226110 25 -12226098
rect -25 -12226238 25 -12226226
rect -25 -12226635 -19 -12226238
rect 19 -12226635 25 -12226238
rect -25 -12226647 25 -12226635
rect -25 -12306669 25 -12306657
rect -25 -12307066 -19 -12306669
rect 19 -12307066 25 -12306669
rect -25 -12307078 25 -12307066
rect -25 -12307206 25 -12307194
rect -25 -12307603 -19 -12307206
rect 19 -12307603 25 -12307206
rect -25 -12307615 25 -12307603
rect -25 -12387637 25 -12387625
rect -25 -12388034 -19 -12387637
rect 19 -12388034 25 -12387637
rect -25 -12388046 25 -12388034
rect -25 -12388174 25 -12388162
rect -25 -12388571 -19 -12388174
rect 19 -12388571 25 -12388174
rect -25 -12388583 25 -12388571
rect -25 -12468605 25 -12468593
rect -25 -12469002 -19 -12468605
rect 19 -12469002 25 -12468605
rect -25 -12469014 25 -12469002
rect -25 -12469142 25 -12469130
rect -25 -12469539 -19 -12469142
rect 19 -12469539 25 -12469142
rect -25 -12469551 25 -12469539
rect -25 -12549573 25 -12549561
rect -25 -12549970 -19 -12549573
rect 19 -12549970 25 -12549573
rect -25 -12549982 25 -12549970
rect -25 -12550110 25 -12550098
rect -25 -12550507 -19 -12550110
rect 19 -12550507 25 -12550110
rect -25 -12550519 25 -12550507
rect -25 -12630541 25 -12630529
rect -25 -12630938 -19 -12630541
rect 19 -12630938 25 -12630541
rect -25 -12630950 25 -12630938
rect -25 -12631078 25 -12631066
rect -25 -12631475 -19 -12631078
rect 19 -12631475 25 -12631078
rect -25 -12631487 25 -12631475
rect -25 -12711509 25 -12711497
rect -25 -12711906 -19 -12711509
rect 19 -12711906 25 -12711509
rect -25 -12711918 25 -12711906
rect -25 -12712046 25 -12712034
rect -25 -12712443 -19 -12712046
rect 19 -12712443 25 -12712046
rect -25 -12712455 25 -12712443
rect -25 -12792477 25 -12792465
rect -25 -12792874 -19 -12792477
rect 19 -12792874 25 -12792477
rect -25 -12792886 25 -12792874
rect -25 -12793014 25 -12793002
rect -25 -12793411 -19 -12793014
rect 19 -12793411 25 -12793014
rect -25 -12793423 25 -12793411
rect -25 -12873445 25 -12873433
rect -25 -12873842 -19 -12873445
rect 19 -12873842 25 -12873445
rect -25 -12873854 25 -12873842
rect -25 -12873982 25 -12873970
rect -25 -12874379 -19 -12873982
rect 19 -12874379 25 -12873982
rect -25 -12874391 25 -12874379
rect -25 -12954413 25 -12954401
rect -25 -12954810 -19 -12954413
rect 19 -12954810 25 -12954413
rect -25 -12954822 25 -12954810
rect -25 -12954950 25 -12954938
rect -25 -12955347 -19 -12954950
rect 19 -12955347 25 -12954950
rect -25 -12955359 25 -12955347
rect -25 -13035381 25 -13035369
rect -25 -13035778 -19 -13035381
rect 19 -13035778 25 -13035381
rect -25 -13035790 25 -13035778
rect -25 -13035918 25 -13035906
rect -25 -13036315 -19 -13035918
rect 19 -13036315 25 -13035918
rect -25 -13036327 25 -13036315
rect -25 -13116349 25 -13116337
rect -25 -13116746 -19 -13116349
rect 19 -13116746 25 -13116349
rect -25 -13116758 25 -13116746
rect -25 -13116886 25 -13116874
rect -25 -13117283 -19 -13116886
rect 19 -13117283 25 -13116886
rect -25 -13117295 25 -13117283
rect -25 -13197317 25 -13197305
rect -25 -13197714 -19 -13197317
rect 19 -13197714 25 -13197317
rect -25 -13197726 25 -13197714
rect -25 -13197854 25 -13197842
rect -25 -13198251 -19 -13197854
rect 19 -13198251 25 -13197854
rect -25 -13198263 25 -13198251
rect -25 -13278285 25 -13278273
rect -25 -13278682 -19 -13278285
rect 19 -13278682 25 -13278285
rect -25 -13278694 25 -13278682
rect -25 -13278822 25 -13278810
rect -25 -13279219 -19 -13278822
rect 19 -13279219 25 -13278822
rect -25 -13279231 25 -13279219
rect -25 -13359253 25 -13359241
rect -25 -13359650 -19 -13359253
rect 19 -13359650 25 -13359253
rect -25 -13359662 25 -13359650
rect -25 -13359790 25 -13359778
rect -25 -13360187 -19 -13359790
rect 19 -13360187 25 -13359790
rect -25 -13360199 25 -13360187
rect -25 -13440221 25 -13440209
rect -25 -13440618 -19 -13440221
rect 19 -13440618 25 -13440221
rect -25 -13440630 25 -13440618
rect -25 -13440758 25 -13440746
rect -25 -13441155 -19 -13440758
rect 19 -13441155 25 -13440758
rect -25 -13441167 25 -13441155
rect -25 -13521189 25 -13521177
rect -25 -13521586 -19 -13521189
rect 19 -13521586 25 -13521189
rect -25 -13521598 25 -13521586
rect -25 -13521726 25 -13521714
rect -25 -13522123 -19 -13521726
rect 19 -13522123 25 -13521726
rect -25 -13522135 25 -13522123
rect -25 -13602157 25 -13602145
rect -25 -13602554 -19 -13602157
rect 19 -13602554 25 -13602157
rect -25 -13602566 25 -13602554
rect -25 -13602694 25 -13602682
rect -25 -13603091 -19 -13602694
rect 19 -13603091 25 -13602694
rect -25 -13603103 25 -13603091
rect -25 -13683125 25 -13683113
rect -25 -13683522 -19 -13683125
rect 19 -13683522 25 -13683125
rect -25 -13683534 25 -13683522
rect -25 -13683662 25 -13683650
rect -25 -13684059 -19 -13683662
rect 19 -13684059 25 -13683662
rect -25 -13684071 25 -13684059
rect -25 -13764093 25 -13764081
rect -25 -13764490 -19 -13764093
rect 19 -13764490 25 -13764093
rect -25 -13764502 25 -13764490
rect -25 -13764630 25 -13764618
rect -25 -13765027 -19 -13764630
rect 19 -13765027 25 -13764630
rect -25 -13765039 25 -13765027
rect -25 -13845061 25 -13845049
rect -25 -13845458 -19 -13845061
rect 19 -13845458 25 -13845061
rect -25 -13845470 25 -13845458
rect -25 -13845598 25 -13845586
rect -25 -13845995 -19 -13845598
rect 19 -13845995 25 -13845598
rect -25 -13846007 25 -13845995
rect -25 -13926029 25 -13926017
rect -25 -13926426 -19 -13926029
rect 19 -13926426 25 -13926029
rect -25 -13926438 25 -13926426
rect -25 -13926566 25 -13926554
rect -25 -13926963 -19 -13926566
rect 19 -13926963 25 -13926566
rect -25 -13926975 25 -13926963
rect -25 -14006997 25 -14006985
rect -25 -14007394 -19 -14006997
rect 19 -14007394 25 -14006997
rect -25 -14007406 25 -14007394
rect -25 -14007534 25 -14007522
rect -25 -14007931 -19 -14007534
rect 19 -14007931 25 -14007534
rect -25 -14007943 25 -14007931
rect -25 -14087965 25 -14087953
rect -25 -14088362 -19 -14087965
rect 19 -14088362 25 -14087965
rect -25 -14088374 25 -14088362
rect -25 -14088502 25 -14088490
rect -25 -14088899 -19 -14088502
rect 19 -14088899 25 -14088502
rect -25 -14088911 25 -14088899
rect -25 -14168933 25 -14168921
rect -25 -14169330 -19 -14168933
rect 19 -14169330 25 -14168933
rect -25 -14169342 25 -14169330
rect -25 -14169470 25 -14169458
rect -25 -14169867 -19 -14169470
rect 19 -14169867 25 -14169470
rect -25 -14169879 25 -14169867
rect -25 -14249901 25 -14249889
rect -25 -14250298 -19 -14249901
rect 19 -14250298 25 -14249901
rect -25 -14250310 25 -14250298
rect -25 -14250438 25 -14250426
rect -25 -14250835 -19 -14250438
rect 19 -14250835 25 -14250438
rect -25 -14250847 25 -14250835
rect -25 -14330869 25 -14330857
rect -25 -14331266 -19 -14330869
rect 19 -14331266 25 -14330869
rect -25 -14331278 25 -14331266
rect -25 -14331406 25 -14331394
rect -25 -14331803 -19 -14331406
rect 19 -14331803 25 -14331406
rect -25 -14331815 25 -14331803
rect -25 -14411837 25 -14411825
rect -25 -14412234 -19 -14411837
rect 19 -14412234 25 -14411837
rect -25 -14412246 25 -14412234
rect -25 -14412374 25 -14412362
rect -25 -14412771 -19 -14412374
rect 19 -14412771 25 -14412374
rect -25 -14412783 25 -14412771
rect -25 -14492805 25 -14492793
rect -25 -14493202 -19 -14492805
rect 19 -14493202 25 -14492805
rect -25 -14493214 25 -14493202
rect -25 -14493342 25 -14493330
rect -25 -14493739 -19 -14493342
rect 19 -14493739 25 -14493342
rect -25 -14493751 25 -14493739
rect -25 -14573773 25 -14573761
rect -25 -14574170 -19 -14573773
rect 19 -14574170 25 -14573773
rect -25 -14574182 25 -14574170
rect -25 -14574310 25 -14574298
rect -25 -14574707 -19 -14574310
rect 19 -14574707 25 -14574310
rect -25 -14574719 25 -14574707
rect -25 -14654741 25 -14654729
rect -25 -14655138 -19 -14654741
rect 19 -14655138 25 -14654741
rect -25 -14655150 25 -14655138
rect -25 -14655278 25 -14655266
rect -25 -14655675 -19 -14655278
rect 19 -14655675 25 -14655278
rect -25 -14655687 25 -14655675
rect -25 -14735709 25 -14735697
rect -25 -14736106 -19 -14735709
rect 19 -14736106 25 -14735709
rect -25 -14736118 25 -14736106
rect -25 -14736246 25 -14736234
rect -25 -14736643 -19 -14736246
rect 19 -14736643 25 -14736246
rect -25 -14736655 25 -14736643
rect -25 -14816677 25 -14816665
rect -25 -14817074 -19 -14816677
rect 19 -14817074 25 -14816677
rect -25 -14817086 25 -14817074
rect -25 -14817214 25 -14817202
rect -25 -14817611 -19 -14817214
rect 19 -14817611 25 -14817214
rect -25 -14817623 25 -14817611
rect -25 -14897645 25 -14897633
rect -25 -14898042 -19 -14897645
rect 19 -14898042 25 -14897645
rect -25 -14898054 25 -14898042
rect -25 -14898182 25 -14898170
rect -25 -14898579 -19 -14898182
rect 19 -14898579 25 -14898182
rect -25 -14898591 25 -14898579
rect -25 -14978613 25 -14978601
rect -25 -14979010 -19 -14978613
rect 19 -14979010 25 -14978613
rect -25 -14979022 25 -14979010
rect -25 -14979150 25 -14979138
rect -25 -14979547 -19 -14979150
rect 19 -14979547 25 -14979150
rect -25 -14979559 25 -14979547
rect -25 -15059581 25 -15059569
rect -25 -15059978 -19 -15059581
rect 19 -15059978 25 -15059581
rect -25 -15059990 25 -15059978
rect -25 -15060118 25 -15060106
rect -25 -15060515 -19 -15060118
rect 19 -15060515 25 -15060118
rect -25 -15060527 25 -15060515
rect -25 -15140549 25 -15140537
rect -25 -15140946 -19 -15140549
rect 19 -15140946 25 -15140549
rect -25 -15140958 25 -15140946
rect -25 -15141086 25 -15141074
rect -25 -15141483 -19 -15141086
rect 19 -15141483 25 -15141086
rect -25 -15141495 25 -15141483
rect -25 -15221517 25 -15221505
rect -25 -15221914 -19 -15221517
rect 19 -15221914 25 -15221517
rect -25 -15221926 25 -15221914
rect -25 -15222054 25 -15222042
rect -25 -15222451 -19 -15222054
rect 19 -15222451 25 -15222054
rect -25 -15222463 25 -15222451
rect -25 -15302485 25 -15302473
rect -25 -15302882 -19 -15302485
rect 19 -15302882 25 -15302485
rect -25 -15302894 25 -15302882
rect -25 -15303022 25 -15303010
rect -25 -15303419 -19 -15303022
rect 19 -15303419 25 -15303022
rect -25 -15303431 25 -15303419
rect -25 -15383453 25 -15383441
rect -25 -15383850 -19 -15383453
rect 19 -15383850 25 -15383453
rect -25 -15383862 25 -15383850
rect -25 -15383990 25 -15383978
rect -25 -15384387 -19 -15383990
rect 19 -15384387 25 -15383990
rect -25 -15384399 25 -15384387
rect -25 -15464421 25 -15464409
rect -25 -15464818 -19 -15464421
rect 19 -15464818 25 -15464421
rect -25 -15464830 25 -15464818
rect -25 -15464958 25 -15464946
rect -25 -15465355 -19 -15464958
rect 19 -15465355 25 -15464958
rect -25 -15465367 25 -15465355
rect -25 -15545389 25 -15545377
rect -25 -15545786 -19 -15545389
rect 19 -15545786 25 -15545389
rect -25 -15545798 25 -15545786
rect -25 -15545926 25 -15545914
rect -25 -15546323 -19 -15545926
rect 19 -15546323 25 -15545926
rect -25 -15546335 25 -15546323
rect -25 -15626357 25 -15626345
rect -25 -15626754 -19 -15626357
rect 19 -15626754 25 -15626357
rect -25 -15626766 25 -15626754
rect -25 -15626894 25 -15626882
rect -25 -15627291 -19 -15626894
rect 19 -15627291 25 -15626894
rect -25 -15627303 25 -15627291
rect -25 -15707325 25 -15707313
rect -25 -15707722 -19 -15707325
rect 19 -15707722 25 -15707325
rect -25 -15707734 25 -15707722
rect -25 -15707862 25 -15707850
rect -25 -15708259 -19 -15707862
rect 19 -15708259 25 -15707862
rect -25 -15708271 25 -15708259
rect -25 -15788293 25 -15788281
rect -25 -15788690 -19 -15788293
rect 19 -15788690 25 -15788293
rect -25 -15788702 25 -15788690
rect -25 -15788830 25 -15788818
rect -25 -15789227 -19 -15788830
rect 19 -15789227 25 -15788830
rect -25 -15789239 25 -15789227
rect -25 -15869261 25 -15869249
rect -25 -15869658 -19 -15869261
rect 19 -15869658 25 -15869261
rect -25 -15869670 25 -15869658
rect -25 -15869798 25 -15869786
rect -25 -15870195 -19 -15869798
rect 19 -15870195 25 -15869798
rect -25 -15870207 25 -15870195
rect -25 -15950229 25 -15950217
rect -25 -15950626 -19 -15950229
rect 19 -15950626 25 -15950229
rect -25 -15950638 25 -15950626
rect -25 -15950766 25 -15950754
rect -25 -15951163 -19 -15950766
rect 19 -15951163 25 -15950766
rect -25 -15951175 25 -15951163
rect -25 -16031197 25 -16031185
rect -25 -16031594 -19 -16031197
rect 19 -16031594 25 -16031197
rect -25 -16031606 25 -16031594
rect -25 -16031734 25 -16031722
rect -25 -16032131 -19 -16031734
rect 19 -16032131 25 -16031734
rect -25 -16032143 25 -16032131
rect -25 -16112165 25 -16112153
rect -25 -16112562 -19 -16112165
rect 19 -16112562 25 -16112165
rect -25 -16112574 25 -16112562
rect -25 -16112702 25 -16112690
rect -25 -16113099 -19 -16112702
rect 19 -16113099 25 -16112702
rect -25 -16113111 25 -16113099
rect -25 -16193133 25 -16193121
rect -25 -16193530 -19 -16193133
rect 19 -16193530 25 -16193133
rect -25 -16193542 25 -16193530
rect -25 -16193670 25 -16193658
rect -25 -16194067 -19 -16193670
rect 19 -16194067 25 -16193670
rect -25 -16194079 25 -16194067
rect -25 -16274101 25 -16274089
rect -25 -16274498 -19 -16274101
rect 19 -16274498 25 -16274101
rect -25 -16274510 25 -16274498
rect -25 -16274638 25 -16274626
rect -25 -16275035 -19 -16274638
rect 19 -16275035 25 -16274638
rect -25 -16275047 25 -16275035
rect -25 -16355069 25 -16355057
rect -25 -16355466 -19 -16355069
rect 19 -16355466 25 -16355069
rect -25 -16355478 25 -16355466
rect -25 -16355606 25 -16355594
rect -25 -16356003 -19 -16355606
rect 19 -16356003 25 -16355606
rect -25 -16356015 25 -16356003
rect -25 -16436037 25 -16436025
rect -25 -16436434 -19 -16436037
rect 19 -16436434 25 -16436037
rect -25 -16436446 25 -16436434
rect -25 -16436574 25 -16436562
rect -25 -16436971 -19 -16436574
rect 19 -16436971 25 -16436574
rect -25 -16436983 25 -16436971
rect -25 -16517005 25 -16516993
rect -25 -16517402 -19 -16517005
rect 19 -16517402 25 -16517005
rect -25 -16517414 25 -16517402
rect -25 -16517542 25 -16517530
rect -25 -16517939 -19 -16517542
rect 19 -16517939 25 -16517542
rect -25 -16517951 25 -16517939
rect -25 -16597973 25 -16597961
rect -25 -16598370 -19 -16597973
rect 19 -16598370 25 -16597973
rect -25 -16598382 25 -16598370
rect -25 -16598510 25 -16598498
rect -25 -16598907 -19 -16598510
rect 19 -16598907 25 -16598510
rect -25 -16598919 25 -16598907
rect -25 -16678941 25 -16678929
rect -25 -16679338 -19 -16678941
rect 19 -16679338 25 -16678941
rect -25 -16679350 25 -16679338
rect -25 -16679478 25 -16679466
rect -25 -16679875 -19 -16679478
rect 19 -16679875 25 -16679478
rect -25 -16679887 25 -16679875
rect -25 -16759909 25 -16759897
rect -25 -16760306 -19 -16759909
rect 19 -16760306 25 -16759909
rect -25 -16760318 25 -16760306
rect -25 -16760446 25 -16760434
rect -25 -16760843 -19 -16760446
rect 19 -16760843 25 -16760446
rect -25 -16760855 25 -16760843
rect -25 -16840877 25 -16840865
rect -25 -16841274 -19 -16840877
rect 19 -16841274 25 -16840877
rect -25 -16841286 25 -16841274
rect -25 -16841414 25 -16841402
rect -25 -16841811 -19 -16841414
rect 19 -16841811 25 -16841414
rect -25 -16841823 25 -16841811
rect -25 -16921845 25 -16921833
rect -25 -16922242 -19 -16921845
rect 19 -16922242 25 -16921845
rect -25 -16922254 25 -16922242
rect -25 -16922382 25 -16922370
rect -25 -16922779 -19 -16922382
rect 19 -16922779 25 -16922382
rect -25 -16922791 25 -16922779
rect -25 -17002813 25 -17002801
rect -25 -17003210 -19 -17002813
rect 19 -17003210 25 -17002813
rect -25 -17003222 25 -17003210
rect -25 -17003350 25 -17003338
rect -25 -17003747 -19 -17003350
rect 19 -17003747 25 -17003350
rect -25 -17003759 25 -17003747
rect -25 -17083781 25 -17083769
rect -25 -17084178 -19 -17083781
rect 19 -17084178 25 -17083781
rect -25 -17084190 25 -17084178
rect -25 -17084318 25 -17084306
rect -25 -17084715 -19 -17084318
rect 19 -17084715 25 -17084318
rect -25 -17084727 25 -17084715
rect -25 -17164749 25 -17164737
rect -25 -17165146 -19 -17164749
rect 19 -17165146 25 -17164749
rect -25 -17165158 25 -17165146
rect -25 -17165286 25 -17165274
rect -25 -17165683 -19 -17165286
rect 19 -17165683 25 -17165286
rect -25 -17165695 25 -17165683
rect -25 -17245717 25 -17245705
rect -25 -17246114 -19 -17245717
rect 19 -17246114 25 -17245717
rect -25 -17246126 25 -17246114
rect -25 -17246254 25 -17246242
rect -25 -17246651 -19 -17246254
rect 19 -17246651 25 -17246254
rect -25 -17246663 25 -17246651
rect -25 -17326685 25 -17326673
rect -25 -17327082 -19 -17326685
rect 19 -17327082 25 -17326685
rect -25 -17327094 25 -17327082
rect -25 -17327222 25 -17327210
rect -25 -17327619 -19 -17327222
rect 19 -17327619 25 -17327222
rect -25 -17327631 25 -17327619
rect -25 -17407653 25 -17407641
rect -25 -17408050 -19 -17407653
rect 19 -17408050 25 -17407653
rect -25 -17408062 25 -17408050
rect -25 -17408190 25 -17408178
rect -25 -17408587 -19 -17408190
rect 19 -17408587 25 -17408190
rect -25 -17408599 25 -17408587
rect -25 -17488621 25 -17488609
rect -25 -17489018 -19 -17488621
rect 19 -17489018 25 -17488621
rect -25 -17489030 25 -17489018
rect -25 -17489158 25 -17489146
rect -25 -17489555 -19 -17489158
rect 19 -17489555 25 -17489158
rect -25 -17489567 25 -17489555
rect -25 -17569589 25 -17569577
rect -25 -17569986 -19 -17569589
rect 19 -17569986 25 -17569589
rect -25 -17569998 25 -17569986
rect -25 -17570126 25 -17570114
rect -25 -17570523 -19 -17570126
rect 19 -17570523 25 -17570126
rect -25 -17570535 25 -17570523
rect -25 -17650557 25 -17650545
rect -25 -17650954 -19 -17650557
rect 19 -17650954 25 -17650557
rect -25 -17650966 25 -17650954
rect -25 -17651094 25 -17651082
rect -25 -17651491 -19 -17651094
rect 19 -17651491 25 -17651094
rect -25 -17651503 25 -17651491
rect -25 -17731525 25 -17731513
rect -25 -17731922 -19 -17731525
rect 19 -17731922 25 -17731525
rect -25 -17731934 25 -17731922
rect -25 -17732062 25 -17732050
rect -25 -17732459 -19 -17732062
rect 19 -17732459 25 -17732062
rect -25 -17732471 25 -17732459
rect -25 -17812493 25 -17812481
rect -25 -17812890 -19 -17812493
rect 19 -17812890 25 -17812493
rect -25 -17812902 25 -17812890
rect -25 -17813030 25 -17813018
rect -25 -17813427 -19 -17813030
rect 19 -17813427 25 -17813030
rect -25 -17813439 25 -17813427
rect -25 -17893461 25 -17893449
rect -25 -17893858 -19 -17893461
rect 19 -17893858 25 -17893461
rect -25 -17893870 25 -17893858
rect -25 -17893998 25 -17893986
rect -25 -17894395 -19 -17893998
rect 19 -17894395 25 -17893998
rect -25 -17894407 25 -17894395
rect -25 -17974429 25 -17974417
rect -25 -17974826 -19 -17974429
rect 19 -17974826 25 -17974429
rect -25 -17974838 25 -17974826
rect -25 -17974966 25 -17974954
rect -25 -17975363 -19 -17974966
rect 19 -17975363 25 -17974966
rect -25 -17975375 25 -17975363
rect -25 -18055397 25 -18055385
rect -25 -18055794 -19 -18055397
rect 19 -18055794 25 -18055397
rect -25 -18055806 25 -18055794
rect -25 -18055934 25 -18055922
rect -25 -18056331 -19 -18055934
rect 19 -18056331 25 -18055934
rect -25 -18056343 25 -18056331
rect -25 -18136365 25 -18136353
rect -25 -18136762 -19 -18136365
rect 19 -18136762 25 -18136365
rect -25 -18136774 25 -18136762
rect -25 -18136902 25 -18136890
rect -25 -18137299 -19 -18136902
rect 19 -18137299 25 -18136902
rect -25 -18137311 25 -18137299
rect -25 -18217333 25 -18217321
rect -25 -18217730 -19 -18217333
rect 19 -18217730 25 -18217333
rect -25 -18217742 25 -18217730
rect -25 -18217870 25 -18217858
rect -25 -18218267 -19 -18217870
rect 19 -18218267 25 -18217870
rect -25 -18218279 25 -18218267
rect -25 -18298301 25 -18298289
rect -25 -18298698 -19 -18298301
rect 19 -18298698 25 -18298301
rect -25 -18298710 25 -18298698
rect -25 -18298838 25 -18298826
rect -25 -18299235 -19 -18298838
rect 19 -18299235 25 -18298838
rect -25 -18299247 25 -18299235
rect -25 -18379269 25 -18379257
rect -25 -18379666 -19 -18379269
rect 19 -18379666 25 -18379269
rect -25 -18379678 25 -18379666
rect -25 -18379806 25 -18379794
rect -25 -18380203 -19 -18379806
rect 19 -18380203 25 -18379806
rect -25 -18380215 25 -18380203
rect -25 -18460237 25 -18460225
rect -25 -18460634 -19 -18460237
rect 19 -18460634 25 -18460237
rect -25 -18460646 25 -18460634
rect -25 -18460774 25 -18460762
rect -25 -18461171 -19 -18460774
rect 19 -18461171 25 -18460774
rect -25 -18461183 25 -18461171
rect -25 -18541205 25 -18541193
rect -25 -18541602 -19 -18541205
rect 19 -18541602 25 -18541205
rect -25 -18541614 25 -18541602
rect -25 -18541742 25 -18541730
rect -25 -18542139 -19 -18541742
rect 19 -18542139 25 -18541742
rect -25 -18542151 25 -18542139
rect -25 -18622173 25 -18622161
rect -25 -18622570 -19 -18622173
rect 19 -18622570 25 -18622173
rect -25 -18622582 25 -18622570
rect -25 -18622710 25 -18622698
rect -25 -18623107 -19 -18622710
rect 19 -18623107 25 -18622710
rect -25 -18623119 25 -18623107
rect -25 -18703141 25 -18703129
rect -25 -18703538 -19 -18703141
rect 19 -18703538 25 -18703141
rect -25 -18703550 25 -18703538
rect -25 -18703678 25 -18703666
rect -25 -18704075 -19 -18703678
rect 19 -18704075 25 -18703678
rect -25 -18704087 25 -18704075
rect -25 -18784109 25 -18784097
rect -25 -18784506 -19 -18784109
rect 19 -18784506 25 -18784109
rect -25 -18784518 25 -18784506
rect -25 -18784646 25 -18784634
rect -25 -18785043 -19 -18784646
rect 19 -18785043 25 -18784646
rect -25 -18785055 25 -18785043
rect -25 -18865077 25 -18865065
rect -25 -18865474 -19 -18865077
rect 19 -18865474 25 -18865077
rect -25 -18865486 25 -18865474
rect -25 -18865614 25 -18865602
rect -25 -18866011 -19 -18865614
rect 19 -18866011 25 -18865614
rect -25 -18866023 25 -18866011
rect -25 -18946045 25 -18946033
rect -25 -18946442 -19 -18946045
rect 19 -18946442 25 -18946045
rect -25 -18946454 25 -18946442
rect -25 -18946582 25 -18946570
rect -25 -18946979 -19 -18946582
rect 19 -18946979 25 -18946582
rect -25 -18946991 25 -18946979
rect -25 -19027013 25 -19027001
rect -25 -19027410 -19 -19027013
rect 19 -19027410 25 -19027013
rect -25 -19027422 25 -19027410
rect -25 -19027550 25 -19027538
rect -25 -19027947 -19 -19027550
rect 19 -19027947 25 -19027550
rect -25 -19027959 25 -19027947
rect -25 -19107981 25 -19107969
rect -25 -19108378 -19 -19107981
rect 19 -19108378 25 -19107981
rect -25 -19108390 25 -19108378
rect -25 -19108518 25 -19108506
rect -25 -19108915 -19 -19108518
rect 19 -19108915 25 -19108518
rect -25 -19108927 25 -19108915
rect -25 -19188949 25 -19188937
rect -25 -19189346 -19 -19188949
rect 19 -19189346 25 -19188949
rect -25 -19189358 25 -19189346
rect -25 -19189486 25 -19189474
rect -25 -19189883 -19 -19189486
rect 19 -19189883 25 -19189486
rect -25 -19189895 25 -19189883
rect -25 -19269917 25 -19269905
rect -25 -19270314 -19 -19269917
rect 19 -19270314 25 -19269917
rect -25 -19270326 25 -19270314
rect -25 -19270454 25 -19270442
rect -25 -19270851 -19 -19270454
rect 19 -19270851 25 -19270454
rect -25 -19270863 25 -19270851
rect -25 -19350885 25 -19350873
rect -25 -19351282 -19 -19350885
rect 19 -19351282 25 -19350885
rect -25 -19351294 25 -19351282
rect -25 -19351422 25 -19351410
rect -25 -19351819 -19 -19351422
rect 19 -19351819 25 -19351422
rect -25 -19351831 25 -19351819
rect -25 -19431853 25 -19431841
rect -25 -19432250 -19 -19431853
rect 19 -19432250 25 -19431853
rect -25 -19432262 25 -19432250
rect -25 -19432390 25 -19432378
rect -25 -19432787 -19 -19432390
rect 19 -19432787 25 -19432390
rect -25 -19432799 25 -19432787
rect -25 -19512821 25 -19512809
rect -25 -19513218 -19 -19512821
rect 19 -19513218 25 -19512821
rect -25 -19513230 25 -19513218
rect -25 -19513358 25 -19513346
rect -25 -19513755 -19 -19513358
rect 19 -19513755 25 -19513358
rect -25 -19513767 25 -19513755
rect -25 -19593789 25 -19593777
rect -25 -19594186 -19 -19593789
rect 19 -19594186 25 -19593789
rect -25 -19594198 25 -19594186
rect -25 -19594326 25 -19594314
rect -25 -19594723 -19 -19594326
rect 19 -19594723 25 -19594326
rect -25 -19594735 25 -19594723
rect -25 -19674757 25 -19674745
rect -25 -19675154 -19 -19674757
rect 19 -19675154 25 -19674757
rect -25 -19675166 25 -19675154
rect -25 -19675294 25 -19675282
rect -25 -19675691 -19 -19675294
rect 19 -19675691 25 -19675294
rect -25 -19675703 25 -19675691
rect -25 -19755725 25 -19755713
rect -25 -19756122 -19 -19755725
rect 19 -19756122 25 -19755725
rect -25 -19756134 25 -19756122
rect -25 -19756262 25 -19756250
rect -25 -19756659 -19 -19756262
rect 19 -19756659 25 -19756262
rect -25 -19756671 25 -19756659
rect -25 -19836693 25 -19836681
rect -25 -19837090 -19 -19836693
rect 19 -19837090 25 -19836693
rect -25 -19837102 25 -19837090
rect -25 -19837230 25 -19837218
rect -25 -19837627 -19 -19837230
rect 19 -19837627 25 -19837230
rect -25 -19837639 25 -19837627
rect -25 -19917661 25 -19917649
rect -25 -19918058 -19 -19917661
rect 19 -19918058 25 -19917661
rect -25 -19918070 25 -19918058
rect -25 -19918198 25 -19918186
rect -25 -19918595 -19 -19918198
rect 19 -19918595 25 -19918198
rect -25 -19918607 25 -19918595
rect -25 -19998629 25 -19998617
rect -25 -19999026 -19 -19998629
rect 19 -19999026 25 -19998629
rect -25 -19999038 25 -19999026
rect -25 -19999166 25 -19999154
rect -25 -19999563 -19 -19999166
rect 19 -19999563 25 -19999166
rect -25 -19999575 25 -19999563
rect -25 -20079597 25 -20079585
rect -25 -20079994 -19 -20079597
rect 19 -20079994 25 -20079597
rect -25 -20080006 25 -20079994
rect -25 -20080134 25 -20080122
rect -25 -20080531 -19 -20080134
rect 19 -20080531 25 -20080134
rect -25 -20080543 25 -20080531
rect -25 -20160565 25 -20160553
rect -25 -20160962 -19 -20160565
rect 19 -20160962 25 -20160565
rect -25 -20160974 25 -20160962
rect -25 -20161102 25 -20161090
rect -25 -20161499 -19 -20161102
rect 19 -20161499 25 -20161102
rect -25 -20161511 25 -20161499
rect -25 -20241533 25 -20241521
rect -25 -20241930 -19 -20241533
rect 19 -20241930 25 -20241533
rect -25 -20241942 25 -20241930
<< res0p35 >>
rect -37 20161514 37 20241518
rect -37 20080546 37 20160550
rect -37 19999578 37 20079582
rect -37 19918610 37 19998614
rect -37 19837642 37 19917646
rect -37 19756674 37 19836678
rect -37 19675706 37 19755710
rect -37 19594738 37 19674742
rect -37 19513770 37 19593774
rect -37 19432802 37 19512806
rect -37 19351834 37 19431838
rect -37 19270866 37 19350870
rect -37 19189898 37 19269902
rect -37 19108930 37 19188934
rect -37 19027962 37 19107966
rect -37 18946994 37 19026998
rect -37 18866026 37 18946030
rect -37 18785058 37 18865062
rect -37 18704090 37 18784094
rect -37 18623122 37 18703126
rect -37 18542154 37 18622158
rect -37 18461186 37 18541190
rect -37 18380218 37 18460222
rect -37 18299250 37 18379254
rect -37 18218282 37 18298286
rect -37 18137314 37 18217318
rect -37 18056346 37 18136350
rect -37 17975378 37 18055382
rect -37 17894410 37 17974414
rect -37 17813442 37 17893446
rect -37 17732474 37 17812478
rect -37 17651506 37 17731510
rect -37 17570538 37 17650542
rect -37 17489570 37 17569574
rect -37 17408602 37 17488606
rect -37 17327634 37 17407638
rect -37 17246666 37 17326670
rect -37 17165698 37 17245702
rect -37 17084730 37 17164734
rect -37 17003762 37 17083766
rect -37 16922794 37 17002798
rect -37 16841826 37 16921830
rect -37 16760858 37 16840862
rect -37 16679890 37 16759894
rect -37 16598922 37 16678926
rect -37 16517954 37 16597958
rect -37 16436986 37 16516990
rect -37 16356018 37 16436022
rect -37 16275050 37 16355054
rect -37 16194082 37 16274086
rect -37 16113114 37 16193118
rect -37 16032146 37 16112150
rect -37 15951178 37 16031182
rect -37 15870210 37 15950214
rect -37 15789242 37 15869246
rect -37 15708274 37 15788278
rect -37 15627306 37 15707310
rect -37 15546338 37 15626342
rect -37 15465370 37 15545374
rect -37 15384402 37 15464406
rect -37 15303434 37 15383438
rect -37 15222466 37 15302470
rect -37 15141498 37 15221502
rect -37 15060530 37 15140534
rect -37 14979562 37 15059566
rect -37 14898594 37 14978598
rect -37 14817626 37 14897630
rect -37 14736658 37 14816662
rect -37 14655690 37 14735694
rect -37 14574722 37 14654726
rect -37 14493754 37 14573758
rect -37 14412786 37 14492790
rect -37 14331818 37 14411822
rect -37 14250850 37 14330854
rect -37 14169882 37 14249886
rect -37 14088914 37 14168918
rect -37 14007946 37 14087950
rect -37 13926978 37 14006982
rect -37 13846010 37 13926014
rect -37 13765042 37 13845046
rect -37 13684074 37 13764078
rect -37 13603106 37 13683110
rect -37 13522138 37 13602142
rect -37 13441170 37 13521174
rect -37 13360202 37 13440206
rect -37 13279234 37 13359238
rect -37 13198266 37 13278270
rect -37 13117298 37 13197302
rect -37 13036330 37 13116334
rect -37 12955362 37 13035366
rect -37 12874394 37 12954398
rect -37 12793426 37 12873430
rect -37 12712458 37 12792462
rect -37 12631490 37 12711494
rect -37 12550522 37 12630526
rect -37 12469554 37 12549558
rect -37 12388586 37 12468590
rect -37 12307618 37 12387622
rect -37 12226650 37 12306654
rect -37 12145682 37 12225686
rect -37 12064714 37 12144718
rect -37 11983746 37 12063750
rect -37 11902778 37 11982782
rect -37 11821810 37 11901814
rect -37 11740842 37 11820846
rect -37 11659874 37 11739878
rect -37 11578906 37 11658910
rect -37 11497938 37 11577942
rect -37 11416970 37 11496974
rect -37 11336002 37 11416006
rect -37 11255034 37 11335038
rect -37 11174066 37 11254070
rect -37 11093098 37 11173102
rect -37 11012130 37 11092134
rect -37 10931162 37 11011166
rect -37 10850194 37 10930198
rect -37 10769226 37 10849230
rect -37 10688258 37 10768262
rect -37 10607290 37 10687294
rect -37 10526322 37 10606326
rect -37 10445354 37 10525358
rect -37 10364386 37 10444390
rect -37 10283418 37 10363422
rect -37 10202450 37 10282454
rect -37 10121482 37 10201486
rect -37 10040514 37 10120518
rect -37 9959546 37 10039550
rect -37 9878578 37 9958582
rect -37 9797610 37 9877614
rect -37 9716642 37 9796646
rect -37 9635674 37 9715678
rect -37 9554706 37 9634710
rect -37 9473738 37 9553742
rect -37 9392770 37 9472774
rect -37 9311802 37 9391806
rect -37 9230834 37 9310838
rect -37 9149866 37 9229870
rect -37 9068898 37 9148902
rect -37 8987930 37 9067934
rect -37 8906962 37 8986966
rect -37 8825994 37 8905998
rect -37 8745026 37 8825030
rect -37 8664058 37 8744062
rect -37 8583090 37 8663094
rect -37 8502122 37 8582126
rect -37 8421154 37 8501158
rect -37 8340186 37 8420190
rect -37 8259218 37 8339222
rect -37 8178250 37 8258254
rect -37 8097282 37 8177286
rect -37 8016314 37 8096318
rect -37 7935346 37 8015350
rect -37 7854378 37 7934382
rect -37 7773410 37 7853414
rect -37 7692442 37 7772446
rect -37 7611474 37 7691478
rect -37 7530506 37 7610510
rect -37 7449538 37 7529542
rect -37 7368570 37 7448574
rect -37 7287602 37 7367606
rect -37 7206634 37 7286638
rect -37 7125666 37 7205670
rect -37 7044698 37 7124702
rect -37 6963730 37 7043734
rect -37 6882762 37 6962766
rect -37 6801794 37 6881798
rect -37 6720826 37 6800830
rect -37 6639858 37 6719862
rect -37 6558890 37 6638894
rect -37 6477922 37 6557926
rect -37 6396954 37 6476958
rect -37 6315986 37 6395990
rect -37 6235018 37 6315022
rect -37 6154050 37 6234054
rect -37 6073082 37 6153086
rect -37 5992114 37 6072118
rect -37 5911146 37 5991150
rect -37 5830178 37 5910182
rect -37 5749210 37 5829214
rect -37 5668242 37 5748246
rect -37 5587274 37 5667278
rect -37 5506306 37 5586310
rect -37 5425338 37 5505342
rect -37 5344370 37 5424374
rect -37 5263402 37 5343406
rect -37 5182434 37 5262438
rect -37 5101466 37 5181470
rect -37 5020498 37 5100502
rect -37 4939530 37 5019534
rect -37 4858562 37 4938566
rect -37 4777594 37 4857598
rect -37 4696626 37 4776630
rect -37 4615658 37 4695662
rect -37 4534690 37 4614694
rect -37 4453722 37 4533726
rect -37 4372754 37 4452758
rect -37 4291786 37 4371790
rect -37 4210818 37 4290822
rect -37 4129850 37 4209854
rect -37 4048882 37 4128886
rect -37 3967914 37 4047918
rect -37 3886946 37 3966950
rect -37 3805978 37 3885982
rect -37 3725010 37 3805014
rect -37 3644042 37 3724046
rect -37 3563074 37 3643078
rect -37 3482106 37 3562110
rect -37 3401138 37 3481142
rect -37 3320170 37 3400174
rect -37 3239202 37 3319206
rect -37 3158234 37 3238238
rect -37 3077266 37 3157270
rect -37 2996298 37 3076302
rect -37 2915330 37 2995334
rect -37 2834362 37 2914366
rect -37 2753394 37 2833398
rect -37 2672426 37 2752430
rect -37 2591458 37 2671462
rect -37 2510490 37 2590494
rect -37 2429522 37 2509526
rect -37 2348554 37 2428558
rect -37 2267586 37 2347590
rect -37 2186618 37 2266622
rect -37 2105650 37 2185654
rect -37 2024682 37 2104686
rect -37 1943714 37 2023718
rect -37 1862746 37 1942750
rect -37 1781778 37 1861782
rect -37 1700810 37 1780814
rect -37 1619842 37 1699846
rect -37 1538874 37 1618878
rect -37 1457906 37 1537910
rect -37 1376938 37 1456942
rect -37 1295970 37 1375974
rect -37 1215002 37 1295006
rect -37 1134034 37 1214038
rect -37 1053066 37 1133070
rect -37 972098 37 1052102
rect -37 891130 37 971134
rect -37 810162 37 890166
rect -37 729194 37 809198
rect -37 648226 37 728230
rect -37 567258 37 647262
rect -37 486290 37 566294
rect -37 405322 37 485326
rect -37 324354 37 404358
rect -37 243386 37 323390
rect -37 162418 37 242422
rect -37 81450 37 161454
rect -37 482 37 80486
rect -37 -80486 37 -482
rect -37 -161454 37 -81450
rect -37 -242422 37 -162418
rect -37 -323390 37 -243386
rect -37 -404358 37 -324354
rect -37 -485326 37 -405322
rect -37 -566294 37 -486290
rect -37 -647262 37 -567258
rect -37 -728230 37 -648226
rect -37 -809198 37 -729194
rect -37 -890166 37 -810162
rect -37 -971134 37 -891130
rect -37 -1052102 37 -972098
rect -37 -1133070 37 -1053066
rect -37 -1214038 37 -1134034
rect -37 -1295006 37 -1215002
rect -37 -1375974 37 -1295970
rect -37 -1456942 37 -1376938
rect -37 -1537910 37 -1457906
rect -37 -1618878 37 -1538874
rect -37 -1699846 37 -1619842
rect -37 -1780814 37 -1700810
rect -37 -1861782 37 -1781778
rect -37 -1942750 37 -1862746
rect -37 -2023718 37 -1943714
rect -37 -2104686 37 -2024682
rect -37 -2185654 37 -2105650
rect -37 -2266622 37 -2186618
rect -37 -2347590 37 -2267586
rect -37 -2428558 37 -2348554
rect -37 -2509526 37 -2429522
rect -37 -2590494 37 -2510490
rect -37 -2671462 37 -2591458
rect -37 -2752430 37 -2672426
rect -37 -2833398 37 -2753394
rect -37 -2914366 37 -2834362
rect -37 -2995334 37 -2915330
rect -37 -3076302 37 -2996298
rect -37 -3157270 37 -3077266
rect -37 -3238238 37 -3158234
rect -37 -3319206 37 -3239202
rect -37 -3400174 37 -3320170
rect -37 -3481142 37 -3401138
rect -37 -3562110 37 -3482106
rect -37 -3643078 37 -3563074
rect -37 -3724046 37 -3644042
rect -37 -3805014 37 -3725010
rect -37 -3885982 37 -3805978
rect -37 -3966950 37 -3886946
rect -37 -4047918 37 -3967914
rect -37 -4128886 37 -4048882
rect -37 -4209854 37 -4129850
rect -37 -4290822 37 -4210818
rect -37 -4371790 37 -4291786
rect -37 -4452758 37 -4372754
rect -37 -4533726 37 -4453722
rect -37 -4614694 37 -4534690
rect -37 -4695662 37 -4615658
rect -37 -4776630 37 -4696626
rect -37 -4857598 37 -4777594
rect -37 -4938566 37 -4858562
rect -37 -5019534 37 -4939530
rect -37 -5100502 37 -5020498
rect -37 -5181470 37 -5101466
rect -37 -5262438 37 -5182434
rect -37 -5343406 37 -5263402
rect -37 -5424374 37 -5344370
rect -37 -5505342 37 -5425338
rect -37 -5586310 37 -5506306
rect -37 -5667278 37 -5587274
rect -37 -5748246 37 -5668242
rect -37 -5829214 37 -5749210
rect -37 -5910182 37 -5830178
rect -37 -5991150 37 -5911146
rect -37 -6072118 37 -5992114
rect -37 -6153086 37 -6073082
rect -37 -6234054 37 -6154050
rect -37 -6315022 37 -6235018
rect -37 -6395990 37 -6315986
rect -37 -6476958 37 -6396954
rect -37 -6557926 37 -6477922
rect -37 -6638894 37 -6558890
rect -37 -6719862 37 -6639858
rect -37 -6800830 37 -6720826
rect -37 -6881798 37 -6801794
rect -37 -6962766 37 -6882762
rect -37 -7043734 37 -6963730
rect -37 -7124702 37 -7044698
rect -37 -7205670 37 -7125666
rect -37 -7286638 37 -7206634
rect -37 -7367606 37 -7287602
rect -37 -7448574 37 -7368570
rect -37 -7529542 37 -7449538
rect -37 -7610510 37 -7530506
rect -37 -7691478 37 -7611474
rect -37 -7772446 37 -7692442
rect -37 -7853414 37 -7773410
rect -37 -7934382 37 -7854378
rect -37 -8015350 37 -7935346
rect -37 -8096318 37 -8016314
rect -37 -8177286 37 -8097282
rect -37 -8258254 37 -8178250
rect -37 -8339222 37 -8259218
rect -37 -8420190 37 -8340186
rect -37 -8501158 37 -8421154
rect -37 -8582126 37 -8502122
rect -37 -8663094 37 -8583090
rect -37 -8744062 37 -8664058
rect -37 -8825030 37 -8745026
rect -37 -8905998 37 -8825994
rect -37 -8986966 37 -8906962
rect -37 -9067934 37 -8987930
rect -37 -9148902 37 -9068898
rect -37 -9229870 37 -9149866
rect -37 -9310838 37 -9230834
rect -37 -9391806 37 -9311802
rect -37 -9472774 37 -9392770
rect -37 -9553742 37 -9473738
rect -37 -9634710 37 -9554706
rect -37 -9715678 37 -9635674
rect -37 -9796646 37 -9716642
rect -37 -9877614 37 -9797610
rect -37 -9958582 37 -9878578
rect -37 -10039550 37 -9959546
rect -37 -10120518 37 -10040514
rect -37 -10201486 37 -10121482
rect -37 -10282454 37 -10202450
rect -37 -10363422 37 -10283418
rect -37 -10444390 37 -10364386
rect -37 -10525358 37 -10445354
rect -37 -10606326 37 -10526322
rect -37 -10687294 37 -10607290
rect -37 -10768262 37 -10688258
rect -37 -10849230 37 -10769226
rect -37 -10930198 37 -10850194
rect -37 -11011166 37 -10931162
rect -37 -11092134 37 -11012130
rect -37 -11173102 37 -11093098
rect -37 -11254070 37 -11174066
rect -37 -11335038 37 -11255034
rect -37 -11416006 37 -11336002
rect -37 -11496974 37 -11416970
rect -37 -11577942 37 -11497938
rect -37 -11658910 37 -11578906
rect -37 -11739878 37 -11659874
rect -37 -11820846 37 -11740842
rect -37 -11901814 37 -11821810
rect -37 -11982782 37 -11902778
rect -37 -12063750 37 -11983746
rect -37 -12144718 37 -12064714
rect -37 -12225686 37 -12145682
rect -37 -12306654 37 -12226650
rect -37 -12387622 37 -12307618
rect -37 -12468590 37 -12388586
rect -37 -12549558 37 -12469554
rect -37 -12630526 37 -12550522
rect -37 -12711494 37 -12631490
rect -37 -12792462 37 -12712458
rect -37 -12873430 37 -12793426
rect -37 -12954398 37 -12874394
rect -37 -13035366 37 -12955362
rect -37 -13116334 37 -13036330
rect -37 -13197302 37 -13117298
rect -37 -13278270 37 -13198266
rect -37 -13359238 37 -13279234
rect -37 -13440206 37 -13360202
rect -37 -13521174 37 -13441170
rect -37 -13602142 37 -13522138
rect -37 -13683110 37 -13603106
rect -37 -13764078 37 -13684074
rect -37 -13845046 37 -13765042
rect -37 -13926014 37 -13846010
rect -37 -14006982 37 -13926978
rect -37 -14087950 37 -14007946
rect -37 -14168918 37 -14088914
rect -37 -14249886 37 -14169882
rect -37 -14330854 37 -14250850
rect -37 -14411822 37 -14331818
rect -37 -14492790 37 -14412786
rect -37 -14573758 37 -14493754
rect -37 -14654726 37 -14574722
rect -37 -14735694 37 -14655690
rect -37 -14816662 37 -14736658
rect -37 -14897630 37 -14817626
rect -37 -14978598 37 -14898594
rect -37 -15059566 37 -14979562
rect -37 -15140534 37 -15060530
rect -37 -15221502 37 -15141498
rect -37 -15302470 37 -15222466
rect -37 -15383438 37 -15303434
rect -37 -15464406 37 -15384402
rect -37 -15545374 37 -15465370
rect -37 -15626342 37 -15546338
rect -37 -15707310 37 -15627306
rect -37 -15788278 37 -15708274
rect -37 -15869246 37 -15789242
rect -37 -15950214 37 -15870210
rect -37 -16031182 37 -15951178
rect -37 -16112150 37 -16032146
rect -37 -16193118 37 -16113114
rect -37 -16274086 37 -16194082
rect -37 -16355054 37 -16275050
rect -37 -16436022 37 -16356018
rect -37 -16516990 37 -16436986
rect -37 -16597958 37 -16517954
rect -37 -16678926 37 -16598922
rect -37 -16759894 37 -16679890
rect -37 -16840862 37 -16760858
rect -37 -16921830 37 -16841826
rect -37 -17002798 37 -16922794
rect -37 -17083766 37 -17003762
rect -37 -17164734 37 -17084730
rect -37 -17245702 37 -17165698
rect -37 -17326670 37 -17246666
rect -37 -17407638 37 -17327634
rect -37 -17488606 37 -17408602
rect -37 -17569574 37 -17489570
rect -37 -17650542 37 -17570538
rect -37 -17731510 37 -17651506
rect -37 -17812478 37 -17732474
rect -37 -17893446 37 -17813442
rect -37 -17974414 37 -17894410
rect -37 -18055382 37 -17975378
rect -37 -18136350 37 -18056346
rect -37 -18217318 37 -18137314
rect -37 -18298286 37 -18218282
rect -37 -18379254 37 -18299250
rect -37 -18460222 37 -18380218
rect -37 -18541190 37 -18461186
rect -37 -18622158 37 -18542154
rect -37 -18703126 37 -18623122
rect -37 -18784094 37 -18704090
rect -37 -18865062 37 -18785058
rect -37 -18946030 37 -18866026
rect -37 -19026998 37 -18946994
rect -37 -19107966 37 -19027962
rect -37 -19188934 37 -19108930
rect -37 -19269902 37 -19189898
rect -37 -19350870 37 -19270866
rect -37 -19431838 37 -19351834
rect -37 -19512806 37 -19432802
rect -37 -19593774 37 -19513770
rect -37 -19674742 37 -19594738
rect -37 -19755710 37 -19675706
rect -37 -19836678 37 -19756674
rect -37 -19917646 37 -19837642
rect -37 -19998614 37 -19918610
rect -37 -20079582 37 -19999578
rect -37 -20160550 37 -20080546
rect -37 -20241518 37 -20161514
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -148 -20242061 148 20242061
string parameters w 0.350 l 400 m 500 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 2.285meg dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
