../results/sar_adc_controller.lef