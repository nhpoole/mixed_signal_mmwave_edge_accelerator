magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect 156064 -189722 386940 -57768
rect 182217 -194592 282291 -189722
<< metal1 >>
rect 256482 -91196 256760 -91192
rect 256482 -91248 256492 -91196
rect 256544 -91248 256760 -91196
rect 256482 -91252 256760 -91248
rect 274292 -96736 274352 -96726
rect 270862 -96746 270922 -96736
rect 270862 -96798 270866 -96746
rect 270918 -96798 270922 -96746
rect 268876 -97826 268948 -97822
rect 268876 -97878 268886 -97826
rect 268938 -97878 268948 -97826
rect 268876 -97882 268948 -97878
rect 270862 -98096 270922 -96798
rect 274292 -96788 274296 -96736
rect 274348 -96788 274352 -96736
rect 272572 -98022 272644 -98018
rect 272572 -98074 272582 -98022
rect 272634 -98074 272644 -98022
rect 272572 -98078 272644 -98074
rect 274292 -98264 274352 -96788
rect 245134 -99454 245206 -99450
rect 245134 -99506 245144 -99454
rect 245196 -99506 245206 -99454
rect 245134 -99510 245206 -99506
rect 245140 -101694 245200 -99510
rect 274292 -100230 274352 -100220
rect 274292 -100282 274296 -100230
rect 274348 -100282 274352 -100230
rect 269018 -100962 269090 -100958
rect 269018 -101014 269028 -100962
rect 269080 -101014 269090 -100962
rect 269018 -101018 269090 -101014
rect 244754 -101754 245200 -101694
rect 274292 -101738 274352 -100282
rect 274294 -103230 274354 -101908
rect 274294 -103282 274298 -103230
rect 274350 -103282 274354 -103230
rect 274294 -103292 274354 -103282
rect 272580 -105012 272640 -103626
rect 272580 -105064 272584 -105012
rect 272636 -105064 272640 -105012
rect 272580 -105074 272640 -105064
rect 193222 -106014 193436 -106010
rect 193222 -106066 193374 -106014
rect 193426 -106066 193436 -106014
rect 193222 -106070 193436 -106066
rect 275244 -107968 275304 -107472
rect 275244 -108020 275248 -107968
rect 275300 -108020 275304 -107968
rect 275244 -108030 275304 -108020
rect 243263 -114661 243425 -114603
rect 244188 -114912 244288 -114882
rect 244188 -114964 244212 -114912
rect 244264 -114964 244288 -114912
rect 244188 -114994 244288 -114964
rect 340572 -115934 340632 -115928
rect 340572 -115938 341848 -115934
rect 340572 -115990 340576 -115938
rect 340628 -115990 341848 -115938
rect 340572 -115994 341848 -115990
rect 340572 -116000 340632 -115994
rect 206548 -133850 206780 -133844
rect 201482 -133876 206780 -133850
rect 201482 -134056 206574 -133876
rect 206754 -134056 206780 -133876
rect 201482 -134082 206780 -134056
rect 201482 -135136 201542 -134082
rect 206548 -134088 206780 -134082
rect 207072 -133870 207216 -133850
rect 207072 -133986 207086 -133870
rect 207202 -133986 207216 -133870
rect 201482 -135196 201624 -135136
rect 199354 -136092 199498 -136086
rect 207072 -136092 207216 -133986
rect 199354 -136106 207216 -136092
rect 199354 -136222 199368 -136106
rect 199484 -136222 207216 -136106
rect 199354 -136236 207216 -136222
rect 207458 -134758 207558 -134728
rect 207458 -134810 207482 -134758
rect 207534 -134810 207558 -134758
rect 199354 -136242 199498 -136236
rect 207458 -136628 207558 -134810
rect 207452 -136652 207564 -136628
rect 207452 -136704 207482 -136652
rect 207534 -136704 207564 -136652
rect 207452 -136728 207564 -136704
rect 204118 -146174 204230 -146150
rect 204118 -146226 204148 -146174
rect 204200 -146226 204230 -146174
rect 204118 -146250 204230 -146226
rect 204124 -148036 204224 -146250
rect 204124 -148088 204148 -148036
rect 204200 -148088 204224 -148036
rect 204124 -148118 204224 -148088
rect 195644 -149028 195704 -149022
rect 193666 -149032 195704 -149028
rect 193666 -149084 195648 -149032
rect 195700 -149084 195704 -149032
rect 193666 -149088 195704 -149084
rect 195644 -149094 195704 -149088
rect 259992 -149032 260052 -149026
rect 259992 -149036 260920 -149032
rect 259992 -149088 259996 -149036
rect 260048 -149088 260920 -149036
rect 259992 -149092 260920 -149088
rect 259992 -149098 260052 -149092
rect 340704 -166944 340764 -166938
rect 340704 -166948 341756 -166944
rect 340704 -167000 340708 -166948
rect 340760 -167000 341756 -166948
rect 340704 -167004 341756 -167000
rect 340704 -167010 340764 -167004
rect 339824 -182370 339896 -182366
rect 339824 -182422 339834 -182370
rect 339886 -182422 339896 -182370
rect 339824 -182426 339896 -182422
rect 259902 -183556 259962 -183550
rect 184660 -183560 185024 -183556
rect 184660 -183612 184962 -183560
rect 185014 -183612 185024 -183560
rect 184660 -183616 185024 -183612
rect 225734 -183560 226020 -183556
rect 225734 -183612 225958 -183560
rect 226010 -183612 226020 -183560
rect 225734 -183616 226020 -183612
rect 259902 -183560 260944 -183556
rect 259902 -183612 259906 -183560
rect 259958 -183612 260944 -183560
rect 259902 -183616 260944 -183612
rect 259902 -183622 259962 -183616
rect 339580 -184698 339676 -184692
rect 333766 -184720 339676 -184698
rect 333766 -184772 333794 -184720
rect 333846 -184772 339602 -184720
rect 339654 -184772 339676 -184720
rect 333766 -184794 339676 -184772
rect 339580 -184800 339676 -184794
rect 339678 -184900 339800 -184896
rect 339678 -184952 339738 -184900
rect 339790 -184952 339800 -184900
rect 339678 -184956 339800 -184952
rect 334778 -185024 334838 -185018
rect 339830 -185020 339890 -182426
rect 334778 -185028 335058 -185024
rect 334778 -185080 334782 -185028
rect 334834 -185080 335058 -185028
rect 339462 -185080 339890 -185020
rect 334778 -185084 335058 -185080
rect 334778 -185090 334838 -185084
rect 334540 -185242 334636 -185236
rect 334540 -185264 339606 -185242
rect 334540 -185316 334562 -185264
rect 334614 -185316 339606 -185264
rect 334540 -185338 339606 -185316
rect 334540 -185344 334636 -185338
rect 333758 -185808 339474 -185786
rect 333758 -185860 333786 -185808
rect 333838 -185860 339474 -185808
rect 333758 -185882 339474 -185860
<< via1 >>
rect 256492 -91248 256544 -91196
rect 270866 -96798 270918 -96746
rect 268886 -97878 268938 -97826
rect 274296 -96788 274348 -96736
rect 272582 -98074 272634 -98022
rect 245144 -99506 245196 -99454
rect 274296 -100282 274348 -100230
rect 269028 -101014 269080 -100962
rect 274298 -103282 274350 -103230
rect 272584 -105064 272636 -105012
rect 193374 -106066 193426 -106014
rect 275248 -108020 275300 -107968
rect 244212 -114964 244264 -114912
rect 340576 -115990 340628 -115938
rect 206574 -134056 206754 -133876
rect 207086 -133986 207202 -133870
rect 199368 -136222 199484 -136106
rect 207482 -134810 207534 -134758
rect 207482 -136704 207534 -136652
rect 204148 -146226 204200 -146174
rect 204148 -148088 204200 -148036
rect 195648 -149084 195700 -149032
rect 259996 -149088 260048 -149036
rect 340708 -167000 340760 -166948
rect 339834 -182422 339886 -182370
rect 184962 -183612 185014 -183560
rect 225958 -183612 226010 -183560
rect 259906 -183612 259958 -183560
rect 333794 -184772 333846 -184720
rect 339602 -184772 339654 -184720
rect 339738 -184952 339790 -184900
rect 334782 -185080 334834 -185028
rect 334562 -185316 334614 -185264
rect 333786 -185860 333838 -185808
<< metal2 >>
rect 199381 -83670 199441 -83504
rect 250374 -91196 256566 -91166
rect 250374 -91248 256492 -91196
rect 256544 -91248 256566 -91196
rect 250374 -91294 256566 -91248
rect 196484 -91585 196584 -91580
rect 196480 -91602 196588 -91585
rect 196480 -91658 196506 -91602
rect 196562 -91658 196588 -91602
rect 196480 -91675 196588 -91658
rect 194320 -91947 194420 -91942
rect 194316 -91964 194424 -91947
rect 194316 -92020 194342 -91964
rect 194398 -92020 194424 -91964
rect 194316 -92037 194424 -92020
rect 193370 -106010 193430 -106004
rect 193361 -106012 193439 -106010
rect 193361 -106068 193372 -106012
rect 193428 -106068 193439 -106012
rect 193361 -106070 193439 -106068
rect 193370 -106076 193430 -106070
rect 194320 -107740 194420 -92037
rect 190376 -107840 194420 -107740
rect 190376 -108711 190476 -107840
rect 190372 -108728 190480 -108711
rect 190372 -108784 190398 -108728
rect 190454 -108784 190480 -108728
rect 190372 -108801 190480 -108784
rect 190376 -108806 190476 -108801
rect 196484 -109367 196584 -91675
rect 250374 -92336 250502 -91294
rect 250374 -92392 250410 -92336
rect 250466 -92392 250502 -92336
rect 250374 -92437 250502 -92392
rect 266828 -96330 266980 -96291
rect 266828 -96386 266876 -96330
rect 266932 -96386 266980 -96330
rect 279692 -96386 280120 -96326
rect 266828 -96425 266980 -96386
rect 265964 -96582 266148 -96567
rect 265964 -96718 265988 -96582
rect 266124 -96718 266148 -96582
rect 265964 -96733 266148 -96718
rect 265471 -97782 265703 -97743
rect 265471 -97918 265519 -97782
rect 265655 -97918 265703 -97782
rect 265471 -97957 265703 -97918
rect 245104 -99452 262677 -99413
rect 245104 -99454 262573 -99452
rect 245104 -99506 245144 -99454
rect 245196 -99506 262573 -99454
rect 245104 -99508 262573 -99506
rect 262629 -99508 262677 -99452
rect 245104 -99546 262677 -99508
rect 265030 -100918 265198 -100911
rect 265030 -101054 265046 -100918
rect 265182 -101054 265198 -100918
rect 265030 -101061 265198 -101054
rect 250374 -101205 250502 -101200
rect 250370 -101236 250506 -101205
rect 250370 -101292 250410 -101236
rect 250466 -101292 250506 -101236
rect 250370 -101323 250506 -101292
rect 197955 -102432 198015 -102238
rect 198780 -107742 198928 -107705
rect 198780 -107798 198826 -107742
rect 198882 -107798 198928 -107742
rect 198780 -107835 198928 -107798
rect 198789 -109177 198919 -107835
rect 210625 -108120 210634 -107984
rect 210770 -108120 210779 -107984
rect 198475 -109307 198919 -109177
rect 196480 -109384 196588 -109367
rect 196480 -109440 196506 -109384
rect 196562 -109440 196588 -109384
rect 196480 -109457 196588 -109440
rect 196484 -109462 196584 -109457
rect 191447 -110136 191525 -110134
rect 191447 -110192 191458 -110136
rect 191514 -110192 191525 -110136
rect 191447 -110194 191525 -110192
rect 191456 -111380 191516 -110194
rect 194516 -110650 194576 -110641
rect 193494 -110652 194576 -110650
rect 193494 -110708 194518 -110652
rect 194574 -110708 194576 -110652
rect 193494 -110710 194576 -110708
rect 194516 -110719 194576 -110710
rect 191456 -111440 192132 -111380
rect 198475 -112253 198605 -109307
rect 210634 -112248 210770 -108120
rect 211052 -108294 211196 -108259
rect 211052 -108350 211096 -108294
rect 211152 -108350 211196 -108294
rect 211052 -108385 211196 -108350
rect 198471 -112285 198609 -112253
rect 196578 -112288 196859 -112286
rect 196578 -112344 196792 -112288
rect 196848 -112344 196859 -112288
rect 196578 -112346 196859 -112344
rect 198471 -112341 198512 -112285
rect 198568 -112341 198609 -112285
rect 208548 -112286 210770 -112248
rect 198471 -112373 198609 -112341
rect 208476 -112346 210770 -112286
rect 198475 -112378 198605 -112373
rect 208548 -112384 210770 -112346
rect 210170 -114691 210286 -114687
rect 211061 -114691 211187 -108385
rect 211294 -108608 211446 -108569
rect 211294 -108664 211342 -108608
rect 211398 -108664 211446 -108608
rect 211294 -108703 211446 -108664
rect 210165 -114726 211187 -114691
rect 210165 -114782 210200 -114726
rect 210256 -114782 211187 -114726
rect 210165 -114817 211187 -114782
rect 210170 -114821 210286 -114817
rect 211303 -115213 211437 -108703
rect 212365 -108906 212527 -108902
rect 212365 -109042 212378 -108906
rect 212514 -109042 212527 -108906
rect 212365 -109046 212527 -109042
rect 211557 -114910 211647 -114906
rect 208557 -115250 211437 -115213
rect 196618 -115252 196857 -115250
rect 196618 -115308 196790 -115252
rect 196846 -115308 196857 -115252
rect 196618 -115310 196857 -115308
rect 208484 -115310 211437 -115250
rect 208557 -115347 211437 -115310
rect 211552 -114932 211652 -114910
rect 211552 -114988 211574 -114932
rect 211630 -114988 211652 -114932
rect 210524 -115768 210624 -115766
rect 211552 -115768 211652 -114988
rect 210522 -115771 211652 -115768
rect 210520 -115788 211652 -115771
rect 210520 -115844 210546 -115788
rect 210602 -115844 211652 -115788
rect 210520 -115861 211652 -115844
rect 210522 -115868 211652 -115861
rect 207458 -120845 207558 -120840
rect 207454 -120862 207562 -120845
rect 207454 -120918 207480 -120862
rect 207536 -120918 207562 -120862
rect 207454 -120935 207562 -120918
rect 207063 -121642 207225 -121638
rect 207063 -121778 207076 -121642
rect 207212 -121778 207225 -121642
rect 207063 -121782 207225 -121778
rect 206548 -121959 206780 -121954
rect 206544 -121962 206784 -121959
rect 206544 -122178 206556 -121962
rect 206772 -122178 206784 -121962
rect 206544 -122181 206784 -122178
rect 206548 -133850 206780 -122181
rect 206542 -133876 206786 -133850
rect 207072 -133856 207216 -121782
rect 206542 -134056 206574 -133876
rect 206754 -134056 206786 -133876
rect 207066 -133870 207222 -133856
rect 207066 -133986 207086 -133870
rect 207202 -133986 207222 -133870
rect 207066 -134000 207222 -133986
rect 206542 -134082 206786 -134056
rect 207458 -134734 207558 -120935
rect 210524 -122264 210624 -115868
rect 210794 -116871 210894 -116866
rect 210790 -116888 210898 -116871
rect 210790 -116944 210816 -116888
rect 210872 -116944 210898 -116888
rect 210790 -116961 210898 -116944
rect 208246 -122364 210624 -122264
rect 207452 -134758 207564 -134734
rect 207452 -134810 207482 -134758
rect 207534 -134810 207564 -134758
rect 207452 -134834 207564 -134810
rect 207458 -134838 207558 -134834
rect 195602 -136106 199504 -136092
rect 195602 -136222 199368 -136106
rect 199484 -136222 199504 -136106
rect 195602 -136236 199504 -136222
rect 195602 -136480 195746 -136236
rect 195602 -136536 195646 -136480
rect 195702 -136536 195746 -136480
rect 195602 -136580 195746 -136536
rect 195607 -136584 195741 -136580
rect 207458 -136652 207558 -136622
rect 207458 -136704 207482 -136652
rect 207534 -136704 207558 -136652
rect 205993 -137496 206083 -137492
rect 207458 -137496 207558 -136704
rect 205988 -137518 207558 -137496
rect 205988 -137574 206010 -137518
rect 206066 -137574 207558 -137518
rect 205988 -137596 207558 -137574
rect 205993 -137600 206083 -137596
rect 204124 -143645 204224 -143640
rect 204120 -143662 204228 -143645
rect 204120 -143718 204146 -143662
rect 204202 -143718 204228 -143662
rect 204120 -143735 204228 -143718
rect 204124 -146174 204224 -143735
rect 204811 -144748 204901 -144744
rect 208246 -144748 208346 -122364
rect 204806 -144770 208346 -144748
rect 204806 -144826 204828 -144770
rect 204884 -144826 208346 -144770
rect 204806 -144848 208346 -144826
rect 204811 -144852 204901 -144848
rect 204124 -146226 204148 -146174
rect 204200 -146226 204224 -146174
rect 204124 -146256 204224 -146226
rect 158376 -146554 158508 -146518
rect 158376 -146614 160676 -146554
rect 158376 -151698 158508 -146614
rect 204124 -148012 204224 -147992
rect 204118 -148036 204230 -148012
rect 204118 -148088 204148 -148036
rect 204200 -148088 204230 -148036
rect 204118 -148112 204230 -148088
rect 195644 -149028 195704 -149019
rect 195638 -149030 195710 -149028
rect 195638 -149086 195646 -149030
rect 195702 -149086 195710 -149030
rect 195638 -149088 195710 -149086
rect 195644 -149097 195704 -149088
rect 204124 -153944 204224 -148112
rect 205627 -149274 205717 -149270
rect 210794 -149274 210894 -116961
rect 212374 -121643 212518 -109046
rect 245669 -109259 245853 -109244
rect 245669 -109395 245693 -109259
rect 245829 -109395 245853 -109259
rect 245669 -109410 245853 -109395
rect 232501 -109650 232657 -109649
rect 232501 -109786 232511 -109650
rect 232647 -109786 232657 -109650
rect 232501 -109787 232657 -109786
rect 218166 -110148 218334 -110141
rect 218166 -110284 218182 -110148
rect 218318 -110284 218334 -110148
rect 218166 -110291 218334 -110284
rect 212802 -110527 213034 -110522
rect 212798 -110530 213038 -110527
rect 212798 -110746 212810 -110530
rect 213026 -110746 213038 -110530
rect 212798 -110749 213038 -110746
rect 212370 -121682 212522 -121643
rect 212370 -121738 212418 -121682
rect 212474 -121738 212522 -121682
rect 212370 -121777 212522 -121738
rect 212374 -121782 212518 -121777
rect 212802 -121954 213034 -110749
rect 212793 -121962 213043 -121954
rect 212793 -122178 212810 -121962
rect 213026 -122178 213043 -121962
rect 212793 -122186 213043 -122178
rect 205622 -149296 210896 -149274
rect 205622 -149352 205644 -149296
rect 205700 -149352 210896 -149296
rect 205622 -149374 210896 -149352
rect 205627 -149378 205717 -149374
rect 204124 -154044 210658 -153944
rect 210258 -155220 210426 -155213
rect 210258 -155356 210274 -155220
rect 210410 -155356 210426 -155220
rect 210258 -155363 210426 -155356
rect 210036 -169589 210136 -169584
rect 210032 -169606 210140 -169589
rect 210032 -169662 210058 -169606
rect 210114 -169662 210140 -169606
rect 210032 -169679 210140 -169662
rect 186411 -183511 186561 -183502
rect 184913 -183518 186561 -183511
rect 184913 -183560 186418 -183518
rect 184913 -183612 184962 -183560
rect 185014 -183612 186418 -183560
rect 184913 -183654 186418 -183612
rect 186554 -183654 186561 -183518
rect 184913 -183661 186561 -183654
rect 186411 -183670 186561 -183661
rect 210036 -184536 210136 -169679
rect 210267 -170068 210417 -155363
rect 210263 -170070 210421 -170068
rect 210263 -170206 210274 -170070
rect 210410 -170206 210421 -170070
rect 210263 -170208 210421 -170206
rect 210267 -170213 210417 -170208
rect 210558 -170706 210658 -154044
rect 218175 -155218 218325 -110291
rect 231559 -113868 231637 -113866
rect 231559 -113924 231570 -113868
rect 231626 -113924 231637 -113868
rect 231559 -113926 231637 -113924
rect 225357 -114930 226682 -114928
rect 225357 -114986 225368 -114930
rect 225424 -114986 226682 -114930
rect 225357 -114988 226682 -114986
rect 225367 -115466 226956 -115464
rect 225367 -115522 225378 -115466
rect 225434 -115522 226956 -115466
rect 225367 -115524 226956 -115522
rect 232510 -116116 232648 -109787
rect 244188 -113851 244288 -113846
rect 244184 -113868 244292 -113851
rect 244184 -113924 244210 -113868
rect 244266 -113924 244292 -113868
rect 244184 -113941 244292 -113924
rect 244188 -114888 244288 -113941
rect 244182 -114912 244294 -114888
rect 244182 -114964 244212 -114912
rect 244264 -114964 244294 -114912
rect 244182 -114988 244294 -114964
rect 231798 -116176 232648 -116116
rect 245678 -116588 245844 -109410
rect 250374 -110560 250502 -101323
rect 264162 -101968 264326 -101963
rect 264162 -102104 264176 -101968
rect 264312 -102104 264326 -101968
rect 264162 -102109 264326 -102104
rect 263725 -105258 263903 -105246
rect 263725 -105394 263746 -105258
rect 263882 -105394 263903 -105258
rect 263725 -105406 263903 -105394
rect 250732 -110550 250908 -110539
rect 250365 -110596 250511 -110560
rect 250365 -110652 250410 -110596
rect 250466 -110652 250511 -110596
rect 250365 -110688 250511 -110652
rect 250732 -110686 250752 -110550
rect 250888 -110686 250908 -110550
rect 250732 -110697 250908 -110686
rect 250329 -111326 250507 -111314
rect 250329 -111462 250350 -111326
rect 250486 -111462 250507 -111326
rect 250329 -111474 250507 -111462
rect 243378 -116648 245844 -116588
rect 234399 -150312 234522 -150280
rect 234276 -150372 234522 -150312
rect 234399 -151436 234522 -150372
rect 234390 -151470 234531 -151436
rect 234390 -151526 234432 -151470
rect 234488 -151526 234531 -151470
rect 234390 -151559 234531 -151526
rect 250338 -151701 250498 -111474
rect 250334 -151708 250502 -151701
rect 250334 -151844 250350 -151708
rect 250486 -151844 250502 -151708
rect 250334 -151851 250502 -151844
rect 250338 -151856 250498 -151851
rect 218171 -155220 218329 -155218
rect 218171 -155356 218182 -155220
rect 218318 -155356 218329 -155220
rect 218171 -155358 218329 -155356
rect 218175 -155363 218325 -155358
rect 250741 -169266 250899 -110697
rect 255262 -110948 255426 -110943
rect 255262 -111084 255276 -110948
rect 255412 -111084 255426 -110948
rect 255262 -111089 255426 -111084
rect 255271 -135621 255417 -111089
rect 263734 -111319 263894 -105406
rect 264171 -110948 264317 -102109
rect 264578 -103382 264754 -103371
rect 264578 -103518 264598 -103382
rect 264734 -103518 264754 -103382
rect 264578 -103529 264754 -103518
rect 264587 -110544 264745 -103529
rect 265039 -110146 265189 -101061
rect 265480 -109621 265694 -97957
rect 265973 -109249 266139 -96733
rect 266427 -100036 266589 -100032
rect 266427 -100172 266440 -100036
rect 266576 -100172 266589 -100036
rect 266427 -100176 266589 -100172
rect 266436 -108907 266580 -100176
rect 266837 -108574 266971 -96425
rect 274292 -96732 274352 -96723
rect 270862 -96742 270922 -96733
rect 274286 -96734 274358 -96732
rect 270856 -96744 270928 -96742
rect 270856 -96800 270864 -96744
rect 270920 -96800 270928 -96744
rect 274286 -96790 274294 -96734
rect 274350 -96790 274358 -96734
rect 274286 -96792 274358 -96790
rect 270856 -96802 270928 -96800
rect 274292 -96801 274352 -96792
rect 270862 -96811 270922 -96802
rect 268882 -97822 268942 -97816
rect 268873 -97824 268951 -97822
rect 268873 -97880 268884 -97824
rect 268940 -97880 268951 -97824
rect 268873 -97882 268951 -97880
rect 268882 -97888 268942 -97882
rect 272578 -98020 272638 -98009
rect 272578 -98076 272580 -98020
rect 272636 -98076 272638 -98020
rect 267503 -98218 267512 -98082
rect 267648 -98218 267657 -98082
rect 272578 -98087 272638 -98076
rect 267190 -98388 267334 -98353
rect 267190 -98444 267234 -98388
rect 267290 -98444 267334 -98388
rect 267190 -98479 267334 -98444
rect 267199 -108264 267325 -98479
rect 267512 -107989 267648 -98218
rect 267842 -98312 269144 -98252
rect 267842 -98316 267971 -98312
rect 267841 -107710 267971 -98316
rect 274283 -98360 274454 -98358
rect 274283 -98416 274296 -98360
rect 274352 -98416 274454 -98360
rect 274283 -98418 274454 -98416
rect 377155 -99057 377301 -99056
rect 377155 -99117 378347 -99057
rect 268407 -99417 268540 -99411
rect 268403 -99451 268544 -99417
rect 268403 -99507 268445 -99451
rect 268501 -99507 268544 -99451
rect 268403 -99540 268544 -99507
rect 268407 -101632 268540 -99540
rect 274292 -100226 274352 -100217
rect 274286 -100228 274358 -100226
rect 274286 -100284 274294 -100228
rect 274350 -100284 274358 -100228
rect 274286 -100286 274358 -100284
rect 274292 -100295 274352 -100286
rect 269024 -100958 269084 -100952
rect 269015 -100960 269093 -100958
rect 269015 -101016 269026 -100960
rect 269082 -101016 269093 -100960
rect 269015 -101018 269093 -101016
rect 269024 -101024 269084 -101018
rect 268407 -101692 270994 -101632
rect 268136 -101736 268276 -101694
rect 268136 -101792 268178 -101736
rect 268234 -101792 268276 -101736
rect 268136 -107404 268276 -101792
rect 272569 -101736 272816 -101734
rect 272569 -101792 272580 -101736
rect 272636 -101792 272816 -101736
rect 272569 -101794 272816 -101792
rect 268882 -101898 269030 -101838
rect 268882 -101998 268942 -101898
rect 268873 -102000 268951 -101998
rect 268873 -102056 268884 -102000
rect 268940 -102056 268951 -102000
rect 268873 -102058 268951 -102056
rect 274294 -103226 274354 -103217
rect 274288 -103228 274360 -103226
rect 274288 -103284 274296 -103228
rect 274352 -103284 274360 -103228
rect 274288 -103286 274360 -103284
rect 274294 -103295 274354 -103286
rect 295787 -103424 296978 -103412
rect 279388 -103540 279556 -103533
rect 279388 -103676 279404 -103540
rect 279540 -103676 279556 -103540
rect 295787 -103560 295808 -103424
rect 295944 -103560 296978 -103424
rect 295787 -103572 296978 -103560
rect 279388 -103683 279556 -103676
rect 272580 -105008 272640 -104999
rect 272574 -105010 272646 -105008
rect 272574 -105066 272582 -105010
rect 272638 -105066 272646 -105010
rect 272574 -105068 272646 -105066
rect 295832 -105068 296000 -105060
rect 272580 -105077 272640 -105068
rect 275896 -105110 276081 -105108
rect 275896 -105166 276014 -105110
rect 276070 -105166 276081 -105110
rect 275896 -105168 276081 -105166
rect 295832 -105204 295850 -105068
rect 295986 -105204 296000 -105068
rect 294183 -107365 294325 -107360
rect 275792 -107402 276231 -107400
rect 268127 -107406 268285 -107404
rect 268127 -107542 268138 -107406
rect 268274 -107542 268285 -107406
rect 275792 -107458 276164 -107402
rect 276220 -107458 276231 -107402
rect 275792 -107460 276231 -107458
rect 294179 -107403 294329 -107365
rect 294179 -107459 294226 -107403
rect 294282 -107459 294329 -107403
rect 294179 -107497 294329 -107459
rect 268127 -107544 268285 -107542
rect 267837 -107742 267975 -107710
rect 267837 -107798 267878 -107742
rect 267934 -107798 267975 -107742
rect 267837 -107830 267975 -107798
rect 267841 -107835 267971 -107830
rect 275244 -107964 275304 -107955
rect 275238 -107966 275310 -107964
rect 267508 -108024 267652 -107989
rect 275238 -108022 275246 -107966
rect 275302 -108022 275310 -107966
rect 275238 -108024 275310 -108022
rect 267508 -108080 267552 -108024
rect 267608 -108080 267652 -108024
rect 275244 -108033 275304 -108024
rect 267508 -108115 267652 -108080
rect 267512 -108120 267648 -108115
rect 275830 -108160 276144 -108100
rect 267195 -108294 267329 -108264
rect 267195 -108350 267234 -108294
rect 267290 -108350 267329 -108294
rect 267195 -108380 267329 -108350
rect 267199 -108385 267325 -108380
rect 266833 -108608 266975 -108574
rect 266833 -108664 266876 -108608
rect 266932 -108664 266975 -108608
rect 266833 -108698 266975 -108664
rect 266837 -108703 266971 -108698
rect 266432 -108946 266584 -108907
rect 266432 -109002 266480 -108946
rect 266536 -109002 266584 -108946
rect 266432 -109041 266584 -109002
rect 266436 -109046 266580 -109041
rect 265969 -109259 266143 -109249
rect 265969 -109395 265988 -109259
rect 266124 -109395 266143 -109259
rect 265969 -109405 266143 -109395
rect 265973 -109410 266139 -109405
rect 265476 -109655 265698 -109621
rect 265476 -109791 265519 -109655
rect 265655 -109791 265698 -109655
rect 265476 -109825 265698 -109791
rect 265480 -109830 265694 -109825
rect 265035 -110148 265193 -110146
rect 265035 -110284 265046 -110148
rect 265182 -110284 265193 -110148
rect 265035 -110286 265193 -110284
rect 265039 -110291 265189 -110286
rect 264583 -110550 264749 -110544
rect 264583 -110686 264598 -110550
rect 264734 -110686 264749 -110550
rect 264583 -110692 264749 -110686
rect 264587 -110697 264745 -110692
rect 264167 -111084 264176 -110948
rect 264312 -111084 264321 -110948
rect 264171 -111089 264317 -111084
rect 263730 -111326 263898 -111319
rect 263730 -111462 263746 -111326
rect 263882 -111462 263898 -111326
rect 263730 -111469 263898 -111462
rect 263734 -111474 263894 -111469
rect 294183 -124565 294325 -107497
rect 294571 -108186 294717 -108181
rect 294567 -108322 294576 -108186
rect 294712 -108322 294721 -108186
rect 294571 -122067 294717 -108322
rect 294562 -122072 294726 -122067
rect 294562 -122208 294576 -122072
rect 294712 -122208 294726 -122072
rect 294562 -122213 294726 -122208
rect 295832 -122784 296000 -105204
rect 296818 -122434 296978 -103572
rect 340522 -115938 340682 -115884
rect 340522 -115990 340576 -115938
rect 340628 -115990 340682 -115938
rect 340080 -118426 340244 -118421
rect 340080 -118562 340094 -118426
rect 340230 -118562 340244 -118426
rect 340080 -118567 340244 -118562
rect 297540 -122067 297676 -122063
rect 340089 -122067 340235 -118567
rect 297535 -122072 340235 -122067
rect 297535 -122208 297540 -122072
rect 297676 -122208 340235 -122072
rect 297535 -122213 340235 -122208
rect 297540 -122217 297676 -122213
rect 340522 -122434 340682 -115990
rect 377155 -118426 377301 -99117
rect 384590 -101032 384986 -100972
rect 377792 -101582 378406 -101522
rect 377151 -118562 377160 -118426
rect 377296 -118562 377305 -118426
rect 377155 -118567 377301 -118562
rect 296818 -122594 340682 -122434
rect 295832 -122952 336052 -122784
rect 294183 -124707 295881 -124565
rect 255271 -135767 260089 -135621
rect 259943 -136115 260089 -135767
rect 259943 -136120 260094 -136115
rect 259943 -136256 259953 -136120
rect 260089 -136256 260094 -136120
rect 259943 -136261 260094 -136256
rect 259943 -136265 260089 -136261
rect 294513 -136612 294603 -136586
rect 294513 -136668 294530 -136612
rect 294586 -136668 294603 -136612
rect 294513 -136694 294603 -136668
rect 295221 -136937 295356 -136906
rect 295221 -136993 295260 -136937
rect 295316 -136993 295356 -136937
rect 295221 -137023 295356 -136993
rect 259992 -149032 260052 -149023
rect 259986 -149034 260058 -149032
rect 259986 -149090 259994 -149034
rect 260050 -149090 260058 -149034
rect 259986 -149092 260058 -149090
rect 259992 -149101 260052 -149092
rect 251432 -149386 254490 -149286
rect 258310 -149306 258370 -149297
rect 256528 -149308 258370 -149306
rect 256528 -149364 258312 -149308
rect 258368 -149364 258370 -149308
rect 256528 -149366 258370 -149364
rect 258310 -149375 258370 -149366
rect 250737 -169272 250903 -169266
rect 250737 -169408 250752 -169272
rect 250888 -169408 250903 -169272
rect 250737 -169414 250903 -169408
rect 250741 -169419 250899 -169414
rect 210558 -170806 214418 -170706
rect 214318 -179624 214418 -170806
rect 214318 -179684 216972 -179624
rect 227633 -183507 227791 -183498
rect 225905 -183518 227791 -183507
rect 225905 -183560 227644 -183518
rect 225905 -183612 225958 -183560
rect 226010 -183612 227644 -183560
rect 225905 -183654 227644 -183612
rect 227780 -183654 227791 -183518
rect 225905 -183665 227791 -183654
rect 227633 -183674 227791 -183665
rect 251432 -183810 251532 -149386
rect 295230 -150297 295347 -137023
rect 295739 -137257 295881 -124707
rect 298051 -126571 298111 -126488
rect 297116 -126947 297216 -126942
rect 297112 -126964 297220 -126947
rect 297112 -127020 297138 -126964
rect 297194 -127020 297220 -126964
rect 297112 -127037 297220 -127020
rect 297116 -136590 297216 -127037
rect 298023 -131005 298140 -126571
rect 297454 -131122 298140 -131005
rect 297107 -136612 297225 -136590
rect 297107 -136668 297138 -136612
rect 297194 -136668 297225 -136612
rect 297107 -136690 297225 -136668
rect 297454 -136910 297571 -131122
rect 298051 -135004 298111 -133004
rect 298042 -135006 298120 -135004
rect 298042 -135062 298053 -135006
rect 298109 -135062 298120 -135006
rect 298042 -135064 298120 -135062
rect 302051 -135296 302111 -132954
rect 302042 -135298 302120 -135296
rect 302042 -135354 302053 -135298
rect 302109 -135354 302120 -135298
rect 302042 -135356 302120 -135354
rect 306051 -135604 306111 -133004
rect 306042 -135606 306120 -135604
rect 306042 -135662 306053 -135606
rect 306109 -135662 306120 -135606
rect 306042 -135664 306120 -135662
rect 310051 -135888 310111 -132804
rect 310042 -135890 310120 -135888
rect 310042 -135946 310053 -135890
rect 310109 -135946 310120 -135890
rect 310042 -135948 310120 -135946
rect 314051 -136184 314111 -132976
rect 314042 -136186 314120 -136184
rect 314042 -136242 314053 -136186
rect 314109 -136242 314120 -136186
rect 314042 -136244 314120 -136242
rect 318051 -136470 318111 -132934
rect 318042 -136472 318120 -136470
rect 318042 -136528 318053 -136472
rect 318109 -136528 318120 -136472
rect 318042 -136530 318120 -136528
rect 326051 -136746 326111 -132948
rect 326042 -136748 326120 -136746
rect 326042 -136804 326053 -136748
rect 326109 -136804 326120 -136748
rect 326042 -136806 326120 -136804
rect 297453 -136936 297578 -136910
rect 297453 -136992 297487 -136936
rect 297543 -136992 297578 -136936
rect 297453 -137017 297578 -136992
rect 297454 -137020 297571 -137017
rect 330051 -137040 330111 -132928
rect 330042 -137042 330120 -137040
rect 330042 -137098 330053 -137042
rect 330109 -137098 330120 -137042
rect 330042 -137100 330120 -137098
rect 295739 -137423 334893 -137257
rect 334727 -138572 334893 -137423
rect 334723 -138582 334897 -138572
rect 334723 -138718 334742 -138582
rect 334878 -138718 334897 -138582
rect 334723 -138728 334897 -138718
rect 334727 -138733 334893 -138728
rect 295221 -150328 295356 -150297
rect 253223 -150380 253336 -150377
rect 253218 -150415 253831 -150380
rect 295221 -150384 295260 -150328
rect 295316 -150384 295356 -150328
rect 295221 -150414 295356 -150384
rect 253218 -150471 253251 -150415
rect 253307 -150471 253831 -150415
rect 253218 -150503 253831 -150471
rect 253223 -150508 253336 -150503
rect 255065 -151708 255243 -151696
rect 255065 -151844 255086 -151708
rect 255222 -151844 255243 -151708
rect 255065 -151856 255243 -151844
rect 255074 -170066 255234 -151856
rect 335884 -154082 336052 -122952
rect 336237 -137362 336355 -137340
rect 336237 -137418 336268 -137362
rect 336324 -137418 336355 -137362
rect 336237 -137440 336355 -137418
rect 336246 -153801 336346 -137440
rect 377792 -152532 377992 -101582
rect 378162 -137362 378346 -137347
rect 378162 -137498 378186 -137362
rect 378322 -137498 378346 -137362
rect 378162 -137513 378346 -137498
rect 378171 -150067 378337 -137513
rect 378171 -150127 378347 -150067
rect 378171 -150180 378337 -150127
rect 384612 -152042 385152 -151982
rect 377792 -152592 378402 -152532
rect 336242 -153818 336350 -153801
rect 336242 -153874 336268 -153818
rect 336324 -153874 336350 -153818
rect 336242 -153891 336350 -153874
rect 336246 -153896 336346 -153891
rect 335884 -154250 340818 -154082
rect 340650 -166948 340818 -154250
rect 340650 -167000 340708 -166948
rect 340760 -167000 340818 -166948
rect 340650 -167058 340818 -167000
rect 255074 -170226 260016 -170066
rect 259856 -170776 260016 -170226
rect 377792 -170574 377992 -152592
rect 377783 -170606 378001 -170574
rect 259854 -170820 260016 -170776
rect 259854 -170956 259866 -170820
rect 260002 -170956 260016 -170820
rect 259854 -170974 260016 -170956
rect 340100 -170658 340210 -170644
rect 340100 -170714 340118 -170658
rect 340174 -170714 340210 -170658
rect 259854 -170977 260014 -170974
rect 294346 -175038 294599 -175036
rect 294346 -175094 294532 -175038
rect 294588 -175094 294599 -175038
rect 294346 -175096 294599 -175094
rect 299029 -178194 299192 -178192
rect 299029 -178250 299040 -178194
rect 299096 -178250 299192 -178194
rect 299029 -178252 299192 -178250
rect 334540 -180272 334636 -180243
rect 334540 -180328 334560 -180272
rect 334616 -180328 334636 -180272
rect 259902 -183556 259962 -183547
rect 259896 -183558 259968 -183556
rect 259896 -183614 259904 -183558
rect 259960 -183614 259968 -183558
rect 259896 -183616 259968 -183614
rect 259902 -183625 259962 -183616
rect 251432 -183830 254488 -183810
rect 258292 -183830 258352 -183821
rect 251432 -183890 254562 -183830
rect 256782 -183832 258352 -183830
rect 256782 -183888 258294 -183832
rect 258350 -183888 258352 -183832
rect 256782 -183890 258352 -183888
rect 251432 -183910 254488 -183890
rect 258292 -183899 258352 -183890
rect 210027 -184558 210145 -184536
rect 210027 -184614 210058 -184558
rect 210114 -184614 210145 -184558
rect 210027 -184636 210145 -184614
rect 173363 -184718 173506 -184705
rect 173138 -184778 173506 -184718
rect 173363 -186046 173506 -184778
rect 253275 -184792 253413 -184760
rect 253275 -184848 253316 -184792
rect 253372 -184848 253413 -184792
rect 253275 -184880 253413 -184848
rect 253284 -184938 253404 -184880
rect 253284 -184998 253882 -184938
rect 253284 -185028 253404 -184998
rect 173359 -186085 173510 -186046
rect 173359 -186141 173406 -186085
rect 173462 -186141 173510 -186085
rect 173359 -186179 173510 -186141
rect 173363 -186183 173506 -186179
rect 298051 -186346 298111 -184146
rect 298042 -186348 298120 -186346
rect 298042 -186404 298053 -186348
rect 298109 -186404 298120 -186348
rect 298042 -186406 298120 -186404
rect 302051 -186638 302111 -184096
rect 302042 -186640 302120 -186638
rect 302042 -186696 302053 -186640
rect 302109 -186696 302120 -186640
rect 302042 -186698 302120 -186696
rect 306051 -186946 306111 -184146
rect 306042 -186948 306120 -186946
rect 306042 -187004 306053 -186948
rect 306109 -187004 306120 -186948
rect 306042 -187006 306120 -187004
rect 310051 -187230 310111 -183946
rect 310042 -187232 310120 -187230
rect 310042 -187288 310053 -187232
rect 310109 -187288 310120 -187232
rect 310042 -187290 310120 -187288
rect 314051 -187526 314111 -184118
rect 314042 -187528 314120 -187526
rect 314042 -187584 314053 -187528
rect 314109 -187584 314120 -187528
rect 314042 -187586 314120 -187584
rect 318051 -187812 318111 -184076
rect 318042 -187814 318120 -187812
rect 318042 -187870 318053 -187814
rect 318109 -187870 318120 -187814
rect 318042 -187872 318120 -187870
rect 326051 -188088 326111 -184090
rect 326042 -188090 326120 -188088
rect 326042 -188146 326053 -188090
rect 326109 -188146 326120 -188090
rect 326042 -188148 326120 -188146
rect 330051 -188382 330111 -184070
rect 333772 -184698 333868 -184692
rect 333763 -184718 333877 -184698
rect 333763 -184774 333792 -184718
rect 333848 -184774 333877 -184718
rect 333763 -184794 333877 -184774
rect 333772 -184800 333868 -184794
rect 334540 -185242 334636 -180328
rect 339830 -182366 339890 -182360
rect 338791 -182368 339890 -182366
rect 338791 -182424 338802 -182368
rect 338858 -182370 339890 -182368
rect 338858 -182422 339834 -182370
rect 339886 -182422 339890 -182370
rect 338858 -182424 339890 -182422
rect 338791 -182426 339890 -182424
rect 339830 -182432 339890 -182426
rect 339574 -184720 339682 -184698
rect 339574 -184772 339602 -184720
rect 339654 -184772 339682 -184720
rect 339574 -184794 339682 -184772
rect 334737 -185028 334880 -184982
rect 334737 -185080 334782 -185028
rect 334834 -185080 334880 -185028
rect 334534 -185264 334642 -185242
rect 334534 -185316 334562 -185264
rect 334614 -185316 334642 -185264
rect 334534 -185338 334642 -185316
rect 333764 -185786 333860 -185780
rect 333755 -185806 333869 -185786
rect 333755 -185862 333784 -185806
rect 333840 -185862 333869 -185806
rect 333755 -185882 333869 -185862
rect 333764 -185888 333860 -185882
rect 334737 -186042 334880 -185080
rect 339580 -185466 339676 -184794
rect 339734 -184896 339794 -184890
rect 340100 -184896 340210 -170714
rect 377783 -170742 377824 -170606
rect 377960 -170742 378001 -170606
rect 377783 -170774 378001 -170742
rect 339734 -184900 340210 -184896
rect 339734 -184952 339738 -184900
rect 339790 -184952 340210 -184900
rect 339734 -184956 340210 -184952
rect 339734 -184962 339794 -184956
rect 334728 -186046 334889 -186042
rect 334728 -186182 334740 -186046
rect 334876 -186182 334889 -186046
rect 334728 -186185 334889 -186182
rect 330042 -188384 330120 -188382
rect 330042 -188440 330053 -188384
rect 330109 -188440 330120 -188384
rect 330042 -188442 330120 -188440
<< via2 >>
rect 196506 -91658 196562 -91602
rect 194342 -92020 194398 -91964
rect 193372 -106014 193428 -106012
rect 193372 -106066 193374 -106014
rect 193374 -106066 193426 -106014
rect 193426 -106066 193428 -106014
rect 193372 -106068 193428 -106066
rect 190398 -108784 190454 -108728
rect 250410 -92392 250466 -92336
rect 266876 -96386 266932 -96330
rect 265988 -96718 266124 -96582
rect 265519 -97918 265655 -97782
rect 262573 -99508 262629 -99452
rect 265046 -101054 265182 -100918
rect 250410 -101292 250466 -101236
rect 198826 -107798 198882 -107742
rect 210634 -108120 210770 -107984
rect 196506 -109440 196562 -109384
rect 191458 -110192 191514 -110136
rect 194518 -110708 194574 -110652
rect 211096 -108350 211152 -108294
rect 196792 -112344 196848 -112288
rect 198512 -112341 198568 -112285
rect 211342 -108664 211398 -108608
rect 210200 -114782 210256 -114726
rect 212378 -109042 212514 -108906
rect 196790 -115308 196846 -115252
rect 211574 -114988 211630 -114932
rect 210546 -115844 210602 -115788
rect 207480 -120918 207536 -120862
rect 207076 -121778 207212 -121642
rect 206556 -122178 206772 -121962
rect 210816 -116944 210872 -116888
rect 195646 -136536 195702 -136480
rect 206010 -137574 206066 -137518
rect 204146 -143718 204202 -143662
rect 204828 -144826 204884 -144770
rect 195646 -149032 195702 -149030
rect 195646 -149084 195648 -149032
rect 195648 -149084 195700 -149032
rect 195700 -149084 195702 -149032
rect 195646 -149086 195702 -149084
rect 245693 -109395 245829 -109259
rect 232511 -109786 232647 -109650
rect 218182 -110284 218318 -110148
rect 212810 -110746 213026 -110530
rect 212418 -121738 212474 -121682
rect 212810 -122178 213026 -121962
rect 205644 -149352 205700 -149296
rect 210274 -155356 210410 -155220
rect 210058 -169662 210114 -169606
rect 186418 -183654 186554 -183518
rect 210274 -170206 210410 -170070
rect 231570 -113924 231626 -113868
rect 225368 -114986 225424 -114930
rect 225378 -115522 225434 -115466
rect 244210 -113924 244266 -113868
rect 264176 -102104 264312 -101968
rect 263746 -105394 263882 -105258
rect 250410 -110652 250466 -110596
rect 250752 -110686 250888 -110550
rect 250350 -111462 250486 -111326
rect 234432 -151526 234488 -151470
rect 250350 -151844 250486 -151708
rect 218182 -155356 218318 -155220
rect 255276 -111084 255412 -110948
rect 264598 -103518 264734 -103382
rect 266440 -100172 266576 -100036
rect 270864 -96746 270920 -96744
rect 270864 -96798 270866 -96746
rect 270866 -96798 270918 -96746
rect 270918 -96798 270920 -96746
rect 270864 -96800 270920 -96798
rect 274294 -96736 274350 -96734
rect 274294 -96788 274296 -96736
rect 274296 -96788 274348 -96736
rect 274348 -96788 274350 -96736
rect 274294 -96790 274350 -96788
rect 268884 -97826 268940 -97824
rect 268884 -97878 268886 -97826
rect 268886 -97878 268938 -97826
rect 268938 -97878 268940 -97826
rect 268884 -97880 268940 -97878
rect 272580 -98022 272636 -98020
rect 272580 -98074 272582 -98022
rect 272582 -98074 272634 -98022
rect 272634 -98074 272636 -98022
rect 272580 -98076 272636 -98074
rect 267512 -98218 267648 -98082
rect 267234 -98444 267290 -98388
rect 274296 -98416 274352 -98360
rect 268445 -99507 268501 -99451
rect 274294 -100230 274350 -100228
rect 274294 -100282 274296 -100230
rect 274296 -100282 274348 -100230
rect 274348 -100282 274350 -100230
rect 274294 -100284 274350 -100282
rect 269026 -100962 269082 -100960
rect 269026 -101014 269028 -100962
rect 269028 -101014 269080 -100962
rect 269080 -101014 269082 -100962
rect 269026 -101016 269082 -101014
rect 268178 -101792 268234 -101736
rect 272580 -101792 272636 -101736
rect 268884 -102056 268940 -102000
rect 274296 -103230 274352 -103228
rect 274296 -103282 274298 -103230
rect 274298 -103282 274350 -103230
rect 274350 -103282 274352 -103230
rect 274296 -103284 274352 -103282
rect 279404 -103676 279540 -103540
rect 295808 -103560 295944 -103424
rect 272582 -105012 272638 -105010
rect 272582 -105064 272584 -105012
rect 272584 -105064 272636 -105012
rect 272636 -105064 272638 -105012
rect 272582 -105066 272638 -105064
rect 276014 -105166 276070 -105110
rect 295850 -105204 295986 -105068
rect 268138 -107542 268274 -107406
rect 276164 -107458 276220 -107402
rect 294226 -107459 294282 -107403
rect 267878 -107798 267934 -107742
rect 275246 -107968 275302 -107966
rect 275246 -108020 275248 -107968
rect 275248 -108020 275300 -107968
rect 275300 -108020 275302 -107968
rect 275246 -108022 275302 -108020
rect 267552 -108080 267608 -108024
rect 267234 -108350 267290 -108294
rect 266876 -108664 266932 -108608
rect 266480 -109002 266536 -108946
rect 265988 -109395 266124 -109259
rect 265519 -109791 265655 -109655
rect 265046 -110284 265182 -110148
rect 264598 -110686 264734 -110550
rect 264176 -111084 264312 -110948
rect 263746 -111462 263882 -111326
rect 294576 -108322 294712 -108186
rect 294576 -122208 294712 -122072
rect 340094 -118562 340230 -118426
rect 297540 -122208 297676 -122072
rect 377160 -118562 377296 -118426
rect 259953 -136256 260089 -136120
rect 294530 -136668 294586 -136612
rect 295260 -136993 295316 -136937
rect 259994 -149036 260050 -149034
rect 259994 -149088 259996 -149036
rect 259996 -149088 260048 -149036
rect 260048 -149088 260050 -149036
rect 259994 -149090 260050 -149088
rect 258312 -149364 258368 -149308
rect 250752 -169408 250888 -169272
rect 227644 -183654 227780 -183518
rect 297138 -127020 297194 -126964
rect 297138 -136668 297194 -136612
rect 298053 -135062 298109 -135006
rect 302053 -135354 302109 -135298
rect 306053 -135662 306109 -135606
rect 310053 -135946 310109 -135890
rect 314053 -136242 314109 -136186
rect 318053 -136528 318109 -136472
rect 326053 -136804 326109 -136748
rect 297487 -136992 297543 -136936
rect 330053 -137098 330109 -137042
rect 334742 -138718 334878 -138582
rect 295260 -150384 295316 -150328
rect 253251 -150471 253307 -150415
rect 255086 -151844 255222 -151708
rect 336268 -137418 336324 -137362
rect 378186 -137498 378322 -137362
rect 336268 -153874 336324 -153818
rect 259866 -170956 260002 -170820
rect 340118 -170714 340174 -170658
rect 294532 -175094 294588 -175038
rect 299040 -178250 299096 -178194
rect 334560 -180328 334616 -180272
rect 259904 -183560 259960 -183558
rect 259904 -183612 259906 -183560
rect 259906 -183612 259958 -183560
rect 259958 -183612 259960 -183560
rect 259904 -183614 259960 -183612
rect 258294 -183888 258350 -183832
rect 210058 -184614 210114 -184558
rect 253316 -184848 253372 -184792
rect 173406 -186141 173462 -186085
rect 298053 -186404 298109 -186348
rect 302053 -186696 302109 -186640
rect 306053 -187004 306109 -186948
rect 310053 -187288 310109 -187232
rect 314053 -187584 314109 -187528
rect 318053 -187870 318109 -187814
rect 326053 -188146 326109 -188090
rect 333792 -184720 333848 -184718
rect 333792 -184772 333794 -184720
rect 333794 -184772 333846 -184720
rect 333846 -184772 333848 -184720
rect 333792 -184774 333848 -184772
rect 338802 -182424 338858 -182368
rect 333784 -185808 333840 -185806
rect 333784 -185860 333786 -185808
rect 333786 -185860 333838 -185808
rect 333838 -185860 333840 -185808
rect 333784 -185862 333840 -185860
rect 377824 -170742 377960 -170606
rect 334740 -186182 334876 -186046
rect 330053 -188440 330109 -188384
<< metal3 >>
rect 196370 -91602 196584 -91580
rect 196370 -91658 196506 -91602
rect 196562 -91658 196584 -91602
rect 196370 -91680 196584 -91658
rect 194320 -91964 194420 -91942
rect 194320 -92020 194342 -91964
rect 194398 -92020 194420 -91964
rect 194320 -92042 194420 -92020
rect 250369 -92336 250507 -92295
rect 250369 -92392 250410 -92336
rect 250466 -92392 250507 -92336
rect 250369 -92433 250507 -92392
rect 200736 -99558 201006 -99458
rect 250374 -101236 250502 -92433
rect 266832 -96295 266976 -96286
rect 266832 -96330 274386 -96295
rect 266832 -96386 266876 -96330
rect 266932 -96386 274386 -96330
rect 266832 -96425 274386 -96386
rect 266832 -96430 266976 -96425
rect 265968 -96580 266144 -96562
rect 265968 -96582 270968 -96580
rect 265968 -96718 265988 -96582
rect 266124 -96718 270968 -96582
rect 265968 -96726 270968 -96718
rect 265968 -96738 266144 -96726
rect 270822 -96744 270968 -96726
rect 270822 -96800 270864 -96744
rect 270920 -96800 270968 -96744
rect 270822 -96826 270968 -96800
rect 274256 -96734 274386 -96425
rect 274256 -96790 274294 -96734
rect 274350 -96790 274386 -96734
rect 274256 -96816 274386 -96790
rect 265475 -97782 265699 -97738
rect 265475 -97918 265519 -97782
rect 265655 -97824 268974 -97782
rect 265655 -97880 268884 -97824
rect 268940 -97880 268974 -97824
rect 265655 -97918 268974 -97880
rect 265475 -97922 268974 -97918
rect 265475 -97962 265699 -97922
rect 272541 -98020 272671 -97995
rect 272541 -98076 272580 -98020
rect 272636 -98076 272671 -98020
rect 267507 -98082 267653 -98077
rect 267507 -98218 267512 -98082
rect 267648 -98086 267653 -98082
rect 272541 -98086 272671 -98076
rect 267648 -98216 272671 -98086
rect 267648 -98218 267653 -98216
rect 267507 -98223 267653 -98218
rect 267194 -98352 267330 -98348
rect 267194 -98353 274356 -98352
rect 267194 -98360 274359 -98353
rect 267194 -98388 274296 -98360
rect 267194 -98444 267234 -98388
rect 267290 -98416 274296 -98388
rect 274352 -98416 274359 -98360
rect 267290 -98423 274359 -98416
rect 267290 -98444 274356 -98423
rect 267194 -98476 274356 -98444
rect 267194 -98484 267330 -98476
rect 262530 -99412 262673 -99408
rect 262530 -99451 268540 -99412
rect 262530 -99452 268445 -99451
rect 262530 -99508 262573 -99452
rect 262629 -99507 268445 -99452
rect 268501 -99507 268540 -99451
rect 262629 -99508 268540 -99507
rect 262530 -99545 268540 -99508
rect 262530 -99551 262673 -99545
rect 266431 -100030 266585 -100027
rect 266431 -100036 274378 -100030
rect 266431 -100172 266440 -100036
rect 266576 -100144 274378 -100036
rect 266576 -100172 266585 -100144
rect 266431 -100181 266585 -100172
rect 274264 -100228 274378 -100144
rect 274264 -100284 274294 -100228
rect 274350 -100284 274378 -100228
rect 274264 -100298 274378 -100284
rect 257354 -100828 257834 -100728
rect 265034 -100914 265194 -100906
rect 265034 -100918 269112 -100914
rect 265034 -101054 265046 -100918
rect 265182 -100960 269112 -100918
rect 265182 -101016 269026 -100960
rect 269082 -101016 269112 -100960
rect 265182 -101054 269112 -101016
rect 265034 -101064 269112 -101054
rect 265034 -101066 265194 -101064
rect 250374 -101292 250410 -101236
rect 250466 -101292 250502 -101236
rect 250374 -101328 250502 -101292
rect 268156 -101736 272660 -101714
rect 268156 -101792 268178 -101736
rect 268234 -101792 272580 -101736
rect 272636 -101792 272660 -101736
rect 268156 -101814 272660 -101792
rect 264166 -101962 264322 -101958
rect 264166 -101968 268970 -101962
rect 264166 -102104 264176 -101968
rect 264312 -102000 268970 -101968
rect 264312 -102056 268884 -102000
rect 268940 -102056 268970 -102000
rect 264312 -102104 268970 -102056
rect 264166 -102110 268970 -102104
rect 264166 -102114 264322 -102110
rect 274254 -103228 274400 -103192
rect 274254 -103284 274296 -103228
rect 274352 -103284 274400 -103228
rect 264582 -103375 264750 -103366
rect 274254 -103375 274400 -103284
rect 264582 -103382 274400 -103375
rect 264582 -103518 264598 -103382
rect 264734 -103518 274400 -103382
rect 295791 -103412 295961 -103407
rect 264582 -103521 274400 -103518
rect 279392 -103424 295961 -103412
rect 264582 -103534 264750 -103521
rect 279392 -103540 295808 -103424
rect 279392 -103676 279404 -103540
rect 279540 -103560 295808 -103540
rect 295944 -103560 295961 -103424
rect 279540 -103572 295961 -103560
rect 279540 -103676 279552 -103572
rect 295791 -103577 295961 -103572
rect 279392 -103688 279552 -103676
rect 272530 -105010 272686 -104986
rect 272530 -105066 272582 -105010
rect 272638 -105066 272686 -105010
rect 263729 -105250 263899 -105241
rect 272530 -105250 272686 -105066
rect 275988 -105068 295992 -105062
rect 275988 -105110 295850 -105068
rect 275988 -105166 276014 -105110
rect 276070 -105166 295850 -105110
rect 275988 -105204 295850 -105166
rect 295986 -105204 295992 -105068
rect 275988 -105210 295992 -105204
rect 257776 -105356 258178 -105256
rect 263729 -105258 272686 -105250
rect 263729 -105394 263746 -105258
rect 263882 -105394 272686 -105258
rect 263729 -105406 272686 -105394
rect 263729 -105411 263899 -105406
rect 193330 -106012 197124 -105970
rect 193330 -106068 193372 -106012
rect 193428 -106068 197124 -106012
rect 193330 -106110 197124 -106068
rect 196984 -107404 197124 -106110
rect 268131 -107404 268281 -107399
rect 196984 -107406 268281 -107404
rect 196984 -107542 268138 -107406
rect 268274 -107542 268281 -107406
rect 276138 -107402 294325 -107360
rect 276138 -107458 276164 -107402
rect 276220 -107403 294325 -107402
rect 276220 -107458 294226 -107403
rect 276138 -107459 294226 -107458
rect 294282 -107459 294325 -107403
rect 276138 -107502 294325 -107459
rect 196984 -107544 268281 -107542
rect 268131 -107549 268281 -107544
rect 198784 -107705 198924 -107700
rect 198784 -107742 267971 -107705
rect 198784 -107798 198826 -107742
rect 198882 -107798 267878 -107742
rect 267934 -107798 267971 -107742
rect 198784 -107835 267971 -107798
rect 198784 -107840 198924 -107835
rect 275204 -107966 275350 -107944
rect 210629 -107984 210775 -107979
rect 210629 -108120 210634 -107984
rect 210770 -108024 267648 -107984
rect 210770 -108080 267552 -108024
rect 267608 -108080 267648 -108024
rect 210770 -108120 267648 -108080
rect 275204 -108022 275246 -107966
rect 275302 -108022 275350 -107966
rect 210629 -108125 210775 -108120
rect 275204 -108181 275350 -108022
rect 275204 -108186 294717 -108181
rect 211056 -108259 211192 -108254
rect 211056 -108294 267325 -108259
rect 211056 -108350 211096 -108294
rect 211152 -108350 267234 -108294
rect 267290 -108350 267325 -108294
rect 275204 -108322 294576 -108186
rect 294712 -108322 294717 -108186
rect 275204 -108327 294717 -108322
rect 211056 -108385 267325 -108350
rect 211056 -108390 211192 -108385
rect 211298 -108569 211442 -108564
rect 211298 -108608 266971 -108569
rect 211298 -108664 211342 -108608
rect 211398 -108664 266876 -108608
rect 266932 -108664 266971 -108608
rect 211298 -108703 266971 -108664
rect 190376 -108728 190476 -108706
rect 211298 -108708 211442 -108703
rect 190376 -108784 190398 -108728
rect 190454 -108784 190476 -108728
rect 190376 -110116 190476 -108784
rect 212369 -108902 212523 -108897
rect 212369 -108906 266580 -108902
rect 212369 -109042 212378 -108906
rect 212514 -108946 266580 -108906
rect 212514 -109002 266480 -108946
rect 266536 -109002 266580 -108946
rect 212514 -109042 266580 -109002
rect 212369 -109046 266580 -109042
rect 212369 -109051 212523 -109046
rect 245673 -109244 245849 -109239
rect 245673 -109259 266139 -109244
rect 196484 -109384 196584 -109362
rect 196484 -109440 196506 -109384
rect 196562 -109440 196584 -109384
rect 245673 -109395 245693 -109259
rect 245829 -109395 265988 -109259
rect 266124 -109395 266139 -109259
rect 245673 -109410 266139 -109395
rect 245673 -109415 245849 -109410
rect 196484 -110116 196584 -109440
rect 232508 -109644 265694 -109616
rect 232505 -109650 265694 -109644
rect 232505 -109786 232511 -109650
rect 232647 -109655 265694 -109650
rect 232647 -109786 265519 -109655
rect 232505 -109791 265519 -109786
rect 265655 -109791 265694 -109655
rect 232505 -109792 265694 -109791
rect 232508 -109830 265694 -109792
rect 190376 -110136 191542 -110116
rect 190376 -110192 191458 -110136
rect 191514 -110192 191542 -110136
rect 190376 -110216 191542 -110192
rect 194496 -110216 196584 -110116
rect 218170 -110141 218330 -110136
rect 218170 -110148 265189 -110141
rect 194496 -110652 194596 -110216
rect 218170 -110284 218182 -110148
rect 218318 -110284 265046 -110148
rect 265182 -110284 265189 -110148
rect 218170 -110291 265189 -110284
rect 218170 -110296 218330 -110291
rect 194496 -110708 194518 -110652
rect 194574 -110708 194596 -110652
rect 194496 -110732 194596 -110708
rect 212802 -110530 250536 -110522
rect 212802 -110746 212810 -110530
rect 213026 -110596 250536 -110530
rect 213026 -110652 250410 -110596
rect 250466 -110652 250536 -110596
rect 213026 -110746 250536 -110652
rect 250736 -110539 250904 -110534
rect 250736 -110550 264745 -110539
rect 250736 -110686 250752 -110550
rect 250888 -110686 264598 -110550
rect 264734 -110686 264745 -110550
rect 250736 -110697 264745 -110686
rect 250736 -110702 250904 -110697
rect 212802 -110754 250536 -110746
rect 255266 -110943 255422 -110938
rect 255266 -110948 264317 -110943
rect 255266 -111084 255276 -110948
rect 255412 -111084 264176 -110948
rect 264312 -111084 264317 -110948
rect 255266 -111089 264317 -111084
rect 255266 -111094 255422 -111089
rect 336284 -111122 336606 -111022
rect 250333 -111314 250503 -111309
rect 250333 -111326 263894 -111314
rect 250333 -111462 250350 -111326
rect 250486 -111462 263746 -111326
rect 263882 -111462 263894 -111326
rect 250333 -111474 263894 -111462
rect 250333 -111479 250503 -111474
rect 186620 -111908 186720 -111614
rect 186882 -111772 186982 -111506
rect 196756 -112285 198605 -112248
rect 196756 -112288 198512 -112285
rect 196756 -112344 196792 -112288
rect 196848 -112341 198512 -112288
rect 198568 -112341 198605 -112285
rect 196848 -112344 198605 -112341
rect 196756 -112378 198605 -112344
rect 231546 -113868 244288 -113846
rect 231546 -113924 231570 -113868
rect 231626 -113924 244210 -113868
rect 244266 -113924 244288 -113868
rect 231546 -113946 244288 -113924
rect 199111 -114726 210291 -114691
rect 199111 -114782 210200 -114726
rect 210256 -114782 210291 -114726
rect 199111 -114817 210291 -114782
rect 199111 -115218 199237 -114817
rect 211552 -114930 225442 -114910
rect 211552 -114932 225368 -114930
rect 211552 -114988 211574 -114932
rect 211630 -114986 225368 -114932
rect 225424 -114986 225442 -114930
rect 211630 -114988 225442 -114986
rect 211552 -115010 225442 -114988
rect 196754 -115252 199237 -115218
rect 196754 -115308 196790 -115252
rect 196846 -115308 199237 -115252
rect 196754 -115344 199237 -115308
rect 210808 -115466 225456 -115442
rect 210808 -115522 225378 -115466
rect 225434 -115522 225456 -115466
rect 210808 -115542 225456 -115522
rect 210524 -115788 210624 -115644
rect 210524 -115844 210546 -115788
rect 210602 -115844 210624 -115788
rect 210524 -115866 210624 -115844
rect 206496 -117378 206596 -116016
rect 210794 -116888 210894 -116692
rect 210794 -116944 210816 -116888
rect 210872 -116944 210894 -116888
rect 210794 -116966 210894 -116944
rect 206496 -117478 207558 -117378
rect 207458 -120862 207558 -117478
rect 340084 -118421 340240 -118416
rect 340084 -118426 377301 -118421
rect 340084 -118562 340094 -118426
rect 340230 -118562 377160 -118426
rect 377296 -118562 377301 -118426
rect 340084 -118567 377301 -118562
rect 340084 -118572 340240 -118567
rect 338785 -119638 338885 -119002
rect 207458 -120918 207480 -120862
rect 207536 -120918 207558 -120862
rect 207458 -120940 207558 -120918
rect 207067 -121638 207221 -121633
rect 207067 -121642 212518 -121638
rect 207067 -121778 207076 -121642
rect 207212 -121682 212518 -121642
rect 207212 -121738 212418 -121682
rect 212474 -121738 212518 -121682
rect 207212 -121778 212518 -121738
rect 207067 -121782 212518 -121778
rect 207067 -121787 207221 -121782
rect 212797 -121954 213039 -121949
rect 206548 -121962 213039 -121954
rect 206548 -122178 206556 -121962
rect 206772 -122178 212810 -121962
rect 213026 -122178 213039 -121962
rect 206548 -122186 213039 -122178
rect 212797 -122191 213039 -122186
rect 294566 -122067 294722 -122062
rect 294566 -122072 297681 -122067
rect 294566 -122208 294576 -122072
rect 294712 -122208 297540 -122072
rect 297676 -122208 297681 -122072
rect 294566 -122213 297681 -122208
rect 294566 -122218 294722 -122213
rect 338785 -124498 338885 -123906
rect 338785 -124562 338803 -124498
rect 338867 -124562 338885 -124498
rect 338785 -124586 338885 -124562
rect 297116 -126964 298230 -126942
rect 297116 -127020 297138 -126964
rect 297194 -127020 298230 -126964
rect 297116 -127042 298230 -127020
rect 297550 -132004 297938 -131904
rect 297746 -133988 298290 -133888
rect 298030 -135006 336458 -134982
rect 298030 -135062 298053 -135006
rect 298109 -135062 336458 -135006
rect 298030 -135082 336458 -135062
rect 302028 -135298 336456 -135274
rect 302028 -135354 302053 -135298
rect 302109 -135354 336456 -135298
rect 302028 -135374 336456 -135354
rect 306032 -135606 336464 -135584
rect 306032 -135662 306053 -135606
rect 306109 -135662 336464 -135606
rect 306032 -135684 336464 -135662
rect 310030 -135890 336472 -135868
rect 310030 -135946 310053 -135890
rect 310109 -135946 336472 -135890
rect 310030 -135968 336472 -135946
rect 259948 -136120 260094 -136115
rect 259948 -136256 259953 -136120
rect 260089 -136256 260094 -136120
rect 195602 -136480 195746 -136436
rect 195602 -136536 195646 -136480
rect 195702 -136536 195746 -136480
rect 195602 -149030 195746 -136536
rect 203960 -137518 206088 -137496
rect 203960 -137574 206010 -137518
rect 206066 -137574 206088 -137518
rect 203960 -137596 206088 -137574
rect 204124 -143641 204224 -143640
rect 204119 -143658 204229 -143641
rect 204119 -143722 204142 -143658
rect 204206 -143722 204229 -143658
rect 204119 -143739 204229 -143722
rect 204124 -143740 204224 -143739
rect 204348 -144770 204906 -144748
rect 204348 -144826 204828 -144770
rect 204884 -144826 204906 -144770
rect 204348 -144848 204906 -144826
rect 195602 -149086 195646 -149030
rect 195702 -149086 195746 -149030
rect 195602 -149116 195746 -149086
rect 259948 -149034 260094 -136256
rect 314026 -136186 336470 -136166
rect 314026 -136242 314053 -136186
rect 314109 -136242 336470 -136186
rect 314026 -136266 336470 -136242
rect 318028 -136472 336472 -136448
rect 318028 -136528 318053 -136472
rect 318109 -136528 336472 -136472
rect 318028 -136548 336472 -136528
rect 297111 -136590 297221 -136585
rect 294508 -136612 297221 -136590
rect 294508 -136668 294530 -136612
rect 294586 -136668 297138 -136612
rect 297194 -136668 297221 -136612
rect 294508 -136690 297221 -136668
rect 297111 -136695 297221 -136690
rect 326026 -136748 336488 -136726
rect 326026 -136804 326053 -136748
rect 326109 -136804 336488 -136748
rect 326026 -136826 336488 -136804
rect 295225 -136905 295352 -136901
rect 295225 -136936 297574 -136905
rect 295225 -136937 297487 -136936
rect 295225 -136993 295260 -136937
rect 295316 -136992 297487 -136937
rect 297543 -136992 297574 -136936
rect 295316 -136993 297574 -136992
rect 295225 -137022 297574 -136993
rect 295225 -137028 295352 -137022
rect 330026 -137042 336500 -137020
rect 330026 -137098 330053 -137042
rect 330109 -137098 336500 -137042
rect 330026 -137120 336500 -137098
rect 336241 -137342 336351 -137335
rect 338786 -137342 338884 -137337
rect 336241 -137360 338885 -137342
rect 378166 -137347 378342 -137342
rect 336241 -137362 338803 -137360
rect 336241 -137418 336268 -137362
rect 336324 -137418 338803 -137362
rect 336241 -137424 338803 -137418
rect 338867 -137424 338885 -137360
rect 336241 -137442 338885 -137424
rect 351353 -137362 378342 -137347
rect 336241 -137445 336351 -137442
rect 338786 -137447 338884 -137442
rect 351353 -137498 378186 -137362
rect 378322 -137498 378342 -137362
rect 351353 -137513 378342 -137498
rect 351353 -138567 351519 -137513
rect 378166 -137518 378342 -137513
rect 334727 -138582 351519 -138567
rect 334727 -138718 334742 -138582
rect 334878 -138718 351519 -138582
rect 334727 -138733 351519 -138718
rect 259948 -149090 259994 -149034
rect 260050 -149090 260094 -149034
rect 259948 -149118 260094 -149090
rect 203784 -149296 205722 -149274
rect 203784 -149352 205644 -149296
rect 205700 -149352 205722 -149296
rect 203784 -149374 205722 -149352
rect 258292 -149308 258409 -149262
rect 258292 -149364 258312 -149308
rect 258368 -149364 258409 -149308
rect 258292 -150296 258409 -149364
rect 295225 -150296 295352 -150292
rect 258292 -150328 295352 -150296
rect 253218 -150415 253341 -150381
rect 258292 -150384 295260 -150328
rect 295316 -150384 295352 -150328
rect 258292 -150413 295352 -150384
rect 253218 -150471 253251 -150415
rect 253307 -150471 253341 -150415
rect 295225 -150419 295352 -150413
rect 234394 -151435 234527 -151431
rect 253218 -151435 253341 -150471
rect 234394 -151470 253341 -151435
rect 234394 -151526 234432 -151470
rect 234488 -151526 253341 -151470
rect 234394 -151558 253341 -151526
rect 234394 -151564 234527 -151558
rect 255069 -151696 255239 -151691
rect 250338 -151708 255239 -151696
rect 250338 -151844 250350 -151708
rect 250486 -151844 255086 -151708
rect 255222 -151844 255239 -151708
rect 250338 -151856 255239 -151844
rect 255069 -151861 255239 -151856
rect 336246 -153818 336346 -153796
rect 336246 -153874 336268 -153818
rect 336324 -153874 336346 -153818
rect 210262 -155213 210422 -155208
rect 210262 -155220 218325 -155213
rect 210262 -155356 210274 -155220
rect 210410 -155356 218182 -155220
rect 218318 -155356 218325 -155220
rect 210262 -155363 218325 -155356
rect 210262 -155368 210422 -155363
rect 336246 -161489 336346 -153874
rect 336241 -161506 336351 -161489
rect 336241 -161570 336264 -161506
rect 336328 -161570 336351 -161506
rect 336241 -161587 336351 -161570
rect 336246 -161588 336346 -161587
rect 336364 -162132 336720 -162032
rect 338785 -166646 338885 -166622
rect 338785 -166710 338803 -166646
rect 338867 -166710 338885 -166646
rect 338785 -167752 338885 -166710
rect 227633 -169272 250899 -169261
rect 227633 -169408 250752 -169272
rect 250888 -169408 250899 -169272
rect 227633 -169419 250899 -169408
rect 187545 -169584 187643 -169579
rect 187544 -169602 210136 -169584
rect 187544 -169666 187562 -169602
rect 187626 -169606 210136 -169602
rect 187626 -169662 210058 -169606
rect 210114 -169662 210136 -169606
rect 187626 -169666 210136 -169662
rect 187544 -169684 210136 -169666
rect 187545 -169689 187643 -169684
rect 186411 -170070 210417 -170063
rect 186411 -170206 210274 -170070
rect 210410 -170206 210417 -170070
rect 186411 -170213 210417 -170206
rect 186411 -183506 186561 -170213
rect 227633 -183502 227791 -169419
rect 377787 -170574 377997 -170569
rect 340092 -170606 377997 -170574
rect 340092 -170658 377824 -170606
rect 340092 -170714 340118 -170658
rect 340174 -170714 377824 -170658
rect 340092 -170742 377824 -170714
rect 377960 -170742 377997 -170606
rect 340092 -170774 377997 -170742
rect 377787 -170779 377997 -170774
rect 259849 -170820 260019 -170803
rect 259849 -170956 259866 -170820
rect 260002 -170956 260019 -170820
rect 259849 -170973 260019 -170956
rect 186406 -183518 186566 -183506
rect 186406 -183654 186418 -183518
rect 186554 -183654 186566 -183518
rect 186406 -183666 186566 -183654
rect 227628 -183518 227796 -183502
rect 227628 -183654 227644 -183518
rect 227780 -183654 227796 -183518
rect 259854 -183558 260014 -170973
rect 294506 -175038 295272 -175012
rect 294506 -175094 294532 -175038
rect 294588 -175094 295272 -175038
rect 294506 -175112 295272 -175094
rect 295172 -177952 295272 -175112
rect 295172 -178052 298374 -177952
rect 259854 -183614 259904 -183558
rect 259960 -183614 260014 -183558
rect 259854 -183646 260014 -183614
rect 296002 -178194 299114 -178170
rect 296002 -178250 299040 -178194
rect 299096 -178250 299114 -178194
rect 296002 -178270 299114 -178250
rect 227628 -183670 227796 -183654
rect 258272 -183832 258372 -183802
rect 258272 -183888 258294 -183832
rect 258350 -183888 258372 -183832
rect 210031 -184536 210141 -184531
rect 210031 -184558 211630 -184536
rect 210031 -184614 210058 -184558
rect 210114 -184614 211630 -184558
rect 210031 -184636 211630 -184614
rect 210031 -184641 210141 -184636
rect 211530 -184760 211630 -184636
rect 253279 -184760 253409 -184755
rect 211530 -184792 253409 -184760
rect 211530 -184848 253316 -184792
rect 253372 -184848 253409 -184792
rect 211530 -184880 253409 -184848
rect 253279 -184885 253409 -184880
rect 258272 -184818 258372 -183888
rect 296002 -184818 296102 -178270
rect 334535 -180263 334641 -180241
rect 334535 -180327 334556 -180263
rect 334620 -180327 334641 -180263
rect 334535 -180328 334560 -180327
rect 334616 -180328 334641 -180327
rect 334535 -180353 334641 -180328
rect 338785 -182368 338885 -175208
rect 338785 -182424 338802 -182368
rect 338858 -182424 338885 -182368
rect 338785 -182438 338885 -182424
rect 297634 -183014 298016 -182914
rect 333761 -184714 333873 -184693
rect 333761 -184778 333783 -184714
rect 333847 -184718 333873 -184714
rect 333848 -184774 333873 -184718
rect 333847 -184778 333873 -184774
rect 333761 -184799 333873 -184778
rect 258272 -184918 296102 -184818
rect 297882 -184998 298348 -184898
rect 333753 -185802 333865 -185781
rect 333753 -185866 333775 -185802
rect 333839 -185806 333865 -185802
rect 333840 -185862 333865 -185806
rect 333839 -185866 333865 -185862
rect 333753 -185887 333865 -185866
rect 334732 -186041 334885 -186037
rect 173363 -186046 334885 -186041
rect 173363 -186085 334740 -186046
rect 173363 -186141 173406 -186085
rect 173462 -186141 334740 -186085
rect 173363 -186182 334740 -186141
rect 334876 -186182 334885 -186046
rect 173363 -186184 334885 -186182
rect 334732 -186190 334885 -186184
rect 298030 -186348 336458 -186324
rect 298030 -186404 298053 -186348
rect 298109 -186404 336458 -186348
rect 298030 -186424 336458 -186404
rect 302028 -186640 336456 -186616
rect 302028 -186696 302053 -186640
rect 302109 -186696 336456 -186640
rect 302028 -186716 336456 -186696
rect 306032 -186948 336464 -186926
rect 306032 -187004 306053 -186948
rect 306109 -187004 336464 -186948
rect 306032 -187026 336464 -187004
rect 310030 -187232 336472 -187210
rect 310030 -187288 310053 -187232
rect 310109 -187288 336472 -187232
rect 310030 -187310 336472 -187288
rect 314026 -187528 336470 -187508
rect 314026 -187584 314053 -187528
rect 314109 -187584 336470 -187528
rect 314026 -187608 336470 -187584
rect 318028 -187814 336472 -187790
rect 318028 -187870 318053 -187814
rect 318109 -187870 336472 -187814
rect 318028 -187890 336472 -187870
rect 326026 -188090 336488 -188068
rect 326026 -188146 326053 -188090
rect 326109 -188146 336488 -188090
rect 326026 -188168 336488 -188146
rect 330026 -188384 336500 -188362
rect 330026 -188440 330053 -188384
rect 330109 -188440 336500 -188384
rect 330026 -188462 336500 -188440
<< via3 >>
rect 338803 -124562 338867 -124498
rect 204142 -143662 204206 -143658
rect 204142 -143718 204146 -143662
rect 204146 -143718 204202 -143662
rect 204202 -143718 204206 -143662
rect 204142 -143722 204206 -143718
rect 338803 -137424 338867 -137360
rect 336264 -161570 336328 -161506
rect 338803 -166710 338867 -166646
rect 187562 -169666 187626 -169602
rect 334556 -180272 334620 -180263
rect 334556 -180327 334560 -180272
rect 334560 -180327 334616 -180272
rect 334616 -180327 334620 -180272
rect 333783 -184718 333847 -184714
rect 333783 -184774 333792 -184718
rect 333792 -184774 333847 -184718
rect 333783 -184778 333847 -184774
rect 333775 -185806 333839 -185802
rect 333775 -185862 333784 -185806
rect 333784 -185862 333839 -185806
rect 333775 -185866 333839 -185862
<< metal4 >>
rect 157844 -78474 160852 -78352
rect 157844 -79030 157966 -78474
rect 158522 -79030 160852 -78474
rect 157844 -79152 160852 -79030
rect 247146 -78462 296782 -78340
rect 247146 -79018 296104 -78462
rect 296660 -79018 296782 -78462
rect 247146 -79140 296782 -79018
rect 280914 -95428 296776 -95306
rect 280914 -95984 296098 -95428
rect 296654 -95984 296776 -95428
rect 280914 -96106 296776 -95984
rect 211286 -106662 212086 -106540
rect 211286 -107218 211408 -106662
rect 211964 -107218 212086 -106662
rect 211286 -107340 212086 -107218
rect 250952 -106662 251704 -106564
rect 250952 -107218 251050 -106662
rect 251606 -107218 251704 -106662
rect 250952 -107316 251704 -107218
rect 258602 -107340 269368 -106540
rect 157844 -108302 187308 -108180
rect 157844 -108858 157966 -108302
rect 158522 -108858 187308 -108302
rect 157844 -108980 187308 -108858
rect 268534 -109174 269368 -107340
rect 268534 -109208 269334 -109174
rect 229772 -112180 236238 -111508
rect 208338 -113518 212086 -113396
rect 208338 -114074 211408 -113518
rect 211964 -114074 212086 -113518
rect 208338 -114196 212086 -114074
rect 225610 -118458 236324 -117514
rect 342116 -117540 385656 -117418
rect 342116 -118096 384978 -117540
rect 385534 -118096 385656 -117540
rect 342116 -118218 385656 -118096
rect 247830 -118396 251770 -118274
rect 190842 -118921 210439 -118846
rect 190842 -118958 208848 -118921
rect 185684 -119838 208848 -118958
rect 185684 -120184 185806 -119838
rect 185708 -120394 185806 -120184
rect 186362 -120184 208848 -119838
rect 186362 -120394 186460 -120184
rect 185708 -120492 186460 -120394
rect 190842 -120437 208848 -120184
rect 210364 -120437 210439 -118921
rect 247830 -118952 251092 -118396
rect 251648 -118952 251770 -118396
rect 247830 -119074 251770 -118952
rect 190842 -120512 210439 -120437
rect 249252 -119838 256954 -119716
rect 249252 -120394 249374 -119838
rect 249930 -120394 256954 -119838
rect 249252 -120516 256954 -120394
rect 293920 -119838 296780 -119716
rect 293920 -120394 296102 -119838
rect 296658 -120394 296780 -119838
rect 293920 -120516 296780 -120394
rect 296080 -123454 302270 -123388
rect 208547 -123749 222055 -123602
rect 208547 -125265 208694 -123749
rect 210210 -125265 222055 -123749
rect 296080 -124010 296146 -123454
rect 296702 -124010 302270 -123454
rect 296080 -124076 302270 -124010
rect 338784 -124498 338886 -124479
rect 338784 -124562 338803 -124498
rect 338867 -124562 338886 -124498
rect 338784 -124581 338886 -124562
rect 208547 -125412 222055 -125265
rect 294496 -128878 302212 -128756
rect 294496 -129434 294618 -128878
rect 295174 -129434 302212 -128878
rect 294496 -129556 302212 -129434
rect 296088 -134266 301586 -134200
rect 296088 -134822 296154 -134266
rect 296710 -134822 301586 -134266
rect 296088 -134888 301586 -134822
rect 338785 -137360 338885 -124581
rect 338785 -137424 338803 -137360
rect 338867 -137424 338885 -137360
rect 338785 -137442 338885 -137424
rect 208535 -141545 221791 -141512
rect 204124 -143658 204224 -141788
rect 208535 -143381 208568 -141545
rect 210404 -143381 221791 -141545
rect 208535 -143414 221791 -143381
rect 204124 -143722 204142 -143658
rect 204206 -143722 204224 -143658
rect 204124 -143740 204224 -143722
rect 200065 -151312 221000 -150512
rect 247926 -150636 261544 -150516
rect 247926 -151192 251050 -150636
rect 251606 -151192 261544 -150636
rect 247926 -151316 261544 -151192
rect 294520 -150668 295272 -150570
rect 294520 -151224 294618 -150668
rect 295174 -151224 295272 -150668
rect 294520 -151322 295272 -151224
rect 380500 -153356 385652 -153234
rect 380500 -153912 384974 -153356
rect 385530 -153912 385652 -153356
rect 380500 -154034 385652 -153912
rect 249184 -154376 256746 -154240
rect 249184 -154932 249398 -154376
rect 249954 -154932 256746 -154376
rect 249184 -155040 256746 -154932
rect 293878 -154362 296776 -154240
rect 293878 -154918 296098 -154362
rect 296654 -154918 296776 -154362
rect 293878 -155040 296776 -154918
rect 336246 -161506 338885 -161488
rect 336246 -161570 336264 -161506
rect 336328 -161570 338885 -161506
rect 336246 -161588 338885 -161570
rect 338785 -166627 338885 -161588
rect 338784 -166646 338886 -166627
rect 338784 -166710 338803 -166646
rect 338867 -166710 338886 -166646
rect 338784 -166729 338886 -166710
rect 186884 -169602 187644 -169584
rect 186884 -169666 187562 -169602
rect 187626 -169666 187644 -169602
rect 186884 -169684 187644 -169666
rect 296088 -174464 301464 -174398
rect 296088 -175020 296154 -174464
rect 296710 -175020 301464 -174464
rect 296088 -175086 301464 -175020
rect 296598 -179888 302070 -179766
rect 296598 -180444 296720 -179888
rect 297276 -180444 302070 -179888
rect 334534 -180263 334642 -180246
rect 334534 -180327 334556 -180263
rect 334620 -180327 334642 -180263
rect 334534 -180344 334642 -180327
rect 296598 -180566 302070 -180444
rect 333766 -184714 333864 -184692
rect 333766 -184778 333783 -184714
rect 333847 -184778 333864 -184714
rect 333766 -184800 333864 -184778
rect 247432 -185162 258624 -185040
rect 247432 -185718 251050 -185162
rect 251606 -185718 258624 -185162
rect 247432 -185840 258624 -185718
rect 295308 -185158 297398 -185036
rect 295308 -185714 296720 -185158
rect 297276 -185714 297398 -185158
rect 295308 -185836 297398 -185714
rect 333758 -185802 333856 -185780
rect 333758 -185866 333775 -185802
rect 333839 -185866 333856 -185802
rect 333758 -185888 333856 -185866
<< via4 >>
rect 157966 -79030 158522 -78474
rect 296104 -79018 296660 -78462
rect 296098 -95984 296654 -95428
rect 211408 -107218 211964 -106662
rect 251050 -107218 251606 -106662
rect 157966 -108858 158522 -108302
rect 211408 -114074 211964 -113518
rect 384978 -118096 385534 -117540
rect 185806 -120394 186362 -119838
rect 208848 -120437 210364 -118921
rect 251092 -118952 251648 -118396
rect 249374 -120394 249930 -119838
rect 296102 -120394 296658 -119838
rect 208694 -125265 210210 -123749
rect 296146 -124010 296702 -123454
rect 294618 -129434 295174 -128878
rect 296154 -134822 296710 -134266
rect 208568 -143381 210404 -141545
rect 251050 -151192 251606 -150636
rect 294618 -151224 295174 -150668
rect 384974 -153912 385530 -153356
rect 249398 -154932 249954 -154376
rect 296098 -154918 296654 -154362
rect 296154 -175020 296710 -174464
rect 296720 -180444 297276 -179888
rect 251050 -185718 251606 -185162
rect 296720 -185714 297276 -185158
<< metal5 >>
rect 296088 -78316 296776 -78314
rect 157844 -78474 158644 -78352
rect 157844 -79030 157966 -78474
rect 158522 -79030 158644 -78474
rect 157844 -108156 158644 -79030
rect 295958 -78462 296806 -78316
rect 295958 -79018 296104 -78462
rect 296660 -79018 296806 -78462
rect 295958 -79164 296806 -79018
rect 296088 -95282 296776 -79164
rect 295952 -95428 296800 -95282
rect 295952 -95984 296098 -95428
rect 296654 -95984 296800 -95428
rect 295952 -96130 296800 -95984
rect 211262 -106662 212110 -106516
rect 211262 -107218 211408 -106662
rect 211964 -107218 212110 -106662
rect 211262 -107364 212110 -107218
rect 250928 -106662 251728 -106540
rect 250928 -107218 251050 -106662
rect 251606 -107218 251728 -106662
rect 157820 -108302 158668 -108156
rect 157820 -108858 157966 -108302
rect 158522 -108858 158668 -108302
rect 157820 -109004 158668 -108858
rect 211286 -113518 212086 -107364
rect 211286 -114074 211408 -113518
rect 211964 -114074 212086 -113518
rect 211286 -114196 212086 -114074
rect 185684 -119838 186484 -117842
rect 250928 -118250 251728 -107218
rect 250928 -118396 251794 -118250
rect 185684 -120394 185806 -119838
rect 186362 -120394 186484 -119838
rect 185684 -120516 186484 -120394
rect 208535 -118822 210437 -118641
rect 208535 -118921 210463 -118822
rect 208535 -120437 208848 -118921
rect 210364 -120437 210463 -118921
rect 250928 -118952 251092 -118396
rect 251648 -118952 251794 -118396
rect 250928 -119098 251794 -118952
rect 208535 -120536 210463 -120437
rect 249228 -119838 250076 -119692
rect 249228 -120394 249374 -119838
rect 249930 -120394 250076 -119838
rect 208535 -123578 210437 -120536
rect 249228 -120540 250076 -120394
rect 208523 -123749 210437 -123578
rect 208523 -125265 208694 -123749
rect 210210 -125265 210437 -123749
rect 208523 -125436 210437 -125265
rect 208535 -141488 210437 -125436
rect 250928 -135242 251728 -119098
rect 296088 -119692 296776 -96130
rect 384832 -117540 385680 -117394
rect 384832 -118096 384978 -117540
rect 385534 -118096 385680 -117540
rect 384832 -118242 385680 -118096
rect 295956 -119838 296804 -119692
rect 295956 -120394 296102 -119838
rect 296658 -120394 296804 -119838
rect 295956 -120540 296804 -120394
rect 296088 -123364 296776 -120540
rect 296056 -123454 296792 -123364
rect 296056 -124010 296146 -123454
rect 296702 -124010 296792 -123454
rect 296056 -124100 296792 -124010
rect 294472 -128878 295320 -128732
rect 294472 -129434 294618 -128878
rect 295174 -129434 295320 -128878
rect 294472 -129580 295320 -129434
rect 250928 -136042 256670 -135242
rect 208511 -141545 210461 -141488
rect 208511 -143381 208568 -141545
rect 210404 -143381 210461 -141545
rect 208511 -143438 210461 -143381
rect 249276 -154376 250076 -149618
rect 249276 -154932 249398 -154376
rect 249954 -154932 250076 -154376
rect 249276 -155054 250076 -154932
rect 250928 -150636 251728 -136042
rect 250928 -151192 251050 -150636
rect 251606 -151192 251728 -150636
rect 250928 -185016 251728 -151192
rect 294496 -150668 295296 -129580
rect 296088 -134176 296776 -124100
rect 296064 -134266 296800 -134176
rect 296064 -134822 296154 -134266
rect 296710 -134822 296800 -134266
rect 296064 -134912 296800 -134822
rect 294496 -151224 294618 -150668
rect 295174 -151224 295296 -150668
rect 294496 -151346 295296 -151224
rect 296088 -154216 296776 -134912
rect 335069 -139430 335869 -122300
rect 384852 -153210 385652 -118242
rect 384828 -153356 385676 -153210
rect 384828 -153912 384974 -153356
rect 385530 -153912 385676 -153356
rect 384828 -154058 385676 -153912
rect 295952 -154362 296800 -154216
rect 295952 -154918 296098 -154362
rect 296654 -154918 296800 -154362
rect 295952 -155064 296800 -154918
rect 296088 -174374 296776 -155064
rect 296064 -174464 296800 -174374
rect 296064 -175020 296154 -174464
rect 296710 -175020 296800 -174464
rect 296064 -175110 296800 -175020
rect 296574 -179888 297422 -179742
rect 296574 -180444 296720 -179888
rect 297276 -180444 297422 -179888
rect 296574 -180590 297422 -180444
rect 250904 -185162 251752 -185016
rect 250904 -185718 251050 -185162
rect 251606 -185718 251752 -185162
rect 250904 -185864 251752 -185718
rect 296598 -185158 297398 -180590
rect 296598 -185714 296720 -185158
rect 297276 -185714 297398 -185158
rect 296598 -185836 297398 -185714
use comparator  comparator_0
timestamp 1626065694
transform 1 0 229012 0 1 -114708
box -3400 -3600 3400 3200
use sample_and_hold  sample_and_hold_0
timestamp 1626065694
transform 1 0 253730 0 1 -183720
box -1766 -2168 42040 29538
use sample_and_hold  sample_and_hold_1
timestamp 1626065694
transform 1 0 253730 0 1 -149196
box -1766 -2168 42040 29538
use peak_detector  peak_detector_0
timestamp 1626065694
transform 1 0 173892 0 1 -185010
box -16568 -878 76950 30828
use diff_to_se_converter  diff_to_se_converter_0
timestamp 1626065694
transform -1 0 194530 0 1 -150652
box -13514 -708 35912 30998
use input_amplifier  input_amplifier_0
timestamp 1626065694
transform -1 0 248960 0 1 -106680
box -13477 -708 90192 28340
use biquad_gm_c_filter  biquad_gm_c_filter_0
timestamp 1626065694
transform 1 0 187212 0 1 -113396
box -1552 -6079 23682 5275
use low_freq_pll  low_freq_pll_0
timestamp 1626065694
transform 1 0 211340 0 1 -129086
box 7294 -22262 38743 17578
use bias_current_distribution  bias_current_distribution_0
timestamp 1626065694
transform 1 0 268974 0 1 -98308
box -440 -10900 12700 3000
use pulse_generator  pulse_generator_0
timestamp 1626065694
transform -1 0 339666 0 1 -185362
box -72 -526 4688 670
use dac_8bit  dac_8bit_0
timestamp 1626065694
transform 1 0 326281 0 1 -110050
box -29235 -75903 58525 12
use dac_8bit  dac_8bit_1
timestamp 1626065694
transform 1 0 326281 0 1 -59040
box -29235 -75903 58525 12
<< labels >>
flabel metal5 s 251350 -185504 251356 -185498 1 FreeSans 600 0 0 0 VSS
flabel metal4 s 252560 -154626 252626 -154538 1 FreeSans 600 0 0 0 VDD
flabel metal3 s 336386 -135042 336406 -135028 1 FreeSans 600 0 0 0 q7A
flabel metal3 s 336392 -135326 336404 -135314 1 FreeSans 600 0 0 0 q6A
flabel metal3 s 336398 -135642 336402 -135632 1 FreeSans 600 0 0 0 q5A
flabel metal3 s 336394 -135924 336410 -135904 1 FreeSans 600 0 0 0 q4A
flabel metal3 s 336392 -136230 336400 -136218 1 FreeSans 600 0 0 0 q3A
flabel metal3 s 336402 -136498 336418 -136486 1 FreeSans 600 0 0 0 q2A
flabel metal3 s 336410 -136792 336422 -136778 1 FreeSans 600 0 0 0 q1A
flabel metal3 s 336388 -137080 336412 -137056 1 FreeSans 600 0 0 0 q0A
flabel metal3 s 297672 -182972 297684 -182956 1 FreeSans 600 0 0 0 vlowB
flabel metal3 s 297928 -184958 297938 -184946 1 FreeSans 600 0 0 0 vrefB
flabel metal3 s 297592 -131956 297600 -131944 1 FreeSans 600 0 0 0 vlowA
flabel metal3 s 297816 -133942 297832 -133926 1 FreeSans 600 0 0 0 vrefA
flabel metal2 s 377876 -131602 377900 -131586 1 FreeSans 600 0 0 0 adc_clk
flabel metal3 s 336360 -186390 336394 -186356 1 FreeSans 600 0 0 0 q7B
flabel metal3 s 336352 -186674 336380 -186650 1 FreeSans 600 0 0 0 q6B
flabel metal3 s 336360 -187004 336384 -186976 1 FreeSans 600 0 0 0 q5B
flabel metal3 s 336346 -187278 336366 -187250 1 FreeSans 600 0 0 0 q4B
flabel metal3 s 336360 -187572 336380 -187544 1 FreeSans 600 0 0 0 q3B
flabel metal3 s 336360 -187860 336384 -187828 1 FreeSans 600 0 0 0 q2B
flabel metal3 s 336380 -188130 336404 -188102 1 FreeSans 600 0 0 0 q1B
flabel metal3 s 336376 -188428 336404 -188404 1 FreeSans 600 0 0 0 q0B
flabel metal2 s 340136 -184296 340154 -184284 1 FreeSans 600 0 0 0 adc_clk
flabel metal1 s 339852 -184050 339870 -184034 1 FreeSans 600 0 0 0 sample
flabel metal3 s 296034 -178004 296042 -178000 1 FreeSans 600 0 0 0 vpeak_sampled
flabel metal2 s 297150 -127600 297164 -127580 1 FreeSans 600 0 0 0 vcp_sampled
flabel metal3 s 252684 -184830 252706 -184802 1 FreeSans 600 0 0 0 vpeak
flabel metal3 s 252302 -151498 252314 -151468 1 FreeSans 600 0 0 0 vcp
flabel metal3 s 233848 -113906 233872 -113882 1 FreeSans 600 0 0 0 vcomp
flabel metal2 s 207498 -136864 207514 -136850 1 FreeSans 600 0 0 0 vocm_filt
flabel metal2 s 190664 -107802 190678 -107782 1 FreeSans 600 0 0 0 vampp
flabel metal2 s 210568 -116246 210592 -116228 1 FreeSans 600 0 0 0 vfiltp
flabel metal2 s 210828 -117166 210854 -117146 1 FreeSans 600 0 0 0 vfiltm
flabel metal3 s 186922 -111650 186936 -111624 1 FreeSans 600 0 0 0 vintm
flabel metal3 s 186656 -111776 186678 -111748 1 FreeSans 600 0 0 0 vintp
flabel metal2 s 197976 -102334 197986 -102326 1 FreeSans 600 0 0 0 gain_ctrl_0
flabel metal3 s 200836 -99526 200866 -99496 1 FreeSans 600 0 0 0 vocm
flabel metal2 s 204160 -152696 204176 -152670 1 FreeSans 600 0 0 0 vse
flabel metal2 s 276048 -108136 276068 -108126 1 FreeSans 600 0 0 0 vbiasn
flabel metal2 s 280014 -96358 280028 -96342 1 FreeSans 600 0 0 0 vbiasp
flabel metal3 s 336424 -111070 336442 -111054 1 FreeSans 600 0 0 0 adc_vcaparrayA
flabel metal3 s 336538 -162098 336560 -162076 1 FreeSans 600 0 0 0 adc_vcaparrayB
flabel metal2 s 384914 -101012 384932 -101002 1 FreeSans 600 0 0 0 adc_compA
flabel metal2 s 384800 -152028 384810 -152024 1 FreeSans 600 0 0 0 adc_compB
flabel metal2 s 196520 -107834 196534 -107828 1 FreeSans 600 0 0 0 vampm
flabel metal2 s 199398 -83588 199416 -83576 1 FreeSans 600 0 0 0 gain_ctrl_1
flabel metal2 s 334794 -185540 334800 -185524 1 FreeSans 600 0 0 0 peak_detector_rst
flabel metal2 s 256268 -91234 256286 -91216 1 FreeSans 600 0 0 0 rst_n
flabel metal3 s 257576 -100770 257584 -100760 1 FreeSans 600 0 0 0 vhpf
flabel metal3 s 257954 -105312 257972 -105298 1 FreeSans 600 0 0 0 vincm
<< end >>
