magic
tech sky130A
magscale 1 2
timestamp 1622610004
<< nwell >>
rect 74185 58508 76094 59026
rect 74185 58187 76419 58508
rect 74185 58186 76094 58187
<< pwell >>
rect 76043 58128 76073 58130
rect 76043 58092 76094 58128
rect 74185 57472 76094 58092
rect 76153 57947 76339 58129
rect 76318 57943 76339 57947
rect 76318 57909 76352 57943
<< nmos >>
rect 74381 57682 74581 57882
rect 74639 57682 74839 57882
rect 74897 57682 75097 57882
rect 75155 57682 75355 57882
rect 75413 57682 75613 57882
rect 75671 57682 75871 57882
<< scnmos >>
rect 76231 57973 76261 58103
<< scpmoshvt >>
rect 76231 58223 76261 58423
<< pmoshvt >>
rect 74381 58406 74581 58806
rect 74639 58406 74839 58806
rect 74897 58406 75097 58806
rect 75155 58406 75355 58806
rect 75413 58406 75613 58806
rect 75671 58406 75871 58806
<< ndiff >>
rect 76179 58091 76231 58103
rect 76179 58057 76187 58091
rect 76221 58057 76231 58091
rect 76179 58023 76231 58057
rect 76179 57989 76187 58023
rect 76221 57989 76231 58023
rect 76179 57973 76231 57989
rect 76261 58091 76313 58103
rect 76261 58057 76271 58091
rect 76305 58057 76313 58091
rect 76261 58023 76313 58057
rect 76261 57989 76271 58023
rect 76305 57989 76313 58023
rect 76261 57973 76313 57989
rect 74323 57870 74381 57882
rect 74323 57694 74335 57870
rect 74369 57694 74381 57870
rect 74323 57682 74381 57694
rect 74581 57870 74639 57882
rect 74581 57694 74593 57870
rect 74627 57694 74639 57870
rect 74581 57682 74639 57694
rect 74839 57870 74897 57882
rect 74839 57694 74851 57870
rect 74885 57694 74897 57870
rect 74839 57682 74897 57694
rect 75097 57870 75155 57882
rect 75097 57694 75109 57870
rect 75143 57694 75155 57870
rect 75097 57682 75155 57694
rect 75355 57870 75413 57882
rect 75355 57694 75367 57870
rect 75401 57694 75413 57870
rect 75355 57682 75413 57694
rect 75613 57870 75671 57882
rect 75613 57694 75625 57870
rect 75659 57694 75671 57870
rect 75613 57682 75671 57694
rect 75871 57870 75929 57882
rect 75871 57694 75883 57870
rect 75917 57694 75929 57870
rect 75871 57682 75929 57694
<< pdiff >>
rect 74323 58794 74381 58806
rect 74323 58418 74335 58794
rect 74369 58418 74381 58794
rect 74323 58406 74381 58418
rect 74581 58794 74639 58806
rect 74581 58418 74593 58794
rect 74627 58418 74639 58794
rect 74581 58406 74639 58418
rect 74839 58794 74897 58806
rect 74839 58418 74851 58794
rect 74885 58418 74897 58794
rect 74839 58406 74897 58418
rect 75097 58794 75155 58806
rect 75097 58418 75109 58794
rect 75143 58418 75155 58794
rect 75097 58406 75155 58418
rect 75355 58794 75413 58806
rect 75355 58418 75367 58794
rect 75401 58418 75413 58794
rect 75355 58406 75413 58418
rect 75613 58794 75671 58806
rect 75613 58418 75625 58794
rect 75659 58418 75671 58794
rect 75613 58406 75671 58418
rect 75871 58794 75929 58806
rect 75871 58418 75883 58794
rect 75917 58418 75929 58794
rect 75871 58406 75929 58418
rect 76179 58411 76231 58423
rect 76179 58377 76187 58411
rect 76221 58377 76231 58411
rect 76179 58343 76231 58377
rect 76179 58309 76187 58343
rect 76221 58309 76231 58343
rect 76179 58275 76231 58309
rect 76179 58241 76187 58275
rect 76221 58241 76231 58275
rect 76179 58223 76231 58241
rect 76261 58411 76313 58423
rect 76261 58377 76271 58411
rect 76305 58377 76313 58411
rect 76261 58343 76313 58377
rect 76261 58309 76271 58343
rect 76305 58309 76313 58343
rect 76261 58275 76313 58309
rect 76261 58241 76271 58275
rect 76305 58241 76313 58275
rect 76261 58223 76313 58241
<< ndiffc >>
rect 76187 58057 76221 58091
rect 76187 57989 76221 58023
rect 76271 58057 76305 58091
rect 76271 57989 76305 58023
rect 74335 57694 74369 57870
rect 74593 57694 74627 57870
rect 74851 57694 74885 57870
rect 75109 57694 75143 57870
rect 75367 57694 75401 57870
rect 75625 57694 75659 57870
rect 75883 57694 75917 57870
<< pdiffc >>
rect 74335 58418 74369 58794
rect 74593 58418 74627 58794
rect 74851 58418 74885 58794
rect 75109 58418 75143 58794
rect 75367 58418 75401 58794
rect 75625 58418 75659 58794
rect 75883 58418 75917 58794
rect 76187 58377 76221 58411
rect 76187 58309 76221 58343
rect 76187 58241 76221 58275
rect 76271 58377 76305 58411
rect 76271 58309 76305 58343
rect 76271 58241 76305 58275
<< psubdiff >>
rect 74221 58022 74317 58056
rect 75935 58022 76031 58056
rect 74221 57960 74255 58022
rect 75997 57960 76031 58022
rect 74221 57542 74255 57604
rect 75997 57542 76031 57604
rect 74221 57508 74317 57542
rect 75935 57508 76031 57542
<< nsubdiff >>
rect 74221 58955 74317 58989
rect 75935 58955 76031 58989
rect 74221 58893 74255 58955
rect 75997 58893 76031 58955
rect 74221 58257 74255 58319
rect 75997 58257 76031 58319
rect 74221 58223 74317 58257
rect 75935 58223 76031 58257
<< psubdiffcont >>
rect 74317 58022 75935 58056
rect 74221 57604 74255 57960
rect 75997 57604 76031 57960
rect 74317 57508 75935 57542
<< nsubdiffcont >>
rect 74317 58955 75935 58989
rect 74221 58319 74255 58893
rect 75997 58319 76031 58893
rect 74317 58223 75935 58257
<< poly >>
rect 74415 58887 74547 58903
rect 74415 58870 74431 58887
rect 74381 58853 74431 58870
rect 74531 58870 74547 58887
rect 74673 58887 74805 58903
rect 74673 58870 74689 58887
rect 74531 58853 74581 58870
rect 74381 58806 74581 58853
rect 74639 58853 74689 58870
rect 74789 58870 74805 58887
rect 74931 58887 75063 58903
rect 74931 58870 74947 58887
rect 74789 58853 74839 58870
rect 74639 58806 74839 58853
rect 74897 58853 74947 58870
rect 75047 58870 75063 58887
rect 75189 58887 75321 58903
rect 75189 58870 75205 58887
rect 75047 58853 75097 58870
rect 74897 58806 75097 58853
rect 75155 58853 75205 58870
rect 75305 58870 75321 58887
rect 75447 58887 75579 58903
rect 75447 58870 75463 58887
rect 75305 58853 75355 58870
rect 75155 58806 75355 58853
rect 75413 58853 75463 58870
rect 75563 58870 75579 58887
rect 75705 58887 75837 58903
rect 75705 58870 75721 58887
rect 75563 58853 75613 58870
rect 75413 58806 75613 58853
rect 75671 58853 75721 58870
rect 75821 58870 75837 58887
rect 75821 58853 75871 58870
rect 75671 58806 75871 58853
rect 74381 58359 74581 58406
rect 74381 58342 74431 58359
rect 74415 58325 74431 58342
rect 74531 58342 74581 58359
rect 74639 58359 74839 58406
rect 74639 58342 74689 58359
rect 74531 58325 74547 58342
rect 74415 58309 74547 58325
rect 74673 58325 74689 58342
rect 74789 58342 74839 58359
rect 74897 58359 75097 58406
rect 74897 58342 74947 58359
rect 74789 58325 74805 58342
rect 74673 58309 74805 58325
rect 74931 58325 74947 58342
rect 75047 58342 75097 58359
rect 75155 58359 75355 58406
rect 75155 58342 75205 58359
rect 75047 58325 75063 58342
rect 74931 58309 75063 58325
rect 75189 58325 75205 58342
rect 75305 58342 75355 58359
rect 75413 58359 75613 58406
rect 75413 58342 75463 58359
rect 75305 58325 75321 58342
rect 75189 58309 75321 58325
rect 75447 58325 75463 58342
rect 75563 58342 75613 58359
rect 75671 58359 75871 58406
rect 75671 58342 75721 58359
rect 75563 58325 75579 58342
rect 75447 58309 75579 58325
rect 75705 58325 75721 58342
rect 75821 58342 75871 58359
rect 75821 58325 75837 58342
rect 75705 58309 75837 58325
rect 76231 58423 76261 58449
rect 76231 58191 76261 58223
rect 76231 58175 76317 58191
rect 76231 58141 76267 58175
rect 76301 58141 76317 58175
rect 76231 58125 76317 58141
rect 76231 58103 76261 58125
rect 74415 57954 74547 57970
rect 74415 57937 74431 57954
rect 74381 57920 74431 57937
rect 74531 57937 74547 57954
rect 74673 57954 74805 57970
rect 74673 57937 74689 57954
rect 74531 57920 74581 57937
rect 74381 57882 74581 57920
rect 74639 57920 74689 57937
rect 74789 57937 74805 57954
rect 74931 57954 75063 57970
rect 74931 57937 74947 57954
rect 74789 57920 74839 57937
rect 74639 57882 74839 57920
rect 74897 57920 74947 57937
rect 75047 57937 75063 57954
rect 75189 57954 75321 57970
rect 75189 57937 75205 57954
rect 75047 57920 75097 57937
rect 74897 57882 75097 57920
rect 75155 57920 75205 57937
rect 75305 57937 75321 57954
rect 75447 57954 75579 57970
rect 75447 57937 75463 57954
rect 75305 57920 75355 57937
rect 75155 57882 75355 57920
rect 75413 57920 75463 57937
rect 75563 57937 75579 57954
rect 75705 57954 75837 57970
rect 75705 57937 75721 57954
rect 75563 57920 75613 57937
rect 75413 57882 75613 57920
rect 75671 57920 75721 57937
rect 75821 57937 75837 57954
rect 75821 57920 75871 57937
rect 75671 57882 75871 57920
rect 74381 57644 74581 57682
rect 74381 57627 74431 57644
rect 74415 57610 74431 57627
rect 74531 57627 74581 57644
rect 74639 57644 74839 57682
rect 74639 57627 74689 57644
rect 74531 57610 74547 57627
rect 74415 57594 74547 57610
rect 74673 57610 74689 57627
rect 74789 57627 74839 57644
rect 74897 57644 75097 57682
rect 74897 57627 74947 57644
rect 74789 57610 74805 57627
rect 74673 57594 74805 57610
rect 74931 57610 74947 57627
rect 75047 57627 75097 57644
rect 75155 57644 75355 57682
rect 75155 57627 75205 57644
rect 75047 57610 75063 57627
rect 74931 57594 75063 57610
rect 75189 57610 75205 57627
rect 75305 57627 75355 57644
rect 75413 57644 75613 57682
rect 75413 57627 75463 57644
rect 75305 57610 75321 57627
rect 75189 57594 75321 57610
rect 75447 57610 75463 57627
rect 75563 57627 75613 57644
rect 75671 57644 75871 57682
rect 75671 57627 75721 57644
rect 75563 57610 75579 57627
rect 75447 57594 75579 57610
rect 75705 57610 75721 57627
rect 75821 57627 75871 57644
rect 75821 57610 75837 57627
rect 75705 57594 75837 57610
rect 76231 57947 76261 57973
<< polycont >>
rect 74431 58853 74531 58887
rect 74689 58853 74789 58887
rect 74947 58853 75047 58887
rect 75205 58853 75305 58887
rect 75463 58853 75563 58887
rect 75721 58853 75821 58887
rect 74431 58325 74531 58359
rect 74689 58325 74789 58359
rect 74947 58325 75047 58359
rect 75205 58325 75305 58359
rect 75463 58325 75563 58359
rect 75721 58325 75821 58359
rect 76267 58141 76301 58175
rect 74431 57920 74531 57954
rect 74689 57920 74789 57954
rect 74947 57920 75047 57954
rect 75205 57920 75305 57954
rect 75463 57920 75563 57954
rect 75721 57920 75821 57954
rect 74431 57610 74531 57644
rect 74689 57610 74789 57644
rect 74947 57610 75047 57644
rect 75205 57610 75305 57644
rect 75463 57610 75563 57644
rect 75721 57610 75821 57644
<< locali >>
rect 74221 58956 74267 58989
rect 75961 58956 76031 58989
rect 74221 58955 74317 58956
rect 75935 58955 76031 58956
rect 74221 58893 74255 58955
rect 75997 58894 76031 58955
rect 74415 58853 74431 58887
rect 74531 58853 74547 58887
rect 74673 58853 74689 58887
rect 74789 58853 74805 58887
rect 74931 58853 74947 58887
rect 75047 58853 75063 58887
rect 75189 58853 75205 58887
rect 75305 58853 75321 58887
rect 75447 58853 75463 58887
rect 75563 58853 75579 58887
rect 75705 58853 75721 58887
rect 75821 58853 75837 58887
rect 74335 58794 74369 58810
rect 74335 58402 74369 58418
rect 74593 58794 74627 58810
rect 74593 58402 74627 58418
rect 74851 58794 74885 58810
rect 74851 58402 74885 58418
rect 75109 58794 75143 58810
rect 75109 58402 75143 58418
rect 75367 58794 75401 58810
rect 75367 58402 75401 58418
rect 75625 58794 75659 58810
rect 75625 58402 75659 58418
rect 75883 58794 75917 58810
rect 75883 58402 75917 58418
rect 74415 58325 74431 58359
rect 74531 58325 74547 58359
rect 74673 58325 74689 58359
rect 74789 58325 74805 58359
rect 74931 58325 74947 58359
rect 75047 58325 75063 58359
rect 75189 58325 75205 58359
rect 75305 58325 75321 58359
rect 75447 58325 75463 58359
rect 75563 58325 75579 58359
rect 75705 58325 75721 58359
rect 75821 58325 75837 58359
rect 74221 58257 74255 58319
rect 76105 58453 76134 58487
rect 76168 58453 76226 58487
rect 76260 58453 76318 58487
rect 76352 58453 76381 58487
rect 75997 58257 76031 58318
rect 74221 58256 74317 58257
rect 74221 58223 74267 58256
rect 75961 58224 76031 58257
rect 75935 58223 76031 58224
rect 76171 58411 76237 58419
rect 76171 58377 76187 58411
rect 76221 58377 76237 58411
rect 76171 58343 76237 58377
rect 76171 58309 76187 58343
rect 76221 58309 76237 58343
rect 76171 58275 76237 58309
rect 76171 58241 76187 58275
rect 76221 58241 76237 58275
rect 76171 58223 76237 58241
rect 76271 58411 76313 58453
rect 76305 58377 76313 58411
rect 76271 58343 76313 58377
rect 76305 58309 76313 58343
rect 76271 58275 76313 58309
rect 76305 58241 76313 58275
rect 76271 58225 76313 58241
rect 76171 58164 76217 58223
rect 76212 58116 76217 58164
rect 76251 58186 76317 58189
rect 76251 58175 76268 58186
rect 76251 58141 76267 58175
rect 76314 58146 76317 58186
rect 76301 58141 76317 58146
rect 76171 58103 76217 58116
rect 76171 58091 76237 58103
rect 76171 58057 76187 58091
rect 76221 58057 76237 58091
rect 74221 58022 74291 58056
rect 75961 58022 76031 58056
rect 74221 57960 74255 58022
rect 75997 57960 76031 58022
rect 76171 58023 76237 58057
rect 76171 57989 76187 58023
rect 76221 57989 76237 58023
rect 76171 57977 76237 57989
rect 76271 58091 76317 58107
rect 76305 58057 76317 58091
rect 76271 58023 76317 58057
rect 76305 57989 76317 58023
rect 74415 57920 74431 57954
rect 74531 57920 74547 57954
rect 74673 57920 74689 57954
rect 74789 57920 74805 57954
rect 74931 57920 74947 57954
rect 75047 57920 75063 57954
rect 75189 57920 75205 57954
rect 75305 57920 75321 57954
rect 75447 57920 75463 57954
rect 75563 57920 75579 57954
rect 75705 57920 75721 57954
rect 75821 57920 75837 57954
rect 74335 57870 74369 57886
rect 74335 57678 74369 57694
rect 74593 57870 74627 57886
rect 74593 57678 74627 57694
rect 74851 57870 74885 57886
rect 74851 57678 74885 57694
rect 75109 57870 75143 57886
rect 75109 57678 75143 57694
rect 75367 57870 75401 57886
rect 75367 57678 75401 57694
rect 75625 57870 75659 57886
rect 75625 57678 75659 57694
rect 75883 57870 75917 57886
rect 75883 57678 75917 57694
rect 74415 57610 74431 57644
rect 74531 57610 74547 57644
rect 74673 57610 74689 57644
rect 74789 57610 74805 57644
rect 74931 57610 74947 57644
rect 75047 57610 75063 57644
rect 75189 57610 75205 57644
rect 75305 57610 75321 57644
rect 75447 57610 75463 57644
rect 75563 57610 75579 57644
rect 75705 57610 75721 57644
rect 75821 57610 75837 57644
rect 76271 57943 76317 57989
rect 76105 57909 76134 57943
rect 76168 57909 76226 57943
rect 76260 57909 76318 57943
rect 76352 57909 76381 57943
rect 74221 57542 74255 57604
rect 75997 57542 76031 57604
rect 74221 57508 74289 57542
rect 75963 57508 76031 57542
<< viali >>
rect 74267 58989 74487 58990
rect 75759 58989 75961 58990
rect 74267 58956 74317 58989
rect 74317 58956 74487 58989
rect 75759 58956 75935 58989
rect 75935 58956 75961 58989
rect 75995 58893 76031 58894
rect 74219 58320 74221 58892
rect 74221 58320 74255 58892
rect 74255 58320 74257 58892
rect 74439 58853 74523 58887
rect 74697 58853 74781 58887
rect 74955 58853 75039 58887
rect 75213 58853 75297 58887
rect 75471 58853 75555 58887
rect 75729 58853 75813 58887
rect 74335 58418 74369 58794
rect 74593 58418 74627 58794
rect 74851 58418 74885 58794
rect 75109 58418 75143 58794
rect 75367 58418 75401 58794
rect 75625 58418 75659 58794
rect 75883 58418 75917 58794
rect 74439 58325 74523 58359
rect 74697 58325 74781 58359
rect 74955 58325 75039 58359
rect 75213 58325 75297 58359
rect 75471 58325 75555 58359
rect 75729 58325 75813 58359
rect 75995 58319 75997 58893
rect 75997 58319 76031 58893
rect 76134 58453 76168 58487
rect 76226 58453 76260 58487
rect 76318 58453 76352 58487
rect 75995 58318 76031 58319
rect 75759 58257 75961 58258
rect 74267 58223 74317 58256
rect 74317 58223 74487 58256
rect 75759 58224 75935 58257
rect 75935 58224 75961 58257
rect 74267 58222 74487 58223
rect 76164 58116 76212 58164
rect 76268 58175 76314 58186
rect 76268 58146 76301 58175
rect 76301 58146 76314 58175
rect 74291 58056 74499 58058
rect 75763 58056 75961 58060
rect 74291 58022 74317 58056
rect 74317 58022 74499 58056
rect 75763 58022 75935 58056
rect 75935 58022 75961 58056
rect 74291 58020 74499 58022
rect 74219 57604 74221 57960
rect 74221 57604 74255 57960
rect 74439 57920 74523 57954
rect 74697 57920 74781 57954
rect 74955 57920 75039 57954
rect 75213 57920 75297 57954
rect 75471 57920 75555 57954
rect 75729 57920 75813 57954
rect 74335 57694 74369 57870
rect 74593 57694 74627 57870
rect 74851 57694 74885 57870
rect 75109 57694 75143 57870
rect 75367 57694 75401 57870
rect 75625 57694 75659 57870
rect 75883 57694 75917 57870
rect 74439 57610 74523 57644
rect 74697 57610 74781 57644
rect 74955 57610 75039 57644
rect 75213 57610 75297 57644
rect 75471 57610 75555 57644
rect 75729 57610 75813 57644
rect 75995 57604 75997 57960
rect 75997 57604 76031 57960
rect 76031 57604 76033 57960
rect 76134 57909 76168 57943
rect 76226 57909 76260 57943
rect 76318 57909 76352 57943
rect 74289 57542 74497 57544
rect 74289 57508 74317 57542
rect 74317 57508 74497 57542
rect 75761 57508 75935 57542
rect 75935 57508 75963 57542
rect 75761 57506 75963 57508
<< metal1 >>
rect 74208 59056 76044 59116
rect 74208 59004 74268 59056
rect 74319 59004 74379 59056
rect 74208 59002 74379 59004
rect 74453 59002 74513 59056
rect 74208 58990 74513 59002
rect 74208 58956 74267 58990
rect 74487 58956 74513 58990
rect 74208 58942 74513 58956
rect 74208 58892 74269 58942
rect 74208 58862 74219 58892
rect 74209 58634 74219 58862
rect 74208 58574 74219 58634
rect 74209 58320 74219 58574
rect 74257 58634 74269 58892
rect 74319 58794 74379 58942
rect 74453 58893 74513 58942
rect 74709 59008 74769 59009
rect 75485 59008 75545 59014
rect 74709 58948 75485 59008
rect 74709 58893 74769 58948
rect 74967 58893 75027 58948
rect 75225 58893 75285 58948
rect 75485 58893 75545 58948
rect 75741 59006 75801 59056
rect 75869 59006 75929 59056
rect 75984 59006 76044 59056
rect 75741 58990 76044 59006
rect 75741 58956 75759 58990
rect 75961 58956 76044 58990
rect 75741 58942 76044 58956
rect 75741 58893 75801 58942
rect 74427 58887 74535 58893
rect 74427 58853 74439 58887
rect 74523 58853 74535 58887
rect 74427 58847 74535 58853
rect 74685 58887 74793 58893
rect 74685 58853 74697 58887
rect 74781 58853 74793 58887
rect 74685 58847 74793 58853
rect 74943 58887 75051 58893
rect 74943 58853 74955 58887
rect 75039 58853 75051 58887
rect 74943 58847 75051 58853
rect 75201 58887 75309 58893
rect 75201 58853 75213 58887
rect 75297 58853 75309 58887
rect 75201 58847 75309 58853
rect 75459 58887 75567 58893
rect 75459 58853 75471 58887
rect 75555 58853 75567 58887
rect 75459 58847 75567 58853
rect 75717 58887 75825 58893
rect 75717 58853 75729 58887
rect 75813 58853 75825 58887
rect 75717 58847 75825 58853
rect 74319 58634 74335 58794
rect 74257 58574 74335 58634
rect 74257 58320 74269 58574
rect 74329 58452 74335 58574
rect 74209 58270 74269 58320
rect 74321 58418 74335 58452
rect 74369 58574 74379 58794
rect 74587 58794 74633 58806
rect 74369 58452 74375 58574
rect 74587 58463 74593 58794
rect 74369 58418 74381 58452
rect 74321 58270 74381 58418
rect 74579 58418 74593 58463
rect 74627 58463 74633 58794
rect 74845 58794 74891 58806
rect 74627 58418 74639 58463
rect 74845 58438 74851 58794
rect 74427 58359 74535 58365
rect 74427 58325 74439 58359
rect 74523 58325 74535 58359
rect 74427 58319 74535 58325
rect 74449 58270 74509 58319
rect 74208 58256 74509 58270
rect 74208 58222 74267 58256
rect 74487 58222 74509 58256
rect 74208 58210 74509 58222
rect 74579 58093 74639 58418
rect 74837 58418 74851 58438
rect 74885 58438 74891 58794
rect 75103 58794 75149 58806
rect 75103 58461 75109 58794
rect 74885 58418 74897 58438
rect 74685 58359 74793 58365
rect 74685 58325 74697 58359
rect 74781 58325 74793 58359
rect 74685 58319 74793 58325
rect 74837 58242 74897 58418
rect 75095 58418 75109 58461
rect 75143 58461 75149 58794
rect 75361 58794 75407 58806
rect 75143 58418 75155 58461
rect 75361 58456 75367 58794
rect 74943 58359 75051 58365
rect 74943 58325 74955 58359
rect 75039 58325 75051 58359
rect 74943 58319 75051 58325
rect 74831 58182 74837 58242
rect 74897 58182 74903 58242
rect 74207 58058 74511 58068
rect 74207 58020 74291 58058
rect 74499 58020 74511 58058
rect 74573 58033 74579 58093
rect 74639 58033 74645 58093
rect 74207 58008 74511 58020
rect 74207 57960 74267 58008
rect 74207 57604 74219 57960
rect 74255 57604 74267 57960
rect 74321 57870 74381 58008
rect 74451 57960 74511 58008
rect 74427 57954 74535 57960
rect 74427 57920 74439 57954
rect 74523 57920 74535 57954
rect 74427 57914 74535 57920
rect 74321 57820 74335 57870
rect 74329 57733 74335 57820
rect 74207 57555 74267 57604
rect 74323 57694 74335 57733
rect 74369 57820 74381 57870
rect 74579 57870 74639 58033
rect 74685 57954 74793 57960
rect 74685 57920 74697 57954
rect 74781 57920 74793 57954
rect 74685 57914 74793 57920
rect 74579 57833 74593 57870
rect 74369 57733 74375 57820
rect 74369 57694 74383 57733
rect 74323 57555 74383 57694
rect 74587 57694 74593 57833
rect 74627 57833 74639 57870
rect 74837 57900 74897 58182
rect 75095 58093 75155 58418
rect 75355 58418 75367 58456
rect 75401 58456 75407 58794
rect 75619 58794 75665 58806
rect 75619 58461 75625 58794
rect 75401 58418 75415 58456
rect 75201 58359 75309 58365
rect 75201 58325 75213 58359
rect 75297 58325 75309 58359
rect 75201 58319 75309 58325
rect 75355 58242 75415 58418
rect 75613 58418 75625 58461
rect 75659 58461 75665 58794
rect 75869 58794 75929 58942
rect 75869 58576 75883 58794
rect 75659 58418 75673 58461
rect 75877 58448 75883 58576
rect 75459 58359 75567 58365
rect 75459 58325 75471 58359
rect 75555 58325 75567 58359
rect 75459 58319 75567 58325
rect 75349 58182 75355 58242
rect 75415 58182 75421 58242
rect 75089 58033 75095 58093
rect 75155 58033 75161 58093
rect 74943 57954 75051 57960
rect 74943 57920 74955 57954
rect 75039 57920 75051 57954
rect 74943 57914 75051 57920
rect 74837 57870 74899 57900
rect 74837 57834 74851 57870
rect 74627 57694 74633 57833
rect 74587 57682 74633 57694
rect 74839 57694 74851 57834
rect 74885 57694 74899 57870
rect 75095 57870 75155 58033
rect 75201 57954 75309 57960
rect 75201 57920 75213 57954
rect 75297 57920 75309 57954
rect 75201 57914 75309 57920
rect 75095 57714 75109 57870
rect 74839 57654 74899 57694
rect 75103 57694 75109 57714
rect 75143 57714 75155 57870
rect 75355 57870 75415 58182
rect 75613 58093 75673 58418
rect 75871 58418 75883 58448
rect 75917 58636 75929 58794
rect 75983 58894 76044 58942
rect 75983 58636 75995 58894
rect 75917 58576 75995 58636
rect 75917 58448 75923 58576
rect 75917 58418 75931 58448
rect 75717 58359 75825 58365
rect 75717 58325 75729 58359
rect 75813 58325 75825 58359
rect 75717 58319 75825 58325
rect 75737 58270 75797 58319
rect 75871 58270 75931 58418
rect 75983 58318 75995 58576
rect 76031 58878 76044 58894
rect 76031 58518 76043 58878
rect 76031 58487 76381 58518
rect 76031 58453 76134 58487
rect 76168 58453 76226 58487
rect 76260 58453 76318 58487
rect 76352 58453 76381 58487
rect 76031 58422 76381 58453
rect 76031 58318 76043 58422
rect 75983 58270 76043 58318
rect 75737 58258 76043 58270
rect 75737 58224 75759 58258
rect 75961 58224 76043 58258
rect 75737 58210 76043 58224
rect 76476 58192 76536 58198
rect 76256 58186 76476 58192
rect 76158 58170 76218 58176
rect 76152 58110 76158 58170
rect 76218 58110 76224 58170
rect 76256 58146 76268 58186
rect 76314 58146 76476 58186
rect 76256 58132 76476 58146
rect 76476 58126 76536 58132
rect 76158 58104 76218 58110
rect 75459 57954 75567 57960
rect 75459 57920 75471 57954
rect 75555 57920 75567 57954
rect 75459 57914 75567 57920
rect 75143 57694 75149 57714
rect 75103 57682 75149 57694
rect 75355 57694 75367 57870
rect 75401 57694 75415 57870
rect 75613 57870 75673 58033
rect 75743 58060 76045 58070
rect 75743 58022 75763 58060
rect 75961 58022 76045 58060
rect 75743 58010 76045 58022
rect 75743 57960 75803 58010
rect 75717 57954 75825 57960
rect 75717 57920 75729 57954
rect 75813 57920 75825 57954
rect 75717 57914 75825 57920
rect 75613 57831 75625 57870
rect 75355 57654 75415 57694
rect 75619 57694 75625 57831
rect 75659 57831 75673 57870
rect 75871 57870 75931 58010
rect 75659 57694 75665 57831
rect 75871 57824 75883 57870
rect 75877 57727 75883 57824
rect 75619 57682 75665 57694
rect 75869 57694 75883 57727
rect 75917 57824 75931 57870
rect 75985 57974 76045 58010
rect 75985 57960 76381 57974
rect 75917 57727 75923 57824
rect 75917 57694 75929 57727
rect 74427 57644 74535 57650
rect 74427 57610 74439 57644
rect 74523 57610 74535 57644
rect 74427 57604 74535 57610
rect 74685 57644 74793 57650
rect 74685 57610 74697 57644
rect 74781 57610 74793 57644
rect 74685 57604 74793 57610
rect 74943 57644 75051 57650
rect 74943 57610 74955 57644
rect 75039 57610 75051 57644
rect 74943 57604 75051 57610
rect 75201 57644 75309 57650
rect 75201 57610 75213 57644
rect 75297 57610 75309 57644
rect 75201 57604 75309 57610
rect 75459 57644 75567 57650
rect 75459 57610 75471 57644
rect 75555 57610 75567 57644
rect 75459 57604 75567 57610
rect 75717 57644 75825 57650
rect 75717 57610 75729 57644
rect 75813 57610 75825 57644
rect 75717 57604 75825 57610
rect 74451 57555 74511 57604
rect 74207 57544 74511 57555
rect 74207 57508 74289 57544
rect 74497 57508 74511 57544
rect 74207 57495 74511 57508
rect 74207 57438 74267 57495
rect 74208 57420 74267 57438
rect 74323 57420 74383 57495
rect 74451 57420 74511 57495
rect 74709 57545 74769 57604
rect 74969 57545 75029 57604
rect 75227 57545 75287 57604
rect 75483 57545 75543 57604
rect 75741 57555 75801 57604
rect 75869 57555 75929 57694
rect 75985 57604 75995 57960
rect 76033 57943 76381 57960
rect 76033 57909 76134 57943
rect 76168 57909 76226 57943
rect 76260 57909 76318 57943
rect 76352 57909 76381 57943
rect 76033 57878 76381 57909
rect 76033 57604 76045 57878
rect 75985 57555 76045 57604
rect 74709 57485 75483 57545
rect 75543 57485 75549 57545
rect 75741 57542 76045 57555
rect 75741 57506 75761 57542
rect 75963 57506 76045 57542
rect 75741 57495 76045 57506
rect 75741 57420 75801 57495
rect 75869 57420 75929 57495
rect 75985 57420 76045 57495
rect 74208 57360 76046 57420
<< via1 >>
rect 75485 58948 75545 59008
rect 74837 58182 74897 58242
rect 74579 58033 74639 58093
rect 75355 58182 75415 58242
rect 75095 58033 75155 58093
rect 76158 58164 76218 58170
rect 76158 58116 76164 58164
rect 76164 58116 76212 58164
rect 76212 58116 76218 58164
rect 76158 58110 76218 58116
rect 76476 58132 76536 58192
rect 75613 58033 75673 58093
rect 75483 57485 75543 57545
<< metal2 >>
rect 75479 58948 75485 59008
rect 75545 58948 76144 59008
rect 74837 58242 74897 58248
rect 75355 58242 75415 58248
rect 74897 58182 75355 58242
rect 74837 58176 74897 58182
rect 75355 58176 75415 58182
rect 76084 58170 76144 58948
rect 76084 58110 76158 58170
rect 76218 58110 76224 58170
rect 76470 58132 76476 58192
rect 76536 58132 76542 58192
rect 74579 58093 74639 58099
rect 75095 58093 75155 58099
rect 74568 58033 74579 58093
rect 74639 58033 75095 58093
rect 75155 58033 75613 58093
rect 75673 58033 75679 58093
rect 74579 58027 74639 58033
rect 75095 58027 75155 58033
rect 75483 57545 75543 57551
rect 76476 57546 76536 58132
rect 75990 57545 76536 57546
rect 75543 57486 76536 57545
rect 75543 57485 76094 57486
rect 75483 57479 75543 57485
<< labels >>
flabel metal1 76416 58154 76424 58160 1 FreeSans 480 0 0 0 tx
port 5 n
flabel metal1 74598 58134 74608 58142 1 FreeSans 480 0 0 0 out
port 2 n
flabel metal1 74860 58140 74870 58148 1 FreeSans 480 0 0 0 in
port 1 n
flabel metal1 75114 59082 75124 59092 1 FreeSans 480 0 0 0 VDD
port 3 n power bidirectional
flabel metal1 75112 57392 75120 57398 1 FreeSans 480 0 0 0 VSS
port 4 n ground bidirectional
flabel metal2 76114 58656 76124 58664 1 FreeSans 480 0 0 0 txb
flabel locali 76183 58215 76217 58249 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 76183 58147 76217 58181 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 76275 58147 76309 58181 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 76318 58453 76352 58487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 76318 57909 76352 57943 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 76318 57909 76352 57943 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 76318 58453 76352 58487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 76381 57926 76381 57926 6 sky130_fd_sc_hd__inv_1_0/inv_1
<< end >>
