magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< poly >>
rect 1671 402 1701 896
rect 2295 526 2325 896
rect 2919 650 2949 896
rect 3543 774 3573 896
rect 4167 402 4197 896
rect 4791 526 4821 896
rect 5415 650 5445 896
rect 6039 774 6069 896
rect 6663 402 6693 896
rect 7287 526 7317 896
rect 7911 650 7941 896
rect 8535 774 8565 896
rect 9159 402 9189 896
rect 9783 526 9813 896
rect 10407 650 10437 896
rect 11031 774 11061 896
rect 11655 402 11685 896
rect 12279 526 12309 896
rect 12903 650 12933 896
rect 13527 774 13557 896
rect 14151 402 14181 896
rect 14775 526 14805 896
rect 15399 650 15429 896
rect 16023 774 16053 896
rect 16647 402 16677 896
rect 17271 526 17301 896
rect 17895 650 17925 896
rect 18519 774 18549 896
rect 19143 402 19173 896
rect 19767 526 19797 896
rect 20391 650 20421 896
rect 21015 774 21045 896
rect 21639 402 21669 896
rect 22263 526 22293 896
rect 22887 650 22917 896
rect 23511 774 23541 896
rect 24135 402 24165 896
rect 24759 526 24789 896
rect 25383 650 25413 896
rect 26007 774 26037 896
rect 26631 402 26661 896
rect 27255 526 27285 896
rect 27879 650 27909 896
rect 28503 774 28533 896
rect 29127 402 29157 896
rect 29751 526 29781 896
rect 30375 650 30405 896
rect 30999 774 31029 896
rect 31623 402 31653 896
rect 32247 526 32277 896
rect 32871 650 32901 896
rect 33495 774 33525 896
rect 34119 402 34149 896
rect 34743 526 34773 896
rect 35367 650 35397 896
rect 35991 774 36021 896
rect 36615 402 36645 896
rect 37239 526 37269 896
rect 37863 650 37893 896
rect 38487 774 38517 896
rect 39111 402 39141 896
rect 39735 526 39765 896
rect 40359 650 40389 896
rect 40983 774 41013 896
rect 41607 402 41637 896
rect 42231 526 42261 896
rect 42855 650 42885 896
rect 43479 774 43509 896
rect 44103 402 44133 896
rect 44727 526 44757 896
rect 45351 650 45381 896
rect 45975 774 46005 896
rect 46599 402 46629 896
rect 47223 526 47253 896
rect 47847 650 47877 896
rect 48471 774 48501 896
rect 49095 402 49125 896
rect 49719 526 49749 896
rect 50343 650 50373 896
rect 50967 774 50997 896
rect 51591 402 51621 896
rect 52215 526 52245 896
rect 52839 650 52869 896
rect 53463 774 53493 896
rect 54087 402 54117 896
rect 54711 526 54741 896
rect 55335 650 55365 896
rect 55959 774 55989 896
rect 56583 402 56613 896
rect 57207 526 57237 896
rect 57831 650 57861 896
rect 58455 774 58485 896
rect 59079 402 59109 896
rect 59703 526 59733 896
rect 60327 650 60357 896
rect 60951 774 60981 896
rect 61575 402 61605 896
rect 62199 526 62229 896
rect 62823 650 62853 896
rect 63447 774 63477 896
rect 64071 402 64101 896
rect 64695 526 64725 896
rect 65319 650 65349 896
rect 65943 774 65973 896
rect 66567 402 66597 896
rect 67191 526 67221 896
rect 67815 650 67845 896
rect 68439 774 68469 896
rect 69063 402 69093 896
rect 69687 526 69717 896
rect 70311 650 70341 896
rect 70935 774 70965 896
rect 71559 402 71589 896
rect 72183 526 72213 896
rect 72807 650 72837 896
rect 73431 774 73461 896
rect 74055 402 74085 896
rect 74679 526 74709 896
rect 75303 650 75333 896
rect 75927 774 75957 896
rect 76551 402 76581 896
rect 77175 526 77205 896
rect 77799 650 77829 896
rect 78423 774 78453 896
rect 79047 402 79077 896
rect 79671 526 79701 896
rect 80295 650 80325 896
rect 80919 774 80949 896
<< metal1 >>
rect 1454 2128 1482 2184
rect 1918 2128 1946 2184
rect 2050 2128 2078 2184
rect 2514 2128 2542 2184
rect 2702 2128 2730 2184
rect 3166 2128 3194 2184
rect 3298 2128 3326 2184
rect 3762 2128 3790 2184
rect 3950 2128 3978 2184
rect 4414 2128 4442 2184
rect 4546 2128 4574 2184
rect 5010 2128 5038 2184
rect 5198 2128 5226 2184
rect 5662 2128 5690 2184
rect 5794 2128 5822 2184
rect 6258 2128 6286 2184
rect 6446 2128 6474 2184
rect 6910 2128 6938 2184
rect 7042 2128 7070 2184
rect 7506 2128 7534 2184
rect 7694 2128 7722 2184
rect 8158 2128 8186 2184
rect 8290 2128 8318 2184
rect 8754 2128 8782 2184
rect 8942 2128 8970 2184
rect 9406 2128 9434 2184
rect 9538 2128 9566 2184
rect 10002 2128 10030 2184
rect 10190 2128 10218 2184
rect 10654 2128 10682 2184
rect 10786 2128 10814 2184
rect 11250 2128 11278 2184
rect 11438 2128 11466 2184
rect 11902 2128 11930 2184
rect 12034 2128 12062 2184
rect 12498 2128 12526 2184
rect 12686 2128 12714 2184
rect 13150 2128 13178 2184
rect 13282 2128 13310 2184
rect 13746 2128 13774 2184
rect 13934 2128 13962 2184
rect 14398 2128 14426 2184
rect 14530 2128 14558 2184
rect 14994 2128 15022 2184
rect 15182 2128 15210 2184
rect 15646 2128 15674 2184
rect 15778 2128 15806 2184
rect 16242 2128 16270 2184
rect 16430 2128 16458 2184
rect 16894 2128 16922 2184
rect 17026 2128 17054 2184
rect 17490 2128 17518 2184
rect 17678 2128 17706 2184
rect 18142 2128 18170 2184
rect 18274 2128 18302 2184
rect 18738 2128 18766 2184
rect 18926 2128 18954 2184
rect 19390 2128 19418 2184
rect 19522 2128 19550 2184
rect 19986 2128 20014 2184
rect 20174 2128 20202 2184
rect 20638 2128 20666 2184
rect 20770 2128 20798 2184
rect 21234 2128 21262 2184
rect 21422 2128 21450 2184
rect 21886 2128 21914 2184
rect 22018 2128 22046 2184
rect 22482 2128 22510 2184
rect 22670 2128 22698 2184
rect 23134 2128 23162 2184
rect 23266 2128 23294 2184
rect 23730 2128 23758 2184
rect 23918 2128 23946 2184
rect 24382 2128 24410 2184
rect 24514 2128 24542 2184
rect 24978 2128 25006 2184
rect 25166 2128 25194 2184
rect 25630 2128 25658 2184
rect 25762 2128 25790 2184
rect 26226 2128 26254 2184
rect 26414 2128 26442 2184
rect 26878 2128 26906 2184
rect 27010 2128 27038 2184
rect 27474 2128 27502 2184
rect 27662 2128 27690 2184
rect 28126 2128 28154 2184
rect 28258 2128 28286 2184
rect 28722 2128 28750 2184
rect 28910 2128 28938 2184
rect 29374 2128 29402 2184
rect 29506 2128 29534 2184
rect 29970 2128 29998 2184
rect 30158 2128 30186 2184
rect 30622 2128 30650 2184
rect 30754 2128 30782 2184
rect 31218 2128 31246 2184
rect 31406 2128 31434 2184
rect 31870 2128 31898 2184
rect 32002 2128 32030 2184
rect 32466 2128 32494 2184
rect 32654 2128 32682 2184
rect 33118 2128 33146 2184
rect 33250 2128 33278 2184
rect 33714 2128 33742 2184
rect 33902 2128 33930 2184
rect 34366 2128 34394 2184
rect 34498 2128 34526 2184
rect 34962 2128 34990 2184
rect 35150 2128 35178 2184
rect 35614 2128 35642 2184
rect 35746 2128 35774 2184
rect 36210 2128 36238 2184
rect 36398 2128 36426 2184
rect 36862 2128 36890 2184
rect 36994 2128 37022 2184
rect 37458 2128 37486 2184
rect 37646 2128 37674 2184
rect 38110 2128 38138 2184
rect 38242 2128 38270 2184
rect 38706 2128 38734 2184
rect 38894 2128 38922 2184
rect 39358 2128 39386 2184
rect 39490 2128 39518 2184
rect 39954 2128 39982 2184
rect 40142 2128 40170 2184
rect 40606 2128 40634 2184
rect 40738 2128 40766 2184
rect 41202 2128 41230 2184
rect 41390 2128 41418 2184
rect 41854 2128 41882 2184
rect 41986 2128 42014 2184
rect 42450 2128 42478 2184
rect 42638 2128 42666 2184
rect 43102 2128 43130 2184
rect 43234 2128 43262 2184
rect 43698 2128 43726 2184
rect 43886 2128 43914 2184
rect 44350 2128 44378 2184
rect 44482 2128 44510 2184
rect 44946 2128 44974 2184
rect 45134 2128 45162 2184
rect 45598 2128 45626 2184
rect 45730 2128 45758 2184
rect 46194 2128 46222 2184
rect 46382 2128 46410 2184
rect 46846 2128 46874 2184
rect 46978 2128 47006 2184
rect 47442 2128 47470 2184
rect 47630 2128 47658 2184
rect 48094 2128 48122 2184
rect 48226 2128 48254 2184
rect 48690 2128 48718 2184
rect 48878 2128 48906 2184
rect 49342 2128 49370 2184
rect 49474 2128 49502 2184
rect 49938 2128 49966 2184
rect 50126 2128 50154 2184
rect 50590 2128 50618 2184
rect 50722 2128 50750 2184
rect 51186 2128 51214 2184
rect 51374 2128 51402 2184
rect 51838 2128 51866 2184
rect 51970 2128 51998 2184
rect 52434 2128 52462 2184
rect 52622 2128 52650 2184
rect 53086 2128 53114 2184
rect 53218 2128 53246 2184
rect 53682 2128 53710 2184
rect 53870 2128 53898 2184
rect 54334 2128 54362 2184
rect 54466 2128 54494 2184
rect 54930 2128 54958 2184
rect 55118 2128 55146 2184
rect 55582 2128 55610 2184
rect 55714 2128 55742 2184
rect 56178 2128 56206 2184
rect 56366 2128 56394 2184
rect 56830 2128 56858 2184
rect 56962 2128 56990 2184
rect 57426 2128 57454 2184
rect 57614 2128 57642 2184
rect 58078 2128 58106 2184
rect 58210 2128 58238 2184
rect 58674 2128 58702 2184
rect 58862 2128 58890 2184
rect 59326 2128 59354 2184
rect 59458 2128 59486 2184
rect 59922 2128 59950 2184
rect 60110 2128 60138 2184
rect 60574 2128 60602 2184
rect 60706 2128 60734 2184
rect 61170 2128 61198 2184
rect 61358 2128 61386 2184
rect 61822 2128 61850 2184
rect 61954 2128 61982 2184
rect 62418 2128 62446 2184
rect 62606 2128 62634 2184
rect 63070 2128 63098 2184
rect 63202 2128 63230 2184
rect 63666 2128 63694 2184
rect 63854 2128 63882 2184
rect 64318 2128 64346 2184
rect 64450 2128 64478 2184
rect 64914 2128 64942 2184
rect 65102 2128 65130 2184
rect 65566 2128 65594 2184
rect 65698 2128 65726 2184
rect 66162 2128 66190 2184
rect 66350 2128 66378 2184
rect 66814 2128 66842 2184
rect 66946 2128 66974 2184
rect 67410 2128 67438 2184
rect 67598 2128 67626 2184
rect 68062 2128 68090 2184
rect 68194 2128 68222 2184
rect 68658 2128 68686 2184
rect 68846 2128 68874 2184
rect 69310 2128 69338 2184
rect 69442 2128 69470 2184
rect 69906 2128 69934 2184
rect 70094 2128 70122 2184
rect 70558 2128 70586 2184
rect 70690 2128 70718 2184
rect 71154 2128 71182 2184
rect 71342 2128 71370 2184
rect 71806 2128 71834 2184
rect 71938 2128 71966 2184
rect 72402 2128 72430 2184
rect 72590 2128 72618 2184
rect 73054 2128 73082 2184
rect 73186 2128 73214 2184
rect 73650 2128 73678 2184
rect 73838 2128 73866 2184
rect 74302 2128 74330 2184
rect 74434 2128 74462 2184
rect 74898 2128 74926 2184
rect 75086 2128 75114 2184
rect 75550 2128 75578 2184
rect 75682 2128 75710 2184
rect 76146 2128 76174 2184
rect 76334 2128 76362 2184
rect 76798 2128 76826 2184
rect 76930 2128 76958 2184
rect 77394 2128 77422 2184
rect 77582 2128 77610 2184
rect 78046 2128 78074 2184
rect 78178 2128 78206 2184
rect 78642 2128 78670 2184
rect 78830 2128 78858 2184
rect 79294 2128 79322 2184
rect 79426 2128 79454 2184
rect 79890 2128 79918 2184
rect 80078 2128 80106 2184
rect 80542 2128 80570 2184
rect 80674 2128 80702 2184
rect 81138 2128 81166 2184
rect 1454 248 1482 868
rect 1654 376 1718 428
rect 1918 124 1946 868
rect 2050 124 2078 868
rect 2278 500 2342 552
rect 2514 248 2542 868
rect 2702 248 2730 868
rect 2902 624 2966 676
rect 3166 124 3194 868
rect 3298 124 3326 868
rect 3526 748 3590 800
rect 3762 248 3790 868
rect 3950 248 3978 868
rect 4150 376 4214 428
rect 4414 124 4442 868
rect 4546 124 4574 868
rect 4774 500 4838 552
rect 5010 248 5038 868
rect 5198 248 5226 868
rect 5398 624 5462 676
rect 5662 124 5690 868
rect 5794 124 5822 868
rect 6022 748 6086 800
rect 6258 248 6286 868
rect 6446 248 6474 868
rect 6646 376 6710 428
rect 6910 124 6938 868
rect 7042 124 7070 868
rect 7270 500 7334 552
rect 7506 248 7534 868
rect 7694 248 7722 868
rect 7894 624 7958 676
rect 8158 124 8186 868
rect 8290 124 8318 868
rect 8518 748 8582 800
rect 8754 248 8782 868
rect 8942 248 8970 868
rect 9142 376 9206 428
rect 9406 124 9434 868
rect 9538 124 9566 868
rect 9766 500 9830 552
rect 10002 248 10030 868
rect 10190 248 10218 868
rect 10390 624 10454 676
rect 10654 124 10682 868
rect 10786 124 10814 868
rect 11014 748 11078 800
rect 11250 248 11278 868
rect 11438 248 11466 868
rect 11638 376 11702 428
rect 11902 124 11930 868
rect 12034 124 12062 868
rect 12262 500 12326 552
rect 12498 248 12526 868
rect 12686 248 12714 868
rect 12886 624 12950 676
rect 13150 124 13178 868
rect 13282 124 13310 868
rect 13510 748 13574 800
rect 13746 248 13774 868
rect 13934 248 13962 868
rect 14134 376 14198 428
rect 14398 124 14426 868
rect 14530 124 14558 868
rect 14758 500 14822 552
rect 14994 248 15022 868
rect 15182 248 15210 868
rect 15382 624 15446 676
rect 15646 124 15674 868
rect 15778 124 15806 868
rect 16006 748 16070 800
rect 16242 248 16270 868
rect 16430 248 16458 868
rect 16630 376 16694 428
rect 16894 124 16922 868
rect 17026 124 17054 868
rect 17254 500 17318 552
rect 17490 248 17518 868
rect 17678 248 17706 868
rect 17878 624 17942 676
rect 18142 124 18170 868
rect 18274 124 18302 868
rect 18502 748 18566 800
rect 18738 248 18766 868
rect 18926 248 18954 868
rect 19126 376 19190 428
rect 19390 124 19418 868
rect 19522 124 19550 868
rect 19750 500 19814 552
rect 19986 248 20014 868
rect 20174 248 20202 868
rect 20374 624 20438 676
rect 20638 124 20666 868
rect 20770 124 20798 868
rect 20998 748 21062 800
rect 21234 248 21262 868
rect 21422 248 21450 868
rect 21622 376 21686 428
rect 21886 124 21914 868
rect 22018 124 22046 868
rect 22246 500 22310 552
rect 22482 248 22510 868
rect 22670 248 22698 868
rect 22870 624 22934 676
rect 23134 124 23162 868
rect 23266 124 23294 868
rect 23494 748 23558 800
rect 23730 248 23758 868
rect 23918 248 23946 868
rect 24118 376 24182 428
rect 24382 124 24410 868
rect 24514 124 24542 868
rect 24742 500 24806 552
rect 24978 248 25006 868
rect 25166 248 25194 868
rect 25366 624 25430 676
rect 25630 124 25658 868
rect 25762 124 25790 868
rect 25990 748 26054 800
rect 26226 248 26254 868
rect 26414 248 26442 868
rect 26614 376 26678 428
rect 26878 124 26906 868
rect 27010 124 27038 868
rect 27238 500 27302 552
rect 27474 248 27502 868
rect 27662 248 27690 868
rect 27862 624 27926 676
rect 28126 124 28154 868
rect 28258 124 28286 868
rect 28486 748 28550 800
rect 28722 248 28750 868
rect 28910 248 28938 868
rect 29110 376 29174 428
rect 29374 124 29402 868
rect 29506 124 29534 868
rect 29734 500 29798 552
rect 29970 248 29998 868
rect 30158 248 30186 868
rect 30358 624 30422 676
rect 30622 124 30650 868
rect 30754 124 30782 868
rect 30982 748 31046 800
rect 31218 248 31246 868
rect 31406 248 31434 868
rect 31606 376 31670 428
rect 31870 124 31898 868
rect 32002 124 32030 868
rect 32230 500 32294 552
rect 32466 248 32494 868
rect 32654 248 32682 868
rect 32854 624 32918 676
rect 33118 124 33146 868
rect 33250 124 33278 868
rect 33478 748 33542 800
rect 33714 248 33742 868
rect 33902 248 33930 868
rect 34102 376 34166 428
rect 34366 124 34394 868
rect 34498 124 34526 868
rect 34726 500 34790 552
rect 34962 248 34990 868
rect 35150 248 35178 868
rect 35350 624 35414 676
rect 35614 124 35642 868
rect 35746 124 35774 868
rect 35974 748 36038 800
rect 36210 248 36238 868
rect 36398 248 36426 868
rect 36598 376 36662 428
rect 36862 124 36890 868
rect 36994 124 37022 868
rect 37222 500 37286 552
rect 37458 248 37486 868
rect 37646 248 37674 868
rect 37846 624 37910 676
rect 38110 124 38138 868
rect 38242 124 38270 868
rect 38470 748 38534 800
rect 38706 248 38734 868
rect 38894 248 38922 868
rect 39094 376 39158 428
rect 39358 124 39386 868
rect 39490 124 39518 868
rect 39718 500 39782 552
rect 39954 248 39982 868
rect 40142 248 40170 868
rect 40342 624 40406 676
rect 40606 124 40634 868
rect 40738 124 40766 868
rect 40966 748 41030 800
rect 41202 248 41230 868
rect 41390 248 41418 868
rect 41590 376 41654 428
rect 41854 124 41882 868
rect 41986 124 42014 868
rect 42214 500 42278 552
rect 42450 248 42478 868
rect 42638 248 42666 868
rect 42838 624 42902 676
rect 43102 124 43130 868
rect 43234 124 43262 868
rect 43462 748 43526 800
rect 43698 248 43726 868
rect 43886 248 43914 868
rect 44086 376 44150 428
rect 44350 124 44378 868
rect 44482 124 44510 868
rect 44710 500 44774 552
rect 44946 248 44974 868
rect 45134 248 45162 868
rect 45334 624 45398 676
rect 45598 124 45626 868
rect 45730 124 45758 868
rect 45958 748 46022 800
rect 46194 248 46222 868
rect 46382 248 46410 868
rect 46582 376 46646 428
rect 46846 124 46874 868
rect 46978 124 47006 868
rect 47206 500 47270 552
rect 47442 248 47470 868
rect 47630 248 47658 868
rect 47830 624 47894 676
rect 48094 124 48122 868
rect 48226 124 48254 868
rect 48454 748 48518 800
rect 48690 248 48718 868
rect 48878 248 48906 868
rect 49078 376 49142 428
rect 49342 124 49370 868
rect 49474 124 49502 868
rect 49702 500 49766 552
rect 49938 248 49966 868
rect 50126 248 50154 868
rect 50326 624 50390 676
rect 50590 124 50618 868
rect 50722 124 50750 868
rect 50950 748 51014 800
rect 51186 248 51214 868
rect 51374 248 51402 868
rect 51574 376 51638 428
rect 51838 124 51866 868
rect 51970 124 51998 868
rect 52198 500 52262 552
rect 52434 248 52462 868
rect 52622 248 52650 868
rect 52822 624 52886 676
rect 53086 124 53114 868
rect 53218 124 53246 868
rect 53446 748 53510 800
rect 53682 248 53710 868
rect 53870 248 53898 868
rect 54070 376 54134 428
rect 54334 124 54362 868
rect 54466 124 54494 868
rect 54694 500 54758 552
rect 54930 248 54958 868
rect 55118 248 55146 868
rect 55318 624 55382 676
rect 55582 124 55610 868
rect 55714 124 55742 868
rect 55942 748 56006 800
rect 56178 248 56206 868
rect 56366 248 56394 868
rect 56566 376 56630 428
rect 56830 124 56858 868
rect 56962 124 56990 868
rect 57190 500 57254 552
rect 57426 248 57454 868
rect 57614 248 57642 868
rect 57814 624 57878 676
rect 58078 124 58106 868
rect 58210 124 58238 868
rect 58438 748 58502 800
rect 58674 248 58702 868
rect 58862 248 58890 868
rect 59062 376 59126 428
rect 59326 124 59354 868
rect 59458 124 59486 868
rect 59686 500 59750 552
rect 59922 248 59950 868
rect 60110 248 60138 868
rect 60310 624 60374 676
rect 60574 124 60602 868
rect 60706 124 60734 868
rect 60934 748 60998 800
rect 61170 248 61198 868
rect 61358 248 61386 868
rect 61558 376 61622 428
rect 61822 124 61850 868
rect 61954 124 61982 868
rect 62182 500 62246 552
rect 62418 248 62446 868
rect 62606 248 62634 868
rect 62806 624 62870 676
rect 63070 124 63098 868
rect 63202 124 63230 868
rect 63430 748 63494 800
rect 63666 248 63694 868
rect 63854 248 63882 868
rect 64054 376 64118 428
rect 64318 124 64346 868
rect 64450 124 64478 868
rect 64678 500 64742 552
rect 64914 248 64942 868
rect 65102 248 65130 868
rect 65302 624 65366 676
rect 65566 124 65594 868
rect 65698 124 65726 868
rect 65926 748 65990 800
rect 66162 248 66190 868
rect 66350 248 66378 868
rect 66550 376 66614 428
rect 66814 124 66842 868
rect 66946 124 66974 868
rect 67174 500 67238 552
rect 67410 248 67438 868
rect 67598 248 67626 868
rect 67798 624 67862 676
rect 68062 124 68090 868
rect 68194 124 68222 868
rect 68422 748 68486 800
rect 68658 248 68686 868
rect 68846 248 68874 868
rect 69046 376 69110 428
rect 69310 124 69338 868
rect 69442 124 69470 868
rect 69670 500 69734 552
rect 69906 248 69934 868
rect 70094 248 70122 868
rect 70294 624 70358 676
rect 70558 124 70586 868
rect 70690 124 70718 868
rect 70918 748 70982 800
rect 71154 248 71182 868
rect 71342 248 71370 868
rect 71542 376 71606 428
rect 71806 124 71834 868
rect 71938 124 71966 868
rect 72166 500 72230 552
rect 72402 248 72430 868
rect 72590 248 72618 868
rect 72790 624 72854 676
rect 73054 124 73082 868
rect 73186 124 73214 868
rect 73414 748 73478 800
rect 73650 248 73678 868
rect 73838 248 73866 868
rect 74038 376 74102 428
rect 74302 124 74330 868
rect 74434 124 74462 868
rect 74662 500 74726 552
rect 74898 248 74926 868
rect 75086 248 75114 868
rect 75286 624 75350 676
rect 75550 124 75578 868
rect 75682 124 75710 868
rect 75910 748 75974 800
rect 76146 248 76174 868
rect 76334 248 76362 868
rect 76534 376 76598 428
rect 76798 124 76826 868
rect 76930 124 76958 868
rect 77158 500 77222 552
rect 77394 248 77422 868
rect 77582 248 77610 868
rect 77782 624 77846 676
rect 78046 124 78074 868
rect 78178 124 78206 868
rect 78406 748 78470 800
rect 78642 248 78670 868
rect 78830 248 78858 868
rect 79030 376 79094 428
rect 79294 124 79322 868
rect 79426 124 79454 868
rect 79654 500 79718 552
rect 79890 248 79918 868
rect 80078 248 80106 868
rect 80278 624 80342 676
rect 80542 124 80570 868
rect 80674 124 80702 868
rect 80902 748 80966 800
rect 81138 248 81166 868
<< metal2 >>
rect 3530 750 3586 798
rect 6026 750 6082 798
rect 8522 750 8578 798
rect 11018 750 11074 798
rect 13514 750 13570 798
rect 16010 750 16066 798
rect 18506 750 18562 798
rect 21002 750 21058 798
rect 23498 750 23554 798
rect 25994 750 26050 798
rect 28490 750 28546 798
rect 30986 750 31042 798
rect 33482 750 33538 798
rect 35978 750 36034 798
rect 38474 750 38530 798
rect 40970 750 41026 798
rect 43466 750 43522 798
rect 45962 750 46018 798
rect 48458 750 48514 798
rect 50954 750 51010 798
rect 53450 750 53506 798
rect 55946 750 56002 798
rect 58442 750 58498 798
rect 60938 750 60994 798
rect 63434 750 63490 798
rect 65930 750 65986 798
rect 68426 750 68482 798
rect 70922 750 70978 798
rect 73418 750 73474 798
rect 75914 750 75970 798
rect 78410 750 78466 798
rect 80906 750 80962 798
rect 2906 626 2962 674
rect 5402 626 5458 674
rect 7898 626 7954 674
rect 10394 626 10450 674
rect 12890 626 12946 674
rect 15386 626 15442 674
rect 17882 626 17938 674
rect 20378 626 20434 674
rect 22874 626 22930 674
rect 25370 626 25426 674
rect 27866 626 27922 674
rect 30362 626 30418 674
rect 32858 626 32914 674
rect 35354 626 35410 674
rect 37850 626 37906 674
rect 40346 626 40402 674
rect 42842 626 42898 674
rect 45338 626 45394 674
rect 47834 626 47890 674
rect 50330 626 50386 674
rect 52826 626 52882 674
rect 55322 626 55378 674
rect 57818 626 57874 674
rect 60314 626 60370 674
rect 62810 626 62866 674
rect 65306 626 65362 674
rect 67802 626 67858 674
rect 70298 626 70354 674
rect 72794 626 72850 674
rect 75290 626 75346 674
rect 77786 626 77842 674
rect 80282 626 80338 674
rect 2282 502 2338 550
rect 4778 502 4834 550
rect 7274 502 7330 550
rect 9770 502 9826 550
rect 12266 502 12322 550
rect 14762 502 14818 550
rect 17258 502 17314 550
rect 19754 502 19810 550
rect 22250 502 22306 550
rect 24746 502 24802 550
rect 27242 502 27298 550
rect 29738 502 29794 550
rect 32234 502 32290 550
rect 34730 502 34786 550
rect 37226 502 37282 550
rect 39722 502 39778 550
rect 42218 502 42274 550
rect 44714 502 44770 550
rect 47210 502 47266 550
rect 49706 502 49762 550
rect 52202 502 52258 550
rect 54698 502 54754 550
rect 57194 502 57250 550
rect 59690 502 59746 550
rect 62186 502 62242 550
rect 64682 502 64738 550
rect 67178 502 67234 550
rect 69674 502 69730 550
rect 72170 502 72226 550
rect 74666 502 74722 550
rect 77162 502 77218 550
rect 79658 502 79714 550
rect 1658 378 1714 426
rect 4154 378 4210 426
rect 6650 378 6706 426
rect 9146 378 9202 426
rect 11642 378 11698 426
rect 14138 378 14194 426
rect 16634 378 16690 426
rect 19130 378 19186 426
rect 21626 378 21682 426
rect 24122 378 24178 426
rect 26618 378 26674 426
rect 29114 378 29170 426
rect 31610 378 31666 426
rect 34106 378 34162 426
rect 36602 378 36658 426
rect 39098 378 39154 426
rect 41594 378 41650 426
rect 44090 378 44146 426
rect 46586 378 46642 426
rect 49082 378 49138 426
rect 51578 378 51634 426
rect 54074 378 54130 426
rect 56570 378 56626 426
rect 59066 378 59122 426
rect 61562 378 61618 426
rect 64058 378 64114 426
rect 66554 378 66610 426
rect 69050 378 69106 426
rect 71546 378 71602 426
rect 74042 378 74098 426
rect 76538 378 76594 426
rect 79034 378 79090 426
rect 1440 224 1496 272
rect 2500 224 2556 272
rect 2688 224 2744 272
rect 3748 224 3804 272
rect 3936 224 3992 272
rect 4996 224 5052 272
rect 5184 224 5240 272
rect 6244 224 6300 272
rect 6432 224 6488 272
rect 7492 224 7548 272
rect 7680 224 7736 272
rect 8740 224 8796 272
rect 8928 224 8984 272
rect 9988 224 10044 272
rect 10176 224 10232 272
rect 11236 224 11292 272
rect 11424 224 11480 272
rect 12484 224 12540 272
rect 12672 224 12728 272
rect 13732 224 13788 272
rect 13920 224 13976 272
rect 14980 224 15036 272
rect 15168 224 15224 272
rect 16228 224 16284 272
rect 16416 224 16472 272
rect 17476 224 17532 272
rect 17664 224 17720 272
rect 18724 224 18780 272
rect 18912 224 18968 272
rect 19972 224 20028 272
rect 20160 224 20216 272
rect 21220 224 21276 272
rect 21408 224 21464 272
rect 22468 224 22524 272
rect 22656 224 22712 272
rect 23716 224 23772 272
rect 23904 224 23960 272
rect 24964 224 25020 272
rect 25152 224 25208 272
rect 26212 224 26268 272
rect 26400 224 26456 272
rect 27460 224 27516 272
rect 27648 224 27704 272
rect 28708 224 28764 272
rect 28896 224 28952 272
rect 29956 224 30012 272
rect 30144 224 30200 272
rect 31204 224 31260 272
rect 31392 224 31448 272
rect 32452 224 32508 272
rect 32640 224 32696 272
rect 33700 224 33756 272
rect 33888 224 33944 272
rect 34948 224 35004 272
rect 35136 224 35192 272
rect 36196 224 36252 272
rect 36384 224 36440 272
rect 37444 224 37500 272
rect 37632 224 37688 272
rect 38692 224 38748 272
rect 38880 224 38936 272
rect 39940 224 39996 272
rect 40128 224 40184 272
rect 41188 224 41244 272
rect 41376 224 41432 272
rect 42436 224 42492 272
rect 42624 224 42680 272
rect 43684 224 43740 272
rect 43872 224 43928 272
rect 44932 224 44988 272
rect 45120 224 45176 272
rect 46180 224 46236 272
rect 46368 224 46424 272
rect 47428 224 47484 272
rect 47616 224 47672 272
rect 48676 224 48732 272
rect 48864 224 48920 272
rect 49924 224 49980 272
rect 50112 224 50168 272
rect 51172 224 51228 272
rect 51360 224 51416 272
rect 52420 224 52476 272
rect 52608 224 52664 272
rect 53668 224 53724 272
rect 53856 224 53912 272
rect 54916 224 54972 272
rect 55104 224 55160 272
rect 56164 224 56220 272
rect 56352 224 56408 272
rect 57412 224 57468 272
rect 57600 224 57656 272
rect 58660 224 58716 272
rect 58848 224 58904 272
rect 59908 224 59964 272
rect 60096 224 60152 272
rect 61156 224 61212 272
rect 61344 224 61400 272
rect 62404 224 62460 272
rect 62592 224 62648 272
rect 63652 224 63708 272
rect 63840 224 63896 272
rect 64900 224 64956 272
rect 65088 224 65144 272
rect 66148 224 66204 272
rect 66336 224 66392 272
rect 67396 224 67452 272
rect 67584 224 67640 272
rect 68644 224 68700 272
rect 68832 224 68888 272
rect 69892 224 69948 272
rect 70080 224 70136 272
rect 71140 224 71196 272
rect 71328 224 71384 272
rect 72388 224 72444 272
rect 72576 224 72632 272
rect 73636 224 73692 272
rect 73824 224 73880 272
rect 74884 224 74940 272
rect 75072 224 75128 272
rect 76132 224 76188 272
rect 76320 224 76376 272
rect 77380 224 77436 272
rect 77568 224 77624 272
rect 78628 224 78684 272
rect 78816 224 78872 272
rect 79876 224 79932 272
rect 80064 224 80120 272
rect 81124 224 81180 272
rect 1904 100 1960 148
rect 2036 100 2092 148
rect 3152 100 3208 148
rect 3284 100 3340 148
rect 4400 100 4456 148
rect 4532 100 4588 148
rect 5648 100 5704 148
rect 5780 100 5836 148
rect 6896 100 6952 148
rect 7028 100 7084 148
rect 8144 100 8200 148
rect 8276 100 8332 148
rect 9392 100 9448 148
rect 9524 100 9580 148
rect 10640 100 10696 148
rect 10772 100 10828 148
rect 11888 100 11944 148
rect 12020 100 12076 148
rect 13136 100 13192 148
rect 13268 100 13324 148
rect 14384 100 14440 148
rect 14516 100 14572 148
rect 15632 100 15688 148
rect 15764 100 15820 148
rect 16880 100 16936 148
rect 17012 100 17068 148
rect 18128 100 18184 148
rect 18260 100 18316 148
rect 19376 100 19432 148
rect 19508 100 19564 148
rect 20624 100 20680 148
rect 20756 100 20812 148
rect 21872 100 21928 148
rect 22004 100 22060 148
rect 23120 100 23176 148
rect 23252 100 23308 148
rect 24368 100 24424 148
rect 24500 100 24556 148
rect 25616 100 25672 148
rect 25748 100 25804 148
rect 26864 100 26920 148
rect 26996 100 27052 148
rect 28112 100 28168 148
rect 28244 100 28300 148
rect 29360 100 29416 148
rect 29492 100 29548 148
rect 30608 100 30664 148
rect 30740 100 30796 148
rect 31856 100 31912 148
rect 31988 100 32044 148
rect 33104 100 33160 148
rect 33236 100 33292 148
rect 34352 100 34408 148
rect 34484 100 34540 148
rect 35600 100 35656 148
rect 35732 100 35788 148
rect 36848 100 36904 148
rect 36980 100 37036 148
rect 38096 100 38152 148
rect 38228 100 38284 148
rect 39344 100 39400 148
rect 39476 100 39532 148
rect 40592 100 40648 148
rect 40724 100 40780 148
rect 41840 100 41896 148
rect 41972 100 42028 148
rect 43088 100 43144 148
rect 43220 100 43276 148
rect 44336 100 44392 148
rect 44468 100 44524 148
rect 45584 100 45640 148
rect 45716 100 45772 148
rect 46832 100 46888 148
rect 46964 100 47020 148
rect 48080 100 48136 148
rect 48212 100 48268 148
rect 49328 100 49384 148
rect 49460 100 49516 148
rect 50576 100 50632 148
rect 50708 100 50764 148
rect 51824 100 51880 148
rect 51956 100 52012 148
rect 53072 100 53128 148
rect 53204 100 53260 148
rect 54320 100 54376 148
rect 54452 100 54508 148
rect 55568 100 55624 148
rect 55700 100 55756 148
rect 56816 100 56872 148
rect 56948 100 57004 148
rect 58064 100 58120 148
rect 58196 100 58252 148
rect 59312 100 59368 148
rect 59444 100 59500 148
rect 60560 100 60616 148
rect 60692 100 60748 148
rect 61808 100 61864 148
rect 61940 100 61996 148
rect 63056 100 63112 148
rect 63188 100 63244 148
rect 64304 100 64360 148
rect 64436 100 64492 148
rect 65552 100 65608 148
rect 65684 100 65740 148
rect 66800 100 66856 148
rect 66932 100 66988 148
rect 68048 100 68104 148
rect 68180 100 68236 148
rect 69296 100 69352 148
rect 69428 100 69484 148
rect 70544 100 70600 148
rect 70676 100 70732 148
rect 71792 100 71848 148
rect 71924 100 71980 148
rect 73040 100 73096 148
rect 73172 100 73228 148
rect 74288 100 74344 148
rect 74420 100 74476 148
rect 75536 100 75592 148
rect 75668 100 75724 148
rect 76784 100 76840 148
rect 76916 100 76972 148
rect 78032 100 78088 148
rect 78164 100 78220 148
rect 79280 100 79336 148
rect 79412 100 79468 148
rect 80528 100 80584 148
rect 80660 100 80716 148
<< metal3 >>
rect 1949 1482 2047 1580
rect 3197 1482 3295 1580
rect 4445 1482 4543 1580
rect 5693 1482 5791 1580
rect 6941 1482 7039 1580
rect 8189 1482 8287 1580
rect 9437 1482 9535 1580
rect 10685 1482 10783 1580
rect 11933 1482 12031 1580
rect 13181 1482 13279 1580
rect 14429 1482 14527 1580
rect 15677 1482 15775 1580
rect 16925 1482 17023 1580
rect 18173 1482 18271 1580
rect 19421 1482 19519 1580
rect 20669 1482 20767 1580
rect 21917 1482 22015 1580
rect 23165 1482 23263 1580
rect 24413 1482 24511 1580
rect 25661 1482 25759 1580
rect 26909 1482 27007 1580
rect 28157 1482 28255 1580
rect 29405 1482 29503 1580
rect 30653 1482 30751 1580
rect 31901 1482 31999 1580
rect 33149 1482 33247 1580
rect 34397 1482 34495 1580
rect 35645 1482 35743 1580
rect 36893 1482 36991 1580
rect 38141 1482 38239 1580
rect 39389 1482 39487 1580
rect 40637 1482 40735 1580
rect 41885 1482 41983 1580
rect 43133 1482 43231 1580
rect 44381 1482 44479 1580
rect 45629 1482 45727 1580
rect 46877 1482 46975 1580
rect 48125 1482 48223 1580
rect 49373 1482 49471 1580
rect 50621 1482 50719 1580
rect 51869 1482 51967 1580
rect 53117 1482 53215 1580
rect 54365 1482 54463 1580
rect 55613 1482 55711 1580
rect 56861 1482 56959 1580
rect 58109 1482 58207 1580
rect 59357 1482 59455 1580
rect 60605 1482 60703 1580
rect 61853 1482 61951 1580
rect 63101 1482 63199 1580
rect 64349 1482 64447 1580
rect 65597 1482 65695 1580
rect 66845 1482 66943 1580
rect 68093 1482 68191 1580
rect 69341 1482 69439 1580
rect 70589 1482 70687 1580
rect 71837 1482 71935 1580
rect 73085 1482 73183 1580
rect 74333 1482 74431 1580
rect 75581 1482 75679 1580
rect 76829 1482 76927 1580
rect 78077 1482 78175 1580
rect 79325 1482 79423 1580
rect 80573 1482 80671 1580
rect 0 744 81246 804
rect 0 620 81246 680
rect 0 496 81246 556
rect 0 372 81246 432
rect 1468 218 3776 278
rect 3964 218 6272 278
rect 6460 218 8768 278
rect 8956 218 11264 278
rect 11452 218 13760 278
rect 13948 218 16256 278
rect 16444 218 18752 278
rect 18940 218 21248 278
rect 21436 218 23744 278
rect 23932 218 26240 278
rect 26428 218 28736 278
rect 28924 218 31232 278
rect 31420 218 33728 278
rect 33916 218 36224 278
rect 36412 218 38720 278
rect 38908 218 41216 278
rect 41404 218 43712 278
rect 43900 218 46208 278
rect 46396 218 48704 278
rect 48892 218 51200 278
rect 51388 218 53696 278
rect 53884 218 56192 278
rect 56380 218 58688 278
rect 58876 218 61184 278
rect 61372 218 63680 278
rect 63868 218 66176 278
rect 66364 218 68672 278
rect 68860 218 71168 278
rect 71356 218 73664 278
rect 73852 218 76160 278
rect 76348 218 78656 278
rect 78844 218 81152 278
rect 1932 94 3312 154
rect 4428 94 5808 154
rect 6924 94 8304 154
rect 9420 94 10800 154
rect 11916 94 13296 154
rect 14412 94 15792 154
rect 16908 94 18288 154
rect 19404 94 20784 154
rect 21900 94 23280 154
rect 24396 94 25776 154
rect 26892 94 28272 154
rect 29388 94 30768 154
rect 31884 94 33264 154
rect 34380 94 35760 154
rect 36876 94 38256 154
rect 39372 94 40752 154
rect 41868 94 43248 154
rect 44364 94 45744 154
rect 46860 94 48240 154
rect 49356 94 50736 154
rect 51852 94 53232 154
rect 54348 94 55728 154
rect 56844 94 58224 154
rect 59340 94 60720 154
rect 61836 94 63216 154
rect 64332 94 65712 154
rect 66828 94 68208 154
rect 69324 94 70704 154
rect 71820 94 73200 154
rect 74316 94 75696 154
rect 76812 94 78192 154
rect 79308 94 80688 154
use contact_25  contact_25_255
timestamp 1624494425
transform 1 0 1436 0 1 216
box 0 0 64 64
use contact_26  contact_26_255
timestamp 1624494425
transform 1 0 1435 0 1 211
box 0 0 66 74
use contact_25  contact_25_254
timestamp 1624494425
transform 1 0 1900 0 1 92
box 0 0 64 64
use contact_26  contact_26_254
timestamp 1624494425
transform 1 0 1899 0 1 87
box 0 0 66 74
use contact_25  contact_25_252
timestamp 1624494425
transform 1 0 2032 0 1 92
box 0 0 64 64
use contact_26  contact_26_252
timestamp 1624494425
transform 1 0 2031 0 1 87
box 0 0 66 74
use contact_23  contact_23_127
timestamp 1624494425
transform 1 0 1653 0 1 369
box 0 0 66 66
use contact_24  contact_24_127
timestamp 1624494425
transform 1 0 1657 0 1 369
box 0 0 58 66
use contact_25  contact_25_383
timestamp 1624494425
transform 1 0 1654 0 1 370
box 0 0 64 64
use contact_26  contact_26_383
timestamp 1624494425
transform 1 0 1653 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_127
timestamp 1624494425
transform 1 0 1374 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_126
timestamp 1624494425
transform -1 0 2622 0 1 868
box 65 0 675 1316
use contact_23  contact_23_126
timestamp 1624494425
transform 1 0 2277 0 1 493
box 0 0 66 66
use contact_24  contact_24_126
timestamp 1624494425
transform 1 0 2281 0 1 493
box 0 0 58 66
use contact_25  contact_25_253
timestamp 1624494425
transform 1 0 2496 0 1 216
box 0 0 64 64
use contact_25  contact_25_382
timestamp 1624494425
transform 1 0 2278 0 1 494
box 0 0 64 64
use contact_26  contact_26_253
timestamp 1624494425
transform 1 0 2495 0 1 211
box 0 0 66 74
use contact_26  contact_26_382
timestamp 1624494425
transform 1 0 2277 0 1 489
box 0 0 66 74
use contact_26  contact_26_381
timestamp 1624494425
transform 1 0 2901 0 1 613
box 0 0 66 74
use contact_26  contact_26_251
timestamp 1624494425
transform 1 0 2683 0 1 211
box 0 0 66 74
use contact_26  contact_26_250
timestamp 1624494425
transform 1 0 3147 0 1 87
box 0 0 66 74
use contact_25  contact_25_381
timestamp 1624494425
transform 1 0 2902 0 1 618
box 0 0 64 64
use contact_25  contact_25_251
timestamp 1624494425
transform 1 0 2684 0 1 216
box 0 0 64 64
use contact_25  contact_25_250
timestamp 1624494425
transform 1 0 3148 0 1 92
box 0 0 64 64
use contact_24  contact_24_125
timestamp 1624494425
transform 1 0 2905 0 1 617
box 0 0 58 66
use contact_23  contact_23_125
timestamp 1624494425
transform 1 0 2901 0 1 617
box 0 0 66 66
use column_mux_0  column_mux_0_125
timestamp 1624494425
transform 1 0 2622 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_124
timestamp 1624494425
transform -1 0 3870 0 1 868
box 65 0 675 1316
use contact_23  contact_23_124
timestamp 1624494425
transform 1 0 3525 0 1 741
box 0 0 66 66
use contact_24  contact_24_124
timestamp 1624494425
transform 1 0 3529 0 1 741
box 0 0 58 66
use contact_25  contact_25_248
timestamp 1624494425
transform 1 0 3280 0 1 92
box 0 0 64 64
use contact_25  contact_25_249
timestamp 1624494425
transform 1 0 3744 0 1 216
box 0 0 64 64
use contact_25  contact_25_380
timestamp 1624494425
transform 1 0 3526 0 1 742
box 0 0 64 64
use contact_26  contact_26_248
timestamp 1624494425
transform 1 0 3279 0 1 87
box 0 0 66 74
use contact_26  contact_26_249
timestamp 1624494425
transform 1 0 3743 0 1 211
box 0 0 66 74
use contact_26  contact_26_380
timestamp 1624494425
transform 1 0 3525 0 1 737
box 0 0 66 74
use contact_26  contact_26_379
timestamp 1624494425
transform 1 0 4149 0 1 365
box 0 0 66 74
use contact_26  contact_26_247
timestamp 1624494425
transform 1 0 3931 0 1 211
box 0 0 66 74
use contact_26  contact_26_246
timestamp 1624494425
transform 1 0 4395 0 1 87
box 0 0 66 74
use contact_25  contact_25_379
timestamp 1624494425
transform 1 0 4150 0 1 370
box 0 0 64 64
use contact_25  contact_25_247
timestamp 1624494425
transform 1 0 3932 0 1 216
box 0 0 64 64
use contact_25  contact_25_246
timestamp 1624494425
transform 1 0 4396 0 1 92
box 0 0 64 64
use contact_24  contact_24_123
timestamp 1624494425
transform 1 0 4153 0 1 369
box 0 0 58 66
use contact_23  contact_23_123
timestamp 1624494425
transform 1 0 4149 0 1 369
box 0 0 66 66
use column_mux_0  column_mux_0_123
timestamp 1624494425
transform 1 0 3870 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_122
timestamp 1624494425
transform -1 0 5118 0 1 868
box 65 0 675 1316
use contact_23  contact_23_122
timestamp 1624494425
transform 1 0 4773 0 1 493
box 0 0 66 66
use contact_24  contact_24_122
timestamp 1624494425
transform 1 0 4777 0 1 493
box 0 0 58 66
use contact_25  contact_25_244
timestamp 1624494425
transform 1 0 4528 0 1 92
box 0 0 64 64
use contact_25  contact_25_245
timestamp 1624494425
transform 1 0 4992 0 1 216
box 0 0 64 64
use contact_25  contact_25_378
timestamp 1624494425
transform 1 0 4774 0 1 494
box 0 0 64 64
use contact_26  contact_26_244
timestamp 1624494425
transform 1 0 4527 0 1 87
box 0 0 66 74
use contact_26  contact_26_245
timestamp 1624494425
transform 1 0 4991 0 1 211
box 0 0 66 74
use contact_26  contact_26_378
timestamp 1624494425
transform 1 0 4773 0 1 489
box 0 0 66 74
use contact_26  contact_26_377
timestamp 1624494425
transform 1 0 5397 0 1 613
box 0 0 66 74
use contact_26  contact_26_243
timestamp 1624494425
transform 1 0 5179 0 1 211
box 0 0 66 74
use contact_26  contact_26_242
timestamp 1624494425
transform 1 0 5643 0 1 87
box 0 0 66 74
use contact_25  contact_25_377
timestamp 1624494425
transform 1 0 5398 0 1 618
box 0 0 64 64
use contact_25  contact_25_243
timestamp 1624494425
transform 1 0 5180 0 1 216
box 0 0 64 64
use contact_25  contact_25_242
timestamp 1624494425
transform 1 0 5644 0 1 92
box 0 0 64 64
use contact_24  contact_24_121
timestamp 1624494425
transform 1 0 5401 0 1 617
box 0 0 58 66
use contact_23  contact_23_121
timestamp 1624494425
transform 1 0 5397 0 1 617
box 0 0 66 66
use column_mux_0  column_mux_0_121
timestamp 1624494425
transform 1 0 5118 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_120
timestamp 1624494425
transform -1 0 6366 0 1 868
box 65 0 675 1316
use contact_23  contact_23_120
timestamp 1624494425
transform 1 0 6021 0 1 741
box 0 0 66 66
use contact_24  contact_24_120
timestamp 1624494425
transform 1 0 6025 0 1 741
box 0 0 58 66
use contact_25  contact_25_240
timestamp 1624494425
transform 1 0 5776 0 1 92
box 0 0 64 64
use contact_25  contact_25_241
timestamp 1624494425
transform 1 0 6240 0 1 216
box 0 0 64 64
use contact_25  contact_25_376
timestamp 1624494425
transform 1 0 6022 0 1 742
box 0 0 64 64
use contact_26  contact_26_240
timestamp 1624494425
transform 1 0 5775 0 1 87
box 0 0 66 74
use contact_26  contact_26_241
timestamp 1624494425
transform 1 0 6239 0 1 211
box 0 0 66 74
use contact_26  contact_26_376
timestamp 1624494425
transform 1 0 6021 0 1 737
box 0 0 66 74
use contact_23  contact_23_119
timestamp 1624494425
transform 1 0 6645 0 1 369
box 0 0 66 66
use contact_24  contact_24_119
timestamp 1624494425
transform 1 0 6649 0 1 369
box 0 0 58 66
use contact_25  contact_25_238
timestamp 1624494425
transform 1 0 6892 0 1 92
box 0 0 64 64
use contact_25  contact_25_239
timestamp 1624494425
transform 1 0 6428 0 1 216
box 0 0 64 64
use contact_25  contact_25_375
timestamp 1624494425
transform 1 0 6646 0 1 370
box 0 0 64 64
use contact_26  contact_26_238
timestamp 1624494425
transform 1 0 6891 0 1 87
box 0 0 66 74
use contact_26  contact_26_239
timestamp 1624494425
transform 1 0 6427 0 1 211
box 0 0 66 74
use contact_26  contact_26_375
timestamp 1624494425
transform 1 0 6645 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_119
timestamp 1624494425
transform 1 0 6366 0 1 868
box 65 0 675 1316
use contact_23  contact_23_118
timestamp 1624494425
transform 1 0 7269 0 1 493
box 0 0 66 66
use contact_24  contact_24_118
timestamp 1624494425
transform 1 0 7273 0 1 493
box 0 0 58 66
use contact_25  contact_25_236
timestamp 1624494425
transform 1 0 7024 0 1 92
box 0 0 64 64
use contact_25  contact_25_237
timestamp 1624494425
transform 1 0 7488 0 1 216
box 0 0 64 64
use contact_25  contact_25_374
timestamp 1624494425
transform 1 0 7270 0 1 494
box 0 0 64 64
use contact_26  contact_26_236
timestamp 1624494425
transform 1 0 7023 0 1 87
box 0 0 66 74
use contact_26  contact_26_237
timestamp 1624494425
transform 1 0 7487 0 1 211
box 0 0 66 74
use contact_26  contact_26_374
timestamp 1624494425
transform 1 0 7269 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_118
timestamp 1624494425
transform -1 0 7614 0 1 868
box 65 0 675 1316
use contact_23  contact_23_117
timestamp 1624494425
transform 1 0 7893 0 1 617
box 0 0 66 66
use contact_24  contact_24_117
timestamp 1624494425
transform 1 0 7897 0 1 617
box 0 0 58 66
use contact_25  contact_25_234
timestamp 1624494425
transform 1 0 8140 0 1 92
box 0 0 64 64
use contact_25  contact_25_235
timestamp 1624494425
transform 1 0 7676 0 1 216
box 0 0 64 64
use contact_25  contact_25_373
timestamp 1624494425
transform 1 0 7894 0 1 618
box 0 0 64 64
use contact_26  contact_26_234
timestamp 1624494425
transform 1 0 8139 0 1 87
box 0 0 66 74
use contact_26  contact_26_235
timestamp 1624494425
transform 1 0 7675 0 1 211
box 0 0 66 74
use contact_26  contact_26_373
timestamp 1624494425
transform 1 0 7893 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_117
timestamp 1624494425
transform 1 0 7614 0 1 868
box 65 0 675 1316
use contact_23  contact_23_116
timestamp 1624494425
transform 1 0 8517 0 1 741
box 0 0 66 66
use contact_24  contact_24_116
timestamp 1624494425
transform 1 0 8521 0 1 741
box 0 0 58 66
use contact_25  contact_25_232
timestamp 1624494425
transform 1 0 8272 0 1 92
box 0 0 64 64
use contact_25  contact_25_233
timestamp 1624494425
transform 1 0 8736 0 1 216
box 0 0 64 64
use contact_25  contact_25_372
timestamp 1624494425
transform 1 0 8518 0 1 742
box 0 0 64 64
use contact_26  contact_26_232
timestamp 1624494425
transform 1 0 8271 0 1 87
box 0 0 66 74
use contact_26  contact_26_233
timestamp 1624494425
transform 1 0 8735 0 1 211
box 0 0 66 74
use contact_26  contact_26_372
timestamp 1624494425
transform 1 0 8517 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_116
timestamp 1624494425
transform -1 0 8862 0 1 868
box 65 0 675 1316
use contact_23  contact_23_115
timestamp 1624494425
transform 1 0 9141 0 1 369
box 0 0 66 66
use contact_24  contact_24_115
timestamp 1624494425
transform 1 0 9145 0 1 369
box 0 0 58 66
use contact_25  contact_25_231
timestamp 1624494425
transform 1 0 8924 0 1 216
box 0 0 64 64
use contact_25  contact_25_371
timestamp 1624494425
transform 1 0 9142 0 1 370
box 0 0 64 64
use contact_26  contact_26_231
timestamp 1624494425
transform 1 0 8923 0 1 211
box 0 0 66 74
use contact_26  contact_26_371
timestamp 1624494425
transform 1 0 9141 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_115
timestamp 1624494425
transform 1 0 8862 0 1 868
box 65 0 675 1316
use contact_25  contact_25_228
timestamp 1624494425
transform 1 0 9520 0 1 92
box 0 0 64 64
use contact_25  contact_25_230
timestamp 1624494425
transform 1 0 9388 0 1 92
box 0 0 64 64
use contact_26  contact_26_228
timestamp 1624494425
transform 1 0 9519 0 1 87
box 0 0 66 74
use contact_26  contact_26_230
timestamp 1624494425
transform 1 0 9387 0 1 87
box 0 0 66 74
use contact_25  contact_25_229
timestamp 1624494425
transform 1 0 9984 0 1 216
box 0 0 64 64
use contact_26  contact_26_229
timestamp 1624494425
transform 1 0 9983 0 1 211
box 0 0 66 74
use contact_23  contact_23_114
timestamp 1624494425
transform 1 0 9765 0 1 493
box 0 0 66 66
use contact_24  contact_24_114
timestamp 1624494425
transform 1 0 9769 0 1 493
box 0 0 58 66
use contact_25  contact_25_370
timestamp 1624494425
transform 1 0 9766 0 1 494
box 0 0 64 64
use contact_26  contact_26_370
timestamp 1624494425
transform 1 0 9765 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_114
timestamp 1624494425
transform -1 0 10110 0 1 868
box 65 0 675 1316
use contact_23  contact_23_113
timestamp 1624494425
transform 1 0 10389 0 1 617
box 0 0 66 66
use contact_24  contact_24_113
timestamp 1624494425
transform 1 0 10393 0 1 617
box 0 0 58 66
use contact_25  contact_25_227
timestamp 1624494425
transform 1 0 10172 0 1 216
box 0 0 64 64
use contact_25  contact_25_369
timestamp 1624494425
transform 1 0 10390 0 1 618
box 0 0 64 64
use contact_26  contact_26_227
timestamp 1624494425
transform 1 0 10171 0 1 211
box 0 0 66 74
use contact_26  contact_26_369
timestamp 1624494425
transform 1 0 10389 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_113
timestamp 1624494425
transform 1 0 10110 0 1 868
box 65 0 675 1316
use contact_23  contact_23_112
timestamp 1624494425
transform 1 0 11013 0 1 741
box 0 0 66 66
use contact_24  contact_24_112
timestamp 1624494425
transform 1 0 11017 0 1 741
box 0 0 58 66
use contact_25  contact_25_224
timestamp 1624494425
transform 1 0 10768 0 1 92
box 0 0 64 64
use contact_25  contact_25_226
timestamp 1624494425
transform 1 0 10636 0 1 92
box 0 0 64 64
use contact_25  contact_25_368
timestamp 1624494425
transform 1 0 11014 0 1 742
box 0 0 64 64
use contact_26  contact_26_224
timestamp 1624494425
transform 1 0 10767 0 1 87
box 0 0 66 74
use contact_26  contact_26_226
timestamp 1624494425
transform 1 0 10635 0 1 87
box 0 0 66 74
use contact_26  contact_26_368
timestamp 1624494425
transform 1 0 11013 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_112
timestamp 1624494425
transform -1 0 11358 0 1 868
box 65 0 675 1316
use contact_23  contact_23_111
timestamp 1624494425
transform 1 0 11637 0 1 369
box 0 0 66 66
use contact_24  contact_24_111
timestamp 1624494425
transform 1 0 11641 0 1 369
box 0 0 58 66
use contact_25  contact_25_223
timestamp 1624494425
transform 1 0 11420 0 1 216
box 0 0 64 64
use contact_25  contact_25_225
timestamp 1624494425
transform 1 0 11232 0 1 216
box 0 0 64 64
use contact_25  contact_25_367
timestamp 1624494425
transform 1 0 11638 0 1 370
box 0 0 64 64
use contact_26  contact_26_223
timestamp 1624494425
transform 1 0 11419 0 1 211
box 0 0 66 74
use contact_26  contact_26_225
timestamp 1624494425
transform 1 0 11231 0 1 211
box 0 0 66 74
use contact_26  contact_26_367
timestamp 1624494425
transform 1 0 11637 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_111
timestamp 1624494425
transform 1 0 11358 0 1 868
box 65 0 675 1316
use contact_23  contact_23_110
timestamp 1624494425
transform 1 0 12261 0 1 493
box 0 0 66 66
use contact_24  contact_24_110
timestamp 1624494425
transform 1 0 12265 0 1 493
box 0 0 58 66
use contact_25  contact_25_220
timestamp 1624494425
transform 1 0 12016 0 1 92
box 0 0 64 64
use contact_25  contact_25_222
timestamp 1624494425
transform 1 0 11884 0 1 92
box 0 0 64 64
use contact_25  contact_25_366
timestamp 1624494425
transform 1 0 12262 0 1 494
box 0 0 64 64
use contact_26  contact_26_220
timestamp 1624494425
transform 1 0 12015 0 1 87
box 0 0 66 74
use contact_26  contact_26_222
timestamp 1624494425
transform 1 0 11883 0 1 87
box 0 0 66 74
use contact_26  contact_26_366
timestamp 1624494425
transform 1 0 12261 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_110
timestamp 1624494425
transform -1 0 12606 0 1 868
box 65 0 675 1316
use contact_23  contact_23_109
timestamp 1624494425
transform 1 0 12885 0 1 617
box 0 0 66 66
use contact_24  contact_24_109
timestamp 1624494425
transform 1 0 12889 0 1 617
box 0 0 58 66
use contact_25  contact_25_219
timestamp 1624494425
transform 1 0 12668 0 1 216
box 0 0 64 64
use contact_25  contact_25_221
timestamp 1624494425
transform 1 0 12480 0 1 216
box 0 0 64 64
use contact_25  contact_25_365
timestamp 1624494425
transform 1 0 12886 0 1 618
box 0 0 64 64
use contact_26  contact_26_219
timestamp 1624494425
transform 1 0 12667 0 1 211
box 0 0 66 74
use contact_26  contact_26_221
timestamp 1624494425
transform 1 0 12479 0 1 211
box 0 0 66 74
use contact_26  contact_26_365
timestamp 1624494425
transform 1 0 12885 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_109
timestamp 1624494425
transform 1 0 12606 0 1 868
box 65 0 675 1316
use contact_23  contact_23_108
timestamp 1624494425
transform 1 0 13509 0 1 741
box 0 0 66 66
use contact_24  contact_24_108
timestamp 1624494425
transform 1 0 13513 0 1 741
box 0 0 58 66
use contact_25  contact_25_216
timestamp 1624494425
transform 1 0 13264 0 1 92
box 0 0 64 64
use contact_25  contact_25_218
timestamp 1624494425
transform 1 0 13132 0 1 92
box 0 0 64 64
use contact_25  contact_25_364
timestamp 1624494425
transform 1 0 13510 0 1 742
box 0 0 64 64
use contact_26  contact_26_216
timestamp 1624494425
transform 1 0 13263 0 1 87
box 0 0 66 74
use contact_26  contact_26_218
timestamp 1624494425
transform 1 0 13131 0 1 87
box 0 0 66 74
use contact_26  contact_26_364
timestamp 1624494425
transform 1 0 13509 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_108
timestamp 1624494425
transform -1 0 13854 0 1 868
box 65 0 675 1316
use contact_23  contact_23_107
timestamp 1624494425
transform 1 0 14133 0 1 369
box 0 0 66 66
use contact_24  contact_24_107
timestamp 1624494425
transform 1 0 14137 0 1 369
box 0 0 58 66
use contact_25  contact_25_215
timestamp 1624494425
transform 1 0 13916 0 1 216
box 0 0 64 64
use contact_25  contact_25_217
timestamp 1624494425
transform 1 0 13728 0 1 216
box 0 0 64 64
use contact_25  contact_25_363
timestamp 1624494425
transform 1 0 14134 0 1 370
box 0 0 64 64
use contact_26  contact_26_215
timestamp 1624494425
transform 1 0 13915 0 1 211
box 0 0 66 74
use contact_26  contact_26_217
timestamp 1624494425
transform 1 0 13727 0 1 211
box 0 0 66 74
use contact_26  contact_26_363
timestamp 1624494425
transform 1 0 14133 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_107
timestamp 1624494425
transform 1 0 13854 0 1 868
box 65 0 675 1316
use contact_23  contact_23_106
timestamp 1624494425
transform 1 0 14757 0 1 493
box 0 0 66 66
use contact_24  contact_24_106
timestamp 1624494425
transform 1 0 14761 0 1 493
box 0 0 58 66
use contact_25  contact_25_212
timestamp 1624494425
transform 1 0 14512 0 1 92
box 0 0 64 64
use contact_25  contact_25_214
timestamp 1624494425
transform 1 0 14380 0 1 92
box 0 0 64 64
use contact_25  contact_25_362
timestamp 1624494425
transform 1 0 14758 0 1 494
box 0 0 64 64
use contact_26  contact_26_212
timestamp 1624494425
transform 1 0 14511 0 1 87
box 0 0 66 74
use contact_26  contact_26_214
timestamp 1624494425
transform 1 0 14379 0 1 87
box 0 0 66 74
use contact_26  contact_26_362
timestamp 1624494425
transform 1 0 14757 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_106
timestamp 1624494425
transform -1 0 15102 0 1 868
box 65 0 675 1316
use contact_23  contact_23_105
timestamp 1624494425
transform 1 0 15381 0 1 617
box 0 0 66 66
use contact_24  contact_24_105
timestamp 1624494425
transform 1 0 15385 0 1 617
box 0 0 58 66
use contact_25  contact_25_211
timestamp 1624494425
transform 1 0 15164 0 1 216
box 0 0 64 64
use contact_25  contact_25_213
timestamp 1624494425
transform 1 0 14976 0 1 216
box 0 0 64 64
use contact_25  contact_25_361
timestamp 1624494425
transform 1 0 15382 0 1 618
box 0 0 64 64
use contact_26  contact_26_211
timestamp 1624494425
transform 1 0 15163 0 1 211
box 0 0 66 74
use contact_26  contact_26_213
timestamp 1624494425
transform 1 0 14975 0 1 211
box 0 0 66 74
use contact_26  contact_26_361
timestamp 1624494425
transform 1 0 15381 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_105
timestamp 1624494425
transform 1 0 15102 0 1 868
box 65 0 675 1316
use contact_23  contact_23_104
timestamp 1624494425
transform 1 0 16005 0 1 741
box 0 0 66 66
use contact_24  contact_24_104
timestamp 1624494425
transform 1 0 16009 0 1 741
box 0 0 58 66
use contact_25  contact_25_208
timestamp 1624494425
transform 1 0 15760 0 1 92
box 0 0 64 64
use contact_25  contact_25_210
timestamp 1624494425
transform 1 0 15628 0 1 92
box 0 0 64 64
use contact_25  contact_25_360
timestamp 1624494425
transform 1 0 16006 0 1 742
box 0 0 64 64
use contact_26  contact_26_208
timestamp 1624494425
transform 1 0 15759 0 1 87
box 0 0 66 74
use contact_26  contact_26_210
timestamp 1624494425
transform 1 0 15627 0 1 87
box 0 0 66 74
use contact_26  contact_26_360
timestamp 1624494425
transform 1 0 16005 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_104
timestamp 1624494425
transform -1 0 16350 0 1 868
box 65 0 675 1316
use contact_23  contact_23_103
timestamp 1624494425
transform 1 0 16629 0 1 369
box 0 0 66 66
use contact_24  contact_24_103
timestamp 1624494425
transform 1 0 16633 0 1 369
box 0 0 58 66
use contact_25  contact_25_207
timestamp 1624494425
transform 1 0 16412 0 1 216
box 0 0 64 64
use contact_25  contact_25_209
timestamp 1624494425
transform 1 0 16224 0 1 216
box 0 0 64 64
use contact_25  contact_25_359
timestamp 1624494425
transform 1 0 16630 0 1 370
box 0 0 64 64
use contact_26  contact_26_207
timestamp 1624494425
transform 1 0 16411 0 1 211
box 0 0 66 74
use contact_26  contact_26_209
timestamp 1624494425
transform 1 0 16223 0 1 211
box 0 0 66 74
use contact_26  contact_26_359
timestamp 1624494425
transform 1 0 16629 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_103
timestamp 1624494425
transform 1 0 16350 0 1 868
box 65 0 675 1316
use contact_23  contact_23_102
timestamp 1624494425
transform 1 0 17253 0 1 493
box 0 0 66 66
use contact_24  contact_24_102
timestamp 1624494425
transform 1 0 17257 0 1 493
box 0 0 58 66
use contact_25  contact_25_204
timestamp 1624494425
transform 1 0 17008 0 1 92
box 0 0 64 64
use contact_25  contact_25_206
timestamp 1624494425
transform 1 0 16876 0 1 92
box 0 0 64 64
use contact_25  contact_25_358
timestamp 1624494425
transform 1 0 17254 0 1 494
box 0 0 64 64
use contact_26  contact_26_204
timestamp 1624494425
transform 1 0 17007 0 1 87
box 0 0 66 74
use contact_26  contact_26_206
timestamp 1624494425
transform 1 0 16875 0 1 87
box 0 0 66 74
use contact_26  contact_26_358
timestamp 1624494425
transform 1 0 17253 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_102
timestamp 1624494425
transform -1 0 17598 0 1 868
box 65 0 675 1316
use contact_23  contact_23_101
timestamp 1624494425
transform 1 0 17877 0 1 617
box 0 0 66 66
use contact_24  contact_24_101
timestamp 1624494425
transform 1 0 17881 0 1 617
box 0 0 58 66
use contact_25  contact_25_203
timestamp 1624494425
transform 1 0 17660 0 1 216
box 0 0 64 64
use contact_25  contact_25_205
timestamp 1624494425
transform 1 0 17472 0 1 216
box 0 0 64 64
use contact_25  contact_25_357
timestamp 1624494425
transform 1 0 17878 0 1 618
box 0 0 64 64
use contact_26  contact_26_203
timestamp 1624494425
transform 1 0 17659 0 1 211
box 0 0 66 74
use contact_26  contact_26_205
timestamp 1624494425
transform 1 0 17471 0 1 211
box 0 0 66 74
use contact_26  contact_26_357
timestamp 1624494425
transform 1 0 17877 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_101
timestamp 1624494425
transform 1 0 17598 0 1 868
box 65 0 675 1316
use contact_23  contact_23_100
timestamp 1624494425
transform 1 0 18501 0 1 741
box 0 0 66 66
use contact_24  contact_24_100
timestamp 1624494425
transform 1 0 18505 0 1 741
box 0 0 58 66
use contact_25  contact_25_200
timestamp 1624494425
transform 1 0 18256 0 1 92
box 0 0 64 64
use contact_25  contact_25_202
timestamp 1624494425
transform 1 0 18124 0 1 92
box 0 0 64 64
use contact_25  contact_25_356
timestamp 1624494425
transform 1 0 18502 0 1 742
box 0 0 64 64
use contact_26  contact_26_200
timestamp 1624494425
transform 1 0 18255 0 1 87
box 0 0 66 74
use contact_26  contact_26_202
timestamp 1624494425
transform 1 0 18123 0 1 87
box 0 0 66 74
use contact_26  contact_26_356
timestamp 1624494425
transform 1 0 18501 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_100
timestamp 1624494425
transform -1 0 18846 0 1 868
box 65 0 675 1316
use contact_23  contact_23_99
timestamp 1624494425
transform 1 0 19125 0 1 369
box 0 0 66 66
use contact_24  contact_24_99
timestamp 1624494425
transform 1 0 19129 0 1 369
box 0 0 58 66
use contact_25  contact_25_199
timestamp 1624494425
transform 1 0 18908 0 1 216
box 0 0 64 64
use contact_25  contact_25_201
timestamp 1624494425
transform 1 0 18720 0 1 216
box 0 0 64 64
use contact_25  contact_25_355
timestamp 1624494425
transform 1 0 19126 0 1 370
box 0 0 64 64
use contact_26  contact_26_199
timestamp 1624494425
transform 1 0 18907 0 1 211
box 0 0 66 74
use contact_26  contact_26_201
timestamp 1624494425
transform 1 0 18719 0 1 211
box 0 0 66 74
use contact_26  contact_26_355
timestamp 1624494425
transform 1 0 19125 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_99
timestamp 1624494425
transform 1 0 18846 0 1 868
box 65 0 675 1316
use contact_23  contact_23_98
timestamp 1624494425
transform 1 0 19749 0 1 493
box 0 0 66 66
use contact_24  contact_24_98
timestamp 1624494425
transform 1 0 19753 0 1 493
box 0 0 58 66
use contact_25  contact_25_196
timestamp 1624494425
transform 1 0 19504 0 1 92
box 0 0 64 64
use contact_25  contact_25_198
timestamp 1624494425
transform 1 0 19372 0 1 92
box 0 0 64 64
use contact_25  contact_25_354
timestamp 1624494425
transform 1 0 19750 0 1 494
box 0 0 64 64
use contact_26  contact_26_196
timestamp 1624494425
transform 1 0 19503 0 1 87
box 0 0 66 74
use contact_26  contact_26_198
timestamp 1624494425
transform 1 0 19371 0 1 87
box 0 0 66 74
use contact_26  contact_26_354
timestamp 1624494425
transform 1 0 19749 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_98
timestamp 1624494425
transform -1 0 20094 0 1 868
box 65 0 675 1316
use contact_23  contact_23_97
timestamp 1624494425
transform 1 0 20373 0 1 617
box 0 0 66 66
use contact_25  contact_25_195
timestamp 1624494425
transform 1 0 20156 0 1 216
box 0 0 64 64
use contact_25  contact_25_197
timestamp 1624494425
transform 1 0 19968 0 1 216
box 0 0 64 64
use contact_25  contact_25_353
timestamp 1624494425
transform 1 0 20374 0 1 618
box 0 0 64 64
use contact_26  contact_26_195
timestamp 1624494425
transform 1 0 20155 0 1 211
box 0 0 66 74
use contact_26  contact_26_197
timestamp 1624494425
transform 1 0 19967 0 1 211
box 0 0 66 74
use contact_26  contact_26_353
timestamp 1624494425
transform 1 0 20373 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_97
timestamp 1624494425
transform 1 0 20094 0 1 868
box 65 0 675 1316
use contact_24  contact_24_97
timestamp 1624494425
transform 1 0 20377 0 1 617
box 0 0 58 66
use contact_25  contact_25_192
timestamp 1624494425
transform 1 0 20752 0 1 92
box 0 0 64 64
use contact_25  contact_25_194
timestamp 1624494425
transform 1 0 20620 0 1 92
box 0 0 64 64
use contact_26  contact_26_192
timestamp 1624494425
transform 1 0 20751 0 1 87
box 0 0 66 74
use contact_26  contact_26_194
timestamp 1624494425
transform 1 0 20619 0 1 87
box 0 0 66 74
use column_mux_0  column_mux_0_96
timestamp 1624494425
transform -1 0 21342 0 1 868
box 65 0 675 1316
use contact_23  contact_23_96
timestamp 1624494425
transform 1 0 20997 0 1 741
box 0 0 66 66
use contact_24  contact_24_96
timestamp 1624494425
transform 1 0 21001 0 1 741
box 0 0 58 66
use contact_25  contact_25_191
timestamp 1624494425
transform 1 0 21404 0 1 216
box 0 0 64 64
use contact_25  contact_25_193
timestamp 1624494425
transform 1 0 21216 0 1 216
box 0 0 64 64
use contact_25  contact_25_352
timestamp 1624494425
transform 1 0 20998 0 1 742
box 0 0 64 64
use contact_26  contact_26_191
timestamp 1624494425
transform 1 0 21403 0 1 211
box 0 0 66 74
use contact_26  contact_26_193
timestamp 1624494425
transform 1 0 21215 0 1 211
box 0 0 66 74
use contact_26  contact_26_352
timestamp 1624494425
transform 1 0 20997 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_95
timestamp 1624494425
transform 1 0 21342 0 1 868
box 65 0 675 1316
use contact_23  contact_23_95
timestamp 1624494425
transform 1 0 21621 0 1 369
box 0 0 66 66
use contact_24  contact_24_95
timestamp 1624494425
transform 1 0 21625 0 1 369
box 0 0 58 66
use contact_25  contact_25_188
timestamp 1624494425
transform 1 0 22000 0 1 92
box 0 0 64 64
use contact_25  contact_25_190
timestamp 1624494425
transform 1 0 21868 0 1 92
box 0 0 64 64
use contact_25  contact_25_351
timestamp 1624494425
transform 1 0 21622 0 1 370
box 0 0 64 64
use contact_26  contact_26_188
timestamp 1624494425
transform 1 0 21999 0 1 87
box 0 0 66 74
use contact_26  contact_26_190
timestamp 1624494425
transform 1 0 21867 0 1 87
box 0 0 66 74
use contact_26  contact_26_351
timestamp 1624494425
transform 1 0 21621 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_94
timestamp 1624494425
transform -1 0 22590 0 1 868
box 65 0 675 1316
use contact_23  contact_23_94
timestamp 1624494425
transform 1 0 22245 0 1 493
box 0 0 66 66
use contact_24  contact_24_94
timestamp 1624494425
transform 1 0 22249 0 1 493
box 0 0 58 66
use contact_25  contact_25_187
timestamp 1624494425
transform 1 0 22652 0 1 216
box 0 0 64 64
use contact_25  contact_25_189
timestamp 1624494425
transform 1 0 22464 0 1 216
box 0 0 64 64
use contact_25  contact_25_350
timestamp 1624494425
transform 1 0 22246 0 1 494
box 0 0 64 64
use contact_26  contact_26_187
timestamp 1624494425
transform 1 0 22651 0 1 211
box 0 0 66 74
use contact_26  contact_26_189
timestamp 1624494425
transform 1 0 22463 0 1 211
box 0 0 66 74
use contact_26  contact_26_350
timestamp 1624494425
transform 1 0 22245 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_93
timestamp 1624494425
transform 1 0 22590 0 1 868
box 65 0 675 1316
use contact_23  contact_23_93
timestamp 1624494425
transform 1 0 22869 0 1 617
box 0 0 66 66
use contact_24  contact_24_93
timestamp 1624494425
transform 1 0 22873 0 1 617
box 0 0 58 66
use contact_25  contact_25_184
timestamp 1624494425
transform 1 0 23248 0 1 92
box 0 0 64 64
use contact_25  contact_25_186
timestamp 1624494425
transform 1 0 23116 0 1 92
box 0 0 64 64
use contact_25  contact_25_349
timestamp 1624494425
transform 1 0 22870 0 1 618
box 0 0 64 64
use contact_26  contact_26_184
timestamp 1624494425
transform 1 0 23247 0 1 87
box 0 0 66 74
use contact_26  contact_26_186
timestamp 1624494425
transform 1 0 23115 0 1 87
box 0 0 66 74
use contact_26  contact_26_349
timestamp 1624494425
transform 1 0 22869 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_92
timestamp 1624494425
transform -1 0 23838 0 1 868
box 65 0 675 1316
use contact_23  contact_23_92
timestamp 1624494425
transform 1 0 23493 0 1 741
box 0 0 66 66
use contact_24  contact_24_92
timestamp 1624494425
transform 1 0 23497 0 1 741
box 0 0 58 66
use contact_25  contact_25_183
timestamp 1624494425
transform 1 0 23900 0 1 216
box 0 0 64 64
use contact_25  contact_25_185
timestamp 1624494425
transform 1 0 23712 0 1 216
box 0 0 64 64
use contact_25  contact_25_348
timestamp 1624494425
transform 1 0 23494 0 1 742
box 0 0 64 64
use contact_26  contact_26_183
timestamp 1624494425
transform 1 0 23899 0 1 211
box 0 0 66 74
use contact_26  contact_26_185
timestamp 1624494425
transform 1 0 23711 0 1 211
box 0 0 66 74
use contact_26  contact_26_348
timestamp 1624494425
transform 1 0 23493 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_91
timestamp 1624494425
transform 1 0 23838 0 1 868
box 65 0 675 1316
use contact_23  contact_23_91
timestamp 1624494425
transform 1 0 24117 0 1 369
box 0 0 66 66
use contact_24  contact_24_91
timestamp 1624494425
transform 1 0 24121 0 1 369
box 0 0 58 66
use contact_25  contact_25_180
timestamp 1624494425
transform 1 0 24496 0 1 92
box 0 0 64 64
use contact_25  contact_25_182
timestamp 1624494425
transform 1 0 24364 0 1 92
box 0 0 64 64
use contact_25  contact_25_347
timestamp 1624494425
transform 1 0 24118 0 1 370
box 0 0 64 64
use contact_26  contact_26_180
timestamp 1624494425
transform 1 0 24495 0 1 87
box 0 0 66 74
use contact_26  contact_26_182
timestamp 1624494425
transform 1 0 24363 0 1 87
box 0 0 66 74
use contact_26  contact_26_347
timestamp 1624494425
transform 1 0 24117 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_90
timestamp 1624494425
transform -1 0 25086 0 1 868
box 65 0 675 1316
use contact_23  contact_23_90
timestamp 1624494425
transform 1 0 24741 0 1 493
box 0 0 66 66
use contact_24  contact_24_90
timestamp 1624494425
transform 1 0 24745 0 1 493
box 0 0 58 66
use contact_25  contact_25_179
timestamp 1624494425
transform 1 0 25148 0 1 216
box 0 0 64 64
use contact_25  contact_25_181
timestamp 1624494425
transform 1 0 24960 0 1 216
box 0 0 64 64
use contact_25  contact_25_346
timestamp 1624494425
transform 1 0 24742 0 1 494
box 0 0 64 64
use contact_26  contact_26_179
timestamp 1624494425
transform 1 0 25147 0 1 211
box 0 0 66 74
use contact_26  contact_26_181
timestamp 1624494425
transform 1 0 24959 0 1 211
box 0 0 66 74
use contact_26  contact_26_346
timestamp 1624494425
transform 1 0 24741 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_89
timestamp 1624494425
transform 1 0 25086 0 1 868
box 65 0 675 1316
use contact_23  contact_23_89
timestamp 1624494425
transform 1 0 25365 0 1 617
box 0 0 66 66
use contact_24  contact_24_89
timestamp 1624494425
transform 1 0 25369 0 1 617
box 0 0 58 66
use contact_25  contact_25_176
timestamp 1624494425
transform 1 0 25744 0 1 92
box 0 0 64 64
use contact_25  contact_25_178
timestamp 1624494425
transform 1 0 25612 0 1 92
box 0 0 64 64
use contact_25  contact_25_345
timestamp 1624494425
transform 1 0 25366 0 1 618
box 0 0 64 64
use contact_26  contact_26_176
timestamp 1624494425
transform 1 0 25743 0 1 87
box 0 0 66 74
use contact_26  contact_26_178
timestamp 1624494425
transform 1 0 25611 0 1 87
box 0 0 66 74
use contact_26  contact_26_345
timestamp 1624494425
transform 1 0 25365 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_88
timestamp 1624494425
transform -1 0 26334 0 1 868
box 65 0 675 1316
use contact_23  contact_23_88
timestamp 1624494425
transform 1 0 25989 0 1 741
box 0 0 66 66
use contact_24  contact_24_88
timestamp 1624494425
transform 1 0 25993 0 1 741
box 0 0 58 66
use contact_25  contact_25_175
timestamp 1624494425
transform 1 0 26396 0 1 216
box 0 0 64 64
use contact_25  contact_25_177
timestamp 1624494425
transform 1 0 26208 0 1 216
box 0 0 64 64
use contact_25  contact_25_344
timestamp 1624494425
transform 1 0 25990 0 1 742
box 0 0 64 64
use contact_26  contact_26_175
timestamp 1624494425
transform 1 0 26395 0 1 211
box 0 0 66 74
use contact_26  contact_26_177
timestamp 1624494425
transform 1 0 26207 0 1 211
box 0 0 66 74
use contact_26  contact_26_344
timestamp 1624494425
transform 1 0 25989 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_87
timestamp 1624494425
transform 1 0 26334 0 1 868
box 65 0 675 1316
use contact_23  contact_23_87
timestamp 1624494425
transform 1 0 26613 0 1 369
box 0 0 66 66
use contact_24  contact_24_87
timestamp 1624494425
transform 1 0 26617 0 1 369
box 0 0 58 66
use contact_25  contact_25_172
timestamp 1624494425
transform 1 0 26992 0 1 92
box 0 0 64 64
use contact_25  contact_25_174
timestamp 1624494425
transform 1 0 26860 0 1 92
box 0 0 64 64
use contact_25  contact_25_343
timestamp 1624494425
transform 1 0 26614 0 1 370
box 0 0 64 64
use contact_26  contact_26_172
timestamp 1624494425
transform 1 0 26991 0 1 87
box 0 0 66 74
use contact_26  contact_26_174
timestamp 1624494425
transform 1 0 26859 0 1 87
box 0 0 66 74
use contact_26  contact_26_343
timestamp 1624494425
transform 1 0 26613 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_86
timestamp 1624494425
transform -1 0 27582 0 1 868
box 65 0 675 1316
use contact_23  contact_23_86
timestamp 1624494425
transform 1 0 27237 0 1 493
box 0 0 66 66
use contact_24  contact_24_86
timestamp 1624494425
transform 1 0 27241 0 1 493
box 0 0 58 66
use contact_25  contact_25_171
timestamp 1624494425
transform 1 0 27644 0 1 216
box 0 0 64 64
use contact_25  contact_25_173
timestamp 1624494425
transform 1 0 27456 0 1 216
box 0 0 64 64
use contact_25  contact_25_342
timestamp 1624494425
transform 1 0 27238 0 1 494
box 0 0 64 64
use contact_26  contact_26_171
timestamp 1624494425
transform 1 0 27643 0 1 211
box 0 0 66 74
use contact_26  contact_26_173
timestamp 1624494425
transform 1 0 27455 0 1 211
box 0 0 66 74
use contact_26  contact_26_342
timestamp 1624494425
transform 1 0 27237 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_85
timestamp 1624494425
transform 1 0 27582 0 1 868
box 65 0 675 1316
use contact_23  contact_23_85
timestamp 1624494425
transform 1 0 27861 0 1 617
box 0 0 66 66
use contact_24  contact_24_85
timestamp 1624494425
transform 1 0 27865 0 1 617
box 0 0 58 66
use contact_25  contact_25_168
timestamp 1624494425
transform 1 0 28240 0 1 92
box 0 0 64 64
use contact_25  contact_25_170
timestamp 1624494425
transform 1 0 28108 0 1 92
box 0 0 64 64
use contact_25  contact_25_341
timestamp 1624494425
transform 1 0 27862 0 1 618
box 0 0 64 64
use contact_26  contact_26_168
timestamp 1624494425
transform 1 0 28239 0 1 87
box 0 0 66 74
use contact_26  contact_26_170
timestamp 1624494425
transform 1 0 28107 0 1 87
box 0 0 66 74
use contact_26  contact_26_341
timestamp 1624494425
transform 1 0 27861 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_84
timestamp 1624494425
transform -1 0 28830 0 1 868
box 65 0 675 1316
use contact_23  contact_23_84
timestamp 1624494425
transform 1 0 28485 0 1 741
box 0 0 66 66
use contact_24  contact_24_84
timestamp 1624494425
transform 1 0 28489 0 1 741
box 0 0 58 66
use contact_25  contact_25_167
timestamp 1624494425
transform 1 0 28892 0 1 216
box 0 0 64 64
use contact_25  contact_25_169
timestamp 1624494425
transform 1 0 28704 0 1 216
box 0 0 64 64
use contact_25  contact_25_340
timestamp 1624494425
transform 1 0 28486 0 1 742
box 0 0 64 64
use contact_26  contact_26_167
timestamp 1624494425
transform 1 0 28891 0 1 211
box 0 0 66 74
use contact_26  contact_26_169
timestamp 1624494425
transform 1 0 28703 0 1 211
box 0 0 66 74
use contact_26  contact_26_340
timestamp 1624494425
transform 1 0 28485 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_83
timestamp 1624494425
transform 1 0 28830 0 1 868
box 65 0 675 1316
use contact_23  contact_23_83
timestamp 1624494425
transform 1 0 29109 0 1 369
box 0 0 66 66
use contact_24  contact_24_83
timestamp 1624494425
transform 1 0 29113 0 1 369
box 0 0 58 66
use contact_25  contact_25_164
timestamp 1624494425
transform 1 0 29488 0 1 92
box 0 0 64 64
use contact_25  contact_25_166
timestamp 1624494425
transform 1 0 29356 0 1 92
box 0 0 64 64
use contact_25  contact_25_339
timestamp 1624494425
transform 1 0 29110 0 1 370
box 0 0 64 64
use contact_26  contact_26_164
timestamp 1624494425
transform 1 0 29487 0 1 87
box 0 0 66 74
use contact_26  contact_26_166
timestamp 1624494425
transform 1 0 29355 0 1 87
box 0 0 66 74
use contact_26  contact_26_339
timestamp 1624494425
transform 1 0 29109 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_82
timestamp 1624494425
transform -1 0 30078 0 1 868
box 65 0 675 1316
use contact_23  contact_23_82
timestamp 1624494425
transform 1 0 29733 0 1 493
box 0 0 66 66
use contact_24  contact_24_82
timestamp 1624494425
transform 1 0 29737 0 1 493
box 0 0 58 66
use contact_25  contact_25_163
timestamp 1624494425
transform 1 0 30140 0 1 216
box 0 0 64 64
use contact_25  contact_25_165
timestamp 1624494425
transform 1 0 29952 0 1 216
box 0 0 64 64
use contact_25  contact_25_338
timestamp 1624494425
transform 1 0 29734 0 1 494
box 0 0 64 64
use contact_26  contact_26_163
timestamp 1624494425
transform 1 0 30139 0 1 211
box 0 0 66 74
use contact_26  contact_26_165
timestamp 1624494425
transform 1 0 29951 0 1 211
box 0 0 66 74
use contact_26  contact_26_338
timestamp 1624494425
transform 1 0 29733 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_81
timestamp 1624494425
transform 1 0 30078 0 1 868
box 65 0 675 1316
use contact_23  contact_23_81
timestamp 1624494425
transform 1 0 30357 0 1 617
box 0 0 66 66
use contact_24  contact_24_81
timestamp 1624494425
transform 1 0 30361 0 1 617
box 0 0 58 66
use contact_25  contact_25_160
timestamp 1624494425
transform 1 0 30736 0 1 92
box 0 0 64 64
use contact_25  contact_25_162
timestamp 1624494425
transform 1 0 30604 0 1 92
box 0 0 64 64
use contact_25  contact_25_337
timestamp 1624494425
transform 1 0 30358 0 1 618
box 0 0 64 64
use contact_26  contact_26_160
timestamp 1624494425
transform 1 0 30735 0 1 87
box 0 0 66 74
use contact_26  contact_26_162
timestamp 1624494425
transform 1 0 30603 0 1 87
box 0 0 66 74
use contact_26  contact_26_337
timestamp 1624494425
transform 1 0 30357 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_80
timestamp 1624494425
transform -1 0 31326 0 1 868
box 65 0 675 1316
use contact_23  contact_23_80
timestamp 1624494425
transform 1 0 30981 0 1 741
box 0 0 66 66
use contact_24  contact_24_80
timestamp 1624494425
transform 1 0 30985 0 1 741
box 0 0 58 66
use contact_25  contact_25_161
timestamp 1624494425
transform 1 0 31200 0 1 216
box 0 0 64 64
use contact_25  contact_25_336
timestamp 1624494425
transform 1 0 30982 0 1 742
box 0 0 64 64
use contact_26  contact_26_161
timestamp 1624494425
transform 1 0 31199 0 1 211
box 0 0 66 74
use contact_26  contact_26_336
timestamp 1624494425
transform 1 0 30981 0 1 737
box 0 0 66 74
use contact_25  contact_25_159
timestamp 1624494425
transform 1 0 31388 0 1 216
box 0 0 64 64
use contact_26  contact_26_159
timestamp 1624494425
transform 1 0 31387 0 1 211
box 0 0 66 74
use contact_25  contact_25_158
timestamp 1624494425
transform 1 0 31852 0 1 92
box 0 0 64 64
use contact_26  contact_26_158
timestamp 1624494425
transform 1 0 31851 0 1 87
box 0 0 66 74
use contact_25  contact_25_156
timestamp 1624494425
transform 1 0 31984 0 1 92
box 0 0 64 64
use contact_26  contact_26_156
timestamp 1624494425
transform 1 0 31983 0 1 87
box 0 0 66 74
use contact_23  contact_23_79
timestamp 1624494425
transform 1 0 31605 0 1 369
box 0 0 66 66
use contact_24  contact_24_79
timestamp 1624494425
transform 1 0 31609 0 1 369
box 0 0 58 66
use contact_25  contact_25_335
timestamp 1624494425
transform 1 0 31606 0 1 370
box 0 0 64 64
use contact_26  contact_26_335
timestamp 1624494425
transform 1 0 31605 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_79
timestamp 1624494425
transform 1 0 31326 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_78
timestamp 1624494425
transform -1 0 32574 0 1 868
box 65 0 675 1316
use contact_23  contact_23_78
timestamp 1624494425
transform 1 0 32229 0 1 493
box 0 0 66 66
use contact_24  contact_24_78
timestamp 1624494425
transform 1 0 32233 0 1 493
box 0 0 58 66
use contact_25  contact_25_157
timestamp 1624494425
transform 1 0 32448 0 1 216
box 0 0 64 64
use contact_25  contact_25_334
timestamp 1624494425
transform 1 0 32230 0 1 494
box 0 0 64 64
use contact_26  contact_26_157
timestamp 1624494425
transform 1 0 32447 0 1 211
box 0 0 66 74
use contact_26  contact_26_334
timestamp 1624494425
transform 1 0 32229 0 1 489
box 0 0 66 74
use contact_26  contact_26_333
timestamp 1624494425
transform 1 0 32853 0 1 613
box 0 0 66 74
use contact_26  contact_26_155
timestamp 1624494425
transform 1 0 32635 0 1 211
box 0 0 66 74
use contact_26  contact_26_154
timestamp 1624494425
transform 1 0 33099 0 1 87
box 0 0 66 74
use contact_25  contact_25_333
timestamp 1624494425
transform 1 0 32854 0 1 618
box 0 0 64 64
use contact_25  contact_25_155
timestamp 1624494425
transform 1 0 32636 0 1 216
box 0 0 64 64
use contact_25  contact_25_154
timestamp 1624494425
transform 1 0 33100 0 1 92
box 0 0 64 64
use contact_24  contact_24_77
timestamp 1624494425
transform 1 0 32857 0 1 617
box 0 0 58 66
use contact_23  contact_23_77
timestamp 1624494425
transform 1 0 32853 0 1 617
box 0 0 66 66
use column_mux_0  column_mux_0_77
timestamp 1624494425
transform 1 0 32574 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_76
timestamp 1624494425
transform -1 0 33822 0 1 868
box 65 0 675 1316
use contact_23  contact_23_76
timestamp 1624494425
transform 1 0 33477 0 1 741
box 0 0 66 66
use contact_24  contact_24_76
timestamp 1624494425
transform 1 0 33481 0 1 741
box 0 0 58 66
use contact_25  contact_25_152
timestamp 1624494425
transform 1 0 33232 0 1 92
box 0 0 64 64
use contact_25  contact_25_153
timestamp 1624494425
transform 1 0 33696 0 1 216
box 0 0 64 64
use contact_25  contact_25_332
timestamp 1624494425
transform 1 0 33478 0 1 742
box 0 0 64 64
use contact_26  contact_26_152
timestamp 1624494425
transform 1 0 33231 0 1 87
box 0 0 66 74
use contact_26  contact_26_153
timestamp 1624494425
transform 1 0 33695 0 1 211
box 0 0 66 74
use contact_26  contact_26_332
timestamp 1624494425
transform 1 0 33477 0 1 737
box 0 0 66 74
use contact_26  contact_26_331
timestamp 1624494425
transform 1 0 34101 0 1 365
box 0 0 66 74
use contact_26  contact_26_151
timestamp 1624494425
transform 1 0 33883 0 1 211
box 0 0 66 74
use contact_26  contact_26_150
timestamp 1624494425
transform 1 0 34347 0 1 87
box 0 0 66 74
use contact_25  contact_25_331
timestamp 1624494425
transform 1 0 34102 0 1 370
box 0 0 64 64
use contact_25  contact_25_151
timestamp 1624494425
transform 1 0 33884 0 1 216
box 0 0 64 64
use contact_25  contact_25_150
timestamp 1624494425
transform 1 0 34348 0 1 92
box 0 0 64 64
use contact_24  contact_24_75
timestamp 1624494425
transform 1 0 34105 0 1 369
box 0 0 58 66
use contact_23  contact_23_75
timestamp 1624494425
transform 1 0 34101 0 1 369
box 0 0 66 66
use column_mux_0  column_mux_0_75
timestamp 1624494425
transform 1 0 33822 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_74
timestamp 1624494425
transform -1 0 35070 0 1 868
box 65 0 675 1316
use contact_23  contact_23_74
timestamp 1624494425
transform 1 0 34725 0 1 493
box 0 0 66 66
use contact_24  contact_24_74
timestamp 1624494425
transform 1 0 34729 0 1 493
box 0 0 58 66
use contact_25  contact_25_148
timestamp 1624494425
transform 1 0 34480 0 1 92
box 0 0 64 64
use contact_25  contact_25_149
timestamp 1624494425
transform 1 0 34944 0 1 216
box 0 0 64 64
use contact_25  contact_25_330
timestamp 1624494425
transform 1 0 34726 0 1 494
box 0 0 64 64
use contact_26  contact_26_148
timestamp 1624494425
transform 1 0 34479 0 1 87
box 0 0 66 74
use contact_26  contact_26_149
timestamp 1624494425
transform 1 0 34943 0 1 211
box 0 0 66 74
use contact_26  contact_26_330
timestamp 1624494425
transform 1 0 34725 0 1 489
box 0 0 66 74
use contact_26  contact_26_329
timestamp 1624494425
transform 1 0 35349 0 1 613
box 0 0 66 74
use contact_26  contact_26_147
timestamp 1624494425
transform 1 0 35131 0 1 211
box 0 0 66 74
use contact_26  contact_26_146
timestamp 1624494425
transform 1 0 35595 0 1 87
box 0 0 66 74
use contact_25  contact_25_329
timestamp 1624494425
transform 1 0 35350 0 1 618
box 0 0 64 64
use contact_25  contact_25_147
timestamp 1624494425
transform 1 0 35132 0 1 216
box 0 0 64 64
use contact_25  contact_25_146
timestamp 1624494425
transform 1 0 35596 0 1 92
box 0 0 64 64
use contact_24  contact_24_73
timestamp 1624494425
transform 1 0 35353 0 1 617
box 0 0 58 66
use contact_23  contact_23_73
timestamp 1624494425
transform 1 0 35349 0 1 617
box 0 0 66 66
use column_mux_0  column_mux_0_73
timestamp 1624494425
transform 1 0 35070 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_72
timestamp 1624494425
transform -1 0 36318 0 1 868
box 65 0 675 1316
use contact_23  contact_23_72
timestamp 1624494425
transform 1 0 35973 0 1 741
box 0 0 66 66
use contact_24  contact_24_72
timestamp 1624494425
transform 1 0 35977 0 1 741
box 0 0 58 66
use contact_25  contact_25_144
timestamp 1624494425
transform 1 0 35728 0 1 92
box 0 0 64 64
use contact_25  contact_25_145
timestamp 1624494425
transform 1 0 36192 0 1 216
box 0 0 64 64
use contact_25  contact_25_328
timestamp 1624494425
transform 1 0 35974 0 1 742
box 0 0 64 64
use contact_26  contact_26_144
timestamp 1624494425
transform 1 0 35727 0 1 87
box 0 0 66 74
use contact_26  contact_26_145
timestamp 1624494425
transform 1 0 36191 0 1 211
box 0 0 66 74
use contact_26  contact_26_328
timestamp 1624494425
transform 1 0 35973 0 1 737
box 0 0 66 74
use contact_23  contact_23_71
timestamp 1624494425
transform 1 0 36597 0 1 369
box 0 0 66 66
use contact_24  contact_24_71
timestamp 1624494425
transform 1 0 36601 0 1 369
box 0 0 58 66
use contact_25  contact_25_142
timestamp 1624494425
transform 1 0 36844 0 1 92
box 0 0 64 64
use contact_25  contact_25_143
timestamp 1624494425
transform 1 0 36380 0 1 216
box 0 0 64 64
use contact_25  contact_25_327
timestamp 1624494425
transform 1 0 36598 0 1 370
box 0 0 64 64
use contact_26  contact_26_142
timestamp 1624494425
transform 1 0 36843 0 1 87
box 0 0 66 74
use contact_26  contact_26_143
timestamp 1624494425
transform 1 0 36379 0 1 211
box 0 0 66 74
use contact_26  contact_26_327
timestamp 1624494425
transform 1 0 36597 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_71
timestamp 1624494425
transform 1 0 36318 0 1 868
box 65 0 675 1316
use contact_23  contact_23_70
timestamp 1624494425
transform 1 0 37221 0 1 493
box 0 0 66 66
use contact_24  contact_24_70
timestamp 1624494425
transform 1 0 37225 0 1 493
box 0 0 58 66
use contact_25  contact_25_140
timestamp 1624494425
transform 1 0 36976 0 1 92
box 0 0 64 64
use contact_25  contact_25_141
timestamp 1624494425
transform 1 0 37440 0 1 216
box 0 0 64 64
use contact_25  contact_25_326
timestamp 1624494425
transform 1 0 37222 0 1 494
box 0 0 64 64
use contact_26  contact_26_140
timestamp 1624494425
transform 1 0 36975 0 1 87
box 0 0 66 74
use contact_26  contact_26_141
timestamp 1624494425
transform 1 0 37439 0 1 211
box 0 0 66 74
use contact_26  contact_26_326
timestamp 1624494425
transform 1 0 37221 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_70
timestamp 1624494425
transform -1 0 37566 0 1 868
box 65 0 675 1316
use contact_23  contact_23_69
timestamp 1624494425
transform 1 0 37845 0 1 617
box 0 0 66 66
use contact_24  contact_24_69
timestamp 1624494425
transform 1 0 37849 0 1 617
box 0 0 58 66
use contact_25  contact_25_138
timestamp 1624494425
transform 1 0 38092 0 1 92
box 0 0 64 64
use contact_25  contact_25_139
timestamp 1624494425
transform 1 0 37628 0 1 216
box 0 0 64 64
use contact_25  contact_25_325
timestamp 1624494425
transform 1 0 37846 0 1 618
box 0 0 64 64
use contact_26  contact_26_138
timestamp 1624494425
transform 1 0 38091 0 1 87
box 0 0 66 74
use contact_26  contact_26_139
timestamp 1624494425
transform 1 0 37627 0 1 211
box 0 0 66 74
use contact_26  contact_26_325
timestamp 1624494425
transform 1 0 37845 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_69
timestamp 1624494425
transform 1 0 37566 0 1 868
box 65 0 675 1316
use contact_23  contact_23_68
timestamp 1624494425
transform 1 0 38469 0 1 741
box 0 0 66 66
use contact_24  contact_24_68
timestamp 1624494425
transform 1 0 38473 0 1 741
box 0 0 58 66
use contact_25  contact_25_136
timestamp 1624494425
transform 1 0 38224 0 1 92
box 0 0 64 64
use contact_25  contact_25_137
timestamp 1624494425
transform 1 0 38688 0 1 216
box 0 0 64 64
use contact_25  contact_25_324
timestamp 1624494425
transform 1 0 38470 0 1 742
box 0 0 64 64
use contact_26  contact_26_136
timestamp 1624494425
transform 1 0 38223 0 1 87
box 0 0 66 74
use contact_26  contact_26_137
timestamp 1624494425
transform 1 0 38687 0 1 211
box 0 0 66 74
use contact_26  contact_26_324
timestamp 1624494425
transform 1 0 38469 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_68
timestamp 1624494425
transform -1 0 38814 0 1 868
box 65 0 675 1316
use contact_23  contact_23_67
timestamp 1624494425
transform 1 0 39093 0 1 369
box 0 0 66 66
use contact_24  contact_24_67
timestamp 1624494425
transform 1 0 39097 0 1 369
box 0 0 58 66
use contact_25  contact_25_135
timestamp 1624494425
transform 1 0 38876 0 1 216
box 0 0 64 64
use contact_25  contact_25_323
timestamp 1624494425
transform 1 0 39094 0 1 370
box 0 0 64 64
use contact_26  contact_26_135
timestamp 1624494425
transform 1 0 38875 0 1 211
box 0 0 66 74
use contact_26  contact_26_323
timestamp 1624494425
transform 1 0 39093 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_67
timestamp 1624494425
transform 1 0 38814 0 1 868
box 65 0 675 1316
use contact_23  contact_23_66
timestamp 1624494425
transform 1 0 39717 0 1 493
box 0 0 66 66
use contact_24  contact_24_66
timestamp 1624494425
transform 1 0 39721 0 1 493
box 0 0 58 66
use contact_25  contact_25_132
timestamp 1624494425
transform 1 0 39472 0 1 92
box 0 0 64 64
use contact_25  contact_25_134
timestamp 1624494425
transform 1 0 39340 0 1 92
box 0 0 64 64
use contact_25  contact_25_322
timestamp 1624494425
transform 1 0 39718 0 1 494
box 0 0 64 64
use contact_26  contact_26_132
timestamp 1624494425
transform 1 0 39471 0 1 87
box 0 0 66 74
use contact_26  contact_26_134
timestamp 1624494425
transform 1 0 39339 0 1 87
box 0 0 66 74
use contact_26  contact_26_322
timestamp 1624494425
transform 1 0 39717 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_66
timestamp 1624494425
transform -1 0 40062 0 1 868
box 65 0 675 1316
use contact_23  contact_23_65
timestamp 1624494425
transform 1 0 40341 0 1 617
box 0 0 66 66
use contact_24  contact_24_65
timestamp 1624494425
transform 1 0 40345 0 1 617
box 0 0 58 66
use contact_25  contact_25_131
timestamp 1624494425
transform 1 0 40124 0 1 216
box 0 0 64 64
use contact_25  contact_25_133
timestamp 1624494425
transform 1 0 39936 0 1 216
box 0 0 64 64
use contact_25  contact_25_321
timestamp 1624494425
transform 1 0 40342 0 1 618
box 0 0 64 64
use contact_26  contact_26_131
timestamp 1624494425
transform 1 0 40123 0 1 211
box 0 0 66 74
use contact_26  contact_26_133
timestamp 1624494425
transform 1 0 39935 0 1 211
box 0 0 66 74
use contact_26  contact_26_321
timestamp 1624494425
transform 1 0 40341 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_65
timestamp 1624494425
transform 1 0 40062 0 1 868
box 65 0 675 1316
use contact_23  contact_23_64
timestamp 1624494425
transform 1 0 40965 0 1 741
box 0 0 66 66
use contact_24  contact_24_64
timestamp 1624494425
transform 1 0 40969 0 1 741
box 0 0 58 66
use contact_25  contact_25_128
timestamp 1624494425
transform 1 0 40720 0 1 92
box 0 0 64 64
use contact_25  contact_25_130
timestamp 1624494425
transform 1 0 40588 0 1 92
box 0 0 64 64
use contact_25  contact_25_320
timestamp 1624494425
transform 1 0 40966 0 1 742
box 0 0 64 64
use contact_26  contact_26_128
timestamp 1624494425
transform 1 0 40719 0 1 87
box 0 0 66 74
use contact_26  contact_26_130
timestamp 1624494425
transform 1 0 40587 0 1 87
box 0 0 66 74
use contact_26  contact_26_320
timestamp 1624494425
transform 1 0 40965 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_64
timestamp 1624494425
transform -1 0 41310 0 1 868
box 65 0 675 1316
use contact_23  contact_23_63
timestamp 1624494425
transform 1 0 41589 0 1 369
box 0 0 66 66
use contact_24  contact_24_63
timestamp 1624494425
transform 1 0 41593 0 1 369
box 0 0 58 66
use contact_25  contact_25_127
timestamp 1624494425
transform 1 0 41372 0 1 216
box 0 0 64 64
use contact_25  contact_25_129
timestamp 1624494425
transform 1 0 41184 0 1 216
box 0 0 64 64
use contact_25  contact_25_319
timestamp 1624494425
transform 1 0 41590 0 1 370
box 0 0 64 64
use contact_26  contact_26_127
timestamp 1624494425
transform 1 0 41371 0 1 211
box 0 0 66 74
use contact_26  contact_26_129
timestamp 1624494425
transform 1 0 41183 0 1 211
box 0 0 66 74
use contact_26  contact_26_319
timestamp 1624494425
transform 1 0 41589 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_63
timestamp 1624494425
transform 1 0 41310 0 1 868
box 65 0 675 1316
use contact_23  contact_23_62
timestamp 1624494425
transform 1 0 42213 0 1 493
box 0 0 66 66
use contact_24  contact_24_62
timestamp 1624494425
transform 1 0 42217 0 1 493
box 0 0 58 66
use contact_25  contact_25_124
timestamp 1624494425
transform 1 0 41968 0 1 92
box 0 0 64 64
use contact_25  contact_25_126
timestamp 1624494425
transform 1 0 41836 0 1 92
box 0 0 64 64
use contact_25  contact_25_318
timestamp 1624494425
transform 1 0 42214 0 1 494
box 0 0 64 64
use contact_26  contact_26_124
timestamp 1624494425
transform 1 0 41967 0 1 87
box 0 0 66 74
use contact_26  contact_26_126
timestamp 1624494425
transform 1 0 41835 0 1 87
box 0 0 66 74
use contact_26  contact_26_318
timestamp 1624494425
transform 1 0 42213 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_62
timestamp 1624494425
transform -1 0 42558 0 1 868
box 65 0 675 1316
use contact_23  contact_23_61
timestamp 1624494425
transform 1 0 42837 0 1 617
box 0 0 66 66
use contact_24  contact_24_61
timestamp 1624494425
transform 1 0 42841 0 1 617
box 0 0 58 66
use contact_25  contact_25_123
timestamp 1624494425
transform 1 0 42620 0 1 216
box 0 0 64 64
use contact_25  contact_25_125
timestamp 1624494425
transform 1 0 42432 0 1 216
box 0 0 64 64
use contact_25  contact_25_317
timestamp 1624494425
transform 1 0 42838 0 1 618
box 0 0 64 64
use contact_26  contact_26_123
timestamp 1624494425
transform 1 0 42619 0 1 211
box 0 0 66 74
use contact_26  contact_26_125
timestamp 1624494425
transform 1 0 42431 0 1 211
box 0 0 66 74
use contact_26  contact_26_317
timestamp 1624494425
transform 1 0 42837 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_61
timestamp 1624494425
transform 1 0 42558 0 1 868
box 65 0 675 1316
use contact_23  contact_23_60
timestamp 1624494425
transform 1 0 43461 0 1 741
box 0 0 66 66
use contact_24  contact_24_60
timestamp 1624494425
transform 1 0 43465 0 1 741
box 0 0 58 66
use contact_25  contact_25_120
timestamp 1624494425
transform 1 0 43216 0 1 92
box 0 0 64 64
use contact_25  contact_25_122
timestamp 1624494425
transform 1 0 43084 0 1 92
box 0 0 64 64
use contact_25  contact_25_316
timestamp 1624494425
transform 1 0 43462 0 1 742
box 0 0 64 64
use contact_26  contact_26_120
timestamp 1624494425
transform 1 0 43215 0 1 87
box 0 0 66 74
use contact_26  contact_26_122
timestamp 1624494425
transform 1 0 43083 0 1 87
box 0 0 66 74
use contact_26  contact_26_316
timestamp 1624494425
transform 1 0 43461 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_60
timestamp 1624494425
transform -1 0 43806 0 1 868
box 65 0 675 1316
use contact_23  contact_23_59
timestamp 1624494425
transform 1 0 44085 0 1 369
box 0 0 66 66
use contact_24  contact_24_59
timestamp 1624494425
transform 1 0 44089 0 1 369
box 0 0 58 66
use contact_25  contact_25_119
timestamp 1624494425
transform 1 0 43868 0 1 216
box 0 0 64 64
use contact_25  contact_25_121
timestamp 1624494425
transform 1 0 43680 0 1 216
box 0 0 64 64
use contact_25  contact_25_315
timestamp 1624494425
transform 1 0 44086 0 1 370
box 0 0 64 64
use contact_26  contact_26_119
timestamp 1624494425
transform 1 0 43867 0 1 211
box 0 0 66 74
use contact_26  contact_26_121
timestamp 1624494425
transform 1 0 43679 0 1 211
box 0 0 66 74
use contact_26  contact_26_315
timestamp 1624494425
transform 1 0 44085 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_59
timestamp 1624494425
transform 1 0 43806 0 1 868
box 65 0 675 1316
use contact_23  contact_23_58
timestamp 1624494425
transform 1 0 44709 0 1 493
box 0 0 66 66
use contact_24  contact_24_58
timestamp 1624494425
transform 1 0 44713 0 1 493
box 0 0 58 66
use contact_25  contact_25_116
timestamp 1624494425
transform 1 0 44464 0 1 92
box 0 0 64 64
use contact_25  contact_25_118
timestamp 1624494425
transform 1 0 44332 0 1 92
box 0 0 64 64
use contact_25  contact_25_314
timestamp 1624494425
transform 1 0 44710 0 1 494
box 0 0 64 64
use contact_26  contact_26_116
timestamp 1624494425
transform 1 0 44463 0 1 87
box 0 0 66 74
use contact_26  contact_26_118
timestamp 1624494425
transform 1 0 44331 0 1 87
box 0 0 66 74
use contact_26  contact_26_314
timestamp 1624494425
transform 1 0 44709 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_58
timestamp 1624494425
transform -1 0 45054 0 1 868
box 65 0 675 1316
use contact_23  contact_23_57
timestamp 1624494425
transform 1 0 45333 0 1 617
box 0 0 66 66
use contact_24  contact_24_57
timestamp 1624494425
transform 1 0 45337 0 1 617
box 0 0 58 66
use contact_25  contact_25_115
timestamp 1624494425
transform 1 0 45116 0 1 216
box 0 0 64 64
use contact_25  contact_25_117
timestamp 1624494425
transform 1 0 44928 0 1 216
box 0 0 64 64
use contact_25  contact_25_313
timestamp 1624494425
transform 1 0 45334 0 1 618
box 0 0 64 64
use contact_26  contact_26_115
timestamp 1624494425
transform 1 0 45115 0 1 211
box 0 0 66 74
use contact_26  contact_26_117
timestamp 1624494425
transform 1 0 44927 0 1 211
box 0 0 66 74
use contact_26  contact_26_313
timestamp 1624494425
transform 1 0 45333 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_57
timestamp 1624494425
transform 1 0 45054 0 1 868
box 65 0 675 1316
use contact_23  contact_23_56
timestamp 1624494425
transform 1 0 45957 0 1 741
box 0 0 66 66
use contact_24  contact_24_56
timestamp 1624494425
transform 1 0 45961 0 1 741
box 0 0 58 66
use contact_25  contact_25_112
timestamp 1624494425
transform 1 0 45712 0 1 92
box 0 0 64 64
use contact_25  contact_25_114
timestamp 1624494425
transform 1 0 45580 0 1 92
box 0 0 64 64
use contact_25  contact_25_312
timestamp 1624494425
transform 1 0 45958 0 1 742
box 0 0 64 64
use contact_26  contact_26_112
timestamp 1624494425
transform 1 0 45711 0 1 87
box 0 0 66 74
use contact_26  contact_26_114
timestamp 1624494425
transform 1 0 45579 0 1 87
box 0 0 66 74
use contact_26  contact_26_312
timestamp 1624494425
transform 1 0 45957 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_56
timestamp 1624494425
transform -1 0 46302 0 1 868
box 65 0 675 1316
use contact_23  contact_23_55
timestamp 1624494425
transform 1 0 46581 0 1 369
box 0 0 66 66
use contact_24  contact_24_55
timestamp 1624494425
transform 1 0 46585 0 1 369
box 0 0 58 66
use contact_25  contact_25_111
timestamp 1624494425
transform 1 0 46364 0 1 216
box 0 0 64 64
use contact_25  contact_25_113
timestamp 1624494425
transform 1 0 46176 0 1 216
box 0 0 64 64
use contact_25  contact_25_311
timestamp 1624494425
transform 1 0 46582 0 1 370
box 0 0 64 64
use contact_26  contact_26_111
timestamp 1624494425
transform 1 0 46363 0 1 211
box 0 0 66 74
use contact_26  contact_26_113
timestamp 1624494425
transform 1 0 46175 0 1 211
box 0 0 66 74
use contact_26  contact_26_311
timestamp 1624494425
transform 1 0 46581 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_55
timestamp 1624494425
transform 1 0 46302 0 1 868
box 65 0 675 1316
use contact_23  contact_23_54
timestamp 1624494425
transform 1 0 47205 0 1 493
box 0 0 66 66
use contact_24  contact_24_54
timestamp 1624494425
transform 1 0 47209 0 1 493
box 0 0 58 66
use contact_25  contact_25_108
timestamp 1624494425
transform 1 0 46960 0 1 92
box 0 0 64 64
use contact_25  contact_25_110
timestamp 1624494425
transform 1 0 46828 0 1 92
box 0 0 64 64
use contact_25  contact_25_310
timestamp 1624494425
transform 1 0 47206 0 1 494
box 0 0 64 64
use contact_26  contact_26_108
timestamp 1624494425
transform 1 0 46959 0 1 87
box 0 0 66 74
use contact_26  contact_26_110
timestamp 1624494425
transform 1 0 46827 0 1 87
box 0 0 66 74
use contact_26  contact_26_310
timestamp 1624494425
transform 1 0 47205 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_54
timestamp 1624494425
transform -1 0 47550 0 1 868
box 65 0 675 1316
use contact_23  contact_23_53
timestamp 1624494425
transform 1 0 47829 0 1 617
box 0 0 66 66
use contact_24  contact_24_53
timestamp 1624494425
transform 1 0 47833 0 1 617
box 0 0 58 66
use contact_25  contact_25_107
timestamp 1624494425
transform 1 0 47612 0 1 216
box 0 0 64 64
use contact_25  contact_25_109
timestamp 1624494425
transform 1 0 47424 0 1 216
box 0 0 64 64
use contact_25  contact_25_309
timestamp 1624494425
transform 1 0 47830 0 1 618
box 0 0 64 64
use contact_26  contact_26_107
timestamp 1624494425
transform 1 0 47611 0 1 211
box 0 0 66 74
use contact_26  contact_26_109
timestamp 1624494425
transform 1 0 47423 0 1 211
box 0 0 66 74
use contact_26  contact_26_309
timestamp 1624494425
transform 1 0 47829 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_53
timestamp 1624494425
transform 1 0 47550 0 1 868
box 65 0 675 1316
use contact_23  contact_23_52
timestamp 1624494425
transform 1 0 48453 0 1 741
box 0 0 66 66
use contact_24  contact_24_52
timestamp 1624494425
transform 1 0 48457 0 1 741
box 0 0 58 66
use contact_25  contact_25_104
timestamp 1624494425
transform 1 0 48208 0 1 92
box 0 0 64 64
use contact_25  contact_25_106
timestamp 1624494425
transform 1 0 48076 0 1 92
box 0 0 64 64
use contact_25  contact_25_308
timestamp 1624494425
transform 1 0 48454 0 1 742
box 0 0 64 64
use contact_26  contact_26_104
timestamp 1624494425
transform 1 0 48207 0 1 87
box 0 0 66 74
use contact_26  contact_26_106
timestamp 1624494425
transform 1 0 48075 0 1 87
box 0 0 66 74
use contact_26  contact_26_308
timestamp 1624494425
transform 1 0 48453 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_52
timestamp 1624494425
transform -1 0 48798 0 1 868
box 65 0 675 1316
use contact_23  contact_23_51
timestamp 1624494425
transform 1 0 49077 0 1 369
box 0 0 66 66
use contact_24  contact_24_51
timestamp 1624494425
transform 1 0 49081 0 1 369
box 0 0 58 66
use contact_25  contact_25_103
timestamp 1624494425
transform 1 0 48860 0 1 216
box 0 0 64 64
use contact_25  contact_25_105
timestamp 1624494425
transform 1 0 48672 0 1 216
box 0 0 64 64
use contact_25  contact_25_307
timestamp 1624494425
transform 1 0 49078 0 1 370
box 0 0 64 64
use contact_26  contact_26_103
timestamp 1624494425
transform 1 0 48859 0 1 211
box 0 0 66 74
use contact_26  contact_26_105
timestamp 1624494425
transform 1 0 48671 0 1 211
box 0 0 66 74
use contact_26  contact_26_307
timestamp 1624494425
transform 1 0 49077 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_51
timestamp 1624494425
transform 1 0 48798 0 1 868
box 65 0 675 1316
use contact_23  contact_23_50
timestamp 1624494425
transform 1 0 49701 0 1 493
box 0 0 66 66
use contact_25  contact_25_100
timestamp 1624494425
transform 1 0 49456 0 1 92
box 0 0 64 64
use contact_25  contact_25_102
timestamp 1624494425
transform 1 0 49324 0 1 92
box 0 0 64 64
use contact_25  contact_25_306
timestamp 1624494425
transform 1 0 49702 0 1 494
box 0 0 64 64
use contact_26  contact_26_100
timestamp 1624494425
transform 1 0 49455 0 1 87
box 0 0 66 74
use contact_26  contact_26_102
timestamp 1624494425
transform 1 0 49323 0 1 87
box 0 0 66 74
use contact_26  contact_26_306
timestamp 1624494425
transform 1 0 49701 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_50
timestamp 1624494425
transform -1 0 50046 0 1 868
box 65 0 675 1316
use contact_24  contact_24_50
timestamp 1624494425
transform 1 0 49705 0 1 493
box 0 0 58 66
use contact_25  contact_25_99
timestamp 1624494425
transform 1 0 50108 0 1 216
box 0 0 64 64
use contact_25  contact_25_101
timestamp 1624494425
transform 1 0 49920 0 1 216
box 0 0 64 64
use contact_26  contact_26_99
timestamp 1624494425
transform 1 0 50107 0 1 211
box 0 0 66 74
use contact_26  contact_26_101
timestamp 1624494425
transform 1 0 49919 0 1 211
box 0 0 66 74
use column_mux_0  column_mux_0_49
timestamp 1624494425
transform 1 0 50046 0 1 868
box 65 0 675 1316
use contact_23  contact_23_49
timestamp 1624494425
transform 1 0 50325 0 1 617
box 0 0 66 66
use contact_24  contact_24_49
timestamp 1624494425
transform 1 0 50329 0 1 617
box 0 0 58 66
use contact_25  contact_25_96
timestamp 1624494425
transform 1 0 50704 0 1 92
box 0 0 64 64
use contact_25  contact_25_98
timestamp 1624494425
transform 1 0 50572 0 1 92
box 0 0 64 64
use contact_25  contact_25_305
timestamp 1624494425
transform 1 0 50326 0 1 618
box 0 0 64 64
use contact_26  contact_26_96
timestamp 1624494425
transform 1 0 50703 0 1 87
box 0 0 66 74
use contact_26  contact_26_98
timestamp 1624494425
transform 1 0 50571 0 1 87
box 0 0 66 74
use contact_26  contact_26_305
timestamp 1624494425
transform 1 0 50325 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_48
timestamp 1624494425
transform -1 0 51294 0 1 868
box 65 0 675 1316
use contact_23  contact_23_48
timestamp 1624494425
transform 1 0 50949 0 1 741
box 0 0 66 66
use contact_24  contact_24_48
timestamp 1624494425
transform 1 0 50953 0 1 741
box 0 0 58 66
use contact_25  contact_25_95
timestamp 1624494425
transform 1 0 51356 0 1 216
box 0 0 64 64
use contact_25  contact_25_97
timestamp 1624494425
transform 1 0 51168 0 1 216
box 0 0 64 64
use contact_25  contact_25_304
timestamp 1624494425
transform 1 0 50950 0 1 742
box 0 0 64 64
use contact_26  contact_26_95
timestamp 1624494425
transform 1 0 51355 0 1 211
box 0 0 66 74
use contact_26  contact_26_97
timestamp 1624494425
transform 1 0 51167 0 1 211
box 0 0 66 74
use contact_26  contact_26_304
timestamp 1624494425
transform 1 0 50949 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_47
timestamp 1624494425
transform 1 0 51294 0 1 868
box 65 0 675 1316
use contact_23  contact_23_47
timestamp 1624494425
transform 1 0 51573 0 1 369
box 0 0 66 66
use contact_24  contact_24_47
timestamp 1624494425
transform 1 0 51577 0 1 369
box 0 0 58 66
use contact_25  contact_25_92
timestamp 1624494425
transform 1 0 51952 0 1 92
box 0 0 64 64
use contact_25  contact_25_94
timestamp 1624494425
transform 1 0 51820 0 1 92
box 0 0 64 64
use contact_25  contact_25_303
timestamp 1624494425
transform 1 0 51574 0 1 370
box 0 0 64 64
use contact_26  contact_26_92
timestamp 1624494425
transform 1 0 51951 0 1 87
box 0 0 66 74
use contact_26  contact_26_94
timestamp 1624494425
transform 1 0 51819 0 1 87
box 0 0 66 74
use contact_26  contact_26_303
timestamp 1624494425
transform 1 0 51573 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_46
timestamp 1624494425
transform -1 0 52542 0 1 868
box 65 0 675 1316
use contact_23  contact_23_46
timestamp 1624494425
transform 1 0 52197 0 1 493
box 0 0 66 66
use contact_24  contact_24_46
timestamp 1624494425
transform 1 0 52201 0 1 493
box 0 0 58 66
use contact_25  contact_25_91
timestamp 1624494425
transform 1 0 52604 0 1 216
box 0 0 64 64
use contact_25  contact_25_93
timestamp 1624494425
transform 1 0 52416 0 1 216
box 0 0 64 64
use contact_25  contact_25_302
timestamp 1624494425
transform 1 0 52198 0 1 494
box 0 0 64 64
use contact_26  contact_26_91
timestamp 1624494425
transform 1 0 52603 0 1 211
box 0 0 66 74
use contact_26  contact_26_93
timestamp 1624494425
transform 1 0 52415 0 1 211
box 0 0 66 74
use contact_26  contact_26_302
timestamp 1624494425
transform 1 0 52197 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_45
timestamp 1624494425
transform 1 0 52542 0 1 868
box 65 0 675 1316
use contact_23  contact_23_45
timestamp 1624494425
transform 1 0 52821 0 1 617
box 0 0 66 66
use contact_24  contact_24_45
timestamp 1624494425
transform 1 0 52825 0 1 617
box 0 0 58 66
use contact_25  contact_25_88
timestamp 1624494425
transform 1 0 53200 0 1 92
box 0 0 64 64
use contact_25  contact_25_90
timestamp 1624494425
transform 1 0 53068 0 1 92
box 0 0 64 64
use contact_25  contact_25_301
timestamp 1624494425
transform 1 0 52822 0 1 618
box 0 0 64 64
use contact_26  contact_26_88
timestamp 1624494425
transform 1 0 53199 0 1 87
box 0 0 66 74
use contact_26  contact_26_90
timestamp 1624494425
transform 1 0 53067 0 1 87
box 0 0 66 74
use contact_26  contact_26_301
timestamp 1624494425
transform 1 0 52821 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_44
timestamp 1624494425
transform -1 0 53790 0 1 868
box 65 0 675 1316
use contact_23  contact_23_44
timestamp 1624494425
transform 1 0 53445 0 1 741
box 0 0 66 66
use contact_24  contact_24_44
timestamp 1624494425
transform 1 0 53449 0 1 741
box 0 0 58 66
use contact_25  contact_25_87
timestamp 1624494425
transform 1 0 53852 0 1 216
box 0 0 64 64
use contact_25  contact_25_89
timestamp 1624494425
transform 1 0 53664 0 1 216
box 0 0 64 64
use contact_25  contact_25_300
timestamp 1624494425
transform 1 0 53446 0 1 742
box 0 0 64 64
use contact_26  contact_26_87
timestamp 1624494425
transform 1 0 53851 0 1 211
box 0 0 66 74
use contact_26  contact_26_89
timestamp 1624494425
transform 1 0 53663 0 1 211
box 0 0 66 74
use contact_26  contact_26_300
timestamp 1624494425
transform 1 0 53445 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_43
timestamp 1624494425
transform 1 0 53790 0 1 868
box 65 0 675 1316
use contact_23  contact_23_43
timestamp 1624494425
transform 1 0 54069 0 1 369
box 0 0 66 66
use contact_24  contact_24_43
timestamp 1624494425
transform 1 0 54073 0 1 369
box 0 0 58 66
use contact_25  contact_25_84
timestamp 1624494425
transform 1 0 54448 0 1 92
box 0 0 64 64
use contact_25  contact_25_86
timestamp 1624494425
transform 1 0 54316 0 1 92
box 0 0 64 64
use contact_25  contact_25_299
timestamp 1624494425
transform 1 0 54070 0 1 370
box 0 0 64 64
use contact_26  contact_26_84
timestamp 1624494425
transform 1 0 54447 0 1 87
box 0 0 66 74
use contact_26  contact_26_86
timestamp 1624494425
transform 1 0 54315 0 1 87
box 0 0 66 74
use contact_26  contact_26_299
timestamp 1624494425
transform 1 0 54069 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_42
timestamp 1624494425
transform -1 0 55038 0 1 868
box 65 0 675 1316
use contact_23  contact_23_42
timestamp 1624494425
transform 1 0 54693 0 1 493
box 0 0 66 66
use contact_24  contact_24_42
timestamp 1624494425
transform 1 0 54697 0 1 493
box 0 0 58 66
use contact_25  contact_25_83
timestamp 1624494425
transform 1 0 55100 0 1 216
box 0 0 64 64
use contact_25  contact_25_85
timestamp 1624494425
transform 1 0 54912 0 1 216
box 0 0 64 64
use contact_25  contact_25_298
timestamp 1624494425
transform 1 0 54694 0 1 494
box 0 0 64 64
use contact_26  contact_26_83
timestamp 1624494425
transform 1 0 55099 0 1 211
box 0 0 66 74
use contact_26  contact_26_85
timestamp 1624494425
transform 1 0 54911 0 1 211
box 0 0 66 74
use contact_26  contact_26_298
timestamp 1624494425
transform 1 0 54693 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_41
timestamp 1624494425
transform 1 0 55038 0 1 868
box 65 0 675 1316
use contact_23  contact_23_41
timestamp 1624494425
transform 1 0 55317 0 1 617
box 0 0 66 66
use contact_24  contact_24_41
timestamp 1624494425
transform 1 0 55321 0 1 617
box 0 0 58 66
use contact_25  contact_25_80
timestamp 1624494425
transform 1 0 55696 0 1 92
box 0 0 64 64
use contact_25  contact_25_82
timestamp 1624494425
transform 1 0 55564 0 1 92
box 0 0 64 64
use contact_25  contact_25_297
timestamp 1624494425
transform 1 0 55318 0 1 618
box 0 0 64 64
use contact_26  contact_26_80
timestamp 1624494425
transform 1 0 55695 0 1 87
box 0 0 66 74
use contact_26  contact_26_82
timestamp 1624494425
transform 1 0 55563 0 1 87
box 0 0 66 74
use contact_26  contact_26_297
timestamp 1624494425
transform 1 0 55317 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_40
timestamp 1624494425
transform -1 0 56286 0 1 868
box 65 0 675 1316
use contact_23  contact_23_40
timestamp 1624494425
transform 1 0 55941 0 1 741
box 0 0 66 66
use contact_24  contact_24_40
timestamp 1624494425
transform 1 0 55945 0 1 741
box 0 0 58 66
use contact_25  contact_25_79
timestamp 1624494425
transform 1 0 56348 0 1 216
box 0 0 64 64
use contact_25  contact_25_81
timestamp 1624494425
transform 1 0 56160 0 1 216
box 0 0 64 64
use contact_25  contact_25_296
timestamp 1624494425
transform 1 0 55942 0 1 742
box 0 0 64 64
use contact_26  contact_26_79
timestamp 1624494425
transform 1 0 56347 0 1 211
box 0 0 66 74
use contact_26  contact_26_81
timestamp 1624494425
transform 1 0 56159 0 1 211
box 0 0 66 74
use contact_26  contact_26_296
timestamp 1624494425
transform 1 0 55941 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_39
timestamp 1624494425
transform 1 0 56286 0 1 868
box 65 0 675 1316
use contact_23  contact_23_39
timestamp 1624494425
transform 1 0 56565 0 1 369
box 0 0 66 66
use contact_24  contact_24_39
timestamp 1624494425
transform 1 0 56569 0 1 369
box 0 0 58 66
use contact_25  contact_25_76
timestamp 1624494425
transform 1 0 56944 0 1 92
box 0 0 64 64
use contact_25  contact_25_78
timestamp 1624494425
transform 1 0 56812 0 1 92
box 0 0 64 64
use contact_25  contact_25_295
timestamp 1624494425
transform 1 0 56566 0 1 370
box 0 0 64 64
use contact_26  contact_26_76
timestamp 1624494425
transform 1 0 56943 0 1 87
box 0 0 66 74
use contact_26  contact_26_78
timestamp 1624494425
transform 1 0 56811 0 1 87
box 0 0 66 74
use contact_26  contact_26_295
timestamp 1624494425
transform 1 0 56565 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_38
timestamp 1624494425
transform -1 0 57534 0 1 868
box 65 0 675 1316
use contact_23  contact_23_38
timestamp 1624494425
transform 1 0 57189 0 1 493
box 0 0 66 66
use contact_24  contact_24_38
timestamp 1624494425
transform 1 0 57193 0 1 493
box 0 0 58 66
use contact_25  contact_25_75
timestamp 1624494425
transform 1 0 57596 0 1 216
box 0 0 64 64
use contact_25  contact_25_77
timestamp 1624494425
transform 1 0 57408 0 1 216
box 0 0 64 64
use contact_25  contact_25_294
timestamp 1624494425
transform 1 0 57190 0 1 494
box 0 0 64 64
use contact_26  contact_26_75
timestamp 1624494425
transform 1 0 57595 0 1 211
box 0 0 66 74
use contact_26  contact_26_77
timestamp 1624494425
transform 1 0 57407 0 1 211
box 0 0 66 74
use contact_26  contact_26_294
timestamp 1624494425
transform 1 0 57189 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_37
timestamp 1624494425
transform 1 0 57534 0 1 868
box 65 0 675 1316
use contact_23  contact_23_37
timestamp 1624494425
transform 1 0 57813 0 1 617
box 0 0 66 66
use contact_24  contact_24_37
timestamp 1624494425
transform 1 0 57817 0 1 617
box 0 0 58 66
use contact_25  contact_25_72
timestamp 1624494425
transform 1 0 58192 0 1 92
box 0 0 64 64
use contact_25  contact_25_74
timestamp 1624494425
transform 1 0 58060 0 1 92
box 0 0 64 64
use contact_25  contact_25_293
timestamp 1624494425
transform 1 0 57814 0 1 618
box 0 0 64 64
use contact_26  contact_26_72
timestamp 1624494425
transform 1 0 58191 0 1 87
box 0 0 66 74
use contact_26  contact_26_74
timestamp 1624494425
transform 1 0 58059 0 1 87
box 0 0 66 74
use contact_26  contact_26_293
timestamp 1624494425
transform 1 0 57813 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_36
timestamp 1624494425
transform -1 0 58782 0 1 868
box 65 0 675 1316
use contact_23  contact_23_36
timestamp 1624494425
transform 1 0 58437 0 1 741
box 0 0 66 66
use contact_24  contact_24_36
timestamp 1624494425
transform 1 0 58441 0 1 741
box 0 0 58 66
use contact_25  contact_25_71
timestamp 1624494425
transform 1 0 58844 0 1 216
box 0 0 64 64
use contact_25  contact_25_73
timestamp 1624494425
transform 1 0 58656 0 1 216
box 0 0 64 64
use contact_25  contact_25_292
timestamp 1624494425
transform 1 0 58438 0 1 742
box 0 0 64 64
use contact_26  contact_26_71
timestamp 1624494425
transform 1 0 58843 0 1 211
box 0 0 66 74
use contact_26  contact_26_73
timestamp 1624494425
transform 1 0 58655 0 1 211
box 0 0 66 74
use contact_26  contact_26_292
timestamp 1624494425
transform 1 0 58437 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_35
timestamp 1624494425
transform 1 0 58782 0 1 868
box 65 0 675 1316
use contact_23  contact_23_35
timestamp 1624494425
transform 1 0 59061 0 1 369
box 0 0 66 66
use contact_24  contact_24_35
timestamp 1624494425
transform 1 0 59065 0 1 369
box 0 0 58 66
use contact_25  contact_25_68
timestamp 1624494425
transform 1 0 59440 0 1 92
box 0 0 64 64
use contact_25  contact_25_70
timestamp 1624494425
transform 1 0 59308 0 1 92
box 0 0 64 64
use contact_25  contact_25_291
timestamp 1624494425
transform 1 0 59062 0 1 370
box 0 0 64 64
use contact_26  contact_26_68
timestamp 1624494425
transform 1 0 59439 0 1 87
box 0 0 66 74
use contact_26  contact_26_70
timestamp 1624494425
transform 1 0 59307 0 1 87
box 0 0 66 74
use contact_26  contact_26_291
timestamp 1624494425
transform 1 0 59061 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_34
timestamp 1624494425
transform -1 0 60030 0 1 868
box 65 0 675 1316
use contact_23  contact_23_34
timestamp 1624494425
transform 1 0 59685 0 1 493
box 0 0 66 66
use contact_24  contact_24_34
timestamp 1624494425
transform 1 0 59689 0 1 493
box 0 0 58 66
use contact_25  contact_25_69
timestamp 1624494425
transform 1 0 59904 0 1 216
box 0 0 64 64
use contact_25  contact_25_290
timestamp 1624494425
transform 1 0 59686 0 1 494
box 0 0 64 64
use contact_26  contact_26_69
timestamp 1624494425
transform 1 0 59903 0 1 211
box 0 0 66 74
use contact_26  contact_26_290
timestamp 1624494425
transform 1 0 59685 0 1 489
box 0 0 66 74
use contact_25  contact_25_67
timestamp 1624494425
transform 1 0 60092 0 1 216
box 0 0 64 64
use contact_26  contact_26_67
timestamp 1624494425
transform 1 0 60091 0 1 211
box 0 0 66 74
use contact_25  contact_25_66
timestamp 1624494425
transform 1 0 60556 0 1 92
box 0 0 64 64
use contact_26  contact_26_66
timestamp 1624494425
transform 1 0 60555 0 1 87
box 0 0 66 74
use contact_25  contact_25_64
timestamp 1624494425
transform 1 0 60688 0 1 92
box 0 0 64 64
use contact_26  contact_26_64
timestamp 1624494425
transform 1 0 60687 0 1 87
box 0 0 66 74
use contact_23  contact_23_33
timestamp 1624494425
transform 1 0 60309 0 1 617
box 0 0 66 66
use contact_24  contact_24_33
timestamp 1624494425
transform 1 0 60313 0 1 617
box 0 0 58 66
use contact_25  contact_25_289
timestamp 1624494425
transform 1 0 60310 0 1 618
box 0 0 64 64
use contact_26  contact_26_289
timestamp 1624494425
transform 1 0 60309 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_33
timestamp 1624494425
transform 1 0 60030 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_32
timestamp 1624494425
transform -1 0 61278 0 1 868
box 65 0 675 1316
use contact_23  contact_23_32
timestamp 1624494425
transform 1 0 60933 0 1 741
box 0 0 66 66
use contact_24  contact_24_32
timestamp 1624494425
transform 1 0 60937 0 1 741
box 0 0 58 66
use contact_25  contact_25_65
timestamp 1624494425
transform 1 0 61152 0 1 216
box 0 0 64 64
use contact_25  contact_25_288
timestamp 1624494425
transform 1 0 60934 0 1 742
box 0 0 64 64
use contact_26  contact_26_65
timestamp 1624494425
transform 1 0 61151 0 1 211
box 0 0 66 74
use contact_26  contact_26_288
timestamp 1624494425
transform 1 0 60933 0 1 737
box 0 0 66 74
use contact_26  contact_26_287
timestamp 1624494425
transform 1 0 61557 0 1 365
box 0 0 66 74
use contact_26  contact_26_63
timestamp 1624494425
transform 1 0 61339 0 1 211
box 0 0 66 74
use contact_26  contact_26_62
timestamp 1624494425
transform 1 0 61803 0 1 87
box 0 0 66 74
use contact_25  contact_25_287
timestamp 1624494425
transform 1 0 61558 0 1 370
box 0 0 64 64
use contact_25  contact_25_63
timestamp 1624494425
transform 1 0 61340 0 1 216
box 0 0 64 64
use contact_25  contact_25_62
timestamp 1624494425
transform 1 0 61804 0 1 92
box 0 0 64 64
use contact_24  contact_24_31
timestamp 1624494425
transform 1 0 61561 0 1 369
box 0 0 58 66
use contact_23  contact_23_31
timestamp 1624494425
transform 1 0 61557 0 1 369
box 0 0 66 66
use column_mux_0  column_mux_0_31
timestamp 1624494425
transform 1 0 61278 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_30
timestamp 1624494425
transform -1 0 62526 0 1 868
box 65 0 675 1316
use contact_23  contact_23_30
timestamp 1624494425
transform 1 0 62181 0 1 493
box 0 0 66 66
use contact_24  contact_24_30
timestamp 1624494425
transform 1 0 62185 0 1 493
box 0 0 58 66
use contact_25  contact_25_60
timestamp 1624494425
transform 1 0 61936 0 1 92
box 0 0 64 64
use contact_25  contact_25_61
timestamp 1624494425
transform 1 0 62400 0 1 216
box 0 0 64 64
use contact_25  contact_25_286
timestamp 1624494425
transform 1 0 62182 0 1 494
box 0 0 64 64
use contact_26  contact_26_60
timestamp 1624494425
transform 1 0 61935 0 1 87
box 0 0 66 74
use contact_26  contact_26_61
timestamp 1624494425
transform 1 0 62399 0 1 211
box 0 0 66 74
use contact_26  contact_26_286
timestamp 1624494425
transform 1 0 62181 0 1 489
box 0 0 66 74
use contact_26  contact_26_285
timestamp 1624494425
transform 1 0 62805 0 1 613
box 0 0 66 74
use contact_26  contact_26_59
timestamp 1624494425
transform 1 0 62587 0 1 211
box 0 0 66 74
use contact_26  contact_26_58
timestamp 1624494425
transform 1 0 63051 0 1 87
box 0 0 66 74
use contact_25  contact_25_285
timestamp 1624494425
transform 1 0 62806 0 1 618
box 0 0 64 64
use contact_25  contact_25_59
timestamp 1624494425
transform 1 0 62588 0 1 216
box 0 0 64 64
use contact_25  contact_25_58
timestamp 1624494425
transform 1 0 63052 0 1 92
box 0 0 64 64
use contact_24  contact_24_29
timestamp 1624494425
transform 1 0 62809 0 1 617
box 0 0 58 66
use contact_23  contact_23_29
timestamp 1624494425
transform 1 0 62805 0 1 617
box 0 0 66 66
use column_mux_0  column_mux_0_29
timestamp 1624494425
transform 1 0 62526 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_28
timestamp 1624494425
transform -1 0 63774 0 1 868
box 65 0 675 1316
use contact_23  contact_23_28
timestamp 1624494425
transform 1 0 63429 0 1 741
box 0 0 66 66
use contact_24  contact_24_28
timestamp 1624494425
transform 1 0 63433 0 1 741
box 0 0 58 66
use contact_25  contact_25_56
timestamp 1624494425
transform 1 0 63184 0 1 92
box 0 0 64 64
use contact_25  contact_25_57
timestamp 1624494425
transform 1 0 63648 0 1 216
box 0 0 64 64
use contact_25  contact_25_284
timestamp 1624494425
transform 1 0 63430 0 1 742
box 0 0 64 64
use contact_26  contact_26_56
timestamp 1624494425
transform 1 0 63183 0 1 87
box 0 0 66 74
use contact_26  contact_26_57
timestamp 1624494425
transform 1 0 63647 0 1 211
box 0 0 66 74
use contact_26  contact_26_284
timestamp 1624494425
transform 1 0 63429 0 1 737
box 0 0 66 74
use contact_26  contact_26_283
timestamp 1624494425
transform 1 0 64053 0 1 365
box 0 0 66 74
use contact_26  contact_26_55
timestamp 1624494425
transform 1 0 63835 0 1 211
box 0 0 66 74
use contact_26  contact_26_54
timestamp 1624494425
transform 1 0 64299 0 1 87
box 0 0 66 74
use contact_25  contact_25_283
timestamp 1624494425
transform 1 0 64054 0 1 370
box 0 0 64 64
use contact_25  contact_25_55
timestamp 1624494425
transform 1 0 63836 0 1 216
box 0 0 64 64
use contact_25  contact_25_54
timestamp 1624494425
transform 1 0 64300 0 1 92
box 0 0 64 64
use contact_24  contact_24_27
timestamp 1624494425
transform 1 0 64057 0 1 369
box 0 0 58 66
use contact_23  contact_23_27
timestamp 1624494425
transform 1 0 64053 0 1 369
box 0 0 66 66
use column_mux_0  column_mux_0_27
timestamp 1624494425
transform 1 0 63774 0 1 868
box 65 0 675 1316
use column_mux_0  column_mux_0_26
timestamp 1624494425
transform -1 0 65022 0 1 868
box 65 0 675 1316
use contact_23  contact_23_26
timestamp 1624494425
transform 1 0 64677 0 1 493
box 0 0 66 66
use contact_24  contact_24_26
timestamp 1624494425
transform 1 0 64681 0 1 493
box 0 0 58 66
use contact_25  contact_25_52
timestamp 1624494425
transform 1 0 64432 0 1 92
box 0 0 64 64
use contact_25  contact_25_53
timestamp 1624494425
transform 1 0 64896 0 1 216
box 0 0 64 64
use contact_25  contact_25_282
timestamp 1624494425
transform 1 0 64678 0 1 494
box 0 0 64 64
use contact_26  contact_26_52
timestamp 1624494425
transform 1 0 64431 0 1 87
box 0 0 66 74
use contact_26  contact_26_53
timestamp 1624494425
transform 1 0 64895 0 1 211
box 0 0 66 74
use contact_26  contact_26_282
timestamp 1624494425
transform 1 0 64677 0 1 489
box 0 0 66 74
use contact_23  contact_23_25
timestamp 1624494425
transform 1 0 65301 0 1 617
box 0 0 66 66
use contact_24  contact_24_25
timestamp 1624494425
transform 1 0 65305 0 1 617
box 0 0 58 66
use contact_25  contact_25_50
timestamp 1624494425
transform 1 0 65548 0 1 92
box 0 0 64 64
use contact_25  contact_25_51
timestamp 1624494425
transform 1 0 65084 0 1 216
box 0 0 64 64
use contact_25  contact_25_281
timestamp 1624494425
transform 1 0 65302 0 1 618
box 0 0 64 64
use contact_26  contact_26_50
timestamp 1624494425
transform 1 0 65547 0 1 87
box 0 0 66 74
use contact_26  contact_26_51
timestamp 1624494425
transform 1 0 65083 0 1 211
box 0 0 66 74
use contact_26  contact_26_281
timestamp 1624494425
transform 1 0 65301 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_25
timestamp 1624494425
transform 1 0 65022 0 1 868
box 65 0 675 1316
use contact_23  contact_23_24
timestamp 1624494425
transform 1 0 65925 0 1 741
box 0 0 66 66
use contact_24  contact_24_24
timestamp 1624494425
transform 1 0 65929 0 1 741
box 0 0 58 66
use contact_25  contact_25_48
timestamp 1624494425
transform 1 0 65680 0 1 92
box 0 0 64 64
use contact_25  contact_25_49
timestamp 1624494425
transform 1 0 66144 0 1 216
box 0 0 64 64
use contact_25  contact_25_280
timestamp 1624494425
transform 1 0 65926 0 1 742
box 0 0 64 64
use contact_26  contact_26_48
timestamp 1624494425
transform 1 0 65679 0 1 87
box 0 0 66 74
use contact_26  contact_26_49
timestamp 1624494425
transform 1 0 66143 0 1 211
box 0 0 66 74
use contact_26  contact_26_280
timestamp 1624494425
transform 1 0 65925 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_24
timestamp 1624494425
transform -1 0 66270 0 1 868
box 65 0 675 1316
use contact_23  contact_23_23
timestamp 1624494425
transform 1 0 66549 0 1 369
box 0 0 66 66
use contact_24  contact_24_23
timestamp 1624494425
transform 1 0 66553 0 1 369
box 0 0 58 66
use contact_25  contact_25_46
timestamp 1624494425
transform 1 0 66796 0 1 92
box 0 0 64 64
use contact_25  contact_25_47
timestamp 1624494425
transform 1 0 66332 0 1 216
box 0 0 64 64
use contact_25  contact_25_279
timestamp 1624494425
transform 1 0 66550 0 1 370
box 0 0 64 64
use contact_26  contact_26_46
timestamp 1624494425
transform 1 0 66795 0 1 87
box 0 0 66 74
use contact_26  contact_26_47
timestamp 1624494425
transform 1 0 66331 0 1 211
box 0 0 66 74
use contact_26  contact_26_279
timestamp 1624494425
transform 1 0 66549 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_23
timestamp 1624494425
transform 1 0 66270 0 1 868
box 65 0 675 1316
use contact_23  contact_23_22
timestamp 1624494425
transform 1 0 67173 0 1 493
box 0 0 66 66
use contact_24  contact_24_22
timestamp 1624494425
transform 1 0 67177 0 1 493
box 0 0 58 66
use contact_25  contact_25_44
timestamp 1624494425
transform 1 0 66928 0 1 92
box 0 0 64 64
use contact_25  contact_25_45
timestamp 1624494425
transform 1 0 67392 0 1 216
box 0 0 64 64
use contact_25  contact_25_278
timestamp 1624494425
transform 1 0 67174 0 1 494
box 0 0 64 64
use contact_26  contact_26_44
timestamp 1624494425
transform 1 0 66927 0 1 87
box 0 0 66 74
use contact_26  contact_26_45
timestamp 1624494425
transform 1 0 67391 0 1 211
box 0 0 66 74
use contact_26  contact_26_278
timestamp 1624494425
transform 1 0 67173 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_22
timestamp 1624494425
transform -1 0 67518 0 1 868
box 65 0 675 1316
use contact_23  contact_23_21
timestamp 1624494425
transform 1 0 67797 0 1 617
box 0 0 66 66
use contact_24  contact_24_21
timestamp 1624494425
transform 1 0 67801 0 1 617
box 0 0 58 66
use contact_25  contact_25_43
timestamp 1624494425
transform 1 0 67580 0 1 216
box 0 0 64 64
use contact_25  contact_25_277
timestamp 1624494425
transform 1 0 67798 0 1 618
box 0 0 64 64
use contact_26  contact_26_43
timestamp 1624494425
transform 1 0 67579 0 1 211
box 0 0 66 74
use contact_26  contact_26_277
timestamp 1624494425
transform 1 0 67797 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_21
timestamp 1624494425
transform 1 0 67518 0 1 868
box 65 0 675 1316
use contact_25  contact_25_40
timestamp 1624494425
transform 1 0 68176 0 1 92
box 0 0 64 64
use contact_25  contact_25_42
timestamp 1624494425
transform 1 0 68044 0 1 92
box 0 0 64 64
use contact_26  contact_26_40
timestamp 1624494425
transform 1 0 68175 0 1 87
box 0 0 66 74
use contact_26  contact_26_42
timestamp 1624494425
transform 1 0 68043 0 1 87
box 0 0 66 74
use contact_25  contact_25_41
timestamp 1624494425
transform 1 0 68640 0 1 216
box 0 0 64 64
use contact_26  contact_26_41
timestamp 1624494425
transform 1 0 68639 0 1 211
box 0 0 66 74
use contact_23  contact_23_20
timestamp 1624494425
transform 1 0 68421 0 1 741
box 0 0 66 66
use contact_24  contact_24_20
timestamp 1624494425
transform 1 0 68425 0 1 741
box 0 0 58 66
use contact_25  contact_25_276
timestamp 1624494425
transform 1 0 68422 0 1 742
box 0 0 64 64
use contact_26  contact_26_276
timestamp 1624494425
transform 1 0 68421 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_20
timestamp 1624494425
transform -1 0 68766 0 1 868
box 65 0 675 1316
use contact_23  contact_23_19
timestamp 1624494425
transform 1 0 69045 0 1 369
box 0 0 66 66
use contact_24  contact_24_19
timestamp 1624494425
transform 1 0 69049 0 1 369
box 0 0 58 66
use contact_25  contact_25_39
timestamp 1624494425
transform 1 0 68828 0 1 216
box 0 0 64 64
use contact_25  contact_25_275
timestamp 1624494425
transform 1 0 69046 0 1 370
box 0 0 64 64
use contact_26  contact_26_39
timestamp 1624494425
transform 1 0 68827 0 1 211
box 0 0 66 74
use contact_26  contact_26_275
timestamp 1624494425
transform 1 0 69045 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_19
timestamp 1624494425
transform 1 0 68766 0 1 868
box 65 0 675 1316
use contact_23  contact_23_18
timestamp 1624494425
transform 1 0 69669 0 1 493
box 0 0 66 66
use contact_24  contact_24_18
timestamp 1624494425
transform 1 0 69673 0 1 493
box 0 0 58 66
use contact_25  contact_25_36
timestamp 1624494425
transform 1 0 69424 0 1 92
box 0 0 64 64
use contact_25  contact_25_38
timestamp 1624494425
transform 1 0 69292 0 1 92
box 0 0 64 64
use contact_25  contact_25_274
timestamp 1624494425
transform 1 0 69670 0 1 494
box 0 0 64 64
use contact_26  contact_26_36
timestamp 1624494425
transform 1 0 69423 0 1 87
box 0 0 66 74
use contact_26  contact_26_38
timestamp 1624494425
transform 1 0 69291 0 1 87
box 0 0 66 74
use contact_26  contact_26_274
timestamp 1624494425
transform 1 0 69669 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_18
timestamp 1624494425
transform -1 0 70014 0 1 868
box 65 0 675 1316
use contact_23  contact_23_17
timestamp 1624494425
transform 1 0 70293 0 1 617
box 0 0 66 66
use contact_24  contact_24_17
timestamp 1624494425
transform 1 0 70297 0 1 617
box 0 0 58 66
use contact_25  contact_25_35
timestamp 1624494425
transform 1 0 70076 0 1 216
box 0 0 64 64
use contact_25  contact_25_37
timestamp 1624494425
transform 1 0 69888 0 1 216
box 0 0 64 64
use contact_25  contact_25_273
timestamp 1624494425
transform 1 0 70294 0 1 618
box 0 0 64 64
use contact_26  contact_26_35
timestamp 1624494425
transform 1 0 70075 0 1 211
box 0 0 66 74
use contact_26  contact_26_37
timestamp 1624494425
transform 1 0 69887 0 1 211
box 0 0 66 74
use contact_26  contact_26_273
timestamp 1624494425
transform 1 0 70293 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_17
timestamp 1624494425
transform 1 0 70014 0 1 868
box 65 0 675 1316
use contact_23  contact_23_16
timestamp 1624494425
transform 1 0 70917 0 1 741
box 0 0 66 66
use contact_24  contact_24_16
timestamp 1624494425
transform 1 0 70921 0 1 741
box 0 0 58 66
use contact_25  contact_25_32
timestamp 1624494425
transform 1 0 70672 0 1 92
box 0 0 64 64
use contact_25  contact_25_34
timestamp 1624494425
transform 1 0 70540 0 1 92
box 0 0 64 64
use contact_25  contact_25_272
timestamp 1624494425
transform 1 0 70918 0 1 742
box 0 0 64 64
use contact_26  contact_26_32
timestamp 1624494425
transform 1 0 70671 0 1 87
box 0 0 66 74
use contact_26  contact_26_34
timestamp 1624494425
transform 1 0 70539 0 1 87
box 0 0 66 74
use contact_26  contact_26_272
timestamp 1624494425
transform 1 0 70917 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_16
timestamp 1624494425
transform -1 0 71262 0 1 868
box 65 0 675 1316
use contact_23  contact_23_15
timestamp 1624494425
transform 1 0 71541 0 1 369
box 0 0 66 66
use contact_24  contact_24_15
timestamp 1624494425
transform 1 0 71545 0 1 369
box 0 0 58 66
use contact_25  contact_25_31
timestamp 1624494425
transform 1 0 71324 0 1 216
box 0 0 64 64
use contact_25  contact_25_33
timestamp 1624494425
transform 1 0 71136 0 1 216
box 0 0 64 64
use contact_25  contact_25_271
timestamp 1624494425
transform 1 0 71542 0 1 370
box 0 0 64 64
use contact_26  contact_26_31
timestamp 1624494425
transform 1 0 71323 0 1 211
box 0 0 66 74
use contact_26  contact_26_33
timestamp 1624494425
transform 1 0 71135 0 1 211
box 0 0 66 74
use contact_26  contact_26_271
timestamp 1624494425
transform 1 0 71541 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_15
timestamp 1624494425
transform 1 0 71262 0 1 868
box 65 0 675 1316
use contact_23  contact_23_14
timestamp 1624494425
transform 1 0 72165 0 1 493
box 0 0 66 66
use contact_24  contact_24_14
timestamp 1624494425
transform 1 0 72169 0 1 493
box 0 0 58 66
use contact_25  contact_25_28
timestamp 1624494425
transform 1 0 71920 0 1 92
box 0 0 64 64
use contact_25  contact_25_30
timestamp 1624494425
transform 1 0 71788 0 1 92
box 0 0 64 64
use contact_25  contact_25_270
timestamp 1624494425
transform 1 0 72166 0 1 494
box 0 0 64 64
use contact_26  contact_26_28
timestamp 1624494425
transform 1 0 71919 0 1 87
box 0 0 66 74
use contact_26  contact_26_30
timestamp 1624494425
transform 1 0 71787 0 1 87
box 0 0 66 74
use contact_26  contact_26_270
timestamp 1624494425
transform 1 0 72165 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_14
timestamp 1624494425
transform -1 0 72510 0 1 868
box 65 0 675 1316
use contact_23  contact_23_13
timestamp 1624494425
transform 1 0 72789 0 1 617
box 0 0 66 66
use contact_24  contact_24_13
timestamp 1624494425
transform 1 0 72793 0 1 617
box 0 0 58 66
use contact_25  contact_25_27
timestamp 1624494425
transform 1 0 72572 0 1 216
box 0 0 64 64
use contact_25  contact_25_29
timestamp 1624494425
transform 1 0 72384 0 1 216
box 0 0 64 64
use contact_25  contact_25_269
timestamp 1624494425
transform 1 0 72790 0 1 618
box 0 0 64 64
use contact_26  contact_26_27
timestamp 1624494425
transform 1 0 72571 0 1 211
box 0 0 66 74
use contact_26  contact_26_29
timestamp 1624494425
transform 1 0 72383 0 1 211
box 0 0 66 74
use contact_26  contact_26_269
timestamp 1624494425
transform 1 0 72789 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_13
timestamp 1624494425
transform 1 0 72510 0 1 868
box 65 0 675 1316
use contact_23  contact_23_12
timestamp 1624494425
transform 1 0 73413 0 1 741
box 0 0 66 66
use contact_24  contact_24_12
timestamp 1624494425
transform 1 0 73417 0 1 741
box 0 0 58 66
use contact_25  contact_25_24
timestamp 1624494425
transform 1 0 73168 0 1 92
box 0 0 64 64
use contact_25  contact_25_26
timestamp 1624494425
transform 1 0 73036 0 1 92
box 0 0 64 64
use contact_25  contact_25_268
timestamp 1624494425
transform 1 0 73414 0 1 742
box 0 0 64 64
use contact_26  contact_26_24
timestamp 1624494425
transform 1 0 73167 0 1 87
box 0 0 66 74
use contact_26  contact_26_26
timestamp 1624494425
transform 1 0 73035 0 1 87
box 0 0 66 74
use contact_26  contact_26_268
timestamp 1624494425
transform 1 0 73413 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_12
timestamp 1624494425
transform -1 0 73758 0 1 868
box 65 0 675 1316
use contact_23  contact_23_11
timestamp 1624494425
transform 1 0 74037 0 1 369
box 0 0 66 66
use contact_24  contact_24_11
timestamp 1624494425
transform 1 0 74041 0 1 369
box 0 0 58 66
use contact_25  contact_25_23
timestamp 1624494425
transform 1 0 73820 0 1 216
box 0 0 64 64
use contact_25  contact_25_25
timestamp 1624494425
transform 1 0 73632 0 1 216
box 0 0 64 64
use contact_25  contact_25_267
timestamp 1624494425
transform 1 0 74038 0 1 370
box 0 0 64 64
use contact_26  contact_26_23
timestamp 1624494425
transform 1 0 73819 0 1 211
box 0 0 66 74
use contact_26  contact_26_25
timestamp 1624494425
transform 1 0 73631 0 1 211
box 0 0 66 74
use contact_26  contact_26_267
timestamp 1624494425
transform 1 0 74037 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_11
timestamp 1624494425
transform 1 0 73758 0 1 868
box 65 0 675 1316
use contact_23  contact_23_10
timestamp 1624494425
transform 1 0 74661 0 1 493
box 0 0 66 66
use contact_24  contact_24_10
timestamp 1624494425
transform 1 0 74665 0 1 493
box 0 0 58 66
use contact_25  contact_25_20
timestamp 1624494425
transform 1 0 74416 0 1 92
box 0 0 64 64
use contact_25  contact_25_22
timestamp 1624494425
transform 1 0 74284 0 1 92
box 0 0 64 64
use contact_25  contact_25_266
timestamp 1624494425
transform 1 0 74662 0 1 494
box 0 0 64 64
use contact_26  contact_26_20
timestamp 1624494425
transform 1 0 74415 0 1 87
box 0 0 66 74
use contact_26  contact_26_22
timestamp 1624494425
transform 1 0 74283 0 1 87
box 0 0 66 74
use contact_26  contact_26_266
timestamp 1624494425
transform 1 0 74661 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_10
timestamp 1624494425
transform -1 0 75006 0 1 868
box 65 0 675 1316
use contact_23  contact_23_9
timestamp 1624494425
transform 1 0 75285 0 1 617
box 0 0 66 66
use contact_24  contact_24_9
timestamp 1624494425
transform 1 0 75289 0 1 617
box 0 0 58 66
use contact_25  contact_25_19
timestamp 1624494425
transform 1 0 75068 0 1 216
box 0 0 64 64
use contact_25  contact_25_21
timestamp 1624494425
transform 1 0 74880 0 1 216
box 0 0 64 64
use contact_25  contact_25_265
timestamp 1624494425
transform 1 0 75286 0 1 618
box 0 0 64 64
use contact_26  contact_26_19
timestamp 1624494425
transform 1 0 75067 0 1 211
box 0 0 66 74
use contact_26  contact_26_21
timestamp 1624494425
transform 1 0 74879 0 1 211
box 0 0 66 74
use contact_26  contact_26_265
timestamp 1624494425
transform 1 0 75285 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_9
timestamp 1624494425
transform 1 0 75006 0 1 868
box 65 0 675 1316
use contact_23  contact_23_8
timestamp 1624494425
transform 1 0 75909 0 1 741
box 0 0 66 66
use contact_24  contact_24_8
timestamp 1624494425
transform 1 0 75913 0 1 741
box 0 0 58 66
use contact_25  contact_25_16
timestamp 1624494425
transform 1 0 75664 0 1 92
box 0 0 64 64
use contact_25  contact_25_18
timestamp 1624494425
transform 1 0 75532 0 1 92
box 0 0 64 64
use contact_25  contact_25_264
timestamp 1624494425
transform 1 0 75910 0 1 742
box 0 0 64 64
use contact_26  contact_26_16
timestamp 1624494425
transform 1 0 75663 0 1 87
box 0 0 66 74
use contact_26  contact_26_18
timestamp 1624494425
transform 1 0 75531 0 1 87
box 0 0 66 74
use contact_26  contact_26_264
timestamp 1624494425
transform 1 0 75909 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_8
timestamp 1624494425
transform -1 0 76254 0 1 868
box 65 0 675 1316
use contact_23  contact_23_7
timestamp 1624494425
transform 1 0 76533 0 1 369
box 0 0 66 66
use contact_24  contact_24_7
timestamp 1624494425
transform 1 0 76537 0 1 369
box 0 0 58 66
use contact_25  contact_25_15
timestamp 1624494425
transform 1 0 76316 0 1 216
box 0 0 64 64
use contact_25  contact_25_17
timestamp 1624494425
transform 1 0 76128 0 1 216
box 0 0 64 64
use contact_25  contact_25_263
timestamp 1624494425
transform 1 0 76534 0 1 370
box 0 0 64 64
use contact_26  contact_26_15
timestamp 1624494425
transform 1 0 76315 0 1 211
box 0 0 66 74
use contact_26  contact_26_17
timestamp 1624494425
transform 1 0 76127 0 1 211
box 0 0 66 74
use contact_26  contact_26_263
timestamp 1624494425
transform 1 0 76533 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_7
timestamp 1624494425
transform 1 0 76254 0 1 868
box 65 0 675 1316
use contact_23  contact_23_6
timestamp 1624494425
transform 1 0 77157 0 1 493
box 0 0 66 66
use contact_24  contact_24_6
timestamp 1624494425
transform 1 0 77161 0 1 493
box 0 0 58 66
use contact_25  contact_25_12
timestamp 1624494425
transform 1 0 76912 0 1 92
box 0 0 64 64
use contact_25  contact_25_14
timestamp 1624494425
transform 1 0 76780 0 1 92
box 0 0 64 64
use contact_25  contact_25_262
timestamp 1624494425
transform 1 0 77158 0 1 494
box 0 0 64 64
use contact_26  contact_26_12
timestamp 1624494425
transform 1 0 76911 0 1 87
box 0 0 66 74
use contact_26  contact_26_14
timestamp 1624494425
transform 1 0 76779 0 1 87
box 0 0 66 74
use contact_26  contact_26_262
timestamp 1624494425
transform 1 0 77157 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_6
timestamp 1624494425
transform -1 0 77502 0 1 868
box 65 0 675 1316
use contact_23  contact_23_5
timestamp 1624494425
transform 1 0 77781 0 1 617
box 0 0 66 66
use contact_24  contact_24_5
timestamp 1624494425
transform 1 0 77785 0 1 617
box 0 0 58 66
use contact_25  contact_25_11
timestamp 1624494425
transform 1 0 77564 0 1 216
box 0 0 64 64
use contact_25  contact_25_13
timestamp 1624494425
transform 1 0 77376 0 1 216
box 0 0 64 64
use contact_25  contact_25_261
timestamp 1624494425
transform 1 0 77782 0 1 618
box 0 0 64 64
use contact_26  contact_26_11
timestamp 1624494425
transform 1 0 77563 0 1 211
box 0 0 66 74
use contact_26  contact_26_13
timestamp 1624494425
transform 1 0 77375 0 1 211
box 0 0 66 74
use contact_26  contact_26_261
timestamp 1624494425
transform 1 0 77781 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_5
timestamp 1624494425
transform 1 0 77502 0 1 868
box 65 0 675 1316
use contact_23  contact_23_4
timestamp 1624494425
transform 1 0 78405 0 1 741
box 0 0 66 66
use contact_24  contact_24_4
timestamp 1624494425
transform 1 0 78409 0 1 741
box 0 0 58 66
use contact_25  contact_25_8
timestamp 1624494425
transform 1 0 78160 0 1 92
box 0 0 64 64
use contact_25  contact_25_10
timestamp 1624494425
transform 1 0 78028 0 1 92
box 0 0 64 64
use contact_25  contact_25_260
timestamp 1624494425
transform 1 0 78406 0 1 742
box 0 0 64 64
use contact_26  contact_26_8
timestamp 1624494425
transform 1 0 78159 0 1 87
box 0 0 66 74
use contact_26  contact_26_10
timestamp 1624494425
transform 1 0 78027 0 1 87
box 0 0 66 74
use contact_26  contact_26_260
timestamp 1624494425
transform 1 0 78405 0 1 737
box 0 0 66 74
use column_mux_0  column_mux_0_4
timestamp 1624494425
transform -1 0 78750 0 1 868
box 65 0 675 1316
use contact_23  contact_23_3
timestamp 1624494425
transform 1 0 79029 0 1 369
box 0 0 66 66
use contact_25  contact_25_7
timestamp 1624494425
transform 1 0 78812 0 1 216
box 0 0 64 64
use contact_25  contact_25_9
timestamp 1624494425
transform 1 0 78624 0 1 216
box 0 0 64 64
use contact_25  contact_25_259
timestamp 1624494425
transform 1 0 79030 0 1 370
box 0 0 64 64
use contact_26  contact_26_7
timestamp 1624494425
transform 1 0 78811 0 1 211
box 0 0 66 74
use contact_26  contact_26_9
timestamp 1624494425
transform 1 0 78623 0 1 211
box 0 0 66 74
use contact_26  contact_26_259
timestamp 1624494425
transform 1 0 79029 0 1 365
box 0 0 66 74
use column_mux_0  column_mux_0_3
timestamp 1624494425
transform 1 0 78750 0 1 868
box 65 0 675 1316
use contact_24  contact_24_3
timestamp 1624494425
transform 1 0 79033 0 1 369
box 0 0 58 66
use contact_25  contact_25_4
timestamp 1624494425
transform 1 0 79408 0 1 92
box 0 0 64 64
use contact_25  contact_25_6
timestamp 1624494425
transform 1 0 79276 0 1 92
box 0 0 64 64
use contact_26  contact_26_4
timestamp 1624494425
transform 1 0 79407 0 1 87
box 0 0 66 74
use contact_26  contact_26_6
timestamp 1624494425
transform 1 0 79275 0 1 87
box 0 0 66 74
use column_mux_0  column_mux_0_2
timestamp 1624494425
transform -1 0 79998 0 1 868
box 65 0 675 1316
use contact_23  contact_23_2
timestamp 1624494425
transform 1 0 79653 0 1 493
box 0 0 66 66
use contact_24  contact_24_2
timestamp 1624494425
transform 1 0 79657 0 1 493
box 0 0 58 66
use contact_25  contact_25_3
timestamp 1624494425
transform 1 0 80060 0 1 216
box 0 0 64 64
use contact_25  contact_25_5
timestamp 1624494425
transform 1 0 79872 0 1 216
box 0 0 64 64
use contact_25  contact_25_258
timestamp 1624494425
transform 1 0 79654 0 1 494
box 0 0 64 64
use contact_26  contact_26_3
timestamp 1624494425
transform 1 0 80059 0 1 211
box 0 0 66 74
use contact_26  contact_26_5
timestamp 1624494425
transform 1 0 79871 0 1 211
box 0 0 66 74
use contact_26  contact_26_258
timestamp 1624494425
transform 1 0 79653 0 1 489
box 0 0 66 74
use column_mux_0  column_mux_0_1
timestamp 1624494425
transform 1 0 79998 0 1 868
box 65 0 675 1316
use contact_23  contact_23_1
timestamp 1624494425
transform 1 0 80277 0 1 617
box 0 0 66 66
use contact_24  contact_24_1
timestamp 1624494425
transform 1 0 80281 0 1 617
box 0 0 58 66
use contact_25  contact_25_0
timestamp 1624494425
transform 1 0 80656 0 1 92
box 0 0 64 64
use contact_25  contact_25_2
timestamp 1624494425
transform 1 0 80524 0 1 92
box 0 0 64 64
use contact_25  contact_25_257
timestamp 1624494425
transform 1 0 80278 0 1 618
box 0 0 64 64
use contact_26  contact_26_0
timestamp 1624494425
transform 1 0 80655 0 1 87
box 0 0 66 74
use contact_26  contact_26_2
timestamp 1624494425
transform 1 0 80523 0 1 87
box 0 0 66 74
use contact_26  contact_26_257
timestamp 1624494425
transform 1 0 80277 0 1 613
box 0 0 66 74
use column_mux_0  column_mux_0_0
timestamp 1624494425
transform -1 0 81246 0 1 868
box 65 0 675 1316
use contact_23  contact_23_0
timestamp 1624494425
transform 1 0 80901 0 1 741
box 0 0 66 66
use contact_24  contact_24_0
timestamp 1624494425
transform 1 0 80905 0 1 741
box 0 0 58 66
use contact_25  contact_25_1
timestamp 1624494425
transform 1 0 81120 0 1 216
box 0 0 64 64
use contact_25  contact_25_256
timestamp 1624494425
transform 1 0 80902 0 1 742
box 0 0 64 64
use contact_26  contact_26_1
timestamp 1624494425
transform 1 0 81119 0 1 211
box 0 0 66 74
use contact_26  contact_26_256
timestamp 1624494425
transform 1 0 80901 0 1 737
box 0 0 66 74
<< labels >>
rlabel metal3 s 0 372 81246 432 4 sel_0
rlabel metal3 s 0 496 81246 556 4 sel_1
rlabel metal3 s 0 620 81246 680 4 sel_2
rlabel metal3 s 0 744 81246 804 4 sel_3
rlabel metal1 s 1454 248 1482 868 4 bl_out_0
rlabel metal1 s 1918 124 1946 868 4 br_out_0
rlabel metal1 s 3950 248 3978 868 4 bl_out_1
rlabel metal1 s 4414 124 4442 868 4 br_out_1
rlabel metal1 s 6446 248 6474 868 4 bl_out_2
rlabel metal1 s 6910 124 6938 868 4 br_out_2
rlabel metal1 s 8942 248 8970 868 4 bl_out_3
rlabel metal1 s 9406 124 9434 868 4 br_out_3
rlabel metal1 s 11438 248 11466 868 4 bl_out_4
rlabel metal1 s 11902 124 11930 868 4 br_out_4
rlabel metal1 s 13934 248 13962 868 4 bl_out_5
rlabel metal1 s 14398 124 14426 868 4 br_out_5
rlabel metal1 s 16430 248 16458 868 4 bl_out_6
rlabel metal1 s 16894 124 16922 868 4 br_out_6
rlabel metal1 s 18926 248 18954 868 4 bl_out_7
rlabel metal1 s 19390 124 19418 868 4 br_out_7
rlabel metal1 s 21422 248 21450 868 4 bl_out_8
rlabel metal1 s 21886 124 21914 868 4 br_out_8
rlabel metal1 s 23918 248 23946 868 4 bl_out_9
rlabel metal1 s 24382 124 24410 868 4 br_out_9
rlabel metal1 s 26414 248 26442 868 4 bl_out_10
rlabel metal1 s 26878 124 26906 868 4 br_out_10
rlabel metal1 s 28910 248 28938 868 4 bl_out_11
rlabel metal1 s 29374 124 29402 868 4 br_out_11
rlabel metal1 s 31406 248 31434 868 4 bl_out_12
rlabel metal1 s 31870 124 31898 868 4 br_out_12
rlabel metal1 s 33902 248 33930 868 4 bl_out_13
rlabel metal1 s 34366 124 34394 868 4 br_out_13
rlabel metal1 s 36398 248 36426 868 4 bl_out_14
rlabel metal1 s 36862 124 36890 868 4 br_out_14
rlabel metal1 s 38894 248 38922 868 4 bl_out_15
rlabel metal1 s 39358 124 39386 868 4 br_out_15
rlabel metal1 s 41390 248 41418 868 4 bl_out_16
rlabel metal1 s 41854 124 41882 868 4 br_out_16
rlabel metal1 s 43886 248 43914 868 4 bl_out_17
rlabel metal1 s 44350 124 44378 868 4 br_out_17
rlabel metal1 s 46382 248 46410 868 4 bl_out_18
rlabel metal1 s 46846 124 46874 868 4 br_out_18
rlabel metal1 s 48878 248 48906 868 4 bl_out_19
rlabel metal1 s 49342 124 49370 868 4 br_out_19
rlabel metal1 s 51374 248 51402 868 4 bl_out_20
rlabel metal1 s 51838 124 51866 868 4 br_out_20
rlabel metal1 s 53870 248 53898 868 4 bl_out_21
rlabel metal1 s 54334 124 54362 868 4 br_out_21
rlabel metal1 s 56366 248 56394 868 4 bl_out_22
rlabel metal1 s 56830 124 56858 868 4 br_out_22
rlabel metal1 s 58862 248 58890 868 4 bl_out_23
rlabel metal1 s 59326 124 59354 868 4 br_out_23
rlabel metal1 s 61358 248 61386 868 4 bl_out_24
rlabel metal1 s 61822 124 61850 868 4 br_out_24
rlabel metal1 s 63854 248 63882 868 4 bl_out_25
rlabel metal1 s 64318 124 64346 868 4 br_out_25
rlabel metal1 s 66350 248 66378 868 4 bl_out_26
rlabel metal1 s 66814 124 66842 868 4 br_out_26
rlabel metal1 s 68846 248 68874 868 4 bl_out_27
rlabel metal1 s 69310 124 69338 868 4 br_out_27
rlabel metal1 s 71342 248 71370 868 4 bl_out_28
rlabel metal1 s 71806 124 71834 868 4 br_out_28
rlabel metal1 s 73838 248 73866 868 4 bl_out_29
rlabel metal1 s 74302 124 74330 868 4 br_out_29
rlabel metal1 s 76334 248 76362 868 4 bl_out_30
rlabel metal1 s 76798 124 76826 868 4 br_out_30
rlabel metal1 s 78830 248 78858 868 4 bl_out_31
rlabel metal1 s 79294 124 79322 868 4 br_out_31
rlabel metal1 s 1454 2128 1482 2184 4 bl_0
rlabel metal1 s 1918 2128 1946 2184 4 br_0
rlabel metal1 s 2514 2128 2542 2184 4 bl_1
rlabel metal1 s 2050 2128 2078 2184 4 br_1
rlabel metal1 s 2702 2128 2730 2184 4 bl_2
rlabel metal1 s 3166 2128 3194 2184 4 br_2
rlabel metal1 s 3762 2128 3790 2184 4 bl_3
rlabel metal1 s 3298 2128 3326 2184 4 br_3
rlabel metal1 s 3950 2128 3978 2184 4 bl_4
rlabel metal1 s 4414 2128 4442 2184 4 br_4
rlabel metal1 s 5010 2128 5038 2184 4 bl_5
rlabel metal1 s 4546 2128 4574 2184 4 br_5
rlabel metal1 s 5198 2128 5226 2184 4 bl_6
rlabel metal1 s 5662 2128 5690 2184 4 br_6
rlabel metal1 s 6258 2128 6286 2184 4 bl_7
rlabel metal1 s 5794 2128 5822 2184 4 br_7
rlabel metal1 s 6446 2128 6474 2184 4 bl_8
rlabel metal1 s 6910 2128 6938 2184 4 br_8
rlabel metal1 s 7506 2128 7534 2184 4 bl_9
rlabel metal1 s 7042 2128 7070 2184 4 br_9
rlabel metal1 s 7694 2128 7722 2184 4 bl_10
rlabel metal1 s 8158 2128 8186 2184 4 br_10
rlabel metal1 s 8754 2128 8782 2184 4 bl_11
rlabel metal1 s 8290 2128 8318 2184 4 br_11
rlabel metal1 s 8942 2128 8970 2184 4 bl_12
rlabel metal1 s 9406 2128 9434 2184 4 br_12
rlabel metal1 s 10002 2128 10030 2184 4 bl_13
rlabel metal1 s 9538 2128 9566 2184 4 br_13
rlabel metal1 s 10190 2128 10218 2184 4 bl_14
rlabel metal1 s 10654 2128 10682 2184 4 br_14
rlabel metal1 s 11250 2128 11278 2184 4 bl_15
rlabel metal1 s 10786 2128 10814 2184 4 br_15
rlabel metal1 s 11438 2128 11466 2184 4 bl_16
rlabel metal1 s 11902 2128 11930 2184 4 br_16
rlabel metal1 s 12498 2128 12526 2184 4 bl_17
rlabel metal1 s 12034 2128 12062 2184 4 br_17
rlabel metal1 s 12686 2128 12714 2184 4 bl_18
rlabel metal1 s 13150 2128 13178 2184 4 br_18
rlabel metal1 s 13746 2128 13774 2184 4 bl_19
rlabel metal1 s 13282 2128 13310 2184 4 br_19
rlabel metal1 s 13934 2128 13962 2184 4 bl_20
rlabel metal1 s 14398 2128 14426 2184 4 br_20
rlabel metal1 s 14994 2128 15022 2184 4 bl_21
rlabel metal1 s 14530 2128 14558 2184 4 br_21
rlabel metal1 s 15182 2128 15210 2184 4 bl_22
rlabel metal1 s 15646 2128 15674 2184 4 br_22
rlabel metal1 s 16242 2128 16270 2184 4 bl_23
rlabel metal1 s 15778 2128 15806 2184 4 br_23
rlabel metal1 s 16430 2128 16458 2184 4 bl_24
rlabel metal1 s 16894 2128 16922 2184 4 br_24
rlabel metal1 s 17490 2128 17518 2184 4 bl_25
rlabel metal1 s 17026 2128 17054 2184 4 br_25
rlabel metal1 s 17678 2128 17706 2184 4 bl_26
rlabel metal1 s 18142 2128 18170 2184 4 br_26
rlabel metal1 s 18738 2128 18766 2184 4 bl_27
rlabel metal1 s 18274 2128 18302 2184 4 br_27
rlabel metal1 s 18926 2128 18954 2184 4 bl_28
rlabel metal1 s 19390 2128 19418 2184 4 br_28
rlabel metal1 s 19986 2128 20014 2184 4 bl_29
rlabel metal1 s 19522 2128 19550 2184 4 br_29
rlabel metal1 s 20174 2128 20202 2184 4 bl_30
rlabel metal1 s 20638 2128 20666 2184 4 br_30
rlabel metal1 s 21234 2128 21262 2184 4 bl_31
rlabel metal1 s 20770 2128 20798 2184 4 br_31
rlabel metal1 s 21422 2128 21450 2184 4 bl_32
rlabel metal1 s 21886 2128 21914 2184 4 br_32
rlabel metal1 s 22482 2128 22510 2184 4 bl_33
rlabel metal1 s 22018 2128 22046 2184 4 br_33
rlabel metal1 s 22670 2128 22698 2184 4 bl_34
rlabel metal1 s 23134 2128 23162 2184 4 br_34
rlabel metal1 s 23730 2128 23758 2184 4 bl_35
rlabel metal1 s 23266 2128 23294 2184 4 br_35
rlabel metal1 s 23918 2128 23946 2184 4 bl_36
rlabel metal1 s 24382 2128 24410 2184 4 br_36
rlabel metal1 s 24978 2128 25006 2184 4 bl_37
rlabel metal1 s 24514 2128 24542 2184 4 br_37
rlabel metal1 s 25166 2128 25194 2184 4 bl_38
rlabel metal1 s 25630 2128 25658 2184 4 br_38
rlabel metal1 s 26226 2128 26254 2184 4 bl_39
rlabel metal1 s 25762 2128 25790 2184 4 br_39
rlabel metal1 s 26414 2128 26442 2184 4 bl_40
rlabel metal1 s 26878 2128 26906 2184 4 br_40
rlabel metal1 s 27474 2128 27502 2184 4 bl_41
rlabel metal1 s 27010 2128 27038 2184 4 br_41
rlabel metal1 s 27662 2128 27690 2184 4 bl_42
rlabel metal1 s 28126 2128 28154 2184 4 br_42
rlabel metal1 s 28722 2128 28750 2184 4 bl_43
rlabel metal1 s 28258 2128 28286 2184 4 br_43
rlabel metal1 s 28910 2128 28938 2184 4 bl_44
rlabel metal1 s 29374 2128 29402 2184 4 br_44
rlabel metal1 s 29970 2128 29998 2184 4 bl_45
rlabel metal1 s 29506 2128 29534 2184 4 br_45
rlabel metal1 s 30158 2128 30186 2184 4 bl_46
rlabel metal1 s 30622 2128 30650 2184 4 br_46
rlabel metal1 s 31218 2128 31246 2184 4 bl_47
rlabel metal1 s 30754 2128 30782 2184 4 br_47
rlabel metal1 s 31406 2128 31434 2184 4 bl_48
rlabel metal1 s 31870 2128 31898 2184 4 br_48
rlabel metal1 s 32466 2128 32494 2184 4 bl_49
rlabel metal1 s 32002 2128 32030 2184 4 br_49
rlabel metal1 s 32654 2128 32682 2184 4 bl_50
rlabel metal1 s 33118 2128 33146 2184 4 br_50
rlabel metal1 s 33714 2128 33742 2184 4 bl_51
rlabel metal1 s 33250 2128 33278 2184 4 br_51
rlabel metal1 s 33902 2128 33930 2184 4 bl_52
rlabel metal1 s 34366 2128 34394 2184 4 br_52
rlabel metal1 s 34962 2128 34990 2184 4 bl_53
rlabel metal1 s 34498 2128 34526 2184 4 br_53
rlabel metal1 s 35150 2128 35178 2184 4 bl_54
rlabel metal1 s 35614 2128 35642 2184 4 br_54
rlabel metal1 s 36210 2128 36238 2184 4 bl_55
rlabel metal1 s 35746 2128 35774 2184 4 br_55
rlabel metal1 s 36398 2128 36426 2184 4 bl_56
rlabel metal1 s 36862 2128 36890 2184 4 br_56
rlabel metal1 s 37458 2128 37486 2184 4 bl_57
rlabel metal1 s 36994 2128 37022 2184 4 br_57
rlabel metal1 s 37646 2128 37674 2184 4 bl_58
rlabel metal1 s 38110 2128 38138 2184 4 br_58
rlabel metal1 s 38706 2128 38734 2184 4 bl_59
rlabel metal1 s 38242 2128 38270 2184 4 br_59
rlabel metal1 s 38894 2128 38922 2184 4 bl_60
rlabel metal1 s 39358 2128 39386 2184 4 br_60
rlabel metal1 s 39954 2128 39982 2184 4 bl_61
rlabel metal1 s 39490 2128 39518 2184 4 br_61
rlabel metal1 s 40142 2128 40170 2184 4 bl_62
rlabel metal1 s 40606 2128 40634 2184 4 br_62
rlabel metal1 s 41202 2128 41230 2184 4 bl_63
rlabel metal1 s 40738 2128 40766 2184 4 br_63
rlabel metal1 s 41390 2128 41418 2184 4 bl_64
rlabel metal1 s 41854 2128 41882 2184 4 br_64
rlabel metal1 s 42450 2128 42478 2184 4 bl_65
rlabel metal1 s 41986 2128 42014 2184 4 br_65
rlabel metal1 s 42638 2128 42666 2184 4 bl_66
rlabel metal1 s 43102 2128 43130 2184 4 br_66
rlabel metal1 s 43698 2128 43726 2184 4 bl_67
rlabel metal1 s 43234 2128 43262 2184 4 br_67
rlabel metal1 s 43886 2128 43914 2184 4 bl_68
rlabel metal1 s 44350 2128 44378 2184 4 br_68
rlabel metal1 s 44946 2128 44974 2184 4 bl_69
rlabel metal1 s 44482 2128 44510 2184 4 br_69
rlabel metal1 s 45134 2128 45162 2184 4 bl_70
rlabel metal1 s 45598 2128 45626 2184 4 br_70
rlabel metal1 s 46194 2128 46222 2184 4 bl_71
rlabel metal1 s 45730 2128 45758 2184 4 br_71
rlabel metal1 s 46382 2128 46410 2184 4 bl_72
rlabel metal1 s 46846 2128 46874 2184 4 br_72
rlabel metal1 s 47442 2128 47470 2184 4 bl_73
rlabel metal1 s 46978 2128 47006 2184 4 br_73
rlabel metal1 s 47630 2128 47658 2184 4 bl_74
rlabel metal1 s 48094 2128 48122 2184 4 br_74
rlabel metal1 s 48690 2128 48718 2184 4 bl_75
rlabel metal1 s 48226 2128 48254 2184 4 br_75
rlabel metal1 s 48878 2128 48906 2184 4 bl_76
rlabel metal1 s 49342 2128 49370 2184 4 br_76
rlabel metal1 s 49938 2128 49966 2184 4 bl_77
rlabel metal1 s 49474 2128 49502 2184 4 br_77
rlabel metal1 s 50126 2128 50154 2184 4 bl_78
rlabel metal1 s 50590 2128 50618 2184 4 br_78
rlabel metal1 s 51186 2128 51214 2184 4 bl_79
rlabel metal1 s 50722 2128 50750 2184 4 br_79
rlabel metal1 s 51374 2128 51402 2184 4 bl_80
rlabel metal1 s 51838 2128 51866 2184 4 br_80
rlabel metal1 s 52434 2128 52462 2184 4 bl_81
rlabel metal1 s 51970 2128 51998 2184 4 br_81
rlabel metal1 s 52622 2128 52650 2184 4 bl_82
rlabel metal1 s 53086 2128 53114 2184 4 br_82
rlabel metal1 s 53682 2128 53710 2184 4 bl_83
rlabel metal1 s 53218 2128 53246 2184 4 br_83
rlabel metal1 s 53870 2128 53898 2184 4 bl_84
rlabel metal1 s 54334 2128 54362 2184 4 br_84
rlabel metal1 s 54930 2128 54958 2184 4 bl_85
rlabel metal1 s 54466 2128 54494 2184 4 br_85
rlabel metal1 s 55118 2128 55146 2184 4 bl_86
rlabel metal1 s 55582 2128 55610 2184 4 br_86
rlabel metal1 s 56178 2128 56206 2184 4 bl_87
rlabel metal1 s 55714 2128 55742 2184 4 br_87
rlabel metal1 s 56366 2128 56394 2184 4 bl_88
rlabel metal1 s 56830 2128 56858 2184 4 br_88
rlabel metal1 s 57426 2128 57454 2184 4 bl_89
rlabel metal1 s 56962 2128 56990 2184 4 br_89
rlabel metal1 s 57614 2128 57642 2184 4 bl_90
rlabel metal1 s 58078 2128 58106 2184 4 br_90
rlabel metal1 s 58674 2128 58702 2184 4 bl_91
rlabel metal1 s 58210 2128 58238 2184 4 br_91
rlabel metal1 s 58862 2128 58890 2184 4 bl_92
rlabel metal1 s 59326 2128 59354 2184 4 br_92
rlabel metal1 s 59922 2128 59950 2184 4 bl_93
rlabel metal1 s 59458 2128 59486 2184 4 br_93
rlabel metal1 s 60110 2128 60138 2184 4 bl_94
rlabel metal1 s 60574 2128 60602 2184 4 br_94
rlabel metal1 s 61170 2128 61198 2184 4 bl_95
rlabel metal1 s 60706 2128 60734 2184 4 br_95
rlabel metal1 s 61358 2128 61386 2184 4 bl_96
rlabel metal1 s 61822 2128 61850 2184 4 br_96
rlabel metal1 s 62418 2128 62446 2184 4 bl_97
rlabel metal1 s 61954 2128 61982 2184 4 br_97
rlabel metal1 s 62606 2128 62634 2184 4 bl_98
rlabel metal1 s 63070 2128 63098 2184 4 br_98
rlabel metal1 s 63666 2128 63694 2184 4 bl_99
rlabel metal1 s 63202 2128 63230 2184 4 br_99
rlabel metal1 s 63854 2128 63882 2184 4 bl_100
rlabel metal1 s 64318 2128 64346 2184 4 br_100
rlabel metal1 s 64914 2128 64942 2184 4 bl_101
rlabel metal1 s 64450 2128 64478 2184 4 br_101
rlabel metal1 s 65102 2128 65130 2184 4 bl_102
rlabel metal1 s 65566 2128 65594 2184 4 br_102
rlabel metal1 s 66162 2128 66190 2184 4 bl_103
rlabel metal1 s 65698 2128 65726 2184 4 br_103
rlabel metal1 s 66350 2128 66378 2184 4 bl_104
rlabel metal1 s 66814 2128 66842 2184 4 br_104
rlabel metal1 s 67410 2128 67438 2184 4 bl_105
rlabel metal1 s 66946 2128 66974 2184 4 br_105
rlabel metal1 s 67598 2128 67626 2184 4 bl_106
rlabel metal1 s 68062 2128 68090 2184 4 br_106
rlabel metal1 s 68658 2128 68686 2184 4 bl_107
rlabel metal1 s 68194 2128 68222 2184 4 br_107
rlabel metal1 s 68846 2128 68874 2184 4 bl_108
rlabel metal1 s 69310 2128 69338 2184 4 br_108
rlabel metal1 s 69906 2128 69934 2184 4 bl_109
rlabel metal1 s 69442 2128 69470 2184 4 br_109
rlabel metal1 s 70094 2128 70122 2184 4 bl_110
rlabel metal1 s 70558 2128 70586 2184 4 br_110
rlabel metal1 s 71154 2128 71182 2184 4 bl_111
rlabel metal1 s 70690 2128 70718 2184 4 br_111
rlabel metal1 s 71342 2128 71370 2184 4 bl_112
rlabel metal1 s 71806 2128 71834 2184 4 br_112
rlabel metal1 s 72402 2128 72430 2184 4 bl_113
rlabel metal1 s 71938 2128 71966 2184 4 br_113
rlabel metal1 s 72590 2128 72618 2184 4 bl_114
rlabel metal1 s 73054 2128 73082 2184 4 br_114
rlabel metal1 s 73650 2128 73678 2184 4 bl_115
rlabel metal1 s 73186 2128 73214 2184 4 br_115
rlabel metal1 s 73838 2128 73866 2184 4 bl_116
rlabel metal1 s 74302 2128 74330 2184 4 br_116
rlabel metal1 s 74898 2128 74926 2184 4 bl_117
rlabel metal1 s 74434 2128 74462 2184 4 br_117
rlabel metal1 s 75086 2128 75114 2184 4 bl_118
rlabel metal1 s 75550 2128 75578 2184 4 br_118
rlabel metal1 s 76146 2128 76174 2184 4 bl_119
rlabel metal1 s 75682 2128 75710 2184 4 br_119
rlabel metal1 s 76334 2128 76362 2184 4 bl_120
rlabel metal1 s 76798 2128 76826 2184 4 br_120
rlabel metal1 s 77394 2128 77422 2184 4 bl_121
rlabel metal1 s 76930 2128 76958 2184 4 br_121
rlabel metal1 s 77582 2128 77610 2184 4 bl_122
rlabel metal1 s 78046 2128 78074 2184 4 br_122
rlabel metal1 s 78642 2128 78670 2184 4 bl_123
rlabel metal1 s 78178 2128 78206 2184 4 br_123
rlabel metal1 s 78830 2128 78858 2184 4 bl_124
rlabel metal1 s 79294 2128 79322 2184 4 br_124
rlabel metal1 s 79890 2128 79918 2184 4 bl_125
rlabel metal1 s 79426 2128 79454 2184 4 br_125
rlabel metal1 s 80078 2128 80106 2184 4 bl_126
rlabel metal1 s 80542 2128 80570 2184 4 br_126
rlabel metal1 s 81138 2128 81166 2184 4 bl_127
rlabel metal1 s 80674 2128 80702 2184 4 br_127
rlabel metal3 s 58109 1482 58207 1580 4 gnd
rlabel metal3 s 10685 1482 10783 1580 4 gnd
rlabel metal3 s 10734 1531 10734 1531 4 gnd
rlabel metal3 s 23165 1482 23263 1580 4 gnd
rlabel metal3 s 13181 1482 13279 1580 4 gnd
rlabel metal3 s 31901 1482 31999 1580 4 gnd
rlabel metal3 s 50621 1482 50719 1580 4 gnd
rlabel metal3 s 44381 1482 44479 1580 4 gnd
rlabel metal3 s 61853 1482 61951 1580 4 gnd
rlabel metal3 s 26909 1482 27007 1580 4 gnd
rlabel metal3 s 26958 1531 26958 1531 4 gnd
rlabel metal3 s 20669 1482 20767 1580 4 gnd
rlabel metal3 s 20718 1531 20718 1531 4 gnd
rlabel metal3 s 71837 1482 71935 1580 4 gnd
rlabel metal3 s 80573 1482 80671 1580 4 gnd
rlabel metal3 s 8189 1482 8287 1580 4 gnd
rlabel metal3 s 21917 1482 22015 1580 4 gnd
rlabel metal3 s 5693 1482 5791 1580 4 gnd
rlabel metal3 s 5742 1531 5742 1531 4 gnd
rlabel metal3 s 19421 1482 19519 1580 4 gnd
rlabel metal3 s 73085 1482 73183 1580 4 gnd
rlabel metal3 s 35645 1482 35743 1580 4 gnd
rlabel metal3 s 3197 1482 3295 1580 4 gnd
rlabel metal3 s 3246 1531 3246 1531 4 gnd
rlabel metal3 s 33149 1482 33247 1580 4 gnd
rlabel metal3 s 64349 1482 64447 1580 4 gnd
rlabel metal3 s 24413 1482 24511 1580 4 gnd
rlabel metal3 s 24462 1531 24462 1531 4 gnd
rlabel metal3 s 39389 1482 39487 1580 4 gnd
rlabel metal3 s 15677 1482 15775 1580 4 gnd
rlabel metal3 s 16925 1482 17023 1580 4 gnd
rlabel metal3 s 49373 1482 49471 1580 4 gnd
rlabel metal3 s 38141 1482 38239 1580 4 gnd
rlabel metal3 s 38190 1531 38190 1531 4 gnd
rlabel metal3 s 45629 1482 45727 1580 4 gnd
rlabel metal3 s 45678 1531 45678 1531 4 gnd
rlabel metal3 s 59357 1482 59455 1580 4 gnd
rlabel metal3 s 9437 1482 9535 1580 4 gnd
rlabel metal3 s 6941 1482 7039 1580 4 gnd
rlabel metal3 s 75581 1482 75679 1580 4 gnd
rlabel metal3 s 75630 1531 75630 1531 4 gnd
rlabel metal3 s 40637 1482 40735 1580 4 gnd
rlabel metal3 s 54365 1482 54463 1580 4 gnd
rlabel metal3 s 65597 1482 65695 1580 4 gnd
rlabel metal3 s 43133 1482 43231 1580 4 gnd
rlabel metal3 s 55613 1482 55711 1580 4 gnd
rlabel metal3 s 63101 1482 63199 1580 4 gnd
rlabel metal3 s 30653 1482 30751 1580 4 gnd
rlabel metal3 s 30702 1531 30702 1531 4 gnd
rlabel metal3 s 74333 1482 74431 1580 4 gnd
rlabel metal3 s 70589 1482 70687 1580 4 gnd
rlabel metal3 s 66845 1482 66943 1580 4 gnd
rlabel metal3 s 76829 1482 76927 1580 4 gnd
rlabel metal3 s 68093 1482 68191 1580 4 gnd
rlabel metal3 s 68142 1531 68142 1531 4 gnd
rlabel metal3 s 79325 1482 79423 1580 4 gnd
rlabel metal3 s 29405 1482 29503 1580 4 gnd
rlabel metal3 s 41885 1482 41983 1580 4 gnd
rlabel metal3 s 41934 1531 41934 1531 4 gnd
rlabel metal3 s 60605 1482 60703 1580 4 gnd
rlabel metal3 s 60654 1531 60654 1531 4 gnd
rlabel metal3 s 53117 1482 53215 1580 4 gnd
rlabel metal3 s 48125 1482 48223 1580 4 gnd
rlabel metal3 s 4445 1482 4543 1580 4 gnd
rlabel metal3 s 4494 1531 4494 1531 4 gnd
rlabel metal3 s 1949 1482 2047 1580 4 gnd
rlabel metal3 s 1998 1531 1998 1531 4 gnd
rlabel metal3 s 28157 1482 28255 1580 4 gnd
rlabel metal3 s 18173 1482 18271 1580 4 gnd
rlabel metal3 s 18222 1531 18222 1531 4 gnd
rlabel metal3 s 69341 1482 69439 1580 4 gnd
rlabel metal3 s 36893 1482 36991 1580 4 gnd
rlabel metal3 s 78077 1482 78175 1580 4 gnd
rlabel metal3 s 51869 1482 51967 1580 4 gnd
rlabel metal3 s 51918 1531 51918 1531 4 gnd
rlabel metal3 s 56861 1482 56959 1580 4 gnd
rlabel metal3 s 14429 1482 14527 1580 4 gnd
rlabel metal3 s 14478 1531 14478 1531 4 gnd
rlabel metal3 s 25661 1482 25759 1580 4 gnd
rlabel metal3 s 34397 1482 34495 1580 4 gnd
rlabel metal3 s 34446 1531 34446 1531 4 gnd
rlabel metal3 s 46877 1482 46975 1580 4 gnd
rlabel metal3 s 11933 1482 12031 1580 4 gnd
<< properties >>
string FIXED_BBOX 0 0 79872 2184
<< end >>
